module tt_um_space_invaders_game (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire clknet_0_clk;
 wire abullet_active;
 wire \abullet_x[0] ;
 wire \abullet_x[1] ;
 wire \abullet_x[2] ;
 wire \abullet_x[3] ;
 wire \abullet_x[4] ;
 wire \abullet_x[5] ;
 wire \abullet_x[6] ;
 wire \abullet_x[7] ;
 wire \abullet_x[8] ;
 wire \abullet_x[9] ;
 wire \abullet_y[1] ;
 wire \abullet_y[2] ;
 wire \abullet_y[3] ;
 wire \abullet_y[4] ;
 wire \abullet_y[5] ;
 wire \abullet_y[6] ;
 wire \abullet_y[7] ;
 wire \abullet_y[8] ;
 wire \abullet_y[9] ;
 wire \aliens_alive[0] ;
 wire \aliens_alive[10] ;
 wire \aliens_alive[11] ;
 wire \aliens_alive[12] ;
 wire \aliens_alive[13] ;
 wire \aliens_alive[14] ;
 wire \aliens_alive[15] ;
 wire \aliens_alive[16] ;
 wire \aliens_alive[17] ;
 wire \aliens_alive[18] ;
 wire \aliens_alive[19] ;
 wire \aliens_alive[1] ;
 wire \aliens_alive[20] ;
 wire \aliens_alive[21] ;
 wire \aliens_alive[22] ;
 wire \aliens_alive[23] ;
 wire \aliens_alive[24] ;
 wire \aliens_alive[25] ;
 wire \aliens_alive[26] ;
 wire \aliens_alive[27] ;
 wire \aliens_alive[28] ;
 wire \aliens_alive[29] ;
 wire \aliens_alive[2] ;
 wire \aliens_alive[30] ;
 wire \aliens_alive[31] ;
 wire \aliens_alive[32] ;
 wire \aliens_alive[33] ;
 wire \aliens_alive[34] ;
 wire \aliens_alive[35] ;
 wire \aliens_alive[36] ;
 wire \aliens_alive[37] ;
 wire \aliens_alive[38] ;
 wire \aliens_alive[39] ;
 wire \aliens_alive[3] ;
 wire \aliens_alive[4] ;
 wire \aliens_alive[5] ;
 wire \aliens_alive[6] ;
 wire \aliens_alive[7] ;
 wire \aliens_alive[8] ;
 wire \aliens_alive[9] ;
 wire \barrier1.bar_rom.row_index[0] ;
 wire \barrier1.bar_rom.row_index[1] ;
 wire \barrier1.bar_rom.row_index[2] ;
 wire \barrier1.bar_rom.row_index[3] ;
 wire \barrier1.col_idx[0] ;
 wire \barrier1.col_idx[1] ;
 wire \barrier1.pix_x[2] ;
 wire \barrier1.pix_x[3] ;
 wire \barrier1.pix_x[4] ;
 wire \barrier1.pix_x[5] ;
 wire \barrier1.pix_x[6] ;
 wire \barrier1.pix_x[7] ;
 wire \barrier1.pix_x[8] ;
 wire \barrier1.pix_x[9] ;
 wire \barrier1.pix_y[4] ;
 wire \barrier1.pix_y[5] ;
 wire \barrier1.pix_y[6] ;
 wire \barrier1.pix_y[7] ;
 wire \barrier1.pix_y[8] ;
 wire \barrier1.pix_y[9] ;
 wire \barrier_health[0][0] ;
 wire \barrier_health[0][1] ;
 wire \barrier_health[0][2] ;
 wire \barrier_health[1][0] ;
 wire \barrier_health[1][1] ;
 wire \barrier_health[1][2] ;
 wire \barrier_health[2][0] ;
 wire \barrier_health[2][1] ;
 wire \barrier_health[2][2] ;
 wire \barrier_health[3][0] ;
 wire \barrier_health[3][1] ;
 wire \barrier_health[3][2] ;
 wire \colRand[0] ;
 wire \colRand[1] ;
 wire \colRand[2] ;
 wire \draw_score_inst.digit_health[0] ;
 wire \draw_score_inst.digit_health[1] ;
 wire \draw_score_inst.score[1] ;
 wire \draw_score_inst.score[2] ;
 wire \draw_score_inst.score[3] ;
 wire \draw_score_inst.score[4] ;
 wire \draw_score_inst.score[5] ;
 wire \draw_score_inst.score[6] ;
 wire \draw_score_inst.score[7] ;
 wire \draw_score_inst.score[8] ;
 wire \draw_score_inst.score[9] ;
 wire \draw_score_inst.segment_rom_health.segments[0] ;
 wire \draw_score_inst.segment_rom_health.segments[2] ;
 wire \draw_score_inst.segment_rom_health.segments[4] ;
 wire \draw_score_inst.segment_rom_health.segments[5] ;
 wire \draw_score_inst.segment_rom_health.segments[6] ;
 wire game_over;
 wire game_won;
 wire \group_x[1] ;
 wire \group_x[2] ;
 wire \group_x[3] ;
 wire \group_x[4] ;
 wire \group_x[5] ;
 wire \group_x[6] ;
 wire \group_x[7] ;
 wire \group_x[8] ;
 wire \group_x[9] ;
 wire hsync;
 wire \lA2_x[1] ;
 wire \lfsr[0] ;
 wire \lfsr[1] ;
 wire \lfsr[2] ;
 wire \lfsr[3] ;
 wire \lfsr[4] ;
 wire \lfsr[5] ;
 wire \lfsr[6] ;
 wire \lfsr[7] ;
 wire \lgA2.rx[0] ;
 wire move_dir;
 wire \movement_dir[1] ;
 wire \movement_dir[2] ;
 wire \myShooter.shooter_left_x[1] ;
 wire \myShooter.shooter_left_x[2] ;
 wire \myShooter.shooter_left_x[3] ;
 wire \myShooter.shooter_left_x[4] ;
 wire \myShooter.shooter_left_x[5] ;
 wire \myShooter.shooter_left_x[6] ;
 wire \myShooter.shooter_left_x[7] ;
 wire \myShooter.shooter_left_x[8] ;
 wire \myShooter.shooter_left_x[9] ;
 wire pb_active;
 wire \pb_x[0] ;
 wire \pb_x[1] ;
 wire \pb_x[2] ;
 wire \pb_x[3] ;
 wire \pb_x[4] ;
 wire \pb_x[5] ;
 wire \pb_x[6] ;
 wire \pb_x[7] ;
 wire \pb_x[8] ;
 wire \pb_x[9] ;
 wire \pb_y[0] ;
 wire \pb_y[1] ;
 wire \pb_y[2] ;
 wire \pb_y[3] ;
 wire \pb_y[4] ;
 wire \pb_y[5] ;
 wire \pb_y[6] ;
 wire \pb_y[7] ;
 wire \pb_y[8] ;
 wire \pb_y[9] ;
 wire prev_button0;
 wire prev_button1;
 wire prev_button2;
 wire \prev_vpos[0] ;
 wire \prev_vpos[1] ;
 wire \prev_vpos[2] ;
 wire \prev_vpos[3] ;
 wire \prev_vpos[4] ;
 wire \prev_vpos[5] ;
 wire \prev_vpos[6] ;
 wire \prev_vpos[7] ;
 wire \prev_vpos[8] ;
 wire \prev_vpos[9] ;
 wire \prev_vpos_shooter[0] ;
 wire \prev_vpos_shooter[1] ;
 wire \prev_vpos_shooter[2] ;
 wire \prev_vpos_shooter[3] ;
 wire \prev_vpos_shooter[4] ;
 wire \prev_vpos_shooter[5] ;
 wire \prev_vpos_shooter[6] ;
 wire \prev_vpos_shooter[7] ;
 wire \prev_vpos_shooter[8] ;
 wire \prev_vpos_shooter[9] ;
 wire \selectedRowRand[0] ;
 wire \selectedRowRand[1] ;
 wire \selectedRowRand[2] ;
 wire \sync_gen.vsync ;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;

 sg13g2_inv_2 _3649_ (.Y(_2820_),
    .A(net1232));
 sg13g2_inv_1 _3650_ (.Y(_2821_),
    .A(\group_x[8] ));
 sg13g2_inv_1 _3651_ (.Y(_2822_),
    .A(net1234));
 sg13g2_inv_2 _3652_ (.Y(_2823_),
    .A(net1238));
 sg13g2_inv_2 _3653_ (.Y(_2824_),
    .A(net1240));
 sg13g2_inv_2 _3654_ (.Y(_2825_),
    .A(net1246));
 sg13g2_inv_4 _3655_ (.A(net1249),
    .Y(_2826_));
 sg13g2_inv_4 _3656_ (.A(net1252),
    .Y(_2827_));
 sg13g2_inv_1 _3657_ (.Y(_2828_),
    .A(\abullet_y[8] ));
 sg13g2_inv_1 _3658_ (.Y(_2829_),
    .A(\abullet_y[7] ));
 sg13g2_inv_1 _3659_ (.Y(_2830_),
    .A(net1254));
 sg13g2_inv_1 _3660_ (.Y(_2831_),
    .A(\abullet_y[5] ));
 sg13g2_inv_1 _3661_ (.Y(_2832_),
    .A(\abullet_y[4] ));
 sg13g2_inv_1 _3662_ (.Y(_2833_),
    .A(\abullet_y[3] ));
 sg13g2_inv_1 _3663_ (.Y(_2834_),
    .A(net1255));
 sg13g2_inv_1 _3664_ (.Y(_2835_),
    .A(net355));
 sg13g2_inv_1 _3665_ (.Y(_2836_),
    .A(\myShooter.shooter_left_x[7] ));
 sg13g2_inv_1 _3666_ (.Y(_2837_),
    .A(net1258));
 sg13g2_inv_1 _3667_ (.Y(_2838_),
    .A(\myShooter.shooter_left_x[5] ));
 sg13g2_inv_2 _3668_ (.Y(_2839_),
    .A(\myShooter.shooter_left_x[1] ));
 sg13g2_inv_1 _3669_ (.Y(_2840_),
    .A(net231));
 sg13g2_inv_1 _3670_ (.Y(_2841_),
    .A(net1264));
 sg13g2_inv_4 _3671_ (.A(net1270),
    .Y(_2842_));
 sg13g2_inv_2 _3672_ (.Y(_2843_),
    .A(net1272));
 sg13g2_inv_4 _3673_ (.A(net1275),
    .Y(_2844_));
 sg13g2_inv_4 _3674_ (.A(net1277),
    .Y(_2845_));
 sg13g2_inv_2 _3675_ (.Y(_2846_),
    .A(net1281));
 sg13g2_inv_1 _3676_ (.Y(_2847_),
    .A(net1289));
 sg13g2_inv_1 _3677_ (.Y(_2848_),
    .A(net1294));
 sg13g2_inv_1 _3678_ (.Y(_2849_),
    .A(net1295));
 sg13g2_inv_2 _3679_ (.Y(_2850_),
    .A(net1299));
 sg13g2_inv_1 _3680_ (.Y(_2851_),
    .A(net1301));
 sg13g2_inv_1 _3681_ (.Y(_2852_),
    .A(net268));
 sg13g2_inv_1 _3682_ (.Y(_2853_),
    .A(net290));
 sg13g2_inv_1 _3683_ (.Y(_2854_),
    .A(net257));
 sg13g2_inv_1 _3684_ (.Y(_2855_),
    .A(net273));
 sg13g2_inv_1 _3685_ (.Y(_2856_),
    .A(net279));
 sg13g2_inv_1 _3686_ (.Y(_2857_),
    .A(net261));
 sg13g2_inv_1 _3687_ (.Y(_2858_),
    .A(net233));
 sg13g2_inv_1 _3688_ (.Y(_2859_),
    .A(\abullet_x[8] ));
 sg13g2_inv_1 _3689_ (.Y(_2860_),
    .A(\abullet_x[6] ));
 sg13g2_inv_1 _3690_ (.Y(_2861_),
    .A(\abullet_x[5] ));
 sg13g2_inv_1 _3691_ (.Y(_2862_),
    .A(net1316));
 sg13g2_inv_1 _3692_ (.Y(_2863_),
    .A(\abullet_x[3] ));
 sg13g2_inv_1 _3693_ (.Y(_2864_),
    .A(net1317));
 sg13g2_inv_1 _3694_ (.Y(_2865_),
    .A(\abullet_x[1] ));
 sg13g2_inv_1 _3695_ (.Y(_2866_),
    .A(net375));
 sg13g2_inv_2 _3696_ (.Y(_2867_),
    .A(net1328));
 sg13g2_inv_1 _3697_ (.Y(_2868_),
    .A(net1333));
 sg13g2_inv_1 _3698_ (.Y(_2869_),
    .A(net1338));
 sg13g2_inv_1 _3699_ (.Y(_2870_),
    .A(net1343));
 sg13g2_inv_1 _3700_ (.Y(_2871_),
    .A(net1344));
 sg13g2_inv_1 _3701_ (.Y(_2872_),
    .A(net1346));
 sg13g2_inv_1 _3702_ (.Y(_2873_),
    .A(net1350));
 sg13g2_inv_1 _3703_ (.Y(_2874_),
    .A(net1397));
 sg13g2_inv_4 _3704_ (.A(net1359),
    .Y(_2875_));
 sg13g2_inv_1 _3705_ (.Y(_2876_),
    .A(net1365));
 sg13g2_inv_2 _3706_ (.Y(_2877_),
    .A(net1353));
 sg13g2_inv_1 _3707_ (.Y(_2878_),
    .A(net1417));
 sg13g2_inv_4 _3708_ (.A(net1395),
    .Y(_2879_));
 sg13g2_inv_1 _3709_ (.Y(_2880_),
    .A(net1392));
 sg13g2_inv_1 _3710_ (.Y(_2881_),
    .A(net1384));
 sg13g2_inv_2 _3711_ (.Y(_2882_),
    .A(net1383));
 sg13g2_inv_2 _3712_ (.Y(_2883_),
    .A(net1377));
 sg13g2_inv_1 _3713_ (.Y(_2884_),
    .A(net1371));
 sg13g2_inv_1 _3714_ (.Y(_2885_),
    .A(net413));
 sg13g2_inv_2 _3715_ (.Y(_2886_),
    .A(_0068_));
 sg13g2_inv_1 _3716_ (.Y(_2887_),
    .A(\pb_y[7] ));
 sg13g2_inv_1 _3717_ (.Y(_2888_),
    .A(\pb_y[6] ));
 sg13g2_inv_1 _3718_ (.Y(_2889_),
    .A(net1323));
 sg13g2_inv_1 _3719_ (.Y(_2890_),
    .A(\pb_y[4] ));
 sg13g2_inv_1 _3720_ (.Y(_2891_),
    .A(net1324));
 sg13g2_inv_1 _3721_ (.Y(_2892_),
    .A(net1325));
 sg13g2_inv_1 _3722_ (.Y(_2893_),
    .A(net1326));
 sg13g2_inv_1 _3723_ (.Y(_2894_),
    .A(\pb_y[0] ));
 sg13g2_inv_1 _3724_ (.Y(_2895_),
    .A(_0074_));
 sg13g2_inv_1 _3725_ (.Y(_2896_),
    .A(_0076_));
 sg13g2_inv_1 _3726_ (.Y(_2897_),
    .A(net1229));
 sg13g2_inv_2 _3727_ (.Y(_2898_),
    .A(\draw_score_inst.score[3] ));
 sg13g2_inv_1 _3728_ (.Y(_2899_),
    .A(\draw_score_inst.score[2] ));
 sg13g2_inv_1 _3729_ (.Y(_2900_),
    .A(net1309));
 sg13g2_inv_4 _3730_ (.A(\draw_score_inst.score[4] ),
    .Y(_2901_));
 sg13g2_inv_1 _3731_ (.Y(_2902_),
    .A(net1306));
 sg13g2_inv_1 _3732_ (.Y(_2903_),
    .A(net1305));
 sg13g2_inv_4 _3733_ (.A(_0010_),
    .Y(_2904_));
 sg13g2_inv_2 _3734_ (.Y(_2905_),
    .A(net1282));
 sg13g2_inv_2 _3735_ (.Y(_2906_),
    .A(_0013_));
 sg13g2_inv_4 _3736_ (.A(_0014_),
    .Y(_2907_));
 sg13g2_inv_1 _3737_ (.Y(_2908_),
    .A(_0015_));
 sg13g2_inv_1 _3738_ (.Y(_2909_),
    .A(_0019_));
 sg13g2_inv_1 _3739_ (.Y(_2910_),
    .A(_0020_));
 sg13g2_inv_1 _3740_ (.Y(_2911_),
    .A(_0021_));
 sg13g2_inv_1 _3741_ (.Y(_2912_),
    .A(_0022_));
 sg13g2_inv_1 _3742_ (.Y(_2913_),
    .A(_0023_));
 sg13g2_inv_1 _3743_ (.Y(_2914_),
    .A(_0026_));
 sg13g2_inv_4 _3744_ (.A(net1373),
    .Y(_2915_));
 sg13g2_inv_1 _3745_ (.Y(_2916_),
    .A(_0042_));
 sg13g2_inv_1 _3746_ (.Y(_2917_),
    .A(_0063_));
 sg13g2_nand2b_1 _3747_ (.Y(_2918_),
    .B(net2),
    .A_N(net351));
 sg13g2_nor2b_1 _3748_ (.A(net328),
    .B_N(net3),
    .Y(_2919_));
 sg13g2_o21ai_1 _3749_ (.B1(\movement_dir[1] ),
    .Y(_2920_),
    .A1(net2),
    .A2(net3));
 sg13g2_o21ai_1 _3750_ (.B1(_2918_),
    .Y(_2921_),
    .A1(_2919_),
    .A2(_2920_));
 sg13g2_and2_1 _3751_ (.A(net1416),
    .B(net352),
    .X(_0003_));
 sg13g2_and2_1 _3752_ (.A(net1416),
    .B(net2),
    .X(_0218_));
 sg13g2_and2_1 _3753_ (.A(net1416),
    .B(net3),
    .X(_0220_));
 sg13g2_nor2_1 _3754_ (.A(_0218_),
    .B(_0220_),
    .Y(_2922_));
 sg13g2_o21ai_1 _3755_ (.B1(_2918_),
    .Y(_2923_),
    .A1(\movement_dir[2] ),
    .A2(_2919_));
 sg13g2_nor2_1 _3756_ (.A(_2922_),
    .B(net329),
    .Y(_0004_));
 sg13g2_nor2_1 _3757_ (.A(\draw_score_inst.score[2] ),
    .B(\draw_score_inst.score[1] ),
    .Y(_2924_));
 sg13g2_nor3_2 _3758_ (.A(net399),
    .B(net335),
    .C(\draw_score_inst.score[1] ),
    .Y(_2925_));
 sg13g2_nand2_1 _3759_ (.Y(_2926_),
    .A(net1307),
    .B(net1308));
 sg13g2_nand3_1 _3760_ (.B(net342),
    .C(net1304),
    .A(_2900_),
    .Y(_2927_));
 sg13g2_nor3_1 _3761_ (.A(net1305),
    .B(_2926_),
    .C(_2927_),
    .Y(_2928_));
 sg13g2_and2_1 _3762_ (.A(net400),
    .B(_2928_),
    .X(_0000_));
 sg13g2_nand2b_1 _3763_ (.Y(_2929_),
    .B(net1416),
    .A_N(game_won));
 sg13g2_nor2_1 _3764_ (.A(game_won),
    .B(game_over),
    .Y(_2930_));
 sg13g2_nor2_1 _3765_ (.A(game_over),
    .B(_2929_),
    .Y(_2931_));
 sg13g2_nand2_1 _3766_ (.Y(_2932_),
    .A(net1416),
    .B(_2930_));
 sg13g2_nand2_2 _3767_ (.Y(_2933_),
    .A(net1317),
    .B(\abullet_x[1] ));
 sg13g2_nand2_1 _3768_ (.Y(_2934_),
    .A(\abullet_x[3] ),
    .B(net1317));
 sg13g2_nand4_1 _3769_ (.B(\abullet_x[3] ),
    .C(net1317),
    .A(net1316),
    .Y(_2935_),
    .D(\abullet_x[1] ));
 sg13g2_nor2_1 _3770_ (.A(_0040_),
    .B(_2935_),
    .Y(_2936_));
 sg13g2_xor2_1 _3771_ (.B(_2936_),
    .A(_0039_),
    .X(_2937_));
 sg13g2_xor2_1 _3772_ (.B(_2935_),
    .A(_0040_),
    .X(_2938_));
 sg13g2_xnor2_1 _3773_ (.Y(_2939_),
    .A(_0040_),
    .B(_2935_));
 sg13g2_nor2_1 _3774_ (.A(_0045_),
    .B(_2933_),
    .Y(_2940_));
 sg13g2_nor2_2 _3775_ (.A(_2862_),
    .B(_2940_),
    .Y(_2941_));
 sg13g2_nor3_2 _3776_ (.A(net1316),
    .B(_0045_),
    .C(_2933_),
    .Y(_2942_));
 sg13g2_nor2_2 _3777_ (.A(_2941_),
    .B(_2942_),
    .Y(_2943_));
 sg13g2_xor2_1 _3778_ (.B(_2933_),
    .A(_0045_),
    .X(_2944_));
 sg13g2_xnor2_1 _3779_ (.Y(_2945_),
    .A(_0045_),
    .B(_2933_));
 sg13g2_nor2_1 _3780_ (.A(\myShooter.shooter_left_x[2] ),
    .B(_2864_),
    .Y(_2946_));
 sg13g2_nor3_1 _3781_ (.A(_2839_),
    .B(\abullet_x[1] ),
    .C(_2946_),
    .Y(_2947_));
 sg13g2_a21o_1 _3782_ (.A2(_2864_),
    .A1(\myShooter.shooter_left_x[2] ),
    .B1(_2947_),
    .X(_2948_));
 sg13g2_nor2b_1 _3783_ (.A(_2948_),
    .B_N(_2933_),
    .Y(_2949_));
 sg13g2_xnor2_1 _3784_ (.Y(_2950_),
    .A(_0046_),
    .B(_2944_));
 sg13g2_a22oi_1 _3785_ (.Y(_2951_),
    .B1(_2945_),
    .B2(net1262),
    .A2(_2943_),
    .A1(net1260));
 sg13g2_o21ai_1 _3786_ (.B1(_2951_),
    .Y(_2952_),
    .A1(_2949_),
    .A2(_2950_));
 sg13g2_o21ai_1 _3787_ (.B1(_2952_),
    .Y(_2953_),
    .A1(net1260),
    .A2(_2943_));
 sg13g2_o21ai_1 _3788_ (.B1(_2953_),
    .Y(_2954_),
    .A1(_0043_),
    .A2(_2938_));
 sg13g2_xnor2_1 _3789_ (.Y(_2955_),
    .A(_0041_),
    .B(_2937_));
 sg13g2_nand2_1 _3790_ (.Y(_2956_),
    .A(_2954_),
    .B(_2955_));
 sg13g2_a21oi_1 _3791_ (.A1(_0043_),
    .A2(_2938_),
    .Y(_2957_),
    .B1(_2956_));
 sg13g2_a21oi_1 _3792_ (.A1(\myShooter.shooter_left_x[6] ),
    .A2(_2937_),
    .Y(_2958_),
    .B1(_2957_));
 sg13g2_nand2_2 _3793_ (.Y(_2959_),
    .A(\abullet_x[6] ),
    .B(\abullet_x[5] ));
 sg13g2_nor3_1 _3794_ (.A(_0035_),
    .B(_2935_),
    .C(_2959_),
    .Y(_2960_));
 sg13g2_o21ai_1 _3795_ (.B1(_0035_),
    .Y(_2961_),
    .A1(_2935_),
    .A2(_2959_));
 sg13g2_nand2b_2 _3796_ (.Y(_2962_),
    .B(_2961_),
    .A_N(_2960_));
 sg13g2_xor2_1 _3797_ (.B(_2962_),
    .A(_0037_),
    .X(_2963_));
 sg13g2_xor2_1 _3798_ (.B(_2960_),
    .A(_0034_),
    .X(_2964_));
 sg13g2_inv_1 _3799_ (.Y(_2965_),
    .A(_2964_));
 sg13g2_a22oi_1 _3800_ (.Y(_2966_),
    .B1(_2964_),
    .B2(net1256),
    .A2(_2962_),
    .A1(net1257));
 sg13g2_o21ai_1 _3801_ (.B1(_2966_),
    .Y(_2967_),
    .A1(_2958_),
    .A2(_2963_));
 sg13g2_nand2_1 _3802_ (.Y(_2968_),
    .A(\abullet_x[8] ),
    .B(net1315));
 sg13g2_nor3_2 _3803_ (.A(_2935_),
    .B(_2959_),
    .C(_2968_),
    .Y(_2969_));
 sg13g2_xnor2_1 _3804_ (.Y(_2970_),
    .A(_0031_),
    .B(_2969_));
 sg13g2_inv_1 _3805_ (.Y(_2971_),
    .A(_2970_));
 sg13g2_xnor2_1 _3806_ (.Y(_2972_),
    .A(_0032_),
    .B(_2970_));
 sg13g2_nor2_1 _3807_ (.A(net1256),
    .B(_2964_),
    .Y(_2973_));
 sg13g2_and2_1 _3808_ (.A(\abullet_x[9] ),
    .B(_2969_),
    .X(_2974_));
 sg13g2_nor3_1 _3809_ (.A(_2972_),
    .B(_2973_),
    .C(_2974_),
    .Y(_2975_));
 sg13g2_nand2_2 _3810_ (.Y(_2976_),
    .A(\myShooter.shooter_left_x[5] ),
    .B(net1260));
 sg13g2_xnor2_1 _3811_ (.Y(_2977_),
    .A(\myShooter.shooter_left_x[5] ),
    .B(net1259));
 sg13g2_nand2_1 _3812_ (.Y(_2978_),
    .A(\abullet_x[5] ),
    .B(_2977_));
 sg13g2_nor2_1 _3813_ (.A(\myShooter.shooter_left_x[1] ),
    .B(_2865_),
    .Y(_2979_));
 sg13g2_nor3_1 _3814_ (.A(\abullet_x[0] ),
    .B(_2946_),
    .C(_2979_),
    .Y(_2980_));
 sg13g2_nand2_1 _3815_ (.Y(_2981_),
    .A(net1262),
    .B(_2863_));
 sg13g2_nand2b_1 _3816_ (.Y(_2982_),
    .B(\abullet_x[3] ),
    .A_N(net1261));
 sg13g2_o21ai_1 _3817_ (.B1(_2982_),
    .Y(_2983_),
    .A1(_2948_),
    .A2(_2980_));
 sg13g2_a22oi_1 _3818_ (.Y(_2984_),
    .B1(_2981_),
    .B2(_2983_),
    .A2(net1316),
    .A1(net1259));
 sg13g2_xnor2_1 _3819_ (.Y(_2985_),
    .A(_0040_),
    .B(_2977_));
 sg13g2_o21ai_1 _3820_ (.B1(_2985_),
    .Y(_2986_),
    .A1(net1259),
    .A2(net1316));
 sg13g2_o21ai_1 _3821_ (.B1(_2978_),
    .Y(_2987_),
    .A1(_2984_),
    .A2(_2986_));
 sg13g2_nor2_1 _3822_ (.A(_0041_),
    .B(_2976_),
    .Y(_2988_));
 sg13g2_xnor2_1 _3823_ (.Y(_2989_),
    .A(_0041_),
    .B(_2976_));
 sg13g2_xnor2_1 _3824_ (.Y(_2990_),
    .A(_0039_),
    .B(_2989_));
 sg13g2_nand2_1 _3825_ (.Y(_2991_),
    .A(_2987_),
    .B(_2990_));
 sg13g2_xor2_1 _3826_ (.B(_2988_),
    .A(_0037_),
    .X(_2992_));
 sg13g2_a22oi_1 _3827_ (.Y(_2993_),
    .B1(_2992_),
    .B2(\abullet_x[7] ),
    .A2(_2989_),
    .A1(\abullet_x[6] ));
 sg13g2_nand4_1 _3828_ (.B(net1258),
    .C(\myShooter.shooter_left_x[5] ),
    .A(net1257),
    .Y(_2994_),
    .D(net1259));
 sg13g2_inv_1 _3829_ (.Y(_2995_),
    .A(_2994_));
 sg13g2_nor2_1 _3830_ (.A(_0047_),
    .B(_2994_),
    .Y(_2996_));
 sg13g2_xor2_1 _3831_ (.B(_2994_),
    .A(_0047_),
    .X(_2997_));
 sg13g2_xor2_1 _3832_ (.B(_2997_),
    .A(_0034_),
    .X(_2998_));
 sg13g2_o21ai_1 _3833_ (.B1(_2998_),
    .Y(_2999_),
    .A1(net1315),
    .A2(_2992_));
 sg13g2_a21o_1 _3834_ (.A2(_2993_),
    .A1(_2991_),
    .B1(_2999_),
    .X(_3000_));
 sg13g2_xor2_1 _3835_ (.B(_2996_),
    .A(_0032_),
    .X(_3001_));
 sg13g2_nor2_1 _3836_ (.A(_2859_),
    .B(_2997_),
    .Y(_3002_));
 sg13g2_a21oi_1 _3837_ (.A1(net1314),
    .A2(_3001_),
    .Y(_3003_),
    .B1(_3002_));
 sg13g2_nand2_1 _3838_ (.Y(_3004_),
    .A(net1256),
    .B(_2995_));
 sg13g2_inv_1 _3839_ (.Y(_3005_),
    .A(_3004_));
 sg13g2_a22oi_1 _3840_ (.Y(_3006_),
    .B1(_3005_),
    .B2(\myShooter.shooter_left_x[9] ),
    .A2(_3003_),
    .A1(_3000_));
 sg13g2_o21ai_1 _3841_ (.B1(_3006_),
    .Y(_3007_),
    .A1(net1314),
    .A2(_3001_));
 sg13g2_nand2_1 _3842_ (.Y(_3008_),
    .A(\abullet_y[5] ),
    .B(\abullet_y[4] ));
 sg13g2_nand4_1 _3843_ (.B(\abullet_y[5] ),
    .C(\abullet_y[4] ),
    .A(net1254),
    .Y(_3009_),
    .D(\abullet_y[3] ));
 sg13g2_nor2_1 _3844_ (.A(\abullet_y[2] ),
    .B(\abullet_y[1] ),
    .Y(_3010_));
 sg13g2_o21ai_1 _3845_ (.B1(\abullet_y[3] ),
    .Y(_3011_),
    .A1(net1255),
    .A2(\abullet_y[1] ));
 sg13g2_nor2_1 _3846_ (.A(_3008_),
    .B(_3011_),
    .Y(_3012_));
 sg13g2_nand2_1 _3847_ (.Y(_3013_),
    .A(net1254),
    .B(_3012_));
 sg13g2_nor2_1 _3848_ (.A(_0050_),
    .B(_3013_),
    .Y(_3014_));
 sg13g2_xnor2_1 _3849_ (.Y(_3015_),
    .A(\abullet_y[8] ),
    .B(_3014_));
 sg13g2_nand2_1 _3850_ (.Y(_3016_),
    .A(\abullet_y[8] ),
    .B(\abullet_y[7] ));
 sg13g2_nor2_1 _3851_ (.A(_3013_),
    .B(_3016_),
    .Y(_3017_));
 sg13g2_xor2_1 _3852_ (.B(_3017_),
    .A(_0049_),
    .X(_3018_));
 sg13g2_inv_1 _3853_ (.Y(_3019_),
    .A(_3018_));
 sg13g2_xor2_1 _3854_ (.B(_3013_),
    .A(_0050_),
    .X(_3020_));
 sg13g2_inv_1 _3855_ (.Y(_3021_),
    .A(_3020_));
 sg13g2_nor3_1 _3856_ (.A(_3015_),
    .B(_3019_),
    .C(_3020_),
    .Y(_3022_));
 sg13g2_o21ai_1 _3857_ (.B1(\abullet_y[6] ),
    .Y(_3023_),
    .A1(\abullet_y[5] ),
    .A2(\abullet_y[4] ));
 sg13g2_o21ai_1 _3858_ (.B1(_2831_),
    .Y(_3024_),
    .A1(_2832_),
    .A2(_3011_));
 sg13g2_nand2b_2 _3859_ (.Y(_3025_),
    .B(_3024_),
    .A_N(_3012_));
 sg13g2_xor2_1 _3860_ (.B(_3011_),
    .A(_0051_),
    .X(_3026_));
 sg13g2_o21ai_1 _3861_ (.B1(_3011_),
    .Y(_3027_),
    .A1(\abullet_y[3] ),
    .A2(net1255));
 sg13g2_inv_1 _3862_ (.Y(_3028_),
    .A(_3027_));
 sg13g2_o21ai_1 _3863_ (.B1(net1254),
    .Y(_3029_),
    .A1(_3026_),
    .A2(_3028_));
 sg13g2_o21ai_1 _3864_ (.B1(_3022_),
    .Y(_3030_),
    .A1(_3025_),
    .A2(_3029_));
 sg13g2_nor2_1 _3865_ (.A(_2970_),
    .B(_2974_),
    .Y(_3031_));
 sg13g2_nor2_1 _3866_ (.A(\abullet_y[9] ),
    .B(\abullet_y[8] ),
    .Y(_3032_));
 sg13g2_nor3_1 _3867_ (.A(\abullet_y[9] ),
    .B(_2828_),
    .C(\abullet_y[7] ),
    .Y(_3033_));
 sg13g2_a21o_1 _3868_ (.A2(_3033_),
    .A1(_3009_),
    .B1(_3032_),
    .X(_3034_));
 sg13g2_nand2_1 _3869_ (.Y(_3035_),
    .A(_3015_),
    .B(_3018_));
 sg13g2_a21oi_1 _3870_ (.A1(\abullet_y[9] ),
    .A2(_3017_),
    .Y(_3036_),
    .B1(_3035_));
 sg13g2_a21oi_1 _3871_ (.A1(\myShooter.shooter_left_x[9] ),
    .A2(_3031_),
    .Y(_3037_),
    .B1(_3036_));
 sg13g2_nand4_1 _3872_ (.B(_3030_),
    .C(_3034_),
    .A(_3007_),
    .Y(_3038_),
    .D(_3037_));
 sg13g2_a21oi_2 _3873_ (.B1(_3038_),
    .Y(_3039_),
    .A2(_2975_),
    .A1(_2967_));
 sg13g2_nor2_1 _3874_ (.A(net1274),
    .B(net1277),
    .Y(_3040_));
 sg13g2_nor2_2 _3875_ (.A(net1272),
    .B(net1274),
    .Y(_3041_));
 sg13g2_nor4_2 _3876_ (.A(net1265),
    .B(net1268),
    .C(net1271),
    .Y(_3042_),
    .D(net1274));
 sg13g2_nor2_1 _3877_ (.A(net1287),
    .B(net1300),
    .Y(_3043_));
 sg13g2_nor2_1 _3878_ (.A(net1290),
    .B(net1296),
    .Y(_3044_));
 sg13g2_inv_1 _3879_ (.Y(_3045_),
    .A(_3044_));
 sg13g2_nor2_2 _3880_ (.A(net1289),
    .B(net1294),
    .Y(_3046_));
 sg13g2_nand2_2 _3881_ (.Y(_3047_),
    .A(net1218),
    .B(net1216));
 sg13g2_nor2_2 _3882_ (.A(net1295),
    .B(net1299),
    .Y(_3048_));
 sg13g2_nand2_1 _3883_ (.Y(_3049_),
    .A(net1213),
    .B(_2850_));
 sg13g2_nor2_1 _3884_ (.A(net1277),
    .B(net1280),
    .Y(_3050_));
 sg13g2_and4_2 _3885_ (.A(_3042_),
    .B(net1193),
    .C(_3048_),
    .D(_3050_),
    .X(_3051_));
 sg13g2_nor4_1 _3886_ (.A(\prev_vpos[7] ),
    .B(\prev_vpos[6] ),
    .C(\prev_vpos[9] ),
    .D(\prev_vpos[8] ),
    .Y(_3052_));
 sg13g2_nor2_1 _3887_ (.A(\prev_vpos[1] ),
    .B(\prev_vpos[0] ),
    .Y(_3053_));
 sg13g2_nor4_1 _3888_ (.A(\prev_vpos[3] ),
    .B(\prev_vpos[2] ),
    .C(\prev_vpos[5] ),
    .D(\prev_vpos[4] ),
    .Y(_3054_));
 sg13g2_nand3_1 _3889_ (.B(_3053_),
    .C(_3054_),
    .A(_3052_),
    .Y(_3055_));
 sg13g2_and2_1 _3890_ (.A(_3051_),
    .B(_3055_),
    .X(_3056_));
 sg13g2_nand2_1 _3891_ (.Y(_3057_),
    .A(_3051_),
    .B(_3055_));
 sg13g2_nor2_1 _3892_ (.A(\draw_score_inst.digit_health[1] ),
    .B(\draw_score_inst.digit_health[0] ),
    .Y(_3058_));
 sg13g2_nor3_1 _3893_ (.A(_0030_),
    .B(net1144),
    .C(_3058_),
    .Y(_3059_));
 sg13g2_nand2_1 _3894_ (.Y(_3060_),
    .A(_3039_),
    .B(_3059_));
 sg13g2_inv_1 _3895_ (.Y(_3061_),
    .A(_3060_));
 sg13g2_a21o_1 _3896_ (.A2(_3060_),
    .A1(net258),
    .B1(net1169),
    .X(_3062_));
 sg13g2_or2_1 _3897_ (.X(_3063_),
    .B(_3060_),
    .A(net258));
 sg13g2_nand2b_2 _3898_ (.Y(_3064_),
    .B(_3063_),
    .A_N(_3062_));
 sg13g2_inv_1 _3899_ (.Y(_0001_),
    .A(_3064_));
 sg13g2_a21o_1 _3900_ (.A2(_3063_),
    .A1(net311),
    .B1(net1169),
    .X(_0002_));
 sg13g2_nor2_2 _3901_ (.A(net1204),
    .B(_2879_),
    .Y(_3065_));
 sg13g2_nand2_2 _3902_ (.Y(_3066_),
    .A(net1411),
    .B(net1396));
 sg13g2_nor2_1 _3903_ (.A(net1198),
    .B(net1196),
    .Y(_3067_));
 sg13g2_nor2_2 _3904_ (.A(_2879_),
    .B(net1200),
    .Y(_3068_));
 sg13g2_nand2_1 _3905_ (.Y(_3069_),
    .A(net1394),
    .B(net1389));
 sg13g2_nand2_2 _3906_ (.Y(_3070_),
    .A(net1388),
    .B(_3065_));
 sg13g2_nor2_1 _3907_ (.A(net1200),
    .B(net1198),
    .Y(_3071_));
 sg13g2_nand2_2 _3908_ (.Y(_3072_),
    .A(net1390),
    .B(net1387));
 sg13g2_nor2_2 _3909_ (.A(_3066_),
    .B(_3072_),
    .Y(_3073_));
 sg13g2_nand2_1 _3910_ (.Y(_3074_),
    .A(net1380),
    .B(_3073_));
 sg13g2_nand2_1 _3911_ (.Y(_3075_),
    .A(net1357),
    .B(net1353));
 sg13g2_nor2_1 _3912_ (.A(net1362),
    .B(net1370),
    .Y(_3076_));
 sg13g2_nand2_1 _3913_ (.Y(_3077_),
    .A(net1202),
    .B(net1194));
 sg13g2_nor4_2 _3914_ (.A(net1375),
    .B(_3074_),
    .C(_3075_),
    .Y(_3078_),
    .D(_3077_));
 sg13g2_nor2_1 _3915_ (.A(net1413),
    .B(_3078_),
    .Y(_3079_));
 sg13g2_nand2b_2 _3916_ (.Y(_3080_),
    .B(net1417),
    .A_N(_3078_));
 sg13g2_and2_1 _3917_ (.A(net220),
    .B(net1088),
    .X(_0081_));
 sg13g2_nor2_1 _3918_ (.A(net1411),
    .B(net1395),
    .Y(_3081_));
 sg13g2_nor3_1 _3919_ (.A(net1414),
    .B(_3065_),
    .C(net1191),
    .Y(_0082_));
 sg13g2_o21ai_1 _3920_ (.B1(net1089),
    .Y(_3082_),
    .A1(net1390),
    .A2(_3065_));
 sg13g2_nor2b_1 _3921_ (.A(_3082_),
    .B_N(_3070_),
    .Y(_0083_));
 sg13g2_nor2_1 _3922_ (.A(_0042_),
    .B(_3066_),
    .Y(_3083_));
 sg13g2_xnor2_1 _3923_ (.Y(_3084_),
    .A(net1386),
    .B(_3083_));
 sg13g2_nor2_1 _3924_ (.A(_3080_),
    .B(net388),
    .Y(_0084_));
 sg13g2_o21ai_1 _3925_ (.B1(net1416),
    .Y(_3085_),
    .A1(net1380),
    .A2(_3073_));
 sg13g2_nor2b_1 _3926_ (.A(_3085_),
    .B_N(_3074_),
    .Y(_0085_));
 sg13g2_nor2_1 _3927_ (.A(net1378),
    .B(_3072_),
    .Y(_3086_));
 sg13g2_xnor2_1 _3928_ (.Y(_3087_),
    .A(net1195),
    .B(_3086_));
 sg13g2_o21ai_1 _3929_ (.B1(net1089),
    .Y(_3088_),
    .A1(_3066_),
    .A2(_3087_));
 sg13g2_a21oi_1 _3930_ (.A1(net1195),
    .A2(net411),
    .Y(_0086_),
    .B1(_3088_));
 sg13g2_nand2_1 _3931_ (.Y(_3089_),
    .A(net1381),
    .B(net1376));
 sg13g2_nand3_1 _3932_ (.B(net1376),
    .C(_3073_),
    .A(net1381),
    .Y(_3090_));
 sg13g2_xnor2_1 _3933_ (.Y(_3091_),
    .A(net1194),
    .B(_3090_));
 sg13g2_nor2_1 _3934_ (.A(_3080_),
    .B(_3091_),
    .Y(_0087_));
 sg13g2_nor2_1 _3935_ (.A(net1368),
    .B(_3090_),
    .Y(_3092_));
 sg13g2_xnor2_1 _3936_ (.Y(_3093_),
    .A(net1363),
    .B(_3092_));
 sg13g2_nor2_1 _3937_ (.A(_3080_),
    .B(net386),
    .Y(_0088_));
 sg13g2_nand2_2 _3938_ (.Y(_3094_),
    .A(net1362),
    .B(net1370));
 sg13g2_nor2_1 _3939_ (.A(_3090_),
    .B(_3094_),
    .Y(_3095_));
 sg13g2_nor2_1 _3940_ (.A(net1357),
    .B(net1202),
    .Y(_3096_));
 sg13g2_o21ai_1 _3941_ (.B1(net1089),
    .Y(_3097_),
    .A1(net1357),
    .A2(_3095_));
 sg13g2_a21oi_1 _3942_ (.A1(net1357),
    .A2(_3095_),
    .Y(_0089_),
    .B1(_3097_));
 sg13g2_nor3_1 _3943_ (.A(net1356),
    .B(_3090_),
    .C(_3094_),
    .Y(_3098_));
 sg13g2_o21ai_1 _3944_ (.B1(net1089),
    .Y(_3099_),
    .A1(net1353),
    .A2(_3098_));
 sg13g2_a21oi_1 _3945_ (.A1(net1353),
    .A2(_3098_),
    .Y(_0090_),
    .B1(_3099_));
 sg13g2_nor2_2 _3946_ (.A(_2843_),
    .B(_2844_),
    .Y(_3100_));
 sg13g2_nand3_1 _3947_ (.B(net1277),
    .C(_3100_),
    .A(net1269),
    .Y(_3101_));
 sg13g2_a21oi_1 _3948_ (.A1(net1363),
    .A2(net1353),
    .Y(_3102_),
    .B1(net1414));
 sg13g2_nand4_1 _3949_ (.B(_3075_),
    .C(_3101_),
    .A(_2841_),
    .Y(_3103_),
    .D(_3102_));
 sg13g2_nand2b_1 _3950_ (.Y(_3104_),
    .B(_2943_),
    .A_N(net1379));
 sg13g2_nand2_1 _3951_ (.Y(_3105_),
    .A(\abullet_x[0] ),
    .B(_3081_));
 sg13g2_xnor2_1 _3952_ (.Y(_3106_),
    .A(net1317),
    .B(\abullet_x[1] ));
 sg13g2_o21ai_1 _3953_ (.B1(_3105_),
    .Y(_3107_),
    .A1(_2916_),
    .A2(_3106_));
 sg13g2_o21ai_1 _3954_ (.B1(net1395),
    .Y(_3108_),
    .A1(_2866_),
    .A2(net1411));
 sg13g2_a221oi_1 _3955_ (.B2(_2865_),
    .C1(_3107_),
    .B1(_3108_),
    .A1(_2916_),
    .Y(_3109_),
    .A2(_3106_));
 sg13g2_a221oi_1 _3956_ (.B2(net1392),
    .C1(_3109_),
    .B1(_3106_),
    .A1(net1384),
    .Y(_3110_),
    .A2(_2945_));
 sg13g2_o21ai_1 _3957_ (.B1(net1379),
    .Y(_3111_),
    .A1(_2941_),
    .A2(_2942_));
 sg13g2_o21ai_1 _3958_ (.B1(_3111_),
    .Y(_3112_),
    .A1(net1384),
    .A2(_2945_));
 sg13g2_o21ai_1 _3959_ (.B1(_3104_),
    .Y(_3113_),
    .A1(_3110_),
    .A2(_3112_));
 sg13g2_xnor2_1 _3960_ (.Y(_3114_),
    .A(_2915_),
    .B(_2938_));
 sg13g2_a22oi_1 _3961_ (.Y(_3115_),
    .B1(_3113_),
    .B2(_3114_),
    .A2(_2939_),
    .A1(net1377));
 sg13g2_xor2_1 _3962_ (.B(_2937_),
    .A(net1368),
    .X(_3116_));
 sg13g2_a22oi_1 _3963_ (.Y(_3117_),
    .B1(_2962_),
    .B2(net1363),
    .A2(_2937_),
    .A1(net1372));
 sg13g2_o21ai_1 _3964_ (.B1(_3117_),
    .Y(_3118_),
    .A1(_3115_),
    .A2(_3116_));
 sg13g2_xor2_1 _3965_ (.B(_2964_),
    .A(net1356),
    .X(_3119_));
 sg13g2_o21ai_1 _3966_ (.B1(_3118_),
    .Y(_3120_),
    .A1(net1363),
    .A2(_2962_));
 sg13g2_a22oi_1 _3967_ (.Y(_3121_),
    .B1(_2971_),
    .B2(net1354),
    .A2(_2964_),
    .A1(net1358));
 sg13g2_o21ai_1 _3968_ (.B1(_3121_),
    .Y(_3122_),
    .A1(_3119_),
    .A2(_3120_));
 sg13g2_o21ai_1 _3969_ (.B1(_3122_),
    .Y(_3123_),
    .A1(net1353),
    .A2(_2971_));
 sg13g2_xnor2_1 _3970_ (.Y(_3124_),
    .A(_2833_),
    .B(_3010_));
 sg13g2_nand2_2 _3971_ (.Y(_3125_),
    .A(net1255),
    .B(\abullet_y[1] ));
 sg13g2_nand2b_2 _3972_ (.Y(_3126_),
    .B(_3125_),
    .A_N(_3010_));
 sg13g2_inv_1 _3973_ (.Y(_3127_),
    .A(_3126_));
 sg13g2_xnor2_1 _3974_ (.Y(_3128_),
    .A(_2904_),
    .B(_3126_));
 sg13g2_o21ai_1 _3975_ (.B1(_3128_),
    .Y(_3129_),
    .A1(\abullet_y[1] ),
    .A2(\barrier1.bar_rom.row_index[1] ));
 sg13g2_a22oi_1 _3976_ (.Y(_3130_),
    .B1(_3127_),
    .B2(net1293),
    .A2(_3124_),
    .A1(net1288));
 sg13g2_nand2_1 _3977_ (.Y(_3131_),
    .A(_3129_),
    .B(_3130_));
 sg13g2_o21ai_1 _3978_ (.B1(_3131_),
    .Y(_3132_),
    .A1(net1288),
    .A2(_3124_));
 sg13g2_o21ai_1 _3979_ (.B1(_3132_),
    .Y(_3133_),
    .A1(net1278),
    .A2(_3026_));
 sg13g2_xnor2_1 _3980_ (.Y(_3134_),
    .A(_2906_),
    .B(_3025_));
 sg13g2_a21oi_1 _3981_ (.A1(net1278),
    .A2(_3026_),
    .Y(_3135_),
    .B1(_3134_));
 sg13g2_a22oi_1 _3982_ (.Y(_3136_),
    .B1(_3133_),
    .B2(_3135_),
    .A2(_3025_),
    .A1(net1277));
 sg13g2_xnor2_1 _3983_ (.Y(_3137_),
    .A(net1254),
    .B(_3012_));
 sg13g2_xnor2_1 _3984_ (.Y(_3138_),
    .A(_2907_),
    .B(_3137_));
 sg13g2_a22oi_1 _3985_ (.Y(_3139_),
    .B1(_3137_),
    .B2(net1275),
    .A2(_3021_),
    .A1(net1272));
 sg13g2_o21ai_1 _3986_ (.B1(_3139_),
    .Y(_3140_),
    .A1(_3136_),
    .A2(_3138_));
 sg13g2_xor2_1 _3987_ (.B(_3015_),
    .A(net1267),
    .X(_3141_));
 sg13g2_a21oi_1 _3988_ (.A1(_2843_),
    .A2(_3020_),
    .Y(_3142_),
    .B1(_3141_));
 sg13g2_nand2_1 _3989_ (.Y(_3143_),
    .A(_3140_),
    .B(_3142_));
 sg13g2_a22oi_1 _3990_ (.Y(_3144_),
    .B1(_3018_),
    .B2(net1264),
    .A2(_3015_),
    .A1(net1270));
 sg13g2_nor2_1 _3991_ (.A(net1264),
    .B(_3018_),
    .Y(_3145_));
 sg13g2_a221oi_1 _3992_ (.B2(_3144_),
    .C1(_3145_),
    .B1(_3143_),
    .A1(\abullet_y[9] ),
    .Y(_3146_),
    .A2(_3017_));
 sg13g2_nand2_1 _3993_ (.Y(_3147_),
    .A(\abullet_x[1] ),
    .B(_3108_));
 sg13g2_a22oi_1 _3994_ (.Y(_3148_),
    .B1(_3105_),
    .B2(_3147_),
    .A2(net1392),
    .A1(_2864_));
 sg13g2_a221oi_1 _3995_ (.B2(\abullet_x[3] ),
    .C1(_3148_),
    .B1(net1199),
    .A1(net1317),
    .Y(_3149_),
    .A2(net1201));
 sg13g2_a221oi_1 _3996_ (.B2(_2862_),
    .C1(_3149_),
    .B1(net1382),
    .A1(_2863_),
    .Y(_3150_),
    .A2(net1386));
 sg13g2_a221oi_1 _3997_ (.B2(\abullet_x[5] ),
    .C1(_3150_),
    .B1(net1195),
    .A1(net1316),
    .Y(_3151_),
    .A2(net1197));
 sg13g2_a221oi_1 _3998_ (.B2(_2860_),
    .C1(_3151_),
    .B1(net1371),
    .A1(_2861_),
    .Y(_3152_),
    .A2(net1377));
 sg13g2_a21o_1 _3999_ (.A2(net1194),
    .A1(\abullet_x[6] ),
    .B1(_3152_),
    .X(_3153_));
 sg13g2_o21ai_1 _4000_ (.B1(_3153_),
    .Y(_3154_),
    .A1(net1315),
    .A2(net1203));
 sg13g2_a22oi_1 _4001_ (.Y(_3155_),
    .B1(net1203),
    .B2(net1315),
    .A2(_2875_),
    .A1(\abullet_x[8] ));
 sg13g2_nor2_1 _4002_ (.A(net1314),
    .B(_2877_),
    .Y(_3156_));
 sg13g2_a221oi_1 _4003_ (.B2(_3155_),
    .C1(_3156_),
    .B1(_3154_),
    .A1(_2859_),
    .Y(_3157_),
    .A2(net1358));
 sg13g2_nor2_1 _4004_ (.A(_2828_),
    .B(net1270),
    .Y(_3158_));
 sg13g2_a22oi_1 _4005_ (.Y(_3159_),
    .B1(net1214),
    .B2(\abullet_y[1] ),
    .A2(net1216),
    .A1(net1255));
 sg13g2_a221oi_1 _4006_ (.B2(_2834_),
    .C1(_3159_),
    .B1(net1293),
    .A1(_2833_),
    .Y(_3160_),
    .A2(net1288));
 sg13g2_a221oi_1 _4007_ (.B2(\abullet_y[3] ),
    .C1(_3160_),
    .B1(net1220),
    .A1(\abullet_y[4] ),
    .Y(_3161_),
    .A2(net1222));
 sg13g2_a221oi_1 _4008_ (.B2(_2832_),
    .C1(_3161_),
    .B1(net1281),
    .A1(_2831_),
    .Y(_3162_),
    .A2(net1277));
 sg13g2_a21oi_1 _4009_ (.A1(\abullet_y[5] ),
    .A2(net1223),
    .Y(_3163_),
    .B1(_3162_));
 sg13g2_a21o_1 _4010_ (.A2(net1275),
    .A1(_2830_),
    .B1(_3163_),
    .X(_3164_));
 sg13g2_a22oi_1 _4011_ (.Y(_3165_),
    .B1(_2844_),
    .B2(net1254),
    .A2(net1224),
    .A1(\abullet_y[7] ));
 sg13g2_nor2_1 _4012_ (.A(\abullet_y[8] ),
    .B(_2842_),
    .Y(_3166_));
 sg13g2_a221oi_1 _4013_ (.B2(_3165_),
    .C1(_3166_),
    .B1(_3164_),
    .A1(_2829_),
    .Y(_3167_),
    .A2(net1272));
 sg13g2_nand2b_1 _4014_ (.Y(_3168_),
    .B(net1264),
    .A_N(\abullet_y[9] ));
 sg13g2_o21ai_1 _4015_ (.B1(_3168_),
    .Y(_3169_),
    .A1(_3158_),
    .A2(_3167_));
 sg13g2_a22oi_1 _4016_ (.Y(_3170_),
    .B1(net1314),
    .B2(_2877_),
    .A2(net1225),
    .A1(\abullet_y[9] ));
 sg13g2_nand3_1 _4017_ (.B(_3169_),
    .C(_3170_),
    .A(net1319),
    .Y(_3171_));
 sg13g2_nor3_1 _4018_ (.A(_3146_),
    .B(_3157_),
    .C(_3171_),
    .Y(_3172_));
 sg13g2_o21ai_1 _4019_ (.B1(_3172_),
    .Y(_3173_),
    .A1(_2974_),
    .A2(_3123_));
 sg13g2_nor2_1 _4020_ (.A(_0033_),
    .B(_3069_),
    .Y(_3174_));
 sg13g2_xor2_1 _4021_ (.B(_3069_),
    .A(_0033_),
    .X(_3175_));
 sg13g2_a22oi_1 _4022_ (.Y(_3176_),
    .B1(net1193),
    .B2(_3048_),
    .A2(_3045_),
    .A1(net1285));
 sg13g2_nand2_2 _4023_ (.Y(_3177_),
    .A(net1216),
    .B(_3048_));
 sg13g2_nand3_1 _4024_ (.B(net1407),
    .C(_3177_),
    .A(net1285),
    .Y(_3178_));
 sg13g2_o21ai_1 _4025_ (.B1(_3178_),
    .Y(_3179_),
    .A1(net1407),
    .A2(_3176_));
 sg13g2_nor2_1 _4026_ (.A(net1394),
    .B(net1389),
    .Y(_3180_));
 sg13g2_nor2_2 _4027_ (.A(net1215),
    .B(_2850_),
    .Y(_3181_));
 sg13g2_nand2_2 _4028_ (.Y(_3182_),
    .A(net1291),
    .B(net1295));
 sg13g2_nand2_2 _4029_ (.Y(_3183_),
    .A(net1295),
    .B(_3181_));
 sg13g2_a21o_1 _4030_ (.A2(_3182_),
    .A1(net1285),
    .B1(net1204),
    .X(_3184_));
 sg13g2_nand3_1 _4031_ (.B(_3183_),
    .C(_3184_),
    .A(net1285),
    .Y(_3185_));
 sg13g2_nand2_1 _4032_ (.Y(_3186_),
    .A(_3180_),
    .B(_3185_));
 sg13g2_o21ai_1 _4033_ (.B1(_3186_),
    .Y(_3187_),
    .A1(_3069_),
    .A2(_3179_));
 sg13g2_nor2_2 _4034_ (.A(net1215),
    .B(net1296),
    .Y(_3188_));
 sg13g2_nand2_2 _4035_ (.Y(_3189_),
    .A(net1292),
    .B(net1213));
 sg13g2_nor2_2 _4036_ (.A(net1290),
    .B(net1213),
    .Y(_3190_));
 sg13g2_nor2_2 _4037_ (.A(_3188_),
    .B(_3190_),
    .Y(_3191_));
 sg13g2_or2_2 _4038_ (.X(_3192_),
    .B(_3190_),
    .A(_3188_));
 sg13g2_nand2_1 _4039_ (.Y(_3193_),
    .A(_0048_),
    .B(_3192_));
 sg13g2_nor2_1 _4040_ (.A(net1293),
    .B(_3048_),
    .Y(_3194_));
 sg13g2_nand2_2 _4041_ (.Y(_3195_),
    .A(net1215),
    .B(net1163));
 sg13g2_nand2_1 _4042_ (.Y(_3196_),
    .A(_3177_),
    .B(_3182_));
 sg13g2_a21oi_2 _4043_ (.B1(_3196_),
    .Y(_3197_),
    .A2(_3192_),
    .A1(_0048_));
 sg13g2_nand2_1 _4044_ (.Y(_3198_),
    .A(net1285),
    .B(_3197_));
 sg13g2_a21oi_1 _4045_ (.A1(net1285),
    .A2(_3197_),
    .Y(_3199_),
    .B1(net1204));
 sg13g2_nor2_2 _4046_ (.A(net1218),
    .B(net1290),
    .Y(_3200_));
 sg13g2_nor2_1 _4047_ (.A(net1219),
    .B(net1163),
    .Y(_3201_));
 sg13g2_nor3_1 _4048_ (.A(net1402),
    .B(_3200_),
    .C(_3201_),
    .Y(_3202_));
 sg13g2_nor3_1 _4049_ (.A(_0044_),
    .B(_3199_),
    .C(_3202_),
    .Y(_3203_));
 sg13g2_nor3_1 _4050_ (.A(_3068_),
    .B(net1190),
    .C(_3203_),
    .Y(_3204_));
 sg13g2_o21ai_1 _4051_ (.B1(_3175_),
    .Y(_3205_),
    .A1(_3187_),
    .A2(_3204_));
 sg13g2_nand3_1 _4052_ (.B(net1191),
    .C(_3183_),
    .A(net1285),
    .Y(_3206_));
 sg13g2_o21ai_1 _4053_ (.B1(_3206_),
    .Y(_3207_),
    .A1(net1394),
    .A2(_3178_));
 sg13g2_nand3b_1 _4054_ (.B(net1394),
    .C(_3184_),
    .Y(_3208_),
    .A_N(_3202_));
 sg13g2_nor2_1 _4055_ (.A(net1290),
    .B(_2905_),
    .Y(_3209_));
 sg13g2_nand2_2 _4056_ (.Y(_3210_),
    .A(net1283),
    .B(_3182_));
 sg13g2_xnor2_1 _4057_ (.Y(_3211_),
    .A(net1279),
    .B(_3210_));
 sg13g2_a21oi_2 _4058_ (.B1(net1288),
    .Y(_3212_),
    .A2(net1295),
    .A1(net1290));
 sg13g2_nand2b_1 _4059_ (.Y(_3213_),
    .B(net1280),
    .A_N(net1189));
 sg13g2_xnor2_1 _4060_ (.Y(_3214_),
    .A(_2845_),
    .B(_3213_));
 sg13g2_nor2_2 _4061_ (.A(_3211_),
    .B(_3214_),
    .Y(_3215_));
 sg13g2_nor2_1 _4062_ (.A(net1198),
    .B(net1380),
    .Y(_3216_));
 sg13g2_nand2_1 _4063_ (.Y(_3217_),
    .A(_3068_),
    .B(_3216_));
 sg13g2_nand2_1 _4064_ (.Y(_3218_),
    .A(net1378),
    .B(_3217_));
 sg13g2_xnor2_1 _4065_ (.Y(_3219_),
    .A(net1196),
    .B(_3174_));
 sg13g2_o21ai_1 _4066_ (.B1(_3219_),
    .Y(_3220_),
    .A1(net1375),
    .A2(_3218_));
 sg13g2_a21oi_1 _4067_ (.A1(net1375),
    .A2(_3218_),
    .Y(_3221_),
    .B1(_3220_));
 sg13g2_or2_1 _4068_ (.X(_3222_),
    .B(_3198_),
    .A(\lgA2.rx[0] ));
 sg13g2_nor2_1 _4069_ (.A(net1190),
    .B(_3207_),
    .Y(_3223_));
 sg13g2_a221oi_1 _4070_ (.B2(_3208_),
    .C1(_3068_),
    .B1(_3223_),
    .A1(net1190),
    .Y(_3224_),
    .A2(_3222_));
 sg13g2_nor4_1 _4071_ (.A(net1370),
    .B(net1360),
    .C(_3041_),
    .D(_3100_),
    .Y(_3225_));
 sg13g2_nand2_1 _4072_ (.Y(_3226_),
    .A(net1358),
    .B(_2877_));
 sg13g2_nand2_1 _4073_ (.Y(_3227_),
    .A(net1362),
    .B(_3226_));
 sg13g2_nor2_1 _4074_ (.A(net1357),
    .B(_2877_),
    .Y(_3228_));
 sg13g2_o21ai_1 _4075_ (.B1(_3227_),
    .Y(_3229_),
    .A1(net1363),
    .A2(_3228_));
 sg13g2_nor4_1 _4076_ (.A(net1265),
    .B(net1268),
    .C(_0014_),
    .D(_3229_),
    .Y(_3230_));
 sg13g2_nand4_1 _4077_ (.B(_3221_),
    .C(_3225_),
    .A(_3215_),
    .Y(_3231_),
    .D(_3230_));
 sg13g2_o21ai_1 _4078_ (.B1(_3205_),
    .Y(_3232_),
    .A1(_3175_),
    .A2(_3224_));
 sg13g2_o21ai_1 _4079_ (.B1(_3173_),
    .Y(_3233_),
    .A1(_3231_),
    .A2(_3232_));
 sg13g2_nand2_2 _4080_ (.Y(_3234_),
    .A(net1349),
    .B(\pb_x[1] ));
 sg13g2_nand4_1 _4081_ (.B(net1346),
    .C(net1348),
    .A(net1344),
    .Y(_3235_),
    .D(net1350));
 sg13g2_nor2_1 _4082_ (.A(net1342),
    .B(_3235_),
    .Y(_3236_));
 sg13g2_xnor2_1 _4083_ (.Y(_3237_),
    .A(net1342),
    .B(_3235_));
 sg13g2_inv_2 _4084_ (.Y(_3238_),
    .A(net1162));
 sg13g2_nor2_1 _4085_ (.A(_0069_),
    .B(_3234_),
    .Y(_3239_));
 sg13g2_xnor2_1 _4086_ (.Y(_3240_),
    .A(_0068_),
    .B(_3239_));
 sg13g2_xnor2_1 _4087_ (.Y(_3241_),
    .A(_2886_),
    .B(_3239_));
 sg13g2_xor2_1 _4088_ (.B(_3234_),
    .A(_0069_),
    .X(_3242_));
 sg13g2_xnor2_1 _4089_ (.Y(_3243_),
    .A(_0069_),
    .B(_3234_));
 sg13g2_a21o_1 _4090_ (.A2(net1210),
    .A1(net1351),
    .B1(_2879_),
    .X(_3244_));
 sg13g2_xnor2_1 _4091_ (.Y(_3245_),
    .A(net1348),
    .B(net1350));
 sg13g2_xor2_1 _4092_ (.B(net1188),
    .A(_0042_),
    .X(_3246_));
 sg13g2_a221oi_1 _4093_ (.B2(_2873_),
    .C1(_3246_),
    .B1(_3244_),
    .A1(net1351),
    .Y(_3247_),
    .A2(net1191));
 sg13g2_a221oi_1 _4094_ (.B2(net1392),
    .C1(_3247_),
    .B1(net1188),
    .A1(net1384),
    .Y(_3248_),
    .A2(_3243_));
 sg13g2_a21o_1 _4095_ (.A2(_3242_),
    .A1(net1199),
    .B1(_3248_),
    .X(_3249_));
 sg13g2_o21ai_1 _4096_ (.B1(_3249_),
    .Y(_3250_),
    .A1(net1379),
    .A2(net1143));
 sg13g2_xnor2_1 _4097_ (.Y(_3251_),
    .A(_2915_),
    .B(net1162));
 sg13g2_a21oi_1 _4098_ (.A1(net1379),
    .A2(net1143),
    .Y(_3252_),
    .B1(_3251_));
 sg13g2_a22oi_1 _4099_ (.Y(_3253_),
    .B1(_3250_),
    .B2(_3252_),
    .A2(net1162),
    .A1(net1377));
 sg13g2_xor2_1 _4100_ (.B(_3236_),
    .A(net1337),
    .X(_3254_));
 sg13g2_xnor2_1 _4101_ (.Y(_3255_),
    .A(net1337),
    .B(_3236_));
 sg13g2_xnor2_1 _4102_ (.Y(_3256_),
    .A(net1366),
    .B(net1140));
 sg13g2_nand2b_1 _4103_ (.Y(_3257_),
    .B(_3256_),
    .A_N(_3253_));
 sg13g2_nand2_2 _4104_ (.Y(_3258_),
    .A(net1338),
    .B(net1343));
 sg13g2_nor2_1 _4105_ (.A(_3235_),
    .B(_3258_),
    .Y(_3259_));
 sg13g2_nor3_2 _4106_ (.A(_0060_),
    .B(_3235_),
    .C(_3258_),
    .Y(_3260_));
 sg13g2_xnor2_1 _4107_ (.Y(_3261_),
    .A(_0060_),
    .B(_3259_));
 sg13g2_xor2_1 _4108_ (.B(_3259_),
    .A(_0060_),
    .X(_3262_));
 sg13g2_a22oi_1 _4109_ (.Y(_3263_),
    .B1(_3262_),
    .B2(net1364),
    .A2(net1140),
    .A1(net1372));
 sg13g2_xor2_1 _4110_ (.B(_3260_),
    .A(net1331),
    .X(_3264_));
 sg13g2_xnor2_1 _4111_ (.Y(_3265_),
    .A(net1331),
    .B(_3260_));
 sg13g2_xnor2_1 _4112_ (.Y(_3266_),
    .A(net1355),
    .B(_3265_));
 sg13g2_a221oi_1 _4113_ (.B2(_3257_),
    .C1(_3266_),
    .B1(_3263_),
    .A1(net1203),
    .Y(_3267_),
    .A2(net1139));
 sg13g2_nand2_1 _4114_ (.Y(_3268_),
    .A(net1333),
    .B(net1334));
 sg13g2_nor3_2 _4115_ (.A(_3235_),
    .B(_3258_),
    .C(_3268_),
    .Y(_3269_));
 sg13g2_xnor2_1 _4116_ (.Y(_3270_),
    .A(_0058_),
    .B(_3269_));
 sg13g2_xor2_1 _4117_ (.B(_3269_),
    .A(_0058_),
    .X(_3271_));
 sg13g2_a221oi_1 _4118_ (.B2(net1354),
    .C1(_3267_),
    .B1(net1134),
    .A1(net1359),
    .Y(_3272_),
    .A2(net1136));
 sg13g2_and2_1 _4119_ (.A(net1329),
    .B(_3269_),
    .X(_3273_));
 sg13g2_nand2_2 _4120_ (.Y(_3274_),
    .A(net1329),
    .B(_3269_));
 sg13g2_o21ai_1 _4121_ (.B1(_3274_),
    .Y(_3275_),
    .A1(net1354),
    .A2(net1134));
 sg13g2_nor2_1 _4122_ (.A(\pb_y[2] ),
    .B(\pb_y[1] ),
    .Y(_3276_));
 sg13g2_o21ai_1 _4123_ (.B1(net1324),
    .Y(_3277_),
    .A1(net1325),
    .A2(\pb_y[1] ));
 sg13g2_nor2_1 _4124_ (.A(_2890_),
    .B(_3277_),
    .Y(_3278_));
 sg13g2_and4_1 _4125_ (.A(\pb_y[7] ),
    .B(net1322),
    .C(net1323),
    .D(_3278_),
    .X(_3279_));
 sg13g2_and2_1 _4126_ (.A(\pb_y[8] ),
    .B(_3279_),
    .X(_3280_));
 sg13g2_nor2_1 _4127_ (.A(net1321),
    .B(_3279_),
    .Y(_3281_));
 sg13g2_nor2_1 _4128_ (.A(_3280_),
    .B(_3281_),
    .Y(_3282_));
 sg13g2_o21ai_1 _4129_ (.B1(net1270),
    .Y(_3283_),
    .A1(_3280_),
    .A2(_3281_));
 sg13g2_xnor2_1 _4130_ (.Y(_3284_),
    .A(net1323),
    .B(_3278_));
 sg13g2_xor2_1 _4131_ (.B(_3277_),
    .A(_0073_),
    .X(_3285_));
 sg13g2_xnor2_1 _4132_ (.Y(_3286_),
    .A(_0073_),
    .B(_3277_));
 sg13g2_nand2_1 _4133_ (.Y(_3287_),
    .A(\pb_y[0] ),
    .B(_3048_));
 sg13g2_nand2_2 _4134_ (.Y(_3288_),
    .A(net1296),
    .B(net1299));
 sg13g2_a21oi_1 _4135_ (.A1(net1212),
    .A2(\pb_y[0] ),
    .Y(_3289_),
    .B1(net1214));
 sg13g2_a21oi_1 _4136_ (.A1(net1326),
    .A2(_3287_),
    .Y(_3290_),
    .B1(_3289_));
 sg13g2_nand2_1 _4137_ (.Y(_3291_),
    .A(net1325),
    .B(net1326));
 sg13g2_nor2b_1 _4138_ (.A(_3276_),
    .B_N(_3291_),
    .Y(_3292_));
 sg13g2_xnor2_1 _4139_ (.Y(_3293_),
    .A(_2904_),
    .B(_3292_));
 sg13g2_nor3_1 _4140_ (.A(net1324),
    .B(net1325),
    .C(\pb_y[1] ),
    .Y(_3294_));
 sg13g2_xnor2_1 _4141_ (.Y(_3295_),
    .A(\pb_y[3] ),
    .B(_3276_));
 sg13g2_inv_1 _4142_ (.Y(_3296_),
    .A(_3295_));
 sg13g2_a22oi_1 _4143_ (.Y(_3297_),
    .B1(_3296_),
    .B2(net1289),
    .A2(_3292_),
    .A1(net1294));
 sg13g2_o21ai_1 _4144_ (.B1(_3297_),
    .Y(_3298_),
    .A1(_3290_),
    .A2(_3293_));
 sg13g2_a22oi_1 _4145_ (.Y(_3299_),
    .B1(_3295_),
    .B2(net1221),
    .A2(_3285_),
    .A1(net1279));
 sg13g2_nand2_1 _4146_ (.Y(_3300_),
    .A(_3298_),
    .B(_3299_));
 sg13g2_o21ai_1 _4147_ (.B1(_3300_),
    .Y(_3301_),
    .A1(net1279),
    .A2(_3285_));
 sg13g2_xnor2_1 _4148_ (.Y(_3302_),
    .A(_0013_),
    .B(_3284_));
 sg13g2_a22oi_1 _4149_ (.Y(_3303_),
    .B1(_3301_),
    .B2(_3302_),
    .A2(_3284_),
    .A1(net1276));
 sg13g2_nor3_1 _4150_ (.A(_2890_),
    .B(_0072_),
    .C(_3277_),
    .Y(_3304_));
 sg13g2_xnor2_1 _4151_ (.Y(_3305_),
    .A(net1322),
    .B(_3304_));
 sg13g2_xnor2_1 _4152_ (.Y(_3306_),
    .A(_2907_),
    .B(_3305_));
 sg13g2_nand3_1 _4153_ (.B(net1323),
    .C(_3278_),
    .A(net1322),
    .Y(_3307_));
 sg13g2_xnor2_1 _4154_ (.Y(_3308_),
    .A(_0071_),
    .B(_3307_));
 sg13g2_inv_1 _4155_ (.Y(_3309_),
    .A(_3308_));
 sg13g2_a22oi_1 _4156_ (.Y(_3310_),
    .B1(_3308_),
    .B2(net1272),
    .A2(_3305_),
    .A1(net1273));
 sg13g2_o21ai_1 _4157_ (.B1(_3310_),
    .Y(_3311_),
    .A1(_3303_),
    .A2(_3306_));
 sg13g2_nand2_1 _4158_ (.Y(_3312_),
    .A(net1224),
    .B(_3309_));
 sg13g2_xor2_1 _4159_ (.B(_3282_),
    .A(net1267),
    .X(_3313_));
 sg13g2_nand3_1 _4160_ (.B(_3312_),
    .C(_3313_),
    .A(_3311_),
    .Y(_3314_));
 sg13g2_nand2b_1 _4161_ (.Y(_3315_),
    .B(net1264),
    .A_N(\pb_y[9] ));
 sg13g2_nand2_1 _4162_ (.Y(_3316_),
    .A(net1225),
    .B(\pb_y[9] ));
 sg13g2_nand2b_1 _4163_ (.Y(_3317_),
    .B(_3316_),
    .A_N(_3280_));
 sg13g2_a22oi_1 _4164_ (.Y(_3318_),
    .B1(_3315_),
    .B2(_3317_),
    .A2(_3314_),
    .A1(_3283_));
 sg13g2_nor2_1 _4165_ (.A(net1275),
    .B(_2888_),
    .Y(_3319_));
 sg13g2_a221oi_1 _4166_ (.B2(_3287_),
    .C1(_3289_),
    .B1(_2893_),
    .A1(net1294),
    .Y(_3320_),
    .A2(_2892_));
 sg13g2_a221oi_1 _4167_ (.B2(net1217),
    .C1(_3320_),
    .B1(net1325),
    .A1(net1221),
    .Y(_3321_),
    .A2(net1324));
 sg13g2_a221oi_1 _4168_ (.B2(net1289),
    .C1(_3321_),
    .B1(_2891_),
    .A1(net1280),
    .Y(_3322_),
    .A2(_2890_));
 sg13g2_a221oi_1 _4169_ (.B2(net1222),
    .C1(_3322_),
    .B1(\pb_y[4] ),
    .A1(net1223),
    .Y(_3323_),
    .A2(net1323));
 sg13g2_a21oi_1 _4170_ (.A1(net1276),
    .A2(_2889_),
    .Y(_3324_),
    .B1(_3323_));
 sg13g2_a22oi_1 _4171_ (.Y(_3325_),
    .B1(_2888_),
    .B2(net1275),
    .A2(_2887_),
    .A1(net1272));
 sg13g2_o21ai_1 _4172_ (.B1(_3325_),
    .Y(_3326_),
    .A1(_3319_),
    .A2(_3324_));
 sg13g2_nand2_1 _4173_ (.Y(_3327_),
    .A(_2842_),
    .B(net1321));
 sg13g2_nand2_1 _4174_ (.Y(_3328_),
    .A(net1224),
    .B(\pb_y[7] ));
 sg13g2_nand4_1 _4175_ (.B(_3326_),
    .C(_3327_),
    .A(_3316_),
    .Y(_3329_),
    .D(_3328_));
 sg13g2_nand2b_1 _4176_ (.Y(_3330_),
    .B(net1270),
    .A_N(net1321));
 sg13g2_nand3_1 _4177_ (.B(_3329_),
    .C(_3330_),
    .A(_3315_),
    .Y(_3331_));
 sg13g2_o21ai_1 _4178_ (.B1(net1327),
    .Y(_3332_),
    .A1(_3316_),
    .A2(_3330_));
 sg13g2_a22oi_1 _4179_ (.Y(_0273_),
    .B1(net1354),
    .B2(_2867_),
    .A2(net1359),
    .A1(_2868_));
 sg13g2_nor2_1 _4180_ (.A(_2867_),
    .B(net1354),
    .Y(_0274_));
 sg13g2_nor2_1 _4181_ (.A(_2869_),
    .B(net1371),
    .Y(_0275_));
 sg13g2_a21oi_1 _4182_ (.A1(net1351),
    .A2(net1191),
    .Y(_0276_),
    .B1(net1350));
 sg13g2_o21ai_1 _4183_ (.B1(_3244_),
    .Y(_0277_),
    .A1(net1348),
    .A2(net1201));
 sg13g2_a22oi_1 _4184_ (.Y(_0278_),
    .B1(net1199),
    .B2(net1346),
    .A2(net1201),
    .A1(net1348));
 sg13g2_o21ai_1 _4185_ (.B1(_0278_),
    .Y(_0279_),
    .A1(_0276_),
    .A2(_0277_));
 sg13g2_a22oi_1 _4186_ (.Y(_0280_),
    .B1(net1382),
    .B2(_2871_),
    .A2(net1384),
    .A1(_2872_));
 sg13g2_nor2_1 _4187_ (.A(_2871_),
    .B(net1382),
    .Y(_0281_));
 sg13g2_a221oi_1 _4188_ (.B2(_0280_),
    .C1(_0281_),
    .B1(_0279_),
    .A1(net1343),
    .Y(_0282_),
    .A2(_2883_));
 sg13g2_a221oi_1 _4189_ (.B2(_2869_),
    .C1(_0282_),
    .B1(net1371),
    .A1(_2870_),
    .Y(_0283_),
    .A2(net1377));
 sg13g2_nand2b_1 _4190_ (.Y(_0284_),
    .B(net1365),
    .A_N(net1334));
 sg13g2_o21ai_1 _4191_ (.B1(_0284_),
    .Y(_0285_),
    .A1(_0275_),
    .A2(_0283_));
 sg13g2_a221oi_1 _4192_ (.B2(net1334),
    .C1(_0274_),
    .B1(net1203),
    .A1(net1333),
    .Y(_0286_),
    .A2(_2875_));
 sg13g2_nand3_1 _4193_ (.B(_0285_),
    .C(_0286_),
    .A(_0273_),
    .Y(_0287_));
 sg13g2_o21ai_1 _4194_ (.B1(_0287_),
    .Y(_0288_),
    .A1(_0273_),
    .A2(_0274_));
 sg13g2_o21ai_1 _4195_ (.B1(_3331_),
    .Y(_0289_),
    .A1(_3280_),
    .A2(_3315_));
 sg13g2_o21ai_1 _4196_ (.B1(_0288_),
    .Y(_0290_),
    .A1(_3272_),
    .A2(_3275_));
 sg13g2_nor4_2 _4197_ (.A(_3318_),
    .B(_3332_),
    .C(_0289_),
    .Y(_0291_),
    .D(_0290_));
 sg13g2_nor3_2 _4198_ (.A(\barrier_health[2][1] ),
    .B(\barrier_health[2][0] ),
    .C(\barrier_health[2][2] ),
    .Y(_0292_));
 sg13g2_inv_1 _4199_ (.Y(_0293_),
    .A(_0292_));
 sg13g2_nor2_2 _4200_ (.A(_2875_),
    .B(net1356),
    .Y(_0294_));
 sg13g2_nand2b_2 _4201_ (.Y(_0295_),
    .B(net1359),
    .A_N(net1355));
 sg13g2_a21oi_1 _4202_ (.A1(_2875_),
    .A2(net1352),
    .Y(_0296_),
    .B1(net1356));
 sg13g2_nand2b_1 _4203_ (.Y(_0297_),
    .B(net1357),
    .A_N(net1352));
 sg13g2_nand3_1 _4204_ (.B(_0296_),
    .C(_0297_),
    .A(net1202),
    .Y(_0298_));
 sg13g2_nand2_1 _4205_ (.Y(_0299_),
    .A(net1378),
    .B(_3072_));
 sg13g2_xnor2_1 _4206_ (.Y(_0300_),
    .A(net1374),
    .B(_0299_));
 sg13g2_a21oi_1 _4207_ (.A1(net1196),
    .A2(net1192),
    .Y(_0301_),
    .B1(net1195));
 sg13g2_xnor2_1 _4208_ (.Y(_0302_),
    .A(net1370),
    .B(_0301_));
 sg13g2_nor4_1 _4209_ (.A(_0292_),
    .B(_0298_),
    .C(_0300_),
    .D(_0302_),
    .Y(_0303_));
 sg13g2_nor2_1 _4210_ (.A(net1388),
    .B(net1387),
    .Y(_0304_));
 sg13g2_nor2_2 _4211_ (.A(_3071_),
    .B(_0304_),
    .Y(_0305_));
 sg13g2_or2_1 _4212_ (.X(_0306_),
    .B(_0304_),
    .A(_3071_));
 sg13g2_nor2b_1 _4213_ (.A(net1394),
    .B_N(\lgA2.rx[0] ),
    .Y(_0307_));
 sg13g2_nor3_1 _4214_ (.A(net1285),
    .B(_2904_),
    .C(net1163),
    .Y(_0308_));
 sg13g2_nor2_2 _4215_ (.A(net1283),
    .B(_3182_),
    .Y(_0309_));
 sg13g2_nor3_2 _4216_ (.A(net1215),
    .B(net1283),
    .C(net1187),
    .Y(_0310_));
 sg13g2_a22oi_1 _4217_ (.Y(_0311_),
    .B1(_0310_),
    .B2(_3065_),
    .A2(_0308_),
    .A1(_0307_));
 sg13g2_nand2_1 _4218_ (.Y(_0312_),
    .A(net1201),
    .B(_0311_));
 sg13g2_nand2_2 _4219_ (.Y(_0313_),
    .A(net1292),
    .B(net1163));
 sg13g2_nand3_1 _4220_ (.B(net1191),
    .C(_0313_),
    .A(net1283),
    .Y(_0314_));
 sg13g2_a21oi_2 _4221_ (.B1(net1292),
    .Y(_0315_),
    .A2(net1300),
    .A1(net1297));
 sg13g2_nand4_1 _4222_ (.B(net1395),
    .C(net1283),
    .A(net1204),
    .Y(_0316_),
    .D(_0315_));
 sg13g2_nand2_1 _4223_ (.Y(_0317_),
    .A(net1297),
    .B(net1395));
 sg13g2_nand3_1 _4224_ (.B(_3046_),
    .C(_0317_),
    .A(net1407),
    .Y(_0318_));
 sg13g2_nand3_1 _4225_ (.B(_0316_),
    .C(_0318_),
    .A(_0314_),
    .Y(_0319_));
 sg13g2_o21ai_1 _4226_ (.B1(_0312_),
    .Y(_0320_),
    .A1(net1200),
    .A2(_0319_));
 sg13g2_xnor2_1 _4227_ (.Y(_0321_),
    .A(net1196),
    .B(net1192));
 sg13g2_nor2_2 _4228_ (.A(net1283),
    .B(_0313_),
    .Y(_0322_));
 sg13g2_nand3_1 _4229_ (.B(_2905_),
    .C(net1163),
    .A(net1291),
    .Y(_0323_));
 sg13g2_nor2_1 _4230_ (.A(net1388),
    .B(_0323_),
    .Y(_0324_));
 sg13g2_nand2_1 _4231_ (.Y(_0325_),
    .A(net1200),
    .B(_0322_));
 sg13g2_nand2_1 _4232_ (.Y(_0326_),
    .A(net1191),
    .B(_0309_));
 sg13g2_o21ai_1 _4233_ (.B1(_0326_),
    .Y(_0327_),
    .A1(net1191),
    .A2(_0323_));
 sg13g2_a21oi_1 _4234_ (.A1(net1388),
    .A2(_0327_),
    .Y(_0328_),
    .B1(_0324_));
 sg13g2_nand4_1 _4235_ (.B(_2879_),
    .C(net1283),
    .A(net1407),
    .Y(_0329_),
    .D(_0315_));
 sg13g2_nor2_1 _4236_ (.A(net1407),
    .B(_3047_),
    .Y(_0330_));
 sg13g2_o21ai_1 _4237_ (.B1(_0330_),
    .Y(_0331_),
    .A1(net1214),
    .A2(net1395));
 sg13g2_nand3_1 _4238_ (.B(_3065_),
    .C(_0313_),
    .A(net1283),
    .Y(_0332_));
 sg13g2_nand3_1 _4239_ (.B(_0331_),
    .C(_0332_),
    .A(_0329_),
    .Y(_0333_));
 sg13g2_a22oi_1 _4240_ (.Y(_0334_),
    .B1(_0310_),
    .B2(_0307_),
    .A2(_0308_),
    .A1(_3065_));
 sg13g2_nand2_1 _4241_ (.Y(_0335_),
    .A(net1388),
    .B(_0334_));
 sg13g2_o21ai_1 _4242_ (.B1(_0335_),
    .Y(_0336_),
    .A1(net1388),
    .A2(_0333_));
 sg13g2_nand2_1 _4243_ (.Y(_0337_),
    .A(net1390),
    .B(_0322_));
 sg13g2_nor2_1 _4244_ (.A(_3065_),
    .B(_0323_),
    .Y(_0338_));
 sg13g2_a21oi_1 _4245_ (.A1(_3065_),
    .A2(_0309_),
    .Y(_0339_),
    .B1(_0338_));
 sg13g2_o21ai_1 _4246_ (.B1(_0337_),
    .Y(_0340_),
    .A1(net1388),
    .A2(_0339_));
 sg13g2_inv_1 _4247_ (.Y(_0341_),
    .A(_0340_));
 sg13g2_mux4_1 _4248_ (.S0(_0305_),
    .A0(_0320_),
    .A1(_0328_),
    .A2(_0341_),
    .A3(_0336_),
    .S1(_0321_),
    .X(_0342_));
 sg13g2_nor2_2 _4249_ (.A(net1387),
    .B(net1381),
    .Y(_0343_));
 sg13g2_nor3_2 _4250_ (.A(net1389),
    .B(net1387),
    .C(net1380),
    .Y(_0344_));
 sg13g2_nor2_2 _4251_ (.A(net1195),
    .B(_0344_),
    .Y(_0345_));
 sg13g2_xor2_1 _4252_ (.B(_0345_),
    .A(net1368),
    .X(_0346_));
 sg13g2_xnor2_1 _4253_ (.Y(_0347_),
    .A(net1374),
    .B(_0344_));
 sg13g2_nand2_2 _4254_ (.Y(_0348_),
    .A(net1369),
    .B(_0345_));
 sg13g2_a21oi_1 _4255_ (.A1(net1362),
    .A2(net1360),
    .Y(_0349_),
    .B1(_2875_));
 sg13g2_nor2_1 _4256_ (.A(net1360),
    .B(_0348_),
    .Y(_0350_));
 sg13g2_o21ai_1 _4257_ (.B1(net1360),
    .Y(_0351_),
    .A1(_3096_),
    .A2(_0348_));
 sg13g2_nand4_1 _4258_ (.B(_0346_),
    .C(_0347_),
    .A(_2877_),
    .Y(_0352_),
    .D(_0351_));
 sg13g2_nor3_2 _4259_ (.A(_0349_),
    .B(_0350_),
    .C(_0352_),
    .Y(_0353_));
 sg13g2_nor3_2 _4260_ (.A(\barrier_health[0][1] ),
    .B(\barrier_health[0][0] ),
    .C(\barrier_health[0][2] ),
    .Y(_0354_));
 sg13g2_xnor2_1 _4261_ (.Y(_0355_),
    .A(net1378),
    .B(_0304_));
 sg13g2_mux2_1 _4262_ (.A0(_0328_),
    .A1(_0336_),
    .S(_0355_),
    .X(_0356_));
 sg13g2_o21ai_1 _4263_ (.B1(_0353_),
    .Y(_0357_),
    .A1(_0305_),
    .A2(_0356_));
 sg13g2_a221oi_1 _4264_ (.B2(_0355_),
    .C1(_0306_),
    .B1(_0341_),
    .A1(net1378),
    .Y(_0358_),
    .A2(_0320_));
 sg13g2_nor3_1 _4265_ (.A(_0354_),
    .B(_0357_),
    .C(_0358_),
    .Y(_0359_));
 sg13g2_nor2_1 _4266_ (.A(net1388),
    .B(_0319_),
    .Y(_0360_));
 sg13g2_a21oi_1 _4267_ (.A1(net1389),
    .A2(_0311_),
    .Y(_0361_),
    .B1(_0360_));
 sg13g2_nor2_1 _4268_ (.A(net1387),
    .B(net1196),
    .Y(_0362_));
 sg13g2_nand2_1 _4269_ (.Y(_0363_),
    .A(net1200),
    .B(_0327_));
 sg13g2_nand2_1 _4270_ (.Y(_0364_),
    .A(_0337_),
    .B(_0363_));
 sg13g2_o21ai_1 _4271_ (.B1(_0325_),
    .Y(_0365_),
    .A1(net1200),
    .A2(_0339_));
 sg13g2_nor3_1 _4272_ (.A(net1380),
    .B(net1375),
    .C(net1369),
    .Y(_0366_));
 sg13g2_nor2_1 _4273_ (.A(net1202),
    .B(_0366_),
    .Y(_0367_));
 sg13g2_a21oi_1 _4274_ (.A1(_0297_),
    .A2(_0367_),
    .Y(_0368_),
    .B1(net1356));
 sg13g2_nor2_1 _4275_ (.A(net1352),
    .B(_0367_),
    .Y(_0369_));
 sg13g2_nor2_1 _4276_ (.A(_0296_),
    .B(_0369_),
    .Y(_0370_));
 sg13g2_nor2_2 _4277_ (.A(_0368_),
    .B(_0370_),
    .Y(_0371_));
 sg13g2_nor3_2 _4278_ (.A(\barrier_health[3][1] ),
    .B(\barrier_health[3][0] ),
    .C(\barrier_health[3][2] ),
    .Y(_0372_));
 sg13g2_xnor2_1 _4279_ (.Y(_0373_),
    .A(net1381),
    .B(net1376));
 sg13g2_nor4_1 _4280_ (.A(net1369),
    .B(net1360),
    .C(_0372_),
    .D(_0373_),
    .Y(_0374_));
 sg13g2_nand2_1 _4281_ (.Y(_0375_),
    .A(_0371_),
    .B(_0374_));
 sg13g2_a221oi_1 _4282_ (.B2(_0343_),
    .C1(_0375_),
    .B1(_0365_),
    .A1(_3067_),
    .Y(_0376_),
    .A2(_0364_));
 sg13g2_nor2_1 _4283_ (.A(net1200),
    .B(_0333_),
    .Y(_0377_));
 sg13g2_a21oi_2 _4284_ (.B1(_0377_),
    .Y(_0378_),
    .A2(_0334_),
    .A1(net1200));
 sg13g2_a22oi_1 _4285_ (.Y(_0379_),
    .B1(_0378_),
    .B2(_3216_),
    .A2(_0362_),
    .A1(_0361_));
 sg13g2_nand2_1 _4286_ (.Y(_0380_),
    .A(_3067_),
    .B(_0365_));
 sg13g2_nand4_1 _4287_ (.B(net1369),
    .C(net1356),
    .A(net1362),
    .Y(_0381_),
    .D(_3226_));
 sg13g2_nand2_1 _4288_ (.Y(_0382_),
    .A(_2877_),
    .B(_3094_));
 sg13g2_o21ai_1 _4289_ (.B1(_0381_),
    .Y(_0383_),
    .A1(net1356),
    .A2(_0382_));
 sg13g2_nor3_2 _4290_ (.A(\barrier_health[1][1] ),
    .B(\barrier_health[1][0] ),
    .C(\barrier_health[1][2] ),
    .Y(_0384_));
 sg13g2_xnor2_1 _4291_ (.Y(_0385_),
    .A(net1369),
    .B(net1360));
 sg13g2_nor4_1 _4292_ (.A(net1368),
    .B(_3228_),
    .C(_0384_),
    .D(_0385_),
    .Y(_0386_));
 sg13g2_nor2_1 _4293_ (.A(net1380),
    .B(net1195),
    .Y(_0387_));
 sg13g2_xnor2_1 _4294_ (.Y(_0388_),
    .A(net1376),
    .B(_0343_));
 sg13g2_nand4_1 _4295_ (.B(_0383_),
    .C(_0386_),
    .A(_0380_),
    .Y(_0389_),
    .D(_0388_));
 sg13g2_a21oi_1 _4296_ (.A1(_0362_),
    .A2(_0364_),
    .Y(_0390_),
    .B1(_0389_));
 sg13g2_a22oi_1 _4297_ (.Y(_0391_),
    .B1(_0378_),
    .B2(_0343_),
    .A2(_0361_),
    .A1(_3216_));
 sg13g2_a22oi_1 _4298_ (.Y(_0392_),
    .B1(_0376_),
    .B2(_0379_),
    .A2(_0342_),
    .A1(_0303_));
 sg13g2_a21oi_1 _4299_ (.A1(_0390_),
    .A2(_0391_),
    .Y(_0393_),
    .B1(_0359_));
 sg13g2_o21ai_1 _4300_ (.B1(net1268),
    .Y(_0394_),
    .A1(net1272),
    .A2(net1273));
 sg13g2_nand2_1 _4301_ (.Y(_0395_),
    .A(net1224),
    .B(net1273));
 sg13g2_nor4_1 _4302_ (.A(net1276),
    .B(net1281),
    .C(net1266),
    .D(_0395_),
    .Y(_0396_));
 sg13g2_o21ai_1 _4303_ (.B1(_0396_),
    .Y(_0397_),
    .A1(_0017_),
    .A2(_0394_));
 sg13g2_a21o_1 _4304_ (.A2(_0394_),
    .A1(_0017_),
    .B1(_0397_),
    .X(_0398_));
 sg13g2_a21o_1 _4305_ (.A2(_0393_),
    .A1(_0392_),
    .B1(_0398_),
    .X(_0399_));
 sg13g2_nand2_1 _4306_ (.Y(_0400_),
    .A(\myShooter.shooter_left_x[8] ),
    .B(_2875_));
 sg13g2_xnor2_1 _4307_ (.Y(_0401_),
    .A(net1256),
    .B(net1358));
 sg13g2_nor2_1 _4308_ (.A(net1258),
    .B(_2884_),
    .Y(_0402_));
 sg13g2_nand2_1 _4309_ (.Y(_0403_),
    .A(net1258),
    .B(net1194));
 sg13g2_nand2b_1 _4310_ (.Y(_0404_),
    .B(_0403_),
    .A_N(_0402_));
 sg13g2_nor2_1 _4311_ (.A(net1261),
    .B(net1198),
    .Y(_0405_));
 sg13g2_nand2b_1 _4312_ (.Y(_0406_),
    .B(net1393),
    .A_N(net1263));
 sg13g2_xor2_1 _4313_ (.B(net1393),
    .A(net1263),
    .X(_0407_));
 sg13g2_xnor2_1 _4314_ (.Y(_0408_),
    .A(\myShooter.shooter_left_x[1] ),
    .B(net1396));
 sg13g2_and2_1 _4315_ (.A(net1411),
    .B(_0408_),
    .X(_0409_));
 sg13g2_nand2_1 _4316_ (.Y(_0410_),
    .A(net1411),
    .B(_0408_));
 sg13g2_a21oi_1 _4317_ (.A1(_2839_),
    .A2(net1395),
    .Y(_0411_),
    .B1(_0409_));
 sg13g2_o21ai_1 _4318_ (.B1(_0406_),
    .Y(_0412_),
    .A1(_0407_),
    .A2(_0411_));
 sg13g2_nand2_1 _4319_ (.Y(_0413_),
    .A(net1261),
    .B(net1198));
 sg13g2_nand2b_1 _4320_ (.Y(_0414_),
    .B(_0413_),
    .A_N(_0405_));
 sg13g2_a21oi_1 _4321_ (.A1(_0412_),
    .A2(_0413_),
    .Y(_0415_),
    .B1(_0405_));
 sg13g2_xor2_1 _4322_ (.B(net1376),
    .A(\myShooter.shooter_left_x[5] ),
    .X(_0416_));
 sg13g2_nor2_1 _4323_ (.A(net1259),
    .B(net1197),
    .Y(_0417_));
 sg13g2_nor2b_1 _4324_ (.A(net1383),
    .B_N(net1259),
    .Y(_0418_));
 sg13g2_nor4_1 _4325_ (.A(_0415_),
    .B(_0416_),
    .C(_0417_),
    .D(_0418_),
    .Y(_0419_));
 sg13g2_nand2b_1 _4326_ (.Y(_0420_),
    .B(_0417_),
    .A_N(_0416_));
 sg13g2_a21oi_1 _4327_ (.A1(_2838_),
    .A2(net1376),
    .Y(_0421_),
    .B1(_0419_));
 sg13g2_nand2_1 _4328_ (.Y(_0422_),
    .A(_0420_),
    .B(_0421_));
 sg13g2_a221oi_1 _4329_ (.B2(_0422_),
    .C1(_0402_),
    .B1(_0403_),
    .A1(_2836_),
    .Y(_0423_),
    .A2(net1363));
 sg13g2_a21o_1 _4330_ (.A2(net1202),
    .A1(\myShooter.shooter_left_x[7] ),
    .B1(_0423_),
    .X(_0424_));
 sg13g2_nand2_1 _4331_ (.Y(_0425_),
    .A(_0401_),
    .B(_0424_));
 sg13g2_or2_1 _4332_ (.X(_0426_),
    .B(_0424_),
    .A(_0401_));
 sg13g2_xnor2_1 _4333_ (.Y(_0427_),
    .A(_0404_),
    .B(_0422_));
 sg13g2_nand2_1 _4334_ (.Y(_0428_),
    .A(_0416_),
    .B(_0418_));
 sg13g2_nand2_1 _4335_ (.Y(_0429_),
    .A(_0420_),
    .B(_0428_));
 sg13g2_a21o_1 _4336_ (.A2(_0429_),
    .A1(_0415_),
    .B1(_0419_),
    .X(_0430_));
 sg13g2_xnor2_1 _4337_ (.Y(_0431_),
    .A(net1265),
    .B(_0394_));
 sg13g2_xnor2_1 _4338_ (.Y(_0432_),
    .A(net1257),
    .B(net1363));
 sg13g2_xor2_1 _4339_ (.B(net1354),
    .A(\myShooter.shooter_left_x[9] ),
    .X(_0433_));
 sg13g2_xor2_1 _4340_ (.B(net1276),
    .A(net1273),
    .X(_0434_));
 sg13g2_xor2_1 _4341_ (.B(_0015_),
    .A(net1273),
    .X(_0435_));
 sg13g2_nand2_1 _4342_ (.Y(_0436_),
    .A(net1280),
    .B(net1289));
 sg13g2_a21o_1 _4343_ (.A2(net1218),
    .A1(_2846_),
    .B1(net1267),
    .X(_0437_));
 sg13g2_nor4_1 _4344_ (.A(_0013_),
    .B(_0434_),
    .C(_0435_),
    .D(_0437_),
    .Y(_0438_));
 sg13g2_xnor2_1 _4345_ (.Y(_0439_),
    .A(_0400_),
    .B(_0433_));
 sg13g2_xnor2_1 _4346_ (.Y(_0440_),
    .A(_0403_),
    .B(_0432_));
 sg13g2_nand4_1 _4347_ (.B(_0436_),
    .C(_0438_),
    .A(_0431_),
    .Y(_0441_),
    .D(_0440_));
 sg13g2_nand2b_1 _4348_ (.Y(_0442_),
    .B(_0430_),
    .A_N(_0441_));
 sg13g2_nor3_1 _4349_ (.A(_0427_),
    .B(_0439_),
    .C(_0442_),
    .Y(_0443_));
 sg13g2_xnor2_1 _4350_ (.Y(_0444_),
    .A(_0407_),
    .B(_0411_));
 sg13g2_a21oi_1 _4351_ (.A1(net1292),
    .A2(net1163),
    .Y(_0445_),
    .B1(net1286));
 sg13g2_nor2_1 _4352_ (.A(net1286),
    .B(_0313_),
    .Y(_0446_));
 sg13g2_a21oi_1 _4353_ (.A1(net1286),
    .A2(_2904_),
    .Y(_0447_),
    .B1(_0445_));
 sg13g2_nor2_1 _4354_ (.A(net1286),
    .B(_3191_),
    .Y(_0448_));
 sg13g2_a21oi_1 _4355_ (.A1(_0444_),
    .A2(_0447_),
    .Y(_0449_),
    .B1(net1211));
 sg13g2_o21ai_1 _4356_ (.B1(_0449_),
    .Y(_0450_),
    .A1(_0444_),
    .A2(_0448_));
 sg13g2_nor2_2 _4357_ (.A(net1287),
    .B(_3189_),
    .Y(_0451_));
 sg13g2_nand2_2 _4358_ (.Y(_0452_),
    .A(net1219),
    .B(_3188_));
 sg13g2_nand3_1 _4359_ (.B(net1300),
    .C(_0010_),
    .A(net1297),
    .Y(_0453_));
 sg13g2_a21oi_1 _4360_ (.A1(_3189_),
    .A2(_0453_),
    .Y(_0454_),
    .B1(net1286));
 sg13g2_a21oi_1 _4361_ (.A1(net1286),
    .A2(_2904_),
    .Y(_0455_),
    .B1(net1189));
 sg13g2_o21ai_1 _4362_ (.B1(_0408_),
    .Y(_0456_),
    .A1(_0444_),
    .A2(_0454_));
 sg13g2_a21o_1 _4363_ (.A2(_0455_),
    .A1(_0444_),
    .B1(_0456_),
    .X(_0457_));
 sg13g2_nor2_2 _4364_ (.A(net1411),
    .B(_0408_),
    .Y(_0458_));
 sg13g2_nor2_1 _4365_ (.A(_0409_),
    .B(_0458_),
    .Y(_0459_));
 sg13g2_nand3_1 _4366_ (.B(_0457_),
    .C(_0459_),
    .A(_0450_),
    .Y(_0460_));
 sg13g2_xnor2_1 _4367_ (.Y(_0461_),
    .A(_0412_),
    .B(_0414_));
 sg13g2_nor2_1 _4368_ (.A(_3177_),
    .B(_0408_),
    .Y(_0462_));
 sg13g2_a21oi_1 _4369_ (.A1(net1286),
    .A2(_0462_),
    .Y(_0463_),
    .B1(_0446_));
 sg13g2_o21ai_1 _4370_ (.B1(net1189),
    .Y(_0464_),
    .A1(_3177_),
    .A2(_0408_));
 sg13g2_a21oi_1 _4371_ (.A1(_0444_),
    .A2(_0463_),
    .Y(_0465_),
    .B1(_0459_));
 sg13g2_o21ai_1 _4372_ (.B1(_0465_),
    .Y(_0466_),
    .A1(_0444_),
    .A2(_0464_));
 sg13g2_nand3_1 _4373_ (.B(_0461_),
    .C(_0466_),
    .A(_0460_),
    .Y(_0467_));
 sg13g2_nor3_1 _4374_ (.A(_0409_),
    .B(_0458_),
    .C(_0463_),
    .Y(_0468_));
 sg13g2_a221oi_1 _4375_ (.B2(_0447_),
    .C1(_0468_),
    .B1(_0458_),
    .A1(_0409_),
    .Y(_0469_),
    .A2(_0455_));
 sg13g2_o21ai_1 _4376_ (.B1(_0458_),
    .Y(_0470_),
    .A1(net1286),
    .A2(_3191_));
 sg13g2_o21ai_1 _4377_ (.B1(_0470_),
    .Y(_0471_),
    .A1(_0410_),
    .A2(_0454_));
 sg13g2_a21o_1 _4378_ (.A2(_0464_),
    .A1(_0459_),
    .B1(_0471_),
    .X(_0472_));
 sg13g2_a21oi_1 _4379_ (.A1(_0444_),
    .A2(_0472_),
    .Y(_0473_),
    .B1(_0461_));
 sg13g2_o21ai_1 _4380_ (.B1(_0473_),
    .Y(_0474_),
    .A1(_0444_),
    .A2(_0469_));
 sg13g2_nand2_1 _4381_ (.Y(_0475_),
    .A(_0467_),
    .B(_0474_));
 sg13g2_nand4_1 _4382_ (.B(_0426_),
    .C(_0443_),
    .A(_0425_),
    .Y(_0476_),
    .D(_0475_));
 sg13g2_nand2_2 _4383_ (.Y(_0477_),
    .A(_0399_),
    .B(_0476_));
 sg13g2_nor2_1 _4384_ (.A(_0291_),
    .B(_0477_),
    .Y(_0478_));
 sg13g2_or2_1 _4385_ (.X(_0479_),
    .B(net1243),
    .A(net1241));
 sg13g2_or3_2 _4386_ (.A(net1241),
    .B(net1242),
    .C(net1246),
    .X(_0480_));
 sg13g2_nor2_1 _4387_ (.A(net1246),
    .B(net1250),
    .Y(_0481_));
 sg13g2_nor3_2 _4388_ (.A(net1242),
    .B(net1246),
    .C(net1251),
    .Y(_0482_));
 sg13g2_nor2_1 _4389_ (.A(net1251),
    .B(_0480_),
    .Y(_0483_));
 sg13g2_nor3_2 _4390_ (.A(net1237),
    .B(net1251),
    .C(_0480_),
    .Y(_0484_));
 sg13g2_nand2_1 _4391_ (.Y(_0485_),
    .A(net1233),
    .B(net1234));
 sg13g2_nor2_1 _4392_ (.A(_0484_),
    .B(_0485_),
    .Y(_0486_));
 sg13g2_o21ai_1 _4393_ (.B1(_2821_),
    .Y(_0487_),
    .A1(net1226),
    .A2(_0484_));
 sg13g2_nand2b_2 _4394_ (.Y(_0488_),
    .B(_0487_),
    .A_N(_0486_));
 sg13g2_xnor2_1 _4395_ (.Y(_0489_),
    .A(_0038_),
    .B(_0488_));
 sg13g2_xnor2_1 _4396_ (.Y(_0490_),
    .A(net1236),
    .B(_0483_));
 sg13g2_nor2_1 _4397_ (.A(net1366),
    .B(_0490_),
    .Y(_0491_));
 sg13g2_nand2_1 _4398_ (.Y(_0492_),
    .A(net1366),
    .B(_0490_));
 sg13g2_nand2b_1 _4399_ (.Y(_0493_),
    .B(_0492_),
    .A_N(_0491_));
 sg13g2_xnor2_1 _4400_ (.Y(_0494_),
    .A(_0075_),
    .B(_0482_));
 sg13g2_xnor2_1 _4401_ (.Y(_0495_),
    .A(_0076_),
    .B(_0481_));
 sg13g2_inv_1 _4402_ (.Y(_0496_),
    .A(net1160));
 sg13g2_nand2_1 _4403_ (.Y(_0497_),
    .A(net1383),
    .B(_0496_));
 sg13g2_xnor2_1 _4404_ (.Y(_0498_),
    .A(net1379),
    .B(net1160));
 sg13g2_xor2_1 _4405_ (.B(net1251),
    .A(net1248),
    .X(_0499_));
 sg13g2_inv_1 _4406_ (.Y(_0500_),
    .A(_0499_));
 sg13g2_xnor2_1 _4407_ (.Y(_0501_),
    .A(_0033_),
    .B(_0499_));
 sg13g2_nand2_1 _4408_ (.Y(_0502_),
    .A(net1249),
    .B(net1391));
 sg13g2_nor2b_2 _4409_ (.A(net1396),
    .B_N(net1252),
    .Y(_0503_));
 sg13g2_nor2_1 _4410_ (.A(net1249),
    .B(net1391),
    .Y(_0504_));
 sg13g2_xor2_1 _4411_ (.B(net1391),
    .A(net1249),
    .X(_0505_));
 sg13g2_o21ai_1 _4412_ (.B1(_0502_),
    .Y(_0506_),
    .A1(_0503_),
    .A2(_0504_));
 sg13g2_a22oi_1 _4413_ (.Y(_0507_),
    .B1(_0501_),
    .B2(_0506_),
    .A2(_0499_),
    .A1(net1385));
 sg13g2_o21ai_1 _4414_ (.B1(_0497_),
    .Y(_0508_),
    .A1(_0498_),
    .A2(_0507_));
 sg13g2_xnor2_1 _4415_ (.Y(_0509_),
    .A(_2915_),
    .B(_0494_));
 sg13g2_nand2_1 _4416_ (.Y(_0510_),
    .A(_0508_),
    .B(_0509_));
 sg13g2_o21ai_1 _4417_ (.B1(_0510_),
    .Y(_0511_),
    .A1(_2883_),
    .A2(_0494_));
 sg13g2_a21oi_1 _4418_ (.A1(_0492_),
    .A2(_0511_),
    .Y(_0512_),
    .B1(_0491_));
 sg13g2_xnor2_1 _4419_ (.Y(_0513_),
    .A(net1227),
    .B(_0484_));
 sg13g2_xor2_1 _4420_ (.B(_0513_),
    .A(net1361),
    .X(_0514_));
 sg13g2_nand2_1 _4421_ (.Y(_0515_),
    .A(net1365),
    .B(_0513_));
 sg13g2_o21ai_1 _4422_ (.B1(_0515_),
    .Y(_0516_),
    .A1(_0512_),
    .A2(_0514_));
 sg13g2_xnor2_1 _4423_ (.Y(_0517_),
    .A(_0512_),
    .B(_0514_));
 sg13g2_xnor2_1 _4424_ (.Y(_0518_),
    .A(_0493_),
    .B(_0511_));
 sg13g2_nor2_1 _4425_ (.A(_0294_),
    .B(_0489_),
    .Y(_0519_));
 sg13g2_xnor2_1 _4426_ (.Y(_0520_),
    .A(_0078_),
    .B(_0486_));
 sg13g2_xor2_1 _4427_ (.B(_0520_),
    .A(_0008_),
    .X(_0521_));
 sg13g2_xor2_1 _4428_ (.B(_0507_),
    .A(_0498_),
    .X(_0522_));
 sg13g2_xor2_1 _4429_ (.B(_0509_),
    .A(_0508_),
    .X(_0523_));
 sg13g2_xnor2_1 _4430_ (.Y(_0524_),
    .A(_0519_),
    .B(_0521_));
 sg13g2_nor4_1 _4431_ (.A(_0518_),
    .B(_0522_),
    .C(_0523_),
    .D(_0524_),
    .Y(_0525_));
 sg13g2_xnor2_1 _4432_ (.Y(_0526_),
    .A(_0489_),
    .B(_0516_));
 sg13g2_and3_2 _4433_ (.X(_0527_),
    .A(_0517_),
    .B(_0525_),
    .C(_0526_));
 sg13g2_xnor2_1 _4434_ (.Y(_0528_),
    .A(_0503_),
    .B(_0505_));
 sg13g2_xor2_1 _4435_ (.B(_0505_),
    .A(_0503_),
    .X(_0529_));
 sg13g2_nor2_2 _4436_ (.A(net1252),
    .B(_2879_),
    .Y(_0530_));
 sg13g2_nor2_2 _4437_ (.A(_0503_),
    .B(_0530_),
    .Y(_0531_));
 sg13g2_or2_1 _4438_ (.X(_0532_),
    .B(_0530_),
    .A(_0503_));
 sg13g2_nor2_2 _4439_ (.A(net1218),
    .B(net1215),
    .Y(_0533_));
 sg13g2_nand2_2 _4440_ (.Y(_0534_),
    .A(net1289),
    .B(net1294));
 sg13g2_nor2_2 _4441_ (.A(_3046_),
    .B(_0533_),
    .Y(_0535_));
 sg13g2_nand2_2 _4442_ (.Y(_0536_),
    .A(_3047_),
    .B(_0534_));
 sg13g2_nor2_2 _4443_ (.A(_2904_),
    .B(_0535_),
    .Y(_0537_));
 sg13g2_o21ai_1 _4444_ (.B1(_0537_),
    .Y(_0538_),
    .A1(net1404),
    .A2(_3049_));
 sg13g2_nand2_1 _4445_ (.Y(_0539_),
    .A(_0452_),
    .B(_0538_));
 sg13g2_nor2_1 _4446_ (.A(_3188_),
    .B(_0535_),
    .Y(_0540_));
 sg13g2_nor2_1 _4447_ (.A(net1213),
    .B(net1299),
    .Y(_0541_));
 sg13g2_nand2_1 _4448_ (.Y(_0542_),
    .A(net1297),
    .B(net1212));
 sg13g2_xnor2_1 _4449_ (.Y(_0543_),
    .A(net1296),
    .B(net1300));
 sg13g2_inv_1 _4450_ (.Y(_0544_),
    .A(_0543_));
 sg13g2_a22oi_1 _4451_ (.Y(_0545_),
    .B1(_0543_),
    .B2(net1193),
    .A2(_0533_),
    .A1(net1297));
 sg13g2_nand2_1 _4452_ (.Y(_0546_),
    .A(net1219),
    .B(net1292));
 sg13g2_nand2_1 _4453_ (.Y(_0547_),
    .A(_0545_),
    .B(_0546_));
 sg13g2_nand3_1 _4454_ (.B(_0545_),
    .C(_0546_),
    .A(net1208),
    .Y(_0548_));
 sg13g2_nor2_1 _4455_ (.A(net1215),
    .B(net1299),
    .Y(_0549_));
 sg13g2_nand2_2 _4456_ (.Y(_0550_),
    .A(net1291),
    .B(net1212));
 sg13g2_nand3_1 _4457_ (.B(_0536_),
    .C(_0550_),
    .A(net1298),
    .Y(_0551_));
 sg13g2_a21oi_2 _4458_ (.B1(_0549_),
    .Y(_0552_),
    .A2(_0048_),
    .A1(net1300));
 sg13g2_nor2_1 _4459_ (.A(_0536_),
    .B(_0552_),
    .Y(_0553_));
 sg13g2_o21ai_1 _4460_ (.B1(_0551_),
    .Y(_0554_),
    .A1(_0536_),
    .A2(_0552_));
 sg13g2_o21ai_1 _4461_ (.B1(_0548_),
    .Y(_0555_),
    .A1(net1209),
    .A2(_0554_));
 sg13g2_nor2_1 _4462_ (.A(net1131),
    .B(_0555_),
    .Y(_0556_));
 sg13g2_a21oi_1 _4463_ (.A1(net1132),
    .A2(_0539_),
    .Y(_0557_),
    .B1(_0556_));
 sg13g2_xor2_1 _4464_ (.B(_0506_),
    .A(_0501_),
    .X(_0558_));
 sg13g2_a22oi_1 _4465_ (.Y(_0559_),
    .B1(_0540_),
    .B2(_0453_),
    .A2(_0535_),
    .A1(_3195_));
 sg13g2_o21ai_1 _4466_ (.B1(_3182_),
    .Y(_0560_),
    .A1(net1297),
    .A2(_2905_));
 sg13g2_nor2_1 _4467_ (.A(net1209),
    .B(_0560_),
    .Y(_0561_));
 sg13g2_a21oi_1 _4468_ (.A1(net1209),
    .A2(_0559_),
    .Y(_0562_),
    .B1(_0561_));
 sg13g2_nand2_1 _4469_ (.Y(_0563_),
    .A(_2904_),
    .B(net1187));
 sg13g2_nand2b_1 _4470_ (.Y(_0564_),
    .B(_0536_),
    .A_N(_0563_));
 sg13g2_nand2_1 _4471_ (.Y(_0565_),
    .A(net1213),
    .B(_0533_));
 sg13g2_o21ai_1 _4472_ (.B1(_0565_),
    .Y(_0566_),
    .A1(_0453_),
    .A2(_0536_));
 sg13g2_nand2_1 _4473_ (.Y(_0567_),
    .A(net1409),
    .B(_0566_));
 sg13g2_o21ai_1 _4474_ (.B1(_0567_),
    .Y(_0568_),
    .A1(net1409),
    .A2(_0564_));
 sg13g2_nor2_1 _4475_ (.A(net1131),
    .B(_0568_),
    .Y(_0569_));
 sg13g2_a21oi_1 _4476_ (.A1(net1131),
    .A2(_0562_),
    .Y(_0570_),
    .B1(_0569_));
 sg13g2_nand2_1 _4477_ (.Y(_0571_),
    .A(_0529_),
    .B(_0570_));
 sg13g2_a21oi_1 _4478_ (.A1(_0528_),
    .A2(_0557_),
    .Y(_0572_),
    .B1(_0558_));
 sg13g2_a21oi_2 _4479_ (.B1(_0451_),
    .Y(_0573_),
    .A2(_0563_),
    .A1(_0536_));
 sg13g2_or2_1 _4480_ (.X(_0574_),
    .B(_0553_),
    .A(_0537_));
 sg13g2_nor2_1 _4481_ (.A(net1408),
    .B(_0574_),
    .Y(_0575_));
 sg13g2_a22oi_1 _4482_ (.Y(_0576_),
    .B1(_3049_),
    .B2(_0537_),
    .A2(net1292),
    .A1(net1219));
 sg13g2_a21oi_1 _4483_ (.A1(net1410),
    .A2(_0576_),
    .Y(_0577_),
    .B1(_0575_));
 sg13g2_nand2_1 _4484_ (.Y(_0578_),
    .A(net1130),
    .B(_0577_));
 sg13g2_o21ai_1 _4485_ (.B1(_0578_),
    .Y(_0579_),
    .A1(net1130),
    .A2(_0573_));
 sg13g2_inv_1 _4486_ (.Y(_0580_),
    .A(_0579_));
 sg13g2_nor2_1 _4487_ (.A(_0528_),
    .B(_0579_),
    .Y(_0581_));
 sg13g2_and2_1 _4488_ (.A(_0546_),
    .B(_0551_),
    .X(_0582_));
 sg13g2_o21ai_1 _4489_ (.B1(_0545_),
    .Y(_0583_),
    .A1(_3194_),
    .A2(_0536_));
 sg13g2_nor2_1 _4490_ (.A(net1408),
    .B(_0582_),
    .Y(_0584_));
 sg13g2_a21oi_1 _4491_ (.A1(net1408),
    .A2(_0583_),
    .Y(_0585_),
    .B1(_0584_));
 sg13g2_a21oi_1 _4492_ (.A1(net1213),
    .A2(_0533_),
    .Y(_0586_),
    .B1(_3190_));
 sg13g2_nor2_1 _4493_ (.A(net1408),
    .B(_0586_),
    .Y(_0587_));
 sg13g2_nand2_2 _4494_ (.Y(_0588_),
    .A(_0453_),
    .B(_0563_));
 sg13g2_and2_1 _4495_ (.A(_0536_),
    .B(_0588_),
    .X(_0589_));
 sg13g2_a21oi_1 _4496_ (.A1(net1408),
    .A2(_0589_),
    .Y(_0590_),
    .B1(_0587_));
 sg13g2_nor2_1 _4497_ (.A(net1130),
    .B(_0585_),
    .Y(_0591_));
 sg13g2_a21oi_1 _4498_ (.A1(net1131),
    .A2(_0590_),
    .Y(_0592_),
    .B1(_0591_));
 sg13g2_a21oi_1 _4499_ (.A1(_0528_),
    .A2(_0592_),
    .Y(_0593_),
    .B1(_0581_));
 sg13g2_a22oi_1 _4500_ (.Y(_0594_),
    .B1(_0593_),
    .B2(_0558_),
    .A2(_0572_),
    .A1(_0571_));
 sg13g2_nand3_1 _4501_ (.B(_0527_),
    .C(_0594_),
    .A(\aliens_alive[12] ),
    .Y(_0595_));
 sg13g2_o21ai_1 _4502_ (.B1(net1241),
    .Y(_0596_),
    .A1(net1242),
    .A2(net1246));
 sg13g2_o21ai_1 _4503_ (.B1(net1235),
    .Y(_0597_),
    .A1(\group_x[6] ),
    .A2(_0596_));
 sg13g2_o21ai_1 _4504_ (.B1(net1233),
    .Y(_0598_),
    .A1(net1234),
    .A2(_0597_));
 sg13g2_nand2_1 _4505_ (.Y(_0599_),
    .A(net1228),
    .B(net1227));
 sg13g2_o21ai_1 _4506_ (.B1(_0598_),
    .Y(_0600_),
    .A1(_0597_),
    .A2(_0599_));
 sg13g2_inv_1 _4507_ (.Y(_0601_),
    .A(_0600_));
 sg13g2_xor2_1 _4508_ (.B(_0600_),
    .A(net1355),
    .X(_0602_));
 sg13g2_nand2_1 _4509_ (.Y(_0603_),
    .A(_0295_),
    .B(_0602_));
 sg13g2_xnor2_1 _4510_ (.Y(_0604_),
    .A(net1231),
    .B(_0598_));
 sg13g2_xor2_1 _4511_ (.B(_0604_),
    .A(_0008_),
    .X(_0605_));
 sg13g2_and2_2 _4512_ (.A(_0480_),
    .B(_0596_),
    .X(_0606_));
 sg13g2_inv_1 _4513_ (.Y(_0607_),
    .A(_0606_));
 sg13g2_nand2_1 _4514_ (.Y(_0608_),
    .A(_2825_),
    .B(net1385));
 sg13g2_xor2_1 _4515_ (.B(net1384),
    .A(net1248),
    .X(_0609_));
 sg13g2_nor2b_1 _4516_ (.A(net1391),
    .B_N(net1249),
    .Y(_0610_));
 sg13g2_nand2_1 _4517_ (.Y(_0611_),
    .A(_2826_),
    .B(net1392));
 sg13g2_a21oi_2 _4518_ (.B1(_0530_),
    .Y(_0612_),
    .A2(_0531_),
    .A1(net1410));
 sg13g2_o21ai_1 _4519_ (.B1(_0611_),
    .Y(_0613_),
    .A1(_0610_),
    .A2(_0612_));
 sg13g2_nor2_1 _4520_ (.A(_2825_),
    .B(net1199),
    .Y(_0614_));
 sg13g2_a21oi_2 _4521_ (.B1(_0614_),
    .Y(_0615_),
    .A2(_0613_),
    .A1(_0609_));
 sg13g2_xor2_1 _4522_ (.B(net1246),
    .A(net1242),
    .X(_0616_));
 sg13g2_xnor2_1 _4523_ (.Y(_0617_),
    .A(net1245),
    .B(net1247));
 sg13g2_xnor2_1 _4524_ (.Y(_0618_),
    .A(net1379),
    .B(_0616_));
 sg13g2_nand2b_1 _4525_ (.Y(_0619_),
    .B(_0618_),
    .A_N(_0615_));
 sg13g2_a22oi_1 _4526_ (.Y(_0620_),
    .B1(_0616_),
    .B2(net1382),
    .A2(_0607_),
    .A1(_2915_));
 sg13g2_a22oi_1 _4527_ (.Y(_0621_),
    .B1(_0619_),
    .B2(_0620_),
    .A2(_0606_),
    .A1(net1374));
 sg13g2_xnor2_1 _4528_ (.Y(_0622_),
    .A(net1237),
    .B(_0596_));
 sg13g2_inv_1 _4529_ (.Y(_0623_),
    .A(_0622_));
 sg13g2_xor2_1 _4530_ (.B(_0622_),
    .A(net1366),
    .X(_0624_));
 sg13g2_nand2_1 _4531_ (.Y(_0625_),
    .A(_0621_),
    .B(_0624_));
 sg13g2_nor2_2 _4532_ (.A(net1194),
    .B(net1367),
    .Y(_0626_));
 sg13g2_nand2b_1 _4533_ (.Y(_0627_),
    .B(_0624_),
    .A_N(_0626_));
 sg13g2_xnor2_1 _4534_ (.Y(_0628_),
    .A(_0061_),
    .B(_0597_));
 sg13g2_xnor2_1 _4535_ (.Y(_0629_),
    .A(net1361),
    .B(_0628_));
 sg13g2_a22oi_1 _4536_ (.Y(_0630_),
    .B1(_0629_),
    .B2(_0627_),
    .A2(_0628_),
    .A1(net1364));
 sg13g2_xor2_1 _4537_ (.B(_0630_),
    .A(_0602_),
    .X(_0631_));
 sg13g2_xnor2_1 _4538_ (.Y(_0632_),
    .A(_0627_),
    .B(_0629_));
 sg13g2_xnor2_1 _4539_ (.Y(_0633_),
    .A(net1374),
    .B(_0606_));
 sg13g2_a21oi_1 _4540_ (.A1(net1382),
    .A2(_0616_),
    .Y(_0634_),
    .B1(_0618_));
 sg13g2_xnor2_1 _4541_ (.Y(_0635_),
    .A(_0633_),
    .B(_0634_));
 sg13g2_xor2_1 _4542_ (.B(_0618_),
    .A(_0615_),
    .X(_0636_));
 sg13g2_xnor2_1 _4543_ (.Y(_0637_),
    .A(_0603_),
    .B(_0605_));
 sg13g2_nand4_1 _4544_ (.B(_0635_),
    .C(_0636_),
    .A(_0625_),
    .Y(_0638_),
    .D(_0637_));
 sg13g2_o21ai_1 _4545_ (.B1(_0632_),
    .Y(_0639_),
    .A1(_0621_),
    .A2(_0624_));
 sg13g2_nor3_2 _4546_ (.A(_0631_),
    .B(_0638_),
    .C(_0639_),
    .Y(_0640_));
 sg13g2_xnor2_1 _4547_ (.Y(_0641_),
    .A(_0505_),
    .B(_0612_));
 sg13g2_xor2_1 _4548_ (.B(_0612_),
    .A(_0505_),
    .X(_0642_));
 sg13g2_xnor2_1 _4549_ (.Y(_0643_),
    .A(net1410),
    .B(_0531_));
 sg13g2_nand2_1 _4550_ (.Y(_0644_),
    .A(net1209),
    .B(_0566_));
 sg13g2_o21ai_1 _4551_ (.B1(_0644_),
    .Y(_0645_),
    .A1(net1209),
    .A2(_0564_));
 sg13g2_nor2_1 _4552_ (.A(net1409),
    .B(_0560_),
    .Y(_0646_));
 sg13g2_a21oi_1 _4553_ (.A1(net1408),
    .A2(_0559_),
    .Y(_0647_),
    .B1(_0646_));
 sg13g2_nand2_1 _4554_ (.Y(_0648_),
    .A(net1110),
    .B(_0645_));
 sg13g2_o21ai_1 _4555_ (.B1(_0648_),
    .Y(_0649_),
    .A1(net1110),
    .A2(_0647_));
 sg13g2_xor2_1 _4556_ (.B(_0613_),
    .A(_0609_),
    .X(_0650_));
 sg13g2_xnor2_1 _4557_ (.Y(_0651_),
    .A(_0609_),
    .B(_0613_));
 sg13g2_mux2_1 _4558_ (.A0(_0547_),
    .A1(_0554_),
    .S(net1209),
    .X(_0652_));
 sg13g2_nand2_1 _4559_ (.Y(_0653_),
    .A(net1404),
    .B(_3048_));
 sg13g2_a21oi_2 _4560_ (.B1(_0451_),
    .Y(_0654_),
    .A2(_0653_),
    .A1(_0537_));
 sg13g2_nor2_1 _4561_ (.A(net1110),
    .B(_0654_),
    .Y(_0655_));
 sg13g2_a21oi_1 _4562_ (.A1(net1110),
    .A2(_0652_),
    .Y(_0656_),
    .B1(_0655_));
 sg13g2_nand2_1 _4563_ (.Y(_0657_),
    .A(net1086),
    .B(_0656_));
 sg13g2_a21oi_1 _4564_ (.A1(net1087),
    .A2(_0649_),
    .Y(_0658_),
    .B1(_0650_));
 sg13g2_nor2_1 _4565_ (.A(net1209),
    .B(_0574_),
    .Y(_0659_));
 sg13g2_a21oi_1 _4566_ (.A1(net1210),
    .A2(_0576_),
    .Y(_0660_),
    .B1(_0659_));
 sg13g2_nand2_1 _4567_ (.Y(_0661_),
    .A(_0573_),
    .B(net1111));
 sg13g2_o21ai_1 _4568_ (.B1(_0661_),
    .Y(_0662_),
    .A1(net1111),
    .A2(_0660_));
 sg13g2_nand2_1 _4569_ (.Y(_0663_),
    .A(_0641_),
    .B(_0662_));
 sg13g2_nand2_1 _4570_ (.Y(_0664_),
    .A(net1408),
    .B(_0582_));
 sg13g2_o21ai_1 _4571_ (.B1(_0664_),
    .Y(_0665_),
    .A1(net1408),
    .A2(_0583_));
 sg13g2_nand2_1 _4572_ (.Y(_0666_),
    .A(net1209),
    .B(_0589_));
 sg13g2_o21ai_1 _4573_ (.B1(_0666_),
    .Y(_0667_),
    .A1(net1210),
    .A2(_0586_));
 sg13g2_mux2_1 _4574_ (.A0(_0667_),
    .A1(_0665_),
    .S(net1110),
    .X(_0668_));
 sg13g2_a21oi_1 _4575_ (.A1(net1086),
    .A2(_0668_),
    .Y(_0669_),
    .B1(_0651_));
 sg13g2_a22oi_1 _4576_ (.Y(_0670_),
    .B1(_0663_),
    .B2(_0669_),
    .A2(_0658_),
    .A1(_0657_));
 sg13g2_nand3_1 _4577_ (.B(_0640_),
    .C(_0670_),
    .A(\aliens_alive[15] ),
    .Y(_0671_));
 sg13g2_nand2b_1 _4578_ (.Y(_0672_),
    .B(net1239),
    .A_N(_0482_));
 sg13g2_and2_1 _4579_ (.A(_2823_),
    .B(_0672_),
    .X(_0673_));
 sg13g2_nor2_1 _4580_ (.A(_0485_),
    .B(_0673_),
    .Y(_0674_));
 sg13g2_o21ai_1 _4581_ (.B1(_2821_),
    .Y(_0675_),
    .A1(net1226),
    .A2(_0673_));
 sg13g2_nand2b_2 _4582_ (.Y(_0676_),
    .B(_0675_),
    .A_N(_0674_));
 sg13g2_xor2_1 _4583_ (.B(_0676_),
    .A(net1355),
    .X(_0677_));
 sg13g2_xnor2_1 _4584_ (.Y(_0678_),
    .A(net1226),
    .B(_0673_));
 sg13g2_xor2_1 _4585_ (.B(_0678_),
    .A(net1361),
    .X(_0679_));
 sg13g2_xnor2_1 _4586_ (.Y(_0680_),
    .A(net1241),
    .B(_0482_));
 sg13g2_inv_1 _4587_ (.Y(_0681_),
    .A(_0680_));
 sg13g2_o21ai_1 _4588_ (.B1(_0502_),
    .Y(_0682_),
    .A1(_0504_),
    .A2(_0612_));
 sg13g2_a22oi_1 _4589_ (.Y(_0683_),
    .B1(_0501_),
    .B2(_0682_),
    .A2(_0499_),
    .A1(net1385));
 sg13g2_nor2_1 _4590_ (.A(_0498_),
    .B(_0683_),
    .Y(_0684_));
 sg13g2_a221oi_1 _4591_ (.B2(_2915_),
    .C1(_0684_),
    .B1(_0681_),
    .A1(net1382),
    .Y(_0685_),
    .A2(_0496_));
 sg13g2_a21oi_1 _4592_ (.A1(net1373),
    .A2(_0680_),
    .Y(_0686_),
    .B1(_0685_));
 sg13g2_xor2_1 _4593_ (.B(_0672_),
    .A(net1236),
    .X(_0687_));
 sg13g2_xnor2_1 _4594_ (.Y(_0688_),
    .A(net1367),
    .B(_0687_));
 sg13g2_a22oi_1 _4595_ (.Y(_0689_),
    .B1(_0688_),
    .B2(_0686_),
    .A2(_0687_),
    .A1(net1371));
 sg13g2_nand2_1 _4596_ (.Y(_0690_),
    .A(net1364),
    .B(_0678_));
 sg13g2_o21ai_1 _4597_ (.B1(_0690_),
    .Y(_0691_),
    .A1(_0679_),
    .A2(_0689_));
 sg13g2_xor2_1 _4598_ (.B(_0688_),
    .A(_0686_),
    .X(_0692_));
 sg13g2_xor2_1 _4599_ (.B(_0674_),
    .A(_0078_),
    .X(_0693_));
 sg13g2_xnor2_1 _4600_ (.Y(_0694_),
    .A(_0008_),
    .B(_0693_));
 sg13g2_a21oi_1 _4601_ (.A1(_0295_),
    .A2(_0677_),
    .Y(_0695_),
    .B1(_0694_));
 sg13g2_xnor2_1 _4602_ (.Y(_0696_),
    .A(_0498_),
    .B(_0683_));
 sg13g2_xnor2_1 _4603_ (.Y(_0697_),
    .A(_2915_),
    .B(_0680_));
 sg13g2_nand2_1 _4604_ (.Y(_0698_),
    .A(_0497_),
    .B(_0498_));
 sg13g2_xnor2_1 _4605_ (.Y(_0699_),
    .A(_0697_),
    .B(_0698_));
 sg13g2_nor2_1 _4606_ (.A(_0626_),
    .B(_0688_),
    .Y(_0700_));
 sg13g2_xnor2_1 _4607_ (.Y(_0701_),
    .A(_0679_),
    .B(_0700_));
 sg13g2_nand3_1 _4608_ (.B(_0677_),
    .C(_0694_),
    .A(_0295_),
    .Y(_0702_));
 sg13g2_nand4_1 _4609_ (.B(_0699_),
    .C(_0701_),
    .A(_0696_),
    .Y(_0703_),
    .D(_0702_));
 sg13g2_xnor2_1 _4610_ (.Y(_0704_),
    .A(_0677_),
    .B(_0691_));
 sg13g2_nor4_2 _4611_ (.A(_0692_),
    .B(_0695_),
    .C(_0703_),
    .Y(_0705_),
    .D(_0704_));
 sg13g2_xor2_1 _4612_ (.B(_0682_),
    .A(_0501_),
    .X(_0706_));
 sg13g2_nand2_1 _4613_ (.Y(_0707_),
    .A(net1086),
    .B(_0649_));
 sg13g2_a21oi_1 _4614_ (.A1(_0641_),
    .A2(_0656_),
    .Y(_0708_),
    .B1(_0706_));
 sg13g2_and2_1 _4615_ (.A(_0641_),
    .B(_0668_),
    .X(_0709_));
 sg13g2_a21oi_1 _4616_ (.A1(net1086),
    .A2(_0662_),
    .Y(_0710_),
    .B1(_0709_));
 sg13g2_a22oi_1 _4617_ (.Y(_0711_),
    .B1(_0710_),
    .B2(_0706_),
    .A2(_0708_),
    .A1(_0707_));
 sg13g2_nand3_1 _4618_ (.B(_0705_),
    .C(_0711_),
    .A(\aliens_alive[11] ),
    .Y(_0712_));
 sg13g2_nand3_1 _4619_ (.B(_0671_),
    .C(_0712_),
    .A(_0595_),
    .Y(_0713_));
 sg13g2_nand2_1 _4620_ (.Y(_0714_),
    .A(net1228),
    .B(net1359));
 sg13g2_xnor2_1 _4621_ (.Y(_0715_),
    .A(net1233),
    .B(net1359));
 sg13g2_xnor2_1 _4622_ (.Y(_0716_),
    .A(net1234),
    .B(net1364));
 sg13g2_xnor2_1 _4623_ (.Y(_0717_),
    .A(net1238),
    .B(net1371));
 sg13g2_xor2_1 _4624_ (.B(net1377),
    .A(net1239),
    .X(_0718_));
 sg13g2_nor2_1 _4625_ (.A(net1245),
    .B(net1197),
    .Y(_0719_));
 sg13g2_nand2_1 _4626_ (.Y(_0720_),
    .A(net1245),
    .B(net1197));
 sg13g2_nand2b_1 _4627_ (.Y(_0721_),
    .B(_0720_),
    .A_N(_0719_));
 sg13g2_nor2_1 _4628_ (.A(_0503_),
    .B(_0610_),
    .Y(_0722_));
 sg13g2_a21oi_2 _4629_ (.B1(_0722_),
    .Y(_0723_),
    .A2(net1391),
    .A1(_2826_));
 sg13g2_o21ai_1 _4630_ (.B1(_0608_),
    .Y(_0724_),
    .A1(_0609_),
    .A2(_0723_));
 sg13g2_a21oi_1 _4631_ (.A1(_0720_),
    .A2(_0724_),
    .Y(_0725_),
    .B1(_0719_));
 sg13g2_nor2_1 _4632_ (.A(_0718_),
    .B(_0725_),
    .Y(_0726_));
 sg13g2_a21oi_1 _4633_ (.A1(_2824_),
    .A2(net1377),
    .Y(_0727_),
    .B1(_0726_));
 sg13g2_nor2b_1 _4634_ (.A(_0727_),
    .B_N(_0717_),
    .Y(_0728_));
 sg13g2_a21oi_1 _4635_ (.A1(_2823_),
    .A2(net1371),
    .Y(_0729_),
    .B1(_0728_));
 sg13g2_nor2b_1 _4636_ (.A(_0729_),
    .B_N(_0716_),
    .Y(_0730_));
 sg13g2_a21oi_1 _4637_ (.A1(net1227),
    .A2(net1364),
    .Y(_0731_),
    .B1(_0730_));
 sg13g2_nand2b_1 _4638_ (.Y(_0732_),
    .B(_0715_),
    .A_N(_0731_));
 sg13g2_xnor2_1 _4639_ (.Y(_0733_),
    .A(net1231),
    .B(net1354));
 sg13g2_a21oi_1 _4640_ (.A1(_0714_),
    .A2(_0732_),
    .Y(_0734_),
    .B1(_0733_));
 sg13g2_and3_1 _4641_ (.X(_0735_),
    .A(_0714_),
    .B(_0732_),
    .C(_0733_));
 sg13g2_xor2_1 _4642_ (.B(_0731_),
    .A(_0715_),
    .X(_0736_));
 sg13g2_xor2_1 _4643_ (.B(_0729_),
    .A(_0716_),
    .X(_0737_));
 sg13g2_xor2_1 _4644_ (.B(_0727_),
    .A(_0717_),
    .X(_0738_));
 sg13g2_xnor2_1 _4645_ (.Y(_0739_),
    .A(_0721_),
    .B(_0724_));
 sg13g2_xnor2_1 _4646_ (.Y(_0740_),
    .A(_0718_),
    .B(_0725_));
 sg13g2_nand4_1 _4647_ (.B(_0737_),
    .C(_0738_),
    .A(_0736_),
    .Y(_0741_),
    .D(_0740_));
 sg13g2_nor4_2 _4648_ (.A(_0734_),
    .B(_0735_),
    .C(_0739_),
    .Y(_0742_),
    .D(_0741_));
 sg13g2_xnor2_1 _4649_ (.Y(_0743_),
    .A(_0609_),
    .B(_0723_));
 sg13g2_mux4_1 _4650_ (.S0(_0529_),
    .A0(_0580_),
    .A1(_0592_),
    .A2(_0570_),
    .A3(_0557_),
    .S1(_0743_),
    .X(_0744_));
 sg13g2_nand2_1 _4651_ (.Y(_0745_),
    .A(_0742_),
    .B(_0744_));
 sg13g2_nor2_1 _4652_ (.A(net1250),
    .B(net1253),
    .Y(_0746_));
 sg13g2_nor3_2 _4653_ (.A(net1247),
    .B(net1250),
    .C(net1253),
    .Y(_0747_));
 sg13g2_nor2b_1 _4654_ (.A(net1242),
    .B_N(_0747_),
    .Y(_0748_));
 sg13g2_nor2_2 _4655_ (.A(_2824_),
    .B(_0748_),
    .Y(_0749_));
 sg13g2_nand2_2 _4656_ (.Y(_0750_),
    .A(\group_x[6] ),
    .B(_0749_));
 sg13g2_nor2_1 _4657_ (.A(_0061_),
    .B(_0750_),
    .Y(_0751_));
 sg13g2_xnor2_1 _4658_ (.Y(_0752_),
    .A(_0074_),
    .B(_0751_));
 sg13g2_xor2_1 _4659_ (.B(_0752_),
    .A(net1355),
    .X(_0753_));
 sg13g2_xnor2_1 _4660_ (.Y(_0754_),
    .A(_0061_),
    .B(_0750_));
 sg13g2_xor2_1 _4661_ (.B(_0754_),
    .A(net1361),
    .X(_0755_));
 sg13g2_nand2b_2 _4662_ (.Y(_0756_),
    .B(_0747_),
    .A_N(_0479_));
 sg13g2_nor2b_2 _4663_ (.A(_0749_),
    .B_N(_0756_),
    .Y(_0757_));
 sg13g2_nand2_1 _4664_ (.Y(_0758_),
    .A(net1373),
    .B(_0757_));
 sg13g2_xnor2_1 _4665_ (.Y(_0759_),
    .A(_2896_),
    .B(_0747_));
 sg13g2_xnor2_1 _4666_ (.Y(_0760_),
    .A(_0076_),
    .B(_0747_));
 sg13g2_xnor2_1 _4667_ (.Y(_0761_),
    .A(net1378),
    .B(_0759_));
 sg13g2_xor2_1 _4668_ (.B(_0746_),
    .A(_0070_),
    .X(_0762_));
 sg13g2_nand2_1 _4669_ (.Y(_0763_),
    .A(net1385),
    .B(_0762_));
 sg13g2_xor2_1 _4670_ (.B(_0762_),
    .A(_0033_),
    .X(_0764_));
 sg13g2_nand2_2 _4671_ (.Y(_0765_),
    .A(net1250),
    .B(net1253));
 sg13g2_xor2_1 _4672_ (.B(net1252),
    .A(net1249),
    .X(_0766_));
 sg13g2_inv_2 _4673_ (.Y(_0767_),
    .A(net1186));
 sg13g2_nand2_1 _4674_ (.Y(_0768_),
    .A(net1391),
    .B(net1186));
 sg13g2_xnor2_1 _4675_ (.Y(_0769_),
    .A(_0042_),
    .B(net1186));
 sg13g2_a21oi_2 _4676_ (.B1(net1191),
    .Y(_0770_),
    .A2(_3066_),
    .A1(_2827_));
 sg13g2_a22oi_1 _4677_ (.Y(_0771_),
    .B1(_0769_),
    .B2(_0770_),
    .A2(net1186),
    .A1(net1391));
 sg13g2_o21ai_1 _4678_ (.B1(_0763_),
    .Y(_0772_),
    .A1(_0764_),
    .A2(_0771_));
 sg13g2_nand2_1 _4679_ (.Y(_0773_),
    .A(_0761_),
    .B(_0772_));
 sg13g2_nand2_1 _4680_ (.Y(_0774_),
    .A(net1382),
    .B(_0759_));
 sg13g2_or2_1 _4681_ (.X(_0775_),
    .B(_0757_),
    .A(net1373));
 sg13g2_nand3_1 _4682_ (.B(_0774_),
    .C(_0775_),
    .A(_0773_),
    .Y(_0776_));
 sg13g2_xor2_1 _4683_ (.B(_0749_),
    .A(net1235),
    .X(_0777_));
 sg13g2_xnor2_1 _4684_ (.Y(_0778_),
    .A(net1366),
    .B(_0777_));
 sg13g2_nand3_1 _4685_ (.B(_0776_),
    .C(_0778_),
    .A(_0758_),
    .Y(_0779_));
 sg13g2_nand2_1 _4686_ (.Y(_0780_),
    .A(net1371),
    .B(_0777_));
 sg13g2_a21oi_1 _4687_ (.A1(_0779_),
    .A2(_0780_),
    .Y(_0781_),
    .B1(_0755_));
 sg13g2_a21oi_1 _4688_ (.A1(net1364),
    .A2(_0754_),
    .Y(_0782_),
    .B1(_0781_));
 sg13g2_a21o_1 _4689_ (.A2(_0776_),
    .A1(_0758_),
    .B1(_0778_),
    .X(_0783_));
 sg13g2_nor2_1 _4690_ (.A(_0294_),
    .B(_0753_),
    .Y(_0784_));
 sg13g2_or2_1 _4691_ (.X(_0785_),
    .B(_0750_),
    .A(_0485_));
 sg13g2_xor2_1 _4692_ (.B(_0785_),
    .A(_0078_),
    .X(_0786_));
 sg13g2_xnor2_1 _4693_ (.Y(_0787_),
    .A(net1352),
    .B(_0786_));
 sg13g2_nor2_1 _4694_ (.A(_0626_),
    .B(_0778_),
    .Y(_0788_));
 sg13g2_xnor2_1 _4695_ (.Y(_0789_),
    .A(_0755_),
    .B(_0788_));
 sg13g2_xnor2_1 _4696_ (.Y(_0790_),
    .A(_0761_),
    .B(_0772_));
 sg13g2_nand2_1 _4697_ (.Y(_0791_),
    .A(_0758_),
    .B(_0775_));
 sg13g2_nor2b_1 _4698_ (.A(_0761_),
    .B_N(_0774_),
    .Y(_0792_));
 sg13g2_xnor2_1 _4699_ (.Y(_0793_),
    .A(_0791_),
    .B(_0792_));
 sg13g2_xnor2_1 _4700_ (.Y(_0794_),
    .A(_0784_),
    .B(_0787_));
 sg13g2_nand4_1 _4701_ (.B(_0790_),
    .C(_0793_),
    .A(_0789_),
    .Y(_0795_),
    .D(_0794_));
 sg13g2_nand2b_1 _4702_ (.Y(_0796_),
    .B(_0782_),
    .A_N(_0753_));
 sg13g2_nand2b_1 _4703_ (.Y(_0797_),
    .B(_0753_),
    .A_N(_0782_));
 sg13g2_a221oi_1 _4704_ (.B2(_0797_),
    .C1(_0795_),
    .B1(_0796_),
    .A1(_0779_),
    .Y(_0798_),
    .A2(_0783_));
 sg13g2_nand2b_1 _4705_ (.Y(_0799_),
    .B(_0770_),
    .A_N(_0769_));
 sg13g2_xor2_1 _4706_ (.B(_0770_),
    .A(_0769_),
    .X(_0800_));
 sg13g2_xnor2_1 _4707_ (.Y(_0801_),
    .A(_0769_),
    .B(_0770_));
 sg13g2_nand2_1 _4708_ (.Y(_0802_),
    .A(net1110),
    .B(_0654_));
 sg13g2_o21ai_1 _4709_ (.B1(_0802_),
    .Y(_0803_),
    .A1(net1113),
    .A2(_0652_));
 sg13g2_xor2_1 _4710_ (.B(_0771_),
    .A(_0764_),
    .X(_0804_));
 sg13g2_nor2_1 _4711_ (.A(net1110),
    .B(_0645_),
    .Y(_0805_));
 sg13g2_a21oi_1 _4712_ (.A1(net1113),
    .A2(_0647_),
    .Y(_0806_),
    .B1(_0805_));
 sg13g2_nand2_1 _4713_ (.Y(_0807_),
    .A(_0801_),
    .B(_0806_));
 sg13g2_a21oi_1 _4714_ (.A1(net1122),
    .A2(_0803_),
    .Y(_0808_),
    .B1(_0804_));
 sg13g2_mux2_1 _4715_ (.A0(_0665_),
    .A1(_0667_),
    .S(net1110),
    .X(_0809_));
 sg13g2_and2_1 _4716_ (.A(net1122),
    .B(_0809_),
    .X(_0810_));
 sg13g2_nor2_1 _4717_ (.A(_0573_),
    .B(net1111),
    .Y(_0811_));
 sg13g2_a21oi_1 _4718_ (.A1(net1111),
    .A2(_0660_),
    .Y(_0812_),
    .B1(_0811_));
 sg13g2_a21oi_1 _4719_ (.A1(_0801_),
    .A2(_0812_),
    .Y(_0813_),
    .B1(_0810_));
 sg13g2_a22oi_1 _4720_ (.Y(_0814_),
    .B1(_0813_),
    .B2(_0804_),
    .A2(_0808_),
    .A1(_0807_));
 sg13g2_nand3_1 _4721_ (.B(_0798_),
    .C(_0814_),
    .A(\aliens_alive[9] ),
    .Y(_0815_));
 sg13g2_o21ai_1 _4722_ (.B1(_0815_),
    .Y(_0816_),
    .A1(_0006_),
    .A2(_0745_));
 sg13g2_nand3b_1 _4723_ (.B(_2825_),
    .C(_0765_),
    .Y(_0817_),
    .A_N(net1245));
 sg13g2_nand2_1 _4724_ (.Y(_0818_),
    .A(net1239),
    .B(_0817_));
 sg13g2_nand3_1 _4725_ (.B(net1239),
    .C(_0817_),
    .A(net1237),
    .Y(_0819_));
 sg13g2_nand2_1 _4726_ (.Y(_0820_),
    .A(_0061_),
    .B(_0819_));
 sg13g2_xnor2_1 _4727_ (.Y(_0821_),
    .A(_2821_),
    .B(_0820_));
 sg13g2_xnor2_1 _4728_ (.Y(_0822_),
    .A(net1355),
    .B(_0821_));
 sg13g2_xnor2_1 _4729_ (.Y(_0823_),
    .A(net1226),
    .B(_0819_));
 sg13g2_inv_1 _4730_ (.Y(_0824_),
    .A(_0823_));
 sg13g2_xor2_1 _4731_ (.B(_0823_),
    .A(net1361),
    .X(_0825_));
 sg13g2_nand2b_1 _4732_ (.Y(_0826_),
    .B(_0765_),
    .A_N(_0480_));
 sg13g2_and2_2 _4733_ (.A(_0818_),
    .B(_0826_),
    .X(_0827_));
 sg13g2_nor2_1 _4734_ (.A(net1373),
    .B(_0827_),
    .Y(_0828_));
 sg13g2_nand2_1 _4735_ (.Y(_0829_),
    .A(net1373),
    .B(_0827_));
 sg13g2_nand2_1 _4736_ (.Y(_0830_),
    .A(_0070_),
    .B(_0765_));
 sg13g2_xnor2_1 _4737_ (.Y(_0831_),
    .A(_2896_),
    .B(_0830_));
 sg13g2_xnor2_1 _4738_ (.Y(_0832_),
    .A(_0076_),
    .B(_0830_));
 sg13g2_nand2_1 _4739_ (.Y(_0833_),
    .A(net1382),
    .B(_0832_));
 sg13g2_xnor2_1 _4740_ (.Y(_0834_),
    .A(net1378),
    .B(net1119));
 sg13g2_xnor2_1 _4741_ (.Y(_0835_),
    .A(net1247),
    .B(_0765_));
 sg13g2_inv_1 _4742_ (.Y(_0836_),
    .A(_0835_));
 sg13g2_xnor2_1 _4743_ (.Y(_0837_),
    .A(_0033_),
    .B(_0835_));
 sg13g2_nand2_1 _4744_ (.Y(_0838_),
    .A(net1391),
    .B(_0767_));
 sg13g2_nand2_1 _4745_ (.Y(_0839_),
    .A(_0799_),
    .B(_0838_));
 sg13g2_a22oi_1 _4746_ (.Y(_0840_),
    .B1(_0837_),
    .B2(_0839_),
    .A2(_0835_),
    .A1(net1385));
 sg13g2_o21ai_1 _4747_ (.B1(_0833_),
    .Y(_0841_),
    .A1(_0834_),
    .A2(_0840_));
 sg13g2_a21oi_1 _4748_ (.A1(_0829_),
    .A2(_0841_),
    .Y(_0842_),
    .B1(_0828_));
 sg13g2_xor2_1 _4749_ (.B(_0818_),
    .A(net1236),
    .X(_0843_));
 sg13g2_xor2_1 _4750_ (.B(_0843_),
    .A(net1367),
    .X(_0844_));
 sg13g2_nand2b_1 _4751_ (.Y(_0845_),
    .B(_0844_),
    .A_N(_0842_));
 sg13g2_o21ai_1 _4752_ (.B1(_0845_),
    .Y(_0846_),
    .A1(net1194),
    .A2(_0843_));
 sg13g2_a22oi_1 _4753_ (.Y(_0847_),
    .B1(_0825_),
    .B2(_0846_),
    .A2(_0824_),
    .A1(net1365));
 sg13g2_xor2_1 _4754_ (.B(_0847_),
    .A(_0822_),
    .X(_0848_));
 sg13g2_xnor2_1 _4755_ (.Y(_0849_),
    .A(_0842_),
    .B(_0844_));
 sg13g2_a21o_1 _4756_ (.A2(_0819_),
    .A1(net1226),
    .B1(net1228),
    .X(_0850_));
 sg13g2_xnor2_1 _4757_ (.Y(_0851_),
    .A(_2820_),
    .B(_0850_));
 sg13g2_xnor2_1 _4758_ (.Y(_0852_),
    .A(net1232),
    .B(_0850_));
 sg13g2_xnor2_1 _4759_ (.Y(_0853_),
    .A(net1352),
    .B(_0851_));
 sg13g2_a21oi_1 _4760_ (.A1(_0295_),
    .A2(_0822_),
    .Y(_0854_),
    .B1(_0853_));
 sg13g2_nor2_1 _4761_ (.A(_0626_),
    .B(_0844_),
    .Y(_0855_));
 sg13g2_xor2_1 _4762_ (.B(_0855_),
    .A(_0825_),
    .X(_0856_));
 sg13g2_xnor2_1 _4763_ (.Y(_0857_),
    .A(_0834_),
    .B(_0840_));
 sg13g2_xnor2_1 _4764_ (.Y(_0858_),
    .A(_2915_),
    .B(_0827_));
 sg13g2_nand2_1 _4765_ (.Y(_0859_),
    .A(_0833_),
    .B(_0834_));
 sg13g2_xnor2_1 _4766_ (.Y(_0860_),
    .A(_0858_),
    .B(_0859_));
 sg13g2_nand3_1 _4767_ (.B(_0822_),
    .C(_0853_),
    .A(_0295_),
    .Y(_0861_));
 sg13g2_nand4_1 _4768_ (.B(_0857_),
    .C(_0860_),
    .A(_0856_),
    .Y(_0862_),
    .D(_0861_));
 sg13g2_nor4_2 _4769_ (.A(_0848_),
    .B(_0849_),
    .C(_0854_),
    .Y(_0863_),
    .D(_0862_));
 sg13g2_xor2_1 _4770_ (.B(_0839_),
    .A(_0837_),
    .X(_0864_));
 sg13g2_mux4_1 _4771_ (.S0(net1122),
    .A0(_0803_),
    .A1(_0806_),
    .A2(_0809_),
    .A3(_0812_),
    .S1(_0864_),
    .X(_0865_));
 sg13g2_nand3_1 _4772_ (.B(_0863_),
    .C(_0865_),
    .A(\aliens_alive[13] ),
    .Y(_0866_));
 sg13g2_and2_1 _4773_ (.A(net1237),
    .B(_0826_),
    .X(_0867_));
 sg13g2_xnor2_1 _4774_ (.Y(_0868_),
    .A(_0061_),
    .B(_0867_));
 sg13g2_nand2_1 _4775_ (.Y(_0869_),
    .A(net1364),
    .B(_0868_));
 sg13g2_xnor2_1 _4776_ (.Y(_0870_),
    .A(_2823_),
    .B(_0826_));
 sg13g2_nor2_1 _4777_ (.A(net1367),
    .B(_0870_),
    .Y(_0871_));
 sg13g2_nand2_1 _4778_ (.Y(_0872_),
    .A(net1366),
    .B(_0870_));
 sg13g2_nand2b_1 _4779_ (.Y(_0873_),
    .B(_0872_),
    .A_N(_0871_));
 sg13g2_xor2_1 _4780_ (.B(_0817_),
    .A(_0075_),
    .X(_0874_));
 sg13g2_nor2_2 _4781_ (.A(net1252),
    .B(net1396),
    .Y(_0875_));
 sg13g2_o21ai_1 _4782_ (.B1(_0838_),
    .Y(_0876_),
    .A1(_0769_),
    .A2(_0875_));
 sg13g2_a22oi_1 _4783_ (.Y(_0877_),
    .B1(_0837_),
    .B2(_0876_),
    .A2(_0835_),
    .A1(net1384));
 sg13g2_o21ai_1 _4784_ (.B1(_0833_),
    .Y(_0878_),
    .A1(_0834_),
    .A2(_0877_));
 sg13g2_xnor2_1 _4785_ (.Y(_0879_),
    .A(net1373),
    .B(_0874_));
 sg13g2_nand2b_1 _4786_ (.Y(_0880_),
    .B(_0878_),
    .A_N(_0879_));
 sg13g2_o21ai_1 _4787_ (.B1(_0880_),
    .Y(_0881_),
    .A1(net1195),
    .A2(_0874_));
 sg13g2_a21oi_1 _4788_ (.A1(_0872_),
    .A2(_0881_),
    .Y(_0882_),
    .B1(_0871_));
 sg13g2_xor2_1 _4789_ (.B(_0868_),
    .A(net1361),
    .X(_0883_));
 sg13g2_o21ai_1 _4790_ (.B1(_0869_),
    .Y(_0884_),
    .A1(_0882_),
    .A2(_0883_));
 sg13g2_nor2_2 _4791_ (.A(\group_x[7] ),
    .B(_0867_),
    .Y(_0885_));
 sg13g2_nor2_1 _4792_ (.A(net1228),
    .B(_0885_),
    .Y(_0886_));
 sg13g2_xnor2_1 _4793_ (.Y(_0887_),
    .A(net1233),
    .B(_0885_));
 sg13g2_xnor2_1 _4794_ (.Y(_0888_),
    .A(net1228),
    .B(_0885_));
 sg13g2_xnor2_1 _4795_ (.Y(_0889_),
    .A(net1355),
    .B(_0887_));
 sg13g2_xor2_1 _4796_ (.B(_0883_),
    .A(_0882_),
    .X(_0890_));
 sg13g2_xnor2_1 _4797_ (.Y(_0891_),
    .A(_0873_),
    .B(_0881_));
 sg13g2_xor2_1 _4798_ (.B(_0879_),
    .A(_0878_),
    .X(_0892_));
 sg13g2_nand2_1 _4799_ (.Y(_0893_),
    .A(_0295_),
    .B(_0889_));
 sg13g2_xnor2_1 _4800_ (.Y(_0894_),
    .A(net1232),
    .B(_0886_));
 sg13g2_xnor2_1 _4801_ (.Y(_0895_),
    .A(net1352),
    .B(_0894_));
 sg13g2_xnor2_1 _4802_ (.Y(_0896_),
    .A(_0834_),
    .B(_0877_));
 sg13g2_xnor2_1 _4803_ (.Y(_0897_),
    .A(_0893_),
    .B(_0895_));
 sg13g2_nand3_1 _4804_ (.B(_0896_),
    .C(_0897_),
    .A(_0892_),
    .Y(_0898_));
 sg13g2_nor3_1 _4805_ (.A(_0890_),
    .B(_0891_),
    .C(_0898_),
    .Y(_0899_));
 sg13g2_o21ai_1 _4806_ (.B1(_0899_),
    .Y(_0900_),
    .A1(_0884_),
    .A2(_0889_));
 sg13g2_a21oi_2 _4807_ (.B1(_0900_),
    .Y(_0901_),
    .A2(_0889_),
    .A1(_0884_));
 sg13g2_nand2b_1 _4808_ (.Y(_0902_),
    .B(_0769_),
    .A_N(_0875_));
 sg13g2_xnor2_1 _4809_ (.Y(_0903_),
    .A(_0769_),
    .B(_0875_));
 sg13g2_xor2_1 _4810_ (.B(_0875_),
    .A(_0769_),
    .X(_0904_));
 sg13g2_nor2_1 _4811_ (.A(_0531_),
    .B(_0555_),
    .Y(_0905_));
 sg13g2_a21oi_1 _4812_ (.A1(_0531_),
    .A2(_0539_),
    .Y(_0906_),
    .B1(_0905_));
 sg13g2_nand2_1 _4813_ (.Y(_0907_),
    .A(net1116),
    .B(_0906_));
 sg13g2_xor2_1 _4814_ (.B(_0876_),
    .A(_0837_),
    .X(_0908_));
 sg13g2_xnor2_1 _4815_ (.Y(_0909_),
    .A(_0837_),
    .B(_0876_));
 sg13g2_nand2_1 _4816_ (.Y(_0910_),
    .A(net1130),
    .B(_0568_));
 sg13g2_o21ai_1 _4817_ (.B1(_0910_),
    .Y(_0911_),
    .A1(net1131),
    .A2(_0562_));
 sg13g2_a21oi_1 _4818_ (.A1(net1118),
    .A2(_0911_),
    .Y(_0912_),
    .B1(_0908_));
 sg13g2_nand2_1 _4819_ (.Y(_0913_),
    .A(_0907_),
    .B(_0912_));
 sg13g2_nand2_1 _4820_ (.Y(_0914_),
    .A(net1130),
    .B(_0585_));
 sg13g2_o21ai_1 _4821_ (.B1(_0914_),
    .Y(_0915_),
    .A1(net1130),
    .A2(_0590_));
 sg13g2_nor2_1 _4822_ (.A(net1130),
    .B(_0577_),
    .Y(_0916_));
 sg13g2_a21oi_1 _4823_ (.A1(net1130),
    .A2(_0573_),
    .Y(_0917_),
    .B1(_0916_));
 sg13g2_inv_1 _4824_ (.Y(_0918_),
    .A(_0917_));
 sg13g2_a21oi_1 _4825_ (.A1(net1116),
    .A2(_0915_),
    .Y(_0919_),
    .B1(_0909_));
 sg13g2_o21ai_1 _4826_ (.B1(_0919_),
    .Y(_0920_),
    .A1(net1116),
    .A2(_0917_));
 sg13g2_nand4_1 _4827_ (.B(_0901_),
    .C(_0913_),
    .A(\aliens_alive[14] ),
    .Y(_0921_),
    .D(_0920_));
 sg13g2_nand2_1 _4828_ (.Y(_0922_),
    .A(net1237),
    .B(_0756_));
 sg13g2_a22oi_1 _4829_ (.Y(_0923_),
    .B1(_0756_),
    .B2(net1237),
    .A2(_0484_),
    .A1(_2827_));
 sg13g2_or2_1 _4830_ (.X(_0924_),
    .B(_0923_),
    .A(net1366));
 sg13g2_xnor2_1 _4831_ (.Y(_0925_),
    .A(net1366),
    .B(_0923_));
 sg13g2_xnor2_1 _4832_ (.Y(_0926_),
    .A(_0075_),
    .B(_0748_));
 sg13g2_a21oi_1 _4833_ (.A1(_0768_),
    .A2(_0902_),
    .Y(_0927_),
    .B1(_0764_));
 sg13g2_a21oi_2 _4834_ (.B1(_0927_),
    .Y(_0928_),
    .A2(_0762_),
    .A1(net1384));
 sg13g2_nand2b_1 _4835_ (.Y(_0929_),
    .B(_0761_),
    .A_N(_0928_));
 sg13g2_xnor2_1 _4836_ (.Y(_0930_),
    .A(net1373),
    .B(_0926_));
 sg13g2_a21o_1 _4837_ (.A2(_0929_),
    .A1(_0774_),
    .B1(_0930_),
    .X(_0931_));
 sg13g2_o21ai_1 _4838_ (.B1(_0931_),
    .Y(_0932_),
    .A1(net1195),
    .A2(_0926_));
 sg13g2_nand2b_1 _4839_ (.Y(_0933_),
    .B(_0932_),
    .A_N(_0925_));
 sg13g2_nor2_1 _4840_ (.A(net1226),
    .B(_0922_),
    .Y(_0934_));
 sg13g2_xnor2_1 _4841_ (.Y(_0935_),
    .A(net1226),
    .B(_0922_));
 sg13g2_xor2_1 _4842_ (.B(_0935_),
    .A(net1360),
    .X(_0936_));
 sg13g2_a21oi_1 _4843_ (.A1(_0924_),
    .A2(_0933_),
    .Y(_0937_),
    .B1(_0936_));
 sg13g2_a21o_1 _4844_ (.A2(_0935_),
    .A1(net1364),
    .B1(_0937_),
    .X(_0938_));
 sg13g2_xnor2_1 _4845_ (.Y(_0939_),
    .A(_0074_),
    .B(_0934_));
 sg13g2_xor2_1 _4846_ (.B(_0939_),
    .A(net1355),
    .X(_0940_));
 sg13g2_inv_1 _4847_ (.Y(_0941_),
    .A(_0940_));
 sg13g2_nor2_1 _4848_ (.A(_0938_),
    .B(_0941_),
    .Y(_0942_));
 sg13g2_nand3_1 _4849_ (.B(_0933_),
    .C(_0936_),
    .A(_0924_),
    .Y(_0943_));
 sg13g2_nand2b_1 _4850_ (.Y(_0944_),
    .B(_0943_),
    .A_N(_0937_));
 sg13g2_xor2_1 _4851_ (.B(_0932_),
    .A(_0925_),
    .X(_0945_));
 sg13g2_nand3_1 _4852_ (.B(_0929_),
    .C(_0930_),
    .A(_0774_),
    .Y(_0946_));
 sg13g2_nand2_1 _4853_ (.Y(_0947_),
    .A(_0931_),
    .B(_0946_));
 sg13g2_xnor2_1 _4854_ (.Y(_0948_),
    .A(_0761_),
    .B(_0928_));
 sg13g2_nor2_1 _4855_ (.A(_0294_),
    .B(_0940_),
    .Y(_0949_));
 sg13g2_nand2_1 _4856_ (.Y(_0950_),
    .A(net1233),
    .B(_0934_));
 sg13g2_xnor2_1 _4857_ (.Y(_0951_),
    .A(_2820_),
    .B(_0950_));
 sg13g2_xor2_1 _4858_ (.B(_0951_),
    .A(net1352),
    .X(_0952_));
 sg13g2_xnor2_1 _4859_ (.Y(_0953_),
    .A(_0949_),
    .B(_0952_));
 sg13g2_nand4_1 _4860_ (.B(_0945_),
    .C(_0947_),
    .A(_0944_),
    .Y(_0954_),
    .D(_0953_));
 sg13g2_a21o_1 _4861_ (.A2(_0941_),
    .A1(_0938_),
    .B1(_0948_),
    .X(_0955_));
 sg13g2_nor3_2 _4862_ (.A(_0942_),
    .B(_0954_),
    .C(_0955_),
    .Y(_0956_));
 sg13g2_nand3_1 _4863_ (.B(_0768_),
    .C(_0902_),
    .A(_0764_),
    .Y(_0957_));
 sg13g2_nand2b_2 _4864_ (.Y(_0958_),
    .B(_0957_),
    .A_N(_0927_));
 sg13g2_mux4_1 _4865_ (.S0(net1116),
    .A0(_0915_),
    .A1(_0918_),
    .A2(_0906_),
    .A3(_0911_),
    .S1(_0958_),
    .X(_0959_));
 sg13g2_nand3_1 _4866_ (.B(_0956_),
    .C(_0959_),
    .A(\aliens_alive[10] ),
    .Y(_0960_));
 sg13g2_nand3_1 _4867_ (.B(_0921_),
    .C(_0960_),
    .A(_0866_),
    .Y(_0961_));
 sg13g2_or3_2 _4868_ (.A(_0713_),
    .B(_0816_),
    .C(_0961_),
    .X(_0962_));
 sg13g2_nor2_1 _4869_ (.A(net1222),
    .B(net1193),
    .Y(_0963_));
 sg13g2_nor3_1 _4870_ (.A(net1223),
    .B(net1222),
    .C(net1193),
    .Y(_0964_));
 sg13g2_o21ai_1 _4871_ (.B1(net1271),
    .Y(_0965_),
    .A1(net1274),
    .A2(_0964_));
 sg13g2_a21o_1 _4872_ (.A2(_2907_),
    .A1(net1223),
    .B1(_0964_),
    .X(_0966_));
 sg13g2_xor2_1 _4873_ (.B(net1193),
    .A(net1279),
    .X(_0967_));
 sg13g2_nor3_1 _4874_ (.A(net1222),
    .B(_0014_),
    .C(net1193),
    .Y(_0968_));
 sg13g2_nor4_1 _4875_ (.A(net1265),
    .B(_0015_),
    .C(_0967_),
    .D(_0968_),
    .Y(_0969_));
 sg13g2_xnor2_1 _4876_ (.Y(_0970_),
    .A(net1269),
    .B(_0965_));
 sg13g2_nand4_1 _4877_ (.B(_0966_),
    .C(_0969_),
    .A(_0962_),
    .Y(_0971_),
    .D(_0970_));
 sg13g2_a21o_1 _4878_ (.A2(_3213_),
    .A1(_3040_),
    .B1(net1224),
    .X(_0972_));
 sg13g2_o21ai_1 _4879_ (.B1(net1266),
    .Y(_0973_),
    .A1(net1268),
    .A2(_0972_));
 sg13g2_xnor2_1 _4880_ (.Y(_0974_),
    .A(net1225),
    .B(_0973_));
 sg13g2_nor2_2 _4881_ (.A(net1295),
    .B(_3047_),
    .Y(_0975_));
 sg13g2_nor2_1 _4882_ (.A(net1222),
    .B(_0975_),
    .Y(_0976_));
 sg13g2_o21ai_1 _4883_ (.B1(net1273),
    .Y(_0977_),
    .A1(net1276),
    .A2(_0976_));
 sg13g2_inv_1 _4884_ (.Y(_0978_),
    .A(_0977_));
 sg13g2_xor2_1 _4885_ (.B(net1266),
    .A(net1271),
    .X(_0979_));
 sg13g2_o21ai_1 _4886_ (.B1(_0978_),
    .Y(_0980_),
    .A1(_0015_),
    .A2(_0979_));
 sg13g2_o21ai_1 _4887_ (.B1(_0977_),
    .Y(_0981_),
    .A1(_2908_),
    .A2(net1266));
 sg13g2_nand2_1 _4888_ (.Y(_0982_),
    .A(net1278),
    .B(_0975_));
 sg13g2_xnor2_1 _4889_ (.Y(_0983_),
    .A(_2906_),
    .B(_0976_));
 sg13g2_xor2_1 _4890_ (.B(_0975_),
    .A(net1278),
    .X(_0984_));
 sg13g2_nor3_1 _4891_ (.A(_0014_),
    .B(_0983_),
    .C(_0984_),
    .Y(_0985_));
 sg13g2_and4_2 _4892_ (.A(_0974_),
    .B(_0980_),
    .C(_0981_),
    .D(_0985_),
    .X(_0986_));
 sg13g2_nand2_2 _4893_ (.Y(_0987_),
    .A(net1282),
    .B(_3192_));
 sg13g2_xnor2_1 _4894_ (.Y(_0988_),
    .A(_2905_),
    .B(_3044_));
 sg13g2_inv_1 _4895_ (.Y(_0989_),
    .A(_0988_));
 sg13g2_a22oi_1 _4896_ (.Y(_0990_),
    .B1(_3191_),
    .B2(_0048_),
    .A2(_3181_),
    .A1(net1213));
 sg13g2_or2_1 _4897_ (.X(_0991_),
    .B(_0990_),
    .A(net1159));
 sg13g2_nand2_1 _4898_ (.Y(_0992_),
    .A(_0987_),
    .B(_0991_));
 sg13g2_nor2_1 _4899_ (.A(net1398),
    .B(_0992_),
    .Y(_0993_));
 sg13g2_nand2_1 _4900_ (.Y(_0994_),
    .A(_3191_),
    .B(_0550_));
 sg13g2_nor2_1 _4901_ (.A(_0552_),
    .B(net1159),
    .Y(_0995_));
 sg13g2_a21oi_1 _4902_ (.A1(net1159),
    .A2(_0994_),
    .Y(_0996_),
    .B1(_0995_));
 sg13g2_a21oi_2 _4903_ (.B1(_0993_),
    .Y(_0997_),
    .A2(_0996_),
    .A1(net1399));
 sg13g2_a21oi_1 _4904_ (.A1(net1297),
    .A2(net1282),
    .Y(_0998_),
    .B1(net1290));
 sg13g2_nand2_1 _4905_ (.Y(_0999_),
    .A(net1207),
    .B(_0998_));
 sg13g2_nand3_1 _4906_ (.B(_0313_),
    .C(_0989_),
    .A(_3177_),
    .Y(_1000_));
 sg13g2_o21ai_1 _4907_ (.B1(_0999_),
    .Y(_1001_),
    .A1(net1207),
    .A2(_1000_));
 sg13g2_nand2_1 _4908_ (.Y(_1002_),
    .A(net1126),
    .B(_1001_));
 sg13g2_o21ai_1 _4909_ (.B1(_1002_),
    .Y(_1003_),
    .A1(net1125),
    .A2(_0997_));
 sg13g2_nor2_1 _4910_ (.A(net1215),
    .B(_0544_),
    .Y(_1004_));
 sg13g2_nand2_1 _4911_ (.Y(_1005_),
    .A(net1292),
    .B(_0543_));
 sg13g2_o21ai_1 _4912_ (.B1(net1282),
    .Y(_1006_),
    .A1(_3190_),
    .A2(_1004_));
 sg13g2_nor2_1 _4913_ (.A(_3192_),
    .B(net1159),
    .Y(_1007_));
 sg13g2_nor2b_1 _4914_ (.A(_1007_),
    .B_N(_1006_),
    .Y(_1008_));
 sg13g2_o21ai_1 _4915_ (.B1(_0987_),
    .Y(_1009_),
    .A1(net1159),
    .A2(_0994_));
 sg13g2_nor2_1 _4916_ (.A(net1205),
    .B(_1009_),
    .Y(_1010_));
 sg13g2_a21oi_2 _4917_ (.B1(_1010_),
    .Y(_1011_),
    .A2(_1008_),
    .A1(net1205));
 sg13g2_nor2_1 _4918_ (.A(_3209_),
    .B(_0322_),
    .Y(_1012_));
 sg13g2_nand2b_2 _4919_ (.Y(_1013_),
    .B(_0323_),
    .A_N(_3209_));
 sg13g2_nor2_1 _4920_ (.A(net1125),
    .B(_1012_),
    .Y(_1014_));
 sg13g2_a21oi_1 _4921_ (.A1(net1125),
    .A2(_1011_),
    .Y(_1015_),
    .B1(_1014_));
 sg13g2_nor2_2 _4922_ (.A(_3209_),
    .B(_0310_),
    .Y(_1016_));
 sg13g2_a21o_1 _4923_ (.A2(_3190_),
    .A1(net1284),
    .B1(_1007_),
    .X(_1017_));
 sg13g2_nor2_1 _4924_ (.A(net1205),
    .B(_1017_),
    .Y(_1018_));
 sg13g2_a21oi_1 _4925_ (.A1(net1205),
    .A2(_1016_),
    .Y(_1019_),
    .B1(_1018_));
 sg13g2_o21ai_1 _4926_ (.B1(_0987_),
    .Y(_1020_),
    .A1(_0552_),
    .A2(net1159));
 sg13g2_and2_1 _4927_ (.A(_0991_),
    .B(_1006_),
    .X(_1021_));
 sg13g2_nand2_1 _4928_ (.Y(_1022_),
    .A(net1397),
    .B(_1021_));
 sg13g2_o21ai_1 _4929_ (.B1(_1022_),
    .Y(_1023_),
    .A1(net1398),
    .A2(_1020_));
 sg13g2_nor2_1 _4930_ (.A(net1124),
    .B(_1023_),
    .Y(_1024_));
 sg13g2_a21oi_1 _4931_ (.A1(net1124),
    .A2(_1019_),
    .Y(_1025_),
    .B1(_1024_));
 sg13g2_nor2_1 _4932_ (.A(_3197_),
    .B(net1159),
    .Y(_1026_));
 sg13g2_a21oi_1 _4933_ (.A1(net1159),
    .A2(_0994_),
    .Y(_1027_),
    .B1(_1026_));
 sg13g2_o21ai_1 _4934_ (.B1(_0987_),
    .Y(_1028_),
    .A1(net1215),
    .A2(net1284));
 sg13g2_nor2_1 _4935_ (.A(net1398),
    .B(_1027_),
    .Y(_1029_));
 sg13g2_a21oi_2 _4936_ (.B1(_1029_),
    .Y(_1030_),
    .A2(_1028_),
    .A1(net1398));
 sg13g2_and3_1 _4937_ (.X(_1031_),
    .A(_2905_),
    .B(_3045_),
    .C(_0313_));
 sg13g2_o21ai_1 _4938_ (.B1(net1402),
    .Y(_1032_),
    .A1(net1282),
    .A2(_3195_));
 sg13g2_o21ai_1 _4939_ (.B1(_1032_),
    .Y(_1033_),
    .A1(net1400),
    .A2(_1031_));
 sg13g2_nand2_1 _4940_ (.Y(_1034_),
    .A(net1125),
    .B(_1030_));
 sg13g2_o21ai_1 _4941_ (.B1(_1034_),
    .Y(_1035_),
    .A1(net1125),
    .A2(_1033_));
 sg13g2_mux4_1 _4942_ (.S0(_0528_),
    .A0(_1035_),
    .A1(_1025_),
    .A2(_1015_),
    .A3(_1003_),
    .S1(_0558_),
    .X(_1036_));
 sg13g2_nand3_1 _4943_ (.B(_0527_),
    .C(_1036_),
    .A(\aliens_alive[20] ),
    .Y(_1037_));
 sg13g2_nor3_1 _4944_ (.A(net1402),
    .B(net1282),
    .C(_3195_),
    .Y(_1038_));
 sg13g2_a21o_1 _4945_ (.A2(_1031_),
    .A1(net1400),
    .B1(_1038_),
    .X(_1039_));
 sg13g2_nor2_1 _4946_ (.A(net1398),
    .B(_1028_),
    .Y(_1040_));
 sg13g2_a21oi_1 _4947_ (.A1(net1397),
    .A2(_1027_),
    .Y(_1041_),
    .B1(_1040_));
 sg13g2_nor2_1 _4948_ (.A(net1102),
    .B(_1041_),
    .Y(_1042_));
 sg13g2_a21oi_2 _4949_ (.B1(_1042_),
    .Y(_1043_),
    .A2(_1039_),
    .A1(net1103));
 sg13g2_nor2_1 _4950_ (.A(net1397),
    .B(_1021_),
    .Y(_1044_));
 sg13g2_a21oi_1 _4951_ (.A1(net1397),
    .A2(_1020_),
    .Y(_1045_),
    .B1(_1044_));
 sg13g2_nor2_1 _4952_ (.A(net1397),
    .B(_1017_),
    .Y(_1046_));
 sg13g2_a21oi_1 _4953_ (.A1(net1397),
    .A2(_1016_),
    .Y(_1047_),
    .B1(_1046_));
 sg13g2_nor2_1 _4954_ (.A(net1102),
    .B(_1047_),
    .Y(_1048_));
 sg13g2_a21oi_2 _4955_ (.B1(_1048_),
    .Y(_1049_),
    .A2(_1045_),
    .A1(net1102));
 sg13g2_nor2_1 _4956_ (.A(net1084),
    .B(_1049_),
    .Y(_1050_));
 sg13g2_nor2_1 _4957_ (.A(_0706_),
    .B(_1050_),
    .Y(_1051_));
 sg13g2_o21ai_1 _4958_ (.B1(_1051_),
    .Y(_1052_),
    .A1(net1087),
    .A2(_1043_));
 sg13g2_nor2_1 _4959_ (.A(net1205),
    .B(_0992_),
    .Y(_1053_));
 sg13g2_a21oi_1 _4960_ (.A1(net1205),
    .A2(_0996_),
    .Y(_1054_),
    .B1(_1053_));
 sg13g2_nand2_1 _4961_ (.Y(_1055_),
    .A(net1400),
    .B(_0998_));
 sg13g2_o21ai_1 _4962_ (.B1(_1055_),
    .Y(_1056_),
    .A1(net1400),
    .A2(_1000_));
 sg13g2_nor2_1 _4963_ (.A(net1105),
    .B(_1056_),
    .Y(_1057_));
 sg13g2_a21oi_1 _4964_ (.A1(net1105),
    .A2(_1054_),
    .Y(_1058_),
    .B1(_1057_));
 sg13g2_nand2_1 _4965_ (.Y(_1059_),
    .A(net1087),
    .B(_1058_));
 sg13g2_nand2_1 _4966_ (.Y(_1060_),
    .A(net1398),
    .B(_1008_));
 sg13g2_o21ai_1 _4967_ (.B1(_1060_),
    .Y(_1061_),
    .A1(net1397),
    .A2(_1009_));
 sg13g2_nor2_1 _4968_ (.A(net1103),
    .B(_1061_),
    .Y(_1062_));
 sg13g2_a21oi_1 _4969_ (.A1(net1105),
    .A2(_1013_),
    .Y(_1063_),
    .B1(_1062_));
 sg13g2_nand2_1 _4970_ (.Y(_1064_),
    .A(net1084),
    .B(_1063_));
 sg13g2_nand3_1 _4971_ (.B(_1059_),
    .C(_1064_),
    .A(_0706_),
    .Y(_1065_));
 sg13g2_nand4_1 _4972_ (.B(_0705_),
    .C(_1052_),
    .A(\aliens_alive[19] ),
    .Y(_1066_),
    .D(_1065_));
 sg13g2_nor2_1 _4973_ (.A(net1087),
    .B(_1049_),
    .Y(_1067_));
 sg13g2_nor2_1 _4974_ (.A(_0650_),
    .B(_1067_),
    .Y(_1068_));
 sg13g2_o21ai_1 _4975_ (.B1(_1068_),
    .Y(_1069_),
    .A1(net1084),
    .A2(_1043_));
 sg13g2_nand2_1 _4976_ (.Y(_1070_),
    .A(net1087),
    .B(_1063_));
 sg13g2_a21oi_1 _4977_ (.A1(net1084),
    .A2(_1058_),
    .Y(_1071_),
    .B1(_0651_));
 sg13g2_nand2_1 _4978_ (.Y(_1072_),
    .A(_1070_),
    .B(_1071_));
 sg13g2_nand4_1 _4979_ (.B(_0640_),
    .C(_1069_),
    .A(\aliens_alive[23] ),
    .Y(_1073_),
    .D(_1072_));
 sg13g2_nand3_1 _4980_ (.B(_1066_),
    .C(_1073_),
    .A(_1037_),
    .Y(_1074_));
 sg13g2_nand2_1 _4981_ (.Y(_1075_),
    .A(_0986_),
    .B(_1074_));
 sg13g2_nand2_1 _4982_ (.Y(_1076_),
    .A(net1102),
    .B(_1041_));
 sg13g2_o21ai_1 _4983_ (.B1(_1076_),
    .Y(_1077_),
    .A1(net1104),
    .A2(_1039_));
 sg13g2_nand2_1 _4984_ (.Y(_1078_),
    .A(net1102),
    .B(_1047_));
 sg13g2_o21ai_1 _4985_ (.B1(_1078_),
    .Y(_1079_),
    .A1(net1102),
    .A2(_1045_));
 sg13g2_nor2_1 _4986_ (.A(net1103),
    .B(_1013_),
    .Y(_1080_));
 sg13g2_a21oi_1 _4987_ (.A1(net1103),
    .A2(_1061_),
    .Y(_1081_),
    .B1(_1080_));
 sg13g2_nor2_1 _4988_ (.A(net1104),
    .B(_1054_),
    .Y(_1082_));
 sg13g2_a21oi_1 _4989_ (.A1(net1106),
    .A2(_1056_),
    .Y(_1083_),
    .B1(_1082_));
 sg13g2_mux4_1 _4990_ (.S0(net1120),
    .A0(_1077_),
    .A1(_1079_),
    .A2(_1081_),
    .A3(_1083_),
    .S1(_0864_),
    .X(_1084_));
 sg13g2_inv_1 _4991_ (.Y(_1085_),
    .A(_1084_));
 sg13g2_nand4_1 _4992_ (.B(_0863_),
    .C(_0986_),
    .A(\aliens_alive[21] ),
    .Y(_1086_),
    .D(_1085_));
 sg13g2_mux4_1 _4993_ (.S0(_0528_),
    .A0(_1003_),
    .A1(_1015_),
    .A2(_1025_),
    .A3(_1035_),
    .S1(_0743_),
    .X(_1087_));
 sg13g2_nand4_1 _4994_ (.B(_0742_),
    .C(_0986_),
    .A(\aliens_alive[16] ),
    .Y(_1088_),
    .D(_1087_));
 sg13g2_mux4_1 _4995_ (.S0(net1121),
    .A0(_1077_),
    .A1(_1079_),
    .A2(_1081_),
    .A3(_1083_),
    .S1(_0804_),
    .X(_1089_));
 sg13g2_inv_1 _4996_ (.Y(_1090_),
    .A(_1089_));
 sg13g2_nand4_1 _4997_ (.B(_0798_),
    .C(_0986_),
    .A(\aliens_alive[17] ),
    .Y(_1091_),
    .D(_1090_));
 sg13g2_and2_1 _4998_ (.A(_1088_),
    .B(_1091_),
    .X(_1092_));
 sg13g2_nor2_1 _4999_ (.A(_0531_),
    .B(_0997_),
    .Y(_1093_));
 sg13g2_a21oi_1 _5000_ (.A1(_0531_),
    .A2(_1001_),
    .Y(_1094_),
    .B1(_1093_));
 sg13g2_nand2_1 _5001_ (.Y(_1095_),
    .A(net1126),
    .B(_1012_));
 sg13g2_o21ai_1 _5002_ (.B1(_1095_),
    .Y(_1096_),
    .A1(net1125),
    .A2(_1011_));
 sg13g2_a21oi_1 _5003_ (.A1(net1117),
    .A2(_1094_),
    .Y(_1097_),
    .B1(_0958_));
 sg13g2_o21ai_1 _5004_ (.B1(_1097_),
    .Y(_1098_),
    .A1(net1117),
    .A2(_1096_));
 sg13g2_nand2_1 _5005_ (.Y(_1099_),
    .A(net1125),
    .B(_1033_));
 sg13g2_o21ai_1 _5006_ (.B1(_1099_),
    .Y(_1100_),
    .A1(net1125),
    .A2(_1030_));
 sg13g2_nand2_1 _5007_ (.Y(_1101_),
    .A(net1115),
    .B(_1100_));
 sg13g2_nor2_1 _5008_ (.A(net1124),
    .B(_1019_),
    .Y(_1102_));
 sg13g2_a21oi_2 _5009_ (.B1(_1102_),
    .Y(_1103_),
    .A2(_1023_),
    .A1(net1124));
 sg13g2_nand2_1 _5010_ (.Y(_1104_),
    .A(net1117),
    .B(_1103_));
 sg13g2_nand3_1 _5011_ (.B(_1101_),
    .C(_1104_),
    .A(_0958_),
    .Y(_1105_));
 sg13g2_nand2_1 _5012_ (.Y(_1106_),
    .A(_1098_),
    .B(_1105_));
 sg13g2_nand4_1 _5013_ (.B(_0956_),
    .C(_0986_),
    .A(\aliens_alive[18] ),
    .Y(_1107_),
    .D(_1106_));
 sg13g2_a21oi_1 _5014_ (.A1(net1115),
    .A2(_1094_),
    .Y(_1108_),
    .B1(_0909_));
 sg13g2_o21ai_1 _5015_ (.B1(_1108_),
    .Y(_1109_),
    .A1(net1115),
    .A2(_1096_));
 sg13g2_mux2_1 _5016_ (.A0(_1100_),
    .A1(_1103_),
    .S(net1115),
    .X(_1110_));
 sg13g2_o21ai_1 _5017_ (.B1(_1109_),
    .Y(_1111_),
    .A1(_0908_),
    .A2(_1110_));
 sg13g2_nand4_1 _5018_ (.B(_0901_),
    .C(_0986_),
    .A(\aliens_alive[22] ),
    .Y(_1112_),
    .D(_1111_));
 sg13g2_nand4_1 _5019_ (.B(_1092_),
    .C(_1107_),
    .A(_1086_),
    .Y(_1113_),
    .D(_1112_));
 sg13g2_nand3b_1 _5020_ (.B(_1075_),
    .C(_0971_),
    .Y(_1114_),
    .A_N(_1113_));
 sg13g2_nor2_2 _5021_ (.A(_0010_),
    .B(net1187),
    .Y(_1115_));
 sg13g2_nor3_2 _5022_ (.A(_0010_),
    .B(_2905_),
    .C(net1187),
    .Y(_1116_));
 sg13g2_nor2_2 _5023_ (.A(net1163),
    .B(_0534_),
    .Y(_1117_));
 sg13g2_a21oi_1 _5024_ (.A1(net1218),
    .A2(_1115_),
    .Y(_1118_),
    .B1(_1117_));
 sg13g2_nor2_1 _5025_ (.A(net1208),
    .B(_1118_),
    .Y(_1119_));
 sg13g2_a21oi_1 _5026_ (.A1(net1208),
    .A2(_1116_),
    .Y(_1120_),
    .B1(_1119_));
 sg13g2_nor2_2 _5027_ (.A(net1218),
    .B(_0315_),
    .Y(_1121_));
 sg13g2_nand2b_1 _5028_ (.Y(_1122_),
    .B(net1287),
    .A_N(_0315_));
 sg13g2_a21oi_1 _5029_ (.A1(_3043_),
    .A2(_3191_),
    .Y(_1123_),
    .B1(_1121_));
 sg13g2_nand2_1 _5030_ (.Y(_1124_),
    .A(net1218),
    .B(_0550_));
 sg13g2_and2_1 _5031_ (.A(net1218),
    .B(_0552_),
    .X(_1125_));
 sg13g2_a21oi_1 _5032_ (.A1(_3200_),
    .A2(_0543_),
    .Y(_1126_),
    .B1(_1125_));
 sg13g2_nand2_1 _5033_ (.Y(_1127_),
    .A(net1405),
    .B(_1123_));
 sg13g2_o21ai_1 _5034_ (.B1(_1127_),
    .Y(_1128_),
    .A1(net1405),
    .A2(_1126_));
 sg13g2_nand2_1 _5035_ (.Y(_1129_),
    .A(net1108),
    .B(_1128_));
 sg13g2_o21ai_1 _5036_ (.B1(_1129_),
    .Y(_1130_),
    .A1(net1109),
    .A2(_1120_));
 sg13g2_nand2b_1 _5037_ (.Y(_1131_),
    .B(_1122_),
    .A_N(_3181_));
 sg13g2_nor2_1 _5038_ (.A(net1403),
    .B(_1131_),
    .Y(_1132_));
 sg13g2_a21oi_2 _5039_ (.B1(_1121_),
    .Y(_1133_),
    .A2(_3046_),
    .A1(net1212));
 sg13g2_inv_1 _5040_ (.Y(_1134_),
    .A(_1133_));
 sg13g2_a21oi_1 _5041_ (.A1(net1403),
    .A2(_1133_),
    .Y(_1135_),
    .B1(_1132_));
 sg13g2_nand2_1 _5042_ (.Y(_1136_),
    .A(net1107),
    .B(_1135_));
 sg13g2_a22oi_1 _5043_ (.Y(_1137_),
    .B1(_0544_),
    .B2(_3200_),
    .A2(_0542_),
    .A1(net1189));
 sg13g2_and2_1 _5044_ (.A(net1208),
    .B(_1137_),
    .X(_1138_));
 sg13g2_a21oi_2 _5045_ (.B1(_0445_),
    .Y(_1139_),
    .A2(_0315_),
    .A1(net1163));
 sg13g2_nor3_2 _5046_ (.A(_3201_),
    .B(_0446_),
    .C(_1121_),
    .Y(_1140_));
 sg13g2_a21oi_1 _5047_ (.A1(net1403),
    .A2(_1139_),
    .Y(_1141_),
    .B1(_1138_));
 sg13g2_o21ai_1 _5048_ (.B1(_1136_),
    .Y(_1142_),
    .A1(net1108),
    .A2(_1141_));
 sg13g2_inv_1 _5049_ (.Y(_1143_),
    .A(_1142_));
 sg13g2_nor2_1 _5050_ (.A(_1117_),
    .B(_1125_),
    .Y(_1144_));
 sg13g2_nand2_1 _5051_ (.Y(_1145_),
    .A(net1403),
    .B(_1144_));
 sg13g2_nor2_1 _5052_ (.A(net1287),
    .B(_3194_),
    .Y(_1146_));
 sg13g2_a22oi_1 _5053_ (.Y(_1147_),
    .B1(_1005_),
    .B2(_1146_),
    .A2(_0453_),
    .A1(net1287));
 sg13g2_o21ai_1 _5054_ (.B1(_1145_),
    .Y(_1148_),
    .A1(net1403),
    .A2(_1147_));
 sg13g2_nand2_1 _5055_ (.Y(_1149_),
    .A(net1107),
    .B(_1116_));
 sg13g2_o21ai_1 _5056_ (.B1(_1149_),
    .Y(_1150_),
    .A1(net1108),
    .A2(_1148_));
 sg13g2_o21ai_1 _5057_ (.B1(_1122_),
    .Y(_1151_),
    .A1(_3194_),
    .A2(_1124_));
 sg13g2_mux2_1 _5058_ (.A0(_1137_),
    .A1(_1151_),
    .S(net1208),
    .X(_1152_));
 sg13g2_nor2_1 _5059_ (.A(net1107),
    .B(_1152_),
    .Y(_1153_));
 sg13g2_a21oi_1 _5060_ (.A1(net1107),
    .A2(_1140_),
    .Y(_1154_),
    .B1(_1153_));
 sg13g2_inv_1 _5061_ (.Y(_1155_),
    .A(_1154_));
 sg13g2_mux4_1 _5062_ (.S0(net1085),
    .A0(_1143_),
    .A1(_1150_),
    .A2(_1130_),
    .A3(_1155_),
    .S1(_0706_),
    .X(_1156_));
 sg13g2_nand3_1 _5063_ (.B(_0705_),
    .C(_1156_),
    .A(\aliens_alive[27] ),
    .Y(_1157_));
 sg13g2_a21oi_1 _5064_ (.A1(net1085),
    .A2(_1130_),
    .Y(_1158_),
    .B1(_0651_));
 sg13g2_o21ai_1 _5065_ (.B1(_1158_),
    .Y(_1159_),
    .A1(net1085),
    .A2(_1154_));
 sg13g2_o21ai_1 _5066_ (.B1(_0651_),
    .Y(_1160_),
    .A1(net1087),
    .A2(_1142_));
 sg13g2_a21o_1 _5067_ (.A2(_1150_),
    .A1(net1087),
    .B1(_1160_),
    .X(_1161_));
 sg13g2_nand4_1 _5068_ (.B(_0640_),
    .C(_1159_),
    .A(\aliens_alive[31] ),
    .Y(_1162_),
    .D(_1161_));
 sg13g2_nor2_1 _5069_ (.A(net1405),
    .B(_1144_),
    .Y(_1163_));
 sg13g2_a21oi_1 _5070_ (.A1(net1403),
    .A2(_1147_),
    .Y(_1164_),
    .B1(_1163_));
 sg13g2_nand2_1 _5071_ (.Y(_1165_),
    .A(net1127),
    .B(_1164_));
 sg13g2_o21ai_1 _5072_ (.B1(_1165_),
    .Y(_1166_),
    .A1(net1127),
    .A2(_1116_));
 sg13g2_nor2_1 _5073_ (.A(net1404),
    .B(_1140_),
    .Y(_1167_));
 sg13g2_a21oi_1 _5074_ (.A1(net1403),
    .A2(_1137_),
    .Y(_1168_),
    .B1(_1167_));
 sg13g2_nor2_1 _5075_ (.A(net1208),
    .B(_1131_),
    .Y(_1169_));
 sg13g2_a21oi_1 _5076_ (.A1(net1208),
    .A2(_1133_),
    .Y(_1170_),
    .B1(_1169_));
 sg13g2_nor2_1 _5077_ (.A(net1127),
    .B(_1170_),
    .Y(_1171_));
 sg13g2_a21oi_1 _5078_ (.A1(net1128),
    .A2(_1168_),
    .Y(_1172_),
    .B1(_1171_));
 sg13g2_nor2_1 _5079_ (.A(net1128),
    .B(_1139_),
    .Y(_1173_));
 sg13g2_a21oi_1 _5080_ (.A1(net1403),
    .A2(_1151_),
    .Y(_1174_),
    .B1(_1138_));
 sg13g2_a21oi_1 _5081_ (.A1(net1127),
    .A2(_1174_),
    .Y(_1175_),
    .B1(_1173_));
 sg13g2_nor2_1 _5082_ (.A(net1405),
    .B(_1123_),
    .Y(_1176_));
 sg13g2_a21oi_1 _5083_ (.A1(net1405),
    .A2(_1126_),
    .Y(_1177_),
    .B1(_1176_));
 sg13g2_nand2_1 _5084_ (.Y(_1178_),
    .A(net1406),
    .B(_1116_));
 sg13g2_o21ai_1 _5085_ (.B1(_1178_),
    .Y(_1179_),
    .A1(net1406),
    .A2(_1118_));
 sg13g2_and2_1 _5086_ (.A(net1127),
    .B(_1179_),
    .X(_1180_));
 sg13g2_a21oi_1 _5087_ (.A1(_0531_),
    .A2(_1177_),
    .Y(_1181_),
    .B1(_1180_));
 sg13g2_mux4_1 _5088_ (.S0(_0528_),
    .A0(_1166_),
    .A1(_1172_),
    .A2(_1175_),
    .A3(_1181_),
    .S1(_0558_),
    .X(_1182_));
 sg13g2_inv_1 _5089_ (.Y(_1183_),
    .A(_1182_));
 sg13g2_nand3_1 _5090_ (.B(_0527_),
    .C(_1183_),
    .A(\aliens_alive[28] ),
    .Y(_1184_));
 sg13g2_nand3_1 _5091_ (.B(_1162_),
    .C(_1184_),
    .A(_1157_),
    .Y(_1185_));
 sg13g2_mux4_1 _5092_ (.S0(_0529_),
    .A0(_1175_),
    .A1(_1181_),
    .A2(_1166_),
    .A3(_1172_),
    .S1(_0743_),
    .X(_1186_));
 sg13g2_inv_1 _5093_ (.Y(_1187_),
    .A(_1186_));
 sg13g2_and3_1 _5094_ (.X(_1188_),
    .A(\aliens_alive[24] ),
    .B(_0742_),
    .C(_1187_));
 sg13g2_nor2_1 _5095_ (.A(net1109),
    .B(_1140_),
    .Y(_1189_));
 sg13g2_a21oi_1 _5096_ (.A1(net1107),
    .A2(_1152_),
    .Y(_1190_),
    .B1(_1189_));
 sg13g2_nand2_1 _5097_ (.Y(_1191_),
    .A(_0801_),
    .B(_1190_));
 sg13g2_nor2_1 _5098_ (.A(net1109),
    .B(_1128_),
    .Y(_1192_));
 sg13g2_a21oi_1 _5099_ (.A1(net1109),
    .A2(_1120_),
    .Y(_1193_),
    .B1(_1192_));
 sg13g2_nand2_1 _5100_ (.Y(_1194_),
    .A(net1122),
    .B(_1193_));
 sg13g2_nand3_1 _5101_ (.B(_1191_),
    .C(_1194_),
    .A(_0804_),
    .Y(_1195_));
 sg13g2_nor2_1 _5102_ (.A(net1108),
    .B(_1116_),
    .Y(_1196_));
 sg13g2_a21oi_1 _5103_ (.A1(net1107),
    .A2(_1148_),
    .Y(_1197_),
    .B1(_1196_));
 sg13g2_nor2_1 _5104_ (.A(net1107),
    .B(_1135_),
    .Y(_1198_));
 sg13g2_a21oi_1 _5105_ (.A1(net1107),
    .A2(_1141_),
    .Y(_1199_),
    .B1(_1198_));
 sg13g2_a21oi_1 _5106_ (.A1(net1120),
    .A2(_1197_),
    .Y(_1200_),
    .B1(_0804_));
 sg13g2_o21ai_1 _5107_ (.B1(_1200_),
    .Y(_1201_),
    .A1(net1120),
    .A2(_1199_));
 sg13g2_and4_1 _5108_ (.A(\aliens_alive[25] ),
    .B(_0798_),
    .C(_1195_),
    .D(_1201_),
    .X(_1202_));
 sg13g2_nor2_1 _5109_ (.A(net1127),
    .B(_1174_),
    .Y(_1203_));
 sg13g2_a21oi_1 _5110_ (.A1(net1127),
    .A2(_1139_),
    .Y(_1204_),
    .B1(_1203_));
 sg13g2_nand2_1 _5111_ (.Y(_1205_),
    .A(net1117),
    .B(_1204_));
 sg13g2_mux2_1 _5112_ (.A0(_1177_),
    .A1(_1179_),
    .S(_0531_),
    .X(_1206_));
 sg13g2_a21oi_1 _5113_ (.A1(net1115),
    .A2(_1206_),
    .Y(_1207_),
    .B1(_0909_));
 sg13g2_nor2_1 _5114_ (.A(net1127),
    .B(_1164_),
    .Y(_1208_));
 sg13g2_a21oi_1 _5115_ (.A1(net1128),
    .A2(_1116_),
    .Y(_1209_),
    .B1(_1208_));
 sg13g2_inv_1 _5116_ (.Y(_1210_),
    .A(_1209_));
 sg13g2_nand2_1 _5117_ (.Y(_1211_),
    .A(net1128),
    .B(_1170_));
 sg13g2_o21ai_1 _5118_ (.B1(_1211_),
    .Y(_1212_),
    .A1(net1128),
    .A2(_1168_));
 sg13g2_inv_1 _5119_ (.Y(_1213_),
    .A(_1212_));
 sg13g2_nor2_1 _5120_ (.A(net1117),
    .B(_1212_),
    .Y(_1214_));
 sg13g2_a21oi_1 _5121_ (.A1(net1117),
    .A2(_1210_),
    .Y(_1215_),
    .B1(_1214_));
 sg13g2_a22oi_1 _5122_ (.Y(_1216_),
    .B1(_1215_),
    .B2(_0909_),
    .A2(_1207_),
    .A1(_1205_));
 sg13g2_nand3_1 _5123_ (.B(_0901_),
    .C(_1216_),
    .A(\aliens_alive[30] ),
    .Y(_1217_));
 sg13g2_mux4_1 _5124_ (.S0(net1117),
    .A0(_1204_),
    .A1(_1206_),
    .A2(_1210_),
    .A3(_1213_),
    .S1(_0958_),
    .X(_1218_));
 sg13g2_nand3_1 _5125_ (.B(_0956_),
    .C(_1218_),
    .A(\aliens_alive[26] ),
    .Y(_1219_));
 sg13g2_nand2_1 _5126_ (.Y(_1220_),
    .A(net1120),
    .B(_1193_));
 sg13g2_nand2_1 _5127_ (.Y(_1221_),
    .A(net1121),
    .B(_1190_));
 sg13g2_nand3_1 _5128_ (.B(_1220_),
    .C(_1221_),
    .A(_0864_),
    .Y(_1222_));
 sg13g2_a21oi_1 _5129_ (.A1(net1121),
    .A2(_1197_),
    .Y(_1223_),
    .B1(_0864_));
 sg13g2_o21ai_1 _5130_ (.B1(_1223_),
    .Y(_1224_),
    .A1(net1121),
    .A2(_1199_));
 sg13g2_nand4_1 _5131_ (.B(_0863_),
    .C(_1222_),
    .A(\aliens_alive[29] ),
    .Y(_1225_),
    .D(_1224_));
 sg13g2_nand3_1 _5132_ (.B(_1219_),
    .C(_1225_),
    .A(_1217_),
    .Y(_1226_));
 sg13g2_nor4_2 _5133_ (.A(_1185_),
    .B(_1188_),
    .C(_1202_),
    .Y(_1227_),
    .D(_1226_));
 sg13g2_a21oi_2 _5134_ (.B1(_0014_),
    .Y(_1228_),
    .A2(net1266),
    .A1(net1271));
 sg13g2_o21ai_1 _5135_ (.B1(_0014_),
    .Y(_1229_),
    .A1(net1271),
    .A2(net1266));
 sg13g2_nor2_1 _5136_ (.A(net1265),
    .B(net1222),
    .Y(_1230_));
 sg13g2_nand4_1 _5137_ (.B(net1276),
    .C(_1229_),
    .A(net1274),
    .Y(_1231_),
    .D(_1230_));
 sg13g2_nor3_1 _5138_ (.A(_1227_),
    .B(_1228_),
    .C(_1231_),
    .Y(_1232_));
 sg13g2_a21oi_1 _5139_ (.A1(net1295),
    .A2(_0533_),
    .Y(_1233_),
    .B1(net1280));
 sg13g2_o21ai_1 _5140_ (.B1(_0013_),
    .Y(_1234_),
    .A1(net1271),
    .A2(_1233_));
 sg13g2_nand2_1 _5141_ (.Y(_1235_),
    .A(net1223),
    .B(_3041_));
 sg13g2_a21oi_1 _5142_ (.A1(_1233_),
    .A2(_1235_),
    .Y(_1236_),
    .B1(_0013_));
 sg13g2_nor2_1 _5143_ (.A(_3040_),
    .B(_3041_),
    .Y(_1237_));
 sg13g2_xnor2_1 _5144_ (.Y(_1238_),
    .A(net1264),
    .B(net1269));
 sg13g2_xnor2_1 _5145_ (.Y(_1239_),
    .A(net1278),
    .B(_0309_));
 sg13g2_nor4_1 _5146_ (.A(net1267),
    .B(_1236_),
    .C(_1237_),
    .D(_1238_),
    .Y(_1240_));
 sg13g2_and3_2 _5147_ (.X(_1241_),
    .A(_1234_),
    .B(_1239_),
    .C(_1240_));
 sg13g2_nor2b_2 _5148_ (.A(_0309_),
    .B_N(_3210_),
    .Y(_1242_));
 sg13g2_nand2b_2 _5149_ (.Y(_1243_),
    .B(_3210_),
    .A_N(_0309_));
 sg13g2_nand2b_1 _5150_ (.Y(_1244_),
    .B(_1005_),
    .A_N(_0315_));
 sg13g2_a21oi_1 _5151_ (.A1(_1243_),
    .A2(_1244_),
    .Y(_1245_),
    .B1(_3196_));
 sg13g2_nand2_1 _5152_ (.Y(_1246_),
    .A(net1401),
    .B(_1245_));
 sg13g2_nor2_1 _5153_ (.A(net1282),
    .B(_3196_),
    .Y(_1247_));
 sg13g2_inv_1 _5154_ (.Y(_1248_),
    .A(_1247_));
 sg13g2_a21oi_1 _5155_ (.A1(net1212),
    .A2(_1007_),
    .Y(_1249_),
    .B1(_1247_));
 sg13g2_o21ai_1 _5156_ (.B1(_1246_),
    .Y(_1250_),
    .A1(net1400),
    .A2(_1249_));
 sg13g2_and3_1 _5157_ (.X(_1251_),
    .A(_3177_),
    .B(_3183_),
    .C(_1242_));
 sg13g2_a21oi_1 _5158_ (.A1(_3177_),
    .A2(_3193_),
    .Y(_1252_),
    .B1(_1242_));
 sg13g2_nor2_1 _5159_ (.A(_1251_),
    .B(_1252_),
    .Y(_1253_));
 sg13g2_nor2_1 _5160_ (.A(net1206),
    .B(_1253_),
    .Y(_1254_));
 sg13g2_nor2_1 _5161_ (.A(_0541_),
    .B(_0987_),
    .Y(_1255_));
 sg13g2_or2_2 _5162_ (.X(_1256_),
    .B(_1255_),
    .A(_1251_));
 sg13g2_a21oi_1 _5163_ (.A1(net1207),
    .A2(_1256_),
    .Y(_1257_),
    .B1(_1254_));
 sg13g2_nor2_1 _5164_ (.A(net1123),
    .B(_1257_),
    .Y(_1258_));
 sg13g2_a21oi_2 _5165_ (.B1(_1258_),
    .Y(_1259_),
    .A2(_1250_),
    .A1(net1126));
 sg13g2_a21oi_1 _5166_ (.A1(net1212),
    .A2(_3190_),
    .Y(_1260_),
    .B1(_1243_));
 sg13g2_o21ai_1 _5167_ (.B1(_1243_),
    .Y(_1261_),
    .A1(_3190_),
    .A2(_1004_));
 sg13g2_nor2b_1 _5168_ (.A(_1260_),
    .B_N(_1261_),
    .Y(_1262_));
 sg13g2_nand2_1 _5169_ (.Y(_1263_),
    .A(net1206),
    .B(_1262_));
 sg13g2_o21ai_1 _5170_ (.B1(_1242_),
    .Y(_1264_),
    .A1(_3192_),
    .A2(_0543_));
 sg13g2_o21ai_1 _5171_ (.B1(_1264_),
    .Y(_1265_),
    .A1(_3181_),
    .A2(_0315_));
 sg13g2_o21ai_1 _5172_ (.B1(_1263_),
    .Y(_1266_),
    .A1(net1207),
    .A2(_1265_));
 sg13g2_nor2_1 _5173_ (.A(net1123),
    .B(_1266_),
    .Y(_1267_));
 sg13g2_nand3_1 _5174_ (.B(net1282),
    .C(_3188_),
    .A(net1300),
    .Y(_1268_));
 sg13g2_a21oi_2 _5175_ (.B1(_1267_),
    .Y(_1269_),
    .A2(_1268_),
    .A1(net1126));
 sg13g2_nand2_1 _5176_ (.Y(_1270_),
    .A(net1117),
    .B(_1269_));
 sg13g2_a21oi_1 _5177_ (.A1(net1115),
    .A2(_1259_),
    .Y(_1271_),
    .B1(_0908_));
 sg13g2_nor2_1 _5178_ (.A(net1401),
    .B(_1253_),
    .Y(_1272_));
 sg13g2_o21ai_1 _5179_ (.B1(_1248_),
    .Y(_1273_),
    .A1(_1242_),
    .A2(_1244_));
 sg13g2_a21oi_1 _5180_ (.A1(net1400),
    .A2(_1273_),
    .Y(_1274_),
    .B1(_1272_));
 sg13g2_nor2_1 _5181_ (.A(net1123),
    .B(_1274_),
    .Y(_1275_));
 sg13g2_a21oi_2 _5182_ (.B1(_1275_),
    .Y(_1276_),
    .A2(_1256_),
    .A1(net1126));
 sg13g2_a21oi_1 _5183_ (.A1(net1213),
    .A2(_3181_),
    .Y(_1277_),
    .B1(_1242_));
 sg13g2_nor2_1 _5184_ (.A(_1260_),
    .B(_1277_),
    .Y(_1278_));
 sg13g2_nor2_1 _5185_ (.A(net1399),
    .B(_1278_),
    .Y(_1279_));
 sg13g2_a21oi_1 _5186_ (.A1(net1400),
    .A2(_1268_),
    .Y(_1280_),
    .B1(_1279_));
 sg13g2_nor2_1 _5187_ (.A(net1124),
    .B(_1280_),
    .Y(_1281_));
 sg13g2_a21oi_1 _5188_ (.A1(_0549_),
    .A2(_1243_),
    .Y(_1282_),
    .B1(_1247_));
 sg13g2_nand2_1 _5189_ (.Y(_1283_),
    .A(_1261_),
    .B(_1264_));
 sg13g2_nor2_1 _5190_ (.A(net1205),
    .B(_1283_),
    .Y(_1284_));
 sg13g2_a21oi_1 _5191_ (.A1(net1205),
    .A2(_1282_),
    .Y(_1285_),
    .B1(_1284_));
 sg13g2_a21oi_2 _5192_ (.B1(_1281_),
    .Y(_1286_),
    .A2(_1285_),
    .A1(net1123));
 sg13g2_mux2_1 _5193_ (.A0(_1276_),
    .A1(_1286_),
    .S(net1115),
    .X(_1287_));
 sg13g2_o21ai_1 _5194_ (.B1(\aliens_alive[38] ),
    .Y(_1288_),
    .A1(_0909_),
    .A2(_1287_));
 sg13g2_a21oi_1 _5195_ (.A1(_1270_),
    .A2(_1271_),
    .Y(_1289_),
    .B1(_1288_));
 sg13g2_and2_1 _5196_ (.A(net1115),
    .B(_1269_),
    .X(_1290_));
 sg13g2_a21oi_1 _5197_ (.A1(net1118),
    .A2(_1259_),
    .Y(_1291_),
    .B1(_1290_));
 sg13g2_mux2_1 _5198_ (.A0(_1276_),
    .A1(_1286_),
    .S(net1118),
    .X(_1292_));
 sg13g2_o21ai_1 _5199_ (.B1(\aliens_alive[34] ),
    .Y(_1293_),
    .A1(_0958_),
    .A2(_1292_));
 sg13g2_a21oi_1 _5200_ (.A1(_0958_),
    .A2(_1291_),
    .Y(_1294_),
    .B1(_1293_));
 sg13g2_a21oi_1 _5201_ (.A1(net1207),
    .A2(_1273_),
    .Y(_1295_),
    .B1(_1254_));
 sg13g2_nand2_1 _5202_ (.Y(_1296_),
    .A(net1106),
    .B(_1256_));
 sg13g2_o21ai_1 _5203_ (.B1(_1296_),
    .Y(_1297_),
    .A1(net1106),
    .A2(_1295_));
 sg13g2_nand2_1 _5204_ (.Y(_1298_),
    .A(net1399),
    .B(_1278_));
 sg13g2_o21ai_1 _5205_ (.B1(_1298_),
    .Y(_1299_),
    .A1(net1399),
    .A2(_1268_));
 sg13g2_nor2_1 _5206_ (.A(net1399),
    .B(_1283_),
    .Y(_1300_));
 sg13g2_a21oi_1 _5207_ (.A1(net1399),
    .A2(_1282_),
    .Y(_1301_),
    .B1(_1300_));
 sg13g2_nor2_1 _5208_ (.A(net1102),
    .B(_1299_),
    .Y(_1302_));
 sg13g2_a21oi_2 _5209_ (.B1(_1302_),
    .Y(_1303_),
    .A2(_1301_),
    .A1(net1103));
 sg13g2_o21ai_1 _5210_ (.B1(_0706_),
    .Y(_1304_),
    .A1(net1084),
    .A2(_1303_));
 sg13g2_a21oi_1 _5211_ (.A1(net1085),
    .A2(_1297_),
    .Y(_1305_),
    .B1(_1304_));
 sg13g2_nand2_1 _5212_ (.Y(_1306_),
    .A(net1206),
    .B(_1245_));
 sg13g2_o21ai_1 _5213_ (.B1(_1306_),
    .Y(_1307_),
    .A1(net1206),
    .A2(_1249_));
 sg13g2_a21oi_1 _5214_ (.A1(net1400),
    .A2(_1256_),
    .Y(_1308_),
    .B1(_1272_));
 sg13g2_nor2_1 _5215_ (.A(net1103),
    .B(_1308_),
    .Y(_1309_));
 sg13g2_a21oi_1 _5216_ (.A1(net1105),
    .A2(_1307_),
    .Y(_1310_),
    .B1(_1309_));
 sg13g2_nand2_1 _5217_ (.Y(_1311_),
    .A(net1401),
    .B(_1262_));
 sg13g2_o21ai_1 _5218_ (.B1(_1311_),
    .Y(_1312_),
    .A1(net1401),
    .A2(_1265_));
 sg13g2_nand2_1 _5219_ (.Y(_1313_),
    .A(net1106),
    .B(_1268_));
 sg13g2_o21ai_1 _5220_ (.B1(_1313_),
    .Y(_1314_),
    .A1(net1106),
    .A2(_1312_));
 sg13g2_a21oi_1 _5221_ (.A1(net1084),
    .A2(_1314_),
    .Y(_1315_),
    .B1(_0706_));
 sg13g2_o21ai_1 _5222_ (.B1(_1315_),
    .Y(_1316_),
    .A1(net1084),
    .A2(_1310_));
 sg13g2_nand2b_1 _5223_ (.Y(_1317_),
    .B(_1316_),
    .A_N(_1305_));
 sg13g2_nand3_1 _5224_ (.B(_0705_),
    .C(_1317_),
    .A(\aliens_alive[35] ),
    .Y(_1318_));
 sg13g2_nand2_1 _5225_ (.Y(_1319_),
    .A(_0650_),
    .B(_1297_));
 sg13g2_a21oi_1 _5226_ (.A1(_0651_),
    .A2(_1314_),
    .Y(_1320_),
    .B1(net1084));
 sg13g2_mux2_1 _5227_ (.A0(_1303_),
    .A1(_1310_),
    .S(_0651_),
    .X(_1321_));
 sg13g2_a22oi_1 _5228_ (.Y(_1322_),
    .B1(_1321_),
    .B2(net1085),
    .A2(_1320_),
    .A1(_1319_));
 sg13g2_nand3b_1 _5229_ (.B(_0640_),
    .C(\aliens_alive[39] ),
    .Y(_1323_),
    .A_N(_1322_));
 sg13g2_nand2_1 _5230_ (.Y(_1324_),
    .A(net1124),
    .B(_1274_));
 sg13g2_o21ai_1 _5231_ (.B1(_1324_),
    .Y(_1325_),
    .A1(net1123),
    .A2(_1256_));
 sg13g2_nand2_1 _5232_ (.Y(_1326_),
    .A(net1124),
    .B(_1280_));
 sg13g2_o21ai_1 _5233_ (.B1(_1326_),
    .Y(_1327_),
    .A1(net1123),
    .A2(_1285_));
 sg13g2_nand2_1 _5234_ (.Y(_1328_),
    .A(net1123),
    .B(_1266_));
 sg13g2_o21ai_1 _5235_ (.B1(_1328_),
    .Y(_1329_),
    .A1(net1126),
    .A2(_1268_));
 sg13g2_nand2_1 _5236_ (.Y(_1330_),
    .A(net1123),
    .B(_1257_));
 sg13g2_o21ai_1 _5237_ (.B1(_1330_),
    .Y(_1331_),
    .A1(net1126),
    .A2(_1250_));
 sg13g2_mux4_1 _5238_ (.S0(_0528_),
    .A0(_1329_),
    .A1(_1331_),
    .A2(_1325_),
    .A3(_1327_),
    .S1(_0558_),
    .X(_1332_));
 sg13g2_nand3_1 _5239_ (.B(_0527_),
    .C(_1332_),
    .A(\aliens_alive[36] ),
    .Y(_1333_));
 sg13g2_nand3_1 _5240_ (.B(_1323_),
    .C(_1333_),
    .A(_1318_),
    .Y(_1334_));
 sg13g2_a221oi_1 _5241_ (.B2(_0956_),
    .C1(_1334_),
    .B1(_1294_),
    .A1(_0901_),
    .Y(_1335_),
    .A2(_1289_));
 sg13g2_nor2b_1 _5242_ (.A(_1335_),
    .B_N(_1241_),
    .Y(_1336_));
 sg13g2_nor2_1 _5243_ (.A(net1105),
    .B(_1256_),
    .Y(_1337_));
 sg13g2_a21oi_1 _5244_ (.A1(net1105),
    .A2(_1295_),
    .Y(_1338_),
    .B1(_1337_));
 sg13g2_and2_1 _5245_ (.A(net1121),
    .B(_1338_),
    .X(_1339_));
 sg13g2_nor2_1 _5246_ (.A(net1102),
    .B(_1301_),
    .Y(_1340_));
 sg13g2_a21oi_1 _5247_ (.A1(net1103),
    .A2(_1299_),
    .Y(_1341_),
    .B1(_1340_));
 sg13g2_nand2_1 _5248_ (.Y(_1342_),
    .A(net1120),
    .B(_1341_));
 sg13g2_nand2_1 _5249_ (.Y(_1343_),
    .A(_0864_),
    .B(_1342_));
 sg13g2_nand2_1 _5250_ (.Y(_1344_),
    .A(net1103),
    .B(_1308_));
 sg13g2_o21ai_1 _5251_ (.B1(_1344_),
    .Y(_1345_),
    .A1(net1104),
    .A2(_1307_));
 sg13g2_nor2_1 _5252_ (.A(net1105),
    .B(_1268_),
    .Y(_1346_));
 sg13g2_a21oi_1 _5253_ (.A1(net1105),
    .A2(_1312_),
    .Y(_1347_),
    .B1(_1346_));
 sg13g2_a21oi_1 _5254_ (.A1(net1121),
    .A2(_1347_),
    .Y(_1348_),
    .B1(_0864_));
 sg13g2_o21ai_1 _5255_ (.B1(_1348_),
    .Y(_1349_),
    .A1(net1121),
    .A2(_1345_));
 sg13g2_o21ai_1 _5256_ (.B1(_1349_),
    .Y(_1350_),
    .A1(_1339_),
    .A2(_1343_));
 sg13g2_nand4_1 _5257_ (.B(_0863_),
    .C(_1241_),
    .A(\aliens_alive[37] ),
    .Y(_1351_),
    .D(_1350_));
 sg13g2_nand2_1 _5258_ (.Y(_1352_),
    .A(net1120),
    .B(_1338_));
 sg13g2_nand2_1 _5259_ (.Y(_1353_),
    .A(net1121),
    .B(_1341_));
 sg13g2_nand3_1 _5260_ (.B(_1352_),
    .C(_1353_),
    .A(_0804_),
    .Y(_1354_));
 sg13g2_a21oi_1 _5261_ (.A1(net1120),
    .A2(_1347_),
    .Y(_1355_),
    .B1(_0804_));
 sg13g2_o21ai_1 _5262_ (.B1(_1355_),
    .Y(_1356_),
    .A1(net1120),
    .A2(_1345_));
 sg13g2_nand2_1 _5263_ (.Y(_1357_),
    .A(_1354_),
    .B(_1356_));
 sg13g2_nand4_1 _5264_ (.B(_0798_),
    .C(_1241_),
    .A(\aliens_alive[33] ),
    .Y(_1358_),
    .D(_1357_));
 sg13g2_mux4_1 _5265_ (.S0(_0529_),
    .A0(_1325_),
    .A1(_1327_),
    .A2(_1329_),
    .A3(_1331_),
    .S1(_0743_),
    .X(_1359_));
 sg13g2_nand4_1 _5266_ (.B(_0742_),
    .C(_1241_),
    .A(\aliens_alive[32] ),
    .Y(_1360_),
    .D(_1359_));
 sg13g2_nand3_1 _5267_ (.B(_1358_),
    .C(_1360_),
    .A(_1351_),
    .Y(_1361_));
 sg13g2_nor3_2 _5268_ (.A(_1232_),
    .B(_1336_),
    .C(_1361_),
    .Y(_1362_));
 sg13g2_nand2_1 _5269_ (.Y(_1363_),
    .A(_1114_),
    .B(_1362_));
 sg13g2_a21oi_1 _5270_ (.A1(_0478_),
    .A2(_1363_),
    .Y(_1364_),
    .B1(_3233_));
 sg13g2_nor3_1 _5271_ (.A(net1204),
    .B(_0305_),
    .C(_1121_),
    .Y(_1365_));
 sg13g2_nand2_1 _5272_ (.Y(_1366_),
    .A(_3288_),
    .B(_0533_));
 sg13g2_o21ai_1 _5273_ (.B1(_0533_),
    .Y(_1367_),
    .A1(_3288_),
    .A2(_0306_));
 sg13g2_a21o_1 _5274_ (.A2(_1367_),
    .A1(net1204),
    .B1(_1365_),
    .X(_1368_));
 sg13g2_nor3_1 _5275_ (.A(net1220),
    .B(net1407),
    .C(_3288_),
    .Y(_1369_));
 sg13g2_nand2_2 _5276_ (.Y(_1370_),
    .A(net1389),
    .B(net1198));
 sg13g2_nor4_1 _5277_ (.A(_0044_),
    .B(_0533_),
    .C(_1369_),
    .D(_1370_),
    .Y(_1371_));
 sg13g2_a221oi_1 _5278_ (.B2(net1190),
    .C1(_1371_),
    .B1(_1368_),
    .A1(_3073_),
    .Y(_1372_),
    .A2(_1366_));
 sg13g2_nand2_1 _5279_ (.Y(_1373_),
    .A(net1204),
    .B(net1190));
 sg13g2_nand4_1 _5280_ (.B(_3070_),
    .C(_3210_),
    .A(net1387),
    .Y(_1374_),
    .D(_1373_));
 sg13g2_o21ai_1 _5281_ (.B1(_1374_),
    .Y(_1375_),
    .A1(net1189),
    .A2(_1372_));
 sg13g2_o21ai_1 _5282_ (.B1(_0015_),
    .Y(_1376_),
    .A1(_3050_),
    .A2(_0395_));
 sg13g2_nand3_1 _5283_ (.B(_2907_),
    .C(_1230_),
    .A(net1223),
    .Y(_1377_));
 sg13g2_nor3_1 _5284_ (.A(_0355_),
    .B(_0435_),
    .C(_1377_),
    .Y(_1378_));
 sg13g2_o21ai_1 _5285_ (.B1(_1378_),
    .Y(_1379_),
    .A1(net1268),
    .A2(_1376_));
 sg13g2_a21oi_1 _5286_ (.A1(net1268),
    .A2(_1376_),
    .Y(_1380_),
    .B1(_1379_));
 sg13g2_nand3_1 _5287_ (.B(_1375_),
    .C(_1380_),
    .A(_0353_),
    .Y(_1381_));
 sg13g2_inv_1 _5288_ (.Y(_1382_),
    .A(_1381_));
 sg13g2_nor2_1 _5289_ (.A(_1364_),
    .B(_1382_),
    .Y(_1383_));
 sg13g2_nor2_1 _5290_ (.A(net1223),
    .B(net1280),
    .Y(_1384_));
 sg13g2_and2_1 _5291_ (.A(net1193),
    .B(_1384_),
    .X(_1385_));
 sg13g2_a21oi_1 _5292_ (.A1(net1187),
    .A2(_1385_),
    .Y(_1386_),
    .B1(_0013_));
 sg13g2_a21oi_1 _5293_ (.A1(_0541_),
    .A2(_1385_),
    .Y(_1387_),
    .B1(_1386_));
 sg13g2_nand2_1 _5294_ (.Y(_1388_),
    .A(_3042_),
    .B(_1387_));
 sg13g2_nor4_2 _5295_ (.A(net1264),
    .B(net1268),
    .C(_0963_),
    .Y(_1389_),
    .D(_1235_));
 sg13g2_or4_1 _5296_ (.A(net1357),
    .B(net1353),
    .C(_1388_),
    .D(_1389_),
    .X(_1390_));
 sg13g2_nand2_1 _5297_ (.Y(_1391_),
    .A(net1394),
    .B(net1387));
 sg13g2_nor3_2 _5298_ (.A(net1198),
    .B(net1196),
    .C(net1190),
    .Y(_1392_));
 sg13g2_o21ai_1 _5299_ (.B1(net1369),
    .Y(_1393_),
    .A1(net1375),
    .A2(_1392_));
 sg13g2_nand2_1 _5300_ (.Y(_1394_),
    .A(_0348_),
    .B(_1370_));
 sg13g2_nor4_1 _5301_ (.A(net1362),
    .B(_1390_),
    .C(_1393_),
    .D(_1394_),
    .Y(_1395_));
 sg13g2_nor3_1 _5302_ (.A(net1271),
    .B(_2906_),
    .C(_0434_),
    .Y(_1396_));
 sg13g2_nand4_1 _5303_ (.B(_2842_),
    .C(_0963_),
    .A(net1225),
    .Y(_1397_),
    .D(_1396_));
 sg13g2_nand2b_1 _5304_ (.Y(_1398_),
    .B(_3042_),
    .A_N(_0013_));
 sg13g2_o21ai_1 _5305_ (.B1(_1397_),
    .Y(_1399_),
    .A1(_0963_),
    .A2(_1398_));
 sg13g2_nand2b_2 _5306_ (.Y(_1400_),
    .B(_1399_),
    .A_N(_0967_));
 sg13g2_nor2_1 _5307_ (.A(_0452_),
    .B(_1400_),
    .Y(_1401_));
 sg13g2_nor2_1 _5308_ (.A(_0982_),
    .B(_1400_),
    .Y(_1402_));
 sg13g2_a21oi_2 _5309_ (.B1(_1400_),
    .Y(_1403_),
    .A2(_0982_),
    .A1(_0452_));
 sg13g2_inv_1 _5310_ (.Y(_1404_),
    .A(_1403_));
 sg13g2_and2_1 _5311_ (.A(net1303),
    .B(net1305),
    .X(_1405_));
 sg13g2_nand2_2 _5312_ (.Y(_1406_),
    .A(net1304),
    .B(\draw_score_inst.score[8] ));
 sg13g2_nand3b_1 _5313_ (.B(net1303),
    .C(net1305),
    .Y(_1407_),
    .A_N(net1306));
 sg13g2_xnor2_1 _5314_ (.Y(_1408_),
    .A(_0020_),
    .B(_1407_));
 sg13g2_nor2_1 _5315_ (.A(net1306),
    .B(net1305),
    .Y(_1409_));
 sg13g2_o21ai_1 _5316_ (.B1(net1303),
    .Y(_1410_),
    .A1(_0019_),
    .A2(_1409_));
 sg13g2_inv_1 _5317_ (.Y(_1411_),
    .A(_1410_));
 sg13g2_nor2b_1 _5318_ (.A(_1409_),
    .B_N(net1303),
    .Y(_1412_));
 sg13g2_o21ai_1 _5319_ (.B1(net1303),
    .Y(_1413_),
    .A1(net1306),
    .A2(net1305));
 sg13g2_a22oi_1 _5320_ (.Y(_1414_),
    .B1(_1413_),
    .B2(_2911_),
    .A2(_1405_),
    .A1(_2902_));
 sg13g2_a221oi_1 _5321_ (.B2(_2911_),
    .C1(_2912_),
    .B1(_1413_),
    .A1(_2902_),
    .Y(_1415_),
    .A2(_1405_));
 sg13g2_nor2_1 _5322_ (.A(_1408_),
    .B(_1415_),
    .Y(_1416_));
 sg13g2_or2_1 _5323_ (.X(_1417_),
    .B(_1415_),
    .A(_1408_));
 sg13g2_nor2_1 _5324_ (.A(_1410_),
    .B(_1417_),
    .Y(_1418_));
 sg13g2_nor2_1 _5325_ (.A(_1411_),
    .B(_1416_),
    .Y(_1419_));
 sg13g2_o21ai_1 _5326_ (.B1(_1410_),
    .Y(_1420_),
    .A1(_1408_),
    .A2(_1415_));
 sg13g2_xnor2_1 _5327_ (.Y(_1421_),
    .A(_2912_),
    .B(_1420_));
 sg13g2_xnor2_1 _5328_ (.Y(_1422_),
    .A(_0022_),
    .B(_1420_));
 sg13g2_nor2_1 _5329_ (.A(_2913_),
    .B(_1422_),
    .Y(_1423_));
 sg13g2_nand2_1 _5330_ (.Y(_1424_),
    .A(_0023_),
    .B(_1421_));
 sg13g2_a21oi_1 _5331_ (.A1(_0022_),
    .A2(_1420_),
    .Y(_1425_),
    .B1(_1414_));
 sg13g2_a21o_1 _5332_ (.A2(_1415_),
    .A1(_1411_),
    .B1(_1425_),
    .X(_1426_));
 sg13g2_o21ai_1 _5333_ (.B1(_1408_),
    .Y(_1427_),
    .A1(_1410_),
    .A2(_1415_));
 sg13g2_and2_1 _5334_ (.A(_1417_),
    .B(_1427_),
    .X(_1428_));
 sg13g2_a221oi_1 _5335_ (.B2(_1426_),
    .C1(_1428_),
    .B1(_1424_),
    .A1(_1411_),
    .Y(_1429_),
    .A2(_1416_));
 sg13g2_xnor2_1 _5336_ (.Y(_1430_),
    .A(_0023_),
    .B(_1429_));
 sg13g2_o21ai_1 _5337_ (.B1(_1422_),
    .Y(_1431_),
    .A1(_2913_),
    .A2(_1429_));
 sg13g2_nand3b_1 _5338_ (.B(_1421_),
    .C(_0023_),
    .Y(_1432_),
    .A_N(_1429_));
 sg13g2_and2_1 _5339_ (.A(_1431_),
    .B(_1432_),
    .X(_1433_));
 sg13g2_a22oi_1 _5340_ (.Y(_1434_),
    .B1(_1431_),
    .B2(_1432_),
    .A2(_1430_),
    .A1(_2901_));
 sg13g2_mux2_1 _5341_ (.A0(_1426_),
    .A1(_1428_),
    .S(_1424_),
    .X(_1435_));
 sg13g2_nor2_1 _5342_ (.A(_1423_),
    .B(_1429_),
    .Y(_1436_));
 sg13g2_mux2_1 _5343_ (.A0(_1436_),
    .A1(_1423_),
    .S(_1426_),
    .X(_1437_));
 sg13g2_nand3_1 _5344_ (.B(_1426_),
    .C(_1428_),
    .A(_1424_),
    .Y(_1438_));
 sg13g2_nand2b_1 _5345_ (.Y(_1439_),
    .B(_1438_),
    .A_N(_1418_));
 sg13g2_nor2_2 _5346_ (.A(_1418_),
    .B(_1435_),
    .Y(_1440_));
 sg13g2_or2_1 _5347_ (.X(_1441_),
    .B(_1435_),
    .A(_1418_));
 sg13g2_nor2_1 _5348_ (.A(net1080),
    .B(_1441_),
    .Y(_1442_));
 sg13g2_nand2b_1 _5349_ (.Y(_1443_),
    .B(_1440_),
    .A_N(net1080));
 sg13g2_o21ai_1 _5350_ (.B1(_2901_),
    .Y(_1444_),
    .A1(_1434_),
    .A2(_1441_));
 sg13g2_nand3b_1 _5351_ (.B(_1440_),
    .C(\draw_score_inst.score[4] ),
    .Y(_1445_),
    .A_N(net1080));
 sg13g2_and2_1 _5352_ (.A(_1444_),
    .B(_1445_),
    .X(_1446_));
 sg13g2_nand3_1 _5353_ (.B(_1444_),
    .C(_1445_),
    .A(_2898_),
    .Y(_1447_));
 sg13g2_o21ai_1 _5354_ (.B1(_0024_),
    .Y(_1448_),
    .A1(net1080),
    .A2(_1441_));
 sg13g2_xor2_1 _5355_ (.B(_1448_),
    .A(_1430_),
    .X(_1449_));
 sg13g2_and3_1 _5356_ (.X(_1450_),
    .A(_2901_),
    .B(_1421_),
    .C(_1430_));
 sg13g2_nor3_1 _5357_ (.A(net1080),
    .B(_1440_),
    .C(_1450_),
    .Y(_1451_));
 sg13g2_nor3_1 _5358_ (.A(_1433_),
    .B(net1080),
    .C(_1441_),
    .Y(_1452_));
 sg13g2_a21o_1 _5359_ (.A2(_1437_),
    .A1(net1080),
    .B1(_1439_),
    .X(_1453_));
 sg13g2_nor3_1 _5360_ (.A(_1451_),
    .B(_1452_),
    .C(_1453_),
    .Y(_1454_));
 sg13g2_or3_1 _5361_ (.A(_1451_),
    .B(_1452_),
    .C(_1453_),
    .X(_1455_));
 sg13g2_a21o_2 _5362_ (.A2(_1449_),
    .A1(_1447_),
    .B1(_1455_),
    .X(_1456_));
 sg13g2_xor2_1 _5363_ (.B(_1456_),
    .A(_0018_),
    .X(_1457_));
 sg13g2_nand2_1 _5364_ (.Y(_1458_),
    .A(_0026_),
    .B(_1457_));
 sg13g2_a21o_1 _5365_ (.A2(_1456_),
    .A1(_2898_),
    .B1(_1446_),
    .X(_1459_));
 sg13g2_nand2b_1 _5366_ (.Y(_1460_),
    .B(_1455_),
    .A_N(_1447_));
 sg13g2_a22oi_1 _5367_ (.Y(_1461_),
    .B1(_1459_),
    .B2(_1460_),
    .A2(_1457_),
    .A1(_0026_));
 sg13g2_a21oi_1 _5368_ (.A1(_1447_),
    .A2(_1449_),
    .Y(_1462_),
    .B1(_1453_));
 sg13g2_nor2_1 _5369_ (.A(_1454_),
    .B(_1462_),
    .Y(_1463_));
 sg13g2_a21oi_1 _5370_ (.A1(_1447_),
    .A2(_1455_),
    .Y(_1464_),
    .B1(_1449_));
 sg13g2_a21o_1 _5371_ (.A2(_1449_),
    .A1(_1447_),
    .B1(_1464_),
    .X(_1465_));
 sg13g2_nand2b_2 _5372_ (.Y(_1466_),
    .B(_1465_),
    .A_N(_1463_));
 sg13g2_nor2_1 _5373_ (.A(_1461_),
    .B(_1466_),
    .Y(_1467_));
 sg13g2_o21ai_1 _5374_ (.B1(_2899_),
    .Y(_1468_),
    .A1(_1461_),
    .A2(_1466_));
 sg13g2_or3_1 _5375_ (.A(_2899_),
    .B(_1461_),
    .C(_1466_),
    .X(_1469_));
 sg13g2_and2_1 _5376_ (.A(_1468_),
    .B(_1469_),
    .X(_1470_));
 sg13g2_and3_1 _5377_ (.X(_1471_),
    .A(_0025_),
    .B(_1468_),
    .C(_1469_));
 sg13g2_nand3_1 _5378_ (.B(_1468_),
    .C(_1469_),
    .A(_0025_),
    .Y(_1472_));
 sg13g2_xor2_1 _5379_ (.B(_1468_),
    .A(_1457_),
    .X(_1473_));
 sg13g2_xnor2_1 _5380_ (.Y(_1474_),
    .A(_1457_),
    .B(_1468_));
 sg13g2_nand2_1 _5381_ (.Y(_1475_),
    .A(_1472_),
    .B(_1473_));
 sg13g2_a21oi_1 _5382_ (.A1(_0026_),
    .A2(_1457_),
    .Y(_1476_),
    .B1(_1465_));
 sg13g2_a21oi_1 _5383_ (.A1(_1459_),
    .A2(_1460_),
    .Y(_1477_),
    .B1(_1458_));
 sg13g2_nor3_1 _5384_ (.A(_1463_),
    .B(_1476_),
    .C(_1477_),
    .Y(_1478_));
 sg13g2_or3_1 _5385_ (.A(_1463_),
    .B(_1476_),
    .C(_1477_),
    .X(_1479_));
 sg13g2_a21oi_1 _5386_ (.A1(_1472_),
    .A2(_1473_),
    .Y(_1480_),
    .B1(_1479_));
 sg13g2_o21ai_1 _5387_ (.B1(_1478_),
    .Y(_1481_),
    .A1(_1471_),
    .A2(_1474_));
 sg13g2_a21oi_1 _5388_ (.A1(_1474_),
    .A2(_1478_),
    .Y(_1482_),
    .B1(_1471_));
 sg13g2_or2_1 _5389_ (.X(_1483_),
    .B(_1470_),
    .A(_0025_));
 sg13g2_a22oi_1 _5390_ (.Y(_1484_),
    .B1(_1482_),
    .B2(_1483_),
    .A2(_1480_),
    .A1(_1470_));
 sg13g2_o21ai_1 _5391_ (.B1(_1475_),
    .Y(_1485_),
    .A1(_1473_),
    .A2(_1482_));
 sg13g2_xnor2_1 _5392_ (.Y(_1486_),
    .A(\draw_score_inst.score[1] ),
    .B(_1481_));
 sg13g2_xnor2_1 _5393_ (.Y(_1487_),
    .A(\draw_score_inst.score[1] ),
    .B(_1480_));
 sg13g2_nand2_1 _5394_ (.Y(_1488_),
    .A(_1485_),
    .B(_1486_));
 sg13g2_nand3_1 _5395_ (.B(_1485_),
    .C(_1486_),
    .A(_1484_),
    .Y(_1489_));
 sg13g2_nand2_1 _5396_ (.Y(_1490_),
    .A(_1403_),
    .B(_1489_));
 sg13g2_or2_1 _5397_ (.X(_1491_),
    .B(_1400_),
    .A(_0540_));
 sg13g2_nor3_2 _5398_ (.A(_3181_),
    .B(_1133_),
    .C(_1491_),
    .Y(_1492_));
 sg13g2_inv_1 _5399_ (.Y(_1493_),
    .A(_1492_));
 sg13g2_o21ai_1 _5400_ (.B1(_1492_),
    .Y(_1494_),
    .A1(_1484_),
    .A2(_1488_));
 sg13g2_xnor2_1 _5401_ (.Y(_1495_),
    .A(net1202),
    .B(_1393_));
 sg13g2_xnor2_1 _5402_ (.Y(_1496_),
    .A(net1374),
    .B(_1392_));
 sg13g2_nand3_1 _5403_ (.B(_2877_),
    .C(_1496_),
    .A(_2875_),
    .Y(_1497_));
 sg13g2_and3_1 _5404_ (.X(_1498_),
    .A(net1196),
    .B(net1192),
    .C(_1391_));
 sg13g2_nor3_1 _5405_ (.A(net1368),
    .B(_1495_),
    .C(_1497_),
    .Y(_1499_));
 sg13g2_o21ai_1 _5406_ (.B1(_1499_),
    .Y(_1500_),
    .A1(_1392_),
    .A2(_1498_));
 sg13g2_nand2_1 _5407_ (.Y(_1501_),
    .A(net1198),
    .B(net1190));
 sg13g2_a221oi_1 _5408_ (.B2(net1192),
    .C1(_1500_),
    .B1(_1501_),
    .A1(_1490_),
    .Y(_1502_),
    .A2(_1494_));
 sg13g2_nor2_1 _5409_ (.A(_1134_),
    .B(_1491_),
    .Y(_1503_));
 sg13g2_nor3_2 _5410_ (.A(_0451_),
    .B(_1134_),
    .C(_1491_),
    .Y(_1504_));
 sg13g2_nand3b_1 _5411_ (.B(_1485_),
    .C(_1487_),
    .Y(_1505_),
    .A_N(_1484_));
 sg13g2_nor3_2 _5412_ (.A(net1278),
    .B(_1400_),
    .C(_1503_),
    .Y(_1506_));
 sg13g2_inv_1 _5413_ (.Y(_1507_),
    .A(_1506_));
 sg13g2_a22oi_1 _5414_ (.Y(_1508_),
    .B1(_1506_),
    .B2(_1489_),
    .A2(_1505_),
    .A1(_1504_));
 sg13g2_nor4_1 _5415_ (.A(net1389),
    .B(_1391_),
    .C(_1500_),
    .D(_1508_),
    .Y(_1509_));
 sg13g2_nand3_1 _5416_ (.B(_1485_),
    .C(_1487_),
    .A(_1484_),
    .Y(_1510_));
 sg13g2_a22oi_1 _5417_ (.Y(_1511_),
    .B1(_1510_),
    .B2(_1504_),
    .A2(_1506_),
    .A1(_1505_));
 sg13g2_nand3_1 _5418_ (.B(_1391_),
    .C(_1501_),
    .A(net1192),
    .Y(_1512_));
 sg13g2_nor3_1 _5419_ (.A(net1387),
    .B(net1380),
    .C(net1375),
    .Y(_1513_));
 sg13g2_a21oi_1 _5420_ (.A1(_3070_),
    .A2(_1513_),
    .Y(_1514_),
    .B1(net1194));
 sg13g2_o21ai_1 _5421_ (.B1(_3076_),
    .Y(_1515_),
    .A1(net1192),
    .A2(_3089_));
 sg13g2_nor3_1 _5422_ (.A(net1407),
    .B(_2879_),
    .C(_1370_),
    .Y(_1516_));
 sg13g2_nor2_1 _5423_ (.A(net1362),
    .B(_1516_),
    .Y(_1517_));
 sg13g2_nand2_1 _5424_ (.Y(_1518_),
    .A(_1515_),
    .B(_1517_));
 sg13g2_nor3_1 _5425_ (.A(_1390_),
    .B(_1514_),
    .C(_1518_),
    .Y(_1519_));
 sg13g2_a21oi_1 _5426_ (.A1(_1419_),
    .A2(_1429_),
    .Y(_1520_),
    .B1(_1413_));
 sg13g2_a21oi_1 _5427_ (.A1(_1412_),
    .A2(_1429_),
    .Y(_1521_),
    .B1(_1419_));
 sg13g2_xor2_1 _5428_ (.B(_1520_),
    .A(_1429_),
    .X(_1522_));
 sg13g2_inv_1 _5429_ (.Y(_1523_),
    .A(_1522_));
 sg13g2_nand3b_1 _5430_ (.B(_1440_),
    .C(_1522_),
    .Y(_1524_),
    .A_N(net1080));
 sg13g2_nor2_1 _5431_ (.A(_1413_),
    .B(_1520_),
    .Y(_1525_));
 sg13g2_a21oi_1 _5432_ (.A1(_1521_),
    .A2(_1524_),
    .Y(_1526_),
    .B1(_1525_));
 sg13g2_xnor2_1 _5433_ (.Y(_1527_),
    .A(_1443_),
    .B(_1526_));
 sg13g2_nor2_1 _5434_ (.A(_1456_),
    .B(_1527_),
    .Y(_1528_));
 sg13g2_a21oi_1 _5435_ (.A1(_1442_),
    .A2(_1525_),
    .Y(_1529_),
    .B1(_1523_));
 sg13g2_nor4_1 _5436_ (.A(_1412_),
    .B(_1419_),
    .C(_1429_),
    .D(_1443_),
    .Y(_1530_));
 sg13g2_nor2_1 _5437_ (.A(_1529_),
    .B(_1530_),
    .Y(_1531_));
 sg13g2_o21ai_1 _5438_ (.B1(_1531_),
    .Y(_1532_),
    .A1(_1456_),
    .A2(_1527_));
 sg13g2_a21oi_1 _5439_ (.A1(_1524_),
    .A2(_1525_),
    .Y(_1533_),
    .B1(_1521_));
 sg13g2_a21o_1 _5440_ (.A2(_1524_),
    .A1(_1521_),
    .B1(_1533_),
    .X(_1534_));
 sg13g2_a21oi_2 _5441_ (.B1(_1456_),
    .Y(_1535_),
    .A2(_1534_),
    .A1(_1532_));
 sg13g2_and3_1 _5442_ (.X(_1536_),
    .A(_1456_),
    .B(_1532_),
    .C(_1534_));
 sg13g2_nor2_2 _5443_ (.A(_1535_),
    .B(_1536_),
    .Y(_1537_));
 sg13g2_nor4_2 _5444_ (.A(_1461_),
    .B(_1466_),
    .C(_1535_),
    .Y(_1538_),
    .D(_1536_));
 sg13g2_xnor2_1 _5445_ (.Y(_1539_),
    .A(_1527_),
    .B(_1535_));
 sg13g2_mux2_1 _5446_ (.A0(_1534_),
    .A1(_1522_),
    .S(_1528_),
    .X(_1540_));
 sg13g2_o21ai_1 _5447_ (.B1(_1540_),
    .Y(_1541_),
    .A1(_1538_),
    .A2(_1539_));
 sg13g2_nand2_1 _5448_ (.Y(_1542_),
    .A(_1467_),
    .B(_1541_));
 sg13g2_xnor2_1 _5449_ (.Y(_1543_),
    .A(_1467_),
    .B(_1541_));
 sg13g2_or2_1 _5450_ (.X(_1544_),
    .B(_1543_),
    .A(_1481_));
 sg13g2_xor2_1 _5451_ (.B(_1542_),
    .A(_1537_),
    .X(_1545_));
 sg13g2_nand2_1 _5452_ (.Y(_1546_),
    .A(_1481_),
    .B(_1543_));
 sg13g2_nand3_1 _5453_ (.B(_1545_),
    .C(_1546_),
    .A(_1544_),
    .Y(_1547_));
 sg13g2_nand4_1 _5454_ (.B(_1544_),
    .C(_1545_),
    .A(_1402_),
    .Y(_1548_),
    .D(_1546_));
 sg13g2_nor2b_1 _5455_ (.A(_1546_),
    .B_N(_1545_),
    .Y(_1549_));
 sg13g2_o21ai_1 _5456_ (.B1(_1539_),
    .Y(_1550_),
    .A1(_1538_),
    .A2(_1540_));
 sg13g2_o21ai_1 _5457_ (.B1(_1550_),
    .Y(_1551_),
    .A1(_1538_),
    .A2(_1539_));
 sg13g2_nor2b_1 _5458_ (.A(_1543_),
    .B_N(_1551_),
    .Y(_1552_));
 sg13g2_a21o_1 _5459_ (.A2(_1552_),
    .A1(_1537_),
    .B1(_1493_),
    .X(_1553_));
 sg13g2_nand3_1 _5460_ (.B(_1544_),
    .C(_1545_),
    .A(_1401_),
    .Y(_1554_));
 sg13g2_o21ai_1 _5461_ (.B1(_1554_),
    .Y(_1555_),
    .A1(_1549_),
    .A2(_1553_));
 sg13g2_a21o_1 _5462_ (.A2(_1552_),
    .A1(_1481_),
    .B1(_1404_),
    .X(_1556_));
 sg13g2_o21ai_1 _5463_ (.B1(_1548_),
    .Y(_1557_),
    .A1(_1545_),
    .A2(_1556_));
 sg13g2_nand3_1 _5464_ (.B(_2877_),
    .C(_0321_),
    .A(net1202),
    .Y(_1558_));
 sg13g2_xnor2_1 _5465_ (.Y(_1559_),
    .A(net1357),
    .B(_1515_));
 sg13g2_nor4_2 _5466_ (.A(_3087_),
    .B(_0346_),
    .C(_1558_),
    .Y(_1560_),
    .D(_1559_));
 sg13g2_inv_1 _5467_ (.Y(_1561_),
    .A(_1560_));
 sg13g2_nor2_1 _5468_ (.A(net1394),
    .B(net1192),
    .Y(_1562_));
 sg13g2_nor3_1 _5469_ (.A(_0305_),
    .B(_1561_),
    .C(_1562_),
    .Y(_1563_));
 sg13g2_o21ai_1 _5470_ (.B1(_1563_),
    .Y(_1564_),
    .A1(_1555_),
    .A2(_1557_));
 sg13g2_nor2_1 _5471_ (.A(_1481_),
    .B(_1545_),
    .Y(_1565_));
 sg13g2_a21oi_1 _5472_ (.A1(_1543_),
    .A2(_1565_),
    .Y(_1566_),
    .B1(_1507_));
 sg13g2_and2_1 _5473_ (.A(_1504_),
    .B(_1547_),
    .X(_1567_));
 sg13g2_nor2_1 _5474_ (.A(net1394),
    .B(_1370_),
    .Y(_1568_));
 sg13g2_and2_1 _5475_ (.A(_1560_),
    .B(_1568_),
    .X(_1569_));
 sg13g2_o21ai_1 _5476_ (.B1(_1569_),
    .Y(_1570_),
    .A1(_1566_),
    .A2(_1567_));
 sg13g2_o21ai_1 _5477_ (.B1(_1551_),
    .Y(_1571_),
    .A1(_1481_),
    .A2(_1543_));
 sg13g2_a21oi_1 _5478_ (.A1(_1545_),
    .A2(_1546_),
    .Y(_1572_),
    .B1(_1571_));
 sg13g2_nor2b_1 _5479_ (.A(_1572_),
    .B_N(_1504_),
    .Y(_1573_));
 sg13g2_nor2b_1 _5480_ (.A(_1537_),
    .B_N(_1552_),
    .Y(_1574_));
 sg13g2_nor3_1 _5481_ (.A(_1481_),
    .B(_1507_),
    .C(_1574_),
    .Y(_1575_));
 sg13g2_and2_1 _5482_ (.A(_1560_),
    .B(_1562_),
    .X(_1576_));
 sg13g2_o21ai_1 _5483_ (.B1(_1576_),
    .Y(_1577_),
    .A1(_1573_),
    .A2(_1575_));
 sg13g2_nand3_1 _5484_ (.B(net1190),
    .C(_0387_),
    .A(net1204),
    .Y(_1578_));
 sg13g2_a22oi_1 _5485_ (.Y(_1579_),
    .B1(_1578_),
    .B2(net1374),
    .A2(_0343_),
    .A1(net1375));
 sg13g2_a21oi_1 _5486_ (.A1(_3067_),
    .A2(_3068_),
    .Y(_1580_),
    .B1(net1375));
 sg13g2_nor4_1 _5487_ (.A(_3077_),
    .B(_1390_),
    .C(_1579_),
    .D(_1580_),
    .Y(_1581_));
 sg13g2_nor2_1 _5488_ (.A(net1307),
    .B(net1308),
    .Y(_1582_));
 sg13g2_nor3_1 _5489_ (.A(\draw_score_inst.score[5] ),
    .B(net1307),
    .C(net1308),
    .Y(_1583_));
 sg13g2_or3_1 _5490_ (.A(net1309),
    .B(net1306),
    .C(net1308),
    .X(_1584_));
 sg13g2_nor2_2 _5491_ (.A(_1406_),
    .B(_1583_),
    .Y(_1585_));
 sg13g2_nor3_2 _5492_ (.A(net1309),
    .B(_1406_),
    .C(_1582_),
    .Y(_1586_));
 sg13g2_a21oi_2 _5493_ (.B1(_0023_),
    .Y(_1587_),
    .A2(_1584_),
    .A1(_1405_));
 sg13g2_nor2_1 _5494_ (.A(_1586_),
    .B(_1587_),
    .Y(_1588_));
 sg13g2_nor2b_1 _5495_ (.A(\draw_score_inst.score[6] ),
    .B_N(_1586_),
    .Y(_1589_));
 sg13g2_xnor2_1 _5496_ (.Y(_1590_),
    .A(_2911_),
    .B(_1589_));
 sg13g2_nor3_1 _5497_ (.A(\draw_score_inst.score[4] ),
    .B(_1586_),
    .C(_1587_),
    .Y(_1591_));
 sg13g2_nor4_1 _5498_ (.A(\draw_score_inst.score[4] ),
    .B(_2912_),
    .C(_1586_),
    .D(_1587_),
    .Y(_1592_));
 sg13g2_nand2_1 _5499_ (.Y(_1593_),
    .A(_0022_),
    .B(_1591_));
 sg13g2_o21ai_1 _5500_ (.B1(_2910_),
    .Y(_1594_),
    .A1(_1406_),
    .A2(_1583_));
 sg13g2_nor4_2 _5501_ (.A(_0020_),
    .B(_0021_),
    .C(_1585_),
    .Y(_1595_),
    .D(_1592_));
 sg13g2_xnor2_1 _5502_ (.Y(_1596_),
    .A(_0019_),
    .B(_1585_));
 sg13g2_nor2_2 _5503_ (.A(_1595_),
    .B(_1596_),
    .Y(_1597_));
 sg13g2_o21ai_1 _5504_ (.B1(_0024_),
    .Y(_1598_),
    .A1(_1595_),
    .A2(_1596_));
 sg13g2_xnor2_1 _5505_ (.Y(_1599_),
    .A(_1588_),
    .B(_1598_));
 sg13g2_xnor2_1 _5506_ (.Y(_1600_),
    .A(_2901_),
    .B(_1597_));
 sg13g2_nand3_1 _5507_ (.B(_1599_),
    .C(_1600_),
    .A(_2898_),
    .Y(_1601_));
 sg13g2_xnor2_1 _5508_ (.Y(_1602_),
    .A(_0022_),
    .B(_1586_));
 sg13g2_o21ai_1 _5509_ (.B1(_1591_),
    .Y(_1603_),
    .A1(_1595_),
    .A2(_1596_));
 sg13g2_xnor2_1 _5510_ (.Y(_1604_),
    .A(_1602_),
    .B(_1603_));
 sg13g2_inv_1 _5511_ (.Y(_1605_),
    .A(_1604_));
 sg13g2_o21ai_1 _5512_ (.B1(_1593_),
    .Y(_1606_),
    .A1(_1595_),
    .A2(_1596_));
 sg13g2_xor2_1 _5513_ (.B(_1606_),
    .A(_1590_),
    .X(_1607_));
 sg13g2_and2_1 _5514_ (.A(_1604_),
    .B(_1607_),
    .X(_1608_));
 sg13g2_nand2_1 _5515_ (.Y(_1609_),
    .A(_1601_),
    .B(_1608_));
 sg13g2_o21ai_1 _5516_ (.B1(_1594_),
    .Y(_1610_),
    .A1(_1590_),
    .A2(_1606_));
 sg13g2_nand2_1 _5517_ (.Y(_1611_),
    .A(_2909_),
    .B(_1595_));
 sg13g2_mux2_1 _5518_ (.A0(_1610_),
    .A1(_2909_),
    .S(_1595_),
    .X(_1612_));
 sg13g2_nand2_1 _5519_ (.Y(_1613_),
    .A(_1609_),
    .B(_1611_));
 sg13g2_a21o_2 _5520_ (.A2(_1608_),
    .A1(_1601_),
    .B1(_1612_),
    .X(_1614_));
 sg13g2_inv_1 _5521_ (.Y(_1615_),
    .A(_1614_));
 sg13g2_and2_1 _5522_ (.A(_2898_),
    .B(_1614_),
    .X(_1616_));
 sg13g2_nand2_1 _5523_ (.Y(_1617_),
    .A(_1600_),
    .B(_1616_));
 sg13g2_a21oi_1 _5524_ (.A1(_0025_),
    .A2(_2914_),
    .Y(_1618_),
    .B1(\draw_score_inst.score[2] ));
 sg13g2_xor2_1 _5525_ (.B(_1614_),
    .A(_0018_),
    .X(_1619_));
 sg13g2_a22oi_1 _5526_ (.Y(_1620_),
    .B1(_1618_),
    .B2(_1619_),
    .A2(_1616_),
    .A1(_1600_));
 sg13g2_nor2_1 _5527_ (.A(_1600_),
    .B(_1616_),
    .Y(_1621_));
 sg13g2_nor3_1 _5528_ (.A(_1599_),
    .B(_1620_),
    .C(_1621_),
    .Y(_1622_));
 sg13g2_nand2_1 _5529_ (.Y(_1623_),
    .A(_1601_),
    .B(_1614_));
 sg13g2_a221oi_1 _5530_ (.B2(_1605_),
    .C1(_1622_),
    .B1(_1623_),
    .A1(_1599_),
    .Y(_1624_),
    .A2(_1617_));
 sg13g2_nor2_1 _5531_ (.A(_1605_),
    .B(_1623_),
    .Y(_1625_));
 sg13g2_or3_1 _5532_ (.A(_1607_),
    .B(_1624_),
    .C(_1625_),
    .X(_1626_));
 sg13g2_a22oi_1 _5533_ (.Y(_1627_),
    .B1(_1626_),
    .B2(_1609_),
    .A2(_1613_),
    .A1(_1612_));
 sg13g2_xor2_1 _5534_ (.B(_1614_),
    .A(_1585_),
    .X(_1628_));
 sg13g2_a21o_1 _5535_ (.A2(_1615_),
    .A1(_1585_),
    .B1(_1597_),
    .X(_1629_));
 sg13g2_inv_1 _5536_ (.Y(_1630_),
    .A(_1629_));
 sg13g2_or2_1 _5537_ (.X(_1631_),
    .B(_1628_),
    .A(_1597_));
 sg13g2_xnor2_1 _5538_ (.Y(_1632_),
    .A(net1202),
    .B(_1580_));
 sg13g2_nor4_1 _5539_ (.A(net1369),
    .B(_3219_),
    .C(_1497_),
    .D(_1632_),
    .Y(_1633_));
 sg13g2_inv_1 _5540_ (.Y(_1634_),
    .A(_1633_));
 sg13g2_nor2_2 _5541_ (.A(net1196),
    .B(_1634_),
    .Y(_1635_));
 sg13g2_inv_1 _5542_ (.Y(_1636_),
    .A(_1635_));
 sg13g2_nand4_1 _5543_ (.B(_1627_),
    .C(_1631_),
    .A(_1506_),
    .Y(_1637_),
    .D(_1635_));
 sg13g2_o21ai_1 _5544_ (.B1(_2909_),
    .Y(_1638_),
    .A1(_1585_),
    .A2(_1615_));
 sg13g2_nand2_1 _5545_ (.Y(_1639_),
    .A(_1628_),
    .B(_1638_));
 sg13g2_nand2_1 _5546_ (.Y(_1640_),
    .A(_1627_),
    .B(_1639_));
 sg13g2_nor2_1 _5547_ (.A(_1627_),
    .B(_1639_),
    .Y(_1641_));
 sg13g2_nand2b_1 _5548_ (.Y(_1642_),
    .B(_1641_),
    .A_N(_1401_));
 sg13g2_nor3_2 _5549_ (.A(net1380),
    .B(_3175_),
    .C(_1634_),
    .Y(_1643_));
 sg13g2_a22oi_1 _5550_ (.Y(_1644_),
    .B1(_1643_),
    .B2(_1492_),
    .A2(_1635_),
    .A1(_1504_));
 sg13g2_nor2_1 _5551_ (.A(_1629_),
    .B(_1641_),
    .Y(_1645_));
 sg13g2_nand2_1 _5552_ (.Y(_1646_),
    .A(_1635_),
    .B(_1638_));
 sg13g2_nand2_1 _5553_ (.Y(_1647_),
    .A(_1628_),
    .B(_1646_));
 sg13g2_o21ai_1 _5554_ (.B1(_1647_),
    .Y(_1648_),
    .A1(_1636_),
    .A2(_1640_));
 sg13g2_a21oi_1 _5555_ (.A1(_1629_),
    .A2(_1648_),
    .Y(_1649_),
    .B1(_1645_));
 sg13g2_or2_1 _5556_ (.X(_1650_),
    .B(_1649_),
    .A(_1644_));
 sg13g2_nand2_1 _5557_ (.Y(_1651_),
    .A(_1640_),
    .B(_1645_));
 sg13g2_nand4_1 _5558_ (.B(_1628_),
    .C(_1629_),
    .A(_1627_),
    .Y(_1652_),
    .D(_1638_));
 sg13g2_a22oi_1 _5559_ (.Y(_1653_),
    .B1(_1652_),
    .B2(_1506_),
    .A2(_1651_),
    .A1(_1504_));
 sg13g2_nand3_1 _5560_ (.B(_3068_),
    .C(_1633_),
    .A(_0033_),
    .Y(_1654_));
 sg13g2_or2_1 _5561_ (.X(_1655_),
    .B(_1654_),
    .A(_1653_));
 sg13g2_a21oi_1 _5562_ (.A1(\draw_score_inst.segment_rom_health.segments[2] ),
    .A2(_1506_),
    .Y(_1656_),
    .B1(_1504_));
 sg13g2_nand2b_1 _5563_ (.Y(_1657_),
    .B(_1562_),
    .A_N(_1656_));
 sg13g2_a22oi_1 _5564_ (.Y(_1658_),
    .B1(_1492_),
    .B2(\draw_score_inst.segment_rom_health.segments[6] ),
    .A2(_1403_),
    .A1(\draw_score_inst.segment_rom_health.segments[0] ));
 sg13g2_a22oi_1 _5565_ (.Y(_1659_),
    .B1(_1506_),
    .B2(\draw_score_inst.segment_rom_health.segments[4] ),
    .A2(_1504_),
    .A1(\draw_score_inst.segment_rom_health.segments[5] ));
 sg13g2_nand4_1 _5566_ (.B(_1630_),
    .C(_1640_),
    .A(_1403_),
    .Y(_1660_),
    .D(_1642_));
 sg13g2_o21ai_1 _5567_ (.B1(_1629_),
    .Y(_1661_),
    .A1(_1627_),
    .A2(_1628_));
 sg13g2_o21ai_1 _5568_ (.B1(_1660_),
    .Y(_1662_),
    .A1(_1404_),
    .A2(_1661_));
 sg13g2_nand2_1 _5569_ (.Y(_1663_),
    .A(_0371_),
    .B(_1568_));
 sg13g2_o21ai_1 _5570_ (.B1(_0347_),
    .Y(_1664_),
    .A1(net1369),
    .A2(_0345_));
 sg13g2_nor2_1 _5571_ (.A(net1360),
    .B(_0355_),
    .Y(_1665_));
 sg13g2_nand2_1 _5572_ (.Y(_1666_),
    .A(_0348_),
    .B(_1665_));
 sg13g2_nor2_1 _5573_ (.A(_1664_),
    .B(_1666_),
    .Y(_1667_));
 sg13g2_nand3_1 _5574_ (.B(net1194),
    .C(_0387_),
    .A(net1362),
    .Y(_1668_));
 sg13g2_nor3_1 _5575_ (.A(_3073_),
    .B(_3226_),
    .C(_1668_),
    .Y(_1669_));
 sg13g2_nand3_1 _5576_ (.B(_1570_),
    .C(_1577_),
    .A(_1564_),
    .Y(_1670_));
 sg13g2_nand2_1 _5577_ (.Y(_1671_),
    .A(_1643_),
    .B(_1662_));
 sg13g2_nand4_1 _5578_ (.B(_1650_),
    .C(_1655_),
    .A(_1637_),
    .Y(_1672_),
    .D(_1671_));
 sg13g2_nor4_1 _5579_ (.A(_1659_),
    .B(_1663_),
    .C(_1664_),
    .D(_1666_),
    .Y(_1673_));
 sg13g2_nand2_1 _5580_ (.Y(_1674_),
    .A(net1192),
    .B(_1663_));
 sg13g2_o21ai_1 _5581_ (.B1(_1657_),
    .Y(_1675_),
    .A1(_1658_),
    .A2(_1674_));
 sg13g2_nand4_1 _5582_ (.B(_0371_),
    .C(_1667_),
    .A(net1378),
    .Y(_1676_),
    .D(_1675_));
 sg13g2_nor2b_1 _5583_ (.A(_1673_),
    .B_N(_1676_),
    .Y(_1677_));
 sg13g2_nand3_1 _5584_ (.B(_0345_),
    .C(_1669_),
    .A(_3217_),
    .Y(_1678_));
 sg13g2_nor4_1 _5585_ (.A(_1388_),
    .B(_1389_),
    .C(_1677_),
    .D(_1678_),
    .Y(_1679_));
 sg13g2_a21o_1 _5586_ (.A2(_1672_),
    .A1(_1581_),
    .B1(_1679_),
    .X(_1680_));
 sg13g2_nor4_1 _5587_ (.A(_0347_),
    .B(_1500_),
    .C(_1511_),
    .D(_1512_),
    .Y(_1681_));
 sg13g2_or3_1 _5588_ (.A(_1502_),
    .B(_1509_),
    .C(_1681_),
    .X(_1682_));
 sg13g2_a221oi_1 _5589_ (.B2(_1395_),
    .C1(_1680_),
    .B1(_1682_),
    .A1(_1519_),
    .Y(_1683_),
    .A2(_1670_));
 sg13g2_a21oi_1 _5590_ (.A1(_1383_),
    .A2(_1683_),
    .Y(_0091_),
    .B1(_3103_));
 sg13g2_nor2_1 _5591_ (.A(_0477_),
    .B(_1363_),
    .Y(_1684_));
 sg13g2_nand2b_1 _5592_ (.Y(_1685_),
    .B(_1381_),
    .A_N(_3233_));
 sg13g2_inv_1 _5593_ (.Y(_1686_),
    .A(_1685_));
 sg13g2_o21ai_1 _5594_ (.B1(_1686_),
    .Y(_1687_),
    .A1(_0291_),
    .A2(_1684_));
 sg13g2_a21oi_1 _5595_ (.A1(_1683_),
    .A2(_1687_),
    .Y(_0092_),
    .B1(_3103_));
 sg13g2_and2_1 _5596_ (.A(_0478_),
    .B(_1362_),
    .X(_1688_));
 sg13g2_a21oi_2 _5597_ (.B1(_3188_),
    .Y(_1689_),
    .A2(net1284),
    .A1(net1297));
 sg13g2_nand2_1 _5598_ (.Y(_1690_),
    .A(net1112),
    .B(_1689_));
 sg13g2_o21ai_1 _5599_ (.B1(_1690_),
    .Y(_1691_),
    .A1(_3212_),
    .A2(net1111));
 sg13g2_nand2_2 _5600_ (.Y(_1692_),
    .A(_3189_),
    .B(_0534_));
 sg13g2_nor2_1 _5601_ (.A(net1290),
    .B(_0048_),
    .Y(_1693_));
 sg13g2_a21oi_2 _5602_ (.B1(_1693_),
    .Y(_1694_),
    .A2(_2905_),
    .A1(net1290));
 sg13g2_nand2_1 _5603_ (.Y(_1695_),
    .A(net1111),
    .B(_1692_));
 sg13g2_o21ai_1 _5604_ (.B1(_1695_),
    .Y(_1696_),
    .A1(net1112),
    .A2(_1694_));
 sg13g2_nor2_1 _5605_ (.A(net1112),
    .B(_1689_),
    .Y(_1697_));
 sg13g2_a21oi_2 _5606_ (.B1(_1697_),
    .Y(_1698_),
    .A2(net1111),
    .A1(net1189));
 sg13g2_nor2_1 _5607_ (.A(net1111),
    .B(_1692_),
    .Y(_1699_));
 sg13g2_a21oi_2 _5608_ (.B1(_1699_),
    .Y(_1700_),
    .A2(_1694_),
    .A1(net1112));
 sg13g2_mux4_1 _5609_ (.S0(net1086),
    .A0(_1691_),
    .A1(_1696_),
    .A2(_1700_),
    .A3(_1698_),
    .S1(_0706_),
    .X(_1701_));
 sg13g2_nand3_1 _5610_ (.B(_0705_),
    .C(_1701_),
    .A(\aliens_alive[3] ),
    .Y(_1702_));
 sg13g2_mux4_1 _5611_ (.S0(net1087),
    .A0(_1691_),
    .A1(_1696_),
    .A2(_1700_),
    .A3(_1698_),
    .S1(_0650_),
    .X(_1703_));
 sg13g2_nand3_1 _5612_ (.B(_0640_),
    .C(_1703_),
    .A(\aliens_alive[7] ),
    .Y(_1704_));
 sg13g2_nand2_1 _5613_ (.Y(_1705_),
    .A(net1133),
    .B(_1689_));
 sg13g2_o21ai_1 _5614_ (.B1(_1705_),
    .Y(_1706_),
    .A1(net1189),
    .A2(net1133));
 sg13g2_nor2_1 _5615_ (.A(net1132),
    .B(_1692_),
    .Y(_1707_));
 sg13g2_a21oi_2 _5616_ (.B1(_1707_),
    .Y(_1708_),
    .A2(_1694_),
    .A1(net1133));
 sg13g2_nor2_1 _5617_ (.A(net1133),
    .B(_1689_),
    .Y(_1709_));
 sg13g2_a21oi_2 _5618_ (.B1(_1709_),
    .Y(_1710_),
    .A2(net1133),
    .A1(net1189));
 sg13g2_nand2_1 _5619_ (.Y(_1711_),
    .A(net1132),
    .B(_1692_));
 sg13g2_o21ai_1 _5620_ (.B1(_1711_),
    .Y(_1712_),
    .A1(net1133),
    .A2(_1694_));
 sg13g2_mux4_1 _5621_ (.S0(_0528_),
    .A0(_1708_),
    .A1(_1710_),
    .A2(_1706_),
    .A3(_1712_),
    .S1(_0558_),
    .X(_1713_));
 sg13g2_nand3_1 _5622_ (.B(_0527_),
    .C(_1713_),
    .A(\aliens_alive[4] ),
    .Y(_1714_));
 sg13g2_mux4_1 _5623_ (.S0(_0743_),
    .A0(_1706_),
    .A1(_1708_),
    .A2(_1712_),
    .A3(_1710_),
    .S1(_0529_),
    .X(_1715_));
 sg13g2_nand3_1 _5624_ (.B(_0742_),
    .C(_1715_),
    .A(\aliens_alive[0] ),
    .Y(_1716_));
 sg13g2_mux4_1 _5625_ (.S0(net1122),
    .A0(_1700_),
    .A1(_1698_),
    .A2(_1691_),
    .A3(_1696_),
    .S1(_0804_),
    .X(_1717_));
 sg13g2_nand3_1 _5626_ (.B(_0798_),
    .C(_1717_),
    .A(\aliens_alive[1] ),
    .Y(_1718_));
 sg13g2_mux4_1 _5627_ (.S0(net1122),
    .A0(_1698_),
    .A1(_1700_),
    .A2(_1696_),
    .A3(_1691_),
    .S1(_0864_),
    .X(_1719_));
 sg13g2_nand3_1 _5628_ (.B(_0863_),
    .C(_1719_),
    .A(\aliens_alive[5] ),
    .Y(_1720_));
 sg13g2_mux4_1 _5629_ (.S0(_0908_),
    .A0(_1706_),
    .A1(_1708_),
    .A2(_1712_),
    .A3(_1710_),
    .S1(net1118),
    .X(_1721_));
 sg13g2_nand3_1 _5630_ (.B(_0901_),
    .C(_1721_),
    .A(\aliens_alive[6] ),
    .Y(_1722_));
 sg13g2_mux4_1 _5631_ (.S0(net1116),
    .A0(_1708_),
    .A1(_1710_),
    .A2(_1706_),
    .A3(_1712_),
    .S1(_0958_),
    .X(_1723_));
 sg13g2_nand3_1 _5632_ (.B(_0956_),
    .C(_1723_),
    .A(\aliens_alive[2] ),
    .Y(_1724_));
 sg13g2_nand4_1 _5633_ (.B(_1704_),
    .C(_1714_),
    .A(_1702_),
    .Y(_1725_),
    .D(_1720_));
 sg13g2_nor2b_1 _5634_ (.A(_1725_),
    .B_N(_1722_),
    .Y(_1726_));
 sg13g2_nand4_1 _5635_ (.B(_1718_),
    .C(_1724_),
    .A(_1716_),
    .Y(_1727_),
    .D(_1726_));
 sg13g2_nor3_1 _5636_ (.A(net1273),
    .B(_0015_),
    .C(_0979_),
    .Y(_1728_));
 sg13g2_nand4_1 _5637_ (.B(_0974_),
    .C(_1727_),
    .A(_3215_),
    .Y(_1729_),
    .D(_1728_));
 sg13g2_o21ai_1 _5638_ (.B1(_1688_),
    .Y(_1730_),
    .A1(_1114_),
    .A2(_1729_));
 sg13g2_nor2b_1 _5639_ (.A(_3233_),
    .B_N(_1730_),
    .Y(_1731_));
 sg13g2_nand2_1 _5640_ (.Y(_1732_),
    .A(_1381_),
    .B(_1731_));
 sg13g2_a21oi_1 _5641_ (.A1(_1683_),
    .A2(_1732_),
    .Y(_0093_),
    .B1(_3103_));
 sg13g2_nor2_1 _5642_ (.A(_1382_),
    .B(_1731_),
    .Y(_1733_));
 sg13g2_a21oi_1 _5643_ (.A1(_1683_),
    .A2(_1733_),
    .Y(_0094_),
    .B1(_3103_));
 sg13g2_a21o_1 _5644_ (.A2(_3061_),
    .A1(net218),
    .B1(_3062_),
    .X(_0095_));
 sg13g2_nor2b_1 _5645_ (.A(_3233_),
    .B_N(_0478_),
    .Y(_1734_));
 sg13g2_nor2b_1 _5646_ (.A(_1114_),
    .B_N(_1362_),
    .Y(_1735_));
 sg13g2_a21o_1 _5647_ (.A2(_1735_),
    .A1(_1734_),
    .B1(_1382_),
    .X(_1736_));
 sg13g2_a21oi_1 _5648_ (.A1(_1683_),
    .A2(_1736_),
    .Y(_0097_),
    .B1(_3103_));
 sg13g2_nor2_1 _5649_ (.A(_0477_),
    .B(_1735_),
    .Y(_1737_));
 sg13g2_nor3_1 _5650_ (.A(_0291_),
    .B(_1685_),
    .C(_1737_),
    .Y(_1738_));
 sg13g2_a21oi_1 _5651_ (.A1(_1683_),
    .A2(_1738_),
    .Y(_0098_),
    .B1(_3103_));
 sg13g2_nand2b_2 _5652_ (.Y(_1739_),
    .B(net4),
    .A_N(prev_button2));
 sg13g2_nor2_1 _5653_ (.A(net1327),
    .B(_1739_),
    .Y(_1740_));
 sg13g2_o21ai_1 _5654_ (.B1(net1178),
    .Y(_1741_),
    .A1(net297),
    .A2(net1155));
 sg13g2_inv_1 _5655_ (.Y(_0099_),
    .A(_1741_));
 sg13g2_o21ai_1 _5656_ (.B1(net1179),
    .Y(_1742_),
    .A1(net1350),
    .A2(net1155));
 sg13g2_a21oi_1 _5657_ (.A1(_2840_),
    .A2(net1155),
    .Y(_0100_),
    .B1(_1742_));
 sg13g2_nor2_2 _5658_ (.A(net379),
    .B(\myShooter.shooter_left_x[1] ),
    .Y(_1743_));
 sg13g2_nand2_1 _5659_ (.Y(_1744_),
    .A(net1263),
    .B(\myShooter.shooter_left_x[1] ));
 sg13g2_nor2b_1 _5660_ (.A(_1743_),
    .B_N(_1744_),
    .Y(_1745_));
 sg13g2_o21ai_1 _5661_ (.B1(net1179),
    .Y(_1746_),
    .A1(net1348),
    .A2(net1155));
 sg13g2_a21oi_1 _5662_ (.A1(net1155),
    .A2(_1745_),
    .Y(_0101_),
    .B1(_1746_));
 sg13g2_xnor2_1 _5663_ (.Y(_1747_),
    .A(net293),
    .B(_1743_));
 sg13g2_o21ai_1 _5664_ (.B1(net1178),
    .Y(_1748_),
    .A1(net1346),
    .A2(net1155));
 sg13g2_a21oi_1 _5665_ (.A1(net1155),
    .A2(net294),
    .Y(_0102_),
    .B1(_1748_));
 sg13g2_o21ai_1 _5666_ (.B1(net1261),
    .Y(_1749_),
    .A1(net1263),
    .A2(\myShooter.shooter_left_x[1] ));
 sg13g2_nand3b_1 _5667_ (.B(net1261),
    .C(net1260),
    .Y(_1750_),
    .A_N(_1743_));
 sg13g2_xor2_1 _5668_ (.B(_1749_),
    .A(net1260),
    .X(_1751_));
 sg13g2_o21ai_1 _5669_ (.B1(net1178),
    .Y(_1752_),
    .A1(net1344),
    .A2(net1155));
 sg13g2_a21oi_1 _5670_ (.A1(net1157),
    .A2(_1751_),
    .Y(_0103_),
    .B1(_1752_));
 sg13g2_xnor2_1 _5671_ (.Y(_1753_),
    .A(_2838_),
    .B(_1750_));
 sg13g2_o21ai_1 _5672_ (.B1(net1178),
    .Y(_1754_),
    .A1(net1343),
    .A2(net1156));
 sg13g2_a21oi_1 _5673_ (.A1(net1156),
    .A2(_1753_),
    .Y(_0104_),
    .B1(_1754_));
 sg13g2_nor2_1 _5674_ (.A(net377),
    .B(_1750_),
    .Y(_1755_));
 sg13g2_xnor2_1 _5675_ (.Y(_1756_),
    .A(net1258),
    .B(_1755_));
 sg13g2_o21ai_1 _5676_ (.B1(net1178),
    .Y(_1757_),
    .A1(net1338),
    .A2(net1156));
 sg13g2_a21oi_1 _5677_ (.A1(net1156),
    .A2(_1756_),
    .Y(_0105_),
    .B1(_1757_));
 sg13g2_nor3_1 _5678_ (.A(_2837_),
    .B(_2976_),
    .C(_1749_),
    .Y(_1758_));
 sg13g2_xnor2_1 _5679_ (.Y(_1759_),
    .A(net1257),
    .B(_1758_));
 sg13g2_o21ai_1 _5680_ (.B1(net1178),
    .Y(_1760_),
    .A1(net1334),
    .A2(net1156));
 sg13g2_a21oi_1 _5681_ (.A1(net1156),
    .A2(_1759_),
    .Y(_0106_),
    .B1(_1760_));
 sg13g2_nor2b_1 _5682_ (.A(net406),
    .B_N(_1758_),
    .Y(_1761_));
 sg13g2_xnor2_1 _5683_ (.Y(_1762_),
    .A(net1256),
    .B(_1761_));
 sg13g2_o21ai_1 _5684_ (.B1(net1178),
    .Y(_1763_),
    .A1(net1333),
    .A2(net1156));
 sg13g2_a21oi_1 _5685_ (.A1(net1157),
    .A2(_1762_),
    .Y(_0107_),
    .B1(_1763_));
 sg13g2_nor2_1 _5686_ (.A(_3004_),
    .B(_1749_),
    .Y(_1764_));
 sg13g2_xnor2_1 _5687_ (.Y(_1765_),
    .A(net355),
    .B(_1764_));
 sg13g2_o21ai_1 _5688_ (.B1(net1175),
    .Y(_1766_),
    .A1(net1330),
    .A2(net1157));
 sg13g2_a21oi_2 _5689_ (.B1(_1766_),
    .Y(_0108_),
    .A2(_1765_),
    .A1(net1157));
 sg13g2_nand2_2 _5690_ (.Y(_1767_),
    .A(net1327),
    .B(net1151));
 sg13g2_nand2_1 _5691_ (.Y(_1768_),
    .A(_0827_),
    .B(net1119));
 sg13g2_nor2_2 _5692_ (.A(net1236),
    .B(_1768_),
    .Y(_1769_));
 sg13g2_nand3_1 _5693_ (.B(_0823_),
    .C(_1769_),
    .A(_0821_),
    .Y(_1770_));
 sg13g2_nor2_1 _5694_ (.A(_0851_),
    .B(_1770_),
    .Y(_1771_));
 sg13g2_nand2_1 _5695_ (.Y(_1772_),
    .A(_0851_),
    .B(_1770_));
 sg13g2_nand3_1 _5696_ (.B(_0851_),
    .C(_1770_),
    .A(net1330),
    .Y(_1773_));
 sg13g2_xnor2_1 _5697_ (.Y(_1774_),
    .A(_0823_),
    .B(_1769_));
 sg13g2_nor2_1 _5698_ (.A(net1334),
    .B(_1774_),
    .Y(_1775_));
 sg13g2_xnor2_1 _5699_ (.Y(_1776_),
    .A(_0827_),
    .B(net1119));
 sg13g2_nand2_1 _5700_ (.Y(_1777_),
    .A(net1343),
    .B(_1776_));
 sg13g2_nand2_1 _5701_ (.Y(_1778_),
    .A(_2886_),
    .B(_0831_));
 sg13g2_nand2_1 _5702_ (.Y(_1779_),
    .A(net1347),
    .B(_0835_));
 sg13g2_nor2_2 _5703_ (.A(net1253),
    .B(\pb_x[1] ),
    .Y(_1780_));
 sg13g2_inv_1 _5704_ (.Y(_1781_),
    .A(_1780_));
 sg13g2_xnor2_1 _5705_ (.Y(_1782_),
    .A(_0005_),
    .B(_0766_));
 sg13g2_nand2_1 _5706_ (.Y(_1783_),
    .A(net1349),
    .B(_0767_));
 sg13g2_o21ai_1 _5707_ (.B1(_1783_),
    .Y(_1784_),
    .A1(_1780_),
    .A2(_1782_));
 sg13g2_xnor2_1 _5708_ (.Y(_1785_),
    .A(_0069_),
    .B(_0835_));
 sg13g2_nand2_1 _5709_ (.Y(_1786_),
    .A(_1784_),
    .B(_1785_));
 sg13g2_xnor2_1 _5710_ (.Y(_1787_),
    .A(net1344),
    .B(net1119));
 sg13g2_a21oi_2 _5711_ (.B1(_1787_),
    .Y(_1788_),
    .A2(_1786_),
    .A1(_1779_));
 sg13g2_a21oi_1 _5712_ (.A1(net1253),
    .A2(net1350),
    .Y(_1789_),
    .B1(net1351));
 sg13g2_nand3_1 _5713_ (.B(_1783_),
    .C(_1789_),
    .A(_1779_),
    .Y(_1790_));
 sg13g2_a22oi_1 _5714_ (.Y(_1791_),
    .B1(_1788_),
    .B2(_1790_),
    .A2(net1119),
    .A1(_2886_));
 sg13g2_xor2_1 _5715_ (.B(_1776_),
    .A(net1342),
    .X(_1792_));
 sg13g2_o21ai_1 _5716_ (.B1(_1777_),
    .Y(_1793_),
    .A1(_1791_),
    .A2(_1792_));
 sg13g2_a21oi_1 _5717_ (.A1(_0827_),
    .A2(net1119),
    .Y(_1794_),
    .B1(_0843_));
 sg13g2_nor2_1 _5718_ (.A(_1769_),
    .B(_1794_),
    .Y(_1795_));
 sg13g2_inv_1 _5719_ (.Y(_1796_),
    .A(_1795_));
 sg13g2_xor2_1 _5720_ (.B(_1795_),
    .A(net1337),
    .X(_1797_));
 sg13g2_nand2_1 _5721_ (.Y(_1798_),
    .A(_1793_),
    .B(_1797_));
 sg13g2_a21o_1 _5722_ (.A2(_1769_),
    .A1(_0823_),
    .B1(_0821_),
    .X(_1799_));
 sg13g2_and2_1 _5723_ (.A(_1770_),
    .B(_1799_),
    .X(_1800_));
 sg13g2_nor2_1 _5724_ (.A(net1331),
    .B(_1800_),
    .Y(_1801_));
 sg13g2_a22oi_1 _5725_ (.Y(_1802_),
    .B1(_1796_),
    .B2(net1338),
    .A2(_1774_),
    .A1(net1336));
 sg13g2_a221oi_1 _5726_ (.B2(_1798_),
    .C1(_1775_),
    .B1(_1802_),
    .A1(net1331),
    .Y(_1803_),
    .A2(_1800_));
 sg13g2_xor2_1 _5727_ (.B(_1772_),
    .A(_0058_),
    .X(_1804_));
 sg13g2_o21ai_1 _5728_ (.B1(_1804_),
    .Y(_1805_),
    .A1(_1801_),
    .A2(_1803_));
 sg13g2_a21oi_2 _5729_ (.B1(_1771_),
    .Y(_1806_),
    .A2(_1805_),
    .A1(_1773_));
 sg13g2_nor2_1 _5730_ (.A(net1162),
    .B(_0827_),
    .Y(_1807_));
 sg13g2_a22oi_1 _5731_ (.Y(_1808_),
    .B1(_0835_),
    .B2(_3242_),
    .A2(_0832_),
    .A1(net1143));
 sg13g2_a22oi_1 _5732_ (.Y(_1809_),
    .B1(_0836_),
    .B2(_3243_),
    .A2(net1186),
    .A1(_3245_));
 sg13g2_nor2_2 _5733_ (.A(_2827_),
    .B(net1350),
    .Y(_1810_));
 sg13g2_inv_1 _5734_ (.Y(_1811_),
    .A(_1810_));
 sg13g2_xor2_1 _5735_ (.B(net1186),
    .A(_3245_),
    .X(_1812_));
 sg13g2_inv_1 _5736_ (.Y(_1813_),
    .A(_1812_));
 sg13g2_o21ai_1 _5737_ (.B1(_1809_),
    .Y(_1814_),
    .A1(_1810_),
    .A2(_1813_));
 sg13g2_a22oi_1 _5738_ (.Y(_1815_),
    .B1(_1808_),
    .B2(_1814_),
    .A2(net1119),
    .A1(net1142));
 sg13g2_nand2_1 _5739_ (.Y(_1816_),
    .A(net1162),
    .B(_0827_));
 sg13g2_o21ai_1 _5740_ (.B1(_1816_),
    .Y(_1817_),
    .A1(_1807_),
    .A2(_1815_));
 sg13g2_o21ai_1 _5741_ (.B1(_1817_),
    .Y(_1818_),
    .A1(net1140),
    .A2(_0843_));
 sg13g2_a22oi_1 _5742_ (.Y(_1819_),
    .B1(_0843_),
    .B2(net1141),
    .A2(_0823_),
    .A1(_3262_));
 sg13g2_a22oi_1 _5743_ (.Y(_1820_),
    .B1(_1818_),
    .B2(_1819_),
    .A2(_0824_),
    .A1(net1139));
 sg13g2_o21ai_1 _5744_ (.B1(_1820_),
    .Y(_1821_),
    .A1(net1136),
    .A2(_0821_));
 sg13g2_a22oi_1 _5745_ (.Y(_1822_),
    .B1(_0852_),
    .B2(net1135),
    .A2(_0821_),
    .A1(net1137));
 sg13g2_a221oi_1 _5746_ (.B2(_1822_),
    .C1(_3273_),
    .B1(_1821_),
    .A1(_3270_),
    .Y(_1823_),
    .A2(_0851_));
 sg13g2_nor2_2 _5747_ (.A(net1321),
    .B(\pb_y[9] ),
    .Y(_1824_));
 sg13g2_or2_1 _5748_ (.X(_1825_),
    .B(\pb_y[9] ),
    .A(net1321));
 sg13g2_nor2_1 _5749_ (.A(_3279_),
    .B(_1825_),
    .Y(_1826_));
 sg13g2_o21ai_1 _5750_ (.B1(_1826_),
    .Y(_1827_),
    .A1(_3305_),
    .A2(_3308_));
 sg13g2_nor3_1 _5751_ (.A(_0071_),
    .B(_3284_),
    .C(_3286_),
    .Y(_1828_));
 sg13g2_nor2_1 _5752_ (.A(_2893_),
    .B(_2894_),
    .Y(_1829_));
 sg13g2_a21oi_1 _5753_ (.A1(net1325),
    .A2(_1829_),
    .Y(_1830_),
    .B1(_3277_));
 sg13g2_nor2b_1 _5754_ (.A(_1830_),
    .B_N(_1828_),
    .Y(_1831_));
 sg13g2_or2_1 _5755_ (.X(_1832_),
    .B(_1831_),
    .A(_1827_));
 sg13g2_inv_1 _5756_ (.Y(_1833_),
    .A(_1832_));
 sg13g2_nand2_1 _5757_ (.Y(_1834_),
    .A(_3284_),
    .B(_3286_));
 sg13g2_nor2_1 _5758_ (.A(net1326),
    .B(_2894_),
    .Y(_1835_));
 sg13g2_a21oi_1 _5759_ (.A1(_2892_),
    .A2(_1835_),
    .Y(_1836_),
    .B1(_3295_));
 sg13g2_o21ai_1 _5760_ (.B1(_3284_),
    .Y(_1837_),
    .A1(_3286_),
    .A2(_1836_));
 sg13g2_a21oi_1 _5761_ (.A1(_3309_),
    .A2(_1837_),
    .Y(_1838_),
    .B1(_1832_));
 sg13g2_o21ai_1 _5762_ (.B1(_1824_),
    .Y(_1839_),
    .A1(_2887_),
    .A2(_2888_));
 sg13g2_nor3_1 _5763_ (.A(_2889_),
    .B(\pb_y[4] ),
    .C(net1324),
    .Y(_1840_));
 sg13g2_nand2_1 _5764_ (.Y(_1841_),
    .A(_2894_),
    .B(_1840_));
 sg13g2_a221oi_1 _5765_ (.B2(_0072_),
    .C1(_2887_),
    .B1(_1841_),
    .A1(_3291_),
    .Y(_1842_),
    .A2(_1840_));
 sg13g2_nor3_2 _5766_ (.A(_1838_),
    .B(_1839_),
    .C(_1842_),
    .Y(_1843_));
 sg13g2_nand2_1 _5767_ (.Y(_1844_),
    .A(\aliens_alive[5] ),
    .B(_1843_));
 sg13g2_or3_2 _5768_ (.A(_1806_),
    .B(_1823_),
    .C(_1844_),
    .X(_1845_));
 sg13g2_and3_1 _5769_ (.X(_1846_),
    .A(_0760_),
    .B(_0923_),
    .C(_0926_));
 sg13g2_nand2b_1 _5770_ (.Y(_1847_),
    .B(_1846_),
    .A_N(_0935_));
 sg13g2_inv_1 _5771_ (.Y(_1848_),
    .A(_1847_));
 sg13g2_nand2_1 _5772_ (.Y(_1849_),
    .A(_2895_),
    .B(_1848_));
 sg13g2_and2_1 _5773_ (.A(_0951_),
    .B(_1849_),
    .X(_1850_));
 sg13g2_nand2_1 _5774_ (.Y(_1851_),
    .A(net1329),
    .B(_1850_));
 sg13g2_a21oi_1 _5775_ (.A1(_0760_),
    .A2(_0926_),
    .Y(_1852_),
    .B1(_0923_));
 sg13g2_or2_1 _5776_ (.X(_1853_),
    .B(_1852_),
    .A(_1846_));
 sg13g2_nand2_1 _5777_ (.Y(_1854_),
    .A(net1339),
    .B(_1853_));
 sg13g2_xnor2_1 _5778_ (.Y(_1855_),
    .A(_0759_),
    .B(_0926_));
 sg13g2_nand2_1 _5779_ (.Y(_1856_),
    .A(_2886_),
    .B(_0760_));
 sg13g2_nand2_1 _5780_ (.Y(_1857_),
    .A(net1347),
    .B(_0762_));
 sg13g2_nand2_1 _5781_ (.Y(_1858_),
    .A(net1349),
    .B(net1186));
 sg13g2_a22oi_1 _5782_ (.Y(_1859_),
    .B1(_1781_),
    .B2(_1782_),
    .A2(net1186),
    .A1(net1349));
 sg13g2_xor2_1 _5783_ (.B(_0762_),
    .A(_0069_),
    .X(_1860_));
 sg13g2_o21ai_1 _5784_ (.B1(_1857_),
    .Y(_1861_),
    .A1(_1859_),
    .A2(_1860_));
 sg13g2_xnor2_1 _5785_ (.Y(_1862_),
    .A(net1345),
    .B(_0759_));
 sg13g2_a22oi_1 _5786_ (.Y(_1863_),
    .B1(_1861_),
    .B2(_1862_),
    .A2(_0760_),
    .A1(_2886_));
 sg13g2_xnor2_1 _5787_ (.Y(_1864_),
    .A(_0065_),
    .B(_1853_));
 sg13g2_nand2_1 _5788_ (.Y(_1865_),
    .A(net1340),
    .B(_1855_));
 sg13g2_o21ai_1 _5789_ (.B1(_1863_),
    .Y(_1866_),
    .A1(net1341),
    .A2(_1855_));
 sg13g2_nand3_1 _5790_ (.B(_1865_),
    .C(_1866_),
    .A(_1864_),
    .Y(_1867_));
 sg13g2_xor2_1 _5791_ (.B(_1846_),
    .A(_0935_),
    .X(_1868_));
 sg13g2_xor2_1 _5792_ (.B(_1868_),
    .A(_0060_),
    .X(_1869_));
 sg13g2_a21oi_1 _5793_ (.A1(_1854_),
    .A2(_1867_),
    .Y(_1870_),
    .B1(_1869_));
 sg13g2_o21ai_1 _5794_ (.B1(_1849_),
    .Y(_1871_),
    .A1(_0939_),
    .A2(_1848_));
 sg13g2_a221oi_1 _5795_ (.B2(\pb_x[8] ),
    .C1(_1870_),
    .B1(_1871_),
    .A1(net1336),
    .Y(_1872_),
    .A2(_1868_));
 sg13g2_xnor2_1 _5796_ (.Y(_1873_),
    .A(_0058_),
    .B(_1850_));
 sg13g2_o21ai_1 _5797_ (.B1(_1873_),
    .Y(_1874_),
    .A1(net1333),
    .A2(_1871_));
 sg13g2_o21ai_1 _5798_ (.B1(_1851_),
    .Y(_1875_),
    .A1(_1872_),
    .A2(_1874_));
 sg13g2_o21ai_1 _5799_ (.B1(_1875_),
    .Y(_1876_),
    .A1(_0951_),
    .A2(_1849_));
 sg13g2_nor2_1 _5800_ (.A(net1139),
    .B(_0935_),
    .Y(_1877_));
 sg13g2_nor2_1 _5801_ (.A(net1141),
    .B(_0923_),
    .Y(_1878_));
 sg13g2_a22oi_1 _5802_ (.Y(_1879_),
    .B1(_0762_),
    .B2(_3242_),
    .A2(_0759_),
    .A1(net1143));
 sg13g2_nor2_1 _5803_ (.A(_3242_),
    .B(_0762_),
    .Y(_1880_));
 sg13g2_a21oi_1 _5804_ (.A1(net1188),
    .A2(_0767_),
    .Y(_1881_),
    .B1(_1880_));
 sg13g2_nor2_1 _5805_ (.A(net1252),
    .B(_2873_),
    .Y(_1882_));
 sg13g2_o21ai_1 _5806_ (.B1(_1811_),
    .Y(_1883_),
    .A1(_0077_),
    .A2(_1882_));
 sg13g2_o21ai_1 _5807_ (.B1(_1881_),
    .Y(_1884_),
    .A1(_1812_),
    .A2(_1883_));
 sg13g2_nand2_1 _5808_ (.Y(_1885_),
    .A(net1161),
    .B(_0926_));
 sg13g2_a22oi_1 _5809_ (.Y(_1886_),
    .B1(_1879_),
    .B2(_1884_),
    .A2(_0760_),
    .A1(_3241_));
 sg13g2_a21oi_1 _5810_ (.A1(_1885_),
    .A2(_1886_),
    .Y(_1887_),
    .B1(_1878_));
 sg13g2_o21ai_1 _5811_ (.B1(_1887_),
    .Y(_1888_),
    .A1(_3237_),
    .A2(_0926_));
 sg13g2_a21oi_1 _5812_ (.A1(net1141),
    .A2(_0923_),
    .Y(_1889_),
    .B1(_1877_));
 sg13g2_nor2_1 _5813_ (.A(net1137),
    .B(_0939_),
    .Y(_1890_));
 sg13g2_a221oi_1 _5814_ (.B2(_1889_),
    .C1(_1890_),
    .B1(_1888_),
    .A1(net1139),
    .Y(_1891_),
    .A2(_0935_));
 sg13g2_nand2_1 _5815_ (.Y(_1892_),
    .A(net1136),
    .B(_0939_));
 sg13g2_o21ai_1 _5816_ (.B1(_1892_),
    .Y(_1893_),
    .A1(_3270_),
    .A2(_0951_));
 sg13g2_a21oi_1 _5817_ (.A1(_3270_),
    .A2(_0951_),
    .Y(_1894_),
    .B1(_3273_));
 sg13g2_o21ai_1 _5818_ (.B1(_1894_),
    .Y(_1895_),
    .A1(_1891_),
    .A2(_1893_));
 sg13g2_nand4_1 _5819_ (.B(_1843_),
    .C(_1876_),
    .A(net239),
    .Y(_1896_),
    .D(_1895_));
 sg13g2_nand2_1 _5820_ (.Y(_1897_),
    .A(_0757_),
    .B(_0760_));
 sg13g2_xnor2_1 _5821_ (.Y(_1898_),
    .A(_0757_),
    .B(_0759_));
 sg13g2_nor2b_1 _5822_ (.A(_1898_),
    .B_N(\pb_x[5] ),
    .Y(_1899_));
 sg13g2_and4_1 _5823_ (.A(_1789_),
    .B(_1856_),
    .C(_1857_),
    .D(_1858_),
    .X(_1900_));
 sg13g2_xnor2_1 _5824_ (.Y(_1901_),
    .A(net1340),
    .B(_1898_));
 sg13g2_nor3_1 _5825_ (.A(_1863_),
    .B(_1900_),
    .C(_1901_),
    .Y(_1902_));
 sg13g2_nor2_1 _5826_ (.A(_1899_),
    .B(_1902_),
    .Y(_1903_));
 sg13g2_nor2_1 _5827_ (.A(net1235),
    .B(_1897_),
    .Y(_1904_));
 sg13g2_a21o_1 _5828_ (.A2(_1897_),
    .A1(_0777_),
    .B1(_1904_),
    .X(_1905_));
 sg13g2_xor2_1 _5829_ (.B(_1905_),
    .A(_0065_),
    .X(_1906_));
 sg13g2_nor3_1 _5830_ (.A(net1235),
    .B(_0754_),
    .C(_1897_),
    .Y(_1907_));
 sg13g2_xor2_1 _5831_ (.B(_1904_),
    .A(_0754_),
    .X(_1908_));
 sg13g2_a22oi_1 _5832_ (.Y(_1909_),
    .B1(_1908_),
    .B2(net1336),
    .A2(_1905_),
    .A1(net1339));
 sg13g2_o21ai_1 _5833_ (.B1(_1909_),
    .Y(_1910_),
    .A1(_1903_),
    .A2(_1906_));
 sg13g2_and2_1 _5834_ (.A(_2895_),
    .B(_1907_),
    .X(_1911_));
 sg13g2_inv_1 _5835_ (.Y(_1912_),
    .A(_1911_));
 sg13g2_o21ai_1 _5836_ (.B1(_1912_),
    .Y(_1913_),
    .A1(_0752_),
    .A2(_1907_));
 sg13g2_xor2_1 _5837_ (.B(_1913_),
    .A(net1331),
    .X(_1914_));
 sg13g2_o21ai_1 _5838_ (.B1(_1910_),
    .Y(_1915_),
    .A1(net1335),
    .A2(_1908_));
 sg13g2_nor2_1 _5839_ (.A(_0786_),
    .B(_1911_),
    .Y(_1916_));
 sg13g2_a22oi_1 _5840_ (.Y(_1917_),
    .B1(_1916_),
    .B2(net1328),
    .A2(_1913_),
    .A1(net1332));
 sg13g2_o21ai_1 _5841_ (.B1(_1917_),
    .Y(_1918_),
    .A1(_1914_),
    .A2(_1915_));
 sg13g2_nor2_1 _5842_ (.A(net1328),
    .B(_1916_),
    .Y(_1919_));
 sg13g2_a21oi_1 _5843_ (.A1(_0786_),
    .A2(_1911_),
    .Y(_1920_),
    .B1(_1919_));
 sg13g2_nand2_2 _5844_ (.Y(_1921_),
    .A(_1918_),
    .B(_1920_));
 sg13g2_nor2_1 _5845_ (.A(net1161),
    .B(_0757_),
    .Y(_1922_));
 sg13g2_o21ai_1 _5846_ (.B1(_1881_),
    .Y(_1923_),
    .A1(_1810_),
    .A2(_1812_));
 sg13g2_a22oi_1 _5847_ (.Y(_1924_),
    .B1(_1879_),
    .B2(_1923_),
    .A2(_0760_),
    .A1(_3241_));
 sg13g2_nor2_1 _5848_ (.A(_3255_),
    .B(_0777_),
    .Y(_1925_));
 sg13g2_a21oi_1 _5849_ (.A1(net1161),
    .A2(_0757_),
    .Y(_1926_),
    .B1(_1925_));
 sg13g2_o21ai_1 _5850_ (.B1(_1926_),
    .Y(_1927_),
    .A1(_1922_),
    .A2(_1924_));
 sg13g2_a22oi_1 _5851_ (.Y(_1928_),
    .B1(_0777_),
    .B2(_3255_),
    .A2(_0754_),
    .A1(net1138));
 sg13g2_nand2_1 _5852_ (.Y(_1929_),
    .A(_1927_),
    .B(_1928_));
 sg13g2_o21ai_1 _5853_ (.B1(_1929_),
    .Y(_1930_),
    .A1(net1138),
    .A2(_0754_));
 sg13g2_o21ai_1 _5854_ (.B1(_1930_),
    .Y(_1931_),
    .A1(net1136),
    .A2(_0752_));
 sg13g2_a22oi_1 _5855_ (.Y(_1932_),
    .B1(_0786_),
    .B2(net1135),
    .A2(_0752_),
    .A1(net1136));
 sg13g2_a21oi_1 _5856_ (.A1(_1931_),
    .A2(_1932_),
    .Y(_1933_),
    .B1(_3273_));
 sg13g2_o21ai_1 _5857_ (.B1(_1933_),
    .Y(_1934_),
    .A1(net1135),
    .A2(_0786_));
 sg13g2_nand4_1 _5858_ (.B(_1843_),
    .C(_1921_),
    .A(net267),
    .Y(_1935_),
    .D(_1934_));
 sg13g2_nor2_2 _5859_ (.A(_0607_),
    .B(_0616_),
    .Y(_1936_));
 sg13g2_nand2_2 _5860_ (.Y(_1937_),
    .A(_2823_),
    .B(_1936_));
 sg13g2_nor2_1 _5861_ (.A(_0628_),
    .B(_1937_),
    .Y(_1938_));
 sg13g2_nor3_1 _5862_ (.A(_0600_),
    .B(_0628_),
    .C(_1937_),
    .Y(_1939_));
 sg13g2_xnor2_1 _5863_ (.Y(_1940_),
    .A(_0601_),
    .B(_1938_));
 sg13g2_nand2_1 _5864_ (.Y(_1941_),
    .A(net1332),
    .B(_1940_));
 sg13g2_xor2_1 _5865_ (.B(_1940_),
    .A(_0059_),
    .X(_1942_));
 sg13g2_xnor2_1 _5866_ (.Y(_1943_),
    .A(_0628_),
    .B(_1937_));
 sg13g2_a21o_1 _5867_ (.A2(_0616_),
    .A1(net1240),
    .B1(_1936_),
    .X(_1944_));
 sg13g2_nand2_1 _5868_ (.Y(_1945_),
    .A(_2826_),
    .B(net1349));
 sg13g2_nor2_1 _5869_ (.A(_2826_),
    .B(net1349),
    .Y(_1946_));
 sg13g2_nor2_1 _5870_ (.A(net1351),
    .B(_1882_),
    .Y(_1947_));
 sg13g2_a21oi_1 _5871_ (.A1(_1810_),
    .A2(_1945_),
    .Y(_1948_),
    .B1(_1946_));
 sg13g2_o21ai_1 _5872_ (.B1(_1948_),
    .Y(_1949_),
    .A1(net1247),
    .A2(net1347));
 sg13g2_a21oi_1 _5873_ (.A1(_1945_),
    .A2(_1947_),
    .Y(_1950_),
    .B1(_1949_));
 sg13g2_a221oi_1 _5874_ (.B2(net1345),
    .C1(_1950_),
    .B1(_0617_),
    .A1(net1247),
    .Y(_1951_),
    .A2(net1347));
 sg13g2_o21ai_1 _5875_ (.B1(_1937_),
    .Y(_1952_),
    .A1(_0623_),
    .A2(_1936_));
 sg13g2_xor2_1 _5876_ (.B(_1952_),
    .A(net1337),
    .X(_1953_));
 sg13g2_xnor2_1 _5877_ (.Y(_1954_),
    .A(net1340),
    .B(_1944_));
 sg13g2_a21oi_1 _5878_ (.A1(_2871_),
    .A2(_0616_),
    .Y(_1955_),
    .B1(_1951_));
 sg13g2_a22oi_1 _5879_ (.Y(_1956_),
    .B1(_1954_),
    .B2(_1955_),
    .A2(_1944_),
    .A1(net1343));
 sg13g2_a22oi_1 _5880_ (.Y(_1957_),
    .B1(_1952_),
    .B2(net1338),
    .A2(_1943_),
    .A1(net1335));
 sg13g2_o21ai_1 _5881_ (.B1(_1957_),
    .Y(_1958_),
    .A1(_1953_),
    .A2(_1956_));
 sg13g2_o21ai_1 _5882_ (.B1(_1958_),
    .Y(_1959_),
    .A1(net1335),
    .A2(_1943_));
 sg13g2_o21ai_1 _5883_ (.B1(_1941_),
    .Y(_1960_),
    .A1(_1942_),
    .A2(_1959_));
 sg13g2_nor2_1 _5884_ (.A(_0604_),
    .B(_1939_),
    .Y(_1961_));
 sg13g2_inv_1 _5885_ (.Y(_1962_),
    .A(_1961_));
 sg13g2_a22oi_1 _5886_ (.Y(_1963_),
    .B1(_1962_),
    .B2(_2867_),
    .A2(_1939_),
    .A1(net1231));
 sg13g2_nor2_1 _5887_ (.A(net1138),
    .B(_0628_),
    .Y(_1964_));
 sg13g2_xnor2_1 _5888_ (.Y(_1965_),
    .A(net1247),
    .B(_3242_));
 sg13g2_a21oi_1 _5889_ (.A1(_3234_),
    .A2(_1948_),
    .Y(_1966_),
    .B1(_1965_));
 sg13g2_a221oi_1 _5890_ (.B2(net1142),
    .C1(_1966_),
    .B1(_0617_),
    .A1(_0070_),
    .Y(_1967_),
    .A2(_3243_));
 sg13g2_a21oi_1 _5891_ (.A1(net1143),
    .A2(_0616_),
    .Y(_1968_),
    .B1(_1967_));
 sg13g2_o21ai_1 _5892_ (.B1(_1968_),
    .Y(_1969_),
    .A1(net1161),
    .A2(_0606_));
 sg13g2_a22oi_1 _5893_ (.Y(_1970_),
    .B1(_0623_),
    .B2(_3254_),
    .A2(_0606_),
    .A1(net1161));
 sg13g2_a22oi_1 _5894_ (.Y(_1971_),
    .B1(_1969_),
    .B2(_1970_),
    .A2(_0622_),
    .A1(_3255_));
 sg13g2_a22oi_1 _5895_ (.Y(_1972_),
    .B1(_0628_),
    .B2(net1138),
    .A2(_0600_),
    .A1(_3265_));
 sg13g2_o21ai_1 _5896_ (.B1(_1972_),
    .Y(_1973_),
    .A1(_1964_),
    .A2(_1971_));
 sg13g2_a22oi_1 _5897_ (.Y(_1974_),
    .B1(_0604_),
    .B2(net1135),
    .A2(_0601_),
    .A1(net1137));
 sg13g2_o21ai_1 _5898_ (.B1(_3274_),
    .Y(_1975_),
    .A1(net1135),
    .A2(_0604_));
 sg13g2_a21oi_1 _5899_ (.A1(_1973_),
    .A2(_1974_),
    .Y(_1976_),
    .B1(_1975_));
 sg13g2_a221oi_1 _5900_ (.B2(_1960_),
    .C1(_1976_),
    .B1(_1963_),
    .A1(net1328),
    .Y(_1977_),
    .A2(_1961_));
 sg13g2_nand3_1 _5901_ (.B(_1843_),
    .C(_1977_),
    .A(net243),
    .Y(_1978_));
 sg13g2_nand3_1 _5902_ (.B(_0495_),
    .C(_0680_),
    .A(net1235),
    .Y(_1979_));
 sg13g2_nor2_1 _5903_ (.A(_0678_),
    .B(_1979_),
    .Y(_1980_));
 sg13g2_nand2b_1 _5904_ (.Y(_1981_),
    .B(_1980_),
    .A_N(_0676_));
 sg13g2_and2_1 _5905_ (.A(_0693_),
    .B(_1981_),
    .X(_1982_));
 sg13g2_xnor2_1 _5906_ (.Y(_1983_),
    .A(_0676_),
    .B(_1980_));
 sg13g2_xor2_1 _5907_ (.B(_0680_),
    .A(net1160),
    .X(_1984_));
 sg13g2_nand2b_1 _5908_ (.Y(_1985_),
    .B(\pb_x[5] ),
    .A_N(_1984_));
 sg13g2_nand2_1 _5909_ (.Y(_1986_),
    .A(_2886_),
    .B(net1160));
 sg13g2_nand2_1 _5910_ (.Y(_1987_),
    .A(net1347),
    .B(_0499_));
 sg13g2_nor2_1 _5911_ (.A(net1250),
    .B(net1349),
    .Y(_1988_));
 sg13g2_nand2_1 _5912_ (.Y(_1989_),
    .A(net1250),
    .B(net1349));
 sg13g2_o21ai_1 _5913_ (.B1(_1989_),
    .Y(_1990_),
    .A1(_1810_),
    .A2(_1988_));
 sg13g2_xnor2_1 _5914_ (.Y(_1991_),
    .A(_0069_),
    .B(_0499_));
 sg13g2_a22oi_1 _5915_ (.Y(_1992_),
    .B1(_1990_),
    .B2(_1991_),
    .A2(_0499_),
    .A1(net1346));
 sg13g2_xnor2_1 _5916_ (.Y(_1993_),
    .A(net1345),
    .B(net1160));
 sg13g2_o21ai_1 _5917_ (.B1(_1986_),
    .Y(_1994_),
    .A1(_1992_),
    .A2(_1993_));
 sg13g2_nand4_1 _5918_ (.B(_1986_),
    .C(_1987_),
    .A(_1947_),
    .Y(_1995_),
    .D(_1989_));
 sg13g2_o21ai_1 _5919_ (.B1(_0687_),
    .Y(_1996_),
    .A1(_0496_),
    .A2(_0681_));
 sg13g2_nand2_1 _5920_ (.Y(_1997_),
    .A(_1979_),
    .B(_1996_));
 sg13g2_xor2_1 _5921_ (.B(_1984_),
    .A(net1341),
    .X(_1998_));
 sg13g2_nand3_1 _5922_ (.B(_1995_),
    .C(_1998_),
    .A(_1994_),
    .Y(_1999_));
 sg13g2_xor2_1 _5923_ (.B(_1997_),
    .A(net1337),
    .X(_2000_));
 sg13g2_a21oi_1 _5924_ (.A1(_1985_),
    .A2(_1999_),
    .Y(_2001_),
    .B1(_2000_));
 sg13g2_xnor2_1 _5925_ (.Y(_2002_),
    .A(_0678_),
    .B(_1979_));
 sg13g2_a221oi_1 _5926_ (.B2(net1335),
    .C1(_2001_),
    .B1(_2002_),
    .A1(net1339),
    .Y(_2003_),
    .A2(_1997_));
 sg13g2_nor2_1 _5927_ (.A(net1335),
    .B(_2002_),
    .Y(_2004_));
 sg13g2_a21oi_1 _5928_ (.A1(net1331),
    .A2(_1983_),
    .Y(_2005_),
    .B1(_2004_));
 sg13g2_nand2b_1 _5929_ (.Y(_2006_),
    .B(_2005_),
    .A_N(_2003_));
 sg13g2_o21ai_1 _5930_ (.B1(_2006_),
    .Y(_2007_),
    .A1(net1331),
    .A2(_1983_));
 sg13g2_xnor2_1 _5931_ (.Y(_2008_),
    .A(_0058_),
    .B(_1982_));
 sg13g2_a22oi_1 _5932_ (.Y(_2009_),
    .B1(_2007_),
    .B2(_2008_),
    .A2(_1982_),
    .A1(net1328));
 sg13g2_inv_1 _5933_ (.Y(_2010_),
    .A(_2009_));
 sg13g2_o21ai_1 _5934_ (.B1(_2010_),
    .Y(_2011_),
    .A1(_0078_),
    .A2(_1981_));
 sg13g2_nand2_1 _5935_ (.Y(_2012_),
    .A(net1142),
    .B(net1160));
 sg13g2_a22oi_1 _5936_ (.Y(_2013_),
    .B1(_0500_),
    .B2(_3243_),
    .A2(net1188),
    .A1(_2826_));
 sg13g2_xnor2_1 _5937_ (.Y(_2014_),
    .A(_2826_),
    .B(net1188));
 sg13g2_o21ai_1 _5938_ (.B1(_2013_),
    .Y(_2015_),
    .A1(_1780_),
    .A2(_2014_));
 sg13g2_a22oi_1 _5939_ (.Y(_2016_),
    .B1(_0499_),
    .B2(_3242_),
    .A2(_0496_),
    .A1(_3240_));
 sg13g2_a22oi_1 _5940_ (.Y(_2017_),
    .B1(_2015_),
    .B2(_2016_),
    .A2(net1160),
    .A1(net1142));
 sg13g2_o21ai_1 _5941_ (.B1(_3238_),
    .Y(_2018_),
    .A1(_0681_),
    .A2(_2017_));
 sg13g2_a22oi_1 _5942_ (.Y(_2019_),
    .B1(_2017_),
    .B2(_0681_),
    .A2(_0687_),
    .A1(_3255_));
 sg13g2_nand2_1 _5943_ (.Y(_2020_),
    .A(_2018_),
    .B(_2019_));
 sg13g2_nand2b_1 _5944_ (.Y(_2021_),
    .B(net1140),
    .A_N(_0687_));
 sg13g2_nand2b_1 _5945_ (.Y(_2022_),
    .B(_3262_),
    .A_N(_0678_));
 sg13g2_a22oi_1 _5946_ (.Y(_2023_),
    .B1(_2020_),
    .B2(_2021_),
    .A2(_0678_),
    .A1(net1139));
 sg13g2_o21ai_1 _5947_ (.B1(_2022_),
    .Y(_2024_),
    .A1(_3265_),
    .A2(_0676_));
 sg13g2_a22oi_1 _5948_ (.Y(_2025_),
    .B1(_0693_),
    .B2(_3270_),
    .A2(_0676_),
    .A1(_3265_));
 sg13g2_o21ai_1 _5949_ (.B1(_2025_),
    .Y(_2026_),
    .A1(_2023_),
    .A2(_2024_));
 sg13g2_o21ai_1 _5950_ (.B1(_2026_),
    .Y(_2027_),
    .A1(_3270_),
    .A2(_0693_));
 sg13g2_nand2_2 _5951_ (.Y(_2028_),
    .A(_3274_),
    .B(_2027_));
 sg13g2_nand4_1 _5952_ (.B(_1843_),
    .C(_2011_),
    .A(net280),
    .Y(_2029_),
    .D(_2028_));
 sg13g2_nand3_1 _5953_ (.B(_0494_),
    .C(net1160),
    .A(_0490_),
    .Y(_2030_));
 sg13g2_nor2_1 _5954_ (.A(_0513_),
    .B(_2030_),
    .Y(_2031_));
 sg13g2_nand2b_1 _5955_ (.Y(_2032_),
    .B(_2031_),
    .A_N(_0488_));
 sg13g2_nor2b_1 _5956_ (.A(_0520_),
    .B_N(_2032_),
    .Y(_2033_));
 sg13g2_nand2_1 _5957_ (.Y(_2034_),
    .A(net1328),
    .B(_2033_));
 sg13g2_a21o_1 _5958_ (.A2(_0495_),
    .A1(_0494_),
    .B1(_0490_),
    .X(_2035_));
 sg13g2_nand2_1 _5959_ (.Y(_2036_),
    .A(_2030_),
    .B(_2035_));
 sg13g2_xnor2_1 _5960_ (.Y(_2037_),
    .A(net1337),
    .B(_2036_));
 sg13g2_xor2_1 _5961_ (.B(_0495_),
    .A(_0494_),
    .X(_2038_));
 sg13g2_nand2_1 _5962_ (.Y(_2039_),
    .A(net1340),
    .B(_2038_));
 sg13g2_nand2_1 _5963_ (.Y(_2040_),
    .A(_1994_),
    .B(_2039_));
 sg13g2_o21ai_1 _5964_ (.B1(_2040_),
    .Y(_2041_),
    .A1(net1340),
    .A2(_2038_));
 sg13g2_a22oi_1 _5965_ (.Y(_2042_),
    .B1(_2037_),
    .B2(_2041_),
    .A2(_2036_),
    .A1(net1339));
 sg13g2_xnor2_1 _5966_ (.Y(_2043_),
    .A(_0513_),
    .B(_2030_));
 sg13g2_xor2_1 _5967_ (.B(_2043_),
    .A(_0060_),
    .X(_2044_));
 sg13g2_xor2_1 _5968_ (.B(_2031_),
    .A(_0488_),
    .X(_2045_));
 sg13g2_a22oi_1 _5969_ (.Y(_2046_),
    .B1(_2045_),
    .B2(net1332),
    .A2(_2043_),
    .A1(net1335));
 sg13g2_o21ai_1 _5970_ (.B1(_2046_),
    .Y(_2047_),
    .A1(_2042_),
    .A2(_2044_));
 sg13g2_o21ai_1 _5971_ (.B1(_2047_),
    .Y(_2048_),
    .A1(net1332),
    .A2(_2045_));
 sg13g2_xor2_1 _5972_ (.B(_2033_),
    .A(_0058_),
    .X(_2049_));
 sg13g2_o21ai_1 _5973_ (.B1(_2034_),
    .Y(_2050_),
    .A1(_2048_),
    .A2(_2049_));
 sg13g2_o21ai_1 _5974_ (.B1(_2050_),
    .Y(_2051_),
    .A1(_0078_),
    .A2(_2032_));
 sg13g2_nand2_1 _5975_ (.Y(_2052_),
    .A(net1161),
    .B(_0494_));
 sg13g2_a21oi_1 _5976_ (.A1(net1253),
    .A2(net1350),
    .Y(_2053_),
    .B1(_0077_));
 sg13g2_nand3_1 _5977_ (.B(_2013_),
    .C(_2053_),
    .A(_2012_),
    .Y(_2054_));
 sg13g2_o21ai_1 _5978_ (.B1(_2054_),
    .Y(_2055_),
    .A1(_3237_),
    .A2(_0494_));
 sg13g2_o21ai_1 _5979_ (.B1(_2052_),
    .Y(_2056_),
    .A1(_2017_),
    .A2(_2055_));
 sg13g2_o21ai_1 _5980_ (.B1(_2056_),
    .Y(_2057_),
    .A1(net1141),
    .A2(_0490_));
 sg13g2_nor2_1 _5981_ (.A(net1138),
    .B(_0513_),
    .Y(_2058_));
 sg13g2_a21oi_1 _5982_ (.A1(net1141),
    .A2(_0490_),
    .Y(_2059_),
    .B1(_2058_));
 sg13g2_nand2_1 _5983_ (.Y(_2060_),
    .A(net1138),
    .B(_0513_));
 sg13g2_a22oi_1 _5984_ (.Y(_2061_),
    .B1(_2057_),
    .B2(_2059_),
    .A2(_0488_),
    .A1(_3265_));
 sg13g2_nor2_1 _5985_ (.A(_3265_),
    .B(_0488_),
    .Y(_2062_));
 sg13g2_a221oi_1 _5986_ (.B2(_2061_),
    .C1(_2062_),
    .B1(_2060_),
    .A1(net1134),
    .Y(_2063_),
    .A2(_0520_));
 sg13g2_nor2_1 _5987_ (.A(_3273_),
    .B(_2063_),
    .Y(_2064_));
 sg13g2_o21ai_1 _5988_ (.B1(_2064_),
    .Y(_2065_),
    .A1(net1134),
    .A2(_0520_));
 sg13g2_nand4_1 _5989_ (.B(_1843_),
    .C(_2051_),
    .A(net272),
    .Y(_2066_),
    .D(_2065_));
 sg13g2_and4_1 _5990_ (.A(_1935_),
    .B(_1978_),
    .C(_2029_),
    .D(_2066_),
    .X(_2067_));
 sg13g2_nand2_2 _5991_ (.Y(_2068_),
    .A(net1240),
    .B(net1243));
 sg13g2_nand4_1 _5992_ (.B(net1237),
    .C(net1240),
    .A(net1234),
    .Y(_2069_),
    .D(net1242));
 sg13g2_or3_1 _5993_ (.A(_2820_),
    .B(net1228),
    .C(_2069_),
    .X(_2070_));
 sg13g2_nor2_1 _5994_ (.A(_0074_),
    .B(_2069_),
    .Y(_2071_));
 sg13g2_xor2_1 _5995_ (.B(_2071_),
    .A(_0078_),
    .X(_2072_));
 sg13g2_nand2_1 _5996_ (.Y(_2073_),
    .A(net1328),
    .B(_2072_));
 sg13g2_nor2_1 _5997_ (.A(net1235),
    .B(_2068_),
    .Y(_2074_));
 sg13g2_xnor2_1 _5998_ (.Y(_2075_),
    .A(net1235),
    .B(_2068_));
 sg13g2_a21oi_1 _5999_ (.A1(_0479_),
    .A2(_2068_),
    .Y(_2076_),
    .B1(net1340));
 sg13g2_a21oi_1 _6000_ (.A1(_2825_),
    .A2(net1346),
    .Y(_2077_),
    .B1(_1948_));
 sg13g2_a21oi_1 _6001_ (.A1(net1247),
    .A2(_2872_),
    .Y(_2078_),
    .B1(_2077_));
 sg13g2_o21ai_1 _6002_ (.B1(_2078_),
    .Y(_2079_),
    .A1(net1242),
    .A2(net1345));
 sg13g2_a21oi_1 _6003_ (.A1(net1243),
    .A2(net1344),
    .Y(_2080_),
    .B1(_2076_));
 sg13g2_xor2_1 _6004_ (.B(_2075_),
    .A(_0065_),
    .X(_2081_));
 sg13g2_nand3_1 _6005_ (.B(_0479_),
    .C(_2068_),
    .A(net1340),
    .Y(_2082_));
 sg13g2_a21oi_1 _6006_ (.A1(_2079_),
    .A2(_2080_),
    .Y(_2083_),
    .B1(_2081_));
 sg13g2_a22oi_1 _6007_ (.Y(_2084_),
    .B1(_2082_),
    .B2(_2083_),
    .A2(_2075_),
    .A1(net1339));
 sg13g2_xor2_1 _6008_ (.B(_2074_),
    .A(_0061_),
    .X(_2085_));
 sg13g2_xor2_1 _6009_ (.B(_2085_),
    .A(_0060_),
    .X(_2086_));
 sg13g2_xnor2_1 _6010_ (.Y(_2087_),
    .A(_0074_),
    .B(_2069_));
 sg13g2_a22oi_1 _6011_ (.Y(_2088_),
    .B1(_2087_),
    .B2(net1332),
    .A2(_2085_),
    .A1(net1335));
 sg13g2_o21ai_1 _6012_ (.B1(_2088_),
    .Y(_2089_),
    .A1(_2084_),
    .A2(_2086_));
 sg13g2_o21ai_1 _6013_ (.B1(_2089_),
    .Y(_2090_),
    .A1(net1332),
    .A2(_2087_));
 sg13g2_xor2_1 _6014_ (.B(_2072_),
    .A(_0058_),
    .X(_2091_));
 sg13g2_o21ai_1 _6015_ (.B1(_2073_),
    .Y(_2092_),
    .A1(_2090_),
    .A2(_2091_));
 sg13g2_xnor2_1 _6016_ (.Y(_2093_),
    .A(_0070_),
    .B(_3242_));
 sg13g2_and2_1 _6017_ (.A(net1250),
    .B(net1188),
    .X(_2094_));
 sg13g2_nor2_1 _6018_ (.A(_1780_),
    .B(_2053_),
    .Y(_2095_));
 sg13g2_a21oi_1 _6019_ (.A1(_2014_),
    .A2(_2095_),
    .Y(_2096_),
    .B1(_2094_));
 sg13g2_or2_1 _6020_ (.X(_2097_),
    .B(_2096_),
    .A(_2093_));
 sg13g2_a22oi_1 _6021_ (.Y(_2098_),
    .B1(_3243_),
    .B2(net1246),
    .A2(net1142),
    .A1(_2896_));
 sg13g2_xor2_1 _6022_ (.B(net1161),
    .A(_0075_),
    .X(_2099_));
 sg13g2_a221oi_1 _6023_ (.B2(_2098_),
    .C1(_2099_),
    .B1(_2097_),
    .A1(_0076_),
    .Y(_2100_),
    .A2(net1143));
 sg13g2_a21oi_1 _6024_ (.A1(net1239),
    .A2(net1161),
    .Y(_2101_),
    .B1(_2100_));
 sg13g2_xnor2_1 _6025_ (.Y(_2102_),
    .A(net1235),
    .B(_3255_));
 sg13g2_a22oi_1 _6026_ (.Y(_2103_),
    .B1(_3262_),
    .B2(net1234),
    .A2(net1141),
    .A1(net1237));
 sg13g2_o21ai_1 _6027_ (.B1(_2103_),
    .Y(_2104_),
    .A1(_2101_),
    .A2(_2102_));
 sg13g2_nand2_1 _6028_ (.Y(_2105_),
    .A(_0074_),
    .B(_3265_));
 sg13g2_a22oi_1 _6029_ (.Y(_2106_),
    .B1(net1137),
    .B2(_2895_),
    .A2(net1138),
    .A1(net1226));
 sg13g2_nand3_1 _6030_ (.B(_2105_),
    .C(_2106_),
    .A(_2104_),
    .Y(_2107_));
 sg13g2_a22oi_1 _6031_ (.Y(_2108_),
    .B1(net1134),
    .B2(net1231),
    .A2(net1136),
    .A1(net1233));
 sg13g2_a22oi_1 _6032_ (.Y(_2109_),
    .B1(_2107_),
    .B2(_2108_),
    .A2(_3270_),
    .A1(_2820_));
 sg13g2_a22oi_1 _6033_ (.Y(_2110_),
    .B1(_2109_),
    .B2(_3274_),
    .A2(_2092_),
    .A1(_2070_));
 sg13g2_nand3_1 _6034_ (.B(_1843_),
    .C(_2110_),
    .A(net296),
    .Y(_2111_));
 sg13g2_nand3_1 _6035_ (.B(_0870_),
    .C(_0874_),
    .A(_0831_),
    .Y(_2112_));
 sg13g2_or2_1 _6036_ (.X(_2113_),
    .B(_2112_),
    .A(_0868_));
 sg13g2_or2_1 _6037_ (.X(_2114_),
    .B(_2113_),
    .A(_0888_));
 sg13g2_inv_1 _6038_ (.Y(_2115_),
    .A(_2114_));
 sg13g2_nand2_1 _6039_ (.Y(_2116_),
    .A(_0894_),
    .B(_2114_));
 sg13g2_nand3_1 _6040_ (.B(_0894_),
    .C(_2114_),
    .A(net1328),
    .Y(_2117_));
 sg13g2_a21o_1 _6041_ (.A2(_0874_),
    .A1(_0831_),
    .B1(_0870_),
    .X(_2118_));
 sg13g2_and2_1 _6042_ (.A(_2112_),
    .B(_2118_),
    .X(_2119_));
 sg13g2_nand2b_1 _6043_ (.Y(_2120_),
    .B(net1338),
    .A_N(_2119_));
 sg13g2_xnor2_1 _6044_ (.Y(_2121_),
    .A(_0832_),
    .B(_0874_));
 sg13g2_o21ai_1 _6045_ (.B1(_1778_),
    .Y(_2122_),
    .A1(net1341),
    .A2(_2121_));
 sg13g2_xnor2_1 _6046_ (.Y(_2123_),
    .A(net1337),
    .B(_2119_));
 sg13g2_a21oi_1 _6047_ (.A1(net1340),
    .A2(_2121_),
    .Y(_2124_),
    .B1(_2123_));
 sg13g2_o21ai_1 _6048_ (.B1(_2124_),
    .Y(_2125_),
    .A1(_1788_),
    .A2(_2122_));
 sg13g2_xnor2_1 _6049_ (.Y(_2126_),
    .A(_0868_),
    .B(_2112_));
 sg13g2_xor2_1 _6050_ (.B(_2126_),
    .A(_0060_),
    .X(_2127_));
 sg13g2_a21oi_1 _6051_ (.A1(_2120_),
    .A2(_2125_),
    .Y(_2128_),
    .B1(_2127_));
 sg13g2_xnor2_1 _6052_ (.Y(_2129_),
    .A(_0888_),
    .B(_2113_));
 sg13g2_a221oi_1 _6053_ (.B2(net1332),
    .C1(_2128_),
    .B1(_2129_),
    .A1(net1335),
    .Y(_2130_),
    .A2(_2126_));
 sg13g2_xnor2_1 _6054_ (.Y(_2131_),
    .A(_0058_),
    .B(_2116_));
 sg13g2_nor2_1 _6055_ (.A(_2130_),
    .B(_2131_),
    .Y(_2132_));
 sg13g2_o21ai_1 _6056_ (.B1(_2132_),
    .Y(_2133_),
    .A1(net1332),
    .A2(_2129_));
 sg13g2_a22oi_1 _6057_ (.Y(_2134_),
    .B1(_2117_),
    .B2(_2133_),
    .A2(_2115_),
    .A1(net1232));
 sg13g2_nor2_1 _6058_ (.A(net1141),
    .B(_0870_),
    .Y(_2135_));
 sg13g2_o21ai_1 _6059_ (.B1(_1809_),
    .Y(_2136_),
    .A1(_1813_),
    .A2(_1883_));
 sg13g2_nand2_1 _6060_ (.Y(_2137_),
    .A(net1162),
    .B(_0874_));
 sg13g2_a22oi_1 _6061_ (.Y(_2138_),
    .B1(_1808_),
    .B2(_2136_),
    .A2(net1119),
    .A1(net1142));
 sg13g2_nand2b_1 _6062_ (.Y(_2139_),
    .B(_3238_),
    .A_N(_0874_));
 sg13g2_a21oi_1 _6063_ (.A1(_2137_),
    .A2(_2138_),
    .Y(_2140_),
    .B1(_2135_));
 sg13g2_a22oi_1 _6064_ (.Y(_2141_),
    .B1(_2139_),
    .B2(_2140_),
    .A2(_0870_),
    .A1(net1140));
 sg13g2_o21ai_1 _6065_ (.B1(_2141_),
    .Y(_2142_),
    .A1(net1139),
    .A2(_0868_));
 sg13g2_a22oi_1 _6066_ (.Y(_2143_),
    .B1(_0888_),
    .B2(_3265_),
    .A2(_0868_),
    .A1(net1138));
 sg13g2_a22oi_1 _6067_ (.Y(_2144_),
    .B1(_2142_),
    .B2(_2143_),
    .A2(_0887_),
    .A1(net1136));
 sg13g2_o21ai_1 _6068_ (.B1(_2144_),
    .Y(_2145_),
    .A1(_3270_),
    .A2(_0894_));
 sg13g2_nand2_1 _6069_ (.Y(_2146_),
    .A(_3274_),
    .B(_2145_));
 sg13g2_a21oi_2 _6070_ (.B1(_2146_),
    .Y(_2147_),
    .A2(_0894_),
    .A1(_3270_));
 sg13g2_nand2_1 _6071_ (.Y(_2148_),
    .A(net277),
    .B(_1843_));
 sg13g2_or3_1 _6072_ (.A(_2134_),
    .B(_2147_),
    .C(_2148_),
    .X(_2149_));
 sg13g2_and4_2 _6073_ (.A(_1896_),
    .B(_2067_),
    .C(_2111_),
    .D(_2149_),
    .X(_2150_));
 sg13g2_nand2_1 _6074_ (.Y(_2151_),
    .A(_2889_),
    .B(_2890_));
 sg13g2_nor4_2 _6075_ (.A(\pb_y[3] ),
    .B(net1325),
    .C(_1825_),
    .Y(_2152_),
    .D(_2151_));
 sg13g2_inv_1 _6076_ (.Y(_2153_),
    .A(_2152_));
 sg13g2_a21oi_2 _6077_ (.B1(_1833_),
    .Y(_2154_),
    .A2(_2153_),
    .A1(_1839_));
 sg13g2_nand4_1 _6078_ (.B(_2011_),
    .C(_2028_),
    .A(net292),
    .Y(_2155_),
    .D(_2154_));
 sg13g2_nand2_1 _6079_ (.Y(_2156_),
    .A(_2890_),
    .B(_3294_));
 sg13g2_nand4_1 _6080_ (.B(\pb_y[6] ),
    .C(net1323),
    .A(\pb_y[7] ),
    .Y(_2157_),
    .D(_2156_));
 sg13g2_nand2_1 _6081_ (.Y(_2158_),
    .A(net1324),
    .B(_3292_));
 sg13g2_o21ai_1 _6082_ (.B1(_3285_),
    .Y(_2159_),
    .A1(_1835_),
    .A2(_2158_));
 sg13g2_nand3_1 _6083_ (.B(_1826_),
    .C(_2159_),
    .A(_3284_),
    .Y(_2160_));
 sg13g2_and4_2 _6084_ (.A(_1824_),
    .B(_1827_),
    .C(_2157_),
    .D(_2160_),
    .X(_2161_));
 sg13g2_nand4_1 _6085_ (.B(_2051_),
    .C(_2065_),
    .A(net238),
    .Y(_2162_),
    .D(_2161_));
 sg13g2_nand4_1 _6086_ (.B(_2051_),
    .C(_2065_),
    .A(net283),
    .Y(_2163_),
    .D(_2154_));
 sg13g2_nand4_1 _6087_ (.B(_2011_),
    .C(_2028_),
    .A(net318),
    .Y(_2164_),
    .D(_2161_));
 sg13g2_nand3_1 _6088_ (.B(_1977_),
    .C(_2161_),
    .A(net307),
    .Y(_2165_));
 sg13g2_nand3_1 _6089_ (.B(_1977_),
    .C(_2154_),
    .A(net298),
    .Y(_2166_));
 sg13g2_nand4_1 _6090_ (.B(_1921_),
    .C(_1934_),
    .A(net256),
    .Y(_2167_),
    .D(_2161_));
 sg13g2_nand4_1 _6091_ (.B(_1921_),
    .C(_1934_),
    .A(net250),
    .Y(_2168_),
    .D(_2154_));
 sg13g2_nand4_1 _6092_ (.B(_1876_),
    .C(_1895_),
    .A(net270),
    .Y(_2169_),
    .D(_2161_));
 sg13g2_nand4_1 _6093_ (.B(_1876_),
    .C(_1895_),
    .A(net255),
    .Y(_2170_),
    .D(_2154_));
 sg13g2_nand2_1 _6094_ (.Y(_2171_),
    .A(net257),
    .B(_2154_));
 sg13g2_nor3_1 _6095_ (.A(_1806_),
    .B(_1823_),
    .C(_2171_),
    .Y(_2172_));
 sg13g2_nand2_1 _6096_ (.Y(_2173_),
    .A(net290),
    .B(_2161_));
 sg13g2_nor3_1 _6097_ (.A(_1806_),
    .B(_1823_),
    .C(_2173_),
    .Y(_2174_));
 sg13g2_nand2_1 _6098_ (.Y(_2175_),
    .A(net268),
    .B(_2161_));
 sg13g2_nor3_1 _6099_ (.A(_2134_),
    .B(_2147_),
    .C(_2175_),
    .Y(_2176_));
 sg13g2_nand3b_1 _6100_ (.B(_2110_),
    .C(_2154_),
    .Y(_2177_),
    .A_N(_0006_));
 sg13g2_nand3_1 _6101_ (.B(_2110_),
    .C(_2161_),
    .A(net275),
    .Y(_2178_));
 sg13g2_nand2_1 _6102_ (.Y(_2179_),
    .A(\aliens_alive[14] ),
    .B(_2154_));
 sg13g2_or3_1 _6103_ (.A(_2134_),
    .B(_2147_),
    .C(_2179_),
    .X(_2180_));
 sg13g2_nand4_1 _6104_ (.B(_2165_),
    .C(_2167_),
    .A(_2162_),
    .Y(_2181_),
    .D(_2178_));
 sg13g2_nand2_1 _6105_ (.Y(_2182_),
    .A(_2164_),
    .B(_2169_));
 sg13g2_nand4_1 _6106_ (.B(_2166_),
    .C(_2168_),
    .A(_2163_),
    .Y(_2183_),
    .D(_2177_));
 sg13g2_nand3_1 _6107_ (.B(_2170_),
    .C(_2180_),
    .A(_2155_),
    .Y(_2184_));
 sg13g2_or4_1 _6108_ (.A(_2172_),
    .B(_2174_),
    .C(_2183_),
    .D(_2184_),
    .X(_2185_));
 sg13g2_nor4_2 _6109_ (.A(_2176_),
    .B(_2181_),
    .C(_2182_),
    .Y(_2186_),
    .D(_2185_));
 sg13g2_or3_1 _6110_ (.A(\pb_y[9] ),
    .B(_3280_),
    .C(_3309_),
    .X(_2187_));
 sg13g2_inv_1 _6111_ (.Y(_2188_),
    .A(_2187_));
 sg13g2_a21oi_1 _6112_ (.A1(_3305_),
    .A2(_2188_),
    .Y(_2189_),
    .B1(_1826_));
 sg13g2_inv_1 _6113_ (.Y(_2190_),
    .A(_2189_));
 sg13g2_nor3_2 _6114_ (.A(net1325),
    .B(net1326),
    .C(net415),
    .Y(_2191_));
 sg13g2_nor2_1 _6115_ (.A(_2891_),
    .B(_2191_),
    .Y(_2192_));
 sg13g2_xnor2_1 _6116_ (.Y(_2193_),
    .A(_0073_),
    .B(_2192_));
 sg13g2_or2_1 _6117_ (.X(_2194_),
    .B(_2193_),
    .A(_1834_));
 sg13g2_nand2b_1 _6118_ (.Y(_2195_),
    .B(_2194_),
    .A_N(_3281_));
 sg13g2_nor3_1 _6119_ (.A(\pb_y[7] ),
    .B(net1322),
    .C(net401),
    .Y(_2196_));
 sg13g2_nand2_1 _6120_ (.Y(_2197_),
    .A(\pb_y[4] ),
    .B(net1324));
 sg13g2_o21ai_1 _6121_ (.B1(_2196_),
    .Y(_2198_),
    .A1(_3291_),
    .A2(_2197_));
 sg13g2_nand2_2 _6122_ (.Y(_2199_),
    .A(net323),
    .B(_2192_));
 sg13g2_a221oi_1 _6123_ (.B2(net1321),
    .C1(\pb_y[9] ),
    .B1(_2198_),
    .A1(_2190_),
    .Y(_2200_),
    .A2(_2195_));
 sg13g2_nand2_1 _6124_ (.Y(_2201_),
    .A(\aliens_alive[38] ),
    .B(_2200_));
 sg13g2_nor3_1 _6125_ (.A(_2134_),
    .B(_2147_),
    .C(_2201_),
    .Y(_2202_));
 sg13g2_inv_1 _6126_ (.Y(_2203_),
    .A(_2202_));
 sg13g2_nand3_1 _6127_ (.B(_1977_),
    .C(_2200_),
    .A(net309),
    .Y(_2204_));
 sg13g2_nand2_2 _6128_ (.Y(_2205_),
    .A(_2203_),
    .B(_2204_));
 sg13g2_nand4_1 _6129_ (.B(_2011_),
    .C(_2028_),
    .A(net278),
    .Y(_2206_),
    .D(_2200_));
 sg13g2_nand4_1 _6130_ (.B(_2051_),
    .C(_2065_),
    .A(net301),
    .Y(_2207_),
    .D(_2200_));
 sg13g2_nand4_1 _6131_ (.B(_2892_),
    .C(net1326),
    .A(\pb_y[3] ),
    .Y(_2208_),
    .D(_2894_));
 sg13g2_nor2b_1 _6132_ (.A(_3305_),
    .B_N(_2208_),
    .Y(_2209_));
 sg13g2_a21oi_1 _6133_ (.A1(_1828_),
    .A2(_2209_),
    .Y(_2210_),
    .B1(_3279_));
 sg13g2_nor2_2 _6134_ (.A(_1825_),
    .B(_2210_),
    .Y(_2211_));
 sg13g2_nand4_1 _6135_ (.B(_1921_),
    .C(_1934_),
    .A(net242),
    .Y(_2212_),
    .D(_2211_));
 sg13g2_nand4_1 _6136_ (.B(_1921_),
    .C(_1934_),
    .A(net300),
    .Y(_2213_),
    .D(_2200_));
 sg13g2_nand3_1 _6137_ (.B(_1977_),
    .C(_2211_),
    .A(net289),
    .Y(_2214_));
 sg13g2_nand4_1 _6138_ (.B(_2011_),
    .C(_2028_),
    .A(net271),
    .Y(_2215_),
    .D(_2211_));
 sg13g2_nand4_1 _6139_ (.B(_2051_),
    .C(_2065_),
    .A(net269),
    .Y(_2216_),
    .D(_2211_));
 sg13g2_nand4_1 _6140_ (.B(_1876_),
    .C(_1895_),
    .A(net244),
    .Y(_2217_),
    .D(_2211_));
 sg13g2_nand4_1 _6141_ (.B(_1876_),
    .C(_1895_),
    .A(net286),
    .Y(_2218_),
    .D(_2200_));
 sg13g2_nand2_1 _6142_ (.Y(_2219_),
    .A(\aliens_alive[37] ),
    .B(_2200_));
 sg13g2_nor3_1 _6143_ (.A(_1806_),
    .B(_1823_),
    .C(_2219_),
    .Y(_2220_));
 sg13g2_inv_1 _6144_ (.Y(_2221_),
    .A(_2220_));
 sg13g2_nand2_1 _6145_ (.Y(_2222_),
    .A(net265),
    .B(_2211_));
 sg13g2_nor3_1 _6146_ (.A(_1806_),
    .B(_1823_),
    .C(_2222_),
    .Y(_2223_));
 sg13g2_inv_1 _6147_ (.Y(_2224_),
    .A(_2223_));
 sg13g2_nand3_1 _6148_ (.B(_2110_),
    .C(_2200_),
    .A(net276),
    .Y(_2225_));
 sg13g2_nand2_1 _6149_ (.Y(_2226_),
    .A(\aliens_alive[30] ),
    .B(_2211_));
 sg13g2_or3_1 _6150_ (.A(_2134_),
    .B(_2147_),
    .C(_2226_),
    .X(_2227_));
 sg13g2_nand3_1 _6151_ (.B(_2110_),
    .C(_2211_),
    .A(net310),
    .Y(_2228_));
 sg13g2_nand4_1 _6152_ (.B(_2215_),
    .C(_2217_),
    .A(_2206_),
    .Y(_2229_),
    .D(_2227_));
 sg13g2_nand4_1 _6153_ (.B(_2212_),
    .C(_2213_),
    .A(_2207_),
    .Y(_2230_),
    .D(_2216_));
 sg13g2_nand4_1 _6154_ (.B(_2218_),
    .C(_2225_),
    .A(_2214_),
    .Y(_2231_),
    .D(_2228_));
 sg13g2_nor3_1 _6155_ (.A(_2229_),
    .B(_2230_),
    .C(_2231_),
    .Y(_2232_));
 sg13g2_nand3_1 _6156_ (.B(_2224_),
    .C(_2232_),
    .A(_2221_),
    .Y(_2233_));
 sg13g2_nor2_2 _6157_ (.A(_2205_),
    .B(_2233_),
    .Y(_2234_));
 sg13g2_nand4_1 _6158_ (.B(_2150_),
    .C(_2186_),
    .A(_1845_),
    .Y(_2235_),
    .D(_2234_));
 sg13g2_nand2_1 _6159_ (.Y(_2236_),
    .A(net1322),
    .B(_2151_));
 sg13g2_nor2_1 _6160_ (.A(\pb_y[7] ),
    .B(\pb_y[9] ),
    .Y(_2237_));
 sg13g2_a21oi_1 _6161_ (.A1(_2236_),
    .A2(_2237_),
    .Y(_2238_),
    .B1(_1824_));
 sg13g2_nor3_1 _6162_ (.A(_1834_),
    .B(_2187_),
    .C(_2208_),
    .Y(_2239_));
 sg13g2_nor3_2 _6163_ (.A(_2190_),
    .B(_2238_),
    .C(_2239_),
    .Y(_2240_));
 sg13g2_inv_1 _6164_ (.Y(_2241_),
    .A(_2240_));
 sg13g2_nand2_1 _6165_ (.Y(_2242_),
    .A(net1136),
    .B(net1134));
 sg13g2_o21ai_1 _6166_ (.B1(_3242_),
    .Y(_2243_),
    .A1(net1351),
    .A2(_3234_));
 sg13g2_nand3_1 _6167_ (.B(net1142),
    .C(_2243_),
    .A(net1162),
    .Y(_2244_));
 sg13g2_nor2_1 _6168_ (.A(net1140),
    .B(_3262_),
    .Y(_2245_));
 sg13g2_a21oi_1 _6169_ (.A1(_2244_),
    .A2(_2245_),
    .Y(_2246_),
    .B1(_2242_));
 sg13g2_nor3_1 _6170_ (.A(net1330),
    .B(net1333),
    .C(_0384_),
    .Y(_2247_));
 sg13g2_o21ai_1 _6171_ (.B1(net1334),
    .Y(_2248_),
    .A1(net1344),
    .A2(net1346));
 sg13g2_o21ai_1 _6172_ (.B1(_2247_),
    .Y(_2249_),
    .A1(_3258_),
    .A2(_2248_));
 sg13g2_nor3_2 _6173_ (.A(_2241_),
    .B(_2246_),
    .C(_2249_),
    .Y(_2250_));
 sg13g2_nor2_1 _6174_ (.A(net1348),
    .B(net1351),
    .Y(_2251_));
 sg13g2_o21ai_1 _6175_ (.B1(_3243_),
    .Y(_2252_),
    .A1(net1188),
    .A2(_2251_));
 sg13g2_o21ai_1 _6176_ (.B1(_3238_),
    .Y(_2253_),
    .A1(net1143),
    .A2(_2252_));
 sg13g2_nor2_1 _6177_ (.A(net1337),
    .B(_2253_),
    .Y(_2254_));
 sg13g2_nor3_1 _6178_ (.A(net1139),
    .B(_2242_),
    .C(_2254_),
    .Y(_2255_));
 sg13g2_nor3_1 _6179_ (.A(net1338),
    .B(net1343),
    .C(net1348),
    .Y(_2256_));
 sg13g2_nand2b_1 _6180_ (.Y(_2257_),
    .B(net1334),
    .A_N(_2256_));
 sg13g2_nor4_1 _6181_ (.A(net1330),
    .B(net1333),
    .C(_0354_),
    .D(_2255_),
    .Y(_2258_));
 sg13g2_nand4_1 _6182_ (.B(_2248_),
    .C(_2257_),
    .A(_2240_),
    .Y(_2259_),
    .D(_2258_));
 sg13g2_nor3_1 _6183_ (.A(_0069_),
    .B(net1188),
    .C(_2251_),
    .Y(_2260_));
 sg13g2_o21ai_1 _6184_ (.B1(_3238_),
    .Y(_2261_),
    .A1(net1143),
    .A2(_2260_));
 sg13g2_nand4_1 _6185_ (.B(_3262_),
    .C(net1134),
    .A(net1140),
    .Y(_2262_),
    .D(_2261_));
 sg13g2_a21oi_1 _6186_ (.A1(net1346),
    .A2(net1348),
    .Y(_2263_),
    .B1(net1344));
 sg13g2_o21ai_1 _6187_ (.B1(_3258_),
    .Y(_2264_),
    .A1(_2869_),
    .A2(_2263_));
 sg13g2_o21ai_1 _6188_ (.B1(net1333),
    .Y(_2265_),
    .A1(net1334),
    .A2(_2264_));
 sg13g2_nor2_1 _6189_ (.A(net1330),
    .B(_0292_),
    .Y(_2266_));
 sg13g2_nand4_1 _6190_ (.B(_2262_),
    .C(_2265_),
    .A(_2242_),
    .Y(_2267_),
    .D(_2266_));
 sg13g2_nor2_2 _6191_ (.A(_2241_),
    .B(_2267_),
    .Y(_2268_));
 sg13g2_nor3_1 _6192_ (.A(_2235_),
    .B(_2250_),
    .C(_2268_),
    .Y(_2269_));
 sg13g2_a21oi_1 _6193_ (.A1(_2259_),
    .A2(_2269_),
    .Y(_2270_),
    .B1(_1767_));
 sg13g2_nor3_1 _6194_ (.A(net1351),
    .B(_0069_),
    .C(_3234_),
    .Y(_2271_));
 sg13g2_o21ai_1 _6195_ (.B1(net1140),
    .Y(_2272_),
    .A1(net1142),
    .A2(_2271_));
 sg13g2_nor2_1 _6196_ (.A(net1331),
    .B(_3262_),
    .Y(_2273_));
 sg13g2_o21ai_1 _6197_ (.B1(_2273_),
    .Y(_2274_),
    .A1(_3238_),
    .A2(_2272_));
 sg13g2_nor3_1 _6198_ (.A(net1330),
    .B(_2885_),
    .C(_0372_),
    .Y(_2275_));
 sg13g2_a21oi_1 _6199_ (.A1(net1343),
    .A2(net1344),
    .Y(_2276_),
    .B1(net1338));
 sg13g2_nor2_1 _6200_ (.A(_3268_),
    .B(_2276_),
    .Y(_2277_));
 sg13g2_a21oi_2 _6201_ (.B1(_2277_),
    .Y(_2278_),
    .A2(_2274_),
    .A1(net1134));
 sg13g2_nand3_1 _6202_ (.B(_2275_),
    .C(_2278_),
    .A(_2240_),
    .Y(_2279_));
 sg13g2_nor2_2 _6203_ (.A(net1144),
    .B(_2279_),
    .Y(_2280_));
 sg13g2_and2_1 _6204_ (.A(_2885_),
    .B(_1739_),
    .X(_2281_));
 sg13g2_nor2_1 _6205_ (.A(net1322),
    .B(_1829_),
    .Y(_2282_));
 sg13g2_a22oi_1 _6206_ (.Y(_2283_),
    .B1(_2152_),
    .B2(_2282_),
    .A2(_1824_),
    .A1(_2887_));
 sg13g2_o21ai_1 _6207_ (.B1(net1171),
    .Y(_2284_),
    .A1(_1767_),
    .A2(_2283_));
 sg13g2_nor4_1 _6208_ (.A(_2270_),
    .B(_2280_),
    .C(_2281_),
    .D(_2284_),
    .Y(_0109_));
 sg13g2_nor2b_1 _6209_ (.A(_1767_),
    .B_N(_2283_),
    .Y(_2285_));
 sg13g2_nand2b_2 _6210_ (.Y(_2286_),
    .B(_2283_),
    .A_N(_1767_));
 sg13g2_nor2_1 _6211_ (.A(net1158),
    .B(_2285_),
    .Y(_2287_));
 sg13g2_o21ai_1 _6212_ (.B1(net1171),
    .Y(_2288_),
    .A1(net223),
    .A2(_2286_));
 sg13g2_a21oi_1 _6213_ (.A1(_2894_),
    .A2(_2287_),
    .Y(_0110_),
    .B1(_2288_));
 sg13g2_nor2_1 _6214_ (.A(net1326),
    .B(net1158),
    .Y(_2289_));
 sg13g2_o21ai_1 _6215_ (.B1(_2289_),
    .Y(_2290_),
    .A1(net393),
    .A2(_2286_));
 sg13g2_nor3_1 _6216_ (.A(net393),
    .B(_2286_),
    .C(_2289_),
    .Y(_2291_));
 sg13g2_nand2_1 _6217_ (.Y(_2292_),
    .A(net1173),
    .B(_2290_));
 sg13g2_nor2_1 _6218_ (.A(_2291_),
    .B(_2292_),
    .Y(_0111_));
 sg13g2_o21ai_1 _6219_ (.B1(_2892_),
    .Y(_2293_),
    .A1(net1327),
    .A2(_1739_));
 sg13g2_nor3_1 _6220_ (.A(net1326),
    .B(net393),
    .C(_2286_),
    .Y(_2294_));
 sg13g2_o21ai_1 _6221_ (.B1(net1173),
    .Y(_2295_),
    .A1(_2293_),
    .A2(_2294_));
 sg13g2_a21oi_1 _6222_ (.A1(_2293_),
    .A2(_2294_),
    .Y(_0112_),
    .B1(_2295_));
 sg13g2_nor2_1 _6223_ (.A(net1324),
    .B(net1158),
    .Y(_2296_));
 sg13g2_o21ai_1 _6224_ (.B1(_2296_),
    .Y(_2297_),
    .A1(_2191_),
    .A2(_2286_));
 sg13g2_nor3_1 _6225_ (.A(_2191_),
    .B(_2286_),
    .C(_2296_),
    .Y(_2298_));
 sg13g2_nand2_1 _6226_ (.Y(_2299_),
    .A(net1173),
    .B(_2297_));
 sg13g2_nor2_1 _6227_ (.A(_2298_),
    .B(_2299_),
    .Y(_0113_));
 sg13g2_a22oi_1 _6228_ (.Y(_2300_),
    .B1(_2287_),
    .B2(net323),
    .A2(_2285_),
    .A1(_2193_));
 sg13g2_nor2_1 _6229_ (.A(net1165),
    .B(net324),
    .Y(_0114_));
 sg13g2_xnor2_1 _6230_ (.Y(_2301_),
    .A(net359),
    .B(_2199_));
 sg13g2_a22oi_1 _6231_ (.Y(_2302_),
    .B1(_2301_),
    .B2(_2285_),
    .A2(_2287_),
    .A1(net1323));
 sg13g2_nor2_1 _6232_ (.A(net1165),
    .B(net360),
    .Y(_0115_));
 sg13g2_nor2_1 _6233_ (.A(net1322),
    .B(net1158),
    .Y(_2303_));
 sg13g2_o21ai_1 _6234_ (.B1(net359),
    .Y(_2304_),
    .A1(net1323),
    .A2(_2199_));
 sg13g2_or2_1 _6235_ (.X(_2305_),
    .B(_2304_),
    .A(_2286_));
 sg13g2_o21ai_1 _6236_ (.B1(net1171),
    .Y(_2306_),
    .A1(_2303_),
    .A2(_2305_));
 sg13g2_a21oi_1 _6237_ (.A1(_2303_),
    .A2(_2305_),
    .Y(_0116_),
    .B1(_2306_));
 sg13g2_nor2_1 _6238_ (.A(net1322),
    .B(_2305_),
    .Y(_2307_));
 sg13g2_nor2_1 _6239_ (.A(_2887_),
    .B(net1158),
    .Y(_2308_));
 sg13g2_o21ai_1 _6240_ (.B1(net1171),
    .Y(_2309_),
    .A1(_2307_),
    .A2(_2308_));
 sg13g2_a21oi_1 _6241_ (.A1(net312),
    .A2(_2307_),
    .Y(_0117_),
    .B1(_2309_));
 sg13g2_nor2_1 _6242_ (.A(net1321),
    .B(net1158),
    .Y(_2310_));
 sg13g2_nand4_1 _6243_ (.B(net1151),
    .C(_2196_),
    .A(net1327),
    .Y(_2311_),
    .D(_2199_));
 sg13g2_xnor2_1 _6244_ (.Y(_2312_),
    .A(_2310_),
    .B(_2311_));
 sg13g2_nor2_1 _6245_ (.A(_2284_),
    .B(_2312_),
    .Y(_0118_));
 sg13g2_nand2_1 _6246_ (.Y(_2313_),
    .A(net321),
    .B(net1171));
 sg13g2_nor2_1 _6247_ (.A(net1321),
    .B(_2311_),
    .Y(_2314_));
 sg13g2_nor3_1 _6248_ (.A(net1158),
    .B(_2313_),
    .C(_2314_),
    .Y(_0119_));
 sg13g2_nor2_1 _6249_ (.A(net1255),
    .B(_0051_),
    .Y(_2315_));
 sg13g2_nand4_1 _6250_ (.B(\abullet_y[1] ),
    .C(_3025_),
    .A(\abullet_y[3] ),
    .Y(_2316_),
    .D(_2315_));
 sg13g2_nand2b_1 _6251_ (.Y(_2317_),
    .B(_2316_),
    .A_N(_3137_));
 sg13g2_a21o_2 _6252_ (.A2(_2317_),
    .A1(_3022_),
    .B1(_3036_),
    .X(_2318_));
 sg13g2_a21oi_1 _6253_ (.A1(\abullet_x[0] ),
    .A2(_2942_),
    .Y(_2319_),
    .B1(_2938_));
 sg13g2_nand2_1 _6254_ (.Y(_2320_),
    .A(_2937_),
    .B(_2319_));
 sg13g2_nor2_1 _6255_ (.A(_2941_),
    .B(_2320_),
    .Y(_2321_));
 sg13g2_nor3_1 _6256_ (.A(_0034_),
    .B(_2962_),
    .C(_2321_),
    .Y(_2322_));
 sg13g2_a21oi_1 _6257_ (.A1(\abullet_x[5] ),
    .A2(net1316),
    .Y(_2323_),
    .B1(\abullet_x[6] ));
 sg13g2_nor2_1 _6258_ (.A(net1314),
    .B(_0372_),
    .Y(_2324_));
 sg13g2_o21ai_1 _6259_ (.B1(_2324_),
    .Y(_2325_),
    .A1(_2968_),
    .A2(_2323_));
 sg13g2_a21o_2 _6260_ (.A2(_3033_),
    .A1(_3023_),
    .B1(_3032_),
    .X(_2326_));
 sg13g2_o21ai_1 _6261_ (.B1(_2326_),
    .Y(_2327_),
    .A1(_2970_),
    .A2(_2322_));
 sg13g2_nor3_2 _6262_ (.A(_2318_),
    .B(_2325_),
    .C(_2327_),
    .Y(_2328_));
 sg13g2_a21oi_2 _6263_ (.B1(\abullet_y[3] ),
    .Y(_2329_),
    .A2(\abullet_y[1] ),
    .A1(net1255));
 sg13g2_nor3_1 _6264_ (.A(net1254),
    .B(\abullet_y[5] ),
    .C(\abullet_y[4] ),
    .Y(_2330_));
 sg13g2_a21o_1 _6265_ (.A2(_2330_),
    .A1(_2329_),
    .B1(_3016_),
    .X(_2331_));
 sg13g2_nand3b_1 _6266_ (.B(net1319),
    .C(_2331_),
    .Y(_2332_),
    .A_N(\abullet_y[9] ));
 sg13g2_nand2_1 _6267_ (.Y(_2333_),
    .A(_2964_),
    .B(_3031_));
 sg13g2_nor2_1 _6268_ (.A(net1317),
    .B(\abullet_x[0] ),
    .Y(_2334_));
 sg13g2_o21ai_1 _6269_ (.B1(_2943_),
    .Y(_2335_),
    .A1(_3106_),
    .A2(_2334_));
 sg13g2_nor2_1 _6270_ (.A(_0039_),
    .B(_2939_),
    .Y(_2336_));
 sg13g2_o21ai_1 _6271_ (.B1(_2336_),
    .Y(_2337_),
    .A1(_2944_),
    .A2(_2335_));
 sg13g2_and4_1 _6272_ (.A(_2962_),
    .B(_2964_),
    .C(_3031_),
    .D(_2337_),
    .X(_2338_));
 sg13g2_nor3_1 _6273_ (.A(\abullet_x[6] ),
    .B(\abullet_x[5] ),
    .C(net1317),
    .Y(_2339_));
 sg13g2_nand2b_1 _6274_ (.Y(_2340_),
    .B(net1315),
    .A_N(_2339_));
 sg13g2_o21ai_1 _6275_ (.B1(net1315),
    .Y(_2341_),
    .A1(net1316),
    .A2(\abullet_x[3] ));
 sg13g2_nor2_1 _6276_ (.A(net1314),
    .B(\abullet_x[8] ),
    .Y(_2342_));
 sg13g2_nand4_1 _6277_ (.B(_2340_),
    .C(_2341_),
    .A(_2326_),
    .Y(_2343_),
    .D(_2342_));
 sg13g2_nor4_1 _6278_ (.A(_0354_),
    .B(_2318_),
    .C(_2338_),
    .D(_2343_),
    .Y(_2344_));
 sg13g2_o21ai_1 _6279_ (.B1(_2342_),
    .Y(_2345_),
    .A1(_2959_),
    .A2(_2341_));
 sg13g2_nand2b_1 _6280_ (.Y(_2346_),
    .B(_2326_),
    .A_N(_0384_));
 sg13g2_o21ai_1 _6281_ (.B1(_2944_),
    .Y(_2347_),
    .A1(\abullet_x[0] ),
    .A2(_2933_));
 sg13g2_nand3_1 _6282_ (.B(_2943_),
    .C(_2347_),
    .A(_2939_),
    .Y(_2348_));
 sg13g2_nor2_1 _6283_ (.A(_2937_),
    .B(_2962_),
    .Y(_2349_));
 sg13g2_a21oi_1 _6284_ (.A1(_2348_),
    .A2(_2349_),
    .Y(_2350_),
    .B1(_2333_));
 sg13g2_nor4_2 _6285_ (.A(_2318_),
    .B(_2345_),
    .C(_2346_),
    .Y(_2351_),
    .D(_2350_));
 sg13g2_nand3_1 _6286_ (.B(_2862_),
    .C(_2934_),
    .A(_2861_),
    .Y(_2352_));
 sg13g2_nand3_1 _6287_ (.B(\abullet_x[6] ),
    .C(_2352_),
    .A(\abullet_x[8] ),
    .Y(_2353_));
 sg13g2_a21oi_1 _6288_ (.A1(\abullet_x[8] ),
    .A2(net1315),
    .Y(_2354_),
    .B1(net1314));
 sg13g2_nand4_1 _6289_ (.B(_2326_),
    .C(_2353_),
    .A(_0293_),
    .Y(_2355_),
    .D(_2354_));
 sg13g2_a21oi_1 _6290_ (.A1(_2862_),
    .A2(_0045_),
    .Y(_2356_),
    .B1(_2939_));
 sg13g2_nand2_1 _6291_ (.Y(_2357_),
    .A(_2335_),
    .B(_2356_));
 sg13g2_nand3_1 _6292_ (.B(_2962_),
    .C(_2357_),
    .A(_2937_),
    .Y(_2358_));
 sg13g2_a21oi_1 _6293_ (.A1(_2965_),
    .A2(_2358_),
    .Y(_2359_),
    .B1(_2970_));
 sg13g2_nor3_1 _6294_ (.A(_2318_),
    .B(_2355_),
    .C(_2359_),
    .Y(_2360_));
 sg13g2_or4_1 _6295_ (.A(_2328_),
    .B(_2332_),
    .C(_2344_),
    .D(_2360_),
    .X(_2361_));
 sg13g2_nor3_1 _6296_ (.A(_3039_),
    .B(_2351_),
    .C(_2361_),
    .Y(_2362_));
 sg13g2_nand2b_1 _6297_ (.Y(_2363_),
    .B(net345),
    .A_N(net1318));
 sg13g2_nand2_1 _6298_ (.Y(_2364_),
    .A(net1150),
    .B(_2363_));
 sg13g2_nor2_1 _6299_ (.A(_2362_),
    .B(_2364_),
    .Y(_2365_));
 sg13g2_o21ai_1 _6300_ (.B1(net1174),
    .Y(_2366_),
    .A1(net1319),
    .A2(net1149));
 sg13g2_nor2_1 _6301_ (.A(_2365_),
    .B(_2366_),
    .Y(_0120_));
 sg13g2_nand2_1 _6302_ (.Y(_2367_),
    .A(\lfsr[0] ),
    .B(net1149));
 sg13g2_and3_1 _6303_ (.X(_2368_),
    .A(\lfsr[0] ),
    .B(_0030_),
    .C(net1149));
 sg13g2_nand3_1 _6304_ (.B(_0030_),
    .C(net1149),
    .A(net345),
    .Y(_2369_));
 sg13g2_o21ai_1 _6305_ (.B1(net1176),
    .Y(_2370_),
    .A1(net1313),
    .A2(_2369_));
 sg13g2_a21oi_1 _6306_ (.A1(_2866_),
    .A2(_2369_),
    .Y(_0121_),
    .B1(_2370_));
 sg13g2_nand2_1 _6307_ (.Y(_2371_),
    .A(net1252),
    .B(net1311));
 sg13g2_xor2_1 _6308_ (.B(net1311),
    .A(net1252),
    .X(_2372_));
 sg13g2_nand2_1 _6309_ (.Y(_2373_),
    .A(\colRand[0] ),
    .B(_2372_));
 sg13g2_xnor2_1 _6310_ (.Y(_2374_),
    .A(net266),
    .B(_2372_));
 sg13g2_o21ai_1 _6311_ (.B1(net1177),
    .Y(_2375_),
    .A1(net330),
    .A2(net1098));
 sg13g2_a21oi_1 _6312_ (.A1(net1098),
    .A2(_2374_),
    .Y(_0122_),
    .B1(_2375_));
 sg13g2_o21ai_1 _6313_ (.B1(net1177),
    .Y(_2376_),
    .A1(net284),
    .A2(net1099));
 sg13g2_and2_1 _6314_ (.A(net1249),
    .B(net1311),
    .X(_2377_));
 sg13g2_xor2_1 _6315_ (.B(net1311),
    .A(net1249),
    .X(_2378_));
 sg13g2_xnor2_1 _6316_ (.Y(_2379_),
    .A(net1313),
    .B(_2378_));
 sg13g2_and3_1 _6317_ (.X(_2380_),
    .A(_2371_),
    .B(_2373_),
    .C(_2379_));
 sg13g2_a21oi_1 _6318_ (.A1(_2371_),
    .A2(_2373_),
    .Y(_2381_),
    .B1(_2379_));
 sg13g2_nor2_1 _6319_ (.A(_2380_),
    .B(_2381_),
    .Y(_2382_));
 sg13g2_xor2_1 _6320_ (.B(_2382_),
    .A(_0067_),
    .X(_2383_));
 sg13g2_a21oi_1 _6321_ (.A1(net1099),
    .A2(_2383_),
    .Y(_0123_),
    .B1(_2376_));
 sg13g2_o21ai_1 _6322_ (.B1(net1176),
    .Y(_2384_),
    .A1(\abullet_x[3] ),
    .A2(net1099));
 sg13g2_a21oi_1 _6323_ (.A1(net1313),
    .A2(_2378_),
    .Y(_2385_),
    .B1(_2377_));
 sg13g2_nor2_1 _6324_ (.A(net1248),
    .B(net1312),
    .Y(_2386_));
 sg13g2_xor2_1 _6325_ (.B(net1311),
    .A(net1248),
    .X(_2387_));
 sg13g2_nor2_1 _6326_ (.A(_2385_),
    .B(_2387_),
    .Y(_2388_));
 sg13g2_xnor2_1 _6327_ (.Y(_2389_),
    .A(_2385_),
    .B(_2387_));
 sg13g2_inv_1 _6328_ (.Y(_2390_),
    .A(_2389_));
 sg13g2_xor2_1 _6329_ (.B(_2389_),
    .A(net1313),
    .X(_2391_));
 sg13g2_nor2_1 _6330_ (.A(net1310),
    .B(_2381_),
    .Y(_2392_));
 sg13g2_o21ai_1 _6331_ (.B1(_2391_),
    .Y(_2393_),
    .A1(_2380_),
    .A2(_2392_));
 sg13g2_nor3_1 _6332_ (.A(_2380_),
    .B(_2391_),
    .C(_2392_),
    .Y(_2394_));
 sg13g2_inv_1 _6333_ (.Y(_2395_),
    .A(_2394_));
 sg13g2_nand2_1 _6334_ (.Y(_2396_),
    .A(_2393_),
    .B(_2395_));
 sg13g2_xnor2_1 _6335_ (.Y(_2397_),
    .A(net319),
    .B(_2396_));
 sg13g2_a21oi_1 _6336_ (.A1(net1099),
    .A2(_2397_),
    .Y(_0124_),
    .B1(_2384_));
 sg13g2_a21oi_1 _6337_ (.A1(net1313),
    .A2(_2390_),
    .Y(_2398_),
    .B1(_2388_));
 sg13g2_and2_1 _6338_ (.A(net1245),
    .B(net1312),
    .X(_2399_));
 sg13g2_xor2_1 _6339_ (.B(net1312),
    .A(net1245),
    .X(_2400_));
 sg13g2_and2_1 _6340_ (.A(net1313),
    .B(_2400_),
    .X(_2401_));
 sg13g2_xnor2_1 _6341_ (.Y(_2402_),
    .A(net1313),
    .B(_2400_));
 sg13g2_xor2_1 _6342_ (.B(_2402_),
    .A(_2386_),
    .X(_2403_));
 sg13g2_nand2_1 _6343_ (.Y(_2404_),
    .A(\colRand[2] ),
    .B(_2403_));
 sg13g2_xnor2_1 _6344_ (.Y(_2405_),
    .A(net1310),
    .B(_2403_));
 sg13g2_nor2_1 _6345_ (.A(_2398_),
    .B(_2405_),
    .Y(_2406_));
 sg13g2_xor2_1 _6346_ (.B(_2405_),
    .A(_2398_),
    .X(_2407_));
 sg13g2_a21oi_1 _6347_ (.A1(net1310),
    .A2(_2393_),
    .Y(_2408_),
    .B1(_2394_));
 sg13g2_inv_1 _6348_ (.Y(_2409_),
    .A(_2408_));
 sg13g2_xor2_1 _6349_ (.B(_2408_),
    .A(_2407_),
    .X(_2410_));
 sg13g2_o21ai_1 _6350_ (.B1(net1177),
    .Y(_2411_),
    .A1(net288),
    .A2(net1098));
 sg13g2_a21oi_1 _6351_ (.A1(net1098),
    .A2(_2410_),
    .Y(_0125_),
    .B1(_2411_));
 sg13g2_o21ai_1 _6352_ (.B1(_2404_),
    .Y(_2412_),
    .A1(_2386_),
    .A2(_2402_));
 sg13g2_nand2_1 _6353_ (.Y(_2413_),
    .A(net1239),
    .B(net1311));
 sg13g2_xor2_1 _6354_ (.B(net1312),
    .A(net1239),
    .X(_2414_));
 sg13g2_o21ai_1 _6355_ (.B1(_2414_),
    .Y(_2415_),
    .A1(_2399_),
    .A2(_2401_));
 sg13g2_or3_1 _6356_ (.A(_2399_),
    .B(_2401_),
    .C(_2414_),
    .X(_2416_));
 sg13g2_and2_1 _6357_ (.A(_2415_),
    .B(_2416_),
    .X(_2417_));
 sg13g2_nand2_1 _6358_ (.Y(_2418_),
    .A(net1310),
    .B(_2417_));
 sg13g2_xnor2_1 _6359_ (.Y(_2419_),
    .A(net1310),
    .B(_2417_));
 sg13g2_nand2b_1 _6360_ (.Y(_2420_),
    .B(_2412_),
    .A_N(_2419_));
 sg13g2_xor2_1 _6361_ (.B(_2419_),
    .A(_2412_),
    .X(_2421_));
 sg13g2_a21oi_1 _6362_ (.A1(_2407_),
    .A2(_2409_),
    .Y(_2422_),
    .B1(_2406_));
 sg13g2_xnor2_1 _6363_ (.Y(_2423_),
    .A(_2421_),
    .B(_2422_));
 sg13g2_o21ai_1 _6364_ (.B1(net1176),
    .Y(_2424_),
    .A1(net365),
    .A2(net1100));
 sg13g2_a21oi_1 _6365_ (.A1(net1100),
    .A2(_2423_),
    .Y(_0126_),
    .B1(_2424_));
 sg13g2_xor2_1 _6366_ (.B(_2413_),
    .A(net1236),
    .X(_2425_));
 sg13g2_nand2_1 _6367_ (.Y(_2426_),
    .A(net1310),
    .B(_2425_));
 sg13g2_xnor2_1 _6368_ (.Y(_2427_),
    .A(net1310),
    .B(_2425_));
 sg13g2_a21oi_1 _6369_ (.A1(_2415_),
    .A2(_2418_),
    .Y(_2428_),
    .B1(_2427_));
 sg13g2_nand3_1 _6370_ (.B(_2418_),
    .C(_2427_),
    .A(_2415_),
    .Y(_2429_));
 sg13g2_nor2b_1 _6371_ (.A(_2428_),
    .B_N(_2429_),
    .Y(_2430_));
 sg13g2_o21ai_1 _6372_ (.B1(_2420_),
    .Y(_2431_),
    .A1(_2421_),
    .A2(_2422_));
 sg13g2_xnor2_1 _6373_ (.Y(_2432_),
    .A(_2430_),
    .B(_2431_));
 sg13g2_o21ai_1 _6374_ (.B1(net1176),
    .Y(_2433_),
    .A1(net380),
    .A2(net1100));
 sg13g2_a21oi_1 _6375_ (.A1(net1100),
    .A2(_2432_),
    .Y(_0127_),
    .B1(_2433_));
 sg13g2_nand3_1 _6376_ (.B(net1239),
    .C(net1311),
    .A(net1238),
    .Y(_2434_));
 sg13g2_a21oi_2 _6377_ (.B1(net1227),
    .Y(_2435_),
    .A2(_2434_),
    .A1(_2426_));
 sg13g2_nand3_1 _6378_ (.B(_2426_),
    .C(_2434_),
    .A(net1227),
    .Y(_2436_));
 sg13g2_nor2b_1 _6379_ (.A(_2435_),
    .B_N(_2436_),
    .Y(_2437_));
 sg13g2_a21o_1 _6380_ (.A2(_2431_),
    .A1(_2430_),
    .B1(_2428_),
    .X(_2438_));
 sg13g2_and2_1 _6381_ (.A(_2437_),
    .B(_2438_),
    .X(_2439_));
 sg13g2_xnor2_1 _6382_ (.Y(_2440_),
    .A(_2437_),
    .B(_2438_));
 sg13g2_o21ai_1 _6383_ (.B1(net1174),
    .Y(_2441_),
    .A1(net1315),
    .A2(net1100));
 sg13g2_a21oi_1 _6384_ (.A1(net1100),
    .A2(_2440_),
    .Y(_0128_),
    .B1(_2441_));
 sg13g2_xnor2_1 _6385_ (.Y(_2442_),
    .A(_0074_),
    .B(_2435_));
 sg13g2_xnor2_1 _6386_ (.Y(_2443_),
    .A(_2439_),
    .B(_2442_));
 sg13g2_o21ai_1 _6387_ (.B1(net1174),
    .Y(_2444_),
    .A1(net367),
    .A2(net1101));
 sg13g2_a21oi_1 _6388_ (.A1(net1101),
    .A2(_2443_),
    .Y(_0129_),
    .B1(_2444_));
 sg13g2_o21ai_1 _6389_ (.B1(net1174),
    .Y(_2445_),
    .A1(net1314),
    .A2(net1101));
 sg13g2_a22oi_1 _6390_ (.Y(_2446_),
    .B1(_2439_),
    .B2(_2442_),
    .A2(_2435_),
    .A1(net1233));
 sg13g2_xnor2_1 _6391_ (.Y(_2447_),
    .A(_0078_),
    .B(_2446_));
 sg13g2_a21oi_1 _6392_ (.A1(net1101),
    .A2(_2447_),
    .Y(_0130_),
    .B1(_2445_));
 sg13g2_xor2_1 _6393_ (.B(net261),
    .A(net279),
    .X(_2448_));
 sg13g2_xor2_1 _6394_ (.B(\lfsr[3] ),
    .A(net302),
    .X(_2449_));
 sg13g2_xnor2_1 _6395_ (.Y(_2450_),
    .A(_2448_),
    .B(_2449_));
 sg13g2_a21oi_1 _6396_ (.A1(net345),
    .A2(net1146),
    .Y(_2451_),
    .B1(net1168));
 sg13g2_o21ai_1 _6397_ (.B1(_2451_),
    .Y(_0131_),
    .A1(net1146),
    .A2(_2450_));
 sg13g2_nand2_1 _6398_ (.Y(_2452_),
    .A(net248),
    .B(net1144));
 sg13g2_a21oi_1 _6399_ (.A1(_2367_),
    .A2(_2452_),
    .Y(_0132_),
    .B1(net1166));
 sg13g2_a21oi_1 _6400_ (.A1(net248),
    .A2(net1149),
    .Y(_2453_),
    .B1(net1167));
 sg13g2_o21ai_1 _6401_ (.B1(_2453_),
    .Y(_0133_),
    .A1(_2858_),
    .A2(net1149));
 sg13g2_o21ai_1 _6402_ (.B1(net1170),
    .Y(_2454_),
    .A1(\lfsr[3] ),
    .A2(net1149));
 sg13g2_a21oi_1 _6403_ (.A1(_2858_),
    .A2(net1149),
    .Y(_0134_),
    .B1(_2454_));
 sg13g2_o21ai_1 _6404_ (.B1(net1176),
    .Y(_2455_),
    .A1(\lfsr[3] ),
    .A2(net1146));
 sg13g2_a21oi_1 _6405_ (.A1(_2857_),
    .A2(net1146),
    .Y(_0135_),
    .B1(_2455_));
 sg13g2_a21oi_1 _6406_ (.A1(net261),
    .A2(net1154),
    .Y(_2456_),
    .B1(net1168));
 sg13g2_o21ai_1 _6407_ (.B1(_2456_),
    .Y(_0136_),
    .A1(_2856_),
    .A2(net1154));
 sg13g2_o21ai_1 _6408_ (.B1(net1177),
    .Y(_2457_),
    .A1(net273),
    .A2(net1154));
 sg13g2_a21oi_1 _6409_ (.A1(_2856_),
    .A2(net1154),
    .Y(_0137_),
    .B1(_2457_));
 sg13g2_a21oi_1 _6410_ (.A1(net302),
    .A2(net1146),
    .Y(_2458_),
    .B1(net1168));
 sg13g2_o21ai_1 _6411_ (.B1(_2458_),
    .Y(_0138_),
    .A1(_2855_),
    .A2(net1146));
 sg13g2_o21ai_1 _6412_ (.B1(net313),
    .Y(_2459_),
    .A1(net245),
    .A2(net305));
 sg13g2_a21oi_1 _6413_ (.A1(net248),
    .A2(_2459_),
    .Y(_2460_),
    .B1(_2369_));
 sg13g2_o21ai_1 _6414_ (.B1(net1170),
    .Y(_2461_),
    .A1(net305),
    .A2(net1101));
 sg13g2_nor2_1 _6415_ (.A(_2460_),
    .B(_2461_),
    .Y(_0139_));
 sg13g2_a21oi_1 _6416_ (.A1(net233),
    .A2(_2459_),
    .Y(_2462_),
    .B1(_2369_));
 sg13g2_o21ai_1 _6417_ (.B1(net1170),
    .Y(_2463_),
    .A1(net245),
    .A2(net1101));
 sg13g2_nor2_1 _6418_ (.A(_2462_),
    .B(_2463_),
    .Y(_0140_));
 sg13g2_nor2b_1 _6419_ (.A(\lfsr[3] ),
    .B_N(_2459_),
    .Y(_2464_));
 sg13g2_o21ai_1 _6420_ (.B1(net1170),
    .Y(_2465_),
    .A1(net313),
    .A2(net1101));
 sg13g2_a21oi_1 _6421_ (.A1(net1101),
    .A2(_2464_),
    .Y(_0141_),
    .B1(_2465_));
 sg13g2_o21ai_1 _6422_ (.B1(net1177),
    .Y(_2466_),
    .A1(net1313),
    .A2(net1099));
 sg13g2_a21oi_1 _6423_ (.A1(_2857_),
    .A2(net1099),
    .Y(_0142_),
    .B1(_2466_));
 sg13g2_o21ai_1 _6424_ (.B1(net1177),
    .Y(_2467_),
    .A1(net1311),
    .A2(net1098));
 sg13g2_a21oi_1 _6425_ (.A1(_2856_),
    .A2(net1098),
    .Y(_0143_),
    .B1(_2467_));
 sg13g2_o21ai_1 _6426_ (.B1(net1177),
    .Y(_2468_),
    .A1(net1310),
    .A2(net1098));
 sg13g2_a21oi_1 _6427_ (.A1(_2855_),
    .A2(net1098),
    .Y(_0144_),
    .B1(_2468_));
 sg13g2_nand3_1 _6428_ (.B(_2930_),
    .C(net1151),
    .A(net1327),
    .Y(_2469_));
 sg13g2_o21ai_1 _6429_ (.B1(net1416),
    .Y(_2470_),
    .A1(_2235_),
    .A2(_2469_));
 sg13g2_a21o_1 _6430_ (.A2(_1767_),
    .A1(net254),
    .B1(_2470_),
    .X(_2471_));
 sg13g2_or2_1 _6431_ (.X(_2472_),
    .B(_2470_),
    .A(_2469_));
 sg13g2_o21ai_1 _6432_ (.B1(net383),
    .Y(_2473_),
    .A1(_2205_),
    .A2(_2233_));
 sg13g2_xor2_1 _6433_ (.B(net1079),
    .A(\draw_score_inst.score[1] ),
    .X(_2474_));
 sg13g2_nand2_1 _6434_ (.Y(_2475_),
    .A(net1077),
    .B(_2474_));
 sg13g2_a21oi_1 _6435_ (.A1(_2473_),
    .A2(_2475_),
    .Y(_2476_),
    .B1(net1074));
 sg13g2_a21o_1 _6436_ (.A2(net1075),
    .A1(\draw_score_inst.score[1] ),
    .B1(_2476_),
    .X(_0145_));
 sg13g2_nand2_1 _6437_ (.Y(_2477_),
    .A(net335),
    .B(net1075));
 sg13g2_nand2_2 _6438_ (.Y(_2478_),
    .A(\draw_score_inst.score[2] ),
    .B(\draw_score_inst.score[1] ));
 sg13g2_nand2b_1 _6439_ (.Y(_2479_),
    .B(_2478_),
    .A_N(_2924_));
 sg13g2_nor2_1 _6440_ (.A(net1077),
    .B(_2479_),
    .Y(_2480_));
 sg13g2_mux2_1 _6441_ (.A0(_0026_),
    .A1(_2479_),
    .S(net1079),
    .X(_2481_));
 sg13g2_a21oi_1 _6442_ (.A1(net1077),
    .A2(_2481_),
    .Y(_2482_),
    .B1(_2480_));
 sg13g2_o21ai_1 _6443_ (.B1(_2477_),
    .Y(_0146_),
    .A1(net1074),
    .A2(_2482_));
 sg13g2_and2_1 _6444_ (.A(net399),
    .B(net1075),
    .X(_2483_));
 sg13g2_nand2_1 _6445_ (.Y(_2484_),
    .A(_2924_),
    .B(net1079));
 sg13g2_o21ai_1 _6446_ (.B1(_2484_),
    .Y(_2485_),
    .A1(_2899_),
    .A2(net1079));
 sg13g2_xnor2_1 _6447_ (.Y(_2486_),
    .A(\draw_score_inst.score[3] ),
    .B(_2485_));
 sg13g2_nand2_1 _6448_ (.Y(_2487_),
    .A(_0018_),
    .B(_2478_));
 sg13g2_xor2_1 _6449_ (.B(_2478_),
    .A(_0018_),
    .X(_2488_));
 sg13g2_mux2_1 _6450_ (.A0(_2486_),
    .A1(_2488_),
    .S(_2233_),
    .X(_2489_));
 sg13g2_nand2b_1 _6451_ (.Y(_2490_),
    .B(_2489_),
    .A_N(_2205_));
 sg13g2_a21oi_1 _6452_ (.A1(_2205_),
    .A2(_2488_),
    .Y(_2491_),
    .B1(net1074));
 sg13g2_a21o_1 _6453_ (.A2(_2491_),
    .A1(_2490_),
    .B1(_2483_),
    .X(_0147_));
 sg13g2_nand2_1 _6454_ (.Y(_2492_),
    .A(net342),
    .B(_2471_));
 sg13g2_nand2_1 _6455_ (.Y(_2493_),
    .A(_2901_),
    .B(_2925_));
 sg13g2_and2_1 _6456_ (.A(net1078),
    .B(_2493_),
    .X(_2494_));
 sg13g2_o21ai_1 _6457_ (.B1(_2494_),
    .Y(_2495_),
    .A1(_2901_),
    .A2(_2925_));
 sg13g2_nand2_2 _6458_ (.Y(_2496_),
    .A(\draw_score_inst.score[3] ),
    .B(\draw_score_inst.score[2] ));
 sg13g2_a21oi_1 _6459_ (.A1(_0024_),
    .A2(_2496_),
    .Y(_2497_),
    .B1(net1078));
 sg13g2_o21ai_1 _6460_ (.B1(_2497_),
    .Y(_2498_),
    .A1(_0024_),
    .A2(_2496_));
 sg13g2_nand2_1 _6461_ (.Y(_2499_),
    .A(_2495_),
    .B(_2498_));
 sg13g2_xnor2_1 _6462_ (.Y(_2500_),
    .A(_0024_),
    .B(_2487_));
 sg13g2_nand2_1 _6463_ (.Y(_2501_),
    .A(net1077),
    .B(_2499_));
 sg13g2_o21ai_1 _6464_ (.B1(_2501_),
    .Y(_2502_),
    .A1(net1077),
    .A2(_2500_));
 sg13g2_o21ai_1 _6465_ (.B1(_2492_),
    .Y(_0148_),
    .A1(_2472_),
    .A2(_2502_));
 sg13g2_nand2_1 _6466_ (.Y(_2503_),
    .A(net1309),
    .B(net1075));
 sg13g2_a21oi_2 _6467_ (.B1(_2901_),
    .Y(_2504_),
    .A2(_2478_),
    .A1(_2898_));
 sg13g2_or2_1 _6468_ (.X(_2505_),
    .B(_2497_),
    .A(_2494_));
 sg13g2_mux2_1 _6469_ (.A0(_2504_),
    .A1(_2505_),
    .S(net1076),
    .X(_2506_));
 sg13g2_xnor2_1 _6470_ (.Y(_2507_),
    .A(_2913_),
    .B(_2506_));
 sg13g2_o21ai_1 _6471_ (.B1(_2503_),
    .Y(_0149_),
    .A1(net1074),
    .A2(_2507_));
 sg13g2_nand2_1 _6472_ (.Y(_2508_),
    .A(net232),
    .B(net1075));
 sg13g2_nand3_1 _6473_ (.B(net1308),
    .C(_2504_),
    .A(net1309),
    .Y(_2509_));
 sg13g2_a21o_1 _6474_ (.A2(_2504_),
    .A1(net1309),
    .B1(net1308),
    .X(_2510_));
 sg13g2_and2_1 _6475_ (.A(_2509_),
    .B(_2510_),
    .X(_2511_));
 sg13g2_nand3_1 _6476_ (.B(net1308),
    .C(_2493_),
    .A(net1309),
    .Y(_2512_));
 sg13g2_a21o_1 _6477_ (.A2(_2493_),
    .A1(net1309),
    .B1(net1308),
    .X(_2513_));
 sg13g2_nand3_1 _6478_ (.B(_2512_),
    .C(_2513_),
    .A(net1078),
    .Y(_2514_));
 sg13g2_a21oi_2 _6479_ (.B1(_2900_),
    .Y(_2515_),
    .A2(_2496_),
    .A1(_2901_));
 sg13g2_xnor2_1 _6480_ (.Y(_2516_),
    .A(_0022_),
    .B(_2515_));
 sg13g2_nand2b_1 _6481_ (.Y(_2517_),
    .B(_2516_),
    .A_N(net1078));
 sg13g2_nand3_1 _6482_ (.B(_2514_),
    .C(_2517_),
    .A(net1076),
    .Y(_2518_));
 sg13g2_o21ai_1 _6483_ (.B1(_2518_),
    .Y(_2519_),
    .A1(net1077),
    .A2(_2511_));
 sg13g2_o21ai_1 _6484_ (.B1(_2508_),
    .Y(_0150_),
    .A1(net1074),
    .A2(_2519_));
 sg13g2_nand2_1 _6485_ (.Y(_2520_),
    .A(net1307),
    .B(net1075));
 sg13g2_nor2_1 _6486_ (.A(net1306),
    .B(_2515_),
    .Y(_2521_));
 sg13g2_nor2b_1 _6487_ (.A(_2926_),
    .B_N(_2515_),
    .Y(_2522_));
 sg13g2_or4_1 _6488_ (.A(_1582_),
    .B(net1078),
    .C(_2521_),
    .D(_2522_),
    .X(_2523_));
 sg13g2_xnor2_1 _6489_ (.Y(_2524_),
    .A(net1306),
    .B(_2512_));
 sg13g2_nand2_1 _6490_ (.Y(_2525_),
    .A(net1078),
    .B(_2524_));
 sg13g2_nand3_1 _6491_ (.B(_2523_),
    .C(_2525_),
    .A(net1076),
    .Y(_2526_));
 sg13g2_xnor2_1 _6492_ (.Y(_2527_),
    .A(net1306),
    .B(_2509_));
 sg13g2_o21ai_1 _6493_ (.B1(_2526_),
    .Y(_2528_),
    .A1(net1076),
    .A2(_2527_));
 sg13g2_o21ai_1 _6494_ (.B1(_2520_),
    .Y(_0151_),
    .A1(net1074),
    .A2(_2528_));
 sg13g2_nor2b_1 _6495_ (.A(net1078),
    .B_N(_2522_),
    .Y(_2529_));
 sg13g2_nor2_1 _6496_ (.A(_0021_),
    .B(_2512_),
    .Y(_2530_));
 sg13g2_a21o_1 _6497_ (.A2(_2530_),
    .A1(net1078),
    .B1(_2529_),
    .X(_2531_));
 sg13g2_nor3_1 _6498_ (.A(_0021_),
    .B(net1076),
    .C(_2509_),
    .Y(_2532_));
 sg13g2_a21o_1 _6499_ (.A2(_2531_),
    .A1(net1076),
    .B1(_2532_),
    .X(_2533_));
 sg13g2_nand2_1 _6500_ (.Y(_2534_),
    .A(net1305),
    .B(net1075));
 sg13g2_xnor2_1 _6501_ (.Y(_2535_),
    .A(net1305),
    .B(_2533_));
 sg13g2_o21ai_1 _6502_ (.B1(_2534_),
    .Y(_0152_),
    .A1(net1074),
    .A2(_2535_));
 sg13g2_nor3_2 _6503_ (.A(_2900_),
    .B(_2903_),
    .C(_2926_),
    .Y(_2536_));
 sg13g2_a22oi_1 _6504_ (.Y(_2537_),
    .B1(_2536_),
    .B2(_2494_),
    .A2(_2529_),
    .A1(_2910_));
 sg13g2_o21ai_1 _6505_ (.B1(net1076),
    .Y(_2538_),
    .A1(net1304),
    .A2(_2537_));
 sg13g2_a21oi_1 _6506_ (.A1(net1304),
    .A2(_2537_),
    .Y(_2539_),
    .B1(_2538_));
 sg13g2_nand3_1 _6507_ (.B(_2504_),
    .C(_2536_),
    .A(net1303),
    .Y(_2540_));
 sg13g2_a21o_1 _6508_ (.A2(_2536_),
    .A1(_2504_),
    .B1(net1303),
    .X(_2541_));
 sg13g2_a21oi_1 _6509_ (.A1(_2540_),
    .A2(_2541_),
    .Y(_2542_),
    .B1(net1076));
 sg13g2_nor3_1 _6510_ (.A(net1074),
    .B(_2539_),
    .C(_2542_),
    .Y(_2543_));
 sg13g2_a21o_1 _6511_ (.A2(net1075),
    .A1(net1303),
    .B1(_2543_),
    .X(_0153_));
 sg13g2_nor4_1 _6512_ (.A(\draw_score_inst.digit_health[1] ),
    .B(net258),
    .C(net1166),
    .D(net1144),
    .Y(_2544_));
 sg13g2_a21o_1 _6513_ (.A2(_2929_),
    .A1(net253),
    .B1(net259),
    .X(_0154_));
 sg13g2_nand2b_1 _6514_ (.Y(_2545_),
    .B(net1151),
    .A_N(_0054_));
 sg13g2_o21ai_1 _6515_ (.B1(net296),
    .Y(_2546_),
    .A1(_2111_),
    .A2(net1096));
 sg13g2_nand2_1 _6516_ (.Y(_0155_),
    .A(net1183),
    .B(_2546_));
 sg13g2_o21ai_1 _6517_ (.B1(net267),
    .Y(_2547_),
    .A1(_1935_),
    .A2(net1097));
 sg13g2_nand2_1 _6518_ (.Y(_0156_),
    .A(net1183),
    .B(_2547_));
 sg13g2_o21ai_1 _6519_ (.B1(net239),
    .Y(_2548_),
    .A1(_1896_),
    .A2(net1096));
 sg13g2_nand2_1 _6520_ (.Y(_0157_),
    .A(net1183),
    .B(_2548_));
 sg13g2_o21ai_1 _6521_ (.B1(net280),
    .Y(_2549_),
    .A1(_2029_),
    .A2(net1096));
 sg13g2_nand2_1 _6522_ (.Y(_0158_),
    .A(net1183),
    .B(_2549_));
 sg13g2_o21ai_1 _6523_ (.B1(net272),
    .Y(_2550_),
    .A1(_2066_),
    .A2(net1097));
 sg13g2_nand2_1 _6524_ (.Y(_0159_),
    .A(net1183),
    .B(_2550_));
 sg13g2_o21ai_1 _6525_ (.B1(net247),
    .Y(_2551_),
    .A1(_1845_),
    .A2(net1096));
 sg13g2_nand2_1 _6526_ (.Y(_0160_),
    .A(net1182),
    .B(_2551_));
 sg13g2_o21ai_1 _6527_ (.B1(net277),
    .Y(_2552_),
    .A1(_2149_),
    .A2(net1096));
 sg13g2_nand2_1 _6528_ (.Y(_0161_),
    .A(net1183),
    .B(_2552_));
 sg13g2_o21ai_1 _6529_ (.B1(net243),
    .Y(_2553_),
    .A1(_1978_),
    .A2(net1096));
 sg13g2_nand2_1 _6530_ (.Y(_0162_),
    .A(net1183),
    .B(_2553_));
 sg13g2_o21ai_1 _6531_ (.B1(net227),
    .Y(_2554_),
    .A1(_2177_),
    .A2(net1096));
 sg13g2_nand2_1 _6532_ (.Y(_0163_),
    .A(net1182),
    .B(net228));
 sg13g2_o21ai_1 _6533_ (.B1(net250),
    .Y(_2555_),
    .A1(_2168_),
    .A2(net1095));
 sg13g2_nand2_1 _6534_ (.Y(_0164_),
    .A(net1182),
    .B(_2555_));
 sg13g2_o21ai_1 _6535_ (.B1(net255),
    .Y(_2556_),
    .A1(_2170_),
    .A2(net1095));
 sg13g2_nand2_1 _6536_ (.Y(_0165_),
    .A(net1182),
    .B(_2556_));
 sg13g2_o21ai_1 _6537_ (.B1(net292),
    .Y(_2557_),
    .A1(_2155_),
    .A2(net1095));
 sg13g2_nand2_1 _6538_ (.Y(_0166_),
    .A(net1180),
    .B(_2557_));
 sg13g2_o21ai_1 _6539_ (.B1(net283),
    .Y(_2558_),
    .A1(_2163_),
    .A2(net1095));
 sg13g2_nand2_1 _6540_ (.Y(_0167_),
    .A(net1182),
    .B(_2558_));
 sg13g2_nor4_1 _6541_ (.A(_1806_),
    .B(_1823_),
    .C(_2171_),
    .D(net1095),
    .Y(_2559_));
 sg13g2_o21ai_1 _6542_ (.B1(net1182),
    .Y(_0168_),
    .A1(_2854_),
    .A2(_2559_));
 sg13g2_o21ai_1 _6543_ (.B1(net299),
    .Y(_2560_),
    .A1(_2180_),
    .A2(net1095));
 sg13g2_nand2_1 _6544_ (.Y(_0169_),
    .A(net1182),
    .B(_2560_));
 sg13g2_o21ai_1 _6545_ (.B1(net298),
    .Y(_2561_),
    .A1(_2166_),
    .A2(net1095));
 sg13g2_nand2_1 _6546_ (.Y(_0170_),
    .A(net1182),
    .B(_2561_));
 sg13g2_o21ai_1 _6547_ (.B1(net275),
    .Y(_2562_),
    .A1(_2178_),
    .A2(net1091));
 sg13g2_nand2_1 _6548_ (.Y(_0171_),
    .A(net1172),
    .B(_2562_));
 sg13g2_o21ai_1 _6549_ (.B1(net256),
    .Y(_2563_),
    .A1(_2167_),
    .A2(net1091));
 sg13g2_nand2_1 _6550_ (.Y(_0172_),
    .A(net1172),
    .B(_2563_));
 sg13g2_o21ai_1 _6551_ (.B1(net270),
    .Y(_2564_),
    .A1(_2169_),
    .A2(net1093));
 sg13g2_nand2_1 _6552_ (.Y(_0173_),
    .A(net1180),
    .B(_2564_));
 sg13g2_o21ai_1 _6553_ (.B1(net318),
    .Y(_2565_),
    .A1(_2164_),
    .A2(net1093));
 sg13g2_nand2_1 _6554_ (.Y(_0174_),
    .A(net1180),
    .B(_2565_));
 sg13g2_o21ai_1 _6555_ (.B1(net238),
    .Y(_2566_),
    .A1(_2162_),
    .A2(net1092));
 sg13g2_nand2_1 _6556_ (.Y(_0175_),
    .A(net1172),
    .B(_2566_));
 sg13g2_nor4_1 _6557_ (.A(_1806_),
    .B(_1823_),
    .C(_2173_),
    .D(net1095),
    .Y(_2567_));
 sg13g2_o21ai_1 _6558_ (.B1(net1180),
    .Y(_0176_),
    .A1(_2853_),
    .A2(_2567_));
 sg13g2_nor4_1 _6559_ (.A(_2134_),
    .B(_2147_),
    .C(_2175_),
    .D(net1093),
    .Y(_2568_));
 sg13g2_o21ai_1 _6560_ (.B1(net1180),
    .Y(_0177_),
    .A1(_2852_),
    .A2(_2568_));
 sg13g2_o21ai_1 _6561_ (.B1(net307),
    .Y(_2569_),
    .A1(_2165_),
    .A2(net1091));
 sg13g2_nand2_1 _6562_ (.Y(_0178_),
    .A(net1173),
    .B(_2569_));
 sg13g2_o21ai_1 _6563_ (.B1(net310),
    .Y(_2570_),
    .A1(_2228_),
    .A2(net1091));
 sg13g2_nand2_1 _6564_ (.Y(_0179_),
    .A(net1172),
    .B(_2570_));
 sg13g2_o21ai_1 _6565_ (.B1(net242),
    .Y(_2571_),
    .A1(_2212_),
    .A2(net1092));
 sg13g2_nand2_1 _6566_ (.Y(_0180_),
    .A(net1172),
    .B(_2571_));
 sg13g2_o21ai_1 _6567_ (.B1(net244),
    .Y(_2572_),
    .A1(_2217_),
    .A2(net1093));
 sg13g2_nand2_1 _6568_ (.Y(_0181_),
    .A(net1180),
    .B(_2572_));
 sg13g2_o21ai_1 _6569_ (.B1(net271),
    .Y(_2573_),
    .A1(_2215_),
    .A2(net1093));
 sg13g2_nand2_1 _6570_ (.Y(_0182_),
    .A(net1181),
    .B(_2573_));
 sg13g2_o21ai_1 _6571_ (.B1(net269),
    .Y(_2574_),
    .A1(_2216_),
    .A2(net1092));
 sg13g2_nand2_1 _6572_ (.Y(_0183_),
    .A(net1181),
    .B(_2574_));
 sg13g2_o21ai_1 _6573_ (.B1(net265),
    .Y(_2575_),
    .A1(_2224_),
    .A2(net1094));
 sg13g2_nand2_1 _6574_ (.Y(_0184_),
    .A(net1181),
    .B(_2575_));
 sg13g2_o21ai_1 _6575_ (.B1(net291),
    .Y(_2576_),
    .A1(_2227_),
    .A2(net1093));
 sg13g2_nand2_1 _6576_ (.Y(_0185_),
    .A(net1180),
    .B(_2576_));
 sg13g2_o21ai_1 _6577_ (.B1(net289),
    .Y(_2577_),
    .A1(_2214_),
    .A2(net1091));
 sg13g2_nand2_1 _6578_ (.Y(_0186_),
    .A(net1172),
    .B(_2577_));
 sg13g2_o21ai_1 _6579_ (.B1(net276),
    .Y(_2578_),
    .A1(_2225_),
    .A2(net1091));
 sg13g2_nand2_1 _6580_ (.Y(_0187_),
    .A(net1172),
    .B(_2578_));
 sg13g2_o21ai_1 _6581_ (.B1(net300),
    .Y(_2579_),
    .A1(_2213_),
    .A2(net1091));
 sg13g2_nand2_1 _6582_ (.Y(_0188_),
    .A(net1172),
    .B(_2579_));
 sg13g2_o21ai_1 _6583_ (.B1(net286),
    .Y(_2580_),
    .A1(_2218_),
    .A2(net1094));
 sg13g2_nand2_1 _6584_ (.Y(_0189_),
    .A(net1181),
    .B(_2580_));
 sg13g2_o21ai_1 _6585_ (.B1(net278),
    .Y(_2581_),
    .A1(_2206_),
    .A2(net1093));
 sg13g2_nand2_1 _6586_ (.Y(_0190_),
    .A(net1180),
    .B(_2581_));
 sg13g2_o21ai_1 _6587_ (.B1(net301),
    .Y(_2582_),
    .A1(_2207_),
    .A2(net1091));
 sg13g2_nand2_1 _6588_ (.Y(_0191_),
    .A(net1181),
    .B(_2582_));
 sg13g2_o21ai_1 _6589_ (.B1(net303),
    .Y(_2583_),
    .A1(_2221_),
    .A2(net1093));
 sg13g2_nand2_1 _6590_ (.Y(_0192_),
    .A(net1181),
    .B(_2583_));
 sg13g2_o21ai_1 _6591_ (.B1(net287),
    .Y(_2584_),
    .A1(_2203_),
    .A2(net1097));
 sg13g2_nand2_1 _6592_ (.Y(_0193_),
    .A(net1184),
    .B(_2584_));
 sg13g2_o21ai_1 _6593_ (.B1(net309),
    .Y(_2585_),
    .A1(_2204_),
    .A2(net1097));
 sg13g2_nand2_1 _6594_ (.Y(_0194_),
    .A(net1184),
    .B(_2585_));
 sg13g2_and2_1 _6595_ (.A(net4),
    .B(net1181),
    .X(_0195_));
 sg13g2_nand2_1 _6596_ (.Y(_2586_),
    .A(net1320),
    .B(_2344_));
 sg13g2_or2_1 _6597_ (.X(_2587_),
    .B(_2259_),
    .A(_2885_));
 sg13g2_xor2_1 _6598_ (.B(_2586_),
    .A(\barrier_health[0][0] ),
    .X(_2588_));
 sg13g2_nand3_1 _6599_ (.B(_2587_),
    .C(_2588_),
    .A(net1150),
    .Y(_2589_));
 sg13g2_nor3_1 _6600_ (.A(net263),
    .B(_1767_),
    .C(_2259_),
    .Y(_2590_));
 sg13g2_o21ai_1 _6601_ (.B1(_2589_),
    .Y(_2591_),
    .A1(\barrier_health[0][0] ),
    .A2(net1150));
 sg13g2_o21ai_1 _6602_ (.B1(net1174),
    .Y(_0196_),
    .A1(_2590_),
    .A2(_2591_));
 sg13g2_a21o_1 _6603_ (.A2(_2587_),
    .A1(_2586_),
    .B1(net1144),
    .X(_2592_));
 sg13g2_o21ai_1 _6604_ (.B1(net315),
    .Y(_2593_),
    .A1(\barrier_health[0][0] ),
    .A2(_2592_));
 sg13g2_or3_1 _6605_ (.A(net315),
    .B(\barrier_health[0][0] ),
    .C(_2592_),
    .X(_2594_));
 sg13g2_a21oi_1 _6606_ (.A1(net316),
    .A2(_2594_),
    .Y(_0197_),
    .B1(net1167));
 sg13g2_a21o_1 _6607_ (.A2(_2594_),
    .A1(net251),
    .B1(net1167),
    .X(_0198_));
 sg13g2_nand2_1 _6608_ (.Y(_2595_),
    .A(net1320),
    .B(_2351_));
 sg13g2_nor2_1 _6609_ (.A(net1145),
    .B(_2595_),
    .Y(_2596_));
 sg13g2_nor2b_2 _6610_ (.A(_1767_),
    .B_N(_2250_),
    .Y(_2597_));
 sg13g2_xnor2_1 _6611_ (.Y(_2598_),
    .A(\barrier_health[1][0] ),
    .B(_2596_));
 sg13g2_a21oi_1 _6612_ (.A1(net221),
    .A2(_2597_),
    .Y(_2599_),
    .B1(net1167));
 sg13g2_o21ai_1 _6613_ (.B1(_2599_),
    .Y(_0199_),
    .A1(_2597_),
    .A2(_2598_));
 sg13g2_xor2_1 _6614_ (.B(\barrier_health[1][0] ),
    .A(net353),
    .X(_2600_));
 sg13g2_or2_1 _6615_ (.X(_2601_),
    .B(_2600_),
    .A(_2595_));
 sg13g2_a221oi_1 _6616_ (.B2(net353),
    .C1(net1144),
    .B1(_2595_),
    .A1(pb_active),
    .Y(_2602_),
    .A2(_2250_));
 sg13g2_o21ai_1 _6617_ (.B1(net1174),
    .Y(_2603_),
    .A1(net353),
    .A2(net1150));
 sg13g2_a221oi_1 _6618_ (.B2(_2602_),
    .C1(_2603_),
    .B1(_2601_),
    .A1(_2597_),
    .Y(_0200_),
    .A2(_2600_));
 sg13g2_or2_1 _6619_ (.X(_2604_),
    .B(_2597_),
    .A(_2596_));
 sg13g2_or2_1 _6620_ (.X(_2605_),
    .B(_2604_),
    .A(net392));
 sg13g2_o21ai_1 _6621_ (.B1(net392),
    .Y(_2606_),
    .A1(\barrier_health[1][1] ),
    .A2(\barrier_health[1][0] ));
 sg13g2_nand3b_1 _6622_ (.B(_2604_),
    .C(_2606_),
    .Y(_2607_),
    .A_N(_0384_));
 sg13g2_a21o_1 _6623_ (.A2(_2607_),
    .A1(_2605_),
    .B1(net1168),
    .X(_0201_));
 sg13g2_nand2_1 _6624_ (.Y(_2608_),
    .A(net1327),
    .B(_2268_));
 sg13g2_nand2_1 _6625_ (.Y(_2609_),
    .A(net1154),
    .B(_2608_));
 sg13g2_nand2_2 _6626_ (.Y(_2610_),
    .A(net1320),
    .B(_2360_));
 sg13g2_xnor2_1 _6627_ (.Y(_2611_),
    .A(\barrier_health[2][0] ),
    .B(_2610_));
 sg13g2_nor2_1 _6628_ (.A(_2609_),
    .B(_2611_),
    .Y(_2612_));
 sg13g2_nand2b_1 _6629_ (.Y(_2613_),
    .B(net1145),
    .A_N(\barrier_health[2][0] ));
 sg13g2_nand3_1 _6630_ (.B(net1150),
    .C(_2268_),
    .A(net1327),
    .Y(_2614_));
 sg13g2_o21ai_1 _6631_ (.B1(_2613_),
    .Y(_2615_),
    .A1(net240),
    .A2(_2614_));
 sg13g2_o21ai_1 _6632_ (.B1(net1175),
    .Y(_0202_),
    .A1(_2612_),
    .A2(net241));
 sg13g2_xnor2_1 _6633_ (.Y(_2616_),
    .A(net361),
    .B(\barrier_health[2][0] ));
 sg13g2_mux2_1 _6634_ (.A0(_2616_),
    .A1(net361),
    .S(_2610_),
    .X(_2617_));
 sg13g2_nor2_1 _6635_ (.A(_2609_),
    .B(_2617_),
    .Y(_2618_));
 sg13g2_o21ai_1 _6636_ (.B1(net1176),
    .Y(_2619_),
    .A1(net361),
    .A2(net1154));
 sg13g2_nor2_1 _6637_ (.A(_2614_),
    .B(_2616_),
    .Y(_2620_));
 sg13g2_nor3_1 _6638_ (.A(_2618_),
    .B(_2619_),
    .C(_2620_),
    .Y(_0203_));
 sg13g2_a21oi_1 _6639_ (.A1(_2608_),
    .A2(_2610_),
    .Y(_2621_),
    .B1(net1145));
 sg13g2_o21ai_1 _6640_ (.B1(\barrier_health[2][2] ),
    .Y(_2622_),
    .A1(\barrier_health[2][1] ),
    .A2(\barrier_health[2][0] ));
 sg13g2_nand2_1 _6641_ (.Y(_2623_),
    .A(_0293_),
    .B(_2622_));
 sg13g2_mux2_1 _6642_ (.A0(net363),
    .A1(_2623_),
    .S(_2621_),
    .X(_2624_));
 sg13g2_nand2b_1 _6643_ (.Y(_0204_),
    .B(net1176),
    .A_N(_2624_));
 sg13g2_nand2_2 _6644_ (.Y(_2625_),
    .A(net1320),
    .B(_2328_));
 sg13g2_nor2_1 _6645_ (.A(net1145),
    .B(_2625_),
    .Y(_2626_));
 sg13g2_xnor2_1 _6646_ (.Y(_2627_),
    .A(\barrier_health[3][0] ),
    .B(_2626_));
 sg13g2_a21oi_1 _6647_ (.A1(net225),
    .A2(_2280_),
    .Y(_2628_),
    .B1(net1167));
 sg13g2_o21ai_1 _6648_ (.B1(_2628_),
    .Y(_0205_),
    .A1(_2280_),
    .A2(_2627_));
 sg13g2_o21ai_1 _6649_ (.B1(net1174),
    .Y(_2629_),
    .A1(net348),
    .A2(net1151));
 sg13g2_xor2_1 _6650_ (.B(\barrier_health[3][0] ),
    .A(net348),
    .X(_2630_));
 sg13g2_nand2_1 _6651_ (.Y(_2631_),
    .A(net1150),
    .B(_2279_));
 sg13g2_or2_1 _6652_ (.X(_2632_),
    .B(_2630_),
    .A(_2625_));
 sg13g2_a21oi_1 _6653_ (.A1(net348),
    .A2(_2625_),
    .Y(_2633_),
    .B1(_2631_));
 sg13g2_a221oi_1 _6654_ (.B2(_2633_),
    .C1(_2629_),
    .B1(_2632_),
    .A1(_2280_),
    .Y(_0206_),
    .A2(_2630_));
 sg13g2_o21ai_1 _6655_ (.B1(\barrier_health[3][2] ),
    .Y(_2634_),
    .A1(\barrier_health[3][1] ),
    .A2(\barrier_health[3][0] ));
 sg13g2_nor2b_1 _6656_ (.A(_0372_),
    .B_N(_2634_),
    .Y(_2635_));
 sg13g2_a21oi_1 _6657_ (.A1(net364),
    .A2(_2625_),
    .Y(_2636_),
    .B1(_2631_));
 sg13g2_o21ai_1 _6658_ (.B1(_2636_),
    .Y(_2637_),
    .A1(_2625_),
    .A2(_2635_));
 sg13g2_and2_1 _6659_ (.A(_2280_),
    .B(_2635_),
    .X(_2638_));
 sg13g2_o21ai_1 _6660_ (.B1(_2637_),
    .Y(_2639_),
    .A1(net364),
    .A2(net1150));
 sg13g2_o21ai_1 _6661_ (.B1(net1174),
    .Y(_0207_),
    .A1(_2638_),
    .A2(_2639_));
 sg13g2_nor2_1 _6662_ (.A(net1212),
    .B(net1413),
    .Y(_0263_));
 sg13g2_nor2_1 _6663_ (.A(net1212),
    .B(net1165),
    .Y(_0208_));
 sg13g2_nor2_1 _6664_ (.A(net1214),
    .B(net1412),
    .Y(_0264_));
 sg13g2_nor2_1 _6665_ (.A(net1214),
    .B(net1165),
    .Y(_0209_));
 sg13g2_nor2_1 _6666_ (.A(net1217),
    .B(net1412),
    .Y(_0265_));
 sg13g2_nor2_1 _6667_ (.A(net1217),
    .B(net1164),
    .Y(_0210_));
 sg13g2_nor2_1 _6668_ (.A(net1221),
    .B(net1412),
    .Y(_0266_));
 sg13g2_nor2_1 _6669_ (.A(net1221),
    .B(net1164),
    .Y(_0211_));
 sg13g2_nor2_1 _6670_ (.A(_2846_),
    .B(net1412),
    .Y(_0267_));
 sg13g2_nor2_1 _6671_ (.A(net1222),
    .B(net1164),
    .Y(_0212_));
 sg13g2_nor2_1 _6672_ (.A(_2845_),
    .B(net1412),
    .Y(_0268_));
 sg13g2_nor2_1 _6673_ (.A(net1223),
    .B(net1164),
    .Y(_0213_));
 sg13g2_nor2_1 _6674_ (.A(_2844_),
    .B(net1412),
    .Y(_0269_));
 sg13g2_nor2_1 _6675_ (.A(_2844_),
    .B(net1164),
    .Y(_0214_));
 sg13g2_nor2_1 _6676_ (.A(net1224),
    .B(net1412),
    .Y(_0270_));
 sg13g2_nor2_1 _6677_ (.A(net1224),
    .B(net1164),
    .Y(_0215_));
 sg13g2_nor2_1 _6678_ (.A(_2842_),
    .B(net1413),
    .Y(_0271_));
 sg13g2_nor2_1 _6679_ (.A(_2842_),
    .B(net1164),
    .Y(_0216_));
 sg13g2_nor2_1 _6680_ (.A(net1225),
    .B(net1412),
    .Y(_0272_));
 sg13g2_nor2_1 _6681_ (.A(net1225),
    .B(net1164),
    .Y(_0217_));
 sg13g2_and4_1 _6682_ (.A(_2824_),
    .B(net1242),
    .C(net1246),
    .D(_0746_),
    .X(_2640_));
 sg13g2_nor4_1 _6683_ (.A(_0628_),
    .B(_1940_),
    .C(_1952_),
    .D(_2640_),
    .Y(_2641_));
 sg13g2_nor3_2 _6684_ (.A(net1231),
    .B(_1962_),
    .C(_2641_),
    .Y(_2642_));
 sg13g2_o21ai_1 _6685_ (.B1(net1302),
    .Y(_2643_),
    .A1(net1147),
    .A2(_2642_));
 sg13g2_nor2b_1 _6686_ (.A(_0747_),
    .B_N(net1243),
    .Y(_2644_));
 sg13g2_o21ai_1 _6687_ (.B1(net1238),
    .Y(_2645_),
    .A1(net1240),
    .A2(_2644_));
 sg13g2_nor2b_1 _6688_ (.A(net1231),
    .B_N(net1244),
    .Y(_2646_));
 sg13g2_a21oi_1 _6689_ (.A1(net1238),
    .A2(_2646_),
    .Y(_2647_),
    .B1(_0078_));
 sg13g2_nor2_1 _6690_ (.A(_0599_),
    .B(_2647_),
    .Y(_2648_));
 sg13g2_nand4_1 _6691_ (.B(net1152),
    .C(_2645_),
    .A(net229),
    .Y(_2649_),
    .D(_2648_));
 sg13g2_nand3_1 _6692_ (.B(_2643_),
    .C(_2649_),
    .A(net1),
    .Y(_0219_));
 sg13g2_or2_1 _6693_ (.X(_2650_),
    .B(_3094_),
    .A(_3089_));
 sg13g2_a21oi_1 _6694_ (.A1(_3228_),
    .A2(_2650_),
    .Y(_2651_),
    .B1(net1352));
 sg13g2_o21ai_1 _6695_ (.B1(net1353),
    .Y(_2652_),
    .A1(net1358),
    .A2(_0367_));
 sg13g2_nor3_2 _6696_ (.A(net1414),
    .B(_2651_),
    .C(_2652_),
    .Y(_0221_));
 sg13g2_nand2_1 _6697_ (.Y(_2653_),
    .A(net1299),
    .B(_3080_));
 sg13g2_nand2_1 _6698_ (.Y(_2654_),
    .A(net1417),
    .B(_3078_));
 sg13g2_nor4_1 _6699_ (.A(net1225),
    .B(net1268),
    .C(net1281),
    .D(_1235_),
    .Y(_2655_));
 sg13g2_a21oi_2 _6700_ (.B1(_2654_),
    .Y(_2656_),
    .A2(_2655_),
    .A1(_1117_));
 sg13g2_nor2_1 _6701_ (.A(net1299),
    .B(net1083),
    .Y(_2657_));
 sg13g2_a21oi_1 _6702_ (.A1(net1299),
    .A2(_3080_),
    .Y(_0222_),
    .B1(_2657_));
 sg13g2_nand2_1 _6703_ (.Y(_2658_),
    .A(net1416),
    .B(net1187));
 sg13g2_a22oi_1 _6704_ (.Y(_0223_),
    .B1(_2658_),
    .B2(_3080_),
    .A2(_2653_),
    .A1(net1214));
 sg13g2_a22oi_1 _6705_ (.Y(_2659_),
    .B1(_0588_),
    .B2(net1083),
    .A2(net1088),
    .A1(net1294));
 sg13g2_inv_1 _6706_ (.Y(_0224_),
    .A(_2659_));
 sg13g2_xnor2_1 _6707_ (.Y(_2660_),
    .A(net1284),
    .B(_1115_));
 sg13g2_a22oi_1 _6708_ (.Y(_2661_),
    .B1(net1083),
    .B2(_2660_),
    .A2(net1088),
    .A1(net1289));
 sg13g2_inv_1 _6709_ (.Y(_0225_),
    .A(net370));
 sg13g2_nor2_1 _6710_ (.A(net1187),
    .B(_0534_),
    .Y(_2662_));
 sg13g2_nor3_1 _6711_ (.A(net1278),
    .B(net1187),
    .C(_0534_),
    .Y(_2663_));
 sg13g2_xnor2_1 _6712_ (.Y(_2664_),
    .A(net1278),
    .B(_2662_));
 sg13g2_a22oi_1 _6713_ (.Y(_2665_),
    .B1(net1083),
    .B2(_2664_),
    .A2(net1088),
    .A1(net1280));
 sg13g2_inv_1 _6714_ (.Y(_0226_),
    .A(_2665_));
 sg13g2_xnor2_1 _6715_ (.Y(_2666_),
    .A(net414),
    .B(_2663_));
 sg13g2_a22oi_1 _6716_ (.Y(_2667_),
    .B1(net1083),
    .B2(_2666_),
    .A2(net1088),
    .A1(net1276));
 sg13g2_inv_1 _6717_ (.Y(_0227_),
    .A(_2667_));
 sg13g2_nand3_1 _6718_ (.B(net1280),
    .C(_2662_),
    .A(net1276),
    .Y(_2668_));
 sg13g2_nor2_1 _6719_ (.A(_0014_),
    .B(_2668_),
    .Y(_2669_));
 sg13g2_xnor2_1 _6720_ (.Y(_2670_),
    .A(_2907_),
    .B(_2668_));
 sg13g2_a22oi_1 _6721_ (.Y(_2671_),
    .B1(net1083),
    .B2(_2670_),
    .A2(net1088),
    .A1(net1273));
 sg13g2_inv_1 _6722_ (.Y(_0228_),
    .A(_2671_));
 sg13g2_xnor2_1 _6723_ (.Y(_2672_),
    .A(net405),
    .B(_2669_));
 sg13g2_a22oi_1 _6724_ (.Y(_2673_),
    .B1(_2656_),
    .B2(_2672_),
    .A2(net1088),
    .A1(net1271));
 sg13g2_inv_1 _6725_ (.Y(_0229_),
    .A(_2673_));
 sg13g2_nor3_1 _6726_ (.A(net1224),
    .B(_2844_),
    .C(_2668_),
    .Y(_2674_));
 sg13g2_nand2b_1 _6727_ (.Y(_2675_),
    .B(_2674_),
    .A_N(net1266));
 sg13g2_xnor2_1 _6728_ (.Y(_2676_),
    .A(net1266),
    .B(_2674_));
 sg13g2_a22oi_1 _6729_ (.Y(_2677_),
    .B1(net1083),
    .B2(_2676_),
    .A2(net1088),
    .A1(net1269));
 sg13g2_inv_1 _6730_ (.Y(_0230_),
    .A(_2677_));
 sg13g2_o21ai_1 _6731_ (.B1(net1083),
    .Y(_2678_),
    .A1(net341),
    .A2(_2675_));
 sg13g2_a21o_1 _6732_ (.A2(_2675_),
    .A1(net341),
    .B1(_2678_),
    .X(_2679_));
 sg13g2_o21ai_1 _6733_ (.B1(_2679_),
    .Y(_0231_),
    .A1(net1225),
    .A2(_3080_));
 sg13g2_nand4_1 _6734_ (.B(_3100_),
    .C(_3200_),
    .A(net1295),
    .Y(_2680_),
    .D(_1384_));
 sg13g2_nor4_1 _6735_ (.A(net1264),
    .B(_2842_),
    .C(_2654_),
    .D(_2680_),
    .Y(_2681_));
 sg13g2_a21o_1 _6736_ (.A2(net1089),
    .A1(net235),
    .B1(_2681_),
    .X(_0232_));
 sg13g2_o21ai_1 _6737_ (.B1(_3005_),
    .Y(_2682_),
    .A1(net1261),
    .A2(net1263));
 sg13g2_nor2_1 _6738_ (.A(\myShooter.shooter_left_x[9] ),
    .B(_2897_),
    .Y(_2683_));
 sg13g2_a22oi_1 _6739_ (.Y(_2684_),
    .B1(_2682_),
    .B2(_2683_),
    .A2(\movement_dir[2] ),
    .A1(_2897_));
 sg13g2_nor4_1 _6740_ (.A(\prev_vpos_shooter[7] ),
    .B(\prev_vpos_shooter[6] ),
    .C(\prev_vpos_shooter[9] ),
    .D(\prev_vpos_shooter[8] ),
    .Y(_2685_));
 sg13g2_nor2_1 _6741_ (.A(\prev_vpos_shooter[1] ),
    .B(\prev_vpos_shooter[0] ),
    .Y(_2686_));
 sg13g2_nor4_1 _6742_ (.A(\prev_vpos_shooter[3] ),
    .B(\prev_vpos_shooter[2] ),
    .C(\prev_vpos_shooter[5] ),
    .D(\prev_vpos_shooter[4] ),
    .Y(_2687_));
 sg13g2_nand3_1 _6743_ (.B(_2686_),
    .C(_2687_),
    .A(_2685_),
    .Y(_2688_));
 sg13g2_nor4_1 _6744_ (.A(net1256),
    .B(net1257),
    .C(net1258),
    .D(\myShooter.shooter_left_x[5] ),
    .Y(_2689_));
 sg13g2_o21ai_1 _6745_ (.B1(net1259),
    .Y(_2690_),
    .A1(net1261),
    .A2(net1263));
 sg13g2_nand4_1 _6746_ (.B(\movement_dir[2] ),
    .C(_2689_),
    .A(_2835_),
    .Y(_2691_),
    .D(_2690_));
 sg13g2_nand3_1 _6747_ (.B(_2688_),
    .C(_2691_),
    .A(_3051_),
    .Y(_2692_));
 sg13g2_or2_1 _6748_ (.X(_2693_),
    .B(_2692_),
    .A(_2684_));
 sg13g2_a21oi_1 _6749_ (.A1(net237),
    .A2(net1082),
    .Y(_2694_),
    .B1(net1168));
 sg13g2_o21ai_1 _6750_ (.B1(_2694_),
    .Y(_0233_),
    .A1(_2840_),
    .A2(net1082));
 sg13g2_xnor2_1 _6751_ (.Y(_2695_),
    .A(net231),
    .B(net1230));
 sg13g2_o21ai_1 _6752_ (.B1(net1263),
    .Y(_2696_),
    .A1(net1082),
    .A2(_2695_));
 sg13g2_or3_1 _6753_ (.A(net1263),
    .B(net1082),
    .C(_2695_),
    .X(_2697_));
 sg13g2_nand3_1 _6754_ (.B(_2696_),
    .C(_2697_),
    .A(net1176),
    .Y(_0234_));
 sg13g2_xor2_1 _6755_ (.B(net1230),
    .A(net1262),
    .X(_2698_));
 sg13g2_a21oi_1 _6756_ (.A1(net1230),
    .A2(_1744_),
    .Y(_2699_),
    .B1(_1743_));
 sg13g2_and2_1 _6757_ (.A(_2698_),
    .B(_2699_),
    .X(_2700_));
 sg13g2_xnor2_1 _6758_ (.Y(_2701_),
    .A(_2698_),
    .B(_2699_));
 sg13g2_a21oi_1 _6759_ (.A1(net1262),
    .A2(net1082),
    .Y(_2702_),
    .B1(net1168));
 sg13g2_o21ai_1 _6760_ (.B1(_2702_),
    .Y(_0235_),
    .A1(net1082),
    .A2(_2701_));
 sg13g2_xnor2_1 _6761_ (.Y(_2703_),
    .A(net1260),
    .B(net1230));
 sg13g2_a21oi_1 _6762_ (.A1(net1262),
    .A2(net1230),
    .Y(_2704_),
    .B1(_2700_));
 sg13g2_xor2_1 _6763_ (.B(_2704_),
    .A(_2703_),
    .X(_2705_));
 sg13g2_a21oi_1 _6764_ (.A1(net1260),
    .A2(net1082),
    .Y(_2706_),
    .B1(net1168));
 sg13g2_o21ai_1 _6765_ (.B1(_2706_),
    .Y(_0236_),
    .A1(net1082),
    .A2(_2705_));
 sg13g2_xor2_1 _6766_ (.B(net1229),
    .A(\myShooter.shooter_left_x[5] ),
    .X(_2707_));
 sg13g2_nand2_1 _6767_ (.Y(_2708_),
    .A(_2700_),
    .B(_2703_));
 sg13g2_o21ai_1 _6768_ (.B1(net1259),
    .Y(_2709_),
    .A1(net1261),
    .A2(_2897_));
 sg13g2_nand2_2 _6769_ (.Y(_2710_),
    .A(_2708_),
    .B(_2709_));
 sg13g2_nand2b_1 _6770_ (.Y(_2711_),
    .B(_2710_),
    .A_N(_2707_));
 sg13g2_xor2_1 _6771_ (.B(_2710_),
    .A(_2707_),
    .X(_2712_));
 sg13g2_o21ai_1 _6772_ (.B1(net1178),
    .Y(_2713_),
    .A1(net1081),
    .A2(_2712_));
 sg13g2_a21o_1 _6773_ (.A2(net1081),
    .A1(net396),
    .B1(_2713_),
    .X(_0237_));
 sg13g2_o21ai_1 _6774_ (.B1(_2711_),
    .Y(_2714_),
    .A1(_2838_),
    .A2(net1229));
 sg13g2_xnor2_1 _6775_ (.Y(_2715_),
    .A(net1258),
    .B(net1229));
 sg13g2_xnor2_1 _6776_ (.Y(_2716_),
    .A(_2714_),
    .B(_2715_));
 sg13g2_a21oi_1 _6777_ (.A1(net304),
    .A2(net1081),
    .Y(_2717_),
    .B1(net1167));
 sg13g2_o21ai_1 _6778_ (.B1(_2717_),
    .Y(_0238_),
    .A1(net1081),
    .A2(_2716_));
 sg13g2_xnor2_1 _6779_ (.Y(_2718_),
    .A(net1257),
    .B(net1229));
 sg13g2_a21oi_1 _6780_ (.A1(net1258),
    .A2(_2897_),
    .Y(_2719_),
    .B1(_2714_));
 sg13g2_a21oi_1 _6781_ (.A1(_2837_),
    .A2(net1229),
    .Y(_2720_),
    .B1(_2719_));
 sg13g2_xnor2_1 _6782_ (.Y(_2721_),
    .A(_2718_),
    .B(_2720_));
 sg13g2_a21oi_1 _6783_ (.A1(net1257),
    .A2(net1081),
    .Y(_2722_),
    .B1(net1167));
 sg13g2_o21ai_1 _6784_ (.B1(_2722_),
    .Y(_0239_),
    .A1(net1081),
    .A2(_2721_));
 sg13g2_nand3_1 _6785_ (.B(_2897_),
    .C(_2719_),
    .A(_2836_),
    .Y(_2723_));
 sg13g2_nand3_1 _6786_ (.B(net1229),
    .C(_2720_),
    .A(net1257),
    .Y(_2724_));
 sg13g2_a21oi_1 _6787_ (.A1(_2723_),
    .A2(_2724_),
    .Y(_2725_),
    .B1(net1081));
 sg13g2_o21ai_1 _6788_ (.B1(net1175),
    .Y(_2726_),
    .A1(net1256),
    .A2(_2725_));
 sg13g2_a21oi_1 _6789_ (.A1(net1256),
    .A2(_2725_),
    .Y(_0240_),
    .B1(_2726_));
 sg13g2_nor2_1 _6790_ (.A(net1229),
    .B(_2689_),
    .Y(_2727_));
 sg13g2_nor3_1 _6791_ (.A(net1081),
    .B(_2710_),
    .C(_2727_),
    .Y(_2728_));
 sg13g2_nor3_1 _6792_ (.A(_2835_),
    .B(net1167),
    .C(_2728_),
    .Y(_0241_));
 sg13g2_a21oi_2 _6793_ (.B1(net1144),
    .Y(_2729_),
    .A2(_2363_),
    .A1(_2332_));
 sg13g2_a21o_2 _6794_ (.A2(_2363_),
    .A1(_2332_),
    .B1(net1144),
    .X(_2730_));
 sg13g2_nand2b_1 _6795_ (.Y(_2731_),
    .B(\selectedRowRand[0] ),
    .A_N(\selectedRowRand[1] ));
 sg13g2_nor3_1 _6796_ (.A(net1318),
    .B(_2917_),
    .C(_2731_),
    .Y(_2732_));
 sg13g2_nor2_1 _6797_ (.A(\selectedRowRand[2] ),
    .B(net1318),
    .Y(_2733_));
 sg13g2_nand2_1 _6798_ (.Y(_2734_),
    .A(net245),
    .B(_2733_));
 sg13g2_inv_1 _6799_ (.Y(_2735_),
    .A(_2734_));
 sg13g2_a21oi_1 _6800_ (.A1(\selectedRowRand[0] ),
    .A2(_2735_),
    .Y(_2736_),
    .B1(_2732_));
 sg13g2_nor2b_1 _6801_ (.A(net325),
    .B_N(net1318),
    .Y(_2737_));
 sg13g2_o21ai_1 _6802_ (.B1(_2736_),
    .Y(_2738_),
    .A1(_0063_),
    .A2(_2734_));
 sg13g2_o21ai_1 _6803_ (.B1(net1090),
    .Y(_2739_),
    .A1(_2737_),
    .A2(_2738_));
 sg13g2_o21ai_1 _6804_ (.B1(net326),
    .Y(_2740_),
    .A1(\abullet_y[1] ),
    .A2(net1090));
 sg13g2_nor2_1 _6805_ (.A(net1166),
    .B(net327),
    .Y(_0242_));
 sg13g2_a21o_1 _6806_ (.A2(_3126_),
    .A1(net1318),
    .B1(_2735_),
    .X(_2741_));
 sg13g2_o21ai_1 _6807_ (.B1(net1170),
    .Y(_2742_),
    .A1(net1255),
    .A2(net1090));
 sg13g2_a21oi_1 _6808_ (.A1(net1090),
    .A2(_2741_),
    .Y(_0243_),
    .B1(_2742_));
 sg13g2_nand2_1 _6809_ (.Y(_2743_),
    .A(net338),
    .B(_3125_));
 sg13g2_xnor2_1 _6810_ (.Y(_2744_),
    .A(net338),
    .B(_3125_));
 sg13g2_a21oi_1 _6811_ (.A1(_2731_),
    .A2(_2733_),
    .Y(_2745_),
    .B1(_2732_));
 sg13g2_nand2_1 _6812_ (.Y(_2746_),
    .A(net1090),
    .B(_2745_));
 sg13g2_a21oi_1 _6813_ (.A1(net1318),
    .A2(_2744_),
    .Y(_2747_),
    .B1(_2746_));
 sg13g2_o21ai_1 _6814_ (.B1(net1170),
    .Y(_2748_),
    .A1(\abullet_y[3] ),
    .A2(net1090));
 sg13g2_nor2_1 _6815_ (.A(_2747_),
    .B(_2748_),
    .Y(_0244_));
 sg13g2_a21oi_1 _6816_ (.A1(net372),
    .A2(_2743_),
    .Y(_2749_),
    .B1(_0030_));
 sg13g2_o21ai_1 _6817_ (.B1(_2749_),
    .Y(_2750_),
    .A1(net372),
    .A2(_2743_));
 sg13g2_o21ai_1 _6818_ (.B1(net1170),
    .Y(_2751_),
    .A1(_2730_),
    .A2(net373));
 sg13g2_a21oi_1 _6819_ (.A1(_2832_),
    .A2(_2730_),
    .Y(_0245_),
    .B1(_2751_));
 sg13g2_o21ai_1 _6820_ (.B1(_2736_),
    .Y(_2752_),
    .A1(_2832_),
    .A2(_2329_));
 sg13g2_a21oi_1 _6821_ (.A1(_2729_),
    .A2(_2752_),
    .Y(_2753_),
    .B1(net331));
 sg13g2_or2_1 _6822_ (.X(_2754_),
    .B(_2329_),
    .A(_3008_));
 sg13g2_nand2_1 _6823_ (.Y(_2755_),
    .A(net1318),
    .B(_2754_));
 sg13g2_and3_1 _6824_ (.X(_2756_),
    .A(_2729_),
    .B(_2736_),
    .C(_2755_));
 sg13g2_nor3_1 _6825_ (.A(net1166),
    .B(_2753_),
    .C(_2756_),
    .Y(_0246_));
 sg13g2_a21oi_1 _6826_ (.A1(_2734_),
    .A2(_2754_),
    .Y(_2757_),
    .B1(_2730_));
 sg13g2_or2_2 _6827_ (.X(_2758_),
    .B(_2754_),
    .A(_2830_));
 sg13g2_a21oi_1 _6828_ (.A1(net1318),
    .A2(_2758_),
    .Y(_2759_),
    .B1(_2735_));
 sg13g2_o21ai_1 _6829_ (.B1(net1171),
    .Y(_2760_),
    .A1(net1254),
    .A2(_2757_));
 sg13g2_a21oi_1 _6830_ (.A1(_2729_),
    .A2(_2759_),
    .Y(_0247_),
    .B1(_2760_));
 sg13g2_o21ai_1 _6831_ (.B1(net1319),
    .Y(_2761_),
    .A1(_2829_),
    .A2(_2758_));
 sg13g2_nor2b_1 _6832_ (.A(_2746_),
    .B_N(_2761_),
    .Y(_2762_));
 sg13g2_a21oi_1 _6833_ (.A1(_2745_),
    .A2(_2758_),
    .Y(_2763_),
    .B1(_2730_));
 sg13g2_o21ai_1 _6834_ (.B1(net1171),
    .Y(_2764_),
    .A1(net340),
    .A2(_2763_));
 sg13g2_nor2_1 _6835_ (.A(_2762_),
    .B(_2764_),
    .Y(_0248_));
 sg13g2_o21ai_1 _6836_ (.B1(net346),
    .Y(_2765_),
    .A1(_0050_),
    .A2(_2758_));
 sg13g2_nor3_1 _6837_ (.A(\abullet_y[8] ),
    .B(_0050_),
    .C(_2758_),
    .Y(_2766_));
 sg13g2_nor2b_1 _6838_ (.A(_2766_),
    .B_N(net1319),
    .Y(_2767_));
 sg13g2_a21oi_1 _6839_ (.A1(_2765_),
    .A2(_2767_),
    .Y(_2768_),
    .B1(_2746_));
 sg13g2_a21oi_1 _6840_ (.A1(net346),
    .A2(_2730_),
    .Y(_2769_),
    .B1(_2768_));
 sg13g2_nor2_1 _6841_ (.A(net1166),
    .B(net347),
    .Y(_0249_));
 sg13g2_or3_1 _6842_ (.A(net333),
    .B(_3016_),
    .C(_2758_),
    .X(_2770_));
 sg13g2_o21ai_1 _6843_ (.B1(net333),
    .Y(_2771_),
    .A1(_3016_),
    .A2(_2758_));
 sg13g2_nand3_1 _6844_ (.B(_2770_),
    .C(_2771_),
    .A(net1319),
    .Y(_2772_));
 sg13g2_o21ai_1 _6845_ (.B1(net1170),
    .Y(_2773_),
    .A1(\abullet_y[9] ),
    .A2(net1090));
 sg13g2_a21oi_1 _6846_ (.A1(net1090),
    .A2(_2772_),
    .Y(_0250_),
    .B1(_2773_));
 sg13g2_nor2_1 _6847_ (.A(_3064_),
    .B(_0002_),
    .Y(_0251_));
 sg13g2_nand2_1 _6848_ (.Y(_0252_),
    .A(_0001_),
    .B(_0002_));
 sg13g2_o21ai_1 _6849_ (.B1(net1),
    .Y(_2774_),
    .A1(net281),
    .A2(net1147));
 sg13g2_a21oi_1 _6850_ (.A1(_2827_),
    .A2(net1147),
    .Y(_0253_),
    .B1(_2774_));
 sg13g2_xor2_1 _6851_ (.B(net281),
    .A(net1250),
    .X(_2775_));
 sg13g2_xnor2_1 _6852_ (.Y(_2776_),
    .A(_2851_),
    .B(_2775_));
 sg13g2_a21oi_1 _6853_ (.A1(net1152),
    .A2(_2776_),
    .Y(_2777_),
    .B1(net1415));
 sg13g2_o21ai_1 _6854_ (.B1(_2777_),
    .Y(_0254_),
    .A1(_2826_),
    .A2(net1153));
 sg13g2_xnor2_1 _6855_ (.Y(_2778_),
    .A(net1248),
    .B(net1302));
 sg13g2_a21oi_1 _6856_ (.A1(net1302),
    .A2(_0765_),
    .Y(_2779_),
    .B1(_0746_));
 sg13g2_nand2_1 _6857_ (.Y(_2780_),
    .A(_2778_),
    .B(_2779_));
 sg13g2_xnor2_1 _6858_ (.Y(_2781_),
    .A(_2778_),
    .B(_2779_));
 sg13g2_o21ai_1 _6859_ (.B1(net1),
    .Y(_2782_),
    .A1(net1248),
    .A2(net1153));
 sg13g2_a21oi_1 _6860_ (.A1(net1152),
    .A2(_2781_),
    .Y(_0255_),
    .B1(_2782_));
 sg13g2_o21ai_1 _6861_ (.B1(_2780_),
    .Y(_2783_),
    .A1(_2825_),
    .A2(net1302));
 sg13g2_nand2b_1 _6862_ (.Y(_2784_),
    .B(net1302),
    .A_N(net1244));
 sg13g2_xnor2_1 _6863_ (.Y(_2785_),
    .A(net1244),
    .B(net368));
 sg13g2_xnor2_1 _6864_ (.Y(_2786_),
    .A(_2783_),
    .B(_2785_));
 sg13g2_o21ai_1 _6865_ (.B1(net1417),
    .Y(_2787_),
    .A1(net1244),
    .A2(net1152));
 sg13g2_a21oi_1 _6866_ (.A1(net1153),
    .A2(_2786_),
    .Y(_0256_),
    .B1(_2787_));
 sg13g2_xnor2_1 _6867_ (.Y(_2788_),
    .A(net1240),
    .B(net1302));
 sg13g2_inv_1 _6868_ (.Y(_2789_),
    .A(_2788_));
 sg13g2_a21o_1 _6869_ (.A2(_2851_),
    .A1(net1244),
    .B1(_2783_),
    .X(_2790_));
 sg13g2_nand2_1 _6870_ (.Y(_2791_),
    .A(_2784_),
    .B(_2790_));
 sg13g2_nand3_1 _6871_ (.B(_2788_),
    .C(_2790_),
    .A(_2784_),
    .Y(_2792_));
 sg13g2_a21oi_1 _6872_ (.A1(_2789_),
    .A2(_2791_),
    .Y(_2793_),
    .B1(net1147));
 sg13g2_a22oi_1 _6873_ (.Y(_2794_),
    .B1(_2792_),
    .B2(_2793_),
    .A2(net1147),
    .A1(net1240));
 sg13g2_nand2_1 _6874_ (.Y(_0257_),
    .A(net1417),
    .B(_2794_));
 sg13g2_o21ai_1 _6875_ (.B1(net1417),
    .Y(_2795_),
    .A1(_2823_),
    .A2(net1152));
 sg13g2_xor2_1 _6876_ (.B(net1302),
    .A(net1238),
    .X(_2796_));
 sg13g2_o21ai_1 _6877_ (.B1(_2792_),
    .Y(_2797_),
    .A1(_2824_),
    .A2(net1301));
 sg13g2_xnor2_1 _6878_ (.Y(_2798_),
    .A(_2796_),
    .B(_2797_));
 sg13g2_a21o_1 _6879_ (.A2(_2798_),
    .A1(net1152),
    .B1(_2795_),
    .X(_0258_));
 sg13g2_nor2_1 _6880_ (.A(net1227),
    .B(net1301),
    .Y(_2799_));
 sg13g2_xor2_1 _6881_ (.B(net1301),
    .A(net1234),
    .X(_2800_));
 sg13g2_or2_1 _6882_ (.X(_2801_),
    .B(_2796_),
    .A(_2792_));
 sg13g2_o21ai_1 _6883_ (.B1(_2851_),
    .Y(_2802_),
    .A1(net1238),
    .A2(net1240));
 sg13g2_a21oi_1 _6884_ (.A1(_2823_),
    .A2(_2824_),
    .Y(_2803_),
    .B1(net1301));
 sg13g2_and3_1 _6885_ (.X(_2804_),
    .A(_2800_),
    .B(_2801_),
    .C(_2802_));
 sg13g2_a21oi_1 _6886_ (.A1(_2801_),
    .A2(_2802_),
    .Y(_2805_),
    .B1(_2800_));
 sg13g2_o21ai_1 _6887_ (.B1(net1152),
    .Y(_2806_),
    .A1(_2804_),
    .A2(_2805_));
 sg13g2_o21ai_1 _6888_ (.B1(_2806_),
    .Y(_2807_),
    .A1(net1234),
    .A2(net1152));
 sg13g2_nor2_1 _6889_ (.A(net1415),
    .B(_2807_),
    .Y(_0259_));
 sg13g2_nor2_1 _6890_ (.A(net1233),
    .B(_2851_),
    .Y(_2808_));
 sg13g2_nor2_1 _6891_ (.A(net1228),
    .B(net1301),
    .Y(_2809_));
 sg13g2_or2_1 _6892_ (.X(_2810_),
    .B(_2809_),
    .A(_2808_));
 sg13g2_o21ai_1 _6893_ (.B1(_2810_),
    .Y(_2811_),
    .A1(_2799_),
    .A2(_2805_));
 sg13g2_nor3_1 _6894_ (.A(_2799_),
    .B(_2805_),
    .C(_2810_),
    .Y(_2812_));
 sg13g2_nor2_1 _6895_ (.A(net1146),
    .B(_2812_),
    .Y(_2813_));
 sg13g2_a221oi_1 _6896_ (.B2(_2813_),
    .C1(net1415),
    .B1(_2811_),
    .A1(net1228),
    .Y(_0260_),
    .A2(net1146));
 sg13g2_nor3_1 _6897_ (.A(_2800_),
    .B(_2801_),
    .C(_2808_),
    .Y(_2814_));
 sg13g2_nor4_1 _6898_ (.A(_2799_),
    .B(_2803_),
    .C(_2809_),
    .D(_2814_),
    .Y(_2815_));
 sg13g2_nor2_1 _6899_ (.A(net1301),
    .B(_2815_),
    .Y(_2816_));
 sg13g2_a21oi_1 _6900_ (.A1(net1301),
    .A2(_2815_),
    .Y(_2817_),
    .B1(net1147));
 sg13g2_nor2b_1 _6901_ (.A(_2816_),
    .B_N(_2817_),
    .Y(_2818_));
 sg13g2_o21ai_1 _6902_ (.B1(net1417),
    .Y(_2819_),
    .A1(net1231),
    .A2(_2818_));
 sg13g2_a21oi_1 _6903_ (.A1(net1231),
    .A2(_2818_),
    .Y(_0261_),
    .B1(_2819_));
 sg13g2_nand2b_1 _6904_ (.Y(_0262_),
    .B(_3064_),
    .A_N(_0002_));
 sg13g2_a21o_1 _6905_ (.A2(_3063_),
    .A1(net311),
    .B1(net1166),
    .X(_0096_));
 sg13g2_dfrbp_1 _6906_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net95),
    .D(_0081_),
    .Q_N(\lgA2.rx[0] ),
    .Q(\barrier1.col_idx[0] ));
 sg13g2_dfrbp_1 _6907_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net94),
    .D(_0082_),
    .Q_N(_0044_),
    .Q(\barrier1.col_idx[1] ));
 sg13g2_dfrbp_1 _6908_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net93),
    .D(_0083_),
    .Q_N(_0042_),
    .Q(\barrier1.pix_x[2] ));
 sg13g2_dfrbp_1 _6909_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net92),
    .D(_0084_),
    .Q_N(_0033_),
    .Q(\barrier1.pix_x[3] ));
 sg13g2_dfrbp_1 _6910_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net91),
    .D(_0085_),
    .Q_N(_0029_),
    .Q(\barrier1.pix_x[4] ));
 sg13g2_dfrbp_1 _6911_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net90),
    .D(_0086_),
    .Q_N(_0028_),
    .Q(\barrier1.pix_x[5] ));
 sg13g2_dfrbp_1 _6912_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net89),
    .D(_0087_),
    .Q_N(_0027_),
    .Q(\barrier1.pix_x[6] ));
 sg13g2_dfrbp_1 _6913_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net88),
    .D(_0088_),
    .Q_N(_0036_),
    .Q(\barrier1.pix_x[7] ));
 sg13g2_dfrbp_1 _6914_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net87),
    .D(_0089_),
    .Q_N(_0038_),
    .Q(\barrier1.pix_x[8] ));
 sg13g2_dfrbp_1 _6915_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net86),
    .D(_0090_),
    .Q_N(_0008_),
    .Q(\barrier1.pix_x[9] ));
 sg13g2_dfrbp_1 _6916_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net85),
    .D(_0091_),
    .Q_N(_3447_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _6917_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net84),
    .D(_0092_),
    .Q_N(_3446_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _6918_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net83),
    .D(_0093_),
    .Q_N(_3445_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _6919_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net82),
    .D(_0094_),
    .Q_N(_3444_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _6920_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net81),
    .D(net219),
    .Q_N(_0080_),
    .Q(\draw_score_inst.digit_health[0] ));
 sg13g2_dfrbp_1 _6921_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net79),
    .D(_0096_),
    .Q_N(_3443_),
    .Q(\draw_score_inst.digit_health[1] ));
 sg13g2_dfrbp_1 _6922_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net77),
    .D(_0097_),
    .Q_N(_3442_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _6923_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net76),
    .D(_0098_),
    .Q_N(_3441_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _6924_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net75),
    .D(_0099_),
    .Q_N(_0077_),
    .Q(\pb_x[0] ));
 sg13g2_dfrbp_1 _6925_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net73),
    .D(_0100_),
    .Q_N(_3440_),
    .Q(\pb_x[1] ));
 sg13g2_dfrbp_1 _6926_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net71),
    .D(_0101_),
    .Q_N(_0005_),
    .Q(\pb_x[2] ));
 sg13g2_dfrbp_1 _6927_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net69),
    .D(net295),
    .Q_N(_0069_),
    .Q(\pb_x[3] ));
 sg13g2_dfrbp_1 _6928_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net67),
    .D(_0103_),
    .Q_N(_0068_),
    .Q(\pb_x[4] ));
 sg13g2_dfrbp_1 _6929_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net65),
    .D(_0104_),
    .Q_N(_0066_),
    .Q(\pb_x[5] ));
 sg13g2_dfrbp_1 _6930_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net63),
    .D(net378),
    .Q_N(_0065_),
    .Q(\pb_x[6] ));
 sg13g2_dfrbp_1 _6931_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net61),
    .D(_0106_),
    .Q_N(_0060_),
    .Q(\pb_x[7] ));
 sg13g2_dfrbp_1 _6932_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net59),
    .D(_0107_),
    .Q_N(_0059_),
    .Q(\pb_x[8] ));
 sg13g2_dfrbp_1 _6933_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net57),
    .D(_0108_),
    .Q_N(_0058_),
    .Q(\pb_x[9] ));
 sg13g2_dfrbp_1 _6934_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net55),
    .D(_0109_),
    .Q_N(_0054_),
    .Q(pb_active));
 sg13g2_dfrbp_1 _6935_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net54),
    .D(net224),
    .Q_N(_0009_),
    .Q(\pb_y[0] ));
 sg13g2_dfrbp_1 _6936_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net53),
    .D(_0111_),
    .Q_N(_3439_),
    .Q(\pb_y[1] ));
 sg13g2_dfrbp_1 _6937_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net52),
    .D(_0112_),
    .Q_N(_3438_),
    .Q(\pb_y[2] ));
 sg13g2_dfrbp_1 _6938_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net51),
    .D(_0113_),
    .Q_N(_3437_),
    .Q(\pb_y[3] ));
 sg13g2_dfrbp_1 _6939_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net50),
    .D(_0114_),
    .Q_N(_0073_),
    .Q(\pb_y[4] ));
 sg13g2_dfrbp_1 _6940_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net49),
    .D(_0115_),
    .Q_N(_0072_),
    .Q(\pb_y[5] ));
 sg13g2_dfrbp_1 _6941_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net48),
    .D(_0116_),
    .Q_N(_3436_),
    .Q(\pb_y[6] ));
 sg13g2_dfrbp_1 _6942_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net47),
    .D(_0117_),
    .Q_N(_0071_),
    .Q(\pb_y[7] ));
 sg13g2_dfrbp_1 _6943_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net46),
    .D(_0118_),
    .Q_N(_3435_),
    .Q(\pb_y[8] ));
 sg13g2_dfrbp_1 _6944_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net45),
    .D(net322),
    .Q_N(_3434_),
    .Q(\pb_y[9] ));
 sg13g2_dfrbp_1 _6945_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net44),
    .D(_0120_),
    .Q_N(_0030_),
    .Q(abullet_active));
 sg13g2_dfrbp_1 _6946_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net42),
    .D(net376),
    .Q_N(_3433_),
    .Q(\abullet_x[0] ));
 sg13g2_dfrbp_1 _6947_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net40),
    .D(_0122_),
    .Q_N(_3432_),
    .Q(\abullet_x[1] ));
 sg13g2_dfrbp_1 _6948_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net38),
    .D(net285),
    .Q_N(_3431_),
    .Q(\abullet_x[2] ));
 sg13g2_dfrbp_1 _6949_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net36),
    .D(net320),
    .Q_N(_0045_),
    .Q(\abullet_x[3] ));
 sg13g2_dfrbp_1 _6950_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net34),
    .D(_0125_),
    .Q_N(_3430_),
    .Q(\abullet_x[4] ));
 sg13g2_dfrbp_1 _6951_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net32),
    .D(_0126_),
    .Q_N(_0040_),
    .Q(\abullet_x[5] ));
 sg13g2_dfrbp_1 _6952_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net30),
    .D(_0127_),
    .Q_N(_0039_),
    .Q(\abullet_x[6] ));
 sg13g2_dfrbp_1 _6953_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net28),
    .D(_0128_),
    .Q_N(_0035_),
    .Q(\abullet_x[7] ));
 sg13g2_dfrbp_1 _6954_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net26),
    .D(_0129_),
    .Q_N(_0034_),
    .Q(\abullet_x[8] ));
 sg13g2_dfrbp_1 _6955_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net24),
    .D(_0130_),
    .Q_N(_0031_),
    .Q(\abullet_x[9] ));
 sg13g2_dfrbp_1 _6956_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net22),
    .D(_0131_),
    .Q_N(_3429_),
    .Q(\lfsr[0] ));
 sg13g2_dfrbp_1 _6957_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net217),
    .D(net249),
    .Q_N(_3428_),
    .Q(\lfsr[1] ));
 sg13g2_dfrbp_1 _6958_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net215),
    .D(_0133_),
    .Q_N(_3427_),
    .Q(\lfsr[2] ));
 sg13g2_dfrbp_1 _6959_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net213),
    .D(net234),
    .Q_N(_3426_),
    .Q(\lfsr[3] ));
 sg13g2_dfrbp_1 _6960_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net211),
    .D(net262),
    .Q_N(_3425_),
    .Q(\lfsr[4] ));
 sg13g2_dfrbp_1 _6961_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net209),
    .D(_0136_),
    .Q_N(_3424_),
    .Q(\lfsr[5] ));
 sg13g2_dfrbp_1 _6962_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net205),
    .D(_0137_),
    .Q_N(_3423_),
    .Q(\lfsr[6] ));
 sg13g2_dfrbp_1 _6963_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net203),
    .D(_0138_),
    .Q_N(_3422_),
    .Q(\lfsr[7] ));
 sg13g2_dfrbp_1 _6964_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net201),
    .D(net306),
    .Q_N(_3421_),
    .Q(\selectedRowRand[0] ));
 sg13g2_dfrbp_1 _6965_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net199),
    .D(net246),
    .Q_N(_3420_),
    .Q(\selectedRowRand[1] ));
 sg13g2_dfrbp_1 _6966_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net197),
    .D(net314),
    .Q_N(_0063_),
    .Q(\selectedRowRand[2] ));
 sg13g2_dfrbp_1 _6967_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net195),
    .D(_0142_),
    .Q_N(_3419_),
    .Q(\colRand[0] ));
 sg13g2_dfrbp_1 _6968_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net193),
    .D(_0143_),
    .Q_N(_3418_),
    .Q(\colRand[1] ));
 sg13g2_dfrbp_1 _6969_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net191),
    .D(net274),
    .Q_N(_0067_),
    .Q(\colRand[2] ));
 sg13g2_dfrbp_1 _6970_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net189),
    .D(net384),
    .Q_N(_0025_),
    .Q(\draw_score_inst.score[1] ));
 sg13g2_dfrbp_1 _6971_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net187),
    .D(net336),
    .Q_N(_0026_),
    .Q(\draw_score_inst.score[2] ));
 sg13g2_dfrbp_1 _6972_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net185),
    .D(_0147_),
    .Q_N(_0018_),
    .Q(\draw_score_inst.score[3] ));
 sg13g2_dfrbp_1 _6973_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net181),
    .D(net343),
    .Q_N(_0024_),
    .Q(\draw_score_inst.score[4] ));
 sg13g2_dfrbp_1 _6974_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net179),
    .D(_0149_),
    .Q_N(_0023_),
    .Q(\draw_score_inst.score[5] ));
 sg13g2_dfrbp_1 _6975_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net177),
    .D(_0150_),
    .Q_N(_0022_),
    .Q(\draw_score_inst.score[6] ));
 sg13g2_dfrbp_1 _6976_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net175),
    .D(_0151_),
    .Q_N(_0021_),
    .Q(\draw_score_inst.score[7] ));
 sg13g2_dfrbp_1 _6977_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net173),
    .D(_0152_),
    .Q_N(_0020_),
    .Q(\draw_score_inst.score[8] ));
 sg13g2_dfrbp_1 _6978_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net171),
    .D(_0153_),
    .Q_N(_0019_),
    .Q(\draw_score_inst.score[9] ));
 sg13g2_dfrbp_1 _6979_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net183),
    .D(net260),
    .Q_N(_3448_),
    .Q(game_over));
 sg13g2_dfrbp_1 _6980_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net169),
    .D(_0000_),
    .Q_N(_3417_),
    .Q(game_won));
 sg13g2_dfrbp_1 _6981_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net167),
    .D(_0155_),
    .Q_N(_3416_),
    .Q(\aliens_alive[0] ));
 sg13g2_dfrbp_1 _6982_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net165),
    .D(_0156_),
    .Q_N(_3415_),
    .Q(\aliens_alive[1] ));
 sg13g2_dfrbp_1 _6983_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net163),
    .D(_0157_),
    .Q_N(_3414_),
    .Q(\aliens_alive[2] ));
 sg13g2_dfrbp_1 _6984_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net161),
    .D(_0158_),
    .Q_N(_3413_),
    .Q(\aliens_alive[3] ));
 sg13g2_dfrbp_1 _6985_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net159),
    .D(_0159_),
    .Q_N(_3412_),
    .Q(\aliens_alive[4] ));
 sg13g2_dfrbp_1 _6986_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net157),
    .D(_0160_),
    .Q_N(_3411_),
    .Q(\aliens_alive[5] ));
 sg13g2_dfrbp_1 _6987_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net155),
    .D(_0161_),
    .Q_N(_3410_),
    .Q(\aliens_alive[6] ));
 sg13g2_dfrbp_1 _6988_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net153),
    .D(_0162_),
    .Q_N(_3409_),
    .Q(\aliens_alive[7] ));
 sg13g2_dfrbp_1 _6989_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net151),
    .D(_0163_),
    .Q_N(_0006_),
    .Q(\aliens_alive[8] ));
 sg13g2_dfrbp_1 _6990_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net149),
    .D(_0164_),
    .Q_N(_3408_),
    .Q(\aliens_alive[9] ));
 sg13g2_dfrbp_1 _6991_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net147),
    .D(_0165_),
    .Q_N(_3407_),
    .Q(\aliens_alive[10] ));
 sg13g2_dfrbp_1 _6992_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net145),
    .D(_0166_),
    .Q_N(_3406_),
    .Q(\aliens_alive[11] ));
 sg13g2_dfrbp_1 _6993_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net143),
    .D(_0167_),
    .Q_N(_3405_),
    .Q(\aliens_alive[12] ));
 sg13g2_dfrbp_1 _6994_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net141),
    .D(_0168_),
    .Q_N(_3404_),
    .Q(\aliens_alive[13] ));
 sg13g2_dfrbp_1 _6995_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net139),
    .D(_0169_),
    .Q_N(_3403_),
    .Q(\aliens_alive[14] ));
 sg13g2_dfrbp_1 _6996_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net137),
    .D(_0170_),
    .Q_N(_3402_),
    .Q(\aliens_alive[15] ));
 sg13g2_dfrbp_1 _6997_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net135),
    .D(_0171_),
    .Q_N(_3401_),
    .Q(\aliens_alive[16] ));
 sg13g2_dfrbp_1 _6998_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net133),
    .D(_0172_),
    .Q_N(_3400_),
    .Q(\aliens_alive[17] ));
 sg13g2_dfrbp_1 _6999_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net131),
    .D(_0173_),
    .Q_N(_3399_),
    .Q(\aliens_alive[18] ));
 sg13g2_dfrbp_1 _7000_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net129),
    .D(_0174_),
    .Q_N(_3398_),
    .Q(\aliens_alive[19] ));
 sg13g2_dfrbp_1 _7001_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net127),
    .D(_0175_),
    .Q_N(_3397_),
    .Q(\aliens_alive[20] ));
 sg13g2_dfrbp_1 _7002_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net125),
    .D(_0176_),
    .Q_N(_3396_),
    .Q(\aliens_alive[21] ));
 sg13g2_dfrbp_1 _7003_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net123),
    .D(_0177_),
    .Q_N(_3395_),
    .Q(\aliens_alive[22] ));
 sg13g2_dfrbp_1 _7004_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net121),
    .D(_0178_),
    .Q_N(_3394_),
    .Q(\aliens_alive[23] ));
 sg13g2_dfrbp_1 _7005_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net119),
    .D(_0179_),
    .Q_N(_3393_),
    .Q(\aliens_alive[24] ));
 sg13g2_dfrbp_1 _7006_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net117),
    .D(_0180_),
    .Q_N(_3392_),
    .Q(\aliens_alive[25] ));
 sg13g2_dfrbp_1 _7007_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net115),
    .D(_0181_),
    .Q_N(_3391_),
    .Q(\aliens_alive[26] ));
 sg13g2_dfrbp_1 _7008_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net113),
    .D(_0182_),
    .Q_N(_3390_),
    .Q(\aliens_alive[27] ));
 sg13g2_dfrbp_1 _7009_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net111),
    .D(_0183_),
    .Q_N(_3389_),
    .Q(\aliens_alive[28] ));
 sg13g2_dfrbp_1 _7010_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net109),
    .D(_0184_),
    .Q_N(_3388_),
    .Q(\aliens_alive[29] ));
 sg13g2_dfrbp_1 _7011_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net107),
    .D(_0185_),
    .Q_N(_3387_),
    .Q(\aliens_alive[30] ));
 sg13g2_dfrbp_1 _7012_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net105),
    .D(_0186_),
    .Q_N(_3386_),
    .Q(\aliens_alive[31] ));
 sg13g2_dfrbp_1 _7013_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net103),
    .D(_0187_),
    .Q_N(_3385_),
    .Q(\aliens_alive[32] ));
 sg13g2_dfrbp_1 _7014_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net101),
    .D(_0188_),
    .Q_N(_3384_),
    .Q(\aliens_alive[33] ));
 sg13g2_dfrbp_1 _7015_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net99),
    .D(_0189_),
    .Q_N(_3383_),
    .Q(\aliens_alive[34] ));
 sg13g2_dfrbp_1 _7016_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net97),
    .D(_0190_),
    .Q_N(_3382_),
    .Q(\aliens_alive[35] ));
 sg13g2_dfrbp_1 _7017_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net80),
    .D(_0191_),
    .Q_N(_3381_),
    .Q(\aliens_alive[36] ));
 sg13g2_dfrbp_1 _7018_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net74),
    .D(_0192_),
    .Q_N(_3380_),
    .Q(\aliens_alive[37] ));
 sg13g2_dfrbp_1 _7019_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net70),
    .D(_0193_),
    .Q_N(_3379_),
    .Q(\aliens_alive[38] ));
 sg13g2_dfrbp_1 _7020_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net66),
    .D(_0194_),
    .Q_N(_3378_),
    .Q(\aliens_alive[39] ));
 sg13g2_dfrbp_1 _7021_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net62),
    .D(_0195_),
    .Q_N(_3377_),
    .Q(prev_button2));
 sg13g2_dfrbp_1 _7022_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net60),
    .D(net264),
    .Q_N(_0056_),
    .Q(\barrier_health[0][0] ));
 sg13g2_dfrbp_1 _7023_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net58),
    .D(net317),
    .Q_N(_3376_),
    .Q(\barrier_health[0][1] ));
 sg13g2_dfrbp_1 _7024_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net56),
    .D(net252),
    .Q_N(_3375_),
    .Q(\barrier_health[0][2] ));
 sg13g2_dfrbp_1 _7025_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net43),
    .D(net222),
    .Q_N(_0055_),
    .Q(\barrier_health[1][0] ));
 sg13g2_dfrbp_1 _7026_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net41),
    .D(net354),
    .Q_N(_3374_),
    .Q(\barrier_health[1][1] ));
 sg13g2_dfrbp_1 _7027_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net39),
    .D(_0201_),
    .Q_N(_3373_),
    .Q(\barrier_health[1][2] ));
 sg13g2_dfrbp_1 _7028_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net37),
    .D(_0202_),
    .Q_N(_0053_),
    .Q(\barrier_health[2][0] ));
 sg13g2_dfrbp_1 _7029_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net35),
    .D(net362),
    .Q_N(_3372_),
    .Q(\barrier_health[2][1] ));
 sg13g2_dfrbp_1 _7030_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net33),
    .D(_0204_),
    .Q_N(_3371_),
    .Q(\barrier_health[2][2] ));
 sg13g2_dfrbp_1 _7031_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net31),
    .D(net226),
    .Q_N(_0052_),
    .Q(\barrier_health[3][0] ));
 sg13g2_dfrbp_1 _7032_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net29),
    .D(net349),
    .Q_N(_3370_),
    .Q(\barrier_health[3][1] ));
 sg13g2_dfrbp_1 _7033_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net27),
    .D(_0207_),
    .Q_N(_3369_),
    .Q(\barrier_health[3][2] ));
 sg13g2_dfrbp_1 _7034_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net25),
    .D(_0208_),
    .Q_N(_3368_),
    .Q(\prev_vpos_shooter[0] ));
 sg13g2_dfrbp_1 _7035_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net23),
    .D(_0209_),
    .Q_N(_3367_),
    .Q(\prev_vpos_shooter[1] ));
 sg13g2_dfrbp_1 _7036_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net21),
    .D(_0210_),
    .Q_N(_3366_),
    .Q(\prev_vpos_shooter[2] ));
 sg13g2_dfrbp_1 _7037_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net216),
    .D(_0211_),
    .Q_N(_3365_),
    .Q(\prev_vpos_shooter[3] ));
 sg13g2_dfrbp_1 _7038_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net214),
    .D(_0212_),
    .Q_N(_3364_),
    .Q(\prev_vpos_shooter[4] ));
 sg13g2_dfrbp_1 _7039_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net212),
    .D(_0213_),
    .Q_N(_3363_),
    .Q(\prev_vpos_shooter[5] ));
 sg13g2_dfrbp_1 _7040_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net210),
    .D(_0214_),
    .Q_N(_3362_),
    .Q(\prev_vpos_shooter[6] ));
 sg13g2_dfrbp_1 _7041_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net208),
    .D(_0215_),
    .Q_N(_3361_),
    .Q(\prev_vpos_shooter[7] ));
 sg13g2_dfrbp_1 _7042_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net204),
    .D(_0216_),
    .Q_N(_3360_),
    .Q(\prev_vpos_shooter[8] ));
 sg13g2_dfrbp_1 _7043_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net202),
    .D(_0217_),
    .Q_N(_3359_),
    .Q(\prev_vpos_shooter[9] ));
 sg13g2_dfrbp_1 _7044_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net200),
    .D(_0218_),
    .Q_N(_3358_),
    .Q(prev_button0));
 sg13g2_dfrbp_1 _7045_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net198),
    .D(net230),
    .Q_N(_0007_),
    .Q(move_dir));
 sg13g2_dfrbp_1 _7046_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net194),
    .D(_0220_),
    .Q_N(_3357_),
    .Q(prev_button1));
 sg13g2_dfrbp_1 _7047_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net192),
    .D(_0221_),
    .Q_N(_3356_),
    .Q(hsync));
 sg13g2_dfrbp_1 _7048_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net190),
    .D(_0222_),
    .Q_N(_3355_),
    .Q(\barrier1.bar_rom.row_index[0] ));
 sg13g2_dfrbp_1 _7049_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net186),
    .D(_0223_),
    .Q_N(_0048_),
    .Q(\barrier1.bar_rom.row_index[1] ));
 sg13g2_dfrbp_1 _7050_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net180),
    .D(_0224_),
    .Q_N(_0010_),
    .Q(\barrier1.bar_rom.row_index[2] ));
 sg13g2_dfrbp_1 _7051_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net176),
    .D(_0225_),
    .Q_N(_0011_),
    .Q(\barrier1.bar_rom.row_index[3] ));
 sg13g2_dfrbp_1 _7052_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net172),
    .D(_0226_),
    .Q_N(_0012_),
    .Q(\barrier1.pix_y[4] ));
 sg13g2_dfrbp_1 _7053_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net168),
    .D(_0227_),
    .Q_N(_0013_),
    .Q(\barrier1.pix_y[5] ));
 sg13g2_dfrbp_1 _7054_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net164),
    .D(_0228_),
    .Q_N(_0014_),
    .Q(\barrier1.pix_y[6] ));
 sg13g2_dfrbp_1 _7055_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net160),
    .D(_0229_),
    .Q_N(_0015_),
    .Q(\barrier1.pix_y[7] ));
 sg13g2_dfrbp_1 _7056_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net156),
    .D(_0230_),
    .Q_N(_0016_),
    .Q(\barrier1.pix_y[8] ));
 sg13g2_dfrbp_1 _7057_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net152),
    .D(_0231_),
    .Q_N(_0017_),
    .Q(\barrier1.pix_y[9] ));
 sg13g2_dfrbp_1 _7058_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net148),
    .D(net236),
    .Q_N(_3354_),
    .Q(\sync_gen.vsync ));
 sg13g2_dfrbp_1 _7059_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net144),
    .D(_0233_),
    .Q_N(_0079_),
    .Q(\myShooter.shooter_left_x[1] ));
 sg13g2_dfrbp_1 _7060_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net140),
    .D(_0234_),
    .Q_N(_3353_),
    .Q(\myShooter.shooter_left_x[2] ));
 sg13g2_dfrbp_1 _7061_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net136),
    .D(_0235_),
    .Q_N(_0046_),
    .Q(\myShooter.shooter_left_x[3] ));
 sg13g2_dfrbp_1 _7062_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net132),
    .D(_0236_),
    .Q_N(_3352_),
    .Q(\myShooter.shooter_left_x[4] ));
 sg13g2_dfrbp_1 _7063_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net128),
    .D(_0237_),
    .Q_N(_0043_),
    .Q(\myShooter.shooter_left_x[5] ));
 sg13g2_dfrbp_1 _7064_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net124),
    .D(_0238_),
    .Q_N(_0041_),
    .Q(\myShooter.shooter_left_x[6] ));
 sg13g2_dfrbp_1 _7065_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net120),
    .D(_0239_),
    .Q_N(_0037_),
    .Q(\myShooter.shooter_left_x[7] ));
 sg13g2_dfrbp_1 _7066_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net116),
    .D(_0240_),
    .Q_N(_0047_),
    .Q(\myShooter.shooter_left_x[8] ));
 sg13g2_dfrbp_1 _7067_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net184),
    .D(_0241_),
    .Q_N(_0032_),
    .Q(\myShooter.shooter_left_x[9] ));
 sg13g2_dfrbp_1 _7068_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net206),
    .D(_0001_),
    .Q_N(_3449_),
    .Q(\draw_score_inst.segment_rom_health.segments[4] ));
 sg13g2_dfrbp_1 _7069_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net112),
    .D(_0002_),
    .Q_N(_3351_),
    .Q(\draw_score_inst.segment_rom_health.segments[6] ));
 sg13g2_dfrbp_1 _7070_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net108),
    .D(_0242_),
    .Q_N(_0062_),
    .Q(\abullet_y[1] ));
 sg13g2_dfrbp_1 _7071_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net104),
    .D(_0243_),
    .Q_N(_3350_),
    .Q(\abullet_y[2] ));
 sg13g2_dfrbp_1 _7072_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net100),
    .D(net339),
    .Q_N(_0064_),
    .Q(\abullet_y[3] ));
 sg13g2_dfrbp_1 _7073_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net96),
    .D(net374),
    .Q_N(_0051_),
    .Q(\abullet_y[4] ));
 sg13g2_dfrbp_1 _7074_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net72),
    .D(net332),
    .Q_N(_3349_),
    .Q(\abullet_y[5] ));
 sg13g2_dfrbp_1 _7075_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net64),
    .D(_0247_),
    .Q_N(_3348_),
    .Q(\abullet_y[6] ));
 sg13g2_dfrbp_1 _7076_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net188),
    .D(_0248_),
    .Q_N(_0050_),
    .Q(\abullet_y[7] ));
 sg13g2_dfrbp_1 _7077_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net178),
    .D(_0249_),
    .Q_N(_3347_),
    .Q(\abullet_y[8] ));
 sg13g2_dfrbp_1 _7078_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net170),
    .D(net334),
    .Q_N(_0049_),
    .Q(\abullet_y[9] ));
 sg13g2_dfrbp_1 _7079_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net162),
    .D(_0251_),
    .Q_N(_3346_),
    .Q(\draw_score_inst.segment_rom_health.segments[5] ));
 sg13g2_dfrbp_1 _7080_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net158),
    .D(_0252_),
    .Q_N(_3345_),
    .Q(\draw_score_inst.segment_rom_health.segments[2] ));
 sg13g2_dfrbp_1 _7081_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net154),
    .D(net282),
    .Q_N(\lA2_x[1] ),
    .Q(\group_x[1] ));
 sg13g2_dfrbp_1 _7082_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net146),
    .D(_0254_),
    .Q_N(_3344_),
    .Q(\group_x[2] ));
 sg13g2_dfrbp_1 _7083_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net138),
    .D(_0255_),
    .Q_N(_0070_),
    .Q(\group_x[3] ));
 sg13g2_dfrbp_1 _7084_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net130),
    .D(_0256_),
    .Q_N(_0076_),
    .Q(\group_x[4] ));
 sg13g2_dfrbp_1 _7085_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net122),
    .D(_0257_),
    .Q_N(_0075_),
    .Q(\group_x[5] ));
 sg13g2_dfrbp_1 _7086_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net114),
    .D(_0258_),
    .Q_N(_0057_),
    .Q(\group_x[6] ));
 sg13g2_dfrbp_1 _7087_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net106),
    .D(_0259_),
    .Q_N(_0061_),
    .Q(\group_x[7] ));
 sg13g2_dfrbp_1 _7088_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net98),
    .D(_0260_),
    .Q_N(_0074_),
    .Q(\group_x[8] ));
 sg13g2_dfrbp_1 _7089_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net68),
    .D(_0261_),
    .Q_N(_0078_),
    .Q(\group_x[9] ));
 sg13g2_dfrbp_1 _7090_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net207),
    .D(_0262_),
    .Q_N(_3450_),
    .Q(\draw_score_inst.segment_rom_health.segments[0] ));
 sg13g2_dfrbp_1 _7091_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net196),
    .D(_0003_),
    .Q_N(_3451_),
    .Q(\movement_dir[1] ));
 sg13g2_dfrbp_1 _7092_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net182),
    .D(_0004_),
    .Q_N(_3343_),
    .Q(\movement_dir[2] ));
 sg13g2_dfrbp_1 _7093_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net174),
    .D(_0263_),
    .Q_N(_3342_),
    .Q(\prev_vpos[0] ));
 sg13g2_dfrbp_1 _7094_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net166),
    .D(_0264_),
    .Q_N(_3341_),
    .Q(\prev_vpos[1] ));
 sg13g2_dfrbp_1 _7095_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net150),
    .D(_0265_),
    .Q_N(_3340_),
    .Q(\prev_vpos[2] ));
 sg13g2_dfrbp_1 _7096_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net142),
    .D(_0266_),
    .Q_N(_3339_),
    .Q(\prev_vpos[3] ));
 sg13g2_dfrbp_1 _7097_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net134),
    .D(_0267_),
    .Q_N(_3338_),
    .Q(\prev_vpos[4] ));
 sg13g2_dfrbp_1 _7098_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net126),
    .D(_0268_),
    .Q_N(_3337_),
    .Q(\prev_vpos[5] ));
 sg13g2_dfrbp_1 _7099_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net118),
    .D(_0269_),
    .Q_N(_3336_),
    .Q(\prev_vpos[6] ));
 sg13g2_dfrbp_1 _7100_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net110),
    .D(_0270_),
    .Q_N(_3335_),
    .Q(\prev_vpos[7] ));
 sg13g2_dfrbp_1 _7101_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net102),
    .D(_0271_),
    .Q_N(_3334_),
    .Q(\prev_vpos[8] ));
 sg13g2_dfrbp_1 _7102_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net78),
    .D(_0272_),
    .Q_N(_3333_),
    .Q(\prev_vpos[9] ));
 sg13g2_tiehi _6956__22 (.L_HI(net22));
 sg13g2_tiehi _7035__23 (.L_HI(net23));
 sg13g2_tiehi _6955__24 (.L_HI(net24));
 sg13g2_tiehi _7034__25 (.L_HI(net25));
 sg13g2_tiehi _6954__26 (.L_HI(net26));
 sg13g2_tiehi _7033__27 (.L_HI(net27));
 sg13g2_tiehi _6953__28 (.L_HI(net28));
 sg13g2_tiehi _7032__29 (.L_HI(net29));
 sg13g2_tiehi _6952__30 (.L_HI(net30));
 sg13g2_tiehi _7031__31 (.L_HI(net31));
 sg13g2_tiehi _6951__32 (.L_HI(net32));
 sg13g2_tiehi _7030__33 (.L_HI(net33));
 sg13g2_tiehi _6950__34 (.L_HI(net34));
 sg13g2_tiehi _7029__35 (.L_HI(net35));
 sg13g2_tiehi _6949__36 (.L_HI(net36));
 sg13g2_tiehi _7028__37 (.L_HI(net37));
 sg13g2_tiehi _6948__38 (.L_HI(net38));
 sg13g2_tiehi _7027__39 (.L_HI(net39));
 sg13g2_tiehi _6947__40 (.L_HI(net40));
 sg13g2_tiehi _7026__41 (.L_HI(net41));
 sg13g2_tiehi _6946__42 (.L_HI(net42));
 sg13g2_tiehi _7025__43 (.L_HI(net43));
 sg13g2_tiehi _6945__44 (.L_HI(net44));
 sg13g2_tiehi _6944__45 (.L_HI(net45));
 sg13g2_tiehi _6943__46 (.L_HI(net46));
 sg13g2_tiehi _6942__47 (.L_HI(net47));
 sg13g2_tiehi _6941__48 (.L_HI(net48));
 sg13g2_tiehi _6940__49 (.L_HI(net49));
 sg13g2_tiehi _6939__50 (.L_HI(net50));
 sg13g2_tiehi _6938__51 (.L_HI(net51));
 sg13g2_tiehi _6937__52 (.L_HI(net52));
 sg13g2_tiehi _6936__53 (.L_HI(net53));
 sg13g2_tiehi _6935__54 (.L_HI(net54));
 sg13g2_tiehi _6934__55 (.L_HI(net55));
 sg13g2_tiehi _7024__56 (.L_HI(net56));
 sg13g2_tiehi _6933__57 (.L_HI(net57));
 sg13g2_tiehi _7023__58 (.L_HI(net58));
 sg13g2_tiehi _6932__59 (.L_HI(net59));
 sg13g2_tiehi _7022__60 (.L_HI(net60));
 sg13g2_tiehi _6931__61 (.L_HI(net61));
 sg13g2_tiehi _7021__62 (.L_HI(net62));
 sg13g2_tiehi _6930__63 (.L_HI(net63));
 sg13g2_tiehi _7075__64 (.L_HI(net64));
 sg13g2_tiehi _6929__65 (.L_HI(net65));
 sg13g2_tiehi _7020__66 (.L_HI(net66));
 sg13g2_tiehi _6928__67 (.L_HI(net67));
 sg13g2_tiehi _7089__68 (.L_HI(net68));
 sg13g2_tiehi _6927__69 (.L_HI(net69));
 sg13g2_tiehi _7019__70 (.L_HI(net70));
 sg13g2_tiehi _6926__71 (.L_HI(net71));
 sg13g2_tiehi _7074__72 (.L_HI(net72));
 sg13g2_tiehi _6925__73 (.L_HI(net73));
 sg13g2_tiehi _7018__74 (.L_HI(net74));
 sg13g2_tiehi _6924__75 (.L_HI(net75));
 sg13g2_tiehi _6923__76 (.L_HI(net76));
 sg13g2_tiehi _6922__77 (.L_HI(net77));
 sg13g2_tiehi _7102__78 (.L_HI(net78));
 sg13g2_tiehi _6921__79 (.L_HI(net79));
 sg13g2_tiehi _7017__80 (.L_HI(net80));
 sg13g2_tiehi _6920__81 (.L_HI(net81));
 sg13g2_tiehi _6919__82 (.L_HI(net82));
 sg13g2_tiehi _6918__83 (.L_HI(net83));
 sg13g2_tiehi _6917__84 (.L_HI(net84));
 sg13g2_tiehi _6916__85 (.L_HI(net85));
 sg13g2_tiehi _6915__86 (.L_HI(net86));
 sg13g2_tiehi _6914__87 (.L_HI(net87));
 sg13g2_tiehi _6913__88 (.L_HI(net88));
 sg13g2_tiehi _6912__89 (.L_HI(net89));
 sg13g2_tiehi _6911__90 (.L_HI(net90));
 sg13g2_tiehi _6910__91 (.L_HI(net91));
 sg13g2_tiehi _6909__92 (.L_HI(net92));
 sg13g2_tiehi _6908__93 (.L_HI(net93));
 sg13g2_tiehi _6907__94 (.L_HI(net94));
 sg13g2_tiehi _6906__95 (.L_HI(net95));
 sg13g2_tiehi _7073__96 (.L_HI(net96));
 sg13g2_tiehi _7016__97 (.L_HI(net97));
 sg13g2_tiehi _7088__98 (.L_HI(net98));
 sg13g2_tiehi _7015__99 (.L_HI(net99));
 sg13g2_tiehi _7072__100 (.L_HI(net100));
 sg13g2_tiehi _7014__101 (.L_HI(net101));
 sg13g2_tiehi _7101__102 (.L_HI(net102));
 sg13g2_tiehi _7013__103 (.L_HI(net103));
 sg13g2_tiehi _7071__104 (.L_HI(net104));
 sg13g2_tiehi _7012__105 (.L_HI(net105));
 sg13g2_tiehi _7087__106 (.L_HI(net106));
 sg13g2_tiehi _7011__107 (.L_HI(net107));
 sg13g2_tiehi _7070__108 (.L_HI(net108));
 sg13g2_tiehi _7010__109 (.L_HI(net109));
 sg13g2_tiehi _7100__110 (.L_HI(net110));
 sg13g2_tiehi _7009__111 (.L_HI(net111));
 sg13g2_tiehi _7069__112 (.L_HI(net112));
 sg13g2_tiehi _7008__113 (.L_HI(net113));
 sg13g2_tiehi _7086__114 (.L_HI(net114));
 sg13g2_tiehi _7007__115 (.L_HI(net115));
 sg13g2_tiehi _7066__116 (.L_HI(net116));
 sg13g2_tiehi _7006__117 (.L_HI(net117));
 sg13g2_tiehi _7099__118 (.L_HI(net118));
 sg13g2_tiehi _7005__119 (.L_HI(net119));
 sg13g2_tiehi _7065__120 (.L_HI(net120));
 sg13g2_tiehi _7004__121 (.L_HI(net121));
 sg13g2_tiehi _7085__122 (.L_HI(net122));
 sg13g2_tiehi _7003__123 (.L_HI(net123));
 sg13g2_tiehi _7064__124 (.L_HI(net124));
 sg13g2_tiehi _7002__125 (.L_HI(net125));
 sg13g2_tiehi _7098__126 (.L_HI(net126));
 sg13g2_tiehi _7001__127 (.L_HI(net127));
 sg13g2_tiehi _7063__128 (.L_HI(net128));
 sg13g2_tiehi _7000__129 (.L_HI(net129));
 sg13g2_tiehi _7084__130 (.L_HI(net130));
 sg13g2_tiehi _6999__131 (.L_HI(net131));
 sg13g2_tiehi _7062__132 (.L_HI(net132));
 sg13g2_tiehi _6998__133 (.L_HI(net133));
 sg13g2_tiehi _7097__134 (.L_HI(net134));
 sg13g2_tiehi _6997__135 (.L_HI(net135));
 sg13g2_tiehi _7061__136 (.L_HI(net136));
 sg13g2_tiehi _6996__137 (.L_HI(net137));
 sg13g2_tiehi _7083__138 (.L_HI(net138));
 sg13g2_tiehi _6995__139 (.L_HI(net139));
 sg13g2_tiehi _7060__140 (.L_HI(net140));
 sg13g2_tiehi _6994__141 (.L_HI(net141));
 sg13g2_tiehi _7096__142 (.L_HI(net142));
 sg13g2_tiehi _6993__143 (.L_HI(net143));
 sg13g2_tiehi _7059__144 (.L_HI(net144));
 sg13g2_tiehi _6992__145 (.L_HI(net145));
 sg13g2_tiehi _7082__146 (.L_HI(net146));
 sg13g2_tiehi _6991__147 (.L_HI(net147));
 sg13g2_tiehi _7058__148 (.L_HI(net148));
 sg13g2_tiehi _6990__149 (.L_HI(net149));
 sg13g2_tiehi _7095__150 (.L_HI(net150));
 sg13g2_tiehi _6989__151 (.L_HI(net151));
 sg13g2_tiehi _7057__152 (.L_HI(net152));
 sg13g2_tiehi _6988__153 (.L_HI(net153));
 sg13g2_tiehi _7081__154 (.L_HI(net154));
 sg13g2_tiehi _6987__155 (.L_HI(net155));
 sg13g2_tiehi _7056__156 (.L_HI(net156));
 sg13g2_tiehi _6986__157 (.L_HI(net157));
 sg13g2_tiehi _7080__158 (.L_HI(net158));
 sg13g2_tiehi _6985__159 (.L_HI(net159));
 sg13g2_tiehi _7055__160 (.L_HI(net160));
 sg13g2_tiehi _6984__161 (.L_HI(net161));
 sg13g2_tiehi _7079__162 (.L_HI(net162));
 sg13g2_tiehi _6983__163 (.L_HI(net163));
 sg13g2_tiehi _7054__164 (.L_HI(net164));
 sg13g2_tiehi _6982__165 (.L_HI(net165));
 sg13g2_tiehi _7094__166 (.L_HI(net166));
 sg13g2_tiehi _6981__167 (.L_HI(net167));
 sg13g2_tiehi _7053__168 (.L_HI(net168));
 sg13g2_tiehi _6980__169 (.L_HI(net169));
 sg13g2_tiehi _7078__170 (.L_HI(net170));
 sg13g2_tiehi _6978__171 (.L_HI(net171));
 sg13g2_tiehi _7052__172 (.L_HI(net172));
 sg13g2_tiehi _6977__173 (.L_HI(net173));
 sg13g2_tiehi _7093__174 (.L_HI(net174));
 sg13g2_tiehi _6976__175 (.L_HI(net175));
 sg13g2_tiehi _7051__176 (.L_HI(net176));
 sg13g2_tiehi _6975__177 (.L_HI(net177));
 sg13g2_tiehi _7077__178 (.L_HI(net178));
 sg13g2_tiehi _6974__179 (.L_HI(net179));
 sg13g2_tiehi _7050__180 (.L_HI(net180));
 sg13g2_tiehi _6973__181 (.L_HI(net181));
 sg13g2_tiehi _7092__182 (.L_HI(net182));
 sg13g2_tiehi _6979__183 (.L_HI(net183));
 sg13g2_tiehi _7067__184 (.L_HI(net184));
 sg13g2_tiehi _6972__185 (.L_HI(net185));
 sg13g2_tiehi _7049__186 (.L_HI(net186));
 sg13g2_tiehi _6971__187 (.L_HI(net187));
 sg13g2_tiehi _7076__188 (.L_HI(net188));
 sg13g2_tiehi _6970__189 (.L_HI(net189));
 sg13g2_tiehi _7048__190 (.L_HI(net190));
 sg13g2_tiehi _6969__191 (.L_HI(net191));
 sg13g2_tiehi _7047__192 (.L_HI(net192));
 sg13g2_tiehi _6968__193 (.L_HI(net193));
 sg13g2_tiehi _7046__194 (.L_HI(net194));
 sg13g2_tiehi _6967__195 (.L_HI(net195));
 sg13g2_tiehi _7091__196 (.L_HI(net196));
 sg13g2_tiehi _6966__197 (.L_HI(net197));
 sg13g2_tiehi _7045__198 (.L_HI(net198));
 sg13g2_tiehi _6965__199 (.L_HI(net199));
 sg13g2_tiehi _7044__200 (.L_HI(net200));
 sg13g2_tiehi _6964__201 (.L_HI(net201));
 sg13g2_tiehi _7043__202 (.L_HI(net202));
 sg13g2_tiehi _6963__203 (.L_HI(net203));
 sg13g2_tiehi _7042__204 (.L_HI(net204));
 sg13g2_tiehi _6962__205 (.L_HI(net205));
 sg13g2_tiehi _7068__206 (.L_HI(net206));
 sg13g2_tiehi _7090__207 (.L_HI(net207));
 sg13g2_tiehi _7041__208 (.L_HI(net208));
 sg13g2_tiehi _6961__209 (.L_HI(net209));
 sg13g2_tiehi _7040__210 (.L_HI(net210));
 sg13g2_tiehi _6960__211 (.L_HI(net211));
 sg13g2_tiehi _7039__212 (.L_HI(net212));
 sg13g2_tiehi _6959__213 (.L_HI(net213));
 sg13g2_tiehi _7038__214 (.L_HI(net214));
 sg13g2_tiehi _6958__215 (.L_HI(net215));
 sg13g2_tiehi _7037__216 (.L_HI(net216));
 sg13g2_tiehi _6957__217 (.L_HI(net217));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_space_invaders_game_6 (.L_LO(net6));
 sg13g2_tielo tt_um_space_invaders_game_7 (.L_LO(net7));
 sg13g2_tielo tt_um_space_invaders_game_8 (.L_LO(net8));
 sg13g2_tielo tt_um_space_invaders_game_9 (.L_LO(net9));
 sg13g2_tielo tt_um_space_invaders_game_10 (.L_LO(net10));
 sg13g2_tielo tt_um_space_invaders_game_11 (.L_LO(net11));
 sg13g2_tielo tt_um_space_invaders_game_12 (.L_LO(net12));
 sg13g2_tielo tt_um_space_invaders_game_13 (.L_LO(net13));
 sg13g2_tielo tt_um_space_invaders_game_14 (.L_LO(net14));
 sg13g2_tielo tt_um_space_invaders_game_15 (.L_LO(net15));
 sg13g2_tielo tt_um_space_invaders_game_16 (.L_LO(net16));
 sg13g2_tielo tt_um_space_invaders_game_17 (.L_LO(net17));
 sg13g2_tielo tt_um_space_invaders_game_18 (.L_LO(net18));
 sg13g2_tielo tt_um_space_invaders_game_19 (.L_LO(net19));
 sg13g2_tielo tt_um_space_invaders_game_20 (.L_LO(net20));
 sg13g2_tiehi _7036__21 (.L_HI(net21));
 sg13g2_buf_2 _7316_ (.A(\sync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_2 _7317_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout1074 (.X(net1074),
    .A(_2472_));
 sg13g2_buf_4 fanout1075 (.X(net1075),
    .A(_2471_));
 sg13g2_buf_2 fanout1076 (.A(net1077),
    .X(net1076));
 sg13g2_buf_2 fanout1077 (.A(_2234_),
    .X(net1077));
 sg13g2_buf_2 fanout1078 (.A(_2186_),
    .X(net1078));
 sg13g2_buf_1 fanout1079 (.A(_2186_),
    .X(net1079));
 sg13g2_buf_2 fanout1080 (.A(_1434_),
    .X(net1080));
 sg13g2_buf_2 fanout1081 (.A(_2693_),
    .X(net1081));
 sg13g2_buf_2 fanout1082 (.A(_2693_),
    .X(net1082));
 sg13g2_buf_4 fanout1083 (.X(net1083),
    .A(_2656_));
 sg13g2_buf_2 fanout1084 (.A(net1085),
    .X(net1084));
 sg13g2_buf_2 fanout1085 (.A(net1086),
    .X(net1085));
 sg13g2_buf_2 fanout1086 (.A(_0642_),
    .X(net1086));
 sg13g2_buf_4 fanout1087 (.X(net1087),
    .A(_0641_));
 sg13g2_buf_4 fanout1088 (.X(net1088),
    .A(_3079_));
 sg13g2_buf_2 fanout1089 (.A(_3079_),
    .X(net1089));
 sg13g2_buf_2 fanout1090 (.A(_2729_),
    .X(net1090));
 sg13g2_buf_2 fanout1091 (.A(net1092),
    .X(net1091));
 sg13g2_buf_1 fanout1092 (.A(net1094),
    .X(net1092));
 sg13g2_buf_2 fanout1093 (.A(net1094),
    .X(net1093));
 sg13g2_buf_1 fanout1094 (.A(net1097),
    .X(net1094));
 sg13g2_buf_2 fanout1095 (.A(net1096),
    .X(net1095));
 sg13g2_buf_2 fanout1096 (.A(net1097),
    .X(net1096));
 sg13g2_buf_4 fanout1097 (.X(net1097),
    .A(_2545_));
 sg13g2_buf_2 fanout1098 (.A(net1099),
    .X(net1098));
 sg13g2_buf_2 fanout1099 (.A(net1100),
    .X(net1099));
 sg13g2_buf_2 fanout1100 (.A(_2368_),
    .X(net1100));
 sg13g2_buf_2 fanout1101 (.A(_2368_),
    .X(net1101));
 sg13g2_buf_2 fanout1102 (.A(net1104),
    .X(net1102));
 sg13g2_buf_2 fanout1103 (.A(net1104),
    .X(net1103));
 sg13g2_buf_1 fanout1104 (.A(net1114),
    .X(net1104));
 sg13g2_buf_2 fanout1105 (.A(net1106),
    .X(net1105));
 sg13g2_buf_1 fanout1106 (.A(net1114),
    .X(net1106));
 sg13g2_buf_2 fanout1107 (.A(net1108),
    .X(net1107));
 sg13g2_buf_1 fanout1108 (.A(net1109),
    .X(net1108));
 sg13g2_buf_1 fanout1109 (.A(net1114),
    .X(net1109));
 sg13g2_buf_2 fanout1110 (.A(net1113),
    .X(net1110));
 sg13g2_buf_2 fanout1111 (.A(net1113),
    .X(net1111));
 sg13g2_buf_1 fanout1112 (.A(net1113),
    .X(net1112));
 sg13g2_buf_1 fanout1113 (.A(net1114),
    .X(net1113));
 sg13g2_buf_2 fanout1114 (.A(_0643_),
    .X(net1114));
 sg13g2_buf_2 fanout1115 (.A(_0904_),
    .X(net1115));
 sg13g2_buf_2 fanout1116 (.A(_0904_),
    .X(net1116));
 sg13g2_buf_2 fanout1117 (.A(net1118),
    .X(net1117));
 sg13g2_buf_2 fanout1118 (.A(_0903_),
    .X(net1118));
 sg13g2_buf_4 fanout1119 (.X(net1119),
    .A(_0831_));
 sg13g2_buf_2 fanout1120 (.A(_0801_),
    .X(net1120));
 sg13g2_buf_2 fanout1121 (.A(net1122),
    .X(net1121));
 sg13g2_buf_4 fanout1122 (.X(net1122),
    .A(_0800_));
 sg13g2_buf_2 fanout1123 (.A(net1124),
    .X(net1123));
 sg13g2_buf_2 fanout1124 (.A(net1129),
    .X(net1124));
 sg13g2_buf_2 fanout1125 (.A(net1126),
    .X(net1125));
 sg13g2_buf_2 fanout1126 (.A(net1129),
    .X(net1126));
 sg13g2_buf_2 fanout1127 (.A(net1129),
    .X(net1127));
 sg13g2_buf_1 fanout1128 (.A(net1129),
    .X(net1128));
 sg13g2_buf_2 fanout1129 (.A(_0532_),
    .X(net1129));
 sg13g2_buf_2 fanout1130 (.A(net1132),
    .X(net1130));
 sg13g2_buf_1 fanout1131 (.A(net1132),
    .X(net1131));
 sg13g2_buf_1 fanout1132 (.A(net1133),
    .X(net1132));
 sg13g2_buf_2 fanout1133 (.A(_0532_),
    .X(net1133));
 sg13g2_buf_4 fanout1134 (.X(net1134),
    .A(_3271_));
 sg13g2_buf_2 fanout1135 (.A(_3271_),
    .X(net1135));
 sg13g2_buf_4 fanout1136 (.X(net1136),
    .A(_3264_));
 sg13g2_buf_2 fanout1137 (.A(_3264_),
    .X(net1137));
 sg13g2_buf_2 fanout1138 (.A(net1139),
    .X(net1138));
 sg13g2_buf_2 fanout1139 (.A(_3261_),
    .X(net1139));
 sg13g2_buf_2 fanout1140 (.A(net1141),
    .X(net1140));
 sg13g2_buf_2 fanout1141 (.A(_3254_),
    .X(net1141));
 sg13g2_buf_2 fanout1142 (.A(_3241_),
    .X(net1142));
 sg13g2_buf_2 fanout1143 (.A(_3240_),
    .X(net1143));
 sg13g2_buf_4 fanout1144 (.X(net1144),
    .A(net1148));
 sg13g2_buf_1 fanout1145 (.A(net1148),
    .X(net1145));
 sg13g2_buf_4 fanout1146 (.X(net1146),
    .A(net1148));
 sg13g2_buf_2 fanout1147 (.A(net1148),
    .X(net1147));
 sg13g2_buf_4 fanout1148 (.X(net1148),
    .A(_3057_));
 sg13g2_buf_2 fanout1149 (.A(net1150),
    .X(net1149));
 sg13g2_buf_2 fanout1150 (.A(net1151),
    .X(net1150));
 sg13g2_buf_4 fanout1151 (.X(net1151),
    .A(_3056_));
 sg13g2_buf_2 fanout1152 (.A(net1153),
    .X(net1152));
 sg13g2_buf_1 fanout1153 (.A(net1154),
    .X(net1153));
 sg13g2_buf_4 fanout1154 (.X(net1154),
    .A(_3056_));
 sg13g2_buf_2 fanout1155 (.A(net1156),
    .X(net1155));
 sg13g2_buf_2 fanout1156 (.A(net1157),
    .X(net1156));
 sg13g2_buf_2 fanout1157 (.A(net1158),
    .X(net1157));
 sg13g2_buf_4 fanout1158 (.X(net1158),
    .A(_1740_));
 sg13g2_buf_2 fanout1159 (.A(_0988_),
    .X(net1159));
 sg13g2_buf_4 fanout1160 (.X(net1160),
    .A(_0495_));
 sg13g2_buf_2 fanout1161 (.A(net1162),
    .X(net1161));
 sg13g2_buf_2 fanout1162 (.A(_3237_),
    .X(net1162));
 sg13g2_buf_4 fanout1163 (.X(net1163),
    .A(_3049_));
 sg13g2_buf_2 fanout1164 (.A(net1166),
    .X(net1164));
 sg13g2_buf_1 fanout1165 (.A(net1166),
    .X(net1165));
 sg13g2_buf_4 fanout1166 (.X(net1166),
    .A(net1169));
 sg13g2_buf_4 fanout1167 (.X(net1167),
    .A(net1169));
 sg13g2_buf_2 fanout1168 (.A(net1169),
    .X(net1168));
 sg13g2_buf_2 fanout1169 (.A(_2932_),
    .X(net1169));
 sg13g2_buf_2 fanout1170 (.A(net1171),
    .X(net1170));
 sg13g2_buf_4 fanout1171 (.X(net1171),
    .A(net1185));
 sg13g2_buf_2 fanout1172 (.A(net1173),
    .X(net1172));
 sg13g2_buf_2 fanout1173 (.A(net1185),
    .X(net1173));
 sg13g2_buf_4 fanout1174 (.X(net1174),
    .A(net1175));
 sg13g2_buf_2 fanout1175 (.A(net1185),
    .X(net1175));
 sg13g2_buf_4 fanout1176 (.X(net1176),
    .A(net1179));
 sg13g2_buf_2 fanout1177 (.A(net1179),
    .X(net1177));
 sg13g2_buf_2 fanout1178 (.A(net1179),
    .X(net1178));
 sg13g2_buf_2 fanout1179 (.A(net1185),
    .X(net1179));
 sg13g2_buf_2 fanout1180 (.A(net1181),
    .X(net1180));
 sg13g2_buf_2 fanout1181 (.A(net1184),
    .X(net1181));
 sg13g2_buf_2 fanout1182 (.A(net1184),
    .X(net1182));
 sg13g2_buf_2 fanout1183 (.A(net1184),
    .X(net1183));
 sg13g2_buf_2 fanout1184 (.A(net1185),
    .X(net1184));
 sg13g2_buf_4 fanout1185 (.X(net1185),
    .A(_2931_));
 sg13g2_buf_4 fanout1186 (.X(net1186),
    .A(_0766_));
 sg13g2_buf_4 fanout1187 (.X(net1187),
    .A(_3288_));
 sg13g2_buf_2 fanout1188 (.A(_3245_),
    .X(net1188));
 sg13g2_buf_4 fanout1189 (.X(net1189),
    .A(_3212_));
 sg13g2_buf_2 fanout1190 (.A(_3180_),
    .X(net1190));
 sg13g2_buf_4 fanout1191 (.X(net1191),
    .A(_3081_));
 sg13g2_buf_2 fanout1192 (.A(_3072_),
    .X(net1192));
 sg13g2_buf_4 fanout1193 (.X(net1193),
    .A(_3046_));
 sg13g2_buf_4 fanout1194 (.X(net1194),
    .A(_2884_));
 sg13g2_buf_4 fanout1195 (.X(net1195),
    .A(_2883_));
 sg13g2_buf_4 fanout1196 (.X(net1196),
    .A(_2882_));
 sg13g2_buf_2 fanout1197 (.A(_2882_),
    .X(net1197));
 sg13g2_buf_4 fanout1198 (.X(net1198),
    .A(_2881_));
 sg13g2_buf_2 fanout1199 (.A(_2881_),
    .X(net1199));
 sg13g2_buf_2 fanout1200 (.A(net1201),
    .X(net1200));
 sg13g2_buf_2 fanout1201 (.A(_2880_),
    .X(net1201));
 sg13g2_buf_4 fanout1202 (.X(net1202),
    .A(_2876_));
 sg13g2_buf_2 fanout1203 (.A(_2876_),
    .X(net1203));
 sg13g2_buf_2 fanout1204 (.A(net1211),
    .X(net1204));
 sg13g2_buf_2 fanout1205 (.A(net1207),
    .X(net1205));
 sg13g2_buf_1 fanout1206 (.A(net1207),
    .X(net1206));
 sg13g2_buf_2 fanout1207 (.A(net1208),
    .X(net1207));
 sg13g2_buf_2 fanout1208 (.A(net1211),
    .X(net1208));
 sg13g2_buf_2 fanout1209 (.A(net1210),
    .X(net1209));
 sg13g2_buf_2 fanout1210 (.A(net1211),
    .X(net1210));
 sg13g2_buf_2 fanout1211 (.A(_2874_),
    .X(net1211));
 sg13g2_buf_4 fanout1212 (.X(net1212),
    .A(_2850_));
 sg13g2_buf_4 fanout1213 (.X(net1213),
    .A(net1214));
 sg13g2_buf_4 fanout1214 (.X(net1214),
    .A(_2849_));
 sg13g2_buf_4 fanout1215 (.X(net1215),
    .A(net1216));
 sg13g2_buf_4 fanout1216 (.X(net1216),
    .A(net1217));
 sg13g2_buf_2 fanout1217 (.A(_2848_),
    .X(net1217));
 sg13g2_buf_4 fanout1218 (.X(net1218),
    .A(net1220));
 sg13g2_buf_1 fanout1219 (.A(net1220),
    .X(net1219));
 sg13g2_buf_2 fanout1220 (.A(net1221),
    .X(net1220));
 sg13g2_buf_2 fanout1221 (.A(_2847_),
    .X(net1221));
 sg13g2_buf_4 fanout1222 (.X(net1222),
    .A(_2846_));
 sg13g2_buf_4 fanout1223 (.X(net1223),
    .A(_2845_));
 sg13g2_buf_4 fanout1224 (.X(net1224),
    .A(_2843_));
 sg13g2_buf_4 fanout1225 (.X(net1225),
    .A(_2841_));
 sg13g2_buf_2 fanout1226 (.A(net1227),
    .X(net1226));
 sg13g2_buf_4 fanout1227 (.X(net1227),
    .A(_2822_));
 sg13g2_buf_4 fanout1228 (.X(net1228),
    .A(_2821_));
 sg13g2_buf_2 fanout1229 (.A(\movement_dir[1] ),
    .X(net1229));
 sg13g2_buf_2 fanout1230 (.A(\movement_dir[1] ),
    .X(net1230));
 sg13g2_buf_4 fanout1231 (.X(net1231),
    .A(net412));
 sg13g2_buf_2 fanout1232 (.A(\group_x[9] ),
    .X(net1232));
 sg13g2_buf_4 fanout1233 (.X(net1233),
    .A(\group_x[8] ));
 sg13g2_buf_4 fanout1234 (.X(net1234),
    .A(\group_x[7] ));
 sg13g2_buf_2 fanout1235 (.A(net1236),
    .X(net1235));
 sg13g2_buf_4 fanout1236 (.X(net1236),
    .A(_0057_));
 sg13g2_buf_2 fanout1237 (.A(net1238),
    .X(net1237));
 sg13g2_buf_4 fanout1238 (.X(net1238),
    .A(\group_x[6] ));
 sg13g2_buf_4 fanout1239 (.X(net1239),
    .A(net1241));
 sg13g2_buf_4 fanout1240 (.X(net1240),
    .A(net1241));
 sg13g2_buf_2 fanout1241 (.A(\group_x[5] ),
    .X(net1241));
 sg13g2_buf_2 fanout1242 (.A(net1244),
    .X(net1242));
 sg13g2_buf_1 fanout1243 (.A(net1244),
    .X(net1243));
 sg13g2_buf_2 fanout1244 (.A(net1245),
    .X(net1244));
 sg13g2_buf_4 fanout1245 (.X(net1245),
    .A(\group_x[4] ));
 sg13g2_buf_2 fanout1246 (.A(net1247),
    .X(net1246));
 sg13g2_buf_2 fanout1247 (.A(net1248),
    .X(net1247));
 sg13g2_buf_4 fanout1248 (.X(net1248),
    .A(net397));
 sg13g2_buf_4 fanout1249 (.X(net1249),
    .A(net1251));
 sg13g2_buf_4 fanout1250 (.X(net1250),
    .A(net1251));
 sg13g2_buf_4 fanout1251 (.X(net1251),
    .A(\group_x[2] ));
 sg13g2_buf_4 fanout1252 (.X(net1252),
    .A(\group_x[1] ));
 sg13g2_buf_2 fanout1253 (.A(\group_x[1] ),
    .X(net1253));
 sg13g2_buf_2 fanout1254 (.A(net402),
    .X(net1254));
 sg13g2_buf_2 fanout1255 (.A(net408),
    .X(net1255));
 sg13g2_buf_4 fanout1256 (.X(net1256),
    .A(net371));
 sg13g2_buf_4 fanout1257 (.X(net1257),
    .A(net407));
 sg13g2_buf_2 fanout1258 (.A(\myShooter.shooter_left_x[6] ),
    .X(net1258));
 sg13g2_buf_2 fanout1259 (.A(net1260),
    .X(net1259));
 sg13g2_buf_4 fanout1260 (.X(net1260),
    .A(net366));
 sg13g2_buf_4 fanout1261 (.X(net1261),
    .A(\myShooter.shooter_left_x[3] ));
 sg13g2_buf_2 fanout1262 (.A(net389),
    .X(net1262));
 sg13g2_buf_4 fanout1263 (.X(net1263),
    .A(net379));
 sg13g2_buf_4 fanout1264 (.X(net1264),
    .A(\barrier1.pix_y[9] ));
 sg13g2_buf_2 fanout1265 (.A(\barrier1.pix_y[9] ),
    .X(net1265));
 sg13g2_buf_4 fanout1266 (.X(net1266),
    .A(net1267));
 sg13g2_buf_2 fanout1267 (.A(_0016_),
    .X(net1267));
 sg13g2_buf_2 fanout1268 (.A(net1269),
    .X(net1268));
 sg13g2_buf_2 fanout1269 (.A(net1270),
    .X(net1269));
 sg13g2_buf_4 fanout1270 (.X(net1270),
    .A(net344));
 sg13g2_buf_4 fanout1271 (.X(net1271),
    .A(net1272));
 sg13g2_buf_4 fanout1272 (.X(net1272),
    .A(\barrier1.pix_y[7] ));
 sg13g2_buf_4 fanout1273 (.X(net1273),
    .A(net1274));
 sg13g2_buf_2 fanout1274 (.A(net1275),
    .X(net1274));
 sg13g2_buf_4 fanout1275 (.X(net1275),
    .A(net356));
 sg13g2_buf_4 fanout1276 (.X(net1276),
    .A(net1277));
 sg13g2_buf_4 fanout1277 (.X(net1277),
    .A(net337));
 sg13g2_buf_4 fanout1278 (.X(net1278),
    .A(net409));
 sg13g2_buf_2 fanout1279 (.A(_0012_),
    .X(net1279));
 sg13g2_buf_4 fanout1280 (.X(net1280),
    .A(net1281));
 sg13g2_buf_4 fanout1281 (.X(net1281),
    .A(net350));
 sg13g2_buf_2 fanout1282 (.A(net1284),
    .X(net1282));
 sg13g2_buf_4 fanout1283 (.X(net1283),
    .A(net1284));
 sg13g2_buf_2 fanout1284 (.A(_0011_),
    .X(net1284));
 sg13g2_buf_2 fanout1285 (.A(net1288),
    .X(net1285));
 sg13g2_buf_2 fanout1286 (.A(net1287),
    .X(net1286));
 sg13g2_buf_2 fanout1287 (.A(net1288),
    .X(net1287));
 sg13g2_buf_2 fanout1288 (.A(net1289),
    .X(net1288));
 sg13g2_buf_4 fanout1289 (.X(net1289),
    .A(net369));
 sg13g2_buf_2 fanout1290 (.A(net1291),
    .X(net1290));
 sg13g2_buf_1 fanout1291 (.A(net1292),
    .X(net1291));
 sg13g2_buf_2 fanout1292 (.A(net1293),
    .X(net1292));
 sg13g2_buf_2 fanout1293 (.A(net1294),
    .X(net1293));
 sg13g2_buf_4 fanout1294 (.X(net1294),
    .A(net358));
 sg13g2_buf_4 fanout1295 (.X(net1295),
    .A(net1298));
 sg13g2_buf_2 fanout1296 (.A(net1298),
    .X(net1296));
 sg13g2_buf_2 fanout1297 (.A(net1298),
    .X(net1297));
 sg13g2_buf_1 fanout1298 (.A(\barrier1.bar_rom.row_index[1] ),
    .X(net1298));
 sg13g2_buf_2 fanout1299 (.A(net382),
    .X(net1299));
 sg13g2_buf_2 fanout1300 (.A(\barrier1.bar_rom.row_index[0] ),
    .X(net1300));
 sg13g2_buf_2 fanout1301 (.A(net1302),
    .X(net1301));
 sg13g2_buf_2 fanout1302 (.A(move_dir),
    .X(net1302));
 sg13g2_buf_2 fanout1303 (.A(net391),
    .X(net1303));
 sg13g2_buf_1 fanout1304 (.A(\draw_score_inst.score[9] ),
    .X(net1304));
 sg13g2_buf_2 fanout1305 (.A(net395),
    .X(net1305));
 sg13g2_buf_2 fanout1306 (.A(\draw_score_inst.score[7] ),
    .X(net1306));
 sg13g2_buf_1 fanout1307 (.A(net357),
    .X(net1307));
 sg13g2_buf_2 fanout1308 (.A(\draw_score_inst.score[6] ),
    .X(net1308));
 sg13g2_buf_2 fanout1309 (.A(net381),
    .X(net1309));
 sg13g2_buf_2 fanout1310 (.A(\colRand[2] ),
    .X(net1310));
 sg13g2_buf_4 fanout1311 (.X(net1311),
    .A(net308));
 sg13g2_buf_1 fanout1312 (.A(\colRand[1] ),
    .X(net1312));
 sg13g2_buf_4 fanout1313 (.X(net1313),
    .A(net266));
 sg13g2_buf_2 fanout1314 (.A(net403),
    .X(net1314));
 sg13g2_buf_2 fanout1315 (.A(net404),
    .X(net1315));
 sg13g2_buf_2 fanout1316 (.A(\abullet_x[4] ),
    .X(net1316));
 sg13g2_buf_4 fanout1317 (.X(net1317),
    .A(\abullet_x[2] ));
 sg13g2_buf_2 fanout1318 (.A(net1319),
    .X(net1318));
 sg13g2_buf_2 fanout1319 (.A(net1320),
    .X(net1319));
 sg13g2_buf_2 fanout1320 (.A(abullet_active),
    .X(net1320));
 sg13g2_buf_2 fanout1321 (.A(\pb_y[8] ),
    .X(net1321));
 sg13g2_buf_2 fanout1322 (.A(\pb_y[6] ),
    .X(net1322));
 sg13g2_buf_2 fanout1323 (.A(\pb_y[5] ),
    .X(net1323));
 sg13g2_buf_2 fanout1324 (.A(\pb_y[3] ),
    .X(net1324));
 sg13g2_buf_2 fanout1325 (.A(\pb_y[2] ),
    .X(net1325));
 sg13g2_buf_2 fanout1326 (.A(\pb_y[1] ),
    .X(net1326));
 sg13g2_buf_4 fanout1327 (.X(net1327),
    .A(pb_active));
 sg13g2_buf_4 fanout1328 (.X(net1328),
    .A(net1329));
 sg13g2_buf_2 fanout1329 (.A(net1330),
    .X(net1329));
 sg13g2_buf_4 fanout1330 (.X(net1330),
    .A(net398));
 sg13g2_buf_4 fanout1331 (.X(net1331),
    .A(_0059_));
 sg13g2_buf_4 fanout1332 (.X(net1332),
    .A(\pb_x[8] ));
 sg13g2_buf_4 fanout1333 (.X(net1333),
    .A(\pb_x[8] ));
 sg13g2_buf_2 fanout1334 (.A(net1336),
    .X(net1334));
 sg13g2_buf_2 fanout1335 (.A(net1336),
    .X(net1335));
 sg13g2_buf_2 fanout1336 (.A(\pb_x[7] ),
    .X(net1336));
 sg13g2_buf_4 fanout1337 (.X(net1337),
    .A(_0065_));
 sg13g2_buf_4 fanout1338 (.X(net1338),
    .A(\pb_x[6] ));
 sg13g2_buf_2 fanout1339 (.A(\pb_x[6] ),
    .X(net1339));
 sg13g2_buf_2 fanout1340 (.A(net1341),
    .X(net1340));
 sg13g2_buf_2 fanout1341 (.A(net1342),
    .X(net1341));
 sg13g2_buf_2 fanout1342 (.A(_0066_),
    .X(net1342));
 sg13g2_buf_4 fanout1343 (.X(net1343),
    .A(\pb_x[5] ));
 sg13g2_buf_4 fanout1344 (.X(net1344),
    .A(net394));
 sg13g2_buf_2 fanout1345 (.A(\pb_x[4] ),
    .X(net1345));
 sg13g2_buf_2 fanout1346 (.A(\pb_x[3] ),
    .X(net1346));
 sg13g2_buf_2 fanout1347 (.A(\pb_x[3] ),
    .X(net1347));
 sg13g2_buf_2 fanout1348 (.A(net390),
    .X(net1348));
 sg13g2_buf_2 fanout1349 (.A(\pb_x[2] ),
    .X(net1349));
 sg13g2_buf_2 fanout1350 (.A(\pb_x[1] ),
    .X(net1350));
 sg13g2_buf_2 fanout1351 (.A(\pb_x[0] ),
    .X(net1351));
 sg13g2_buf_4 fanout1352 (.X(net1352),
    .A(_0008_));
 sg13g2_buf_4 fanout1353 (.X(net1353),
    .A(net1354));
 sg13g2_buf_4 fanout1354 (.X(net1354),
    .A(\barrier1.pix_x[9] ));
 sg13g2_buf_4 fanout1355 (.X(net1355),
    .A(net1356));
 sg13g2_buf_4 fanout1356 (.X(net1356),
    .A(_0038_));
 sg13g2_buf_4 fanout1357 (.X(net1357),
    .A(net1358));
 sg13g2_buf_2 fanout1358 (.A(net1359),
    .X(net1358));
 sg13g2_buf_4 fanout1359 (.X(net1359),
    .A(\barrier1.pix_x[8] ));
 sg13g2_buf_4 fanout1360 (.X(net1360),
    .A(_0036_));
 sg13g2_buf_4 fanout1361 (.X(net1361),
    .A(_0036_));
 sg13g2_buf_2 fanout1362 (.A(net1363),
    .X(net1362));
 sg13g2_buf_4 fanout1363 (.X(net1363),
    .A(net385));
 sg13g2_buf_4 fanout1364 (.X(net1364),
    .A(net1365));
 sg13g2_buf_2 fanout1365 (.A(\barrier1.pix_x[7] ),
    .X(net1365));
 sg13g2_buf_4 fanout1366 (.X(net1366),
    .A(net1367));
 sg13g2_buf_2 fanout1367 (.A(net1368),
    .X(net1367));
 sg13g2_buf_4 fanout1368 (.X(net1368),
    .A(_0027_));
 sg13g2_buf_2 fanout1369 (.A(net1370),
    .X(net1369));
 sg13g2_buf_2 fanout1370 (.A(net1372),
    .X(net1370));
 sg13g2_buf_4 fanout1371 (.X(net1371),
    .A(net1372));
 sg13g2_buf_2 fanout1372 (.A(\barrier1.pix_x[6] ),
    .X(net1372));
 sg13g2_buf_4 fanout1373 (.X(net1373),
    .A(net1374));
 sg13g2_buf_4 fanout1374 (.X(net1374),
    .A(_0028_));
 sg13g2_buf_2 fanout1375 (.A(net1376),
    .X(net1375));
 sg13g2_buf_2 fanout1376 (.A(net1377),
    .X(net1376));
 sg13g2_buf_4 fanout1377 (.X(net1377),
    .A(\barrier1.pix_x[5] ));
 sg13g2_buf_4 fanout1378 (.X(net1378),
    .A(_0029_));
 sg13g2_buf_4 fanout1379 (.X(net1379),
    .A(_0029_));
 sg13g2_buf_4 fanout1380 (.X(net1380),
    .A(net1383));
 sg13g2_buf_2 fanout1381 (.A(net1383),
    .X(net1381));
 sg13g2_buf_4 fanout1382 (.X(net1382),
    .A(net1383));
 sg13g2_buf_2 fanout1383 (.A(\barrier1.pix_x[4] ),
    .X(net1383));
 sg13g2_buf_4 fanout1384 (.X(net1384),
    .A(net1386));
 sg13g2_buf_2 fanout1385 (.A(net1386),
    .X(net1385));
 sg13g2_buf_2 fanout1386 (.A(net387),
    .X(net1386));
 sg13g2_buf_4 fanout1387 (.X(net1387),
    .A(\barrier1.pix_x[3] ));
 sg13g2_buf_2 fanout1388 (.A(net1389),
    .X(net1388));
 sg13g2_buf_2 fanout1389 (.A(net1390),
    .X(net1389));
 sg13g2_buf_2 fanout1390 (.A(net1393),
    .X(net1390));
 sg13g2_buf_2 fanout1391 (.A(net1392),
    .X(net1391));
 sg13g2_buf_2 fanout1392 (.A(net1393),
    .X(net1392));
 sg13g2_buf_2 fanout1393 (.A(\barrier1.pix_x[2] ),
    .X(net1393));
 sg13g2_buf_2 fanout1394 (.A(net1395),
    .X(net1394));
 sg13g2_buf_4 fanout1395 (.X(net1395),
    .A(\barrier1.col_idx[1] ));
 sg13g2_buf_2 fanout1396 (.A(net410),
    .X(net1396));
 sg13g2_buf_2 fanout1397 (.A(net1398),
    .X(net1397));
 sg13g2_buf_2 fanout1398 (.A(net1399),
    .X(net1398));
 sg13g2_buf_2 fanout1399 (.A(net1402),
    .X(net1399));
 sg13g2_buf_2 fanout1400 (.A(net1402),
    .X(net1400));
 sg13g2_buf_1 fanout1401 (.A(net1402),
    .X(net1401));
 sg13g2_buf_2 fanout1402 (.A(net1406),
    .X(net1402));
 sg13g2_buf_2 fanout1403 (.A(net1404),
    .X(net1403));
 sg13g2_buf_1 fanout1404 (.A(net1405),
    .X(net1404));
 sg13g2_buf_1 fanout1405 (.A(net1406),
    .X(net1405));
 sg13g2_buf_1 fanout1406 (.A(net1407),
    .X(net1406));
 sg13g2_buf_2 fanout1407 (.A(\barrier1.col_idx[0] ),
    .X(net1407));
 sg13g2_buf_2 fanout1408 (.A(net1409),
    .X(net1408));
 sg13g2_buf_1 fanout1409 (.A(net1410),
    .X(net1409));
 sg13g2_buf_2 fanout1410 (.A(net1411),
    .X(net1410));
 sg13g2_buf_4 fanout1411 (.X(net1411),
    .A(\barrier1.col_idx[0] ));
 sg13g2_buf_2 fanout1412 (.A(net1413),
    .X(net1412));
 sg13g2_buf_2 fanout1413 (.A(net1414),
    .X(net1413));
 sg13g2_buf_2 fanout1414 (.A(net1415),
    .X(net1414));
 sg13g2_buf_2 fanout1415 (.A(_2878_),
    .X(net1415));
 sg13g2_buf_8 fanout1416 (.A(net1417),
    .X(net1416));
 sg13g2_buf_8 fanout1417 (.A(net1),
    .X(net1417));
 sg13g2_buf_4 input1 (.X(net1),
    .A(rst_n));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_tielo tt_um_space_invaders_game_5 (.L_LO(net5));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_25__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0080_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0095_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold3 (.A(\lgA2.rx[0] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0055_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0199_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0009_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0110_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0052_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0205_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold10 (.A(\aliens_alive[8] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold11 (.A(_2554_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0007_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0219_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0079_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold15 (.A(\draw_score_inst.score[6] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold16 (.A(\lfsr[2] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0134_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold18 (.A(\sync_gen.vsync ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0232_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold20 (.A(\myShooter.shooter_left_x[1] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold21 (.A(\aliens_alive[20] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold22 (.A(\aliens_alive[2] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0053_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold24 (.A(_2615_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold25 (.A(\aliens_alive[25] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold26 (.A(\aliens_alive[7] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold27 (.A(\aliens_alive[26] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold28 (.A(\selectedRowRand[1] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0140_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold30 (.A(\aliens_alive[5] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold31 (.A(\lfsr[1] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0132_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold33 (.A(\aliens_alive[9] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold34 (.A(\barrier_health[0][2] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0198_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold36 (.A(game_over),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold37 (.A(_2930_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold38 (.A(\aliens_alive[10] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold39 (.A(\aliens_alive[17] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold40 (.A(\aliens_alive[13] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold41 (.A(\draw_score_inst.digit_health[0] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold42 (.A(_2544_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0154_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold44 (.A(\lfsr[4] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0135_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0056_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0196_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold48 (.A(\aliens_alive[29] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold49 (.A(\colRand[0] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold50 (.A(\aliens_alive[1] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold51 (.A(\aliens_alive[22] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold52 (.A(\aliens_alive[28] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold53 (.A(\aliens_alive[18] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold54 (.A(\aliens_alive[27] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold55 (.A(\aliens_alive[4] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold56 (.A(\lfsr[6] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0144_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold58 (.A(\aliens_alive[16] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold59 (.A(\aliens_alive[32] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold60 (.A(\aliens_alive[6] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold61 (.A(\aliens_alive[35] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold62 (.A(\lfsr[5] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold63 (.A(\aliens_alive[3] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold64 (.A(\lA2_x[1] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0253_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold66 (.A(\aliens_alive[12] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold67 (.A(\abullet_x[2] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0123_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold69 (.A(\aliens_alive[34] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold70 (.A(\aliens_alive[38] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold71 (.A(\abullet_x[4] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold72 (.A(\aliens_alive[31] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold73 (.A(\aliens_alive[21] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold74 (.A(\aliens_alive[30] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold75 (.A(\aliens_alive[11] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0046_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold77 (.A(_1747_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0102_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold79 (.A(\aliens_alive[0] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold80 (.A(\pb_x[0] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold81 (.A(\aliens_alive[15] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold82 (.A(\aliens_alive[14] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold83 (.A(\aliens_alive[33] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold84 (.A(\aliens_alive[36] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold85 (.A(\lfsr[7] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold86 (.A(\aliens_alive[37] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold87 (.A(\myShooter.shooter_left_x[6] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold88 (.A(\selectedRowRand[0] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0139_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold90 (.A(\aliens_alive[23] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold91 (.A(\colRand[1] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold92 (.A(\aliens_alive[39] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold93 (.A(\aliens_alive[24] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold94 (.A(\draw_score_inst.digit_health[1] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold95 (.A(\pb_y[7] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold96 (.A(\selectedRowRand[2] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0141_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold98 (.A(\barrier_health[0][1] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold99 (.A(_2593_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0197_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold101 (.A(\aliens_alive[19] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0067_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0124_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold104 (.A(\pb_y[9] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0119_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold106 (.A(\pb_y[4] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold107 (.A(_2300_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0062_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold109 (.A(_2739_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold110 (.A(_2740_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold111 (.A(prev_button1),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold112 (.A(_2923_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold113 (.A(\abullet_x[1] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold114 (.A(\abullet_y[5] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0246_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0049_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0250_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold118 (.A(\draw_score_inst.score[2] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0146_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold120 (.A(\barrier1.pix_y[5] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0064_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0244_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold123 (.A(\abullet_y[7] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0017_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold125 (.A(\draw_score_inst.score[4] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0148_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold127 (.A(\barrier1.pix_y[8] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold128 (.A(\lfsr[0] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold129 (.A(\abullet_y[8] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold130 (.A(_2769_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold131 (.A(\barrier_health[3][1] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0206_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold133 (.A(\barrier1.pix_y[4] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold134 (.A(prev_button0),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold135 (.A(_2921_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold136 (.A(\barrier_health[1][1] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0200_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold138 (.A(\myShooter.shooter_left_x[9] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold139 (.A(\barrier1.pix_y[6] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold140 (.A(\draw_score_inst.score[7] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold141 (.A(\barrier1.bar_rom.row_index[2] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0072_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold143 (.A(_2302_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold144 (.A(\barrier_health[2][1] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0203_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold146 (.A(\barrier_health[2][2] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold147 (.A(\barrier_health[3][2] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold148 (.A(\abullet_x[5] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold149 (.A(\myShooter.shooter_left_x[4] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold150 (.A(\abullet_x[8] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold151 (.A(move_dir),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold152 (.A(\barrier1.bar_rom.row_index[3] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold153 (.A(_2661_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold154 (.A(\myShooter.shooter_left_x[8] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0051_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold156 (.A(_2750_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0245_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold158 (.A(\abullet_x[0] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0121_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0043_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0105_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold162 (.A(\myShooter.shooter_left_x[2] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold163 (.A(\abullet_x[6] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold164 (.A(\draw_score_inst.score[5] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold165 (.A(\barrier1.bar_rom.row_index[0] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0025_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0145_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold168 (.A(\barrier1.pix_x[7] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold169 (.A(_3093_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold170 (.A(\barrier1.pix_x[3] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold171 (.A(_3084_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold172 (.A(\myShooter.shooter_left_x[3] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold173 (.A(\pb_x[2] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold174 (.A(\draw_score_inst.score[9] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold175 (.A(\barrier_health[1][2] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold176 (.A(\pb_y[0] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold177 (.A(\pb_x[4] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold178 (.A(\draw_score_inst.score[8] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold179 (.A(\myShooter.shooter_left_x[5] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold180 (.A(\group_x[3] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold181 (.A(\pb_x[9] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold182 (.A(\draw_score_inst.score[3] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold183 (.A(_2925_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold184 (.A(\pb_y[5] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold185 (.A(\abullet_y[6] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold186 (.A(\abullet_x[9] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold187 (.A(\abullet_x[7] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0015_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0037_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold190 (.A(\myShooter.shooter_left_x[7] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold191 (.A(\abullet_y[2] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0012_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold193 (.A(\barrier1.col_idx[1] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold194 (.A(_3066_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold195 (.A(\group_x[9] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold196 (.A(pb_active),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0013_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold198 (.A(\pb_y[0] ),
    .X(net415));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_decap_8 FILLER_13_588 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_decap_8 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_637 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_8 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_decap_8 FILLER_13_798 ();
 sg13g2_decap_8 FILLER_13_805 ();
 sg13g2_decap_8 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_833 ();
 sg13g2_decap_8 FILLER_13_840 ();
 sg13g2_decap_8 FILLER_13_847 ();
 sg13g2_decap_8 FILLER_13_854 ();
 sg13g2_fill_1 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_8 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_511 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_574 ();
 sg13g2_decap_8 FILLER_14_581 ();
 sg13g2_decap_8 FILLER_14_588 ();
 sg13g2_decap_8 FILLER_14_595 ();
 sg13g2_decap_8 FILLER_14_602 ();
 sg13g2_decap_8 FILLER_14_609 ();
 sg13g2_decap_8 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_623 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_decap_8 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_decap_8 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_658 ();
 sg13g2_decap_8 FILLER_14_665 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_decap_8 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_decap_8 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_14_840 ();
 sg13g2_decap_8 FILLER_14_847 ();
 sg13g2_decap_8 FILLER_14_854 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_434 ();
 sg13g2_decap_8 FILLER_15_441 ();
 sg13g2_decap_8 FILLER_15_448 ();
 sg13g2_decap_8 FILLER_15_455 ();
 sg13g2_decap_8 FILLER_15_462 ();
 sg13g2_decap_8 FILLER_15_469 ();
 sg13g2_decap_8 FILLER_15_476 ();
 sg13g2_decap_8 FILLER_15_483 ();
 sg13g2_decap_8 FILLER_15_490 ();
 sg13g2_decap_8 FILLER_15_497 ();
 sg13g2_decap_8 FILLER_15_504 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_518 ();
 sg13g2_decap_8 FILLER_15_525 ();
 sg13g2_decap_8 FILLER_15_532 ();
 sg13g2_decap_8 FILLER_15_539 ();
 sg13g2_decap_8 FILLER_15_546 ();
 sg13g2_decap_8 FILLER_15_553 ();
 sg13g2_decap_8 FILLER_15_560 ();
 sg13g2_decap_8 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_574 ();
 sg13g2_decap_8 FILLER_15_581 ();
 sg13g2_decap_8 FILLER_15_588 ();
 sg13g2_decap_8 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_602 ();
 sg13g2_decap_8 FILLER_15_609 ();
 sg13g2_decap_8 FILLER_15_616 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_8 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_644 ();
 sg13g2_decap_8 FILLER_15_651 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_decap_8 FILLER_15_665 ();
 sg13g2_decap_8 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_679 ();
 sg13g2_decap_8 FILLER_15_686 ();
 sg13g2_decap_8 FILLER_15_693 ();
 sg13g2_decap_8 FILLER_15_700 ();
 sg13g2_decap_8 FILLER_15_707 ();
 sg13g2_decap_8 FILLER_15_714 ();
 sg13g2_decap_8 FILLER_15_721 ();
 sg13g2_decap_8 FILLER_15_728 ();
 sg13g2_decap_8 FILLER_15_735 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_decap_8 FILLER_15_749 ();
 sg13g2_decap_8 FILLER_15_756 ();
 sg13g2_decap_8 FILLER_15_763 ();
 sg13g2_decap_8 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_777 ();
 sg13g2_decap_8 FILLER_15_784 ();
 sg13g2_decap_8 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_798 ();
 sg13g2_decap_8 FILLER_15_805 ();
 sg13g2_decap_8 FILLER_15_812 ();
 sg13g2_decap_8 FILLER_15_819 ();
 sg13g2_decap_8 FILLER_15_826 ();
 sg13g2_decap_8 FILLER_15_833 ();
 sg13g2_decap_8 FILLER_15_840 ();
 sg13g2_decap_8 FILLER_15_847 ();
 sg13g2_decap_8 FILLER_15_854 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_8 FILLER_16_455 ();
 sg13g2_decap_8 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_469 ();
 sg13g2_decap_8 FILLER_16_476 ();
 sg13g2_decap_8 FILLER_16_483 ();
 sg13g2_decap_8 FILLER_16_490 ();
 sg13g2_decap_8 FILLER_16_497 ();
 sg13g2_decap_8 FILLER_16_504 ();
 sg13g2_decap_8 FILLER_16_511 ();
 sg13g2_decap_8 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_525 ();
 sg13g2_decap_8 FILLER_16_532 ();
 sg13g2_decap_8 FILLER_16_539 ();
 sg13g2_decap_8 FILLER_16_546 ();
 sg13g2_decap_8 FILLER_16_553 ();
 sg13g2_decap_8 FILLER_16_560 ();
 sg13g2_decap_8 FILLER_16_567 ();
 sg13g2_decap_8 FILLER_16_574 ();
 sg13g2_decap_8 FILLER_16_581 ();
 sg13g2_decap_8 FILLER_16_588 ();
 sg13g2_decap_8 FILLER_16_595 ();
 sg13g2_decap_8 FILLER_16_602 ();
 sg13g2_decap_8 FILLER_16_609 ();
 sg13g2_decap_8 FILLER_16_616 ();
 sg13g2_decap_8 FILLER_16_623 ();
 sg13g2_decap_8 FILLER_16_630 ();
 sg13g2_decap_8 FILLER_16_637 ();
 sg13g2_decap_8 FILLER_16_644 ();
 sg13g2_decap_8 FILLER_16_651 ();
 sg13g2_decap_8 FILLER_16_658 ();
 sg13g2_decap_8 FILLER_16_665 ();
 sg13g2_decap_8 FILLER_16_672 ();
 sg13g2_decap_8 FILLER_16_679 ();
 sg13g2_decap_8 FILLER_16_686 ();
 sg13g2_decap_8 FILLER_16_693 ();
 sg13g2_decap_8 FILLER_16_700 ();
 sg13g2_decap_8 FILLER_16_707 ();
 sg13g2_decap_8 FILLER_16_714 ();
 sg13g2_decap_8 FILLER_16_721 ();
 sg13g2_decap_8 FILLER_16_728 ();
 sg13g2_decap_8 FILLER_16_735 ();
 sg13g2_decap_8 FILLER_16_742 ();
 sg13g2_decap_8 FILLER_16_749 ();
 sg13g2_decap_8 FILLER_16_756 ();
 sg13g2_decap_8 FILLER_16_763 ();
 sg13g2_decap_8 FILLER_16_770 ();
 sg13g2_decap_8 FILLER_16_777 ();
 sg13g2_decap_8 FILLER_16_784 ();
 sg13g2_decap_8 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_798 ();
 sg13g2_decap_8 FILLER_16_805 ();
 sg13g2_decap_8 FILLER_16_812 ();
 sg13g2_decap_8 FILLER_16_819 ();
 sg13g2_decap_8 FILLER_16_826 ();
 sg13g2_decap_8 FILLER_16_833 ();
 sg13g2_decap_8 FILLER_16_840 ();
 sg13g2_decap_8 FILLER_16_847 ();
 sg13g2_decap_8 FILLER_16_854 ();
 sg13g2_fill_1 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_427 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_448 ();
 sg13g2_decap_8 FILLER_17_455 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_497 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_fill_1 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_decap_8 FILLER_18_427 ();
 sg13g2_decap_8 FILLER_18_434 ();
 sg13g2_decap_8 FILLER_18_441 ();
 sg13g2_decap_8 FILLER_18_448 ();
 sg13g2_decap_8 FILLER_18_455 ();
 sg13g2_decap_8 FILLER_18_462 ();
 sg13g2_decap_8 FILLER_18_469 ();
 sg13g2_decap_8 FILLER_18_476 ();
 sg13g2_decap_8 FILLER_18_483 ();
 sg13g2_decap_8 FILLER_18_490 ();
 sg13g2_decap_8 FILLER_18_497 ();
 sg13g2_decap_8 FILLER_18_504 ();
 sg13g2_decap_8 FILLER_18_511 ();
 sg13g2_decap_8 FILLER_18_518 ();
 sg13g2_decap_8 FILLER_18_525 ();
 sg13g2_decap_8 FILLER_18_532 ();
 sg13g2_decap_8 FILLER_18_539 ();
 sg13g2_decap_8 FILLER_18_546 ();
 sg13g2_decap_8 FILLER_18_553 ();
 sg13g2_decap_8 FILLER_18_560 ();
 sg13g2_decap_8 FILLER_18_567 ();
 sg13g2_decap_8 FILLER_18_574 ();
 sg13g2_decap_8 FILLER_18_581 ();
 sg13g2_decap_8 FILLER_18_588 ();
 sg13g2_decap_8 FILLER_18_595 ();
 sg13g2_decap_8 FILLER_18_602 ();
 sg13g2_decap_8 FILLER_18_609 ();
 sg13g2_decap_8 FILLER_18_616 ();
 sg13g2_decap_8 FILLER_18_623 ();
 sg13g2_decap_8 FILLER_18_630 ();
 sg13g2_decap_8 FILLER_18_637 ();
 sg13g2_decap_8 FILLER_18_644 ();
 sg13g2_decap_8 FILLER_18_651 ();
 sg13g2_decap_8 FILLER_18_658 ();
 sg13g2_decap_8 FILLER_18_665 ();
 sg13g2_decap_8 FILLER_18_672 ();
 sg13g2_decap_8 FILLER_18_679 ();
 sg13g2_decap_8 FILLER_18_686 ();
 sg13g2_decap_8 FILLER_18_693 ();
 sg13g2_decap_8 FILLER_18_700 ();
 sg13g2_decap_8 FILLER_18_707 ();
 sg13g2_decap_8 FILLER_18_714 ();
 sg13g2_decap_8 FILLER_18_721 ();
 sg13g2_decap_8 FILLER_18_728 ();
 sg13g2_decap_8 FILLER_18_735 ();
 sg13g2_decap_8 FILLER_18_742 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_decap_8 FILLER_18_756 ();
 sg13g2_decap_8 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_770 ();
 sg13g2_decap_8 FILLER_18_777 ();
 sg13g2_decap_8 FILLER_18_784 ();
 sg13g2_decap_8 FILLER_18_791 ();
 sg13g2_decap_8 FILLER_18_798 ();
 sg13g2_decap_8 FILLER_18_805 ();
 sg13g2_decap_8 FILLER_18_812 ();
 sg13g2_decap_8 FILLER_18_819 ();
 sg13g2_decap_8 FILLER_18_826 ();
 sg13g2_decap_8 FILLER_18_833 ();
 sg13g2_decap_8 FILLER_18_840 ();
 sg13g2_decap_8 FILLER_18_847 ();
 sg13g2_decap_8 FILLER_18_854 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_decap_8 FILLER_19_427 ();
 sg13g2_decap_8 FILLER_19_434 ();
 sg13g2_decap_8 FILLER_19_441 ();
 sg13g2_decap_8 FILLER_19_448 ();
 sg13g2_decap_8 FILLER_19_455 ();
 sg13g2_decap_8 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_490 ();
 sg13g2_decap_8 FILLER_19_497 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_532 ();
 sg13g2_decap_8 FILLER_19_539 ();
 sg13g2_decap_8 FILLER_19_546 ();
 sg13g2_decap_8 FILLER_19_553 ();
 sg13g2_decap_8 FILLER_19_560 ();
 sg13g2_decap_8 FILLER_19_567 ();
 sg13g2_decap_8 FILLER_19_574 ();
 sg13g2_decap_8 FILLER_19_581 ();
 sg13g2_decap_8 FILLER_19_588 ();
 sg13g2_decap_8 FILLER_19_595 ();
 sg13g2_decap_8 FILLER_19_602 ();
 sg13g2_decap_8 FILLER_19_609 ();
 sg13g2_decap_8 FILLER_19_616 ();
 sg13g2_decap_8 FILLER_19_623 ();
 sg13g2_decap_8 FILLER_19_630 ();
 sg13g2_decap_8 FILLER_19_637 ();
 sg13g2_decap_8 FILLER_19_644 ();
 sg13g2_decap_8 FILLER_19_651 ();
 sg13g2_decap_8 FILLER_19_658 ();
 sg13g2_decap_8 FILLER_19_665 ();
 sg13g2_decap_8 FILLER_19_672 ();
 sg13g2_decap_8 FILLER_19_679 ();
 sg13g2_decap_8 FILLER_19_686 ();
 sg13g2_decap_8 FILLER_19_693 ();
 sg13g2_decap_8 FILLER_19_700 ();
 sg13g2_decap_8 FILLER_19_707 ();
 sg13g2_decap_8 FILLER_19_714 ();
 sg13g2_decap_8 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_784 ();
 sg13g2_decap_8 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_798 ();
 sg13g2_decap_8 FILLER_19_805 ();
 sg13g2_decap_8 FILLER_19_812 ();
 sg13g2_decap_8 FILLER_19_819 ();
 sg13g2_decap_8 FILLER_19_826 ();
 sg13g2_decap_8 FILLER_19_833 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_decap_8 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_854 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_decap_8 FILLER_20_427 ();
 sg13g2_decap_8 FILLER_20_434 ();
 sg13g2_decap_8 FILLER_20_441 ();
 sg13g2_decap_8 FILLER_20_448 ();
 sg13g2_decap_8 FILLER_20_455 ();
 sg13g2_decap_8 FILLER_20_462 ();
 sg13g2_decap_8 FILLER_20_469 ();
 sg13g2_decap_8 FILLER_20_476 ();
 sg13g2_decap_8 FILLER_20_483 ();
 sg13g2_decap_8 FILLER_20_490 ();
 sg13g2_decap_8 FILLER_20_497 ();
 sg13g2_decap_8 FILLER_20_504 ();
 sg13g2_decap_8 FILLER_20_511 ();
 sg13g2_decap_8 FILLER_20_518 ();
 sg13g2_decap_8 FILLER_20_525 ();
 sg13g2_decap_8 FILLER_20_532 ();
 sg13g2_decap_8 FILLER_20_539 ();
 sg13g2_decap_8 FILLER_20_546 ();
 sg13g2_decap_8 FILLER_20_553 ();
 sg13g2_decap_8 FILLER_20_560 ();
 sg13g2_decap_8 FILLER_20_567 ();
 sg13g2_decap_8 FILLER_20_574 ();
 sg13g2_decap_8 FILLER_20_581 ();
 sg13g2_decap_8 FILLER_20_588 ();
 sg13g2_decap_8 FILLER_20_595 ();
 sg13g2_decap_8 FILLER_20_602 ();
 sg13g2_decap_8 FILLER_20_609 ();
 sg13g2_decap_8 FILLER_20_616 ();
 sg13g2_decap_8 FILLER_20_623 ();
 sg13g2_decap_8 FILLER_20_630 ();
 sg13g2_decap_8 FILLER_20_637 ();
 sg13g2_decap_8 FILLER_20_644 ();
 sg13g2_decap_8 FILLER_20_651 ();
 sg13g2_decap_8 FILLER_20_658 ();
 sg13g2_decap_8 FILLER_20_665 ();
 sg13g2_decap_8 FILLER_20_672 ();
 sg13g2_decap_8 FILLER_20_679 ();
 sg13g2_decap_8 FILLER_20_686 ();
 sg13g2_decap_8 FILLER_20_693 ();
 sg13g2_decap_8 FILLER_20_700 ();
 sg13g2_decap_8 FILLER_20_707 ();
 sg13g2_decap_8 FILLER_20_714 ();
 sg13g2_decap_8 FILLER_20_721 ();
 sg13g2_decap_8 FILLER_20_728 ();
 sg13g2_decap_8 FILLER_20_735 ();
 sg13g2_decap_8 FILLER_20_742 ();
 sg13g2_decap_8 FILLER_20_749 ();
 sg13g2_decap_8 FILLER_20_756 ();
 sg13g2_decap_8 FILLER_20_763 ();
 sg13g2_decap_8 FILLER_20_770 ();
 sg13g2_decap_8 FILLER_20_777 ();
 sg13g2_decap_8 FILLER_20_784 ();
 sg13g2_decap_8 FILLER_20_791 ();
 sg13g2_decap_8 FILLER_20_798 ();
 sg13g2_decap_8 FILLER_20_805 ();
 sg13g2_decap_8 FILLER_20_812 ();
 sg13g2_decap_8 FILLER_20_819 ();
 sg13g2_decap_8 FILLER_20_826 ();
 sg13g2_decap_8 FILLER_20_833 ();
 sg13g2_decap_8 FILLER_20_840 ();
 sg13g2_decap_8 FILLER_20_847 ();
 sg13g2_decap_8 FILLER_20_854 ();
 sg13g2_fill_1 FILLER_20_861 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_decap_8 FILLER_21_427 ();
 sg13g2_decap_8 FILLER_21_434 ();
 sg13g2_decap_8 FILLER_21_441 ();
 sg13g2_decap_8 FILLER_21_448 ();
 sg13g2_decap_8 FILLER_21_455 ();
 sg13g2_decap_8 FILLER_21_462 ();
 sg13g2_decap_8 FILLER_21_469 ();
 sg13g2_decap_8 FILLER_21_476 ();
 sg13g2_decap_8 FILLER_21_483 ();
 sg13g2_decap_8 FILLER_21_490 ();
 sg13g2_decap_8 FILLER_21_497 ();
 sg13g2_decap_8 FILLER_21_504 ();
 sg13g2_decap_8 FILLER_21_511 ();
 sg13g2_decap_8 FILLER_21_518 ();
 sg13g2_decap_8 FILLER_21_525 ();
 sg13g2_decap_8 FILLER_21_532 ();
 sg13g2_decap_8 FILLER_21_539 ();
 sg13g2_decap_8 FILLER_21_546 ();
 sg13g2_decap_8 FILLER_21_553 ();
 sg13g2_decap_8 FILLER_21_560 ();
 sg13g2_decap_8 FILLER_21_567 ();
 sg13g2_decap_8 FILLER_21_574 ();
 sg13g2_decap_8 FILLER_21_581 ();
 sg13g2_decap_8 FILLER_21_588 ();
 sg13g2_decap_8 FILLER_21_595 ();
 sg13g2_decap_8 FILLER_21_602 ();
 sg13g2_decap_8 FILLER_21_609 ();
 sg13g2_decap_8 FILLER_21_616 ();
 sg13g2_decap_8 FILLER_21_623 ();
 sg13g2_decap_8 FILLER_21_630 ();
 sg13g2_decap_8 FILLER_21_637 ();
 sg13g2_decap_8 FILLER_21_644 ();
 sg13g2_decap_8 FILLER_21_651 ();
 sg13g2_decap_8 FILLER_21_658 ();
 sg13g2_decap_8 FILLER_21_665 ();
 sg13g2_decap_8 FILLER_21_672 ();
 sg13g2_decap_8 FILLER_21_679 ();
 sg13g2_decap_8 FILLER_21_686 ();
 sg13g2_decap_8 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_700 ();
 sg13g2_decap_8 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_714 ();
 sg13g2_decap_8 FILLER_21_721 ();
 sg13g2_decap_8 FILLER_21_728 ();
 sg13g2_decap_8 FILLER_21_735 ();
 sg13g2_decap_8 FILLER_21_742 ();
 sg13g2_decap_8 FILLER_21_749 ();
 sg13g2_decap_8 FILLER_21_756 ();
 sg13g2_decap_8 FILLER_21_763 ();
 sg13g2_decap_8 FILLER_21_770 ();
 sg13g2_decap_8 FILLER_21_777 ();
 sg13g2_decap_8 FILLER_21_784 ();
 sg13g2_decap_8 FILLER_21_791 ();
 sg13g2_decap_8 FILLER_21_798 ();
 sg13g2_decap_8 FILLER_21_805 ();
 sg13g2_decap_8 FILLER_21_812 ();
 sg13g2_decap_8 FILLER_21_819 ();
 sg13g2_decap_8 FILLER_21_826 ();
 sg13g2_decap_8 FILLER_21_833 ();
 sg13g2_decap_8 FILLER_21_840 ();
 sg13g2_decap_8 FILLER_21_847 ();
 sg13g2_decap_8 FILLER_21_854 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_22_406 ();
 sg13g2_decap_8 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_decap_8 FILLER_22_427 ();
 sg13g2_decap_8 FILLER_22_434 ();
 sg13g2_decap_8 FILLER_22_441 ();
 sg13g2_decap_8 FILLER_22_448 ();
 sg13g2_decap_8 FILLER_22_455 ();
 sg13g2_decap_8 FILLER_22_462 ();
 sg13g2_decap_8 FILLER_22_469 ();
 sg13g2_decap_8 FILLER_22_476 ();
 sg13g2_decap_8 FILLER_22_483 ();
 sg13g2_decap_8 FILLER_22_490 ();
 sg13g2_decap_8 FILLER_22_497 ();
 sg13g2_decap_8 FILLER_22_504 ();
 sg13g2_decap_8 FILLER_22_511 ();
 sg13g2_decap_8 FILLER_22_518 ();
 sg13g2_decap_8 FILLER_22_525 ();
 sg13g2_decap_8 FILLER_22_532 ();
 sg13g2_decap_8 FILLER_22_539 ();
 sg13g2_decap_8 FILLER_22_546 ();
 sg13g2_decap_8 FILLER_22_553 ();
 sg13g2_decap_8 FILLER_22_560 ();
 sg13g2_decap_8 FILLER_22_567 ();
 sg13g2_decap_8 FILLER_22_574 ();
 sg13g2_decap_8 FILLER_22_581 ();
 sg13g2_decap_8 FILLER_22_588 ();
 sg13g2_decap_8 FILLER_22_595 ();
 sg13g2_decap_8 FILLER_22_602 ();
 sg13g2_decap_8 FILLER_22_609 ();
 sg13g2_decap_8 FILLER_22_616 ();
 sg13g2_decap_8 FILLER_22_623 ();
 sg13g2_decap_8 FILLER_22_630 ();
 sg13g2_decap_8 FILLER_22_637 ();
 sg13g2_decap_8 FILLER_22_644 ();
 sg13g2_decap_8 FILLER_22_651 ();
 sg13g2_decap_8 FILLER_22_658 ();
 sg13g2_decap_8 FILLER_22_665 ();
 sg13g2_decap_8 FILLER_22_672 ();
 sg13g2_decap_8 FILLER_22_679 ();
 sg13g2_decap_8 FILLER_22_686 ();
 sg13g2_decap_8 FILLER_22_693 ();
 sg13g2_decap_8 FILLER_22_700 ();
 sg13g2_decap_8 FILLER_22_707 ();
 sg13g2_decap_8 FILLER_22_714 ();
 sg13g2_decap_8 FILLER_22_721 ();
 sg13g2_decap_8 FILLER_22_728 ();
 sg13g2_decap_8 FILLER_22_735 ();
 sg13g2_decap_8 FILLER_22_742 ();
 sg13g2_decap_8 FILLER_22_749 ();
 sg13g2_decap_8 FILLER_22_756 ();
 sg13g2_decap_8 FILLER_22_763 ();
 sg13g2_decap_8 FILLER_22_770 ();
 sg13g2_decap_8 FILLER_22_777 ();
 sg13g2_decap_8 FILLER_22_784 ();
 sg13g2_decap_8 FILLER_22_791 ();
 sg13g2_decap_8 FILLER_22_798 ();
 sg13g2_decap_8 FILLER_22_805 ();
 sg13g2_decap_8 FILLER_22_812 ();
 sg13g2_decap_8 FILLER_22_819 ();
 sg13g2_decap_8 FILLER_22_826 ();
 sg13g2_decap_8 FILLER_22_833 ();
 sg13g2_decap_8 FILLER_22_840 ();
 sg13g2_decap_8 FILLER_22_847 ();
 sg13g2_decap_8 FILLER_22_854 ();
 sg13g2_fill_1 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_decap_8 FILLER_23_406 ();
 sg13g2_decap_8 FILLER_23_413 ();
 sg13g2_decap_8 FILLER_23_420 ();
 sg13g2_decap_8 FILLER_23_427 ();
 sg13g2_decap_8 FILLER_23_434 ();
 sg13g2_decap_8 FILLER_23_441 ();
 sg13g2_decap_8 FILLER_23_448 ();
 sg13g2_decap_8 FILLER_23_455 ();
 sg13g2_decap_8 FILLER_23_462 ();
 sg13g2_decap_8 FILLER_23_469 ();
 sg13g2_decap_8 FILLER_23_476 ();
 sg13g2_decap_8 FILLER_23_483 ();
 sg13g2_decap_8 FILLER_23_490 ();
 sg13g2_decap_8 FILLER_23_497 ();
 sg13g2_decap_8 FILLER_23_504 ();
 sg13g2_decap_8 FILLER_23_511 ();
 sg13g2_decap_8 FILLER_23_518 ();
 sg13g2_decap_8 FILLER_23_525 ();
 sg13g2_decap_8 FILLER_23_532 ();
 sg13g2_decap_8 FILLER_23_539 ();
 sg13g2_decap_8 FILLER_23_546 ();
 sg13g2_decap_8 FILLER_23_553 ();
 sg13g2_decap_8 FILLER_23_560 ();
 sg13g2_decap_8 FILLER_23_567 ();
 sg13g2_decap_8 FILLER_23_574 ();
 sg13g2_decap_8 FILLER_23_581 ();
 sg13g2_decap_8 FILLER_23_588 ();
 sg13g2_decap_8 FILLER_23_595 ();
 sg13g2_decap_8 FILLER_23_602 ();
 sg13g2_decap_8 FILLER_23_609 ();
 sg13g2_decap_8 FILLER_23_616 ();
 sg13g2_decap_8 FILLER_23_623 ();
 sg13g2_decap_8 FILLER_23_630 ();
 sg13g2_decap_8 FILLER_23_637 ();
 sg13g2_decap_8 FILLER_23_644 ();
 sg13g2_decap_8 FILLER_23_651 ();
 sg13g2_decap_8 FILLER_23_658 ();
 sg13g2_decap_8 FILLER_23_665 ();
 sg13g2_decap_8 FILLER_23_672 ();
 sg13g2_decap_8 FILLER_23_679 ();
 sg13g2_decap_8 FILLER_23_686 ();
 sg13g2_decap_8 FILLER_23_693 ();
 sg13g2_decap_8 FILLER_23_700 ();
 sg13g2_decap_8 FILLER_23_707 ();
 sg13g2_decap_8 FILLER_23_714 ();
 sg13g2_decap_8 FILLER_23_721 ();
 sg13g2_decap_8 FILLER_23_728 ();
 sg13g2_decap_8 FILLER_23_735 ();
 sg13g2_decap_8 FILLER_23_742 ();
 sg13g2_decap_8 FILLER_23_749 ();
 sg13g2_decap_8 FILLER_23_756 ();
 sg13g2_decap_8 FILLER_23_763 ();
 sg13g2_decap_8 FILLER_23_770 ();
 sg13g2_decap_8 FILLER_23_777 ();
 sg13g2_decap_8 FILLER_23_784 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_798 ();
 sg13g2_decap_8 FILLER_23_805 ();
 sg13g2_decap_8 FILLER_23_812 ();
 sg13g2_decap_8 FILLER_23_819 ();
 sg13g2_decap_8 FILLER_23_826 ();
 sg13g2_decap_8 FILLER_23_833 ();
 sg13g2_decap_8 FILLER_23_840 ();
 sg13g2_decap_8 FILLER_23_847 ();
 sg13g2_decap_8 FILLER_23_854 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_decap_8 FILLER_24_406 ();
 sg13g2_decap_8 FILLER_24_413 ();
 sg13g2_decap_8 FILLER_24_420 ();
 sg13g2_decap_8 FILLER_24_427 ();
 sg13g2_decap_8 FILLER_24_434 ();
 sg13g2_decap_8 FILLER_24_441 ();
 sg13g2_decap_8 FILLER_24_448 ();
 sg13g2_decap_8 FILLER_24_455 ();
 sg13g2_decap_8 FILLER_24_462 ();
 sg13g2_decap_8 FILLER_24_469 ();
 sg13g2_decap_8 FILLER_24_476 ();
 sg13g2_decap_8 FILLER_24_483 ();
 sg13g2_decap_8 FILLER_24_490 ();
 sg13g2_decap_8 FILLER_24_497 ();
 sg13g2_decap_8 FILLER_24_504 ();
 sg13g2_decap_8 FILLER_24_511 ();
 sg13g2_decap_8 FILLER_24_518 ();
 sg13g2_decap_8 FILLER_24_525 ();
 sg13g2_decap_8 FILLER_24_532 ();
 sg13g2_decap_8 FILLER_24_539 ();
 sg13g2_decap_8 FILLER_24_546 ();
 sg13g2_decap_8 FILLER_24_553 ();
 sg13g2_decap_8 FILLER_24_560 ();
 sg13g2_decap_8 FILLER_24_567 ();
 sg13g2_decap_8 FILLER_24_574 ();
 sg13g2_decap_8 FILLER_24_581 ();
 sg13g2_decap_8 FILLER_24_588 ();
 sg13g2_decap_8 FILLER_24_595 ();
 sg13g2_decap_8 FILLER_24_602 ();
 sg13g2_decap_8 FILLER_24_609 ();
 sg13g2_decap_8 FILLER_24_616 ();
 sg13g2_decap_8 FILLER_24_623 ();
 sg13g2_decap_8 FILLER_24_630 ();
 sg13g2_decap_8 FILLER_24_637 ();
 sg13g2_decap_8 FILLER_24_644 ();
 sg13g2_decap_8 FILLER_24_651 ();
 sg13g2_decap_8 FILLER_24_658 ();
 sg13g2_decap_8 FILLER_24_665 ();
 sg13g2_decap_8 FILLER_24_672 ();
 sg13g2_decap_8 FILLER_24_679 ();
 sg13g2_decap_8 FILLER_24_686 ();
 sg13g2_decap_8 FILLER_24_693 ();
 sg13g2_decap_8 FILLER_24_700 ();
 sg13g2_decap_8 FILLER_24_707 ();
 sg13g2_decap_8 FILLER_24_714 ();
 sg13g2_decap_8 FILLER_24_721 ();
 sg13g2_decap_8 FILLER_24_728 ();
 sg13g2_decap_8 FILLER_24_735 ();
 sg13g2_decap_8 FILLER_24_742 ();
 sg13g2_decap_8 FILLER_24_749 ();
 sg13g2_decap_8 FILLER_24_756 ();
 sg13g2_decap_8 FILLER_24_763 ();
 sg13g2_decap_8 FILLER_24_770 ();
 sg13g2_decap_8 FILLER_24_777 ();
 sg13g2_decap_8 FILLER_24_784 ();
 sg13g2_decap_8 FILLER_24_791 ();
 sg13g2_decap_8 FILLER_24_798 ();
 sg13g2_decap_8 FILLER_24_805 ();
 sg13g2_decap_8 FILLER_24_812 ();
 sg13g2_decap_8 FILLER_24_819 ();
 sg13g2_decap_8 FILLER_24_826 ();
 sg13g2_decap_8 FILLER_24_833 ();
 sg13g2_decap_8 FILLER_24_840 ();
 sg13g2_decap_8 FILLER_24_847 ();
 sg13g2_decap_8 FILLER_24_854 ();
 sg13g2_fill_1 FILLER_24_861 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_fill_2 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_279 ();
 sg13g2_decap_8 FILLER_25_286 ();
 sg13g2_decap_8 FILLER_25_293 ();
 sg13g2_decap_8 FILLER_25_300 ();
 sg13g2_decap_8 FILLER_25_307 ();
 sg13g2_decap_8 FILLER_25_314 ();
 sg13g2_decap_8 FILLER_25_321 ();
 sg13g2_decap_8 FILLER_25_328 ();
 sg13g2_decap_8 FILLER_25_335 ();
 sg13g2_decap_8 FILLER_25_342 ();
 sg13g2_decap_8 FILLER_25_349 ();
 sg13g2_decap_8 FILLER_25_356 ();
 sg13g2_decap_8 FILLER_25_363 ();
 sg13g2_fill_1 FILLER_25_370 ();
 sg13g2_decap_8 FILLER_25_375 ();
 sg13g2_decap_4 FILLER_25_382 ();
 sg13g2_fill_2 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_decap_8 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_25_414 ();
 sg13g2_decap_8 FILLER_25_421 ();
 sg13g2_decap_8 FILLER_25_428 ();
 sg13g2_decap_8 FILLER_25_435 ();
 sg13g2_decap_8 FILLER_25_442 ();
 sg13g2_decap_8 FILLER_25_449 ();
 sg13g2_decap_8 FILLER_25_456 ();
 sg13g2_decap_8 FILLER_25_463 ();
 sg13g2_decap_8 FILLER_25_470 ();
 sg13g2_decap_8 FILLER_25_477 ();
 sg13g2_decap_8 FILLER_25_484 ();
 sg13g2_decap_8 FILLER_25_491 ();
 sg13g2_decap_8 FILLER_25_498 ();
 sg13g2_decap_8 FILLER_25_505 ();
 sg13g2_decap_8 FILLER_25_512 ();
 sg13g2_decap_8 FILLER_25_519 ();
 sg13g2_decap_8 FILLER_25_526 ();
 sg13g2_decap_8 FILLER_25_533 ();
 sg13g2_decap_8 FILLER_25_540 ();
 sg13g2_decap_8 FILLER_25_547 ();
 sg13g2_decap_8 FILLER_25_554 ();
 sg13g2_decap_8 FILLER_25_561 ();
 sg13g2_decap_8 FILLER_25_568 ();
 sg13g2_decap_8 FILLER_25_575 ();
 sg13g2_decap_8 FILLER_25_582 ();
 sg13g2_decap_8 FILLER_25_589 ();
 sg13g2_decap_8 FILLER_25_596 ();
 sg13g2_decap_8 FILLER_25_603 ();
 sg13g2_decap_8 FILLER_25_610 ();
 sg13g2_decap_8 FILLER_25_617 ();
 sg13g2_decap_8 FILLER_25_624 ();
 sg13g2_decap_8 FILLER_25_631 ();
 sg13g2_decap_8 FILLER_25_638 ();
 sg13g2_decap_8 FILLER_25_645 ();
 sg13g2_decap_8 FILLER_25_652 ();
 sg13g2_decap_8 FILLER_25_659 ();
 sg13g2_decap_8 FILLER_25_666 ();
 sg13g2_decap_8 FILLER_25_673 ();
 sg13g2_decap_8 FILLER_25_680 ();
 sg13g2_decap_8 FILLER_25_687 ();
 sg13g2_decap_8 FILLER_25_694 ();
 sg13g2_decap_8 FILLER_25_701 ();
 sg13g2_decap_8 FILLER_25_708 ();
 sg13g2_decap_8 FILLER_25_715 ();
 sg13g2_decap_8 FILLER_25_722 ();
 sg13g2_decap_8 FILLER_25_729 ();
 sg13g2_decap_8 FILLER_25_736 ();
 sg13g2_decap_8 FILLER_25_743 ();
 sg13g2_decap_8 FILLER_25_750 ();
 sg13g2_decap_8 FILLER_25_757 ();
 sg13g2_decap_8 FILLER_25_764 ();
 sg13g2_decap_8 FILLER_25_771 ();
 sg13g2_decap_8 FILLER_25_778 ();
 sg13g2_decap_8 FILLER_25_785 ();
 sg13g2_decap_8 FILLER_25_792 ();
 sg13g2_decap_8 FILLER_25_799 ();
 sg13g2_decap_8 FILLER_25_806 ();
 sg13g2_decap_8 FILLER_25_813 ();
 sg13g2_decap_8 FILLER_25_820 ();
 sg13g2_decap_8 FILLER_25_827 ();
 sg13g2_decap_8 FILLER_25_834 ();
 sg13g2_decap_8 FILLER_25_841 ();
 sg13g2_decap_8 FILLER_25_848 ();
 sg13g2_decap_8 FILLER_25_855 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_4 FILLER_26_63 ();
 sg13g2_fill_1 FILLER_26_67 ();
 sg13g2_fill_1 FILLER_26_94 ();
 sg13g2_decap_4 FILLER_26_104 ();
 sg13g2_fill_1 FILLER_26_108 ();
 sg13g2_decap_8 FILLER_26_113 ();
 sg13g2_decap_8 FILLER_26_120 ();
 sg13g2_decap_8 FILLER_26_127 ();
 sg13g2_decap_8 FILLER_26_134 ();
 sg13g2_decap_8 FILLER_26_141 ();
 sg13g2_decap_8 FILLER_26_148 ();
 sg13g2_decap_8 FILLER_26_155 ();
 sg13g2_decap_8 FILLER_26_162 ();
 sg13g2_decap_8 FILLER_26_169 ();
 sg13g2_decap_8 FILLER_26_176 ();
 sg13g2_decap_8 FILLER_26_183 ();
 sg13g2_decap_8 FILLER_26_190 ();
 sg13g2_decap_8 FILLER_26_197 ();
 sg13g2_decap_8 FILLER_26_204 ();
 sg13g2_decap_8 FILLER_26_211 ();
 sg13g2_decap_8 FILLER_26_218 ();
 sg13g2_decap_8 FILLER_26_225 ();
 sg13g2_decap_8 FILLER_26_232 ();
 sg13g2_decap_8 FILLER_26_239 ();
 sg13g2_decap_8 FILLER_26_246 ();
 sg13g2_decap_8 FILLER_26_253 ();
 sg13g2_fill_2 FILLER_26_260 ();
 sg13g2_fill_1 FILLER_26_262 ();
 sg13g2_fill_1 FILLER_26_267 ();
 sg13g2_fill_2 FILLER_26_277 ();
 sg13g2_decap_8 FILLER_26_302 ();
 sg13g2_decap_8 FILLER_26_332 ();
 sg13g2_decap_8 FILLER_26_339 ();
 sg13g2_decap_8 FILLER_26_346 ();
 sg13g2_decap_4 FILLER_26_353 ();
 sg13g2_fill_2 FILLER_26_357 ();
 sg13g2_fill_1 FILLER_26_367 ();
 sg13g2_fill_1 FILLER_26_373 ();
 sg13g2_decap_4 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_402 ();
 sg13g2_decap_8 FILLER_26_409 ();
 sg13g2_decap_4 FILLER_26_416 ();
 sg13g2_fill_1 FILLER_26_420 ();
 sg13g2_decap_8 FILLER_26_430 ();
 sg13g2_decap_8 FILLER_26_437 ();
 sg13g2_decap_8 FILLER_26_444 ();
 sg13g2_decap_8 FILLER_26_451 ();
 sg13g2_decap_8 FILLER_26_458 ();
 sg13g2_decap_8 FILLER_26_465 ();
 sg13g2_decap_8 FILLER_26_472 ();
 sg13g2_decap_8 FILLER_26_479 ();
 sg13g2_decap_8 FILLER_26_486 ();
 sg13g2_decap_8 FILLER_26_493 ();
 sg13g2_decap_8 FILLER_26_500 ();
 sg13g2_decap_8 FILLER_26_507 ();
 sg13g2_decap_8 FILLER_26_514 ();
 sg13g2_decap_8 FILLER_26_521 ();
 sg13g2_decap_8 FILLER_26_528 ();
 sg13g2_decap_8 FILLER_26_535 ();
 sg13g2_decap_8 FILLER_26_542 ();
 sg13g2_decap_8 FILLER_26_549 ();
 sg13g2_decap_8 FILLER_26_556 ();
 sg13g2_decap_8 FILLER_26_563 ();
 sg13g2_decap_8 FILLER_26_570 ();
 sg13g2_decap_8 FILLER_26_577 ();
 sg13g2_decap_8 FILLER_26_584 ();
 sg13g2_decap_8 FILLER_26_591 ();
 sg13g2_decap_8 FILLER_26_598 ();
 sg13g2_decap_8 FILLER_26_605 ();
 sg13g2_decap_8 FILLER_26_612 ();
 sg13g2_decap_8 FILLER_26_619 ();
 sg13g2_decap_8 FILLER_26_626 ();
 sg13g2_decap_8 FILLER_26_633 ();
 sg13g2_decap_8 FILLER_26_640 ();
 sg13g2_decap_8 FILLER_26_647 ();
 sg13g2_decap_8 FILLER_26_654 ();
 sg13g2_decap_8 FILLER_26_661 ();
 sg13g2_decap_8 FILLER_26_668 ();
 sg13g2_decap_8 FILLER_26_675 ();
 sg13g2_decap_8 FILLER_26_682 ();
 sg13g2_decap_8 FILLER_26_689 ();
 sg13g2_decap_8 FILLER_26_696 ();
 sg13g2_decap_8 FILLER_26_703 ();
 sg13g2_decap_8 FILLER_26_710 ();
 sg13g2_decap_8 FILLER_26_717 ();
 sg13g2_decap_8 FILLER_26_724 ();
 sg13g2_decap_8 FILLER_26_731 ();
 sg13g2_decap_8 FILLER_26_738 ();
 sg13g2_decap_8 FILLER_26_745 ();
 sg13g2_decap_8 FILLER_26_752 ();
 sg13g2_decap_8 FILLER_26_759 ();
 sg13g2_decap_8 FILLER_26_766 ();
 sg13g2_decap_8 FILLER_26_773 ();
 sg13g2_decap_8 FILLER_26_780 ();
 sg13g2_decap_8 FILLER_26_787 ();
 sg13g2_decap_8 FILLER_26_794 ();
 sg13g2_decap_8 FILLER_26_801 ();
 sg13g2_decap_8 FILLER_26_808 ();
 sg13g2_decap_8 FILLER_26_815 ();
 sg13g2_decap_8 FILLER_26_822 ();
 sg13g2_decap_8 FILLER_26_829 ();
 sg13g2_decap_8 FILLER_26_836 ();
 sg13g2_decap_8 FILLER_26_843 ();
 sg13g2_decap_8 FILLER_26_850 ();
 sg13g2_decap_4 FILLER_26_857 ();
 sg13g2_fill_1 FILLER_26_861 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_4 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_57 ();
 sg13g2_fill_1 FILLER_27_79 ();
 sg13g2_fill_2 FILLER_27_88 ();
 sg13g2_decap_4 FILLER_27_120 ();
 sg13g2_fill_2 FILLER_27_124 ();
 sg13g2_decap_8 FILLER_27_136 ();
 sg13g2_decap_8 FILLER_27_143 ();
 sg13g2_decap_8 FILLER_27_150 ();
 sg13g2_decap_8 FILLER_27_157 ();
 sg13g2_decap_8 FILLER_27_164 ();
 sg13g2_decap_8 FILLER_27_171 ();
 sg13g2_decap_8 FILLER_27_178 ();
 sg13g2_decap_8 FILLER_27_185 ();
 sg13g2_decap_8 FILLER_27_192 ();
 sg13g2_decap_8 FILLER_27_199 ();
 sg13g2_decap_8 FILLER_27_206 ();
 sg13g2_fill_2 FILLER_27_213 ();
 sg13g2_decap_4 FILLER_27_226 ();
 sg13g2_decap_8 FILLER_27_246 ();
 sg13g2_fill_1 FILLER_27_253 ();
 sg13g2_fill_2 FILLER_27_284 ();
 sg13g2_fill_1 FILLER_27_286 ();
 sg13g2_fill_2 FILLER_27_342 ();
 sg13g2_fill_2 FILLER_27_353 ();
 sg13g2_fill_1 FILLER_27_355 ();
 sg13g2_fill_2 FILLER_27_434 ();
 sg13g2_fill_1 FILLER_27_436 ();
 sg13g2_decap_8 FILLER_27_441 ();
 sg13g2_decap_8 FILLER_27_448 ();
 sg13g2_decap_8 FILLER_27_455 ();
 sg13g2_decap_8 FILLER_27_462 ();
 sg13g2_decap_8 FILLER_27_469 ();
 sg13g2_decap_8 FILLER_27_476 ();
 sg13g2_decap_8 FILLER_27_483 ();
 sg13g2_decap_8 FILLER_27_490 ();
 sg13g2_decap_8 FILLER_27_497 ();
 sg13g2_decap_8 FILLER_27_504 ();
 sg13g2_decap_8 FILLER_27_511 ();
 sg13g2_decap_8 FILLER_27_518 ();
 sg13g2_decap_8 FILLER_27_525 ();
 sg13g2_decap_8 FILLER_27_532 ();
 sg13g2_decap_8 FILLER_27_539 ();
 sg13g2_decap_8 FILLER_27_546 ();
 sg13g2_decap_8 FILLER_27_553 ();
 sg13g2_decap_8 FILLER_27_560 ();
 sg13g2_decap_8 FILLER_27_567 ();
 sg13g2_decap_8 FILLER_27_574 ();
 sg13g2_decap_8 FILLER_27_581 ();
 sg13g2_decap_8 FILLER_27_588 ();
 sg13g2_decap_8 FILLER_27_595 ();
 sg13g2_decap_8 FILLER_27_602 ();
 sg13g2_decap_8 FILLER_27_609 ();
 sg13g2_decap_8 FILLER_27_616 ();
 sg13g2_decap_8 FILLER_27_623 ();
 sg13g2_decap_8 FILLER_27_630 ();
 sg13g2_decap_8 FILLER_27_637 ();
 sg13g2_decap_8 FILLER_27_644 ();
 sg13g2_decap_8 FILLER_27_651 ();
 sg13g2_decap_8 FILLER_27_658 ();
 sg13g2_decap_8 FILLER_27_665 ();
 sg13g2_decap_8 FILLER_27_672 ();
 sg13g2_decap_8 FILLER_27_679 ();
 sg13g2_decap_8 FILLER_27_686 ();
 sg13g2_decap_8 FILLER_27_693 ();
 sg13g2_decap_8 FILLER_27_700 ();
 sg13g2_decap_8 FILLER_27_707 ();
 sg13g2_decap_8 FILLER_27_714 ();
 sg13g2_decap_8 FILLER_27_721 ();
 sg13g2_decap_8 FILLER_27_728 ();
 sg13g2_decap_8 FILLER_27_735 ();
 sg13g2_decap_8 FILLER_27_742 ();
 sg13g2_decap_8 FILLER_27_749 ();
 sg13g2_decap_8 FILLER_27_756 ();
 sg13g2_decap_8 FILLER_27_763 ();
 sg13g2_decap_8 FILLER_27_770 ();
 sg13g2_decap_8 FILLER_27_777 ();
 sg13g2_decap_8 FILLER_27_784 ();
 sg13g2_decap_8 FILLER_27_791 ();
 sg13g2_decap_8 FILLER_27_798 ();
 sg13g2_decap_8 FILLER_27_805 ();
 sg13g2_decap_8 FILLER_27_812 ();
 sg13g2_decap_8 FILLER_27_819 ();
 sg13g2_decap_8 FILLER_27_826 ();
 sg13g2_decap_8 FILLER_27_833 ();
 sg13g2_decap_8 FILLER_27_840 ();
 sg13g2_decap_8 FILLER_27_847 ();
 sg13g2_decap_8 FILLER_27_854 ();
 sg13g2_fill_1 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_fill_2 FILLER_28_68 ();
 sg13g2_fill_2 FILLER_28_88 ();
 sg13g2_fill_2 FILLER_28_106 ();
 sg13g2_fill_1 FILLER_28_108 ();
 sg13g2_fill_2 FILLER_28_114 ();
 sg13g2_fill_2 FILLER_28_140 ();
 sg13g2_fill_1 FILLER_28_142 ();
 sg13g2_decap_8 FILLER_28_160 ();
 sg13g2_decap_8 FILLER_28_193 ();
 sg13g2_decap_8 FILLER_28_200 ();
 sg13g2_fill_2 FILLER_28_207 ();
 sg13g2_fill_1 FILLER_28_209 ();
 sg13g2_fill_1 FILLER_28_248 ();
 sg13g2_fill_2 FILLER_28_275 ();
 sg13g2_fill_1 FILLER_28_295 ();
 sg13g2_fill_2 FILLER_28_310 ();
 sg13g2_fill_1 FILLER_28_312 ();
 sg13g2_fill_2 FILLER_28_331 ();
 sg13g2_fill_2 FILLER_28_376 ();
 sg13g2_fill_1 FILLER_28_378 ();
 sg13g2_fill_1 FILLER_28_388 ();
 sg13g2_decap_4 FILLER_28_452 ();
 sg13g2_fill_2 FILLER_28_456 ();
 sg13g2_decap_8 FILLER_28_484 ();
 sg13g2_decap_8 FILLER_28_491 ();
 sg13g2_decap_8 FILLER_28_498 ();
 sg13g2_decap_8 FILLER_28_505 ();
 sg13g2_decap_8 FILLER_28_512 ();
 sg13g2_decap_8 FILLER_28_519 ();
 sg13g2_decap_8 FILLER_28_526 ();
 sg13g2_decap_8 FILLER_28_533 ();
 sg13g2_decap_8 FILLER_28_540 ();
 sg13g2_decap_8 FILLER_28_547 ();
 sg13g2_decap_8 FILLER_28_554 ();
 sg13g2_decap_8 FILLER_28_584 ();
 sg13g2_decap_8 FILLER_28_591 ();
 sg13g2_decap_8 FILLER_28_598 ();
 sg13g2_decap_8 FILLER_28_605 ();
 sg13g2_decap_8 FILLER_28_612 ();
 sg13g2_decap_8 FILLER_28_619 ();
 sg13g2_decap_8 FILLER_28_626 ();
 sg13g2_decap_8 FILLER_28_633 ();
 sg13g2_decap_8 FILLER_28_640 ();
 sg13g2_decap_8 FILLER_28_647 ();
 sg13g2_decap_8 FILLER_28_654 ();
 sg13g2_decap_8 FILLER_28_661 ();
 sg13g2_decap_8 FILLER_28_668 ();
 sg13g2_decap_8 FILLER_28_675 ();
 sg13g2_decap_8 FILLER_28_682 ();
 sg13g2_decap_8 FILLER_28_689 ();
 sg13g2_decap_8 FILLER_28_696 ();
 sg13g2_decap_8 FILLER_28_703 ();
 sg13g2_decap_8 FILLER_28_710 ();
 sg13g2_decap_8 FILLER_28_717 ();
 sg13g2_decap_8 FILLER_28_724 ();
 sg13g2_decap_8 FILLER_28_731 ();
 sg13g2_decap_8 FILLER_28_738 ();
 sg13g2_decap_8 FILLER_28_745 ();
 sg13g2_decap_8 FILLER_28_752 ();
 sg13g2_decap_8 FILLER_28_759 ();
 sg13g2_decap_8 FILLER_28_766 ();
 sg13g2_decap_8 FILLER_28_773 ();
 sg13g2_decap_8 FILLER_28_780 ();
 sg13g2_decap_8 FILLER_28_787 ();
 sg13g2_decap_8 FILLER_28_794 ();
 sg13g2_decap_8 FILLER_28_801 ();
 sg13g2_decap_8 FILLER_28_808 ();
 sg13g2_decap_8 FILLER_28_815 ();
 sg13g2_decap_8 FILLER_28_822 ();
 sg13g2_decap_8 FILLER_28_829 ();
 sg13g2_decap_8 FILLER_28_836 ();
 sg13g2_decap_8 FILLER_28_843 ();
 sg13g2_decap_8 FILLER_28_850 ();
 sg13g2_decap_4 FILLER_28_857 ();
 sg13g2_fill_1 FILLER_28_861 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_4 FILLER_29_28 ();
 sg13g2_decap_4 FILLER_29_36 ();
 sg13g2_fill_2 FILLER_29_40 ();
 sg13g2_decap_8 FILLER_29_47 ();
 sg13g2_fill_2 FILLER_29_74 ();
 sg13g2_fill_1 FILLER_29_76 ();
 sg13g2_fill_2 FILLER_29_90 ();
 sg13g2_decap_4 FILLER_29_121 ();
 sg13g2_decap_4 FILLER_29_171 ();
 sg13g2_fill_2 FILLER_29_175 ();
 sg13g2_decap_4 FILLER_29_181 ();
 sg13g2_fill_2 FILLER_29_185 ();
 sg13g2_fill_2 FILLER_29_279 ();
 sg13g2_fill_2 FILLER_29_291 ();
 sg13g2_fill_2 FILLER_29_303 ();
 sg13g2_fill_2 FILLER_29_331 ();
 sg13g2_fill_2 FILLER_29_338 ();
 sg13g2_fill_2 FILLER_29_397 ();
 sg13g2_fill_1 FILLER_29_416 ();
 sg13g2_fill_1 FILLER_29_434 ();
 sg13g2_decap_4 FILLER_29_444 ();
 sg13g2_fill_2 FILLER_29_473 ();
 sg13g2_decap_8 FILLER_29_493 ();
 sg13g2_decap_8 FILLER_29_500 ();
 sg13g2_decap_8 FILLER_29_507 ();
 sg13g2_fill_1 FILLER_29_527 ();
 sg13g2_decap_8 FILLER_29_541 ();
 sg13g2_decap_8 FILLER_29_548 ();
 sg13g2_decap_4 FILLER_29_555 ();
 sg13g2_decap_8 FILLER_29_585 ();
 sg13g2_fill_2 FILLER_29_592 ();
 sg13g2_fill_1 FILLER_29_594 ();
 sg13g2_fill_2 FILLER_29_598 ();
 sg13g2_decap_8 FILLER_29_609 ();
 sg13g2_decap_8 FILLER_29_616 ();
 sg13g2_decap_8 FILLER_29_623 ();
 sg13g2_decap_8 FILLER_29_630 ();
 sg13g2_decap_8 FILLER_29_637 ();
 sg13g2_decap_8 FILLER_29_644 ();
 sg13g2_decap_8 FILLER_29_651 ();
 sg13g2_decap_8 FILLER_29_658 ();
 sg13g2_decap_8 FILLER_29_665 ();
 sg13g2_decap_8 FILLER_29_672 ();
 sg13g2_decap_8 FILLER_29_679 ();
 sg13g2_decap_8 FILLER_29_686 ();
 sg13g2_decap_8 FILLER_29_693 ();
 sg13g2_decap_8 FILLER_29_700 ();
 sg13g2_decap_8 FILLER_29_707 ();
 sg13g2_decap_8 FILLER_29_714 ();
 sg13g2_decap_8 FILLER_29_721 ();
 sg13g2_decap_8 FILLER_29_728 ();
 sg13g2_decap_8 FILLER_29_735 ();
 sg13g2_decap_8 FILLER_29_742 ();
 sg13g2_decap_8 FILLER_29_749 ();
 sg13g2_decap_8 FILLER_29_756 ();
 sg13g2_decap_8 FILLER_29_763 ();
 sg13g2_decap_8 FILLER_29_770 ();
 sg13g2_decap_8 FILLER_29_777 ();
 sg13g2_decap_8 FILLER_29_784 ();
 sg13g2_decap_8 FILLER_29_791 ();
 sg13g2_decap_8 FILLER_29_798 ();
 sg13g2_decap_8 FILLER_29_805 ();
 sg13g2_decap_8 FILLER_29_812 ();
 sg13g2_decap_8 FILLER_29_819 ();
 sg13g2_decap_8 FILLER_29_826 ();
 sg13g2_decap_8 FILLER_29_833 ();
 sg13g2_decap_8 FILLER_29_840 ();
 sg13g2_decap_8 FILLER_29_847 ();
 sg13g2_decap_8 FILLER_29_854 ();
 sg13g2_fill_1 FILLER_29_861 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_4 FILLER_30_71 ();
 sg13g2_fill_1 FILLER_30_75 ();
 sg13g2_decap_4 FILLER_30_93 ();
 sg13g2_fill_2 FILLER_30_97 ();
 sg13g2_fill_2 FILLER_30_103 ();
 sg13g2_fill_2 FILLER_30_116 ();
 sg13g2_fill_2 FILLER_30_126 ();
 sg13g2_fill_1 FILLER_30_128 ();
 sg13g2_decap_4 FILLER_30_134 ();
 sg13g2_fill_1 FILLER_30_138 ();
 sg13g2_decap_8 FILLER_30_144 ();
 sg13g2_fill_2 FILLER_30_151 ();
 sg13g2_fill_2 FILLER_30_165 ();
 sg13g2_fill_2 FILLER_30_172 ();
 sg13g2_fill_1 FILLER_30_174 ();
 sg13g2_fill_1 FILLER_30_180 ();
 sg13g2_decap_8 FILLER_30_184 ();
 sg13g2_decap_4 FILLER_30_191 ();
 sg13g2_fill_1 FILLER_30_195 ();
 sg13g2_fill_1 FILLER_30_242 ();
 sg13g2_fill_1 FILLER_30_278 ();
 sg13g2_fill_1 FILLER_30_301 ();
 sg13g2_fill_2 FILLER_30_337 ();
 sg13g2_fill_1 FILLER_30_339 ();
 sg13g2_fill_1 FILLER_30_350 ();
 sg13g2_fill_2 FILLER_30_360 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_fill_2 FILLER_30_373 ();
 sg13g2_decap_4 FILLER_30_391 ();
 sg13g2_fill_2 FILLER_30_410 ();
 sg13g2_fill_2 FILLER_30_424 ();
 sg13g2_fill_1 FILLER_30_426 ();
 sg13g2_fill_2 FILLER_30_440 ();
 sg13g2_fill_1 FILLER_30_442 ();
 sg13g2_fill_1 FILLER_30_448 ();
 sg13g2_fill_2 FILLER_30_465 ();
 sg13g2_decap_4 FILLER_30_498 ();
 sg13g2_fill_2 FILLER_30_502 ();
 sg13g2_decap_4 FILLER_30_530 ();
 sg13g2_fill_1 FILLER_30_603 ();
 sg13g2_decap_8 FILLER_30_630 ();
 sg13g2_decap_8 FILLER_30_637 ();
 sg13g2_decap_8 FILLER_30_644 ();
 sg13g2_decap_8 FILLER_30_651 ();
 sg13g2_decap_8 FILLER_30_658 ();
 sg13g2_decap_8 FILLER_30_665 ();
 sg13g2_decap_8 FILLER_30_672 ();
 sg13g2_decap_8 FILLER_30_679 ();
 sg13g2_decap_8 FILLER_30_686 ();
 sg13g2_decap_8 FILLER_30_693 ();
 sg13g2_decap_8 FILLER_30_700 ();
 sg13g2_decap_8 FILLER_30_707 ();
 sg13g2_decap_8 FILLER_30_714 ();
 sg13g2_decap_8 FILLER_30_721 ();
 sg13g2_decap_8 FILLER_30_728 ();
 sg13g2_decap_8 FILLER_30_735 ();
 sg13g2_decap_8 FILLER_30_742 ();
 sg13g2_decap_8 FILLER_30_749 ();
 sg13g2_decap_8 FILLER_30_756 ();
 sg13g2_decap_8 FILLER_30_763 ();
 sg13g2_decap_8 FILLER_30_770 ();
 sg13g2_decap_8 FILLER_30_777 ();
 sg13g2_decap_8 FILLER_30_784 ();
 sg13g2_decap_8 FILLER_30_791 ();
 sg13g2_decap_8 FILLER_30_798 ();
 sg13g2_decap_8 FILLER_30_805 ();
 sg13g2_decap_8 FILLER_30_812 ();
 sg13g2_decap_8 FILLER_30_819 ();
 sg13g2_decap_8 FILLER_30_826 ();
 sg13g2_decap_8 FILLER_30_833 ();
 sg13g2_decap_8 FILLER_30_840 ();
 sg13g2_decap_8 FILLER_30_847 ();
 sg13g2_decap_8 FILLER_30_854 ();
 sg13g2_fill_1 FILLER_30_861 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_fill_2 FILLER_31_21 ();
 sg13g2_fill_2 FILLER_31_32 ();
 sg13g2_fill_1 FILLER_31_34 ();
 sg13g2_fill_1 FILLER_31_64 ();
 sg13g2_fill_2 FILLER_31_73 ();
 sg13g2_fill_1 FILLER_31_75 ();
 sg13g2_fill_1 FILLER_31_105 ();
 sg13g2_fill_1 FILLER_31_123 ();
 sg13g2_fill_1 FILLER_31_134 ();
 sg13g2_fill_1 FILLER_31_143 ();
 sg13g2_fill_1 FILLER_31_152 ();
 sg13g2_fill_1 FILLER_31_171 ();
 sg13g2_decap_4 FILLER_31_194 ();
 sg13g2_fill_1 FILLER_31_198 ();
 sg13g2_fill_1 FILLER_31_223 ();
 sg13g2_fill_1 FILLER_31_254 ();
 sg13g2_fill_2 FILLER_31_264 ();
 sg13g2_fill_1 FILLER_31_297 ();
 sg13g2_fill_2 FILLER_31_306 ();
 sg13g2_fill_1 FILLER_31_308 ();
 sg13g2_fill_2 FILLER_31_314 ();
 sg13g2_fill_2 FILLER_31_356 ();
 sg13g2_fill_1 FILLER_31_384 ();
 sg13g2_decap_4 FILLER_31_394 ();
 sg13g2_fill_2 FILLER_31_409 ();
 sg13g2_fill_1 FILLER_31_473 ();
 sg13g2_fill_2 FILLER_31_501 ();
 sg13g2_decap_8 FILLER_31_517 ();
 sg13g2_decap_4 FILLER_31_524 ();
 sg13g2_fill_1 FILLER_31_528 ();
 sg13g2_fill_1 FILLER_31_534 ();
 sg13g2_fill_1 FILLER_31_566 ();
 sg13g2_fill_2 FILLER_31_581 ();
 sg13g2_decap_8 FILLER_31_638 ();
 sg13g2_decap_8 FILLER_31_645 ();
 sg13g2_decap_8 FILLER_31_652 ();
 sg13g2_decap_8 FILLER_31_659 ();
 sg13g2_decap_8 FILLER_31_666 ();
 sg13g2_decap_8 FILLER_31_673 ();
 sg13g2_decap_8 FILLER_31_680 ();
 sg13g2_decap_8 FILLER_31_687 ();
 sg13g2_decap_8 FILLER_31_694 ();
 sg13g2_decap_8 FILLER_31_701 ();
 sg13g2_decap_8 FILLER_31_708 ();
 sg13g2_decap_8 FILLER_31_715 ();
 sg13g2_decap_8 FILLER_31_722 ();
 sg13g2_decap_8 FILLER_31_729 ();
 sg13g2_decap_8 FILLER_31_736 ();
 sg13g2_decap_8 FILLER_31_743 ();
 sg13g2_decap_8 FILLER_31_750 ();
 sg13g2_decap_8 FILLER_31_757 ();
 sg13g2_decap_8 FILLER_31_764 ();
 sg13g2_decap_8 FILLER_31_771 ();
 sg13g2_decap_8 FILLER_31_778 ();
 sg13g2_decap_8 FILLER_31_785 ();
 sg13g2_decap_8 FILLER_31_792 ();
 sg13g2_decap_8 FILLER_31_799 ();
 sg13g2_decap_8 FILLER_31_806 ();
 sg13g2_decap_8 FILLER_31_813 ();
 sg13g2_decap_8 FILLER_31_820 ();
 sg13g2_decap_8 FILLER_31_827 ();
 sg13g2_decap_8 FILLER_31_834 ();
 sg13g2_decap_8 FILLER_31_841 ();
 sg13g2_decap_8 FILLER_31_848 ();
 sg13g2_decap_8 FILLER_31_855 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_50 ();
 sg13g2_fill_1 FILLER_32_68 ();
 sg13g2_decap_4 FILLER_32_72 ();
 sg13g2_fill_2 FILLER_32_76 ();
 sg13g2_fill_2 FILLER_32_85 ();
 sg13g2_decap_8 FILLER_32_114 ();
 sg13g2_fill_1 FILLER_32_121 ();
 sg13g2_fill_2 FILLER_32_126 ();
 sg13g2_decap_4 FILLER_32_137 ();
 sg13g2_fill_2 FILLER_32_141 ();
 sg13g2_fill_2 FILLER_32_167 ();
 sg13g2_fill_1 FILLER_32_201 ();
 sg13g2_fill_1 FILLER_32_269 ();
 sg13g2_fill_2 FILLER_32_311 ();
 sg13g2_fill_2 FILLER_32_323 ();
 sg13g2_fill_1 FILLER_32_333 ();
 sg13g2_fill_2 FILLER_32_346 ();
 sg13g2_decap_4 FILLER_32_385 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_fill_2 FILLER_32_415 ();
 sg13g2_fill_1 FILLER_32_417 ();
 sg13g2_fill_1 FILLER_32_462 ();
 sg13g2_fill_1 FILLER_32_473 ();
 sg13g2_fill_1 FILLER_32_505 ();
 sg13g2_fill_2 FILLER_32_554 ();
 sg13g2_fill_2 FILLER_32_561 ();
 sg13g2_fill_1 FILLER_32_606 ();
 sg13g2_fill_1 FILLER_32_619 ();
 sg13g2_decap_8 FILLER_32_663 ();
 sg13g2_decap_8 FILLER_32_670 ();
 sg13g2_decap_8 FILLER_32_677 ();
 sg13g2_decap_8 FILLER_32_684 ();
 sg13g2_decap_8 FILLER_32_691 ();
 sg13g2_decap_8 FILLER_32_698 ();
 sg13g2_decap_8 FILLER_32_705 ();
 sg13g2_decap_8 FILLER_32_712 ();
 sg13g2_decap_8 FILLER_32_719 ();
 sg13g2_decap_8 FILLER_32_726 ();
 sg13g2_decap_8 FILLER_32_733 ();
 sg13g2_decap_8 FILLER_32_740 ();
 sg13g2_decap_8 FILLER_32_747 ();
 sg13g2_decap_8 FILLER_32_754 ();
 sg13g2_decap_8 FILLER_32_761 ();
 sg13g2_decap_8 FILLER_32_768 ();
 sg13g2_decap_8 FILLER_32_775 ();
 sg13g2_decap_8 FILLER_32_782 ();
 sg13g2_decap_8 FILLER_32_789 ();
 sg13g2_decap_8 FILLER_32_796 ();
 sg13g2_decap_8 FILLER_32_803 ();
 sg13g2_decap_8 FILLER_32_810 ();
 sg13g2_decap_8 FILLER_32_817 ();
 sg13g2_decap_8 FILLER_32_824 ();
 sg13g2_decap_8 FILLER_32_831 ();
 sg13g2_decap_8 FILLER_32_838 ();
 sg13g2_decap_8 FILLER_32_845 ();
 sg13g2_decap_8 FILLER_32_852 ();
 sg13g2_fill_2 FILLER_32_859 ();
 sg13g2_fill_1 FILLER_32_861 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_11 ();
 sg13g2_decap_8 FILLER_33_16 ();
 sg13g2_fill_2 FILLER_33_23 ();
 sg13g2_fill_1 FILLER_33_25 ();
 sg13g2_fill_2 FILLER_33_52 ();
 sg13g2_fill_2 FILLER_33_67 ();
 sg13g2_fill_1 FILLER_33_69 ();
 sg13g2_decap_8 FILLER_33_78 ();
 sg13g2_decap_4 FILLER_33_85 ();
 sg13g2_fill_2 FILLER_33_89 ();
 sg13g2_fill_2 FILLER_33_111 ();
 sg13g2_fill_1 FILLER_33_128 ();
 sg13g2_fill_2 FILLER_33_155 ();
 sg13g2_decap_4 FILLER_33_197 ();
 sg13g2_fill_2 FILLER_33_223 ();
 sg13g2_fill_1 FILLER_33_225 ();
 sg13g2_fill_1 FILLER_33_297 ();
 sg13g2_fill_2 FILLER_33_307 ();
 sg13g2_fill_1 FILLER_33_309 ();
 sg13g2_decap_4 FILLER_33_326 ();
 sg13g2_fill_2 FILLER_33_330 ();
 sg13g2_fill_1 FILLER_33_372 ();
 sg13g2_fill_1 FILLER_33_382 ();
 sg13g2_fill_1 FILLER_33_398 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_fill_1 FILLER_33_419 ();
 sg13g2_fill_2 FILLER_33_428 ();
 sg13g2_fill_1 FILLER_33_430 ();
 sg13g2_fill_2 FILLER_33_440 ();
 sg13g2_decap_4 FILLER_33_494 ();
 sg13g2_fill_2 FILLER_33_498 ();
 sg13g2_decap_4 FILLER_33_593 ();
 sg13g2_fill_2 FILLER_33_597 ();
 sg13g2_decap_4 FILLER_33_630 ();
 sg13g2_fill_1 FILLER_33_634 ();
 sg13g2_decap_8 FILLER_33_644 ();
 sg13g2_decap_8 FILLER_33_651 ();
 sg13g2_decap_8 FILLER_33_658 ();
 sg13g2_decap_8 FILLER_33_665 ();
 sg13g2_decap_8 FILLER_33_672 ();
 sg13g2_decap_8 FILLER_33_679 ();
 sg13g2_decap_8 FILLER_33_686 ();
 sg13g2_decap_8 FILLER_33_693 ();
 sg13g2_decap_8 FILLER_33_700 ();
 sg13g2_decap_8 FILLER_33_707 ();
 sg13g2_decap_8 FILLER_33_714 ();
 sg13g2_decap_8 FILLER_33_721 ();
 sg13g2_decap_8 FILLER_33_728 ();
 sg13g2_decap_8 FILLER_33_735 ();
 sg13g2_decap_8 FILLER_33_742 ();
 sg13g2_decap_8 FILLER_33_749 ();
 sg13g2_decap_8 FILLER_33_756 ();
 sg13g2_decap_8 FILLER_33_763 ();
 sg13g2_decap_8 FILLER_33_770 ();
 sg13g2_decap_8 FILLER_33_777 ();
 sg13g2_decap_8 FILLER_33_784 ();
 sg13g2_decap_8 FILLER_33_791 ();
 sg13g2_decap_8 FILLER_33_798 ();
 sg13g2_decap_8 FILLER_33_805 ();
 sg13g2_decap_8 FILLER_33_812 ();
 sg13g2_decap_8 FILLER_33_819 ();
 sg13g2_decap_8 FILLER_33_826 ();
 sg13g2_decap_8 FILLER_33_833 ();
 sg13g2_decap_8 FILLER_33_840 ();
 sg13g2_decap_8 FILLER_33_847 ();
 sg13g2_decap_8 FILLER_33_854 ();
 sg13g2_fill_1 FILLER_33_861 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_fill_2 FILLER_34_28 ();
 sg13g2_fill_1 FILLER_34_30 ();
 sg13g2_fill_1 FILLER_34_55 ();
 sg13g2_decap_8 FILLER_34_78 ();
 sg13g2_decap_4 FILLER_34_85 ();
 sg13g2_fill_1 FILLER_34_89 ();
 sg13g2_decap_8 FILLER_34_96 ();
 sg13g2_decap_8 FILLER_34_103 ();
 sg13g2_decap_4 FILLER_34_110 ();
 sg13g2_fill_2 FILLER_34_140 ();
 sg13g2_decap_4 FILLER_34_199 ();
 sg13g2_fill_2 FILLER_34_203 ();
 sg13g2_decap_4 FILLER_34_213 ();
 sg13g2_fill_1 FILLER_34_217 ();
 sg13g2_fill_1 FILLER_34_261 ();
 sg13g2_fill_2 FILLER_34_313 ();
 sg13g2_fill_1 FILLER_34_315 ();
 sg13g2_decap_4 FILLER_34_323 ();
 sg13g2_fill_1 FILLER_34_327 ();
 sg13g2_decap_8 FILLER_34_332 ();
 sg13g2_decap_4 FILLER_34_339 ();
 sg13g2_fill_2 FILLER_34_373 ();
 sg13g2_fill_1 FILLER_34_402 ();
 sg13g2_fill_2 FILLER_34_414 ();
 sg13g2_fill_2 FILLER_34_426 ();
 sg13g2_fill_1 FILLER_34_428 ();
 sg13g2_fill_2 FILLER_34_553 ();
 sg13g2_fill_1 FILLER_34_555 ();
 sg13g2_fill_2 FILLER_34_591 ();
 sg13g2_fill_2 FILLER_34_609 ();
 sg13g2_fill_2 FILLER_34_628 ();
 sg13g2_decap_4 FILLER_34_642 ();
 sg13g2_decap_8 FILLER_34_659 ();
 sg13g2_decap_8 FILLER_34_666 ();
 sg13g2_decap_8 FILLER_34_673 ();
 sg13g2_decap_8 FILLER_34_680 ();
 sg13g2_decap_8 FILLER_34_687 ();
 sg13g2_decap_8 FILLER_34_694 ();
 sg13g2_decap_8 FILLER_34_701 ();
 sg13g2_decap_8 FILLER_34_708 ();
 sg13g2_decap_8 FILLER_34_715 ();
 sg13g2_decap_8 FILLER_34_722 ();
 sg13g2_decap_8 FILLER_34_729 ();
 sg13g2_decap_8 FILLER_34_736 ();
 sg13g2_decap_8 FILLER_34_743 ();
 sg13g2_decap_8 FILLER_34_750 ();
 sg13g2_decap_8 FILLER_34_757 ();
 sg13g2_decap_8 FILLER_34_764 ();
 sg13g2_decap_8 FILLER_34_771 ();
 sg13g2_decap_8 FILLER_34_778 ();
 sg13g2_decap_8 FILLER_34_785 ();
 sg13g2_decap_8 FILLER_34_792 ();
 sg13g2_decap_8 FILLER_34_799 ();
 sg13g2_decap_8 FILLER_34_806 ();
 sg13g2_decap_8 FILLER_34_813 ();
 sg13g2_decap_8 FILLER_34_820 ();
 sg13g2_decap_8 FILLER_34_827 ();
 sg13g2_decap_8 FILLER_34_834 ();
 sg13g2_decap_8 FILLER_34_841 ();
 sg13g2_decap_8 FILLER_34_848 ();
 sg13g2_decap_8 FILLER_34_855 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_fill_1 FILLER_35_57 ();
 sg13g2_fill_2 FILLER_35_80 ();
 sg13g2_decap_8 FILLER_35_87 ();
 sg13g2_fill_1 FILLER_35_94 ();
 sg13g2_fill_2 FILLER_35_158 ();
 sg13g2_decap_4 FILLER_35_178 ();
 sg13g2_decap_8 FILLER_35_195 ();
 sg13g2_fill_1 FILLER_35_202 ();
 sg13g2_fill_1 FILLER_35_229 ();
 sg13g2_fill_1 FILLER_35_255 ();
 sg13g2_fill_1 FILLER_35_281 ();
 sg13g2_fill_1 FILLER_35_316 ();
 sg13g2_fill_2 FILLER_35_348 ();
 sg13g2_fill_1 FILLER_35_421 ();
 sg13g2_decap_4 FILLER_35_448 ();
 sg13g2_fill_2 FILLER_35_452 ();
 sg13g2_decap_4 FILLER_35_474 ();
 sg13g2_fill_1 FILLER_35_478 ();
 sg13g2_fill_1 FILLER_35_484 ();
 sg13g2_decap_8 FILLER_35_489 ();
 sg13g2_decap_8 FILLER_35_496 ();
 sg13g2_fill_2 FILLER_35_503 ();
 sg13g2_fill_2 FILLER_35_596 ();
 sg13g2_fill_2 FILLER_35_608 ();
 sg13g2_fill_1 FILLER_35_622 ();
 sg13g2_fill_2 FILLER_35_645 ();
 sg13g2_decap_8 FILLER_35_668 ();
 sg13g2_decap_8 FILLER_35_675 ();
 sg13g2_decap_8 FILLER_35_682 ();
 sg13g2_decap_8 FILLER_35_689 ();
 sg13g2_decap_8 FILLER_35_696 ();
 sg13g2_decap_8 FILLER_35_703 ();
 sg13g2_decap_8 FILLER_35_710 ();
 sg13g2_decap_8 FILLER_35_717 ();
 sg13g2_decap_8 FILLER_35_724 ();
 sg13g2_decap_8 FILLER_35_731 ();
 sg13g2_decap_8 FILLER_35_738 ();
 sg13g2_decap_8 FILLER_35_745 ();
 sg13g2_decap_8 FILLER_35_752 ();
 sg13g2_decap_8 FILLER_35_759 ();
 sg13g2_decap_8 FILLER_35_766 ();
 sg13g2_decap_8 FILLER_35_773 ();
 sg13g2_decap_8 FILLER_35_780 ();
 sg13g2_decap_8 FILLER_35_787 ();
 sg13g2_decap_8 FILLER_35_794 ();
 sg13g2_decap_8 FILLER_35_801 ();
 sg13g2_decap_8 FILLER_35_808 ();
 sg13g2_decap_8 FILLER_35_815 ();
 sg13g2_decap_8 FILLER_35_822 ();
 sg13g2_decap_8 FILLER_35_829 ();
 sg13g2_decap_8 FILLER_35_836 ();
 sg13g2_decap_8 FILLER_35_843 ();
 sg13g2_decap_8 FILLER_35_850 ();
 sg13g2_decap_4 FILLER_35_857 ();
 sg13g2_fill_1 FILLER_35_861 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_fill_2 FILLER_36_28 ();
 sg13g2_fill_1 FILLER_36_30 ();
 sg13g2_decap_8 FILLER_36_53 ();
 sg13g2_fill_1 FILLER_36_88 ();
 sg13g2_decap_4 FILLER_36_94 ();
 sg13g2_fill_2 FILLER_36_98 ();
 sg13g2_fill_1 FILLER_36_118 ();
 sg13g2_decap_8 FILLER_36_145 ();
 sg13g2_fill_1 FILLER_36_152 ();
 sg13g2_fill_1 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_197 ();
 sg13g2_decap_8 FILLER_36_204 ();
 sg13g2_fill_2 FILLER_36_211 ();
 sg13g2_fill_2 FILLER_36_217 ();
 sg13g2_fill_1 FILLER_36_219 ();
 sg13g2_fill_2 FILLER_36_273 ();
 sg13g2_fill_2 FILLER_36_305 ();
 sg13g2_fill_2 FILLER_36_337 ();
 sg13g2_fill_1 FILLER_36_370 ();
 sg13g2_fill_2 FILLER_36_405 ();
 sg13g2_fill_2 FILLER_36_417 ();
 sg13g2_fill_1 FILLER_36_419 ();
 sg13g2_fill_2 FILLER_36_425 ();
 sg13g2_fill_1 FILLER_36_456 ();
 sg13g2_fill_2 FILLER_36_463 ();
 sg13g2_decap_4 FILLER_36_494 ();
 sg13g2_fill_2 FILLER_36_498 ();
 sg13g2_decap_8 FILLER_36_521 ();
 sg13g2_fill_1 FILLER_36_528 ();
 sg13g2_fill_2 FILLER_36_535 ();
 sg13g2_fill_2 FILLER_36_593 ();
 sg13g2_fill_1 FILLER_36_595 ();
 sg13g2_fill_1 FILLER_36_608 ();
 sg13g2_fill_2 FILLER_36_627 ();
 sg13g2_fill_1 FILLER_36_653 ();
 sg13g2_decap_8 FILLER_36_674 ();
 sg13g2_decap_8 FILLER_36_681 ();
 sg13g2_decap_8 FILLER_36_688 ();
 sg13g2_decap_8 FILLER_36_695 ();
 sg13g2_decap_8 FILLER_36_702 ();
 sg13g2_decap_8 FILLER_36_709 ();
 sg13g2_decap_8 FILLER_36_716 ();
 sg13g2_decap_8 FILLER_36_723 ();
 sg13g2_decap_8 FILLER_36_730 ();
 sg13g2_decap_8 FILLER_36_737 ();
 sg13g2_decap_8 FILLER_36_744 ();
 sg13g2_decap_8 FILLER_36_751 ();
 sg13g2_decap_8 FILLER_36_758 ();
 sg13g2_decap_8 FILLER_36_765 ();
 sg13g2_decap_8 FILLER_36_772 ();
 sg13g2_decap_8 FILLER_36_779 ();
 sg13g2_decap_8 FILLER_36_786 ();
 sg13g2_decap_8 FILLER_36_793 ();
 sg13g2_decap_8 FILLER_36_800 ();
 sg13g2_decap_8 FILLER_36_807 ();
 sg13g2_decap_8 FILLER_36_814 ();
 sg13g2_decap_8 FILLER_36_821 ();
 sg13g2_decap_8 FILLER_36_828 ();
 sg13g2_decap_8 FILLER_36_835 ();
 sg13g2_decap_8 FILLER_36_842 ();
 sg13g2_decap_8 FILLER_36_849 ();
 sg13g2_decap_4 FILLER_36_856 ();
 sg13g2_fill_2 FILLER_36_860 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_4 FILLER_37_35 ();
 sg13g2_fill_2 FILLER_37_61 ();
 sg13g2_fill_1 FILLER_37_63 ();
 sg13g2_fill_2 FILLER_37_81 ();
 sg13g2_decap_8 FILLER_37_100 ();
 sg13g2_decap_4 FILLER_37_107 ();
 sg13g2_fill_1 FILLER_37_111 ();
 sg13g2_fill_1 FILLER_37_119 ();
 sg13g2_fill_2 FILLER_37_156 ();
 sg13g2_fill_1 FILLER_37_158 ();
 sg13g2_decap_4 FILLER_37_176 ();
 sg13g2_fill_2 FILLER_37_195 ();
 sg13g2_fill_2 FILLER_37_228 ();
 sg13g2_fill_1 FILLER_37_230 ();
 sg13g2_fill_2 FILLER_37_275 ();
 sg13g2_decap_8 FILLER_37_341 ();
 sg13g2_decap_8 FILLER_37_348 ();
 sg13g2_decap_4 FILLER_37_359 ();
 sg13g2_fill_2 FILLER_37_378 ();
 sg13g2_fill_2 FILLER_37_390 ();
 sg13g2_fill_1 FILLER_37_392 ();
 sg13g2_fill_1 FILLER_37_402 ();
 sg13g2_fill_2 FILLER_37_421 ();
 sg13g2_fill_2 FILLER_37_427 ();
 sg13g2_decap_8 FILLER_37_442 ();
 sg13g2_decap_8 FILLER_37_449 ();
 sg13g2_fill_1 FILLER_37_456 ();
 sg13g2_fill_2 FILLER_37_463 ();
 sg13g2_fill_1 FILLER_37_465 ();
 sg13g2_decap_4 FILLER_37_469 ();
 sg13g2_fill_2 FILLER_37_480 ();
 sg13g2_fill_1 FILLER_37_482 ();
 sg13g2_fill_1 FILLER_37_505 ();
 sg13g2_decap_4 FILLER_37_517 ();
 sg13g2_fill_1 FILLER_37_521 ();
 sg13g2_decap_8 FILLER_37_538 ();
 sg13g2_decap_8 FILLER_37_545 ();
 sg13g2_decap_8 FILLER_37_552 ();
 sg13g2_decap_4 FILLER_37_559 ();
 sg13g2_decap_8 FILLER_37_581 ();
 sg13g2_decap_8 FILLER_37_588 ();
 sg13g2_fill_1 FILLER_37_603 ();
 sg13g2_fill_1 FILLER_37_609 ();
 sg13g2_fill_2 FILLER_37_615 ();
 sg13g2_fill_1 FILLER_37_617 ();
 sg13g2_decap_4 FILLER_37_626 ();
 sg13g2_fill_2 FILLER_37_630 ();
 sg13g2_fill_1 FILLER_37_637 ();
 sg13g2_fill_1 FILLER_37_643 ();
 sg13g2_fill_2 FILLER_37_649 ();
 sg13g2_fill_1 FILLER_37_651 ();
 sg13g2_fill_2 FILLER_37_662 ();
 sg13g2_fill_1 FILLER_37_664 ();
 sg13g2_decap_8 FILLER_37_670 ();
 sg13g2_decap_8 FILLER_37_677 ();
 sg13g2_decap_8 FILLER_37_684 ();
 sg13g2_decap_8 FILLER_37_691 ();
 sg13g2_decap_8 FILLER_37_698 ();
 sg13g2_decap_8 FILLER_37_705 ();
 sg13g2_decap_8 FILLER_37_712 ();
 sg13g2_decap_8 FILLER_37_719 ();
 sg13g2_decap_8 FILLER_37_726 ();
 sg13g2_decap_8 FILLER_37_733 ();
 sg13g2_decap_8 FILLER_37_740 ();
 sg13g2_decap_8 FILLER_37_747 ();
 sg13g2_decap_8 FILLER_37_754 ();
 sg13g2_decap_8 FILLER_37_761 ();
 sg13g2_decap_8 FILLER_37_768 ();
 sg13g2_decap_8 FILLER_37_775 ();
 sg13g2_decap_8 FILLER_37_782 ();
 sg13g2_decap_8 FILLER_37_789 ();
 sg13g2_decap_8 FILLER_37_796 ();
 sg13g2_decap_8 FILLER_37_803 ();
 sg13g2_decap_8 FILLER_37_810 ();
 sg13g2_decap_8 FILLER_37_817 ();
 sg13g2_decap_8 FILLER_37_824 ();
 sg13g2_decap_8 FILLER_37_831 ();
 sg13g2_decap_8 FILLER_37_838 ();
 sg13g2_decap_8 FILLER_37_845 ();
 sg13g2_decap_8 FILLER_37_852 ();
 sg13g2_fill_2 FILLER_37_859 ();
 sg13g2_fill_1 FILLER_37_861 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_4 ();
 sg13g2_fill_2 FILLER_38_32 ();
 sg13g2_fill_2 FILLER_38_69 ();
 sg13g2_fill_1 FILLER_38_71 ();
 sg13g2_fill_2 FILLER_38_97 ();
 sg13g2_fill_1 FILLER_38_99 ();
 sg13g2_decap_8 FILLER_38_120 ();
 sg13g2_fill_1 FILLER_38_127 ();
 sg13g2_fill_2 FILLER_38_160 ();
 sg13g2_fill_2 FILLER_38_177 ();
 sg13g2_fill_2 FILLER_38_199 ();
 sg13g2_decap_8 FILLER_38_204 ();
 sg13g2_fill_2 FILLER_38_211 ();
 sg13g2_fill_2 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_223 ();
 sg13g2_fill_2 FILLER_38_239 ();
 sg13g2_fill_2 FILLER_38_254 ();
 sg13g2_fill_1 FILLER_38_261 ();
 sg13g2_fill_2 FILLER_38_272 ();
 sg13g2_decap_8 FILLER_38_345 ();
 sg13g2_decap_4 FILLER_38_352 ();
 sg13g2_fill_1 FILLER_38_385 ();
 sg13g2_fill_1 FILLER_38_395 ();
 sg13g2_fill_2 FILLER_38_404 ();
 sg13g2_fill_1 FILLER_38_406 ();
 sg13g2_decap_4 FILLER_38_431 ();
 sg13g2_fill_2 FILLER_38_435 ();
 sg13g2_fill_1 FILLER_38_446 ();
 sg13g2_fill_1 FILLER_38_467 ();
 sg13g2_fill_2 FILLER_38_476 ();
 sg13g2_fill_1 FILLER_38_478 ();
 sg13g2_decap_8 FILLER_38_483 ();
 sg13g2_decap_8 FILLER_38_490 ();
 sg13g2_fill_2 FILLER_38_497 ();
 sg13g2_fill_1 FILLER_38_503 ();
 sg13g2_fill_2 FILLER_38_519 ();
 sg13g2_fill_1 FILLER_38_521 ();
 sg13g2_fill_2 FILLER_38_527 ();
 sg13g2_fill_2 FILLER_38_537 ();
 sg13g2_fill_1 FILLER_38_539 ();
 sg13g2_fill_2 FILLER_38_576 ();
 sg13g2_fill_1 FILLER_38_578 ();
 sg13g2_decap_4 FILLER_38_593 ();
 sg13g2_fill_2 FILLER_38_597 ();
 sg13g2_fill_2 FILLER_38_607 ();
 sg13g2_fill_1 FILLER_38_609 ();
 sg13g2_fill_2 FILLER_38_626 ();
 sg13g2_fill_1 FILLER_38_636 ();
 sg13g2_fill_2 FILLER_38_644 ();
 sg13g2_fill_1 FILLER_38_646 ();
 sg13g2_fill_2 FILLER_38_655 ();
 sg13g2_fill_1 FILLER_38_657 ();
 sg13g2_decap_4 FILLER_38_663 ();
 sg13g2_fill_1 FILLER_38_667 ();
 sg13g2_decap_8 FILLER_38_676 ();
 sg13g2_decap_8 FILLER_38_683 ();
 sg13g2_decap_8 FILLER_38_690 ();
 sg13g2_decap_8 FILLER_38_697 ();
 sg13g2_decap_8 FILLER_38_704 ();
 sg13g2_decap_8 FILLER_38_711 ();
 sg13g2_decap_8 FILLER_38_718 ();
 sg13g2_decap_8 FILLER_38_725 ();
 sg13g2_decap_8 FILLER_38_732 ();
 sg13g2_decap_8 FILLER_38_739 ();
 sg13g2_decap_8 FILLER_38_746 ();
 sg13g2_decap_8 FILLER_38_753 ();
 sg13g2_decap_8 FILLER_38_760 ();
 sg13g2_decap_8 FILLER_38_767 ();
 sg13g2_decap_8 FILLER_38_774 ();
 sg13g2_decap_8 FILLER_38_781 ();
 sg13g2_decap_8 FILLER_38_788 ();
 sg13g2_decap_8 FILLER_38_795 ();
 sg13g2_decap_8 FILLER_38_802 ();
 sg13g2_decap_8 FILLER_38_809 ();
 sg13g2_decap_8 FILLER_38_816 ();
 sg13g2_decap_8 FILLER_38_823 ();
 sg13g2_decap_8 FILLER_38_830 ();
 sg13g2_decap_8 FILLER_38_837 ();
 sg13g2_decap_8 FILLER_38_844 ();
 sg13g2_decap_8 FILLER_38_851 ();
 sg13g2_decap_4 FILLER_38_858 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_4 ();
 sg13g2_decap_8 FILLER_39_36 ();
 sg13g2_fill_2 FILLER_39_43 ();
 sg13g2_fill_1 FILLER_39_45 ();
 sg13g2_decap_8 FILLER_39_66 ();
 sg13g2_decap_8 FILLER_39_73 ();
 sg13g2_fill_2 FILLER_39_80 ();
 sg13g2_fill_1 FILLER_39_82 ();
 sg13g2_decap_4 FILLER_39_94 ();
 sg13g2_fill_2 FILLER_39_98 ();
 sg13g2_fill_2 FILLER_39_124 ();
 sg13g2_fill_1 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_132 ();
 sg13g2_fill_2 FILLER_39_149 ();
 sg13g2_fill_2 FILLER_39_186 ();
 sg13g2_fill_2 FILLER_39_197 ();
 sg13g2_fill_1 FILLER_39_203 ();
 sg13g2_decap_4 FILLER_39_234 ();
 sg13g2_fill_2 FILLER_39_238 ();
 sg13g2_fill_1 FILLER_39_246 ();
 sg13g2_fill_2 FILLER_39_271 ();
 sg13g2_fill_1 FILLER_39_278 ();
 sg13g2_fill_2 FILLER_39_288 ();
 sg13g2_decap_8 FILLER_39_294 ();
 sg13g2_decap_8 FILLER_39_301 ();
 sg13g2_fill_2 FILLER_39_320 ();
 sg13g2_fill_1 FILLER_39_322 ();
 sg13g2_fill_2 FILLER_39_334 ();
 sg13g2_decap_4 FILLER_39_362 ();
 sg13g2_fill_2 FILLER_39_382 ();
 sg13g2_fill_1 FILLER_39_384 ();
 sg13g2_decap_8 FILLER_39_404 ();
 sg13g2_fill_2 FILLER_39_411 ();
 sg13g2_fill_2 FILLER_39_426 ();
 sg13g2_fill_2 FILLER_39_474 ();
 sg13g2_fill_1 FILLER_39_476 ();
 sg13g2_fill_1 FILLER_39_495 ();
 sg13g2_fill_2 FILLER_39_519 ();
 sg13g2_fill_1 FILLER_39_521 ();
 sg13g2_fill_2 FILLER_39_538 ();
 sg13g2_fill_2 FILLER_39_548 ();
 sg13g2_fill_2 FILLER_39_625 ();
 sg13g2_fill_2 FILLER_39_640 ();
 sg13g2_fill_2 FILLER_39_667 ();
 sg13g2_decap_8 FILLER_39_685 ();
 sg13g2_decap_4 FILLER_39_692 ();
 sg13g2_decap_8 FILLER_39_700 ();
 sg13g2_decap_8 FILLER_39_707 ();
 sg13g2_decap_8 FILLER_39_714 ();
 sg13g2_decap_8 FILLER_39_721 ();
 sg13g2_decap_8 FILLER_39_728 ();
 sg13g2_decap_8 FILLER_39_735 ();
 sg13g2_decap_8 FILLER_39_742 ();
 sg13g2_decap_8 FILLER_39_749 ();
 sg13g2_decap_8 FILLER_39_756 ();
 sg13g2_decap_8 FILLER_39_763 ();
 sg13g2_decap_8 FILLER_39_770 ();
 sg13g2_decap_8 FILLER_39_777 ();
 sg13g2_decap_8 FILLER_39_784 ();
 sg13g2_decap_8 FILLER_39_791 ();
 sg13g2_decap_8 FILLER_39_798 ();
 sg13g2_decap_8 FILLER_39_805 ();
 sg13g2_decap_8 FILLER_39_812 ();
 sg13g2_decap_8 FILLER_39_819 ();
 sg13g2_decap_8 FILLER_39_826 ();
 sg13g2_decap_8 FILLER_39_833 ();
 sg13g2_decap_8 FILLER_39_840 ();
 sg13g2_decap_8 FILLER_39_847 ();
 sg13g2_decap_8 FILLER_39_854 ();
 sg13g2_fill_1 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_7 ();
 sg13g2_decap_4 FILLER_40_12 ();
 sg13g2_fill_1 FILLER_40_16 ();
 sg13g2_fill_1 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_26 ();
 sg13g2_fill_1 FILLER_40_33 ();
 sg13g2_decap_8 FILLER_40_40 ();
 sg13g2_decap_4 FILLER_40_47 ();
 sg13g2_decap_8 FILLER_40_60 ();
 sg13g2_decap_4 FILLER_40_67 ();
 sg13g2_fill_1 FILLER_40_71 ();
 sg13g2_decap_8 FILLER_40_94 ();
 sg13g2_fill_2 FILLER_40_101 ();
 sg13g2_fill_1 FILLER_40_103 ();
 sg13g2_fill_2 FILLER_40_150 ();
 sg13g2_decap_8 FILLER_40_166 ();
 sg13g2_decap_4 FILLER_40_173 ();
 sg13g2_fill_1 FILLER_40_177 ();
 sg13g2_fill_2 FILLER_40_208 ();
 sg13g2_fill_1 FILLER_40_210 ();
 sg13g2_decap_8 FILLER_40_237 ();
 sg13g2_decap_8 FILLER_40_244 ();
 sg13g2_decap_4 FILLER_40_251 ();
 sg13g2_fill_1 FILLER_40_255 ();
 sg13g2_fill_2 FILLER_40_272 ();
 sg13g2_fill_1 FILLER_40_274 ();
 sg13g2_fill_2 FILLER_40_302 ();
 sg13g2_fill_1 FILLER_40_304 ();
 sg13g2_fill_1 FILLER_40_309 ();
 sg13g2_fill_1 FILLER_40_323 ();
 sg13g2_decap_8 FILLER_40_332 ();
 sg13g2_decap_8 FILLER_40_339 ();
 sg13g2_fill_1 FILLER_40_346 ();
 sg13g2_decap_8 FILLER_40_351 ();
 sg13g2_fill_1 FILLER_40_364 ();
 sg13g2_fill_1 FILLER_40_392 ();
 sg13g2_decap_8 FILLER_40_404 ();
 sg13g2_fill_2 FILLER_40_423 ();
 sg13g2_fill_1 FILLER_40_425 ();
 sg13g2_fill_2 FILLER_40_431 ();
 sg13g2_fill_1 FILLER_40_433 ();
 sg13g2_fill_1 FILLER_40_444 ();
 sg13g2_decap_8 FILLER_40_467 ();
 sg13g2_fill_1 FILLER_40_474 ();
 sg13g2_fill_2 FILLER_40_497 ();
 sg13g2_decap_4 FILLER_40_505 ();
 sg13g2_fill_2 FILLER_40_509 ();
 sg13g2_decap_8 FILLER_40_521 ();
 sg13g2_decap_4 FILLER_40_528 ();
 sg13g2_fill_2 FILLER_40_532 ();
 sg13g2_fill_2 FILLER_40_546 ();
 sg13g2_fill_2 FILLER_40_589 ();
 sg13g2_fill_1 FILLER_40_591 ();
 sg13g2_fill_2 FILLER_40_618 ();
 sg13g2_fill_1 FILLER_40_620 ();
 sg13g2_decap_4 FILLER_40_630 ();
 sg13g2_decap_4 FILLER_40_638 ();
 sg13g2_fill_1 FILLER_40_642 ();
 sg13g2_decap_8 FILLER_40_647 ();
 sg13g2_decap_8 FILLER_40_654 ();
 sg13g2_fill_1 FILLER_40_661 ();
 sg13g2_fill_2 FILLER_40_667 ();
 sg13g2_fill_1 FILLER_40_669 ();
 sg13g2_decap_8 FILLER_40_676 ();
 sg13g2_fill_2 FILLER_40_683 ();
 sg13g2_decap_8 FILLER_40_719 ();
 sg13g2_decap_4 FILLER_40_726 ();
 sg13g2_decap_8 FILLER_40_746 ();
 sg13g2_decap_8 FILLER_40_753 ();
 sg13g2_decap_8 FILLER_40_760 ();
 sg13g2_decap_8 FILLER_40_767 ();
 sg13g2_decap_8 FILLER_40_774 ();
 sg13g2_decap_8 FILLER_40_781 ();
 sg13g2_decap_8 FILLER_40_788 ();
 sg13g2_decap_8 FILLER_40_795 ();
 sg13g2_decap_8 FILLER_40_802 ();
 sg13g2_decap_8 FILLER_40_809 ();
 sg13g2_decap_8 FILLER_40_816 ();
 sg13g2_decap_8 FILLER_40_823 ();
 sg13g2_decap_8 FILLER_40_830 ();
 sg13g2_decap_8 FILLER_40_837 ();
 sg13g2_decap_8 FILLER_40_844 ();
 sg13g2_decap_8 FILLER_40_851 ();
 sg13g2_decap_4 FILLER_40_858 ();
 sg13g2_fill_2 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_2 ();
 sg13g2_decap_4 FILLER_41_37 ();
 sg13g2_decap_4 FILLER_41_71 ();
 sg13g2_fill_1 FILLER_41_75 ();
 sg13g2_fill_1 FILLER_41_97 ();
 sg13g2_decap_8 FILLER_41_129 ();
 sg13g2_fill_1 FILLER_41_146 ();
 sg13g2_fill_1 FILLER_41_152 ();
 sg13g2_fill_2 FILLER_41_163 ();
 sg13g2_fill_1 FILLER_41_165 ();
 sg13g2_fill_1 FILLER_41_180 ();
 sg13g2_decap_4 FILLER_41_217 ();
 sg13g2_fill_2 FILLER_41_236 ();
 sg13g2_fill_1 FILLER_41_238 ();
 sg13g2_fill_2 FILLER_41_250 ();
 sg13g2_fill_2 FILLER_41_265 ();
 sg13g2_decap_8 FILLER_41_286 ();
 sg13g2_fill_2 FILLER_41_306 ();
 sg13g2_fill_1 FILLER_41_333 ();
 sg13g2_decap_4 FILLER_41_349 ();
 sg13g2_decap_4 FILLER_41_379 ();
 sg13g2_fill_1 FILLER_41_414 ();
 sg13g2_fill_1 FILLER_41_484 ();
 sg13g2_fill_2 FILLER_41_495 ();
 sg13g2_fill_2 FILLER_41_505 ();
 sg13g2_fill_2 FILLER_41_520 ();
 sg13g2_fill_2 FILLER_41_532 ();
 sg13g2_fill_1 FILLER_41_558 ();
 sg13g2_fill_2 FILLER_41_611 ();
 sg13g2_fill_2 FILLER_41_618 ();
 sg13g2_fill_1 FILLER_41_620 ();
 sg13g2_fill_2 FILLER_41_629 ();
 sg13g2_fill_1 FILLER_41_655 ();
 sg13g2_decap_4 FILLER_41_694 ();
 sg13g2_decap_8 FILLER_41_708 ();
 sg13g2_decap_4 FILLER_41_715 ();
 sg13g2_decap_8 FILLER_41_745 ();
 sg13g2_decap_8 FILLER_41_752 ();
 sg13g2_decap_8 FILLER_41_759 ();
 sg13g2_decap_8 FILLER_41_766 ();
 sg13g2_decap_8 FILLER_41_773 ();
 sg13g2_decap_8 FILLER_41_780 ();
 sg13g2_decap_8 FILLER_41_787 ();
 sg13g2_decap_8 FILLER_41_794 ();
 sg13g2_decap_8 FILLER_41_801 ();
 sg13g2_decap_8 FILLER_41_808 ();
 sg13g2_decap_8 FILLER_41_815 ();
 sg13g2_decap_8 FILLER_41_822 ();
 sg13g2_decap_8 FILLER_41_829 ();
 sg13g2_decap_8 FILLER_41_836 ();
 sg13g2_decap_8 FILLER_41_843 ();
 sg13g2_decap_8 FILLER_41_850 ();
 sg13g2_decap_4 FILLER_41_857 ();
 sg13g2_fill_1 FILLER_41_861 ();
 sg13g2_decap_4 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_4 ();
 sg13g2_decap_4 FILLER_42_31 ();
 sg13g2_fill_1 FILLER_42_35 ();
 sg13g2_fill_2 FILLER_42_67 ();
 sg13g2_decap_8 FILLER_42_95 ();
 sg13g2_decap_4 FILLER_42_102 ();
 sg13g2_fill_1 FILLER_42_106 ();
 sg13g2_decap_8 FILLER_42_134 ();
 sg13g2_decap_4 FILLER_42_156 ();
 sg13g2_fill_1 FILLER_42_160 ();
 sg13g2_decap_8 FILLER_42_166 ();
 sg13g2_decap_8 FILLER_42_173 ();
 sg13g2_fill_2 FILLER_42_196 ();
 sg13g2_fill_2 FILLER_42_232 ();
 sg13g2_fill_1 FILLER_42_234 ();
 sg13g2_decap_4 FILLER_42_254 ();
 sg13g2_fill_1 FILLER_42_258 ();
 sg13g2_decap_8 FILLER_42_262 ();
 sg13g2_fill_2 FILLER_42_269 ();
 sg13g2_fill_1 FILLER_42_271 ();
 sg13g2_decap_4 FILLER_42_284 ();
 sg13g2_fill_2 FILLER_42_288 ();
 sg13g2_decap_8 FILLER_42_297 ();
 sg13g2_decap_8 FILLER_42_318 ();
 sg13g2_fill_1 FILLER_42_325 ();
 sg13g2_decap_8 FILLER_42_331 ();
 sg13g2_decap_8 FILLER_42_348 ();
 sg13g2_decap_8 FILLER_42_355 ();
 sg13g2_fill_1 FILLER_42_362 ();
 sg13g2_fill_1 FILLER_42_366 ();
 sg13g2_fill_1 FILLER_42_396 ();
 sg13g2_fill_2 FILLER_42_417 ();
 sg13g2_fill_1 FILLER_42_419 ();
 sg13g2_fill_1 FILLER_42_425 ();
 sg13g2_decap_8 FILLER_42_431 ();
 sg13g2_decap_4 FILLER_42_438 ();
 sg13g2_fill_2 FILLER_42_445 ();
 sg13g2_fill_1 FILLER_42_447 ();
 sg13g2_decap_4 FILLER_42_453 ();
 sg13g2_fill_2 FILLER_42_457 ();
 sg13g2_decap_8 FILLER_42_464 ();
 sg13g2_decap_4 FILLER_42_471 ();
 sg13g2_decap_8 FILLER_42_491 ();
 sg13g2_decap_4 FILLER_42_498 ();
 sg13g2_fill_2 FILLER_42_513 ();
 sg13g2_fill_1 FILLER_42_515 ();
 sg13g2_fill_1 FILLER_42_558 ();
 sg13g2_decap_4 FILLER_42_562 ();
 sg13g2_fill_1 FILLER_42_566 ();
 sg13g2_decap_4 FILLER_42_580 ();
 sg13g2_fill_1 FILLER_42_584 ();
 sg13g2_decap_8 FILLER_42_594 ();
 sg13g2_fill_1 FILLER_42_601 ();
 sg13g2_decap_8 FILLER_42_623 ();
 sg13g2_fill_2 FILLER_42_630 ();
 sg13g2_fill_1 FILLER_42_632 ();
 sg13g2_fill_2 FILLER_42_656 ();
 sg13g2_decap_4 FILLER_42_677 ();
 sg13g2_fill_2 FILLER_42_681 ();
 sg13g2_fill_1 FILLER_42_707 ();
 sg13g2_decap_4 FILLER_42_726 ();
 sg13g2_decap_8 FILLER_42_747 ();
 sg13g2_decap_8 FILLER_42_754 ();
 sg13g2_decap_8 FILLER_42_761 ();
 sg13g2_decap_8 FILLER_42_768 ();
 sg13g2_decap_8 FILLER_42_775 ();
 sg13g2_decap_8 FILLER_42_782 ();
 sg13g2_decap_8 FILLER_42_789 ();
 sg13g2_decap_8 FILLER_42_796 ();
 sg13g2_decap_8 FILLER_42_803 ();
 sg13g2_decap_8 FILLER_42_810 ();
 sg13g2_decap_8 FILLER_42_817 ();
 sg13g2_decap_8 FILLER_42_824 ();
 sg13g2_decap_8 FILLER_42_831 ();
 sg13g2_decap_8 FILLER_42_838 ();
 sg13g2_decap_8 FILLER_42_845 ();
 sg13g2_decap_8 FILLER_42_852 ();
 sg13g2_fill_2 FILLER_42_859 ();
 sg13g2_fill_1 FILLER_42_861 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_7 ();
 sg13g2_decap_4 FILLER_43_12 ();
 sg13g2_fill_2 FILLER_43_29 ();
 sg13g2_fill_1 FILLER_43_31 ();
 sg13g2_decap_8 FILLER_43_36 ();
 sg13g2_decap_4 FILLER_43_47 ();
 sg13g2_fill_1 FILLER_43_51 ();
 sg13g2_fill_2 FILLER_43_56 ();
 sg13g2_fill_2 FILLER_43_64 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_fill_2 FILLER_43_77 ();
 sg13g2_fill_1 FILLER_43_79 ();
 sg13g2_fill_1 FILLER_43_89 ();
 sg13g2_fill_2 FILLER_43_95 ();
 sg13g2_fill_1 FILLER_43_97 ();
 sg13g2_fill_1 FILLER_43_103 ();
 sg13g2_decap_4 FILLER_43_108 ();
 sg13g2_fill_2 FILLER_43_112 ();
 sg13g2_fill_2 FILLER_43_118 ();
 sg13g2_fill_1 FILLER_43_120 ();
 sg13g2_decap_4 FILLER_43_125 ();
 sg13g2_fill_2 FILLER_43_129 ();
 sg13g2_fill_1 FILLER_43_149 ();
 sg13g2_decap_4 FILLER_43_174 ();
 sg13g2_fill_1 FILLER_43_178 ();
 sg13g2_fill_1 FILLER_43_185 ();
 sg13g2_fill_2 FILLER_43_192 ();
 sg13g2_decap_4 FILLER_43_211 ();
 sg13g2_fill_2 FILLER_43_215 ();
 sg13g2_fill_2 FILLER_43_221 ();
 sg13g2_fill_1 FILLER_43_229 ();
 sg13g2_fill_2 FILLER_43_258 ();
 sg13g2_fill_2 FILLER_43_271 ();
 sg13g2_decap_4 FILLER_43_327 ();
 sg13g2_fill_1 FILLER_43_331 ();
 sg13g2_fill_1 FILLER_43_358 ();
 sg13g2_decap_8 FILLER_43_378 ();
 sg13g2_fill_1 FILLER_43_385 ();
 sg13g2_decap_8 FILLER_43_396 ();
 sg13g2_fill_1 FILLER_43_403 ();
 sg13g2_fill_1 FILLER_43_440 ();
 sg13g2_decap_8 FILLER_43_462 ();
 sg13g2_decap_4 FILLER_43_469 ();
 sg13g2_fill_2 FILLER_43_493 ();
 sg13g2_decap_4 FILLER_43_517 ();
 sg13g2_decap_8 FILLER_43_530 ();
 sg13g2_fill_1 FILLER_43_537 ();
 sg13g2_fill_1 FILLER_43_563 ();
 sg13g2_decap_4 FILLER_43_569 ();
 sg13g2_fill_2 FILLER_43_604 ();
 sg13g2_decap_4 FILLER_43_610 ();
 sg13g2_fill_1 FILLER_43_614 ();
 sg13g2_decap_4 FILLER_43_627 ();
 sg13g2_decap_4 FILLER_43_636 ();
 sg13g2_decap_4 FILLER_43_654 ();
 sg13g2_fill_2 FILLER_43_666 ();
 sg13g2_fill_1 FILLER_43_668 ();
 sg13g2_decap_8 FILLER_43_686 ();
 sg13g2_fill_2 FILLER_43_705 ();
 sg13g2_fill_2 FILLER_43_723 ();
 sg13g2_fill_1 FILLER_43_732 ();
 sg13g2_decap_8 FILLER_43_754 ();
 sg13g2_decap_8 FILLER_43_761 ();
 sg13g2_decap_8 FILLER_43_768 ();
 sg13g2_decap_8 FILLER_43_775 ();
 sg13g2_decap_8 FILLER_43_782 ();
 sg13g2_decap_8 FILLER_43_789 ();
 sg13g2_decap_8 FILLER_43_796 ();
 sg13g2_decap_8 FILLER_43_803 ();
 sg13g2_decap_8 FILLER_43_810 ();
 sg13g2_decap_8 FILLER_43_817 ();
 sg13g2_decap_8 FILLER_43_824 ();
 sg13g2_decap_8 FILLER_43_831 ();
 sg13g2_decap_8 FILLER_43_838 ();
 sg13g2_decap_8 FILLER_43_845 ();
 sg13g2_decap_8 FILLER_43_852 ();
 sg13g2_fill_2 FILLER_43_859 ();
 sg13g2_fill_1 FILLER_43_861 ();
 sg13g2_fill_1 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_31 ();
 sg13g2_fill_1 FILLER_44_33 ();
 sg13g2_decap_4 FILLER_44_64 ();
 sg13g2_fill_1 FILLER_44_102 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_fill_2 FILLER_44_140 ();
 sg13g2_decap_4 FILLER_44_168 ();
 sg13g2_decap_8 FILLER_44_189 ();
 sg13g2_fill_2 FILLER_44_196 ();
 sg13g2_decap_8 FILLER_44_202 ();
 sg13g2_decap_4 FILLER_44_209 ();
 sg13g2_decap_8 FILLER_44_217 ();
 sg13g2_fill_1 FILLER_44_224 ();
 sg13g2_fill_2 FILLER_44_235 ();
 sg13g2_fill_1 FILLER_44_237 ();
 sg13g2_fill_2 FILLER_44_243 ();
 sg13g2_decap_4 FILLER_44_249 ();
 sg13g2_fill_2 FILLER_44_253 ();
 sg13g2_fill_1 FILLER_44_268 ();
 sg13g2_decap_8 FILLER_44_287 ();
 sg13g2_decap_4 FILLER_44_294 ();
 sg13g2_fill_1 FILLER_44_298 ();
 sg13g2_decap_4 FILLER_44_304 ();
 sg13g2_fill_2 FILLER_44_308 ();
 sg13g2_fill_1 FILLER_44_315 ();
 sg13g2_decap_8 FILLER_44_320 ();
 sg13g2_decap_8 FILLER_44_327 ();
 sg13g2_fill_1 FILLER_44_351 ();
 sg13g2_decap_4 FILLER_44_357 ();
 sg13g2_fill_1 FILLER_44_390 ();
 sg13g2_fill_2 FILLER_44_403 ();
 sg13g2_fill_1 FILLER_44_405 ();
 sg13g2_decap_8 FILLER_44_435 ();
 sg13g2_fill_1 FILLER_44_442 ();
 sg13g2_decap_8 FILLER_44_489 ();
 sg13g2_decap_8 FILLER_44_514 ();
 sg13g2_decap_8 FILLER_44_521 ();
 sg13g2_fill_1 FILLER_44_540 ();
 sg13g2_fill_1 FILLER_44_549 ();
 sg13g2_decap_4 FILLER_44_555 ();
 sg13g2_fill_1 FILLER_44_589 ();
 sg13g2_decap_8 FILLER_44_598 ();
 sg13g2_fill_2 FILLER_44_605 ();
 sg13g2_fill_1 FILLER_44_607 ();
 sg13g2_fill_1 FILLER_44_625 ();
 sg13g2_decap_4 FILLER_44_655 ();
 sg13g2_fill_1 FILLER_44_693 ();
 sg13g2_fill_2 FILLER_44_699 ();
 sg13g2_fill_1 FILLER_44_701 ();
 sg13g2_fill_2 FILLER_44_712 ();
 sg13g2_fill_1 FILLER_44_714 ();
 sg13g2_fill_2 FILLER_44_720 ();
 sg13g2_fill_1 FILLER_44_722 ();
 sg13g2_decap_8 FILLER_44_728 ();
 sg13g2_decap_8 FILLER_44_761 ();
 sg13g2_decap_8 FILLER_44_768 ();
 sg13g2_decap_8 FILLER_44_775 ();
 sg13g2_decap_8 FILLER_44_782 ();
 sg13g2_decap_8 FILLER_44_789 ();
 sg13g2_decap_8 FILLER_44_796 ();
 sg13g2_decap_8 FILLER_44_803 ();
 sg13g2_decap_8 FILLER_44_810 ();
 sg13g2_decap_8 FILLER_44_817 ();
 sg13g2_decap_8 FILLER_44_824 ();
 sg13g2_decap_8 FILLER_44_831 ();
 sg13g2_decap_8 FILLER_44_838 ();
 sg13g2_decap_8 FILLER_44_845 ();
 sg13g2_decap_8 FILLER_44_852 ();
 sg13g2_fill_2 FILLER_44_859 ();
 sg13g2_fill_1 FILLER_44_861 ();
 sg13g2_fill_2 FILLER_45_26 ();
 sg13g2_fill_1 FILLER_45_28 ();
 sg13g2_fill_1 FILLER_45_33 ();
 sg13g2_decap_4 FILLER_45_39 ();
 sg13g2_fill_1 FILLER_45_43 ();
 sg13g2_fill_1 FILLER_45_48 ();
 sg13g2_fill_1 FILLER_45_62 ();
 sg13g2_fill_2 FILLER_45_77 ();
 sg13g2_fill_2 FILLER_45_83 ();
 sg13g2_fill_1 FILLER_45_111 ();
 sg13g2_fill_1 FILLER_45_126 ();
 sg13g2_decap_4 FILLER_45_141 ();
 sg13g2_fill_2 FILLER_45_150 ();
 sg13g2_fill_1 FILLER_45_172 ();
 sg13g2_fill_1 FILLER_45_201 ();
 sg13g2_decap_4 FILLER_45_243 ();
 sg13g2_fill_1 FILLER_45_247 ();
 sg13g2_fill_2 FILLER_45_254 ();
 sg13g2_fill_1 FILLER_45_256 ();
 sg13g2_decap_8 FILLER_45_265 ();
 sg13g2_decap_8 FILLER_45_272 ();
 sg13g2_fill_1 FILLER_45_279 ();
 sg13g2_decap_4 FILLER_45_285 ();
 sg13g2_fill_2 FILLER_45_289 ();
 sg13g2_decap_8 FILLER_45_310 ();
 sg13g2_fill_1 FILLER_45_317 ();
 sg13g2_fill_2 FILLER_45_330 ();
 sg13g2_fill_1 FILLER_45_332 ();
 sg13g2_decap_4 FILLER_45_337 ();
 sg13g2_fill_2 FILLER_45_341 ();
 sg13g2_fill_2 FILLER_45_347 ();
 sg13g2_decap_8 FILLER_45_357 ();
 sg13g2_decap_8 FILLER_45_364 ();
 sg13g2_decap_4 FILLER_45_371 ();
 sg13g2_decap_8 FILLER_45_398 ();
 sg13g2_fill_1 FILLER_45_405 ();
 sg13g2_decap_8 FILLER_45_418 ();
 sg13g2_decap_8 FILLER_45_451 ();
 sg13g2_fill_2 FILLER_45_458 ();
 sg13g2_fill_1 FILLER_45_460 ();
 sg13g2_decap_8 FILLER_45_466 ();
 sg13g2_fill_2 FILLER_45_483 ();
 sg13g2_fill_2 FILLER_45_502 ();
 sg13g2_decap_4 FILLER_45_517 ();
 sg13g2_fill_2 FILLER_45_521 ();
 sg13g2_fill_1 FILLER_45_532 ();
 sg13g2_fill_1 FILLER_45_547 ();
 sg13g2_fill_2 FILLER_45_580 ();
 sg13g2_decap_4 FILLER_45_611 ();
 sg13g2_fill_1 FILLER_45_615 ();
 sg13g2_fill_1 FILLER_45_627 ();
 sg13g2_decap_4 FILLER_45_636 ();
 sg13g2_fill_2 FILLER_45_640 ();
 sg13g2_decap_4 FILLER_45_647 ();
 sg13g2_fill_2 FILLER_45_669 ();
 sg13g2_decap_8 FILLER_45_675 ();
 sg13g2_decap_4 FILLER_45_682 ();
 sg13g2_fill_2 FILLER_45_686 ();
 sg13g2_decap_4 FILLER_45_706 ();
 sg13g2_decap_4 FILLER_45_720 ();
 sg13g2_decap_8 FILLER_45_759 ();
 sg13g2_decap_8 FILLER_45_766 ();
 sg13g2_decap_8 FILLER_45_773 ();
 sg13g2_decap_8 FILLER_45_780 ();
 sg13g2_decap_8 FILLER_45_787 ();
 sg13g2_decap_8 FILLER_45_794 ();
 sg13g2_decap_8 FILLER_45_801 ();
 sg13g2_decap_8 FILLER_45_808 ();
 sg13g2_decap_8 FILLER_45_815 ();
 sg13g2_decap_8 FILLER_45_822 ();
 sg13g2_decap_8 FILLER_45_829 ();
 sg13g2_decap_8 FILLER_45_836 ();
 sg13g2_decap_8 FILLER_45_843 ();
 sg13g2_decap_8 FILLER_45_850 ();
 sg13g2_decap_4 FILLER_45_857 ();
 sg13g2_fill_1 FILLER_45_861 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_7 ();
 sg13g2_fill_1 FILLER_46_46 ();
 sg13g2_fill_1 FILLER_46_63 ();
 sg13g2_fill_2 FILLER_46_100 ();
 sg13g2_fill_2 FILLER_46_108 ();
 sg13g2_fill_1 FILLER_46_110 ();
 sg13g2_fill_1 FILLER_46_116 ();
 sg13g2_decap_8 FILLER_46_143 ();
 sg13g2_decap_4 FILLER_46_150 ();
 sg13g2_fill_2 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_166 ();
 sg13g2_decap_4 FILLER_46_173 ();
 sg13g2_fill_1 FILLER_46_177 ();
 sg13g2_decap_8 FILLER_46_205 ();
 sg13g2_decap_8 FILLER_46_212 ();
 sg13g2_fill_2 FILLER_46_219 ();
 sg13g2_fill_2 FILLER_46_256 ();
 sg13g2_fill_1 FILLER_46_258 ();
 sg13g2_fill_2 FILLER_46_264 ();
 sg13g2_fill_1 FILLER_46_266 ();
 sg13g2_fill_2 FILLER_46_272 ();
 sg13g2_decap_8 FILLER_46_280 ();
 sg13g2_fill_2 FILLER_46_330 ();
 sg13g2_fill_1 FILLER_46_332 ();
 sg13g2_decap_4 FILLER_46_347 ();
 sg13g2_fill_2 FILLER_46_361 ();
 sg13g2_fill_1 FILLER_46_363 ();
 sg13g2_decap_4 FILLER_46_381 ();
 sg13g2_fill_2 FILLER_46_385 ();
 sg13g2_fill_2 FILLER_46_392 ();
 sg13g2_fill_1 FILLER_46_394 ();
 sg13g2_fill_2 FILLER_46_434 ();
 sg13g2_fill_2 FILLER_46_440 ();
 sg13g2_fill_2 FILLER_46_491 ();
 sg13g2_fill_1 FILLER_46_516 ();
 sg13g2_fill_2 FILLER_46_546 ();
 sg13g2_fill_1 FILLER_46_548 ();
 sg13g2_fill_2 FILLER_46_575 ();
 sg13g2_fill_1 FILLER_46_577 ();
 sg13g2_fill_1 FILLER_46_583 ();
 sg13g2_decap_4 FILLER_46_589 ();
 sg13g2_fill_1 FILLER_46_593 ();
 sg13g2_decap_4 FILLER_46_628 ();
 sg13g2_fill_1 FILLER_46_632 ();
 sg13g2_fill_1 FILLER_46_659 ();
 sg13g2_decap_8 FILLER_46_703 ();
 sg13g2_decap_4 FILLER_46_715 ();
 sg13g2_fill_2 FILLER_46_724 ();
 sg13g2_fill_1 FILLER_46_726 ();
 sg13g2_fill_1 FILLER_46_732 ();
 sg13g2_fill_2 FILLER_46_738 ();
 sg13g2_decap_8 FILLER_46_765 ();
 sg13g2_decap_8 FILLER_46_772 ();
 sg13g2_decap_8 FILLER_46_779 ();
 sg13g2_decap_8 FILLER_46_786 ();
 sg13g2_decap_8 FILLER_46_793 ();
 sg13g2_decap_8 FILLER_46_800 ();
 sg13g2_decap_8 FILLER_46_807 ();
 sg13g2_decap_8 FILLER_46_814 ();
 sg13g2_decap_8 FILLER_46_821 ();
 sg13g2_decap_8 FILLER_46_828 ();
 sg13g2_decap_8 FILLER_46_835 ();
 sg13g2_decap_8 FILLER_46_842 ();
 sg13g2_decap_8 FILLER_46_849 ();
 sg13g2_decap_4 FILLER_46_856 ();
 sg13g2_fill_2 FILLER_46_860 ();
 sg13g2_fill_2 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_41 ();
 sg13g2_fill_2 FILLER_47_65 ();
 sg13g2_fill_1 FILLER_47_99 ();
 sg13g2_fill_2 FILLER_47_116 ();
 sg13g2_decap_4 FILLER_47_124 ();
 sg13g2_fill_1 FILLER_47_132 ();
 sg13g2_fill_2 FILLER_47_138 ();
 sg13g2_fill_1 FILLER_47_154 ();
 sg13g2_fill_1 FILLER_47_160 ();
 sg13g2_decap_8 FILLER_47_175 ();
 sg13g2_decap_4 FILLER_47_182 ();
 sg13g2_fill_1 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_201 ();
 sg13g2_fill_2 FILLER_47_224 ();
 sg13g2_fill_1 FILLER_47_226 ();
 sg13g2_fill_2 FILLER_47_249 ();
 sg13g2_fill_2 FILLER_47_274 ();
 sg13g2_fill_1 FILLER_47_276 ();
 sg13g2_fill_1 FILLER_47_292 ();
 sg13g2_fill_1 FILLER_47_344 ();
 sg13g2_decap_4 FILLER_47_373 ();
 sg13g2_fill_2 FILLER_47_377 ();
 sg13g2_decap_4 FILLER_47_392 ();
 sg13g2_fill_1 FILLER_47_396 ();
 sg13g2_fill_2 FILLER_47_404 ();
 sg13g2_fill_1 FILLER_47_406 ();
 sg13g2_fill_2 FILLER_47_412 ();
 sg13g2_fill_1 FILLER_47_430 ();
 sg13g2_fill_1 FILLER_47_446 ();
 sg13g2_fill_1 FILLER_47_456 ();
 sg13g2_decap_8 FILLER_47_492 ();
 sg13g2_fill_2 FILLER_47_499 ();
 sg13g2_decap_8 FILLER_47_517 ();
 sg13g2_fill_1 FILLER_47_527 ();
 sg13g2_fill_2 FILLER_47_537 ();
 sg13g2_fill_1 FILLER_47_539 ();
 sg13g2_fill_2 FILLER_47_562 ();
 sg13g2_fill_2 FILLER_47_580 ();
 sg13g2_fill_1 FILLER_47_582 ();
 sg13g2_decap_8 FILLER_47_603 ();
 sg13g2_decap_8 FILLER_47_610 ();
 sg13g2_decap_8 FILLER_47_617 ();
 sg13g2_fill_2 FILLER_47_624 ();
 sg13g2_decap_8 FILLER_47_658 ();
 sg13g2_fill_1 FILLER_47_665 ();
 sg13g2_decap_8 FILLER_47_709 ();
 sg13g2_fill_2 FILLER_47_720 ();
 sg13g2_decap_8 FILLER_47_776 ();
 sg13g2_decap_8 FILLER_47_783 ();
 sg13g2_decap_8 FILLER_47_790 ();
 sg13g2_decap_8 FILLER_47_797 ();
 sg13g2_decap_8 FILLER_47_804 ();
 sg13g2_decap_8 FILLER_47_811 ();
 sg13g2_decap_8 FILLER_47_818 ();
 sg13g2_decap_8 FILLER_47_825 ();
 sg13g2_decap_8 FILLER_47_832 ();
 sg13g2_decap_8 FILLER_47_839 ();
 sg13g2_decap_8 FILLER_47_846 ();
 sg13g2_decap_8 FILLER_47_853 ();
 sg13g2_fill_2 FILLER_47_860 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_37 ();
 sg13g2_fill_2 FILLER_48_80 ();
 sg13g2_fill_2 FILLER_48_107 ();
 sg13g2_decap_4 FILLER_48_114 ();
 sg13g2_fill_2 FILLER_48_118 ();
 sg13g2_fill_2 FILLER_48_129 ();
 sg13g2_fill_1 FILLER_48_131 ();
 sg13g2_decap_8 FILLER_48_141 ();
 sg13g2_decap_8 FILLER_48_176 ();
 sg13g2_decap_4 FILLER_48_183 ();
 sg13g2_fill_2 FILLER_48_210 ();
 sg13g2_decap_4 FILLER_48_225 ();
 sg13g2_fill_1 FILLER_48_229 ();
 sg13g2_decap_8 FILLER_48_248 ();
 sg13g2_decap_4 FILLER_48_255 ();
 sg13g2_decap_4 FILLER_48_269 ();
 sg13g2_decap_8 FILLER_48_277 ();
 sg13g2_decap_4 FILLER_48_284 ();
 sg13g2_fill_1 FILLER_48_288 ();
 sg13g2_decap_4 FILLER_48_298 ();
 sg13g2_decap_4 FILLER_48_307 ();
 sg13g2_fill_1 FILLER_48_311 ();
 sg13g2_decap_4 FILLER_48_325 ();
 sg13g2_fill_2 FILLER_48_347 ();
 sg13g2_fill_1 FILLER_48_354 ();
 sg13g2_decap_8 FILLER_48_359 ();
 sg13g2_decap_4 FILLER_48_371 ();
 sg13g2_fill_1 FILLER_48_375 ();
 sg13g2_decap_8 FILLER_48_400 ();
 sg13g2_decap_4 FILLER_48_407 ();
 sg13g2_fill_2 FILLER_48_411 ();
 sg13g2_decap_4 FILLER_48_434 ();
 sg13g2_fill_2 FILLER_48_438 ();
 sg13g2_decap_8 FILLER_48_465 ();
 sg13g2_decap_8 FILLER_48_472 ();
 sg13g2_fill_2 FILLER_48_479 ();
 sg13g2_decap_4 FILLER_48_530 ();
 sg13g2_fill_1 FILLER_48_534 ();
 sg13g2_fill_2 FILLER_48_572 ();
 sg13g2_decap_4 FILLER_48_584 ();
 sg13g2_fill_1 FILLER_48_588 ();
 sg13g2_fill_2 FILLER_48_593 ();
 sg13g2_fill_1 FILLER_48_595 ();
 sg13g2_decap_4 FILLER_48_602 ();
 sg13g2_decap_8 FILLER_48_623 ();
 sg13g2_fill_1 FILLER_48_630 ();
 sg13g2_fill_1 FILLER_48_646 ();
 sg13g2_fill_1 FILLER_48_653 ();
 sg13g2_decap_8 FILLER_48_667 ();
 sg13g2_fill_2 FILLER_48_682 ();
 sg13g2_fill_1 FILLER_48_684 ();
 sg13g2_fill_2 FILLER_48_696 ();
 sg13g2_fill_2 FILLER_48_703 ();
 sg13g2_fill_2 FILLER_48_736 ();
 sg13g2_decap_8 FILLER_48_766 ();
 sg13g2_decap_8 FILLER_48_773 ();
 sg13g2_decap_8 FILLER_48_780 ();
 sg13g2_decap_8 FILLER_48_787 ();
 sg13g2_decap_8 FILLER_48_794 ();
 sg13g2_decap_8 FILLER_48_801 ();
 sg13g2_decap_8 FILLER_48_808 ();
 sg13g2_decap_8 FILLER_48_815 ();
 sg13g2_decap_8 FILLER_48_822 ();
 sg13g2_decap_8 FILLER_48_829 ();
 sg13g2_decap_8 FILLER_48_836 ();
 sg13g2_decap_8 FILLER_48_843 ();
 sg13g2_decap_8 FILLER_48_850 ();
 sg13g2_decap_4 FILLER_48_857 ();
 sg13g2_fill_1 FILLER_48_861 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_7 ();
 sg13g2_fill_2 FILLER_49_80 ();
 sg13g2_fill_1 FILLER_49_87 ();
 sg13g2_fill_2 FILLER_49_109 ();
 sg13g2_fill_1 FILLER_49_111 ();
 sg13g2_decap_4 FILLER_49_146 ();
 sg13g2_decap_8 FILLER_49_167 ();
 sg13g2_decap_4 FILLER_49_174 ();
 sg13g2_fill_2 FILLER_49_178 ();
 sg13g2_decap_8 FILLER_49_184 ();
 sg13g2_decap_8 FILLER_49_204 ();
 sg13g2_fill_2 FILLER_49_211 ();
 sg13g2_fill_1 FILLER_49_213 ();
 sg13g2_decap_8 FILLER_49_220 ();
 sg13g2_decap_8 FILLER_49_227 ();
 sg13g2_decap_8 FILLER_49_234 ();
 sg13g2_fill_1 FILLER_49_241 ();
 sg13g2_fill_2 FILLER_49_279 ();
 sg13g2_decap_4 FILLER_49_304 ();
 sg13g2_fill_2 FILLER_49_308 ();
 sg13g2_fill_2 FILLER_49_323 ();
 sg13g2_fill_2 FILLER_49_340 ();
 sg13g2_fill_1 FILLER_49_342 ();
 sg13g2_fill_1 FILLER_49_383 ();
 sg13g2_fill_2 FILLER_49_403 ();
 sg13g2_decap_8 FILLER_49_415 ();
 sg13g2_fill_1 FILLER_49_422 ();
 sg13g2_fill_2 FILLER_49_428 ();
 sg13g2_fill_1 FILLER_49_430 ();
 sg13g2_fill_1 FILLER_49_439 ();
 sg13g2_fill_2 FILLER_49_465 ();
 sg13g2_fill_1 FILLER_49_467 ();
 sg13g2_fill_1 FILLER_49_472 ();
 sg13g2_decap_4 FILLER_49_477 ();
 sg13g2_fill_1 FILLER_49_487 ();
 sg13g2_decap_8 FILLER_49_503 ();
 sg13g2_fill_1 FILLER_49_510 ();
 sg13g2_decap_8 FILLER_49_539 ();
 sg13g2_decap_8 FILLER_49_546 ();
 sg13g2_decap_8 FILLER_49_556 ();
 sg13g2_decap_4 FILLER_49_563 ();
 sg13g2_fill_1 FILLER_49_591 ();
 sg13g2_fill_2 FILLER_49_605 ();
 sg13g2_fill_1 FILLER_49_607 ();
 sg13g2_fill_1 FILLER_49_620 ();
 sg13g2_fill_1 FILLER_49_647 ();
 sg13g2_fill_2 FILLER_49_668 ();
 sg13g2_fill_1 FILLER_49_670 ();
 sg13g2_fill_1 FILLER_49_679 ();
 sg13g2_fill_1 FILLER_49_685 ();
 sg13g2_fill_1 FILLER_49_704 ();
 sg13g2_fill_1 FILLER_49_721 ();
 sg13g2_decap_8 FILLER_49_778 ();
 sg13g2_decap_8 FILLER_49_785 ();
 sg13g2_decap_8 FILLER_49_792 ();
 sg13g2_decap_8 FILLER_49_799 ();
 sg13g2_decap_8 FILLER_49_806 ();
 sg13g2_decap_8 FILLER_49_813 ();
 sg13g2_decap_8 FILLER_49_820 ();
 sg13g2_decap_8 FILLER_49_827 ();
 sg13g2_decap_8 FILLER_49_834 ();
 sg13g2_decap_8 FILLER_49_841 ();
 sg13g2_decap_8 FILLER_49_848 ();
 sg13g2_decap_8 FILLER_49_855 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_4 FILLER_50_7 ();
 sg13g2_fill_1 FILLER_50_11 ();
 sg13g2_fill_1 FILLER_50_16 ();
 sg13g2_fill_1 FILLER_50_48 ();
 sg13g2_decap_4 FILLER_50_65 ();
 sg13g2_decap_4 FILLER_50_77 ();
 sg13g2_fill_1 FILLER_50_81 ();
 sg13g2_decap_4 FILLER_50_92 ();
 sg13g2_fill_1 FILLER_50_96 ();
 sg13g2_fill_2 FILLER_50_115 ();
 sg13g2_decap_4 FILLER_50_121 ();
 sg13g2_fill_2 FILLER_50_125 ();
 sg13g2_decap_8 FILLER_50_143 ();
 sg13g2_fill_1 FILLER_50_154 ();
 sg13g2_decap_8 FILLER_50_160 ();
 sg13g2_fill_2 FILLER_50_167 ();
 sg13g2_decap_4 FILLER_50_195 ();
 sg13g2_fill_1 FILLER_50_199 ();
 sg13g2_fill_2 FILLER_50_205 ();
 sg13g2_decap_8 FILLER_50_240 ();
 sg13g2_decap_4 FILLER_50_247 ();
 sg13g2_fill_1 FILLER_50_287 ();
 sg13g2_decap_4 FILLER_50_303 ();
 sg13g2_fill_1 FILLER_50_307 ();
 sg13g2_fill_2 FILLER_50_319 ();
 sg13g2_fill_1 FILLER_50_321 ();
 sg13g2_fill_2 FILLER_50_327 ();
 sg13g2_fill_1 FILLER_50_329 ();
 sg13g2_fill_1 FILLER_50_348 ();
 sg13g2_decap_4 FILLER_50_354 ();
 sg13g2_fill_2 FILLER_50_358 ();
 sg13g2_decap_8 FILLER_50_374 ();
 sg13g2_decap_8 FILLER_50_381 ();
 sg13g2_fill_2 FILLER_50_388 ();
 sg13g2_fill_1 FILLER_50_390 ();
 sg13g2_fill_2 FILLER_50_399 ();
 sg13g2_fill_1 FILLER_50_401 ();
 sg13g2_fill_1 FILLER_50_436 ();
 sg13g2_fill_1 FILLER_50_442 ();
 sg13g2_decap_4 FILLER_50_451 ();
 sg13g2_decap_4 FILLER_50_463 ();
 sg13g2_fill_2 FILLER_50_467 ();
 sg13g2_fill_1 FILLER_50_493 ();
 sg13g2_decap_8 FILLER_50_500 ();
 sg13g2_fill_2 FILLER_50_507 ();
 sg13g2_decap_8 FILLER_50_525 ();
 sg13g2_fill_2 FILLER_50_532 ();
 sg13g2_fill_1 FILLER_50_554 ();
 sg13g2_fill_2 FILLER_50_569 ();
 sg13g2_decap_4 FILLER_50_588 ();
 sg13g2_fill_2 FILLER_50_609 ();
 sg13g2_fill_1 FILLER_50_611 ();
 sg13g2_fill_2 FILLER_50_620 ();
 sg13g2_fill_2 FILLER_50_648 ();
 sg13g2_fill_1 FILLER_50_650 ();
 sg13g2_fill_2 FILLER_50_660 ();
 sg13g2_fill_1 FILLER_50_668 ();
 sg13g2_decap_8 FILLER_50_674 ();
 sg13g2_fill_2 FILLER_50_681 ();
 sg13g2_decap_8 FILLER_50_688 ();
 sg13g2_decap_4 FILLER_50_695 ();
 sg13g2_fill_2 FILLER_50_707 ();
 sg13g2_decap_8 FILLER_50_747 ();
 sg13g2_fill_1 FILLER_50_754 ();
 sg13g2_decap_8 FILLER_50_764 ();
 sg13g2_decap_8 FILLER_50_771 ();
 sg13g2_decap_8 FILLER_50_778 ();
 sg13g2_decap_8 FILLER_50_785 ();
 sg13g2_decap_8 FILLER_50_792 ();
 sg13g2_decap_8 FILLER_50_799 ();
 sg13g2_decap_8 FILLER_50_806 ();
 sg13g2_decap_8 FILLER_50_813 ();
 sg13g2_decap_8 FILLER_50_820 ();
 sg13g2_decap_8 FILLER_50_827 ();
 sg13g2_decap_8 FILLER_50_834 ();
 sg13g2_decap_8 FILLER_50_841 ();
 sg13g2_decap_8 FILLER_50_848 ();
 sg13g2_decap_8 FILLER_50_855 ();
 sg13g2_fill_2 FILLER_51_26 ();
 sg13g2_fill_1 FILLER_51_28 ();
 sg13g2_fill_2 FILLER_51_63 ();
 sg13g2_fill_1 FILLER_51_65 ();
 sg13g2_fill_1 FILLER_51_74 ();
 sg13g2_fill_2 FILLER_51_96 ();
 sg13g2_fill_1 FILLER_51_98 ();
 sg13g2_fill_2 FILLER_51_118 ();
 sg13g2_decap_4 FILLER_51_145 ();
 sg13g2_fill_1 FILLER_51_149 ();
 sg13g2_fill_2 FILLER_51_191 ();
 sg13g2_fill_1 FILLER_51_193 ();
 sg13g2_fill_1 FILLER_51_221 ();
 sg13g2_fill_2 FILLER_51_233 ();
 sg13g2_fill_2 FILLER_51_262 ();
 sg13g2_fill_1 FILLER_51_264 ();
 sg13g2_decap_8 FILLER_51_274 ();
 sg13g2_decap_4 FILLER_51_281 ();
 sg13g2_fill_1 FILLER_51_285 ();
 sg13g2_decap_8 FILLER_51_290 ();
 sg13g2_fill_2 FILLER_51_297 ();
 sg13g2_fill_1 FILLER_51_299 ();
 sg13g2_decap_4 FILLER_51_324 ();
 sg13g2_decap_4 FILLER_51_348 ();
 sg13g2_fill_1 FILLER_51_352 ();
 sg13g2_fill_1 FILLER_51_393 ();
 sg13g2_decap_8 FILLER_51_406 ();
 sg13g2_decap_8 FILLER_51_417 ();
 sg13g2_decap_8 FILLER_51_424 ();
 sg13g2_decap_4 FILLER_51_431 ();
 sg13g2_fill_2 FILLER_51_445 ();
 sg13g2_fill_1 FILLER_51_447 ();
 sg13g2_fill_1 FILLER_51_456 ();
 sg13g2_decap_8 FILLER_51_470 ();
 sg13g2_fill_2 FILLER_51_477 ();
 sg13g2_fill_2 FILLER_51_505 ();
 sg13g2_decap_8 FILLER_51_524 ();
 sg13g2_decap_8 FILLER_51_551 ();
 sg13g2_fill_2 FILLER_51_571 ();
 sg13g2_fill_2 FILLER_51_588 ();
 sg13g2_decap_8 FILLER_51_622 ();
 sg13g2_decap_4 FILLER_51_643 ();
 sg13g2_decap_8 FILLER_51_699 ();
 sg13g2_decap_4 FILLER_51_706 ();
 sg13g2_fill_2 FILLER_51_718 ();
 sg13g2_decap_4 FILLER_51_724 ();
 sg13g2_decap_8 FILLER_51_733 ();
 sg13g2_fill_2 FILLER_51_740 ();
 sg13g2_fill_1 FILLER_51_742 ();
 sg13g2_decap_8 FILLER_51_769 ();
 sg13g2_decap_8 FILLER_51_776 ();
 sg13g2_decap_8 FILLER_51_783 ();
 sg13g2_decap_8 FILLER_51_790 ();
 sg13g2_decap_8 FILLER_51_797 ();
 sg13g2_decap_8 FILLER_51_804 ();
 sg13g2_decap_8 FILLER_51_811 ();
 sg13g2_decap_8 FILLER_51_818 ();
 sg13g2_decap_8 FILLER_51_825 ();
 sg13g2_decap_8 FILLER_51_832 ();
 sg13g2_decap_8 FILLER_51_839 ();
 sg13g2_decap_8 FILLER_51_846 ();
 sg13g2_decap_8 FILLER_51_853 ();
 sg13g2_fill_2 FILLER_51_860 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_4 FILLER_52_7 ();
 sg13g2_fill_2 FILLER_52_15 ();
 sg13g2_fill_1 FILLER_52_17 ();
 sg13g2_decap_8 FILLER_52_40 ();
 sg13g2_decap_4 FILLER_52_47 ();
 sg13g2_fill_2 FILLER_52_51 ();
 sg13g2_decap_4 FILLER_52_62 ();
 sg13g2_fill_1 FILLER_52_66 ();
 sg13g2_fill_2 FILLER_52_91 ();
 sg13g2_fill_2 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_118 ();
 sg13g2_decap_4 FILLER_52_125 ();
 sg13g2_fill_1 FILLER_52_129 ();
 sg13g2_fill_2 FILLER_52_143 ();
 sg13g2_fill_1 FILLER_52_145 ();
 sg13g2_fill_1 FILLER_52_154 ();
 sg13g2_fill_2 FILLER_52_165 ();
 sg13g2_fill_1 FILLER_52_167 ();
 sg13g2_fill_1 FILLER_52_182 ();
 sg13g2_decap_4 FILLER_52_196 ();
 sg13g2_fill_2 FILLER_52_212 ();
 sg13g2_fill_2 FILLER_52_219 ();
 sg13g2_decap_8 FILLER_52_242 ();
 sg13g2_decap_4 FILLER_52_249 ();
 sg13g2_fill_2 FILLER_52_253 ();
 sg13g2_fill_2 FILLER_52_271 ();
 sg13g2_fill_2 FILLER_52_281 ();
 sg13g2_decap_4 FILLER_52_288 ();
 sg13g2_decap_8 FILLER_52_301 ();
 sg13g2_fill_1 FILLER_52_308 ();
 sg13g2_decap_8 FILLER_52_322 ();
 sg13g2_fill_2 FILLER_52_329 ();
 sg13g2_decap_8 FILLER_52_336 ();
 sg13g2_decap_8 FILLER_52_343 ();
 sg13g2_decap_4 FILLER_52_350 ();
 sg13g2_decap_8 FILLER_52_366 ();
 sg13g2_decap_4 FILLER_52_373 ();
 sg13g2_fill_1 FILLER_52_377 ();
 sg13g2_decap_4 FILLER_52_382 ();
 sg13g2_fill_2 FILLER_52_386 ();
 sg13g2_decap_8 FILLER_52_393 ();
 sg13g2_fill_2 FILLER_52_400 ();
 sg13g2_fill_1 FILLER_52_402 ();
 sg13g2_decap_8 FILLER_52_411 ();
 sg13g2_decap_4 FILLER_52_418 ();
 sg13g2_fill_2 FILLER_52_435 ();
 sg13g2_fill_1 FILLER_52_437 ();
 sg13g2_decap_8 FILLER_52_443 ();
 sg13g2_fill_1 FILLER_52_450 ();
 sg13g2_fill_1 FILLER_52_488 ();
 sg13g2_decap_8 FILLER_52_493 ();
 sg13g2_decap_4 FILLER_52_508 ();
 sg13g2_decap_4 FILLER_52_520 ();
 sg13g2_fill_1 FILLER_52_524 ();
 sg13g2_decap_4 FILLER_52_529 ();
 sg13g2_fill_1 FILLER_52_539 ();
 sg13g2_decap_8 FILLER_52_545 ();
 sg13g2_decap_4 FILLER_52_552 ();
 sg13g2_fill_2 FILLER_52_556 ();
 sg13g2_decap_4 FILLER_52_593 ();
 sg13g2_fill_2 FILLER_52_597 ();
 sg13g2_fill_2 FILLER_52_605 ();
 sg13g2_fill_1 FILLER_52_607 ();
 sg13g2_decap_4 FILLER_52_626 ();
 sg13g2_fill_1 FILLER_52_630 ();
 sg13g2_decap_8 FILLER_52_646 ();
 sg13g2_decap_4 FILLER_52_653 ();
 sg13g2_decap_8 FILLER_52_666 ();
 sg13g2_decap_4 FILLER_52_673 ();
 sg13g2_fill_1 FILLER_52_677 ();
 sg13g2_fill_2 FILLER_52_684 ();
 sg13g2_decap_8 FILLER_52_697 ();
 sg13g2_decap_4 FILLER_52_704 ();
 sg13g2_fill_1 FILLER_52_708 ();
 sg13g2_decap_4 FILLER_52_722 ();
 sg13g2_fill_2 FILLER_52_726 ();
 sg13g2_fill_2 FILLER_52_733 ();
 sg13g2_decap_8 FILLER_52_741 ();
 sg13g2_decap_4 FILLER_52_748 ();
 sg13g2_decap_8 FILLER_52_769 ();
 sg13g2_decap_8 FILLER_52_776 ();
 sg13g2_decap_8 FILLER_52_783 ();
 sg13g2_decap_8 FILLER_52_790 ();
 sg13g2_decap_8 FILLER_52_797 ();
 sg13g2_decap_8 FILLER_52_804 ();
 sg13g2_decap_8 FILLER_52_811 ();
 sg13g2_decap_8 FILLER_52_818 ();
 sg13g2_decap_8 FILLER_52_825 ();
 sg13g2_decap_8 FILLER_52_832 ();
 sg13g2_decap_8 FILLER_52_839 ();
 sg13g2_decap_8 FILLER_52_846 ();
 sg13g2_decap_8 FILLER_52_853 ();
 sg13g2_fill_2 FILLER_52_860 ();
 sg13g2_fill_1 FILLER_53_36 ();
 sg13g2_fill_2 FILLER_53_46 ();
 sg13g2_fill_1 FILLER_53_65 ();
 sg13g2_decap_4 FILLER_53_77 ();
 sg13g2_fill_1 FILLER_53_81 ();
 sg13g2_decap_8 FILLER_53_85 ();
 sg13g2_fill_2 FILLER_53_92 ();
 sg13g2_decap_4 FILLER_53_128 ();
 sg13g2_fill_2 FILLER_53_143 ();
 sg13g2_fill_1 FILLER_53_145 ();
 sg13g2_fill_1 FILLER_53_160 ();
 sg13g2_fill_2 FILLER_53_166 ();
 sg13g2_decap_4 FILLER_53_177 ();
 sg13g2_fill_2 FILLER_53_213 ();
 sg13g2_fill_1 FILLER_53_215 ();
 sg13g2_fill_2 FILLER_53_221 ();
 sg13g2_fill_1 FILLER_53_223 ();
 sg13g2_decap_4 FILLER_53_238 ();
 sg13g2_fill_1 FILLER_53_242 ();
 sg13g2_decap_4 FILLER_53_255 ();
 sg13g2_fill_2 FILLER_53_259 ();
 sg13g2_fill_1 FILLER_53_271 ();
 sg13g2_fill_1 FILLER_53_282 ();
 sg13g2_fill_2 FILLER_53_303 ();
 sg13g2_fill_1 FILLER_53_341 ();
 sg13g2_fill_2 FILLER_53_357 ();
 sg13g2_fill_1 FILLER_53_359 ();
 sg13g2_fill_1 FILLER_53_370 ();
 sg13g2_fill_2 FILLER_53_397 ();
 sg13g2_fill_1 FILLER_53_399 ();
 sg13g2_decap_4 FILLER_53_404 ();
 sg13g2_fill_2 FILLER_53_408 ();
 sg13g2_decap_4 FILLER_53_489 ();
 sg13g2_fill_1 FILLER_53_493 ();
 sg13g2_fill_1 FILLER_53_504 ();
 sg13g2_decap_8 FILLER_53_521 ();
 sg13g2_fill_2 FILLER_53_528 ();
 sg13g2_fill_2 FILLER_53_552 ();
 sg13g2_decap_8 FILLER_53_567 ();
 sg13g2_decap_4 FILLER_53_574 ();
 sg13g2_decap_8 FILLER_53_583 ();
 sg13g2_fill_2 FILLER_53_590 ();
 sg13g2_fill_1 FILLER_53_592 ();
 sg13g2_decap_8 FILLER_53_623 ();
 sg13g2_fill_1 FILLER_53_630 ();
 sg13g2_decap_4 FILLER_53_644 ();
 sg13g2_fill_1 FILLER_53_674 ();
 sg13g2_fill_2 FILLER_53_744 ();
 sg13g2_decap_8 FILLER_53_762 ();
 sg13g2_decap_8 FILLER_53_769 ();
 sg13g2_decap_8 FILLER_53_776 ();
 sg13g2_decap_8 FILLER_53_783 ();
 sg13g2_decap_8 FILLER_53_790 ();
 sg13g2_decap_8 FILLER_53_797 ();
 sg13g2_decap_8 FILLER_53_804 ();
 sg13g2_decap_8 FILLER_53_811 ();
 sg13g2_decap_8 FILLER_53_818 ();
 sg13g2_decap_8 FILLER_53_825 ();
 sg13g2_decap_8 FILLER_53_832 ();
 sg13g2_decap_8 FILLER_53_839 ();
 sg13g2_decap_8 FILLER_53_846 ();
 sg13g2_decap_8 FILLER_53_853 ();
 sg13g2_fill_2 FILLER_53_860 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_4 FILLER_54_7 ();
 sg13g2_fill_2 FILLER_54_19 ();
 sg13g2_decap_4 FILLER_54_44 ();
 sg13g2_decap_4 FILLER_54_53 ();
 sg13g2_fill_2 FILLER_54_78 ();
 sg13g2_decap_8 FILLER_54_95 ();
 sg13g2_decap_4 FILLER_54_102 ();
 sg13g2_fill_2 FILLER_54_106 ();
 sg13g2_fill_2 FILLER_54_111 ();
 sg13g2_fill_1 FILLER_54_113 ();
 sg13g2_fill_1 FILLER_54_118 ();
 sg13g2_decap_8 FILLER_54_150 ();
 sg13g2_fill_2 FILLER_54_165 ();
 sg13g2_fill_1 FILLER_54_167 ();
 sg13g2_fill_1 FILLER_54_194 ();
 sg13g2_fill_1 FILLER_54_207 ();
 sg13g2_decap_8 FILLER_54_227 ();
 sg13g2_fill_2 FILLER_54_234 ();
 sg13g2_fill_1 FILLER_54_236 ();
 sg13g2_fill_2 FILLER_54_250 ();
 sg13g2_fill_1 FILLER_54_261 ();
 sg13g2_fill_2 FILLER_54_276 ();
 sg13g2_fill_1 FILLER_54_278 ();
 sg13g2_fill_2 FILLER_54_284 ();
 sg13g2_fill_1 FILLER_54_286 ();
 sg13g2_fill_1 FILLER_54_296 ();
 sg13g2_fill_2 FILLER_54_301 ();
 sg13g2_fill_1 FILLER_54_325 ();
 sg13g2_fill_1 FILLER_54_334 ();
 sg13g2_decap_8 FILLER_54_343 ();
 sg13g2_fill_1 FILLER_54_350 ();
 sg13g2_fill_2 FILLER_54_360 ();
 sg13g2_fill_1 FILLER_54_362 ();
 sg13g2_fill_1 FILLER_54_375 ();
 sg13g2_decap_4 FILLER_54_423 ();
 sg13g2_decap_4 FILLER_54_466 ();
 sg13g2_fill_1 FILLER_54_470 ();
 sg13g2_decap_8 FILLER_54_482 ();
 sg13g2_decap_8 FILLER_54_489 ();
 sg13g2_fill_2 FILLER_54_504 ();
 sg13g2_fill_1 FILLER_54_506 ();
 sg13g2_fill_2 FILLER_54_515 ();
 sg13g2_fill_1 FILLER_54_517 ();
 sg13g2_fill_1 FILLER_54_526 ();
 sg13g2_fill_2 FILLER_54_535 ();
 sg13g2_fill_1 FILLER_54_542 ();
 sg13g2_decap_8 FILLER_54_546 ();
 sg13g2_decap_4 FILLER_54_553 ();
 sg13g2_decap_8 FILLER_54_591 ();
 sg13g2_fill_2 FILLER_54_598 ();
 sg13g2_decap_8 FILLER_54_619 ();
 sg13g2_fill_1 FILLER_54_626 ();
 sg13g2_decap_4 FILLER_54_642 ();
 sg13g2_fill_1 FILLER_54_646 ();
 sg13g2_fill_2 FILLER_54_655 ();
 sg13g2_fill_1 FILLER_54_657 ();
 sg13g2_decap_8 FILLER_54_668 ();
 sg13g2_decap_4 FILLER_54_675 ();
 sg13g2_decap_4 FILLER_54_685 ();
 sg13g2_fill_2 FILLER_54_702 ();
 sg13g2_fill_2 FILLER_54_712 ();
 sg13g2_fill_1 FILLER_54_727 ();
 sg13g2_fill_1 FILLER_54_733 ();
 sg13g2_decap_4 FILLER_54_738 ();
 sg13g2_decap_8 FILLER_54_765 ();
 sg13g2_decap_8 FILLER_54_772 ();
 sg13g2_decap_8 FILLER_54_779 ();
 sg13g2_decap_8 FILLER_54_786 ();
 sg13g2_decap_8 FILLER_54_793 ();
 sg13g2_decap_8 FILLER_54_800 ();
 sg13g2_decap_8 FILLER_54_807 ();
 sg13g2_decap_8 FILLER_54_814 ();
 sg13g2_decap_8 FILLER_54_821 ();
 sg13g2_decap_8 FILLER_54_828 ();
 sg13g2_decap_8 FILLER_54_835 ();
 sg13g2_decap_8 FILLER_54_842 ();
 sg13g2_decap_8 FILLER_54_849 ();
 sg13g2_decap_4 FILLER_54_856 ();
 sg13g2_fill_2 FILLER_54_860 ();
 sg13g2_fill_2 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_2 ();
 sg13g2_fill_2 FILLER_55_29 ();
 sg13g2_fill_1 FILLER_55_31 ();
 sg13g2_decap_4 FILLER_55_58 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_4 FILLER_55_84 ();
 sg13g2_fill_1 FILLER_55_130 ();
 sg13g2_fill_2 FILLER_55_168 ();
 sg13g2_fill_1 FILLER_55_184 ();
 sg13g2_fill_1 FILLER_55_214 ();
 sg13g2_fill_2 FILLER_55_220 ();
 sg13g2_fill_1 FILLER_55_244 ();
 sg13g2_decap_8 FILLER_55_250 ();
 sg13g2_fill_1 FILLER_55_282 ();
 sg13g2_fill_2 FILLER_55_298 ();
 sg13g2_fill_1 FILLER_55_300 ();
 sg13g2_fill_2 FILLER_55_334 ();
 sg13g2_fill_1 FILLER_55_351 ();
 sg13g2_decap_8 FILLER_55_360 ();
 sg13g2_fill_2 FILLER_55_367 ();
 sg13g2_fill_1 FILLER_55_374 ();
 sg13g2_fill_2 FILLER_55_380 ();
 sg13g2_fill_1 FILLER_55_396 ();
 sg13g2_fill_2 FILLER_55_444 ();
 sg13g2_fill_1 FILLER_55_458 ();
 sg13g2_decap_4 FILLER_55_515 ();
 sg13g2_fill_2 FILLER_55_547 ();
 sg13g2_fill_1 FILLER_55_549 ();
 sg13g2_fill_2 FILLER_55_560 ();
 sg13g2_fill_1 FILLER_55_562 ();
 sg13g2_decap_4 FILLER_55_572 ();
 sg13g2_fill_1 FILLER_55_576 ();
 sg13g2_decap_4 FILLER_55_596 ();
 sg13g2_fill_1 FILLER_55_608 ();
 sg13g2_fill_2 FILLER_55_625 ();
 sg13g2_fill_2 FILLER_55_632 ();
 sg13g2_fill_1 FILLER_55_652 ();
 sg13g2_fill_2 FILLER_55_661 ();
 sg13g2_decap_8 FILLER_55_695 ();
 sg13g2_fill_2 FILLER_55_702 ();
 sg13g2_fill_2 FILLER_55_722 ();
 sg13g2_fill_1 FILLER_55_724 ();
 sg13g2_decap_4 FILLER_55_733 ();
 sg13g2_fill_2 FILLER_55_737 ();
 sg13g2_decap_8 FILLER_55_761 ();
 sg13g2_decap_8 FILLER_55_768 ();
 sg13g2_decap_8 FILLER_55_775 ();
 sg13g2_decap_8 FILLER_55_782 ();
 sg13g2_decap_8 FILLER_55_789 ();
 sg13g2_decap_8 FILLER_55_796 ();
 sg13g2_decap_8 FILLER_55_803 ();
 sg13g2_decap_8 FILLER_55_810 ();
 sg13g2_decap_8 FILLER_55_817 ();
 sg13g2_decap_8 FILLER_55_824 ();
 sg13g2_decap_8 FILLER_55_831 ();
 sg13g2_decap_8 FILLER_55_838 ();
 sg13g2_decap_8 FILLER_55_845 ();
 sg13g2_decap_8 FILLER_55_852 ();
 sg13g2_fill_2 FILLER_55_859 ();
 sg13g2_fill_1 FILLER_55_861 ();
 sg13g2_decap_4 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_4 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_fill_1 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_55 ();
 sg13g2_fill_2 FILLER_56_62 ();
 sg13g2_fill_1 FILLER_56_102 ();
 sg13g2_fill_1 FILLER_56_140 ();
 sg13g2_fill_2 FILLER_56_168 ();
 sg13g2_decap_4 FILLER_56_182 ();
 sg13g2_fill_2 FILLER_56_186 ();
 sg13g2_fill_1 FILLER_56_202 ();
 sg13g2_fill_1 FILLER_56_213 ();
 sg13g2_fill_2 FILLER_56_224 ();
 sg13g2_fill_2 FILLER_56_239 ();
 sg13g2_fill_2 FILLER_56_246 ();
 sg13g2_fill_1 FILLER_56_248 ();
 sg13g2_fill_2 FILLER_56_262 ();
 sg13g2_fill_1 FILLER_56_264 ();
 sg13g2_fill_1 FILLER_56_270 ();
 sg13g2_decap_8 FILLER_56_285 ();
 sg13g2_decap_8 FILLER_56_292 ();
 sg13g2_decap_4 FILLER_56_299 ();
 sg13g2_fill_1 FILLER_56_315 ();
 sg13g2_fill_2 FILLER_56_325 ();
 sg13g2_decap_8 FILLER_56_335 ();
 sg13g2_fill_1 FILLER_56_342 ();
 sg13g2_fill_1 FILLER_56_369 ();
 sg13g2_fill_1 FILLER_56_386 ();
 sg13g2_fill_2 FILLER_56_396 ();
 sg13g2_fill_2 FILLER_56_421 ();
 sg13g2_fill_1 FILLER_56_423 ();
 sg13g2_fill_1 FILLER_56_441 ();
 sg13g2_decap_4 FILLER_56_457 ();
 sg13g2_decap_8 FILLER_56_466 ();
 sg13g2_fill_2 FILLER_56_473 ();
 sg13g2_decap_8 FILLER_56_485 ();
 sg13g2_fill_1 FILLER_56_492 ();
 sg13g2_fill_2 FILLER_56_519 ();
 sg13g2_fill_1 FILLER_56_521 ();
 sg13g2_decap_8 FILLER_56_551 ();
 sg13g2_fill_2 FILLER_56_558 ();
 sg13g2_decap_4 FILLER_56_571 ();
 sg13g2_fill_1 FILLER_56_575 ();
 sg13g2_fill_2 FILLER_56_581 ();
 sg13g2_decap_4 FILLER_56_610 ();
 sg13g2_fill_1 FILLER_56_628 ();
 sg13g2_decap_4 FILLER_56_647 ();
 sg13g2_fill_2 FILLER_56_651 ();
 sg13g2_fill_2 FILLER_56_656 ();
 sg13g2_fill_1 FILLER_56_678 ();
 sg13g2_fill_1 FILLER_56_701 ();
 sg13g2_fill_2 FILLER_56_714 ();
 sg13g2_decap_4 FILLER_56_725 ();
 sg13g2_decap_8 FILLER_56_759 ();
 sg13g2_decap_8 FILLER_56_766 ();
 sg13g2_decap_8 FILLER_56_773 ();
 sg13g2_decap_8 FILLER_56_780 ();
 sg13g2_decap_8 FILLER_56_787 ();
 sg13g2_decap_8 FILLER_56_794 ();
 sg13g2_decap_8 FILLER_56_801 ();
 sg13g2_decap_8 FILLER_56_808 ();
 sg13g2_decap_8 FILLER_56_815 ();
 sg13g2_decap_8 FILLER_56_822 ();
 sg13g2_decap_8 FILLER_56_829 ();
 sg13g2_decap_8 FILLER_56_836 ();
 sg13g2_decap_8 FILLER_56_843 ();
 sg13g2_decap_8 FILLER_56_850 ();
 sg13g2_decap_4 FILLER_56_857 ();
 sg13g2_fill_1 FILLER_56_861 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_32 ();
 sg13g2_fill_2 FILLER_57_39 ();
 sg13g2_fill_1 FILLER_57_41 ();
 sg13g2_fill_2 FILLER_57_76 ();
 sg13g2_decap_8 FILLER_57_82 ();
 sg13g2_fill_2 FILLER_57_89 ();
 sg13g2_fill_1 FILLER_57_91 ();
 sg13g2_decap_4 FILLER_57_107 ();
 sg13g2_decap_4 FILLER_57_140 ();
 sg13g2_fill_1 FILLER_57_144 ();
 sg13g2_fill_2 FILLER_57_166 ();
 sg13g2_fill_1 FILLER_57_182 ();
 sg13g2_fill_2 FILLER_57_208 ();
 sg13g2_fill_1 FILLER_57_210 ();
 sg13g2_decap_4 FILLER_57_236 ();
 sg13g2_decap_8 FILLER_57_283 ();
 sg13g2_fill_2 FILLER_57_290 ();
 sg13g2_fill_1 FILLER_57_292 ();
 sg13g2_fill_2 FILLER_57_298 ();
 sg13g2_fill_1 FILLER_57_311 ();
 sg13g2_fill_2 FILLER_57_326 ();
 sg13g2_fill_1 FILLER_57_328 ();
 sg13g2_decap_8 FILLER_57_337 ();
 sg13g2_decap_8 FILLER_57_344 ();
 sg13g2_fill_2 FILLER_57_351 ();
 sg13g2_decap_8 FILLER_57_362 ();
 sg13g2_decap_8 FILLER_57_369 ();
 sg13g2_fill_2 FILLER_57_384 ();
 sg13g2_fill_2 FILLER_57_394 ();
 sg13g2_fill_1 FILLER_57_432 ();
 sg13g2_decap_4 FILLER_57_450 ();
 sg13g2_fill_2 FILLER_57_454 ();
 sg13g2_decap_8 FILLER_57_490 ();
 sg13g2_fill_2 FILLER_57_497 ();
 sg13g2_fill_1 FILLER_57_499 ();
 sg13g2_fill_2 FILLER_57_508 ();
 sg13g2_fill_1 FILLER_57_510 ();
 sg13g2_decap_4 FILLER_57_519 ();
 sg13g2_fill_2 FILLER_57_541 ();
 sg13g2_fill_1 FILLER_57_567 ();
 sg13g2_decap_8 FILLER_57_605 ();
 sg13g2_fill_2 FILLER_57_612 ();
 sg13g2_decap_8 FILLER_57_626 ();
 sg13g2_fill_2 FILLER_57_633 ();
 sg13g2_fill_1 FILLER_57_635 ();
 sg13g2_decap_8 FILLER_57_644 ();
 sg13g2_decap_4 FILLER_57_651 ();
 sg13g2_fill_1 FILLER_57_655 ();
 sg13g2_fill_2 FILLER_57_667 ();
 sg13g2_fill_1 FILLER_57_669 ();
 sg13g2_decap_8 FILLER_57_676 ();
 sg13g2_decap_8 FILLER_57_683 ();
 sg13g2_decap_8 FILLER_57_690 ();
 sg13g2_fill_2 FILLER_57_697 ();
 sg13g2_fill_1 FILLER_57_699 ();
 sg13g2_decap_8 FILLER_57_731 ();
 sg13g2_fill_1 FILLER_57_738 ();
 sg13g2_fill_1 FILLER_57_743 ();
 sg13g2_decap_8 FILLER_57_755 ();
 sg13g2_decap_8 FILLER_57_762 ();
 sg13g2_decap_8 FILLER_57_769 ();
 sg13g2_decap_8 FILLER_57_776 ();
 sg13g2_decap_8 FILLER_57_783 ();
 sg13g2_decap_8 FILLER_57_790 ();
 sg13g2_decap_8 FILLER_57_797 ();
 sg13g2_decap_8 FILLER_57_804 ();
 sg13g2_decap_8 FILLER_57_811 ();
 sg13g2_decap_8 FILLER_57_818 ();
 sg13g2_decap_8 FILLER_57_825 ();
 sg13g2_decap_8 FILLER_57_832 ();
 sg13g2_decap_8 FILLER_57_839 ();
 sg13g2_decap_8 FILLER_57_846 ();
 sg13g2_decap_8 FILLER_57_853 ();
 sg13g2_fill_2 FILLER_57_860 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_7 ();
 sg13g2_decap_4 FILLER_58_12 ();
 sg13g2_fill_1 FILLER_58_16 ();
 sg13g2_decap_8 FILLER_58_25 ();
 sg13g2_decap_8 FILLER_58_32 ();
 sg13g2_decap_8 FILLER_58_48 ();
 sg13g2_fill_1 FILLER_58_55 ();
 sg13g2_decap_4 FILLER_58_65 ();
 sg13g2_fill_1 FILLER_58_69 ();
 sg13g2_decap_4 FILLER_58_81 ();
 sg13g2_fill_1 FILLER_58_117 ();
 sg13g2_fill_2 FILLER_58_126 ();
 sg13g2_fill_2 FILLER_58_143 ();
 sg13g2_fill_1 FILLER_58_156 ();
 sg13g2_fill_2 FILLER_58_175 ();
 sg13g2_fill_2 FILLER_58_185 ();
 sg13g2_fill_2 FILLER_58_203 ();
 sg13g2_decap_4 FILLER_58_212 ();
 sg13g2_decap_8 FILLER_58_227 ();
 sg13g2_fill_2 FILLER_58_234 ();
 sg13g2_decap_8 FILLER_58_242 ();
 sg13g2_decap_4 FILLER_58_249 ();
 sg13g2_fill_2 FILLER_58_258 ();
 sg13g2_decap_8 FILLER_58_291 ();
 sg13g2_fill_1 FILLER_58_298 ();
 sg13g2_fill_1 FILLER_58_304 ();
 sg13g2_decap_8 FILLER_58_315 ();
 sg13g2_decap_4 FILLER_58_326 ();
 sg13g2_fill_2 FILLER_58_330 ();
 sg13g2_decap_4 FILLER_58_341 ();
 sg13g2_fill_1 FILLER_58_345 ();
 sg13g2_fill_2 FILLER_58_358 ();
 sg13g2_decap_4 FILLER_58_379 ();
 sg13g2_decap_8 FILLER_58_421 ();
 sg13g2_fill_2 FILLER_58_445 ();
 sg13g2_fill_1 FILLER_58_447 ();
 sg13g2_decap_4 FILLER_58_470 ();
 sg13g2_decap_4 FILLER_58_482 ();
 sg13g2_fill_2 FILLER_58_486 ();
 sg13g2_fill_2 FILLER_58_493 ();
 sg13g2_fill_1 FILLER_58_495 ();
 sg13g2_fill_1 FILLER_58_520 ();
 sg13g2_decap_8 FILLER_58_525 ();
 sg13g2_fill_1 FILLER_58_532 ();
 sg13g2_decap_8 FILLER_58_558 ();
 sg13g2_decap_8 FILLER_58_571 ();
 sg13g2_fill_2 FILLER_58_578 ();
 sg13g2_fill_2 FILLER_58_584 ();
 sg13g2_fill_2 FILLER_58_604 ();
 sg13g2_decap_8 FILLER_58_612 ();
 sg13g2_decap_4 FILLER_58_619 ();
 sg13g2_fill_2 FILLER_58_633 ();
 sg13g2_fill_1 FILLER_58_635 ();
 sg13g2_decap_4 FILLER_58_647 ();
 sg13g2_fill_2 FILLER_58_651 ();
 sg13g2_fill_1 FILLER_58_673 ();
 sg13g2_fill_2 FILLER_58_706 ();
 sg13g2_fill_1 FILLER_58_708 ();
 sg13g2_decap_4 FILLER_58_726 ();
 sg13g2_fill_2 FILLER_58_730 ();
 sg13g2_decap_8 FILLER_58_759 ();
 sg13g2_decap_8 FILLER_58_766 ();
 sg13g2_decap_8 FILLER_58_773 ();
 sg13g2_decap_8 FILLER_58_780 ();
 sg13g2_decap_8 FILLER_58_787 ();
 sg13g2_decap_8 FILLER_58_794 ();
 sg13g2_decap_8 FILLER_58_801 ();
 sg13g2_decap_8 FILLER_58_808 ();
 sg13g2_decap_8 FILLER_58_815 ();
 sg13g2_decap_8 FILLER_58_822 ();
 sg13g2_decap_8 FILLER_58_829 ();
 sg13g2_decap_8 FILLER_58_836 ();
 sg13g2_decap_8 FILLER_58_843 ();
 sg13g2_decap_8 FILLER_58_850 ();
 sg13g2_decap_4 FILLER_58_857 ();
 sg13g2_fill_1 FILLER_58_861 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_7 ();
 sg13g2_fill_1 FILLER_59_12 ();
 sg13g2_fill_1 FILLER_59_43 ();
 sg13g2_fill_1 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_145 ();
 sg13g2_fill_2 FILLER_59_152 ();
 sg13g2_fill_1 FILLER_59_154 ();
 sg13g2_fill_1 FILLER_59_160 ();
 sg13g2_decap_8 FILLER_59_176 ();
 sg13g2_decap_4 FILLER_59_183 ();
 sg13g2_fill_2 FILLER_59_187 ();
 sg13g2_decap_8 FILLER_59_200 ();
 sg13g2_decap_8 FILLER_59_207 ();
 sg13g2_decap_8 FILLER_59_214 ();
 sg13g2_fill_1 FILLER_59_230 ();
 sg13g2_fill_2 FILLER_59_248 ();
 sg13g2_decap_4 FILLER_59_262 ();
 sg13g2_fill_1 FILLER_59_266 ();
 sg13g2_fill_1 FILLER_59_278 ();
 sg13g2_fill_1 FILLER_59_293 ();
 sg13g2_decap_4 FILLER_59_317 ();
 sg13g2_fill_2 FILLER_59_341 ();
 sg13g2_fill_1 FILLER_59_343 ();
 sg13g2_decap_4 FILLER_59_369 ();
 sg13g2_fill_2 FILLER_59_373 ();
 sg13g2_decap_4 FILLER_59_380 ();
 sg13g2_fill_1 FILLER_59_384 ();
 sg13g2_fill_2 FILLER_59_391 ();
 sg13g2_fill_1 FILLER_59_393 ();
 sg13g2_fill_2 FILLER_59_398 ();
 sg13g2_decap_4 FILLER_59_413 ();
 sg13g2_fill_1 FILLER_59_431 ();
 sg13g2_decap_8 FILLER_59_446 ();
 sg13g2_decap_4 FILLER_59_453 ();
 sg13g2_fill_2 FILLER_59_496 ();
 sg13g2_fill_1 FILLER_59_498 ();
 sg13g2_fill_2 FILLER_59_510 ();
 sg13g2_decap_8 FILLER_59_535 ();
 sg13g2_fill_1 FILLER_59_542 ();
 sg13g2_fill_2 FILLER_59_553 ();
 sg13g2_fill_1 FILLER_59_560 ();
 sg13g2_fill_2 FILLER_59_573 ();
 sg13g2_decap_4 FILLER_59_600 ();
 sg13g2_decap_4 FILLER_59_633 ();
 sg13g2_fill_2 FILLER_59_641 ();
 sg13g2_fill_1 FILLER_59_643 ();
 sg13g2_decap_8 FILLER_59_655 ();
 sg13g2_fill_1 FILLER_59_662 ();
 sg13g2_decap_8 FILLER_59_678 ();
 sg13g2_fill_2 FILLER_59_685 ();
 sg13g2_decap_8 FILLER_59_731 ();
 sg13g2_decap_4 FILLER_59_738 ();
 sg13g2_fill_2 FILLER_59_742 ();
 sg13g2_decap_8 FILLER_59_754 ();
 sg13g2_decap_8 FILLER_59_761 ();
 sg13g2_decap_8 FILLER_59_768 ();
 sg13g2_decap_8 FILLER_59_775 ();
 sg13g2_decap_8 FILLER_59_782 ();
 sg13g2_decap_8 FILLER_59_789 ();
 sg13g2_decap_8 FILLER_59_796 ();
 sg13g2_decap_8 FILLER_59_803 ();
 sg13g2_decap_8 FILLER_59_810 ();
 sg13g2_decap_8 FILLER_59_817 ();
 sg13g2_decap_8 FILLER_59_824 ();
 sg13g2_decap_8 FILLER_59_831 ();
 sg13g2_decap_8 FILLER_59_838 ();
 sg13g2_decap_8 FILLER_59_845 ();
 sg13g2_decap_8 FILLER_59_852 ();
 sg13g2_fill_2 FILLER_59_859 ();
 sg13g2_fill_1 FILLER_59_861 ();
 sg13g2_fill_2 FILLER_60_26 ();
 sg13g2_fill_2 FILLER_60_32 ();
 sg13g2_fill_1 FILLER_60_34 ();
 sg13g2_fill_2 FILLER_60_39 ();
 sg13g2_decap_4 FILLER_60_51 ();
 sg13g2_decap_4 FILLER_60_59 ();
 sg13g2_fill_2 FILLER_60_63 ();
 sg13g2_fill_1 FILLER_60_81 ();
 sg13g2_fill_2 FILLER_60_86 ();
 sg13g2_fill_1 FILLER_60_88 ();
 sg13g2_fill_1 FILLER_60_121 ();
 sg13g2_decap_4 FILLER_60_126 ();
 sg13g2_fill_1 FILLER_60_130 ();
 sg13g2_decap_8 FILLER_60_143 ();
 sg13g2_fill_2 FILLER_60_150 ();
 sg13g2_fill_1 FILLER_60_152 ();
 sg13g2_decap_4 FILLER_60_189 ();
 sg13g2_fill_1 FILLER_60_193 ();
 sg13g2_decap_4 FILLER_60_200 ();
 sg13g2_fill_1 FILLER_60_204 ();
 sg13g2_fill_1 FILLER_60_231 ();
 sg13g2_fill_2 FILLER_60_246 ();
 sg13g2_fill_1 FILLER_60_256 ();
 sg13g2_fill_2 FILLER_60_266 ();
 sg13g2_decap_8 FILLER_60_272 ();
 sg13g2_decap_4 FILLER_60_279 ();
 sg13g2_fill_2 FILLER_60_283 ();
 sg13g2_decap_4 FILLER_60_295 ();
 sg13g2_fill_1 FILLER_60_299 ();
 sg13g2_fill_1 FILLER_60_306 ();
 sg13g2_decap_8 FILLER_60_311 ();
 sg13g2_fill_2 FILLER_60_318 ();
 sg13g2_fill_2 FILLER_60_330 ();
 sg13g2_fill_1 FILLER_60_332 ();
 sg13g2_fill_1 FILLER_60_342 ();
 sg13g2_decap_8 FILLER_60_366 ();
 sg13g2_fill_2 FILLER_60_373 ();
 sg13g2_fill_1 FILLER_60_375 ();
 sg13g2_fill_2 FILLER_60_381 ();
 sg13g2_fill_1 FILLER_60_383 ();
 sg13g2_fill_1 FILLER_60_449 ();
 sg13g2_decap_4 FILLER_60_464 ();
 sg13g2_decap_4 FILLER_60_472 ();
 sg13g2_fill_2 FILLER_60_476 ();
 sg13g2_fill_2 FILLER_60_486 ();
 sg13g2_fill_1 FILLER_60_488 ();
 sg13g2_fill_2 FILLER_60_530 ();
 sg13g2_decap_8 FILLER_60_568 ();
 sg13g2_decap_8 FILLER_60_575 ();
 sg13g2_decap_8 FILLER_60_582 ();
 sg13g2_decap_8 FILLER_60_589 ();
 sg13g2_decap_8 FILLER_60_600 ();
 sg13g2_fill_1 FILLER_60_607 ();
 sg13g2_fill_2 FILLER_60_613 ();
 sg13g2_fill_2 FILLER_60_631 ();
 sg13g2_fill_2 FILLER_60_649 ();
 sg13g2_fill_1 FILLER_60_651 ();
 sg13g2_fill_2 FILLER_60_660 ();
 sg13g2_decap_8 FILLER_60_684 ();
 sg13g2_decap_4 FILLER_60_691 ();
 sg13g2_fill_2 FILLER_60_695 ();
 sg13g2_fill_2 FILLER_60_705 ();
 sg13g2_fill_2 FILLER_60_712 ();
 sg13g2_fill_1 FILLER_60_714 ();
 sg13g2_fill_2 FILLER_60_719 ();
 sg13g2_fill_1 FILLER_60_721 ();
 sg13g2_decap_8 FILLER_60_732 ();
 sg13g2_decap_8 FILLER_60_752 ();
 sg13g2_decap_8 FILLER_60_759 ();
 sg13g2_decap_8 FILLER_60_766 ();
 sg13g2_decap_8 FILLER_60_773 ();
 sg13g2_decap_8 FILLER_60_780 ();
 sg13g2_decap_8 FILLER_60_787 ();
 sg13g2_decap_8 FILLER_60_794 ();
 sg13g2_decap_8 FILLER_60_801 ();
 sg13g2_decap_8 FILLER_60_808 ();
 sg13g2_decap_8 FILLER_60_815 ();
 sg13g2_decap_8 FILLER_60_822 ();
 sg13g2_decap_8 FILLER_60_829 ();
 sg13g2_decap_8 FILLER_60_836 ();
 sg13g2_decap_8 FILLER_60_843 ();
 sg13g2_decap_8 FILLER_60_850 ();
 sg13g2_decap_4 FILLER_60_857 ();
 sg13g2_fill_1 FILLER_60_861 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_fill_1 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_55 ();
 sg13g2_fill_1 FILLER_61_62 ();
 sg13g2_decap_4 FILLER_61_66 ();
 sg13g2_decap_4 FILLER_61_74 ();
 sg13g2_decap_8 FILLER_61_86 ();
 sg13g2_fill_2 FILLER_61_93 ();
 sg13g2_fill_1 FILLER_61_95 ();
 sg13g2_fill_2 FILLER_61_115 ();
 sg13g2_fill_2 FILLER_61_154 ();
 sg13g2_fill_1 FILLER_61_156 ();
 sg13g2_fill_1 FILLER_61_169 ();
 sg13g2_fill_2 FILLER_61_178 ();
 sg13g2_fill_2 FILLER_61_192 ();
 sg13g2_fill_1 FILLER_61_200 ();
 sg13g2_fill_1 FILLER_61_213 ();
 sg13g2_decap_8 FILLER_61_232 ();
 sg13g2_decap_4 FILLER_61_239 ();
 sg13g2_fill_1 FILLER_61_243 ();
 sg13g2_decap_4 FILLER_61_249 ();
 sg13g2_fill_1 FILLER_61_253 ();
 sg13g2_fill_2 FILLER_61_264 ();
 sg13g2_fill_1 FILLER_61_266 ();
 sg13g2_fill_1 FILLER_61_271 ();
 sg13g2_fill_1 FILLER_61_292 ();
 sg13g2_fill_2 FILLER_61_301 ();
 sg13g2_fill_1 FILLER_61_303 ();
 sg13g2_fill_1 FILLER_61_310 ();
 sg13g2_fill_2 FILLER_61_322 ();
 sg13g2_fill_1 FILLER_61_324 ();
 sg13g2_fill_2 FILLER_61_336 ();
 sg13g2_fill_1 FILLER_61_338 ();
 sg13g2_fill_1 FILLER_61_360 ();
 sg13g2_decap_8 FILLER_61_387 ();
 sg13g2_decap_4 FILLER_61_394 ();
 sg13g2_fill_2 FILLER_61_398 ();
 sg13g2_decap_8 FILLER_61_404 ();
 sg13g2_decap_4 FILLER_61_411 ();
 sg13g2_fill_1 FILLER_61_415 ();
 sg13g2_decap_8 FILLER_61_445 ();
 sg13g2_decap_8 FILLER_61_458 ();
 sg13g2_decap_8 FILLER_61_465 ();
 sg13g2_decap_8 FILLER_61_483 ();
 sg13g2_fill_2 FILLER_61_490 ();
 sg13g2_decap_8 FILLER_61_508 ();
 sg13g2_decap_8 FILLER_61_531 ();
 sg13g2_decap_8 FILLER_61_538 ();
 sg13g2_decap_8 FILLER_61_574 ();
 sg13g2_fill_1 FILLER_61_607 ();
 sg13g2_decap_8 FILLER_61_634 ();
 sg13g2_fill_1 FILLER_61_641 ();
 sg13g2_fill_1 FILLER_61_662 ();
 sg13g2_decap_4 FILLER_61_675 ();
 sg13g2_fill_2 FILLER_61_679 ();
 sg13g2_fill_2 FILLER_61_697 ();
 sg13g2_decap_4 FILLER_61_710 ();
 sg13g2_fill_2 FILLER_61_714 ();
 sg13g2_decap_4 FILLER_61_729 ();
 sg13g2_fill_2 FILLER_61_733 ();
 sg13g2_decap_8 FILLER_61_762 ();
 sg13g2_decap_8 FILLER_61_769 ();
 sg13g2_decap_8 FILLER_61_776 ();
 sg13g2_decap_8 FILLER_61_783 ();
 sg13g2_decap_8 FILLER_61_790 ();
 sg13g2_decap_8 FILLER_61_797 ();
 sg13g2_decap_8 FILLER_61_804 ();
 sg13g2_decap_8 FILLER_61_811 ();
 sg13g2_decap_8 FILLER_61_818 ();
 sg13g2_decap_8 FILLER_61_825 ();
 sg13g2_decap_8 FILLER_61_832 ();
 sg13g2_decap_8 FILLER_61_839 ();
 sg13g2_decap_8 FILLER_61_846 ();
 sg13g2_decap_8 FILLER_61_853 ();
 sg13g2_fill_2 FILLER_61_860 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_2 ();
 sg13g2_fill_2 FILLER_62_37 ();
 sg13g2_fill_1 FILLER_62_39 ();
 sg13g2_decap_8 FILLER_62_44 ();
 sg13g2_decap_8 FILLER_62_51 ();
 sg13g2_fill_1 FILLER_62_58 ();
 sg13g2_decap_8 FILLER_62_139 ();
 sg13g2_fill_1 FILLER_62_146 ();
 sg13g2_decap_8 FILLER_62_159 ();
 sg13g2_decap_8 FILLER_62_166 ();
 sg13g2_fill_1 FILLER_62_173 ();
 sg13g2_decap_4 FILLER_62_178 ();
 sg13g2_fill_1 FILLER_62_182 ();
 sg13g2_decap_8 FILLER_62_200 ();
 sg13g2_fill_1 FILLER_62_207 ();
 sg13g2_fill_1 FILLER_62_236 ();
 sg13g2_fill_2 FILLER_62_252 ();
 sg13g2_fill_1 FILLER_62_254 ();
 sg13g2_fill_2 FILLER_62_273 ();
 sg13g2_fill_1 FILLER_62_275 ();
 sg13g2_decap_8 FILLER_62_294 ();
 sg13g2_fill_2 FILLER_62_301 ();
 sg13g2_decap_8 FILLER_62_308 ();
 sg13g2_decap_8 FILLER_62_315 ();
 sg13g2_fill_1 FILLER_62_322 ();
 sg13g2_decap_8 FILLER_62_333 ();
 sg13g2_decap_4 FILLER_62_340 ();
 sg13g2_fill_1 FILLER_62_344 ();
 sg13g2_fill_2 FILLER_62_349 ();
 sg13g2_fill_1 FILLER_62_354 ();
 sg13g2_fill_2 FILLER_62_369 ();
 sg13g2_fill_1 FILLER_62_371 ();
 sg13g2_fill_2 FILLER_62_376 ();
 sg13g2_decap_8 FILLER_62_386 ();
 sg13g2_fill_1 FILLER_62_393 ();
 sg13g2_decap_4 FILLER_62_407 ();
 sg13g2_fill_1 FILLER_62_411 ();
 sg13g2_fill_1 FILLER_62_434 ();
 sg13g2_fill_2 FILLER_62_465 ();
 sg13g2_fill_2 FILLER_62_492 ();
 sg13g2_fill_2 FILLER_62_525 ();
 sg13g2_fill_1 FILLER_62_535 ();
 sg13g2_fill_2 FILLER_62_541 ();
 sg13g2_fill_1 FILLER_62_543 ();
 sg13g2_fill_2 FILLER_62_583 ();
 sg13g2_fill_1 FILLER_62_585 ();
 sg13g2_fill_1 FILLER_62_594 ();
 sg13g2_decap_4 FILLER_62_607 ();
 sg13g2_fill_1 FILLER_62_611 ();
 sg13g2_decap_8 FILLER_62_638 ();
 sg13g2_fill_2 FILLER_62_645 ();
 sg13g2_fill_2 FILLER_62_656 ();
 sg13g2_fill_1 FILLER_62_663 ();
 sg13g2_decap_8 FILLER_62_670 ();
 sg13g2_fill_2 FILLER_62_682 ();
 sg13g2_fill_1 FILLER_62_697 ();
 sg13g2_fill_2 FILLER_62_736 ();
 sg13g2_fill_1 FILLER_62_738 ();
 sg13g2_decap_8 FILLER_62_752 ();
 sg13g2_decap_8 FILLER_62_759 ();
 sg13g2_decap_8 FILLER_62_766 ();
 sg13g2_decap_8 FILLER_62_773 ();
 sg13g2_decap_8 FILLER_62_780 ();
 sg13g2_decap_8 FILLER_62_787 ();
 sg13g2_decap_8 FILLER_62_794 ();
 sg13g2_decap_8 FILLER_62_801 ();
 sg13g2_decap_8 FILLER_62_808 ();
 sg13g2_decap_8 FILLER_62_815 ();
 sg13g2_decap_8 FILLER_62_822 ();
 sg13g2_decap_8 FILLER_62_829 ();
 sg13g2_decap_8 FILLER_62_836 ();
 sg13g2_decap_8 FILLER_62_843 ();
 sg13g2_decap_8 FILLER_62_850 ();
 sg13g2_decap_4 FILLER_62_857 ();
 sg13g2_fill_1 FILLER_62_861 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_33 ();
 sg13g2_decap_4 FILLER_63_40 ();
 sg13g2_fill_1 FILLER_63_44 ();
 sg13g2_fill_2 FILLER_63_82 ();
 sg13g2_fill_1 FILLER_63_84 ();
 sg13g2_fill_2 FILLER_63_102 ();
 sg13g2_fill_1 FILLER_63_108 ();
 sg13g2_fill_2 FILLER_63_118 ();
 sg13g2_fill_2 FILLER_63_126 ();
 sg13g2_fill_1 FILLER_63_148 ();
 sg13g2_decap_8 FILLER_63_169 ();
 sg13g2_fill_1 FILLER_63_176 ();
 sg13g2_decap_8 FILLER_63_200 ();
 sg13g2_fill_2 FILLER_63_207 ();
 sg13g2_fill_1 FILLER_63_209 ();
 sg13g2_decap_8 FILLER_63_215 ();
 sg13g2_decap_8 FILLER_63_246 ();
 sg13g2_fill_1 FILLER_63_253 ();
 sg13g2_decap_4 FILLER_63_258 ();
 sg13g2_fill_1 FILLER_63_262 ();
 sg13g2_decap_4 FILLER_63_267 ();
 sg13g2_fill_1 FILLER_63_271 ();
 sg13g2_fill_2 FILLER_63_290 ();
 sg13g2_fill_2 FILLER_63_302 ();
 sg13g2_fill_2 FILLER_63_317 ();
 sg13g2_fill_1 FILLER_63_319 ();
 sg13g2_fill_1 FILLER_63_343 ();
 sg13g2_fill_1 FILLER_63_393 ();
 sg13g2_decap_4 FILLER_63_426 ();
 sg13g2_fill_1 FILLER_63_430 ();
 sg13g2_decap_4 FILLER_63_436 ();
 sg13g2_decap_8 FILLER_63_466 ();
 sg13g2_fill_2 FILLER_63_473 ();
 sg13g2_decap_8 FILLER_63_481 ();
 sg13g2_fill_2 FILLER_63_496 ();
 sg13g2_fill_2 FILLER_63_510 ();
 sg13g2_fill_1 FILLER_63_516 ();
 sg13g2_fill_2 FILLER_63_525 ();
 sg13g2_fill_1 FILLER_63_527 ();
 sg13g2_decap_4 FILLER_63_563 ();
 sg13g2_decap_8 FILLER_63_572 ();
 sg13g2_fill_1 FILLER_63_579 ();
 sg13g2_decap_8 FILLER_63_603 ();
 sg13g2_fill_2 FILLER_63_610 ();
 sg13g2_decap_4 FILLER_63_616 ();
 sg13g2_fill_1 FILLER_63_620 ();
 sg13g2_decap_4 FILLER_63_631 ();
 sg13g2_fill_2 FILLER_63_635 ();
 sg13g2_fill_2 FILLER_63_645 ();
 sg13g2_fill_1 FILLER_63_647 ();
 sg13g2_fill_2 FILLER_63_656 ();
 sg13g2_fill_1 FILLER_63_658 ();
 sg13g2_fill_2 FILLER_63_675 ();
 sg13g2_fill_1 FILLER_63_677 ();
 sg13g2_fill_2 FILLER_63_686 ();
 sg13g2_decap_8 FILLER_63_704 ();
 sg13g2_fill_2 FILLER_63_711 ();
 sg13g2_decap_8 FILLER_63_749 ();
 sg13g2_decap_8 FILLER_63_756 ();
 sg13g2_decap_8 FILLER_63_763 ();
 sg13g2_decap_8 FILLER_63_770 ();
 sg13g2_decap_8 FILLER_63_777 ();
 sg13g2_decap_8 FILLER_63_784 ();
 sg13g2_decap_8 FILLER_63_791 ();
 sg13g2_decap_8 FILLER_63_798 ();
 sg13g2_decap_8 FILLER_63_805 ();
 sg13g2_decap_8 FILLER_63_812 ();
 sg13g2_decap_8 FILLER_63_819 ();
 sg13g2_decap_8 FILLER_63_826 ();
 sg13g2_decap_8 FILLER_63_833 ();
 sg13g2_decap_8 FILLER_63_840 ();
 sg13g2_decap_8 FILLER_63_847 ();
 sg13g2_decap_8 FILLER_63_854 ();
 sg13g2_fill_1 FILLER_63_861 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_4 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_26 ();
 sg13g2_fill_2 FILLER_64_33 ();
 sg13g2_fill_1 FILLER_64_66 ();
 sg13g2_fill_2 FILLER_64_72 ();
 sg13g2_fill_1 FILLER_64_88 ();
 sg13g2_decap_4 FILLER_64_107 ();
 sg13g2_fill_2 FILLER_64_126 ();
 sg13g2_fill_1 FILLER_64_128 ();
 sg13g2_decap_4 FILLER_64_134 ();
 sg13g2_fill_1 FILLER_64_138 ();
 sg13g2_fill_1 FILLER_64_143 ();
 sg13g2_fill_2 FILLER_64_147 ();
 sg13g2_fill_1 FILLER_64_149 ();
 sg13g2_fill_2 FILLER_64_167 ();
 sg13g2_decap_4 FILLER_64_179 ();
 sg13g2_fill_2 FILLER_64_183 ();
 sg13g2_decap_4 FILLER_64_198 ();
 sg13g2_decap_4 FILLER_64_208 ();
 sg13g2_decap_8 FILLER_64_218 ();
 sg13g2_fill_2 FILLER_64_235 ();
 sg13g2_fill_1 FILLER_64_247 ();
 sg13g2_fill_2 FILLER_64_283 ();
 sg13g2_decap_4 FILLER_64_295 ();
 sg13g2_fill_2 FILLER_64_299 ();
 sg13g2_fill_1 FILLER_64_305 ();
 sg13g2_fill_2 FILLER_64_319 ();
 sg13g2_fill_2 FILLER_64_330 ();
 sg13g2_fill_1 FILLER_64_332 ();
 sg13g2_fill_1 FILLER_64_338 ();
 sg13g2_fill_2 FILLER_64_348 ();
 sg13g2_decap_8 FILLER_64_368 ();
 sg13g2_fill_2 FILLER_64_375 ();
 sg13g2_decap_4 FILLER_64_390 ();
 sg13g2_fill_2 FILLER_64_394 ();
 sg13g2_fill_1 FILLER_64_405 ();
 sg13g2_decap_8 FILLER_64_416 ();
 sg13g2_decap_8 FILLER_64_423 ();
 sg13g2_decap_4 FILLER_64_456 ();
 sg13g2_fill_1 FILLER_64_460 ();
 sg13g2_fill_2 FILLER_64_469 ();
 sg13g2_fill_1 FILLER_64_471 ();
 sg13g2_fill_1 FILLER_64_494 ();
 sg13g2_fill_2 FILLER_64_507 ();
 sg13g2_fill_1 FILLER_64_509 ();
 sg13g2_decap_8 FILLER_64_518 ();
 sg13g2_decap_4 FILLER_64_525 ();
 sg13g2_fill_1 FILLER_64_529 ();
 sg13g2_decap_4 FILLER_64_535 ();
 sg13g2_fill_2 FILLER_64_544 ();
 sg13g2_fill_1 FILLER_64_546 ();
 sg13g2_fill_2 FILLER_64_560 ();
 sg13g2_decap_8 FILLER_64_567 ();
 sg13g2_fill_2 FILLER_64_574 ();
 sg13g2_fill_1 FILLER_64_576 ();
 sg13g2_decap_8 FILLER_64_600 ();
 sg13g2_fill_2 FILLER_64_607 ();
 sg13g2_fill_1 FILLER_64_609 ();
 sg13g2_decap_4 FILLER_64_634 ();
 sg13g2_decap_4 FILLER_64_645 ();
 sg13g2_fill_1 FILLER_64_649 ();
 sg13g2_decap_8 FILLER_64_671 ();
 sg13g2_fill_1 FILLER_64_678 ();
 sg13g2_decap_8 FILLER_64_700 ();
 sg13g2_fill_1 FILLER_64_707 ();
 sg13g2_decap_8 FILLER_64_729 ();
 sg13g2_decap_8 FILLER_64_754 ();
 sg13g2_decap_8 FILLER_64_761 ();
 sg13g2_decap_8 FILLER_64_768 ();
 sg13g2_decap_8 FILLER_64_775 ();
 sg13g2_decap_8 FILLER_64_782 ();
 sg13g2_decap_8 FILLER_64_789 ();
 sg13g2_decap_8 FILLER_64_796 ();
 sg13g2_decap_8 FILLER_64_803 ();
 sg13g2_decap_8 FILLER_64_810 ();
 sg13g2_decap_8 FILLER_64_817 ();
 sg13g2_decap_8 FILLER_64_824 ();
 sg13g2_decap_8 FILLER_64_831 ();
 sg13g2_decap_8 FILLER_64_838 ();
 sg13g2_decap_8 FILLER_64_845 ();
 sg13g2_decap_8 FILLER_64_852 ();
 sg13g2_fill_2 FILLER_64_859 ();
 sg13g2_fill_1 FILLER_64_861 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_fill_1 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_38 ();
 sg13g2_fill_1 FILLER_65_45 ();
 sg13g2_decap_8 FILLER_65_50 ();
 sg13g2_fill_1 FILLER_65_57 ();
 sg13g2_fill_2 FILLER_65_66 ();
 sg13g2_fill_1 FILLER_65_68 ();
 sg13g2_fill_2 FILLER_65_82 ();
 sg13g2_fill_2 FILLER_65_120 ();
 sg13g2_fill_1 FILLER_65_132 ();
 sg13g2_fill_2 FILLER_65_142 ();
 sg13g2_fill_1 FILLER_65_144 ();
 sg13g2_decap_8 FILLER_65_155 ();
 sg13g2_fill_1 FILLER_65_162 ();
 sg13g2_fill_2 FILLER_65_176 ();
 sg13g2_fill_1 FILLER_65_178 ();
 sg13g2_decap_4 FILLER_65_206 ();
 sg13g2_decap_8 FILLER_65_232 ();
 sg13g2_fill_2 FILLER_65_248 ();
 sg13g2_fill_1 FILLER_65_250 ();
 sg13g2_fill_1 FILLER_65_255 ();
 sg13g2_decap_4 FILLER_65_264 ();
 sg13g2_fill_2 FILLER_65_280 ();
 sg13g2_decap_8 FILLER_65_287 ();
 sg13g2_fill_2 FILLER_65_294 ();
 sg13g2_fill_2 FILLER_65_326 ();
 sg13g2_fill_2 FILLER_65_337 ();
 sg13g2_decap_4 FILLER_65_357 ();
 sg13g2_fill_1 FILLER_65_375 ();
 sg13g2_fill_1 FILLER_65_386 ();
 sg13g2_fill_2 FILLER_65_392 ();
 sg13g2_decap_8 FILLER_65_424 ();
 sg13g2_fill_1 FILLER_65_439 ();
 sg13g2_decap_8 FILLER_65_450 ();
 sg13g2_decap_8 FILLER_65_457 ();
 sg13g2_fill_2 FILLER_65_464 ();
 sg13g2_decap_8 FILLER_65_486 ();
 sg13g2_fill_1 FILLER_65_493 ();
 sg13g2_fill_2 FILLER_65_503 ();
 sg13g2_fill_1 FILLER_65_517 ();
 sg13g2_fill_2 FILLER_65_560 ();
 sg13g2_fill_1 FILLER_65_562 ();
 sg13g2_fill_2 FILLER_65_568 ();
 sg13g2_decap_4 FILLER_65_591 ();
 sg13g2_fill_2 FILLER_65_595 ();
 sg13g2_fill_2 FILLER_65_617 ();
 sg13g2_fill_1 FILLER_65_636 ();
 sg13g2_decap_8 FILLER_65_674 ();
 sg13g2_fill_2 FILLER_65_681 ();
 sg13g2_fill_1 FILLER_65_683 ();
 sg13g2_fill_2 FILLER_65_692 ();
 sg13g2_fill_1 FILLER_65_702 ();
 sg13g2_decap_8 FILLER_65_720 ();
 sg13g2_fill_2 FILLER_65_727 ();
 sg13g2_decap_8 FILLER_65_760 ();
 sg13g2_decap_8 FILLER_65_767 ();
 sg13g2_decap_8 FILLER_65_774 ();
 sg13g2_decap_8 FILLER_65_781 ();
 sg13g2_decap_8 FILLER_65_788 ();
 sg13g2_decap_8 FILLER_65_795 ();
 sg13g2_decap_8 FILLER_65_802 ();
 sg13g2_decap_8 FILLER_65_809 ();
 sg13g2_decap_8 FILLER_65_816 ();
 sg13g2_decap_8 FILLER_65_823 ();
 sg13g2_decap_8 FILLER_65_830 ();
 sg13g2_decap_8 FILLER_65_837 ();
 sg13g2_decap_8 FILLER_65_844 ();
 sg13g2_decap_8 FILLER_65_851 ();
 sg13g2_decap_4 FILLER_65_858 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_fill_2 FILLER_66_21 ();
 sg13g2_fill_1 FILLER_66_49 ();
 sg13g2_fill_2 FILLER_66_72 ();
 sg13g2_fill_1 FILLER_66_74 ();
 sg13g2_fill_2 FILLER_66_85 ();
 sg13g2_fill_1 FILLER_66_87 ();
 sg13g2_decap_8 FILLER_66_109 ();
 sg13g2_decap_4 FILLER_66_116 ();
 sg13g2_fill_2 FILLER_66_120 ();
 sg13g2_fill_2 FILLER_66_131 ();
 sg13g2_fill_1 FILLER_66_133 ();
 sg13g2_fill_2 FILLER_66_154 ();
 sg13g2_decap_4 FILLER_66_166 ();
 sg13g2_fill_2 FILLER_66_186 ();
 sg13g2_fill_2 FILLER_66_193 ();
 sg13g2_fill_1 FILLER_66_195 ();
 sg13g2_decap_4 FILLER_66_204 ();
 sg13g2_fill_1 FILLER_66_208 ();
 sg13g2_fill_2 FILLER_66_227 ();
 sg13g2_fill_1 FILLER_66_238 ();
 sg13g2_fill_2 FILLER_66_257 ();
 sg13g2_fill_1 FILLER_66_269 ();
 sg13g2_decap_8 FILLER_66_295 ();
 sg13g2_fill_2 FILLER_66_302 ();
 sg13g2_fill_2 FILLER_66_309 ();
 sg13g2_decap_4 FILLER_66_319 ();
 sg13g2_fill_2 FILLER_66_323 ();
 sg13g2_decap_8 FILLER_66_343 ();
 sg13g2_fill_2 FILLER_66_350 ();
 sg13g2_decap_8 FILLER_66_391 ();
 sg13g2_decap_4 FILLER_66_398 ();
 sg13g2_fill_2 FILLER_66_402 ();
 sg13g2_fill_2 FILLER_66_408 ();
 sg13g2_decap_4 FILLER_66_415 ();
 sg13g2_fill_1 FILLER_66_419 ();
 sg13g2_decap_4 FILLER_66_465 ();
 sg13g2_fill_1 FILLER_66_469 ();
 sg13g2_decap_4 FILLER_66_488 ();
 sg13g2_fill_1 FILLER_66_492 ();
 sg13g2_decap_4 FILLER_66_498 ();
 sg13g2_fill_1 FILLER_66_502 ();
 sg13g2_fill_1 FILLER_66_524 ();
 sg13g2_decap_8 FILLER_66_536 ();
 sg13g2_decap_4 FILLER_66_556 ();
 sg13g2_fill_2 FILLER_66_571 ();
 sg13g2_decap_8 FILLER_66_585 ();
 sg13g2_decap_8 FILLER_66_592 ();
 sg13g2_decap_4 FILLER_66_599 ();
 sg13g2_decap_8 FILLER_66_615 ();
 sg13g2_fill_1 FILLER_66_622 ();
 sg13g2_decap_4 FILLER_66_645 ();
 sg13g2_fill_1 FILLER_66_649 ();
 sg13g2_fill_2 FILLER_66_671 ();
 sg13g2_fill_1 FILLER_66_673 ();
 sg13g2_fill_2 FILLER_66_691 ();
 sg13g2_decap_4 FILLER_66_701 ();
 sg13g2_fill_1 FILLER_66_705 ();
 sg13g2_fill_1 FILLER_66_711 ();
 sg13g2_fill_2 FILLER_66_716 ();
 sg13g2_fill_1 FILLER_66_718 ();
 sg13g2_decap_8 FILLER_66_724 ();
 sg13g2_fill_2 FILLER_66_739 ();
 sg13g2_decap_8 FILLER_66_751 ();
 sg13g2_decap_8 FILLER_66_758 ();
 sg13g2_decap_8 FILLER_66_765 ();
 sg13g2_decap_8 FILLER_66_772 ();
 sg13g2_decap_8 FILLER_66_779 ();
 sg13g2_decap_8 FILLER_66_786 ();
 sg13g2_decap_8 FILLER_66_793 ();
 sg13g2_decap_8 FILLER_66_800 ();
 sg13g2_decap_8 FILLER_66_807 ();
 sg13g2_decap_8 FILLER_66_814 ();
 sg13g2_decap_8 FILLER_66_821 ();
 sg13g2_decap_8 FILLER_66_828 ();
 sg13g2_decap_8 FILLER_66_835 ();
 sg13g2_decap_8 FILLER_66_842 ();
 sg13g2_decap_8 FILLER_66_849 ();
 sg13g2_decap_4 FILLER_66_856 ();
 sg13g2_fill_2 FILLER_66_860 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_fill_1 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_38 ();
 sg13g2_decap_4 FILLER_67_45 ();
 sg13g2_fill_2 FILLER_67_76 ();
 sg13g2_fill_1 FILLER_67_78 ();
 sg13g2_decap_8 FILLER_67_117 ();
 sg13g2_fill_1 FILLER_67_124 ();
 sg13g2_fill_2 FILLER_67_139 ();
 sg13g2_fill_2 FILLER_67_155 ();
 sg13g2_decap_4 FILLER_67_171 ();
 sg13g2_fill_2 FILLER_67_175 ();
 sg13g2_fill_2 FILLER_67_186 ();
 sg13g2_fill_1 FILLER_67_203 ();
 sg13g2_fill_2 FILLER_67_216 ();
 sg13g2_fill_2 FILLER_67_228 ();
 sg13g2_fill_1 FILLER_67_234 ();
 sg13g2_decap_8 FILLER_67_258 ();
 sg13g2_decap_4 FILLER_67_265 ();
 sg13g2_decap_4 FILLER_67_274 ();
 sg13g2_decap_4 FILLER_67_293 ();
 sg13g2_decap_4 FILLER_67_327 ();
 sg13g2_fill_1 FILLER_67_331 ();
 sg13g2_decap_8 FILLER_67_337 ();
 sg13g2_decap_4 FILLER_67_344 ();
 sg13g2_decap_4 FILLER_67_356 ();
 sg13g2_fill_2 FILLER_67_389 ();
 sg13g2_fill_1 FILLER_67_391 ();
 sg13g2_fill_1 FILLER_67_401 ();
 sg13g2_decap_4 FILLER_67_441 ();
 sg13g2_decap_8 FILLER_67_466 ();
 sg13g2_fill_2 FILLER_67_481 ();
 sg13g2_fill_2 FILLER_67_504 ();
 sg13g2_decap_4 FILLER_67_526 ();
 sg13g2_fill_1 FILLER_67_543 ();
 sg13g2_decap_8 FILLER_67_556 ();
 sg13g2_decap_4 FILLER_67_579 ();
 sg13g2_fill_2 FILLER_67_604 ();
 sg13g2_fill_1 FILLER_67_614 ();
 sg13g2_fill_1 FILLER_67_619 ();
 sg13g2_fill_2 FILLER_67_625 ();
 sg13g2_decap_8 FILLER_67_649 ();
 sg13g2_fill_2 FILLER_67_656 ();
 sg13g2_fill_2 FILLER_67_668 ();
 sg13g2_fill_2 FILLER_67_685 ();
 sg13g2_fill_2 FILLER_67_700 ();
 sg13g2_fill_1 FILLER_67_702 ();
 sg13g2_fill_2 FILLER_67_726 ();
 sg13g2_decap_8 FILLER_67_749 ();
 sg13g2_decap_8 FILLER_67_756 ();
 sg13g2_decap_8 FILLER_67_763 ();
 sg13g2_decap_8 FILLER_67_770 ();
 sg13g2_decap_8 FILLER_67_777 ();
 sg13g2_decap_8 FILLER_67_784 ();
 sg13g2_decap_8 FILLER_67_791 ();
 sg13g2_decap_8 FILLER_67_798 ();
 sg13g2_decap_8 FILLER_67_805 ();
 sg13g2_decap_8 FILLER_67_812 ();
 sg13g2_decap_8 FILLER_67_819 ();
 sg13g2_decap_8 FILLER_67_826 ();
 sg13g2_decap_8 FILLER_67_833 ();
 sg13g2_decap_8 FILLER_67_840 ();
 sg13g2_decap_8 FILLER_67_847 ();
 sg13g2_decap_8 FILLER_67_854 ();
 sg13g2_fill_1 FILLER_67_861 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_72 ();
 sg13g2_decap_4 FILLER_68_79 ();
 sg13g2_fill_1 FILLER_68_87 ();
 sg13g2_fill_2 FILLER_68_92 ();
 sg13g2_fill_2 FILLER_68_98 ();
 sg13g2_decap_4 FILLER_68_108 ();
 sg13g2_fill_2 FILLER_68_129 ();
 sg13g2_fill_1 FILLER_68_131 ();
 sg13g2_decap_8 FILLER_68_137 ();
 sg13g2_fill_1 FILLER_68_144 ();
 sg13g2_fill_2 FILLER_68_168 ();
 sg13g2_fill_1 FILLER_68_183 ();
 sg13g2_fill_2 FILLER_68_214 ();
 sg13g2_fill_2 FILLER_68_298 ();
 sg13g2_fill_1 FILLER_68_300 ();
 sg13g2_decap_4 FILLER_68_304 ();
 sg13g2_fill_1 FILLER_68_308 ();
 sg13g2_decap_4 FILLER_68_319 ();
 sg13g2_fill_1 FILLER_68_323 ();
 sg13g2_fill_1 FILLER_68_338 ();
 sg13g2_decap_8 FILLER_68_359 ();
 sg13g2_fill_2 FILLER_68_366 ();
 sg13g2_fill_1 FILLER_68_368 ();
 sg13g2_fill_1 FILLER_68_374 ();
 sg13g2_fill_1 FILLER_68_388 ();
 sg13g2_fill_1 FILLER_68_394 ();
 sg13g2_fill_2 FILLER_68_420 ();
 sg13g2_fill_1 FILLER_68_422 ();
 sg13g2_decap_8 FILLER_68_465 ();
 sg13g2_decap_8 FILLER_68_472 ();
 sg13g2_decap_8 FILLER_68_479 ();
 sg13g2_fill_2 FILLER_68_490 ();
 sg13g2_fill_1 FILLER_68_492 ();
 sg13g2_decap_4 FILLER_68_498 ();
 sg13g2_fill_2 FILLER_68_502 ();
 sg13g2_decap_4 FILLER_68_508 ();
 sg13g2_fill_1 FILLER_68_512 ();
 sg13g2_fill_2 FILLER_68_523 ();
 sg13g2_fill_2 FILLER_68_557 ();
 sg13g2_fill_2 FILLER_68_579 ();
 sg13g2_fill_1 FILLER_68_626 ();
 sg13g2_decap_8 FILLER_68_643 ();
 sg13g2_fill_2 FILLER_68_650 ();
 sg13g2_fill_1 FILLER_68_652 ();
 sg13g2_decap_4 FILLER_68_674 ();
 sg13g2_decap_8 FILLER_68_704 ();
 sg13g2_decap_8 FILLER_68_711 ();
 sg13g2_decap_8 FILLER_68_718 ();
 sg13g2_decap_8 FILLER_68_725 ();
 sg13g2_decap_8 FILLER_68_732 ();
 sg13g2_decap_8 FILLER_68_739 ();
 sg13g2_decap_8 FILLER_68_746 ();
 sg13g2_decap_8 FILLER_68_753 ();
 sg13g2_decap_8 FILLER_68_760 ();
 sg13g2_decap_8 FILLER_68_767 ();
 sg13g2_decap_8 FILLER_68_774 ();
 sg13g2_decap_8 FILLER_68_781 ();
 sg13g2_decap_8 FILLER_68_788 ();
 sg13g2_decap_8 FILLER_68_795 ();
 sg13g2_decap_8 FILLER_68_802 ();
 sg13g2_decap_8 FILLER_68_809 ();
 sg13g2_decap_8 FILLER_68_816 ();
 sg13g2_decap_8 FILLER_68_823 ();
 sg13g2_decap_8 FILLER_68_830 ();
 sg13g2_decap_8 FILLER_68_837 ();
 sg13g2_decap_8 FILLER_68_844 ();
 sg13g2_decap_8 FILLER_68_851 ();
 sg13g2_decap_4 FILLER_68_858 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_4 FILLER_69_28 ();
 sg13g2_fill_1 FILLER_69_32 ();
 sg13g2_fill_2 FILLER_69_47 ();
 sg13g2_decap_4 FILLER_69_53 ();
 sg13g2_decap_8 FILLER_69_71 ();
 sg13g2_fill_1 FILLER_69_78 ();
 sg13g2_fill_2 FILLER_69_99 ();
 sg13g2_fill_1 FILLER_69_125 ();
 sg13g2_fill_2 FILLER_69_144 ();
 sg13g2_decap_8 FILLER_69_214 ();
 sg13g2_decap_4 FILLER_69_221 ();
 sg13g2_decap_8 FILLER_69_233 ();
 sg13g2_decap_4 FILLER_69_240 ();
 sg13g2_fill_2 FILLER_69_244 ();
 sg13g2_decap_8 FILLER_69_267 ();
 sg13g2_fill_1 FILLER_69_274 ();
 sg13g2_decap_8 FILLER_69_287 ();
 sg13g2_decap_4 FILLER_69_294 ();
 sg13g2_fill_1 FILLER_69_318 ();
 sg13g2_fill_2 FILLER_69_344 ();
 sg13g2_decap_8 FILLER_69_350 ();
 sg13g2_decap_4 FILLER_69_375 ();
 sg13g2_fill_2 FILLER_69_379 ();
 sg13g2_fill_2 FILLER_69_387 ();
 sg13g2_fill_2 FILLER_69_398 ();
 sg13g2_decap_4 FILLER_69_412 ();
 sg13g2_fill_1 FILLER_69_416 ();
 sg13g2_decap_4 FILLER_69_422 ();
 sg13g2_fill_2 FILLER_69_426 ();
 sg13g2_decap_8 FILLER_69_433 ();
 sg13g2_decap_8 FILLER_69_440 ();
 sg13g2_decap_8 FILLER_69_447 ();
 sg13g2_decap_8 FILLER_69_454 ();
 sg13g2_decap_4 FILLER_69_461 ();
 sg13g2_fill_1 FILLER_69_475 ();
 sg13g2_fill_1 FILLER_69_511 ();
 sg13g2_fill_1 FILLER_69_517 ();
 sg13g2_decap_4 FILLER_69_522 ();
 sg13g2_fill_2 FILLER_69_526 ();
 sg13g2_decap_8 FILLER_69_533 ();
 sg13g2_decap_4 FILLER_69_540 ();
 sg13g2_decap_4 FILLER_69_553 ();
 sg13g2_fill_1 FILLER_69_557 ();
 sg13g2_decap_8 FILLER_69_569 ();
 sg13g2_decap_4 FILLER_69_576 ();
 sg13g2_fill_2 FILLER_69_602 ();
 sg13g2_decap_8 FILLER_69_624 ();
 sg13g2_fill_1 FILLER_69_631 ();
 sg13g2_decap_8 FILLER_69_637 ();
 sg13g2_decap_8 FILLER_69_644 ();
 sg13g2_decap_8 FILLER_69_651 ();
 sg13g2_decap_8 FILLER_69_665 ();
 sg13g2_decap_8 FILLER_69_672 ();
 sg13g2_decap_8 FILLER_69_679 ();
 sg13g2_fill_1 FILLER_69_686 ();
 sg13g2_decap_8 FILLER_69_696 ();
 sg13g2_decap_8 FILLER_69_703 ();
 sg13g2_decap_8 FILLER_69_710 ();
 sg13g2_decap_8 FILLER_69_717 ();
 sg13g2_decap_8 FILLER_69_724 ();
 sg13g2_decap_8 FILLER_69_731 ();
 sg13g2_decap_8 FILLER_69_738 ();
 sg13g2_decap_8 FILLER_69_745 ();
 sg13g2_decap_8 FILLER_69_752 ();
 sg13g2_decap_8 FILLER_69_759 ();
 sg13g2_decap_8 FILLER_69_766 ();
 sg13g2_decap_8 FILLER_69_773 ();
 sg13g2_decap_8 FILLER_69_780 ();
 sg13g2_decap_8 FILLER_69_787 ();
 sg13g2_decap_8 FILLER_69_794 ();
 sg13g2_decap_8 FILLER_69_801 ();
 sg13g2_decap_8 FILLER_69_808 ();
 sg13g2_decap_8 FILLER_69_815 ();
 sg13g2_decap_8 FILLER_69_822 ();
 sg13g2_decap_8 FILLER_69_829 ();
 sg13g2_decap_8 FILLER_69_836 ();
 sg13g2_decap_8 FILLER_69_843 ();
 sg13g2_decap_8 FILLER_69_850 ();
 sg13g2_decap_4 FILLER_69_857 ();
 sg13g2_fill_1 FILLER_69_861 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_fill_2 FILLER_70_28 ();
 sg13g2_fill_2 FILLER_70_82 ();
 sg13g2_fill_1 FILLER_70_84 ();
 sg13g2_fill_1 FILLER_70_89 ();
 sg13g2_decap_8 FILLER_70_111 ();
 sg13g2_decap_4 FILLER_70_118 ();
 sg13g2_decap_4 FILLER_70_126 ();
 sg13g2_fill_1 FILLER_70_130 ();
 sg13g2_decap_8 FILLER_70_139 ();
 sg13g2_fill_1 FILLER_70_146 ();
 sg13g2_decap_4 FILLER_70_168 ();
 sg13g2_fill_1 FILLER_70_172 ();
 sg13g2_decap_4 FILLER_70_194 ();
 sg13g2_fill_2 FILLER_70_219 ();
 sg13g2_fill_1 FILLER_70_226 ();
 sg13g2_decap_8 FILLER_70_237 ();
 sg13g2_fill_2 FILLER_70_244 ();
 sg13g2_fill_1 FILLER_70_246 ();
 sg13g2_fill_2 FILLER_70_251 ();
 sg13g2_fill_2 FILLER_70_257 ();
 sg13g2_fill_1 FILLER_70_259 ();
 sg13g2_decap_4 FILLER_70_264 ();
 sg13g2_fill_1 FILLER_70_268 ();
 sg13g2_decap_4 FILLER_70_276 ();
 sg13g2_decap_8 FILLER_70_288 ();
 sg13g2_fill_2 FILLER_70_323 ();
 sg13g2_fill_1 FILLER_70_325 ();
 sg13g2_decap_4 FILLER_70_336 ();
 sg13g2_fill_2 FILLER_70_340 ();
 sg13g2_fill_1 FILLER_70_351 ();
 sg13g2_decap_8 FILLER_70_361 ();
 sg13g2_decap_8 FILLER_70_368 ();
 sg13g2_fill_1 FILLER_70_375 ();
 sg13g2_fill_2 FILLER_70_389 ();
 sg13g2_decap_4 FILLER_70_412 ();
 sg13g2_decap_4 FILLER_70_424 ();
 sg13g2_fill_1 FILLER_70_428 ();
 sg13g2_decap_4 FILLER_70_453 ();
 sg13g2_fill_2 FILLER_70_457 ();
 sg13g2_fill_2 FILLER_70_475 ();
 sg13g2_fill_1 FILLER_70_477 ();
 sg13g2_fill_2 FILLER_70_486 ();
 sg13g2_fill_1 FILLER_70_503 ();
 sg13g2_fill_2 FILLER_70_520 ();
 sg13g2_decap_8 FILLER_70_574 ();
 sg13g2_fill_2 FILLER_70_581 ();
 sg13g2_decap_8 FILLER_70_592 ();
 sg13g2_decap_4 FILLER_70_599 ();
 sg13g2_fill_2 FILLER_70_603 ();
 sg13g2_decap_8 FILLER_70_608 ();
 sg13g2_decap_8 FILLER_70_615 ();
 sg13g2_decap_8 FILLER_70_622 ();
 sg13g2_decap_8 FILLER_70_629 ();
 sg13g2_decap_8 FILLER_70_636 ();
 sg13g2_decap_8 FILLER_70_643 ();
 sg13g2_decap_8 FILLER_70_650 ();
 sg13g2_decap_8 FILLER_70_657 ();
 sg13g2_decap_8 FILLER_70_664 ();
 sg13g2_decap_8 FILLER_70_671 ();
 sg13g2_decap_8 FILLER_70_678 ();
 sg13g2_decap_8 FILLER_70_685 ();
 sg13g2_decap_8 FILLER_70_692 ();
 sg13g2_decap_8 FILLER_70_699 ();
 sg13g2_decap_8 FILLER_70_706 ();
 sg13g2_decap_8 FILLER_70_713 ();
 sg13g2_decap_8 FILLER_70_720 ();
 sg13g2_decap_8 FILLER_70_727 ();
 sg13g2_decap_8 FILLER_70_734 ();
 sg13g2_decap_8 FILLER_70_741 ();
 sg13g2_decap_8 FILLER_70_748 ();
 sg13g2_decap_8 FILLER_70_755 ();
 sg13g2_decap_8 FILLER_70_762 ();
 sg13g2_decap_8 FILLER_70_769 ();
 sg13g2_decap_8 FILLER_70_776 ();
 sg13g2_decap_8 FILLER_70_783 ();
 sg13g2_decap_8 FILLER_70_790 ();
 sg13g2_decap_8 FILLER_70_797 ();
 sg13g2_decap_8 FILLER_70_804 ();
 sg13g2_decap_8 FILLER_70_811 ();
 sg13g2_decap_8 FILLER_70_818 ();
 sg13g2_decap_8 FILLER_70_825 ();
 sg13g2_decap_8 FILLER_70_832 ();
 sg13g2_decap_8 FILLER_70_839 ();
 sg13g2_decap_8 FILLER_70_846 ();
 sg13g2_decap_8 FILLER_70_853 ();
 sg13g2_fill_2 FILLER_70_860 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_4 FILLER_71_21 ();
 sg13g2_fill_2 FILLER_71_25 ();
 sg13g2_decap_8 FILLER_71_53 ();
 sg13g2_decap_8 FILLER_71_60 ();
 sg13g2_fill_2 FILLER_71_67 ();
 sg13g2_decap_8 FILLER_71_73 ();
 sg13g2_decap_8 FILLER_71_80 ();
 sg13g2_decap_4 FILLER_71_87 ();
 sg13g2_fill_1 FILLER_71_125 ();
 sg13g2_fill_2 FILLER_71_134 ();
 sg13g2_decap_8 FILLER_71_171 ();
 sg13g2_decap_8 FILLER_71_178 ();
 sg13g2_fill_2 FILLER_71_185 ();
 sg13g2_decap_8 FILLER_71_192 ();
 sg13g2_decap_8 FILLER_71_199 ();
 sg13g2_decap_8 FILLER_71_206 ();
 sg13g2_decap_4 FILLER_71_213 ();
 sg13g2_fill_2 FILLER_71_243 ();
 sg13g2_fill_2 FILLER_71_299 ();
 sg13g2_fill_2 FILLER_71_317 ();
 sg13g2_fill_1 FILLER_71_319 ();
 sg13g2_decap_4 FILLER_71_328 ();
 sg13g2_fill_2 FILLER_71_332 ();
 sg13g2_fill_2 FILLER_71_367 ();
 sg13g2_fill_1 FILLER_71_369 ();
 sg13g2_decap_8 FILLER_71_393 ();
 sg13g2_fill_1 FILLER_71_400 ();
 sg13g2_decap_4 FILLER_71_456 ();
 sg13g2_decap_4 FILLER_71_470 ();
 sg13g2_fill_1 FILLER_71_474 ();
 sg13g2_fill_2 FILLER_71_484 ();
 sg13g2_decap_4 FILLER_71_492 ();
 sg13g2_fill_1 FILLER_71_496 ();
 sg13g2_fill_2 FILLER_71_502 ();
 sg13g2_fill_2 FILLER_71_510 ();
 sg13g2_fill_1 FILLER_71_512 ();
 sg13g2_fill_1 FILLER_71_518 ();
 sg13g2_decap_4 FILLER_71_550 ();
 sg13g2_decap_8 FILLER_71_558 ();
 sg13g2_decap_8 FILLER_71_565 ();
 sg13g2_decap_8 FILLER_71_572 ();
 sg13g2_decap_8 FILLER_71_579 ();
 sg13g2_decap_8 FILLER_71_586 ();
 sg13g2_decap_8 FILLER_71_593 ();
 sg13g2_decap_8 FILLER_71_600 ();
 sg13g2_decap_8 FILLER_71_607 ();
 sg13g2_decap_8 FILLER_71_614 ();
 sg13g2_decap_8 FILLER_71_621 ();
 sg13g2_decap_8 FILLER_71_628 ();
 sg13g2_decap_8 FILLER_71_635 ();
 sg13g2_decap_8 FILLER_71_642 ();
 sg13g2_decap_8 FILLER_71_649 ();
 sg13g2_decap_8 FILLER_71_656 ();
 sg13g2_decap_8 FILLER_71_663 ();
 sg13g2_decap_8 FILLER_71_670 ();
 sg13g2_decap_8 FILLER_71_677 ();
 sg13g2_decap_8 FILLER_71_684 ();
 sg13g2_decap_8 FILLER_71_691 ();
 sg13g2_decap_8 FILLER_71_698 ();
 sg13g2_decap_8 FILLER_71_705 ();
 sg13g2_decap_8 FILLER_71_712 ();
 sg13g2_decap_8 FILLER_71_719 ();
 sg13g2_decap_8 FILLER_71_726 ();
 sg13g2_decap_8 FILLER_71_733 ();
 sg13g2_decap_8 FILLER_71_740 ();
 sg13g2_decap_8 FILLER_71_747 ();
 sg13g2_decap_8 FILLER_71_754 ();
 sg13g2_decap_8 FILLER_71_761 ();
 sg13g2_decap_8 FILLER_71_768 ();
 sg13g2_decap_8 FILLER_71_775 ();
 sg13g2_decap_8 FILLER_71_782 ();
 sg13g2_decap_8 FILLER_71_789 ();
 sg13g2_decap_8 FILLER_71_796 ();
 sg13g2_decap_8 FILLER_71_803 ();
 sg13g2_decap_8 FILLER_71_810 ();
 sg13g2_decap_8 FILLER_71_817 ();
 sg13g2_decap_8 FILLER_71_824 ();
 sg13g2_decap_8 FILLER_71_831 ();
 sg13g2_decap_8 FILLER_71_838 ();
 sg13g2_decap_8 FILLER_71_845 ();
 sg13g2_decap_8 FILLER_71_852 ();
 sg13g2_fill_2 FILLER_71_859 ();
 sg13g2_fill_1 FILLER_71_861 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_fill_2 FILLER_72_35 ();
 sg13g2_fill_1 FILLER_72_37 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_fill_2 FILLER_72_56 ();
 sg13g2_fill_1 FILLER_72_84 ();
 sg13g2_fill_1 FILLER_72_98 ();
 sg13g2_fill_1 FILLER_72_116 ();
 sg13g2_fill_1 FILLER_72_122 ();
 sg13g2_fill_2 FILLER_72_152 ();
 sg13g2_fill_1 FILLER_72_154 ();
 sg13g2_decap_8 FILLER_72_165 ();
 sg13g2_decap_8 FILLER_72_172 ();
 sg13g2_decap_4 FILLER_72_179 ();
 sg13g2_fill_2 FILLER_72_197 ();
 sg13g2_fill_1 FILLER_72_199 ();
 sg13g2_decap_8 FILLER_72_217 ();
 sg13g2_fill_1 FILLER_72_229 ();
 sg13g2_decap_4 FILLER_72_239 ();
 sg13g2_fill_1 FILLER_72_243 ();
 sg13g2_fill_1 FILLER_72_257 ();
 sg13g2_decap_8 FILLER_72_262 ();
 sg13g2_decap_4 FILLER_72_269 ();
 sg13g2_decap_4 FILLER_72_307 ();
 sg13g2_fill_1 FILLER_72_311 ();
 sg13g2_decap_8 FILLER_72_322 ();
 sg13g2_decap_4 FILLER_72_329 ();
 sg13g2_fill_1 FILLER_72_333 ();
 sg13g2_decap_4 FILLER_72_344 ();
 sg13g2_fill_2 FILLER_72_362 ();
 sg13g2_decap_8 FILLER_72_391 ();
 sg13g2_fill_2 FILLER_72_406 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_fill_2 FILLER_72_451 ();
 sg13g2_fill_1 FILLER_72_453 ();
 sg13g2_fill_1 FILLER_72_470 ();
 sg13g2_decap_4 FILLER_72_497 ();
 sg13g2_fill_2 FILLER_72_515 ();
 sg13g2_fill_1 FILLER_72_517 ();
 sg13g2_decap_8 FILLER_72_553 ();
 sg13g2_decap_8 FILLER_72_560 ();
 sg13g2_decap_8 FILLER_72_567 ();
 sg13g2_decap_8 FILLER_72_574 ();
 sg13g2_decap_8 FILLER_72_581 ();
 sg13g2_decap_8 FILLER_72_588 ();
 sg13g2_decap_8 FILLER_72_595 ();
 sg13g2_decap_8 FILLER_72_602 ();
 sg13g2_decap_8 FILLER_72_609 ();
 sg13g2_decap_8 FILLER_72_616 ();
 sg13g2_decap_8 FILLER_72_623 ();
 sg13g2_decap_8 FILLER_72_630 ();
 sg13g2_decap_8 FILLER_72_637 ();
 sg13g2_decap_8 FILLER_72_644 ();
 sg13g2_decap_8 FILLER_72_651 ();
 sg13g2_decap_8 FILLER_72_658 ();
 sg13g2_decap_8 FILLER_72_665 ();
 sg13g2_decap_8 FILLER_72_672 ();
 sg13g2_decap_8 FILLER_72_679 ();
 sg13g2_decap_8 FILLER_72_686 ();
 sg13g2_decap_8 FILLER_72_693 ();
 sg13g2_decap_8 FILLER_72_700 ();
 sg13g2_decap_8 FILLER_72_707 ();
 sg13g2_decap_8 FILLER_72_714 ();
 sg13g2_decap_8 FILLER_72_721 ();
 sg13g2_decap_8 FILLER_72_728 ();
 sg13g2_decap_8 FILLER_72_735 ();
 sg13g2_decap_8 FILLER_72_742 ();
 sg13g2_decap_8 FILLER_72_749 ();
 sg13g2_decap_8 FILLER_72_756 ();
 sg13g2_decap_8 FILLER_72_763 ();
 sg13g2_decap_8 FILLER_72_770 ();
 sg13g2_decap_8 FILLER_72_777 ();
 sg13g2_decap_8 FILLER_72_784 ();
 sg13g2_decap_8 FILLER_72_791 ();
 sg13g2_decap_8 FILLER_72_798 ();
 sg13g2_decap_8 FILLER_72_805 ();
 sg13g2_decap_8 FILLER_72_812 ();
 sg13g2_decap_8 FILLER_72_819 ();
 sg13g2_decap_8 FILLER_72_826 ();
 sg13g2_decap_8 FILLER_72_833 ();
 sg13g2_decap_8 FILLER_72_840 ();
 sg13g2_decap_8 FILLER_72_847 ();
 sg13g2_decap_8 FILLER_72_854 ();
 sg13g2_fill_1 FILLER_72_861 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_4 FILLER_73_84 ();
 sg13g2_fill_1 FILLER_73_88 ();
 sg13g2_fill_2 FILLER_73_106 ();
 sg13g2_fill_2 FILLER_73_129 ();
 sg13g2_fill_1 FILLER_73_131 ();
 sg13g2_fill_2 FILLER_73_138 ();
 sg13g2_decap_4 FILLER_73_144 ();
 sg13g2_fill_2 FILLER_73_148 ();
 sg13g2_decap_8 FILLER_73_163 ();
 sg13g2_decap_4 FILLER_73_170 ();
 sg13g2_fill_2 FILLER_73_174 ();
 sg13g2_fill_1 FILLER_73_215 ();
 sg13g2_fill_2 FILLER_73_225 ();
 sg13g2_fill_1 FILLER_73_227 ();
 sg13g2_fill_2 FILLER_73_233 ();
 sg13g2_fill_1 FILLER_73_235 ();
 sg13g2_fill_1 FILLER_73_250 ();
 sg13g2_fill_1 FILLER_73_272 ();
 sg13g2_decap_4 FILLER_73_278 ();
 sg13g2_fill_1 FILLER_73_282 ();
 sg13g2_fill_2 FILLER_73_299 ();
 sg13g2_decap_8 FILLER_73_329 ();
 sg13g2_decap_8 FILLER_73_336 ();
 sg13g2_decap_8 FILLER_73_369 ();
 sg13g2_decap_4 FILLER_73_376 ();
 sg13g2_decap_4 FILLER_73_422 ();
 sg13g2_fill_1 FILLER_73_426 ();
 sg13g2_decap_8 FILLER_73_431 ();
 sg13g2_decap_8 FILLER_73_438 ();
 sg13g2_decap_4 FILLER_73_445 ();
 sg13g2_fill_1 FILLER_73_461 ();
 sg13g2_fill_1 FILLER_73_471 ();
 sg13g2_fill_2 FILLER_73_476 ();
 sg13g2_fill_2 FILLER_73_496 ();
 sg13g2_fill_2 FILLER_73_512 ();
 sg13g2_decap_8 FILLER_73_549 ();
 sg13g2_decap_8 FILLER_73_556 ();
 sg13g2_decap_8 FILLER_73_563 ();
 sg13g2_decap_8 FILLER_73_570 ();
 sg13g2_decap_8 FILLER_73_577 ();
 sg13g2_decap_8 FILLER_73_584 ();
 sg13g2_decap_8 FILLER_73_591 ();
 sg13g2_decap_8 FILLER_73_598 ();
 sg13g2_decap_8 FILLER_73_605 ();
 sg13g2_decap_8 FILLER_73_612 ();
 sg13g2_decap_8 FILLER_73_619 ();
 sg13g2_decap_8 FILLER_73_626 ();
 sg13g2_decap_8 FILLER_73_633 ();
 sg13g2_decap_8 FILLER_73_640 ();
 sg13g2_decap_8 FILLER_73_647 ();
 sg13g2_decap_8 FILLER_73_654 ();
 sg13g2_decap_8 FILLER_73_661 ();
 sg13g2_decap_8 FILLER_73_668 ();
 sg13g2_decap_8 FILLER_73_675 ();
 sg13g2_decap_8 FILLER_73_682 ();
 sg13g2_decap_8 FILLER_73_689 ();
 sg13g2_decap_8 FILLER_73_696 ();
 sg13g2_decap_8 FILLER_73_703 ();
 sg13g2_decap_8 FILLER_73_710 ();
 sg13g2_decap_8 FILLER_73_717 ();
 sg13g2_decap_8 FILLER_73_724 ();
 sg13g2_decap_8 FILLER_73_731 ();
 sg13g2_decap_8 FILLER_73_738 ();
 sg13g2_decap_8 FILLER_73_745 ();
 sg13g2_decap_8 FILLER_73_752 ();
 sg13g2_decap_8 FILLER_73_759 ();
 sg13g2_decap_8 FILLER_73_766 ();
 sg13g2_decap_8 FILLER_73_773 ();
 sg13g2_decap_8 FILLER_73_780 ();
 sg13g2_decap_8 FILLER_73_787 ();
 sg13g2_decap_8 FILLER_73_794 ();
 sg13g2_decap_8 FILLER_73_801 ();
 sg13g2_decap_8 FILLER_73_808 ();
 sg13g2_decap_8 FILLER_73_815 ();
 sg13g2_decap_8 FILLER_73_822 ();
 sg13g2_decap_8 FILLER_73_829 ();
 sg13g2_decap_8 FILLER_73_836 ();
 sg13g2_decap_8 FILLER_73_843 ();
 sg13g2_decap_8 FILLER_73_850 ();
 sg13g2_decap_4 FILLER_73_857 ();
 sg13g2_fill_1 FILLER_73_861 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_4 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_99 ();
 sg13g2_fill_2 FILLER_74_106 ();
 sg13g2_fill_2 FILLER_74_129 ();
 sg13g2_fill_2 FILLER_74_167 ();
 sg13g2_fill_1 FILLER_74_187 ();
 sg13g2_decap_4 FILLER_74_194 ();
 sg13g2_fill_1 FILLER_74_198 ();
 sg13g2_fill_1 FILLER_74_207 ();
 sg13g2_fill_2 FILLER_74_214 ();
 sg13g2_fill_1 FILLER_74_216 ();
 sg13g2_decap_8 FILLER_74_228 ();
 sg13g2_fill_2 FILLER_74_235 ();
 sg13g2_fill_2 FILLER_74_254 ();
 sg13g2_fill_2 FILLER_74_261 ();
 sg13g2_fill_1 FILLER_74_269 ();
 sg13g2_fill_2 FILLER_74_277 ();
 sg13g2_decap_8 FILLER_74_296 ();
 sg13g2_fill_2 FILLER_74_303 ();
 sg13g2_fill_2 FILLER_74_316 ();
 sg13g2_decap_8 FILLER_74_324 ();
 sg13g2_decap_4 FILLER_74_331 ();
 sg13g2_fill_1 FILLER_74_335 ();
 sg13g2_fill_1 FILLER_74_353 ();
 sg13g2_fill_2 FILLER_74_359 ();
 sg13g2_fill_1 FILLER_74_361 ();
 sg13g2_decap_8 FILLER_74_366 ();
 sg13g2_decap_8 FILLER_74_373 ();
 sg13g2_fill_2 FILLER_74_380 ();
 sg13g2_fill_1 FILLER_74_382 ();
 sg13g2_fill_2 FILLER_74_393 ();
 sg13g2_fill_1 FILLER_74_395 ();
 sg13g2_decap_4 FILLER_74_399 ();
 sg13g2_fill_2 FILLER_74_403 ();
 sg13g2_fill_2 FILLER_74_441 ();
 sg13g2_fill_1 FILLER_74_443 ();
 sg13g2_decap_8 FILLER_74_492 ();
 sg13g2_fill_1 FILLER_74_533 ();
 sg13g2_decap_8 FILLER_74_538 ();
 sg13g2_decap_8 FILLER_74_545 ();
 sg13g2_decap_8 FILLER_74_552 ();
 sg13g2_decap_8 FILLER_74_559 ();
 sg13g2_decap_8 FILLER_74_566 ();
 sg13g2_decap_8 FILLER_74_573 ();
 sg13g2_decap_8 FILLER_74_580 ();
 sg13g2_decap_8 FILLER_74_587 ();
 sg13g2_decap_8 FILLER_74_594 ();
 sg13g2_decap_8 FILLER_74_601 ();
 sg13g2_decap_8 FILLER_74_608 ();
 sg13g2_decap_8 FILLER_74_615 ();
 sg13g2_decap_8 FILLER_74_622 ();
 sg13g2_decap_8 FILLER_74_629 ();
 sg13g2_decap_8 FILLER_74_636 ();
 sg13g2_decap_8 FILLER_74_643 ();
 sg13g2_decap_8 FILLER_74_650 ();
 sg13g2_decap_8 FILLER_74_657 ();
 sg13g2_decap_8 FILLER_74_664 ();
 sg13g2_decap_8 FILLER_74_671 ();
 sg13g2_decap_8 FILLER_74_678 ();
 sg13g2_decap_8 FILLER_74_685 ();
 sg13g2_decap_8 FILLER_74_692 ();
 sg13g2_decap_8 FILLER_74_699 ();
 sg13g2_decap_8 FILLER_74_706 ();
 sg13g2_decap_8 FILLER_74_713 ();
 sg13g2_decap_8 FILLER_74_720 ();
 sg13g2_decap_8 FILLER_74_727 ();
 sg13g2_decap_8 FILLER_74_734 ();
 sg13g2_decap_8 FILLER_74_741 ();
 sg13g2_decap_8 FILLER_74_748 ();
 sg13g2_decap_8 FILLER_74_755 ();
 sg13g2_decap_8 FILLER_74_762 ();
 sg13g2_decap_8 FILLER_74_769 ();
 sg13g2_decap_8 FILLER_74_776 ();
 sg13g2_decap_8 FILLER_74_783 ();
 sg13g2_decap_8 FILLER_74_790 ();
 sg13g2_decap_8 FILLER_74_797 ();
 sg13g2_decap_8 FILLER_74_804 ();
 sg13g2_decap_8 FILLER_74_811 ();
 sg13g2_decap_8 FILLER_74_818 ();
 sg13g2_decap_8 FILLER_74_825 ();
 sg13g2_decap_8 FILLER_74_832 ();
 sg13g2_decap_8 FILLER_74_839 ();
 sg13g2_decap_8 FILLER_74_846 ();
 sg13g2_decap_8 FILLER_74_853 ();
 sg13g2_fill_2 FILLER_74_860 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_117 ();
 sg13g2_decap_8 FILLER_75_124 ();
 sg13g2_fill_1 FILLER_75_131 ();
 sg13g2_fill_2 FILLER_75_137 ();
 sg13g2_fill_1 FILLER_75_148 ();
 sg13g2_decap_8 FILLER_75_164 ();
 sg13g2_fill_2 FILLER_75_171 ();
 sg13g2_fill_1 FILLER_75_173 ();
 sg13g2_decap_4 FILLER_75_195 ();
 sg13g2_fill_1 FILLER_75_199 ();
 sg13g2_fill_1 FILLER_75_208 ();
 sg13g2_decap_8 FILLER_75_213 ();
 sg13g2_fill_2 FILLER_75_220 ();
 sg13g2_decap_8 FILLER_75_239 ();
 sg13g2_fill_2 FILLER_75_246 ();
 sg13g2_fill_1 FILLER_75_248 ();
 sg13g2_fill_1 FILLER_75_254 ();
 sg13g2_decap_8 FILLER_75_268 ();
 sg13g2_fill_1 FILLER_75_275 ();
 sg13g2_decap_8 FILLER_75_280 ();
 sg13g2_fill_2 FILLER_75_287 ();
 sg13g2_fill_1 FILLER_75_289 ();
 sg13g2_decap_8 FILLER_75_377 ();
 sg13g2_fill_1 FILLER_75_384 ();
 sg13g2_decap_8 FILLER_75_405 ();
 sg13g2_decap_4 FILLER_75_412 ();
 sg13g2_decap_4 FILLER_75_420 ();
 sg13g2_fill_1 FILLER_75_424 ();
 sg13g2_fill_1 FILLER_75_429 ();
 sg13g2_fill_2 FILLER_75_434 ();
 sg13g2_fill_1 FILLER_75_436 ();
 sg13g2_fill_2 FILLER_75_444 ();
 sg13g2_fill_2 FILLER_75_452 ();
 sg13g2_fill_2 FILLER_75_464 ();
 sg13g2_fill_1 FILLER_75_466 ();
 sg13g2_decap_4 FILLER_75_507 ();
 sg13g2_fill_2 FILLER_75_511 ();
 sg13g2_fill_2 FILLER_75_517 ();
 sg13g2_decap_8 FILLER_75_528 ();
 sg13g2_decap_8 FILLER_75_535 ();
 sg13g2_decap_8 FILLER_75_542 ();
 sg13g2_decap_8 FILLER_75_549 ();
 sg13g2_decap_8 FILLER_75_556 ();
 sg13g2_decap_8 FILLER_75_563 ();
 sg13g2_decap_8 FILLER_75_570 ();
 sg13g2_decap_8 FILLER_75_577 ();
 sg13g2_decap_8 FILLER_75_584 ();
 sg13g2_decap_8 FILLER_75_591 ();
 sg13g2_decap_8 FILLER_75_598 ();
 sg13g2_decap_8 FILLER_75_605 ();
 sg13g2_decap_8 FILLER_75_612 ();
 sg13g2_decap_8 FILLER_75_619 ();
 sg13g2_decap_8 FILLER_75_626 ();
 sg13g2_decap_8 FILLER_75_633 ();
 sg13g2_decap_8 FILLER_75_640 ();
 sg13g2_decap_8 FILLER_75_647 ();
 sg13g2_decap_8 FILLER_75_654 ();
 sg13g2_decap_8 FILLER_75_661 ();
 sg13g2_decap_8 FILLER_75_668 ();
 sg13g2_decap_8 FILLER_75_675 ();
 sg13g2_decap_8 FILLER_75_682 ();
 sg13g2_decap_8 FILLER_75_689 ();
 sg13g2_decap_8 FILLER_75_696 ();
 sg13g2_decap_8 FILLER_75_703 ();
 sg13g2_decap_8 FILLER_75_710 ();
 sg13g2_decap_8 FILLER_75_717 ();
 sg13g2_decap_8 FILLER_75_724 ();
 sg13g2_decap_8 FILLER_75_731 ();
 sg13g2_decap_8 FILLER_75_738 ();
 sg13g2_decap_8 FILLER_75_745 ();
 sg13g2_decap_8 FILLER_75_752 ();
 sg13g2_decap_8 FILLER_75_759 ();
 sg13g2_decap_8 FILLER_75_766 ();
 sg13g2_decap_8 FILLER_75_773 ();
 sg13g2_decap_8 FILLER_75_780 ();
 sg13g2_decap_8 FILLER_75_787 ();
 sg13g2_decap_8 FILLER_75_794 ();
 sg13g2_decap_8 FILLER_75_801 ();
 sg13g2_decap_8 FILLER_75_808 ();
 sg13g2_decap_8 FILLER_75_815 ();
 sg13g2_decap_8 FILLER_75_822 ();
 sg13g2_decap_8 FILLER_75_829 ();
 sg13g2_decap_8 FILLER_75_836 ();
 sg13g2_decap_8 FILLER_75_843 ();
 sg13g2_decap_8 FILLER_75_850 ();
 sg13g2_decap_4 FILLER_75_857 ();
 sg13g2_fill_1 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_fill_2 FILLER_76_98 ();
 sg13g2_fill_1 FILLER_76_100 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_fill_2 FILLER_76_112 ();
 sg13g2_decap_4 FILLER_76_118 ();
 sg13g2_fill_2 FILLER_76_152 ();
 sg13g2_fill_1 FILLER_76_154 ();
 sg13g2_fill_1 FILLER_76_170 ();
 sg13g2_fill_2 FILLER_76_195 ();
 sg13g2_fill_1 FILLER_76_197 ();
 sg13g2_fill_1 FILLER_76_224 ();
 sg13g2_fill_1 FILLER_76_234 ();
 sg13g2_fill_2 FILLER_76_246 ();
 sg13g2_fill_2 FILLER_76_253 ();
 sg13g2_fill_1 FILLER_76_276 ();
 sg13g2_fill_1 FILLER_76_317 ();
 sg13g2_fill_2 FILLER_76_328 ();
 sg13g2_fill_1 FILLER_76_330 ();
 sg13g2_fill_2 FILLER_76_338 ();
 sg13g2_fill_1 FILLER_76_340 ();
 sg13g2_decap_4 FILLER_76_378 ();
 sg13g2_fill_2 FILLER_76_417 ();
 sg13g2_fill_1 FILLER_76_466 ();
 sg13g2_decap_8 FILLER_76_506 ();
 sg13g2_decap_8 FILLER_76_513 ();
 sg13g2_decap_8 FILLER_76_520 ();
 sg13g2_decap_8 FILLER_76_527 ();
 sg13g2_decap_8 FILLER_76_534 ();
 sg13g2_decap_8 FILLER_76_541 ();
 sg13g2_decap_8 FILLER_76_548 ();
 sg13g2_decap_8 FILLER_76_555 ();
 sg13g2_decap_8 FILLER_76_562 ();
 sg13g2_decap_8 FILLER_76_569 ();
 sg13g2_decap_8 FILLER_76_576 ();
 sg13g2_decap_8 FILLER_76_583 ();
 sg13g2_decap_8 FILLER_76_590 ();
 sg13g2_decap_8 FILLER_76_597 ();
 sg13g2_decap_8 FILLER_76_604 ();
 sg13g2_decap_8 FILLER_76_611 ();
 sg13g2_decap_8 FILLER_76_618 ();
 sg13g2_decap_8 FILLER_76_625 ();
 sg13g2_decap_8 FILLER_76_632 ();
 sg13g2_decap_8 FILLER_76_639 ();
 sg13g2_decap_8 FILLER_76_646 ();
 sg13g2_decap_8 FILLER_76_653 ();
 sg13g2_decap_8 FILLER_76_660 ();
 sg13g2_decap_8 FILLER_76_667 ();
 sg13g2_decap_8 FILLER_76_674 ();
 sg13g2_decap_8 FILLER_76_681 ();
 sg13g2_decap_8 FILLER_76_688 ();
 sg13g2_decap_8 FILLER_76_695 ();
 sg13g2_decap_8 FILLER_76_702 ();
 sg13g2_decap_8 FILLER_76_709 ();
 sg13g2_decap_8 FILLER_76_716 ();
 sg13g2_decap_8 FILLER_76_723 ();
 sg13g2_decap_8 FILLER_76_730 ();
 sg13g2_decap_8 FILLER_76_737 ();
 sg13g2_decap_8 FILLER_76_744 ();
 sg13g2_decap_8 FILLER_76_751 ();
 sg13g2_decap_8 FILLER_76_758 ();
 sg13g2_decap_8 FILLER_76_765 ();
 sg13g2_decap_8 FILLER_76_772 ();
 sg13g2_decap_8 FILLER_76_779 ();
 sg13g2_decap_8 FILLER_76_786 ();
 sg13g2_decap_8 FILLER_76_793 ();
 sg13g2_decap_8 FILLER_76_800 ();
 sg13g2_decap_8 FILLER_76_807 ();
 sg13g2_decap_8 FILLER_76_814 ();
 sg13g2_decap_8 FILLER_76_821 ();
 sg13g2_decap_8 FILLER_76_828 ();
 sg13g2_decap_8 FILLER_76_835 ();
 sg13g2_decap_8 FILLER_76_842 ();
 sg13g2_decap_8 FILLER_76_849 ();
 sg13g2_decap_4 FILLER_76_856 ();
 sg13g2_fill_2 FILLER_76_860 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_4 FILLER_77_98 ();
 sg13g2_fill_1 FILLER_77_102 ();
 sg13g2_fill_2 FILLER_77_165 ();
 sg13g2_fill_1 FILLER_77_167 ();
 sg13g2_fill_1 FILLER_77_178 ();
 sg13g2_fill_1 FILLER_77_184 ();
 sg13g2_fill_2 FILLER_77_195 ();
 sg13g2_fill_2 FILLER_77_206 ();
 sg13g2_decap_4 FILLER_77_258 ();
 sg13g2_fill_2 FILLER_77_272 ();
 sg13g2_fill_1 FILLER_77_274 ();
 sg13g2_fill_2 FILLER_77_301 ();
 sg13g2_fill_1 FILLER_77_303 ();
 sg13g2_fill_2 FILLER_77_313 ();
 sg13g2_fill_1 FILLER_77_315 ();
 sg13g2_fill_2 FILLER_77_333 ();
 sg13g2_fill_2 FILLER_77_346 ();
 sg13g2_fill_2 FILLER_77_386 ();
 sg13g2_fill_2 FILLER_77_438 ();
 sg13g2_decap_8 FILLER_77_498 ();
 sg13g2_decap_8 FILLER_77_505 ();
 sg13g2_decap_8 FILLER_77_512 ();
 sg13g2_decap_8 FILLER_77_519 ();
 sg13g2_decap_8 FILLER_77_526 ();
 sg13g2_decap_8 FILLER_77_533 ();
 sg13g2_decap_8 FILLER_77_540 ();
 sg13g2_decap_8 FILLER_77_547 ();
 sg13g2_decap_8 FILLER_77_554 ();
 sg13g2_decap_8 FILLER_77_561 ();
 sg13g2_decap_8 FILLER_77_568 ();
 sg13g2_decap_8 FILLER_77_575 ();
 sg13g2_decap_8 FILLER_77_582 ();
 sg13g2_decap_8 FILLER_77_589 ();
 sg13g2_decap_8 FILLER_77_596 ();
 sg13g2_decap_8 FILLER_77_603 ();
 sg13g2_decap_8 FILLER_77_610 ();
 sg13g2_decap_8 FILLER_77_617 ();
 sg13g2_decap_8 FILLER_77_624 ();
 sg13g2_decap_8 FILLER_77_631 ();
 sg13g2_decap_8 FILLER_77_638 ();
 sg13g2_decap_8 FILLER_77_645 ();
 sg13g2_decap_8 FILLER_77_652 ();
 sg13g2_decap_8 FILLER_77_659 ();
 sg13g2_decap_8 FILLER_77_666 ();
 sg13g2_decap_8 FILLER_77_673 ();
 sg13g2_decap_8 FILLER_77_680 ();
 sg13g2_decap_8 FILLER_77_687 ();
 sg13g2_decap_8 FILLER_77_694 ();
 sg13g2_decap_8 FILLER_77_701 ();
 sg13g2_decap_8 FILLER_77_708 ();
 sg13g2_decap_8 FILLER_77_715 ();
 sg13g2_decap_8 FILLER_77_722 ();
 sg13g2_decap_8 FILLER_77_729 ();
 sg13g2_decap_8 FILLER_77_736 ();
 sg13g2_decap_8 FILLER_77_743 ();
 sg13g2_decap_8 FILLER_77_750 ();
 sg13g2_decap_8 FILLER_77_757 ();
 sg13g2_decap_8 FILLER_77_764 ();
 sg13g2_decap_8 FILLER_77_771 ();
 sg13g2_decap_8 FILLER_77_778 ();
 sg13g2_decap_8 FILLER_77_785 ();
 sg13g2_decap_8 FILLER_77_792 ();
 sg13g2_decap_8 FILLER_77_799 ();
 sg13g2_decap_8 FILLER_77_806 ();
 sg13g2_decap_8 FILLER_77_813 ();
 sg13g2_decap_8 FILLER_77_820 ();
 sg13g2_decap_8 FILLER_77_827 ();
 sg13g2_decap_8 FILLER_77_834 ();
 sg13g2_decap_8 FILLER_77_841 ();
 sg13g2_decap_8 FILLER_77_848 ();
 sg13g2_decap_8 FILLER_77_855 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_fill_1 FILLER_78_167 ();
 sg13g2_fill_2 FILLER_78_229 ();
 sg13g2_fill_1 FILLER_78_296 ();
 sg13g2_decap_4 FILLER_78_381 ();
 sg13g2_fill_2 FILLER_78_428 ();
 sg13g2_fill_1 FILLER_78_430 ();
 sg13g2_fill_2 FILLER_78_458 ();
 sg13g2_fill_1 FILLER_78_460 ();
 sg13g2_fill_2 FILLER_78_475 ();
 sg13g2_decap_8 FILLER_78_490 ();
 sg13g2_decap_8 FILLER_78_497 ();
 sg13g2_decap_8 FILLER_78_504 ();
 sg13g2_decap_8 FILLER_78_511 ();
 sg13g2_decap_8 FILLER_78_518 ();
 sg13g2_decap_8 FILLER_78_525 ();
 sg13g2_decap_8 FILLER_78_532 ();
 sg13g2_decap_8 FILLER_78_539 ();
 sg13g2_decap_8 FILLER_78_546 ();
 sg13g2_decap_8 FILLER_78_553 ();
 sg13g2_decap_8 FILLER_78_560 ();
 sg13g2_decap_8 FILLER_78_567 ();
 sg13g2_decap_8 FILLER_78_574 ();
 sg13g2_decap_8 FILLER_78_581 ();
 sg13g2_decap_8 FILLER_78_588 ();
 sg13g2_decap_8 FILLER_78_595 ();
 sg13g2_decap_8 FILLER_78_602 ();
 sg13g2_decap_8 FILLER_78_609 ();
 sg13g2_decap_8 FILLER_78_616 ();
 sg13g2_decap_8 FILLER_78_623 ();
 sg13g2_decap_8 FILLER_78_630 ();
 sg13g2_decap_8 FILLER_78_637 ();
 sg13g2_decap_8 FILLER_78_644 ();
 sg13g2_decap_8 FILLER_78_651 ();
 sg13g2_decap_8 FILLER_78_658 ();
 sg13g2_decap_8 FILLER_78_665 ();
 sg13g2_decap_8 FILLER_78_672 ();
 sg13g2_decap_8 FILLER_78_679 ();
 sg13g2_decap_8 FILLER_78_686 ();
 sg13g2_decap_8 FILLER_78_693 ();
 sg13g2_decap_8 FILLER_78_700 ();
 sg13g2_decap_8 FILLER_78_707 ();
 sg13g2_decap_8 FILLER_78_714 ();
 sg13g2_decap_8 FILLER_78_721 ();
 sg13g2_decap_8 FILLER_78_728 ();
 sg13g2_decap_8 FILLER_78_735 ();
 sg13g2_decap_8 FILLER_78_742 ();
 sg13g2_decap_8 FILLER_78_749 ();
 sg13g2_decap_8 FILLER_78_756 ();
 sg13g2_decap_8 FILLER_78_763 ();
 sg13g2_decap_8 FILLER_78_770 ();
 sg13g2_decap_8 FILLER_78_777 ();
 sg13g2_decap_8 FILLER_78_784 ();
 sg13g2_decap_8 FILLER_78_791 ();
 sg13g2_decap_8 FILLER_78_798 ();
 sg13g2_decap_8 FILLER_78_805 ();
 sg13g2_decap_8 FILLER_78_812 ();
 sg13g2_decap_8 FILLER_78_819 ();
 sg13g2_decap_8 FILLER_78_826 ();
 sg13g2_decap_8 FILLER_78_833 ();
 sg13g2_decap_8 FILLER_78_840 ();
 sg13g2_decap_8 FILLER_78_847 ();
 sg13g2_decap_8 FILLER_78_854 ();
 sg13g2_fill_1 FILLER_78_861 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_4 FILLER_79_119 ();
 sg13g2_fill_2 FILLER_79_123 ();
 sg13g2_fill_1 FILLER_79_193 ();
 sg13g2_fill_1 FILLER_79_202 ();
 sg13g2_fill_2 FILLER_79_211 ();
 sg13g2_fill_1 FILLER_79_213 ();
 sg13g2_fill_1 FILLER_79_218 ();
 sg13g2_decap_8 FILLER_79_236 ();
 sg13g2_fill_2 FILLER_79_243 ();
 sg13g2_fill_1 FILLER_79_249 ();
 sg13g2_fill_1 FILLER_79_254 ();
 sg13g2_decap_4 FILLER_79_259 ();
 sg13g2_fill_1 FILLER_79_289 ();
 sg13g2_fill_2 FILLER_79_320 ();
 sg13g2_fill_1 FILLER_79_322 ();
 sg13g2_fill_1 FILLER_79_349 ();
 sg13g2_fill_1 FILLER_79_354 ();
 sg13g2_decap_8 FILLER_79_389 ();
 sg13g2_decap_4 FILLER_79_410 ();
 sg13g2_fill_1 FILLER_79_414 ();
 sg13g2_fill_2 FILLER_79_449 ();
 sg13g2_fill_1 FILLER_79_456 ();
 sg13g2_decap_8 FILLER_79_509 ();
 sg13g2_decap_8 FILLER_79_516 ();
 sg13g2_decap_8 FILLER_79_523 ();
 sg13g2_decap_8 FILLER_79_530 ();
 sg13g2_decap_8 FILLER_79_537 ();
 sg13g2_decap_8 FILLER_79_544 ();
 sg13g2_decap_8 FILLER_79_551 ();
 sg13g2_decap_8 FILLER_79_558 ();
 sg13g2_decap_8 FILLER_79_565 ();
 sg13g2_decap_8 FILLER_79_572 ();
 sg13g2_decap_8 FILLER_79_579 ();
 sg13g2_decap_8 FILLER_79_586 ();
 sg13g2_decap_8 FILLER_79_593 ();
 sg13g2_decap_8 FILLER_79_600 ();
 sg13g2_decap_8 FILLER_79_607 ();
 sg13g2_decap_8 FILLER_79_614 ();
 sg13g2_decap_8 FILLER_79_621 ();
 sg13g2_decap_8 FILLER_79_628 ();
 sg13g2_decap_8 FILLER_79_635 ();
 sg13g2_decap_8 FILLER_79_642 ();
 sg13g2_decap_8 FILLER_79_649 ();
 sg13g2_decap_8 FILLER_79_656 ();
 sg13g2_decap_8 FILLER_79_663 ();
 sg13g2_decap_8 FILLER_79_670 ();
 sg13g2_decap_8 FILLER_79_677 ();
 sg13g2_decap_8 FILLER_79_684 ();
 sg13g2_decap_8 FILLER_79_691 ();
 sg13g2_decap_8 FILLER_79_698 ();
 sg13g2_decap_8 FILLER_79_705 ();
 sg13g2_decap_8 FILLER_79_712 ();
 sg13g2_decap_8 FILLER_79_719 ();
 sg13g2_decap_8 FILLER_79_726 ();
 sg13g2_decap_8 FILLER_79_733 ();
 sg13g2_decap_8 FILLER_79_740 ();
 sg13g2_decap_8 FILLER_79_747 ();
 sg13g2_decap_8 FILLER_79_754 ();
 sg13g2_decap_8 FILLER_79_761 ();
 sg13g2_decap_8 FILLER_79_768 ();
 sg13g2_decap_8 FILLER_79_775 ();
 sg13g2_decap_8 FILLER_79_782 ();
 sg13g2_decap_8 FILLER_79_789 ();
 sg13g2_decap_8 FILLER_79_796 ();
 sg13g2_decap_8 FILLER_79_803 ();
 sg13g2_decap_8 FILLER_79_810 ();
 sg13g2_decap_8 FILLER_79_817 ();
 sg13g2_decap_8 FILLER_79_824 ();
 sg13g2_decap_8 FILLER_79_831 ();
 sg13g2_decap_8 FILLER_79_838 ();
 sg13g2_decap_8 FILLER_79_845 ();
 sg13g2_decap_8 FILLER_79_852 ();
 sg13g2_fill_2 FILLER_79_859 ();
 sg13g2_fill_1 FILLER_79_861 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_fill_2 FILLER_80_116 ();
 sg13g2_fill_2 FILLER_80_160 ();
 sg13g2_fill_1 FILLER_80_162 ();
 sg13g2_fill_2 FILLER_80_171 ();
 sg13g2_fill_2 FILLER_80_177 ();
 sg13g2_fill_1 FILLER_80_179 ();
 sg13g2_decap_4 FILLER_80_211 ();
 sg13g2_fill_2 FILLER_80_215 ();
 sg13g2_fill_1 FILLER_80_243 ();
 sg13g2_decap_4 FILLER_80_270 ();
 sg13g2_decap_8 FILLER_80_278 ();
 sg13g2_fill_1 FILLER_80_285 ();
 sg13g2_fill_2 FILLER_80_312 ();
 sg13g2_fill_2 FILLER_80_340 ();
 sg13g2_fill_1 FILLER_80_342 ();
 sg13g2_fill_2 FILLER_80_372 ();
 sg13g2_fill_2 FILLER_80_404 ();
 sg13g2_fill_1 FILLER_80_432 ();
 sg13g2_fill_2 FILLER_80_457 ();
 sg13g2_fill_2 FILLER_80_469 ();
 sg13g2_fill_1 FILLER_80_471 ();
 sg13g2_decap_8 FILLER_80_494 ();
 sg13g2_decap_8 FILLER_80_501 ();
 sg13g2_decap_8 FILLER_80_508 ();
 sg13g2_decap_8 FILLER_80_515 ();
 sg13g2_decap_8 FILLER_80_522 ();
 sg13g2_decap_8 FILLER_80_529 ();
 sg13g2_decap_8 FILLER_80_536 ();
 sg13g2_decap_8 FILLER_80_543 ();
 sg13g2_decap_8 FILLER_80_550 ();
 sg13g2_decap_8 FILLER_80_557 ();
 sg13g2_decap_8 FILLER_80_564 ();
 sg13g2_decap_8 FILLER_80_571 ();
 sg13g2_decap_8 FILLER_80_578 ();
 sg13g2_decap_8 FILLER_80_585 ();
 sg13g2_decap_8 FILLER_80_592 ();
 sg13g2_decap_8 FILLER_80_599 ();
 sg13g2_decap_8 FILLER_80_606 ();
 sg13g2_decap_8 FILLER_80_613 ();
 sg13g2_decap_8 FILLER_80_620 ();
 sg13g2_decap_8 FILLER_80_627 ();
 sg13g2_decap_8 FILLER_80_634 ();
 sg13g2_decap_8 FILLER_80_641 ();
 sg13g2_decap_8 FILLER_80_648 ();
 sg13g2_decap_8 FILLER_80_655 ();
 sg13g2_decap_8 FILLER_80_662 ();
 sg13g2_decap_8 FILLER_80_669 ();
 sg13g2_decap_8 FILLER_80_676 ();
 sg13g2_decap_8 FILLER_80_683 ();
 sg13g2_decap_8 FILLER_80_690 ();
 sg13g2_decap_8 FILLER_80_697 ();
 sg13g2_decap_8 FILLER_80_704 ();
 sg13g2_decap_8 FILLER_80_711 ();
 sg13g2_decap_8 FILLER_80_718 ();
 sg13g2_decap_8 FILLER_80_725 ();
 sg13g2_decap_8 FILLER_80_732 ();
 sg13g2_decap_8 FILLER_80_739 ();
 sg13g2_decap_8 FILLER_80_746 ();
 sg13g2_decap_8 FILLER_80_753 ();
 sg13g2_decap_8 FILLER_80_760 ();
 sg13g2_decap_8 FILLER_80_767 ();
 sg13g2_decap_8 FILLER_80_774 ();
 sg13g2_decap_8 FILLER_80_781 ();
 sg13g2_decap_8 FILLER_80_788 ();
 sg13g2_decap_8 FILLER_80_795 ();
 sg13g2_decap_8 FILLER_80_802 ();
 sg13g2_decap_8 FILLER_80_809 ();
 sg13g2_decap_8 FILLER_80_816 ();
 sg13g2_decap_8 FILLER_80_823 ();
 sg13g2_decap_8 FILLER_80_830 ();
 sg13g2_decap_8 FILLER_80_837 ();
 sg13g2_decap_8 FILLER_80_844 ();
 sg13g2_decap_8 FILLER_80_851 ();
 sg13g2_decap_4 FILLER_80_858 ();
 assign uio_oe[0] = net5;
 assign uio_oe[1] = net6;
 assign uio_oe[2] = net7;
 assign uio_oe[3] = net8;
 assign uio_oe[4] = net9;
 assign uio_oe[5] = net10;
 assign uio_oe[6] = net11;
 assign uio_oe[7] = net12;
 assign uio_out[0] = net13;
 assign uio_out[1] = net14;
 assign uio_out[2] = net15;
 assign uio_out[3] = net16;
 assign uio_out[4] = net17;
 assign uio_out[5] = net18;
 assign uio_out[6] = net19;
 assign uio_out[7] = net20;
endmodule

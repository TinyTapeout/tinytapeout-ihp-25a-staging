module tt_um_adder_accumulator_sathworld (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire CF;
 wire ZF;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire clknet_0_clk;
 wire net61;
 wire net60;
 wire net59;
 wire net58;
 wire net57;
 wire net56;
 wire net55;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net28;
 wire net29;
 wire net30;
 wire \accumulatorobj.bus[0] ;
 wire \accumulatorobj.bus[1] ;
 wire \accumulatorobj.bus[2] ;
 wire \accumulatorobj.bus[3] ;
 wire \accumulatorobj.bus[4] ;
 wire \accumulatorobj.bus[5] ;
 wire \accumulatorobj.bus[6] ;
 wire \accumulatorobj.bus[7] ;
 wire \aluobj.addsub.genblk1[0].fa.a ;
 wire \aluobj.addsub.genblk1[0].fa.sum ;
 wire \aluobj.addsub.genblk1[1].fa.a ;
 wire \aluobj.addsub.genblk1[1].fa.sum ;
 wire \aluobj.addsub.genblk1[2].fa.a ;
 wire \aluobj.addsub.genblk1[2].fa.sum ;
 wire \aluobj.addsub.genblk1[3].fa.a ;
 wire \aluobj.addsub.genblk1[3].fa.sum ;
 wire \aluobj.addsub.genblk1[4].fa.a ;
 wire \aluobj.addsub.genblk1[4].fa.sum ;
 wire \aluobj.addsub.genblk1[5].fa.a ;
 wire \aluobj.addsub.genblk1[5].fa.sum ;
 wire \aluobj.addsub.genblk1[6].fa.a ;
 wire \aluobj.addsub.genblk1[6].fa.sum ;
 wire \aluobj.addsub.genblk1[7].fa.a ;
 wire \aluobj.addsub.genblk1[7].fa.sum ;
 wire \aluobj.addsub.op_b[0] ;
 wire \aluobj.addsub.op_b[1] ;
 wire \aluobj.addsub.op_b[2] ;
 wire \aluobj.addsub.op_b[3] ;
 wire \aluobj.addsub.op_b[4] ;
 wire \aluobj.addsub.op_b[5] ;
 wire \aluobj.addsub.op_b[6] ;
 wire \aluobj.addsub.op_b[7] ;
 wire \ui_in_buf[0] ;
 wire \ui_in_buf[1] ;
 wire \ui_in_buf[2] ;
 wire \ui_in_buf[3] ;
 wire \ui_in_buf[4] ;
 wire \ui_in_buf[5] ;
 wire \ui_in_buf[6] ;
 wire \ui_in_buf[7] ;
 wire net53;
 wire net54;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;

 sg13g2_inv_2 _144_ (.Y(_085_),
    .A(net11));
 sg13g2_nand2_2 _145_ (.Y(_077_),
    .A(net23),
    .B(net25));
 sg13g2_inv_1 _146_ (.Y(_027_),
    .A(_077_));
 sg13g2_nor2_1 _147_ (.A(net24),
    .B(net10),
    .Y(_028_));
 sg13g2_inv_1 _148_ (.Y(_070_),
    .A(_028_));
 sg13g2_xor2_1 _149_ (.B(\aluobj.addsub.genblk1[0].fa.a ),
    .A(\aluobj.addsub.op_b[0] ),
    .X(\aluobj.addsub.genblk1[0].fa.sum ));
 sg13g2_mux2_1 _150_ (.A0(net9),
    .A1(\aluobj.addsub.genblk1[0].fa.a ),
    .S(\aluobj.addsub.op_b[0] ),
    .X(_029_));
 sg13g2_xnor2_1 _151_ (.Y(_030_),
    .A(\aluobj.addsub.op_b[1] ),
    .B(net9));
 sg13g2_nand2_1 _152_ (.Y(_031_),
    .A(_000_),
    .B(_030_));
 sg13g2_nor2_1 _153_ (.A(_000_),
    .B(_030_),
    .Y(_032_));
 sg13g2_xnor2_1 _154_ (.Y(_033_),
    .A(_000_),
    .B(_030_));
 sg13g2_xnor2_1 _155_ (.Y(\aluobj.addsub.genblk1[1].fa.sum ),
    .A(_029_),
    .B(_033_));
 sg13g2_xor2_1 _156_ (.B(\aluobj.addsub.op_b[2] ),
    .A(net9),
    .X(_034_));
 sg13g2_and2_1 _157_ (.A(\aluobj.addsub.genblk1[2].fa.a ),
    .B(_034_),
    .X(_035_));
 sg13g2_or2_1 _158_ (.X(_036_),
    .B(_034_),
    .A(\aluobj.addsub.genblk1[2].fa.a ));
 sg13g2_nand2b_1 _159_ (.Y(_037_),
    .B(_036_),
    .A_N(_035_));
 sg13g2_a21o_1 _160_ (.A2(_031_),
    .A1(_029_),
    .B1(_032_),
    .X(_038_));
 sg13g2_xnor2_1 _161_ (.Y(\aluobj.addsub.genblk1[2].fa.sum ),
    .A(_037_),
    .B(_038_));
 sg13g2_xor2_1 _162_ (.B(\aluobj.addsub.op_b[3] ),
    .A(net9),
    .X(_039_));
 sg13g2_nand2_1 _163_ (.Y(_040_),
    .A(\aluobj.addsub.genblk1[3].fa.a ),
    .B(_039_));
 sg13g2_nor2_1 _164_ (.A(\aluobj.addsub.genblk1[3].fa.a ),
    .B(_039_),
    .Y(_041_));
 sg13g2_xor2_1 _165_ (.B(_039_),
    .A(\aluobj.addsub.genblk1[3].fa.a ),
    .X(_042_));
 sg13g2_a21oi_1 _166_ (.A1(_036_),
    .A2(_038_),
    .Y(_043_),
    .B1(_035_));
 sg13g2_xnor2_1 _167_ (.Y(\aluobj.addsub.genblk1[3].fa.sum ),
    .A(_042_),
    .B(_043_));
 sg13g2_xor2_1 _168_ (.B(\aluobj.addsub.op_b[4] ),
    .A(net9),
    .X(_044_));
 sg13g2_and2_1 _169_ (.A(\aluobj.addsub.genblk1[4].fa.a ),
    .B(_044_),
    .X(_045_));
 sg13g2_or2_1 _170_ (.X(_046_),
    .B(_044_),
    .A(\aluobj.addsub.genblk1[4].fa.a ));
 sg13g2_nand2b_1 _171_ (.Y(_047_),
    .B(_046_),
    .A_N(_045_));
 sg13g2_o21ai_1 _172_ (.B1(_040_),
    .Y(_048_),
    .A1(_041_),
    .A2(_043_));
 sg13g2_xnor2_1 _173_ (.Y(\aluobj.addsub.genblk1[4].fa.sum ),
    .A(_047_),
    .B(_048_));
 sg13g2_xor2_1 _174_ (.B(\aluobj.addsub.op_b[5] ),
    .A(net9),
    .X(_049_));
 sg13g2_nand2_1 _175_ (.Y(_050_),
    .A(\aluobj.addsub.genblk1[5].fa.a ),
    .B(_049_));
 sg13g2_nor2_1 _176_ (.A(\aluobj.addsub.genblk1[5].fa.a ),
    .B(_049_),
    .Y(_051_));
 sg13g2_xnor2_1 _177_ (.Y(_052_),
    .A(\aluobj.addsub.genblk1[5].fa.a ),
    .B(_049_));
 sg13g2_a21oi_1 _178_ (.A1(_046_),
    .A2(_048_),
    .Y(_053_),
    .B1(_045_));
 sg13g2_xor2_1 _179_ (.B(_053_),
    .A(_052_),
    .X(\aluobj.addsub.genblk1[5].fa.sum ));
 sg13g2_xor2_1 _180_ (.B(\aluobj.addsub.op_b[6] ),
    .A(net9),
    .X(_054_));
 sg13g2_and2_1 _181_ (.A(\aluobj.addsub.genblk1[6].fa.a ),
    .B(_054_),
    .X(_055_));
 sg13g2_or2_1 _182_ (.X(_056_),
    .B(_054_),
    .A(\aluobj.addsub.genblk1[6].fa.a ));
 sg13g2_nand2b_1 _183_ (.Y(_057_),
    .B(_056_),
    .A_N(_055_));
 sg13g2_o21ai_1 _184_ (.B1(_050_),
    .Y(_058_),
    .A1(_051_),
    .A2(_053_));
 sg13g2_xnor2_1 _185_ (.Y(\aluobj.addsub.genblk1[6].fa.sum ),
    .A(_057_),
    .B(_058_));
 sg13g2_xor2_1 _186_ (.B(\aluobj.addsub.op_b[7] ),
    .A(net9),
    .X(_059_));
 sg13g2_nand2_1 _187_ (.Y(_060_),
    .A(\aluobj.addsub.genblk1[7].fa.a ),
    .B(_059_));
 sg13g2_xor2_1 _188_ (.B(_059_),
    .A(\aluobj.addsub.genblk1[7].fa.a ),
    .X(_061_));
 sg13g2_a21oi_1 _189_ (.A1(_056_),
    .A2(_058_),
    .Y(_062_),
    .B1(_055_));
 sg13g2_xnor2_1 _190_ (.Y(\aluobj.addsub.genblk1[7].fa.sum ),
    .A(_061_),
    .B(_062_));
 sg13g2_mux2_1 _191_ (.A0(\aluobj.addsub.genblk1[0].fa.a ),
    .A1(\accumulatorobj.bus[0] ),
    .S(net14),
    .X(uo_out[0]));
 sg13g2_mux2_1 _192_ (.A0(\aluobj.addsub.genblk1[1].fa.a ),
    .A1(\accumulatorobj.bus[1] ),
    .S(net14),
    .X(uo_out[1]));
 sg13g2_mux2_2 _193_ (.A0(\aluobj.addsub.genblk1[2].fa.a ),
    .A1(\accumulatorobj.bus[2] ),
    .S(net14),
    .X(uo_out[2]));
 sg13g2_mux2_2 _194_ (.A0(\aluobj.addsub.genblk1[3].fa.a ),
    .A1(\accumulatorobj.bus[3] ),
    .S(net14),
    .X(uo_out[3]));
 sg13g2_mux2_1 _195_ (.A0(\aluobj.addsub.genblk1[4].fa.a ),
    .A1(\accumulatorobj.bus[4] ),
    .S(net14),
    .X(uo_out[4]));
 sg13g2_mux2_1 _196_ (.A0(\aluobj.addsub.genblk1[5].fa.a ),
    .A1(\accumulatorobj.bus[5] ),
    .S(net14),
    .X(uo_out[5]));
 sg13g2_mux2_1 _197_ (.A0(\aluobj.addsub.genblk1[6].fa.a ),
    .A1(\accumulatorobj.bus[6] ),
    .S(net14),
    .X(uo_out[6]));
 sg13g2_mux2_1 _198_ (.A0(\aluobj.addsub.genblk1[7].fa.a ),
    .A1(\accumulatorobj.bus[7] ),
    .S(net14),
    .X(uo_out[7]));
 sg13g2_and2_1 _199_ (.A(net1),
    .B(net21),
    .X(_001_));
 sg13g2_and2_1 _200_ (.A(net2),
    .B(net21),
    .X(_002_));
 sg13g2_and2_1 _201_ (.A(net3),
    .B(net21),
    .X(_003_));
 sg13g2_and2_1 _202_ (.A(net4),
    .B(net21),
    .X(_004_));
 sg13g2_and2_1 _203_ (.A(net5),
    .B(net22),
    .X(_005_));
 sg13g2_and2_1 _204_ (.A(net6),
    .B(net22),
    .X(_006_));
 sg13g2_and2_1 _205_ (.A(net7),
    .B(net22),
    .X(_007_));
 sg13g2_and2_1 _206_ (.A(net8),
    .B(net22),
    .X(_008_));
 sg13g2_mux2_1 _207_ (.A0(\accumulatorobj.bus[0] ),
    .A1(net81),
    .S(net12),
    .X(_009_));
 sg13g2_mux2_1 _208_ (.A0(\accumulatorobj.bus[1] ),
    .A1(net77),
    .S(net12),
    .X(_010_));
 sg13g2_mux2_1 _209_ (.A0(\accumulatorobj.bus[2] ),
    .A1(net65),
    .S(net12),
    .X(_011_));
 sg13g2_mux2_1 _210_ (.A0(\accumulatorobj.bus[3] ),
    .A1(net75),
    .S(net12),
    .X(_012_));
 sg13g2_mux2_1 _211_ (.A0(\accumulatorobj.bus[4] ),
    .A1(net67),
    .S(net12),
    .X(_013_));
 sg13g2_mux2_1 _212_ (.A0(\accumulatorobj.bus[5] ),
    .A1(net69),
    .S(net12),
    .X(_014_));
 sg13g2_mux2_1 _213_ (.A0(\accumulatorobj.bus[6] ),
    .A1(net73),
    .S(net12),
    .X(_015_));
 sg13g2_mux2_1 _214_ (.A0(\accumulatorobj.bus[7] ),
    .A1(net71),
    .S(net12),
    .X(_016_));
 sg13g2_o21ai_1 _215_ (.B1(_027_),
    .Y(_063_),
    .A1(\aluobj.addsub.genblk1[7].fa.a ),
    .A2(_059_));
 sg13g2_a21oi_1 _216_ (.A1(_060_),
    .A2(_062_),
    .Y(_064_),
    .B1(_063_));
 sg13g2_a21o_1 _217_ (.A2(_077_),
    .A1(net63),
    .B1(_064_),
    .X(_017_));
 sg13g2_mux2_1 _218_ (.A0(\accumulatorobj.bus[0] ),
    .A1(net89),
    .S(net13),
    .X(_018_));
 sg13g2_mux2_1 _219_ (.A0(\accumulatorobj.bus[1] ),
    .A1(net79),
    .S(net13),
    .X(_019_));
 sg13g2_mux2_1 _220_ (.A0(\accumulatorobj.bus[2] ),
    .A1(net87),
    .S(net13),
    .X(_020_));
 sg13g2_mux2_1 _221_ (.A0(\accumulatorobj.bus[3] ),
    .A1(net91),
    .S(net13),
    .X(_021_));
 sg13g2_mux2_1 _222_ (.A0(\accumulatorobj.bus[4] ),
    .A1(net83),
    .S(net13),
    .X(_022_));
 sg13g2_mux2_1 _223_ (.A0(\accumulatorobj.bus[5] ),
    .A1(net95),
    .S(net13),
    .X(_023_));
 sg13g2_mux2_1 _224_ (.A0(\accumulatorobj.bus[6] ),
    .A1(net85),
    .S(net13),
    .X(_024_));
 sg13g2_mux2_1 _225_ (.A0(\accumulatorobj.bus[7] ),
    .A1(net93),
    .S(net13),
    .X(_025_));
 sg13g2_nand2_1 _226_ (.Y(_065_),
    .A(net62),
    .B(_077_));
 sg13g2_nor4_1 _227_ (.A(\aluobj.addsub.genblk1[1].fa.sum ),
    .B(\aluobj.addsub.genblk1[2].fa.sum ),
    .C(\aluobj.addsub.genblk1[3].fa.sum ),
    .D(\aluobj.addsub.genblk1[4].fa.sum ),
    .Y(_066_));
 sg13g2_nand2b_1 _228_ (.Y(_067_),
    .B(_066_),
    .A_N(\aluobj.addsub.genblk1[5].fa.sum ));
 sg13g2_or4_1 _229_ (.A(_077_),
    .B(\aluobj.addsub.genblk1[0].fa.sum ),
    .C(\aluobj.addsub.genblk1[6].fa.sum ),
    .D(_067_),
    .X(_068_));
 sg13g2_o21ai_1 _230_ (.B1(_065_),
    .Y(_026_),
    .A1(\aluobj.addsub.genblk1[7].fa.sum ),
    .A2(_068_));
 sg13g2_nand2_2 _231_ (.Y(_078_),
    .A(net23),
    .B(net25));
 sg13g2_nand2_2 _232_ (.Y(_079_),
    .A(net23),
    .B(net25));
 sg13g2_nand2_2 _233_ (.Y(_080_),
    .A(net23),
    .B(net25));
 sg13g2_nand2_2 _234_ (.Y(_081_),
    .A(net23),
    .B(net25));
 sg13g2_nand2_2 _235_ (.Y(_082_),
    .A(net23),
    .B(net25));
 sg13g2_nand2_2 _236_ (.Y(_083_),
    .A(net23),
    .B(net25));
 sg13g2_nand2_2 _237_ (.Y(_084_),
    .A(net23),
    .B(net25));
 sg13g2_inv_1 _238_ (.Y(_086_),
    .A(net24));
 sg13g2_inv_1 _239_ (.Y(_087_),
    .A(net24));
 sg13g2_inv_1 _240_ (.Y(_088_),
    .A(net24));
 sg13g2_inv_1 _241_ (.Y(_089_),
    .A(net24));
 sg13g2_inv_1 _242_ (.Y(_090_),
    .A(net24));
 sg13g2_inv_1 _243_ (.Y(_091_),
    .A(net24));
 sg13g2_inv_1 _244_ (.Y(_092_),
    .A(net24));
 sg13g2_inv_1 _245_ (.Y(_071_),
    .A(net21));
 sg13g2_inv_1 _246_ (.Y(_072_),
    .A(net21));
 sg13g2_inv_1 _247_ (.Y(_075_),
    .A(net22));
 sg13g2_inv_1 _248_ (.Y(_076_),
    .A(net22));
 sg13g2_inv_1 _249_ (.Y(_069_),
    .A(net21));
 sg13g2_inv_1 _250_ (.Y(_073_),
    .A(net21));
 sg13g2_inv_1 _251_ (.Y(_074_),
    .A(net22));
 sg13g2_dfrbp_1 _252_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net50),
    .D(_001_),
    .Q_N(_125_),
    .Q(\ui_in_buf[0] ));
 sg13g2_dfrbp_1 _253_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net49),
    .D(_002_),
    .Q_N(_124_),
    .Q(\ui_in_buf[1] ));
 sg13g2_dfrbp_1 _254_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net48),
    .D(_003_),
    .Q_N(_123_),
    .Q(\ui_in_buf[2] ));
 sg13g2_dfrbp_1 _255_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net47),
    .D(_004_),
    .Q_N(_122_),
    .Q(\ui_in_buf[3] ));
 sg13g2_dfrbp_1 _256_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net46),
    .D(_005_),
    .Q_N(_121_),
    .Q(\ui_in_buf[4] ));
 sg13g2_dfrbp_1 _257_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net45),
    .D(_006_),
    .Q_N(_120_),
    .Q(\ui_in_buf[5] ));
 sg13g2_dfrbp_1 _258_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net44),
    .D(_007_),
    .Q_N(_119_),
    .Q(\ui_in_buf[6] ));
 sg13g2_dfrbp_1 _259_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net43),
    .D(_008_),
    .Q_N(_118_),
    .Q(\ui_in_buf[7] ));
 sg13g2_dfrbp_1 _260_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net27),
    .D(net82),
    .Q_N(_117_),
    .Q(\aluobj.addsub.op_b[0] ));
 sg13g2_dfrbp_1 _261_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net27),
    .D(net78),
    .Q_N(_116_),
    .Q(\aluobj.addsub.op_b[1] ));
 sg13g2_dfrbp_1 _262_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net27),
    .D(net66),
    .Q_N(_115_),
    .Q(\aluobj.addsub.op_b[2] ));
 sg13g2_dfrbp_1 _263_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net27),
    .D(net76),
    .Q_N(_114_),
    .Q(\aluobj.addsub.op_b[3] ));
 sg13g2_dfrbp_1 _264_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net26),
    .D(net68),
    .Q_N(_113_),
    .Q(\aluobj.addsub.op_b[4] ));
 sg13g2_dfrbp_1 _265_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net26),
    .D(net70),
    .Q_N(_112_),
    .Q(\aluobj.addsub.op_b[5] ));
 sg13g2_dfrbp_1 _266_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net26),
    .D(net74),
    .Q_N(_111_),
    .Q(\aluobj.addsub.op_b[6] ));
 sg13g2_dfrbp_1 _267_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net26),
    .D(net72),
    .Q_N(_110_),
    .Q(\aluobj.addsub.op_b[7] ));
 sg13g2_dfrbp_1 _268_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net42),
    .D(net64),
    .Q_N(_109_),
    .Q(CF));
 sg13g2_dfrbp_1 _269_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net27),
    .D(net90),
    .Q_N(_108_),
    .Q(\aluobj.addsub.genblk1[0].fa.a ));
 sg13g2_dfrbp_1 _270_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net27),
    .D(net80),
    .Q_N(_000_),
    .Q(\aluobj.addsub.genblk1[1].fa.a ));
 sg13g2_dfrbp_1 _271_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net27),
    .D(net88),
    .Q_N(_107_),
    .Q(\aluobj.addsub.genblk1[2].fa.a ));
 sg13g2_dfrbp_1 _272_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net27),
    .D(net92),
    .Q_N(_106_),
    .Q(\aluobj.addsub.genblk1[3].fa.a ));
 sg13g2_dfrbp_1 _273_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net26),
    .D(net84),
    .Q_N(_105_),
    .Q(\aluobj.addsub.genblk1[4].fa.a ));
 sg13g2_dfrbp_1 _274_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net26),
    .D(net96),
    .Q_N(_104_),
    .Q(\aluobj.addsub.genblk1[5].fa.a ));
 sg13g2_dfrbp_1 _275_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net26),
    .D(net86),
    .Q_N(_103_),
    .Q(\aluobj.addsub.genblk1[6].fa.a ));
 sg13g2_dfrbp_1 _276_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net26),
    .D(net94),
    .Q_N(_102_),
    .Q(\aluobj.addsub.genblk1[7].fa.a ));
 sg13g2_dfrbp_1 _277_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net51),
    .D(_026_),
    .Q_N(_101_),
    .Q(ZF));
 sg13g2_tiehi _259__36 (.L_HI(net43));
 sg13g2_tiehi _258__37 (.L_HI(net44));
 sg13g2_tiehi _257__38 (.L_HI(net45));
 sg13g2_tiehi _256__39 (.L_HI(net46));
 sg13g2_tiehi _255__40 (.L_HI(net47));
 sg13g2_tiehi _254__41 (.L_HI(net48));
 sg13g2_tiehi _253__42 (.L_HI(net49));
 sg13g2_tiehi _252__43 (.L_HI(net50));
 sg13g2_tiehi _277__44 (.L_HI(net51));
 sg13g2_tiehi tt_um_adder_accumulator_sathworld_45 (.L_HI(net52));
 sg13g2_tiehi tt_um_adder_accumulator_sathworld_46 (.L_HI(net53));
 sg13g2_tiehi _351__47 (.L_HI(net54));
 sg13g2_tiehi _350__48 (.L_HI(net55));
 sg13g2_tiehi _349__49 (.L_HI(net56));
 sg13g2_tiehi _348__50 (.L_HI(net57));
 sg13g2_tiehi _347__51 (.L_HI(net58));
 sg13g2_tiehi _346__52 (.L_HI(net59));
 sg13g2_tiehi _345__53 (.L_HI(net60));
 sg13g2_tiehi _344__54 (.L_HI(net61));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo _345__16 (.L_LO(net16));
 sg13g2_tielo _346__17 (.L_LO(net17));
 sg13g2_tielo _347__18 (.L_LO(net18));
 sg13g2_tielo _348__19 (.L_LO(net19));
 sg13g2_tielo _349__20 (.L_LO(net20));
 sg13g2_tielo _350__21 (.L_LO(net28));
 sg13g2_tielo _351__22 (.L_LO(net29));
 sg13g2_tielo tt_um_adder_accumulator_sathworld_23 (.L_LO(net30));
 sg13g2_tielo tt_um_adder_accumulator_sathworld_24 (.L_LO(net31));
 sg13g2_tielo tt_um_adder_accumulator_sathworld_25 (.L_LO(net32));
 sg13g2_tielo tt_um_adder_accumulator_sathworld_26 (.L_LO(net33));
 sg13g2_tielo tt_um_adder_accumulator_sathworld_27 (.L_LO(net34));
 sg13g2_tielo tt_um_adder_accumulator_sathworld_28 (.L_LO(net35));
 sg13g2_tielo tt_um_adder_accumulator_sathworld_29 (.L_LO(net36));
 sg13g2_tielo tt_um_adder_accumulator_sathworld_30 (.L_LO(net37));
 sg13g2_tielo tt_um_adder_accumulator_sathworld_31 (.L_LO(net38));
 sg13g2_tielo tt_um_adder_accumulator_sathworld_32 (.L_LO(net39));
 sg13g2_tielo tt_um_adder_accumulator_sathworld_33 (.L_LO(net40));
 sg13g2_tielo tt_um_adder_accumulator_sathworld_34 (.L_LO(net41));
 sg13g2_tiehi _268__35 (.L_HI(net42));
 sg13g2_buf_1 _318_ (.A(ZF),
    .X(uio_out[0]));
 sg13g2_buf_1 _319_ (.A(CF),
    .X(uio_out[1]));
 sg13g2_ebufn_8 _320_ (.Z(\accumulatorobj.bus[0] ),
    .A(\ui_in_buf[0] ),
    .TE_B(_069_));
 sg13g2_ebufn_8 _321_ (.Z(\accumulatorobj.bus[1] ),
    .A(\ui_in_buf[1] ),
    .TE_B(_070_));
 sg13g2_ebufn_8 _322_ (.Z(\accumulatorobj.bus[2] ),
    .A(\ui_in_buf[2] ),
    .TE_B(_071_));
 sg13g2_ebufn_8 _323_ (.Z(\accumulatorobj.bus[3] ),
    .A(\ui_in_buf[3] ),
    .TE_B(_072_));
 sg13g2_ebufn_8 _324_ (.Z(\accumulatorobj.bus[4] ),
    .A(\ui_in_buf[4] ),
    .TE_B(_073_));
 sg13g2_ebufn_8 _325_ (.Z(\accumulatorobj.bus[5] ),
    .A(\ui_in_buf[5] ),
    .TE_B(_074_));
 sg13g2_ebufn_8 _326_ (.Z(\accumulatorobj.bus[6] ),
    .A(\ui_in_buf[6] ),
    .TE_B(_075_));
 sg13g2_ebufn_8 _327_ (.Z(\accumulatorobj.bus[7] ),
    .A(\ui_in_buf[7] ),
    .TE_B(_076_));
 sg13g2_ebufn_8 _328_ (.Z(\accumulatorobj.bus[0] ),
    .A(\aluobj.addsub.genblk1[0].fa.sum ),
    .TE_B(_077_));
 sg13g2_ebufn_8 _329_ (.Z(\accumulatorobj.bus[1] ),
    .A(\aluobj.addsub.genblk1[1].fa.sum ),
    .TE_B(_078_));
 sg13g2_ebufn_8 _330_ (.Z(\accumulatorobj.bus[2] ),
    .A(\aluobj.addsub.genblk1[2].fa.sum ),
    .TE_B(_079_));
 sg13g2_ebufn_8 _331_ (.Z(\accumulatorobj.bus[3] ),
    .A(\aluobj.addsub.genblk1[3].fa.sum ),
    .TE_B(_080_));
 sg13g2_ebufn_8 _332_ (.Z(\accumulatorobj.bus[4] ),
    .A(\aluobj.addsub.genblk1[4].fa.sum ),
    .TE_B(_081_));
 sg13g2_ebufn_8 _333_ (.Z(\accumulatorobj.bus[5] ),
    .A(\aluobj.addsub.genblk1[5].fa.sum ),
    .TE_B(_082_));
 sg13g2_ebufn_8 _334_ (.Z(\accumulatorobj.bus[6] ),
    .A(\aluobj.addsub.genblk1[6].fa.sum ),
    .TE_B(_083_));
 sg13g2_ebufn_8 _335_ (.Z(\accumulatorobj.bus[7] ),
    .A(\aluobj.addsub.genblk1[7].fa.sum ),
    .TE_B(_084_));
 sg13g2_ebufn_8 _336_ (.Z(\accumulatorobj.bus[0] ),
    .A(\aluobj.addsub.genblk1[0].fa.a ),
    .TE_B(_085_));
 sg13g2_ebufn_8 _337_ (.Z(\accumulatorobj.bus[1] ),
    .A(net79),
    .TE_B(_086_));
 sg13g2_ebufn_8 _338_ (.Z(\accumulatorobj.bus[2] ),
    .A(\aluobj.addsub.genblk1[2].fa.a ),
    .TE_B(_087_));
 sg13g2_ebufn_8 _339_ (.Z(\accumulatorobj.bus[3] ),
    .A(\aluobj.addsub.genblk1[3].fa.a ),
    .TE_B(_088_));
 sg13g2_ebufn_8 _340_ (.Z(\accumulatorobj.bus[4] ),
    .A(\aluobj.addsub.genblk1[4].fa.a ),
    .TE_B(_089_));
 sg13g2_ebufn_8 _341_ (.Z(\accumulatorobj.bus[5] ),
    .A(\aluobj.addsub.genblk1[5].fa.a ),
    .TE_B(_090_));
 sg13g2_ebufn_8 _342_ (.Z(\accumulatorobj.bus[6] ),
    .A(\aluobj.addsub.genblk1[6].fa.a ),
    .TE_B(_091_));
 sg13g2_ebufn_8 _343_ (.Z(\accumulatorobj.bus[7] ),
    .A(\aluobj.addsub.genblk1[7].fa.a ),
    .TE_B(_092_));
 sg13g2_ebufn_8 _344_ (.Z(\accumulatorobj.bus[0] ),
    .A(net15),
    .TE_B(net61));
 sg13g2_ebufn_8 _345_ (.Z(\accumulatorobj.bus[1] ),
    .A(net16),
    .TE_B(net60));
 sg13g2_ebufn_8 _346_ (.Z(\accumulatorobj.bus[2] ),
    .A(net17),
    .TE_B(net59));
 sg13g2_ebufn_8 _347_ (.Z(\accumulatorobj.bus[3] ),
    .A(net18),
    .TE_B(net58));
 sg13g2_ebufn_8 _348_ (.Z(\accumulatorobj.bus[4] ),
    .A(net19),
    .TE_B(net57));
 sg13g2_ebufn_8 _349_ (.Z(\accumulatorobj.bus[5] ),
    .A(net20),
    .TE_B(net56));
 sg13g2_ebufn_8 _350_ (.Z(\accumulatorobj.bus[6] ),
    .A(net28),
    .TE_B(net55));
 sg13g2_ebufn_8 _351_ (.Z(\accumulatorobj.bus[7] ),
    .A(net29),
    .TE_B(net54));
 sg13g2_buf_2 fanout21 (.A(net22),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_028_),
    .X(net22));
 sg13g2_buf_4 fanout23 (.X(net23),
    .A(_085_));
 sg13g2_buf_4 fanout24 (.X(net24),
    .A(net11));
 sg13g2_buf_4 fanout25 (.X(net25),
    .A(net10));
 sg13g2_buf_4 fanout26 (.X(net26),
    .A(rst_n));
 sg13g2_buf_4 fanout27 (.X(net27),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_4 input9 (.X(net9),
    .A(uio_in[2]));
 sg13g2_buf_1 input10 (.A(uio_in[3]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[4]),
    .X(net11));
 sg13g2_buf_4 input12 (.X(net12),
    .A(uio_in[5]));
 sg13g2_buf_4 input13 (.X(net13),
    .A(uio_in[6]));
 sg13g2_buf_4 input14 (.X(net14),
    .A(uio_in[7]));
 sg13g2_tielo _344__15 (.L_LO(net15));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(ZF),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold2 (.A(CF),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold3 (.A(_017_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold4 (.A(\aluobj.addsub.op_b[2] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold5 (.A(_011_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold6 (.A(\aluobj.addsub.op_b[4] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold7 (.A(_013_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold8 (.A(\aluobj.addsub.op_b[5] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold9 (.A(_014_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold10 (.A(\aluobj.addsub.op_b[7] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold11 (.A(_016_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold12 (.A(\aluobj.addsub.op_b[6] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold13 (.A(_015_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold14 (.A(\aluobj.addsub.op_b[3] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold15 (.A(_012_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold16 (.A(\aluobj.addsub.op_b[1] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold17 (.A(_010_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold18 (.A(\aluobj.addsub.genblk1[1].fa.a ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold19 (.A(_019_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold20 (.A(\aluobj.addsub.op_b[0] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold21 (.A(_009_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold22 (.A(\aluobj.addsub.genblk1[4].fa.a ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold23 (.A(_022_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold24 (.A(\aluobj.addsub.genblk1[6].fa.a ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold25 (.A(_024_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold26 (.A(\aluobj.addsub.genblk1[2].fa.a ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold27 (.A(_020_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold28 (.A(\aluobj.addsub.genblk1[0].fa.a ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold29 (.A(_018_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold30 (.A(\aluobj.addsub.genblk1[3].fa.a ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold31 (.A(_021_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold32 (.A(\aluobj.addsub.genblk1[7].fa.a ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold33 (.A(_025_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold34 (.A(\aluobj.addsub.genblk1[5].fa.a ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold35 (.A(_023_),
    .X(net96));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_4 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_279 ();
 sg13g2_decap_8 FILLER_22_286 ();
 sg13g2_decap_8 FILLER_22_293 ();
 sg13g2_decap_8 FILLER_22_300 ();
 sg13g2_decap_8 FILLER_22_307 ();
 sg13g2_decap_8 FILLER_22_314 ();
 sg13g2_decap_8 FILLER_22_321 ();
 sg13g2_decap_8 FILLER_22_328 ();
 sg13g2_decap_8 FILLER_22_335 ();
 sg13g2_decap_8 FILLER_22_342 ();
 sg13g2_decap_8 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_decap_8 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_370 ();
 sg13g2_decap_8 FILLER_22_377 ();
 sg13g2_decap_8 FILLER_22_384 ();
 sg13g2_decap_8 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_4 FILLER_23_182 ();
 sg13g2_fill_1 FILLER_23_186 ();
 sg13g2_decap_8 FILLER_23_221 ();
 sg13g2_decap_8 FILLER_23_228 ();
 sg13g2_decap_8 FILLER_23_235 ();
 sg13g2_fill_1 FILLER_23_242 ();
 sg13g2_decap_8 FILLER_23_277 ();
 sg13g2_decap_8 FILLER_23_295 ();
 sg13g2_decap_8 FILLER_23_302 ();
 sg13g2_fill_2 FILLER_23_309 ();
 sg13g2_fill_1 FILLER_23_311 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_4 FILLER_23_322 ();
 sg13g2_fill_2 FILLER_23_326 ();
 sg13g2_fill_2 FILLER_23_353 ();
 sg13g2_fill_1 FILLER_23_355 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_fill_2 FILLER_24_182 ();
 sg13g2_fill_1 FILLER_24_239 ();
 sg13g2_decap_4 FILLER_24_286 ();
 sg13g2_decap_8 FILLER_24_341 ();
 sg13g2_fill_1 FILLER_24_348 ();
 sg13g2_decap_8 FILLER_24_361 ();
 sg13g2_fill_2 FILLER_24_368 ();
 sg13g2_fill_1 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_374 ();
 sg13g2_decap_8 FILLER_24_381 ();
 sg13g2_decap_8 FILLER_24_388 ();
 sg13g2_decap_8 FILLER_24_395 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_4 FILLER_25_182 ();
 sg13g2_fill_1 FILLER_25_186 ();
 sg13g2_fill_1 FILLER_25_196 ();
 sg13g2_decap_4 FILLER_25_220 ();
 sg13g2_fill_1 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_fill_2 FILLER_25_336 ();
 sg13g2_fill_1 FILLER_25_338 ();
 sg13g2_decap_8 FILLER_25_395 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_fill_1 FILLER_26_168 ();
 sg13g2_fill_2 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_242 ();
 sg13g2_fill_1 FILLER_26_257 ();
 sg13g2_fill_2 FILLER_26_266 ();
 sg13g2_fill_1 FILLER_26_368 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_4 FILLER_27_147 ();
 sg13g2_fill_1 FILLER_27_151 ();
 sg13g2_fill_1 FILLER_27_221 ();
 sg13g2_fill_2 FILLER_27_235 ();
 sg13g2_fill_1 FILLER_27_237 ();
 sg13g2_fill_1 FILLER_27_282 ();
 sg13g2_fill_1 FILLER_27_300 ();
 sg13g2_fill_2 FILLER_27_335 ();
 sg13g2_fill_1 FILLER_27_340 ();
 sg13g2_fill_2 FILLER_27_349 ();
 sg13g2_decap_8 FILLER_27_356 ();
 sg13g2_decap_8 FILLER_27_363 ();
 sg13g2_fill_2 FILLER_27_370 ();
 sg13g2_fill_1 FILLER_27_372 ();
 sg13g2_decap_8 FILLER_27_376 ();
 sg13g2_decap_8 FILLER_27_383 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_4 FILLER_28_147 ();
 sg13g2_decap_4 FILLER_28_232 ();
 sg13g2_fill_1 FILLER_28_236 ();
 sg13g2_decap_4 FILLER_28_249 ();
 sg13g2_fill_2 FILLER_28_284 ();
 sg13g2_fill_1 FILLER_28_286 ();
 sg13g2_fill_1 FILLER_28_363 ();
 sg13g2_fill_2 FILLER_28_368 ();
 sg13g2_decap_8 FILLER_28_395 ();
 sg13g2_decap_8 FILLER_28_402 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_fill_1 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_193 ();
 sg13g2_fill_2 FILLER_29_200 ();
 sg13g2_decap_4 FILLER_29_216 ();
 sg13g2_fill_2 FILLER_29_220 ();
 sg13g2_fill_2 FILLER_29_227 ();
 sg13g2_decap_4 FILLER_29_254 ();
 sg13g2_fill_1 FILLER_29_258 ();
 sg13g2_fill_1 FILLER_29_267 ();
 sg13g2_decap_4 FILLER_29_276 ();
 sg13g2_decap_8 FILLER_29_303 ();
 sg13g2_fill_1 FILLER_29_310 ();
 sg13g2_fill_2 FILLER_29_321 ();
 sg13g2_decap_8 FILLER_29_327 ();
 sg13g2_decap_8 FILLER_29_334 ();
 sg13g2_fill_2 FILLER_29_341 ();
 sg13g2_fill_1 FILLER_29_343 ();
 sg13g2_decap_4 FILLER_29_347 ();
 sg13g2_fill_2 FILLER_29_351 ();
 sg13g2_decap_8 FILLER_29_379 ();
 sg13g2_decap_8 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_fill_2 FILLER_30_165 ();
 sg13g2_fill_1 FILLER_30_167 ();
 sg13g2_decap_8 FILLER_30_230 ();
 sg13g2_decap_4 FILLER_30_248 ();
 sg13g2_decap_4 FILLER_30_281 ();
 sg13g2_decap_4 FILLER_30_369 ();
 sg13g2_fill_1 FILLER_30_373 ();
 sg13g2_decap_8 FILLER_30_377 ();
 sg13g2_decap_8 FILLER_30_384 ();
 sg13g2_decap_8 FILLER_30_391 ();
 sg13g2_decap_8 FILLER_30_398 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_fill_1 FILLER_31_191 ();
 sg13g2_decap_4 FILLER_31_202 ();
 sg13g2_fill_1 FILLER_31_229 ();
 sg13g2_decap_4 FILLER_31_255 ();
 sg13g2_fill_2 FILLER_31_259 ();
 sg13g2_fill_1 FILLER_31_278 ();
 sg13g2_fill_2 FILLER_31_305 ();
 sg13g2_fill_1 FILLER_31_307 ();
 sg13g2_decap_8 FILLER_31_316 ();
 sg13g2_decap_4 FILLER_31_323 ();
 sg13g2_fill_2 FILLER_31_327 ();
 sg13g2_decap_4 FILLER_31_333 ();
 sg13g2_fill_1 FILLER_31_337 ();
 sg13g2_decap_8 FILLER_31_343 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_fill_2 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_176 ();
 sg13g2_fill_1 FILLER_32_183 ();
 sg13g2_decap_8 FILLER_32_228 ();
 sg13g2_fill_2 FILLER_32_249 ();
 sg13g2_decap_4 FILLER_32_287 ();
 sg13g2_fill_1 FILLER_32_291 ();
 sg13g2_fill_1 FILLER_32_322 ();
 sg13g2_decap_8 FILLER_32_352 ();
 sg13g2_decap_8 FILLER_32_359 ();
 sg13g2_decap_8 FILLER_32_370 ();
 sg13g2_decap_8 FILLER_32_377 ();
 sg13g2_decap_8 FILLER_32_384 ();
 sg13g2_decap_8 FILLER_32_391 ();
 sg13g2_decap_8 FILLER_32_398 ();
 sg13g2_decap_4 FILLER_32_405 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_fill_1 FILLER_33_147 ();
 sg13g2_decap_4 FILLER_33_151 ();
 sg13g2_fill_1 FILLER_33_155 ();
 sg13g2_fill_1 FILLER_33_235 ();
 sg13g2_decap_8 FILLER_33_242 ();
 sg13g2_fill_1 FILLER_33_283 ();
 sg13g2_fill_2 FILLER_33_312 ();
 sg13g2_fill_1 FILLER_33_314 ();
 sg13g2_fill_1 FILLER_33_318 ();
 sg13g2_decap_8 FILLER_33_327 ();
 sg13g2_fill_2 FILLER_33_334 ();
 sg13g2_fill_1 FILLER_33_336 ();
 sg13g2_decap_8 FILLER_33_363 ();
 sg13g2_decap_8 FILLER_33_370 ();
 sg13g2_decap_8 FILLER_33_377 ();
 sg13g2_decap_8 FILLER_33_384 ();
 sg13g2_decap_8 FILLER_33_391 ();
 sg13g2_decap_8 FILLER_33_398 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_4 FILLER_34_147 ();
 sg13g2_fill_2 FILLER_34_151 ();
 sg13g2_fill_1 FILLER_34_201 ();
 sg13g2_decap_4 FILLER_34_257 ();
 sg13g2_fill_2 FILLER_34_279 ();
 sg13g2_fill_1 FILLER_34_281 ();
 sg13g2_fill_2 FILLER_34_301 ();
 sg13g2_fill_1 FILLER_34_303 ();
 sg13g2_decap_8 FILLER_34_332 ();
 sg13g2_fill_1 FILLER_34_339 ();
 sg13g2_fill_1 FILLER_34_365 ();
 sg13g2_decap_8 FILLER_34_391 ();
 sg13g2_decap_8 FILLER_34_398 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_4 FILLER_35_161 ();
 sg13g2_fill_1 FILLER_35_165 ();
 sg13g2_fill_1 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_185 ();
 sg13g2_decap_8 FILLER_35_192 ();
 sg13g2_fill_2 FILLER_35_199 ();
 sg13g2_fill_2 FILLER_35_221 ();
 sg13g2_decap_4 FILLER_35_230 ();
 sg13g2_fill_2 FILLER_35_234 ();
 sg13g2_decap_4 FILLER_35_241 ();
 sg13g2_fill_1 FILLER_35_245 ();
 sg13g2_fill_2 FILLER_35_250 ();
 sg13g2_fill_1 FILLER_35_252 ();
 sg13g2_decap_4 FILLER_35_320 ();
 sg13g2_decap_8 FILLER_35_353 ();
 sg13g2_decap_8 FILLER_35_360 ();
 sg13g2_decap_8 FILLER_35_367 ();
 sg13g2_decap_8 FILLER_35_374 ();
 sg13g2_decap_8 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_35_396 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_4 FILLER_36_168 ();
 sg13g2_fill_1 FILLER_36_232 ();
 sg13g2_decap_8 FILLER_36_277 ();
 sg13g2_fill_1 FILLER_36_284 ();
 sg13g2_decap_4 FILLER_36_295 ();
 sg13g2_fill_1 FILLER_36_299 ();
 sg13g2_decap_8 FILLER_36_309 ();
 sg13g2_fill_2 FILLER_36_316 ();
 sg13g2_fill_1 FILLER_36_318 ();
 sg13g2_decap_8 FILLER_36_324 ();
 sg13g2_decap_4 FILLER_36_331 ();
 sg13g2_decap_8 FILLER_36_339 ();
 sg13g2_decap_8 FILLER_36_346 ();
 sg13g2_decap_8 FILLER_36_353 ();
 sg13g2_decap_8 FILLER_36_360 ();
 sg13g2_decap_8 FILLER_36_367 ();
 sg13g2_decap_8 FILLER_36_374 ();
 sg13g2_decap_8 FILLER_36_381 ();
 sg13g2_decap_8 FILLER_36_388 ();
 sg13g2_decap_8 FILLER_36_395 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_4 FILLER_37_196 ();
 sg13g2_decap_4 FILLER_37_204 ();
 sg13g2_decap_8 FILLER_37_212 ();
 sg13g2_decap_8 FILLER_37_219 ();
 sg13g2_decap_8 FILLER_37_226 ();
 sg13g2_decap_8 FILLER_37_233 ();
 sg13g2_decap_4 FILLER_37_240 ();
 sg13g2_decap_8 FILLER_37_248 ();
 sg13g2_decap_8 FILLER_37_255 ();
 sg13g2_decap_8 FILLER_37_262 ();
 sg13g2_fill_1 FILLER_37_269 ();
 sg13g2_decap_8 FILLER_37_295 ();
 sg13g2_decap_8 FILLER_37_302 ();
 sg13g2_decap_8 FILLER_37_309 ();
 sg13g2_decap_8 FILLER_37_316 ();
 sg13g2_decap_8 FILLER_37_323 ();
 sg13g2_decap_8 FILLER_37_330 ();
 sg13g2_decap_8 FILLER_37_337 ();
 sg13g2_decap_8 FILLER_37_344 ();
 sg13g2_decap_8 FILLER_37_351 ();
 sg13g2_decap_8 FILLER_37_358 ();
 sg13g2_decap_8 FILLER_37_365 ();
 sg13g2_decap_8 FILLER_37_372 ();
 sg13g2_decap_8 FILLER_37_379 ();
 sg13g2_decap_8 FILLER_37_386 ();
 sg13g2_decap_8 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_8 FILLER_38_164 ();
 sg13g2_decap_8 FILLER_38_171 ();
 sg13g2_decap_8 FILLER_38_178 ();
 sg13g2_decap_8 FILLER_38_185 ();
 sg13g2_decap_8 FILLER_38_192 ();
 sg13g2_decap_8 FILLER_38_199 ();
 sg13g2_decap_8 FILLER_38_206 ();
 sg13g2_decap_8 FILLER_38_213 ();
 sg13g2_decap_8 FILLER_38_220 ();
 sg13g2_decap_8 FILLER_38_227 ();
 sg13g2_decap_8 FILLER_38_234 ();
 sg13g2_decap_8 FILLER_38_241 ();
 sg13g2_fill_1 FILLER_38_272 ();
 sg13g2_fill_2 FILLER_38_286 ();
 sg13g2_decap_4 FILLER_38_308 ();
 sg13g2_decap_4 FILLER_38_316 ();
 sg13g2_decap_4 FILLER_38_324 ();
 sg13g2_decap_4 FILLER_38_332 ();
 sg13g2_decap_4 FILLER_38_340 ();
 sg13g2_decap_4 FILLER_38_348 ();
 sg13g2_decap_4 FILLER_38_356 ();
 sg13g2_decap_4 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net52;
 assign uio_oe[1] = net53;
 assign uio_oe[2] = net30;
 assign uio_oe[3] = net31;
 assign uio_oe[4] = net32;
 assign uio_oe[5] = net33;
 assign uio_oe[6] = net34;
 assign uio_oe[7] = net35;
 assign uio_out[2] = net36;
 assign uio_out[3] = net37;
 assign uio_out[4] = net38;
 assign uio_out[5] = net39;
 assign uio_out[6] = net40;
 assign uio_out[7] = net41;
endmodule

module tt_um_find_the_damn_issue (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire net529;
 wire clk_regs;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire n106_o;
 wire n118_o;
 wire n124_o;
 wire n130_o;
 wire n136_o;
 wire n153_o;
 wire n183_o;
 wire n346_q;
 wire n347_q;
 wire n349_q;
 wire n350_o;
 wire n351_q;
 wire \n352_o[0] ;
 wire \n352_o[10] ;
 wire \n352_o[11] ;
 wire \n352_o[12] ;
 wire \n352_o[13] ;
 wire \n352_o[17] ;
 wire \n352_o[18] ;
 wire \n352_o[19] ;
 wire \n352_o[1] ;
 wire \n352_o[20] ;
 wire \n352_o[21] ;
 wire \n352_o[22] ;
 wire \n352_o[23] ;
 wire \n352_o[2] ;
 wire \n352_o[3] ;
 wire \n352_o[4] ;
 wire \n352_o[5] ;
 wire \n352_o[6] ;
 wire \n352_o[7] ;
 wire \n352_o[8] ;
 wire \n353_q[0] ;
 wire \n353_q[10] ;
 wire \n353_q[11] ;
 wire \n353_q[12] ;
 wire \n353_q[13] ;
 wire \n353_q[14] ;
 wire \n353_q[15] ;
 wire \n353_q[16] ;
 wire \n353_q[17] ;
 wire \n353_q[18] ;
 wire \n353_q[19] ;
 wire \n353_q[1] ;
 wire \n353_q[20] ;
 wire \n353_q[21] ;
 wire \n353_q[22] ;
 wire \n353_q[23] ;
 wire \n353_q[2] ;
 wire \n353_q[3] ;
 wire \n353_q[4] ;
 wire \n353_q[5] ;
 wire \n353_q[6] ;
 wire \n353_q[7] ;
 wire \n353_q[8] ;
 wire \n353_q[9] ;
 wire s_m_io0_en;
 wire s_m_io0_opendrain;
 wire s_m_io0_out;
 wire s_m_io10_out;
 wire s_m_io11_out;
 wire s_m_io12_out;
 wire s_m_io13_out;
 wire s_m_io14_out;
 wire s_m_io15_out;
 wire s_m_io1_en;
 wire s_m_io1_opendrain;
 wire s_m_io1_out;
 wire s_m_io2_en;
 wire s_m_io2_opendrain;
 wire s_m_io2_out;
 wire s_m_io3_en;
 wire s_m_io3_opendrain;
 wire s_m_io3_out;
 wire s_m_io4_en;
 wire s_m_io4_opendrain;
 wire s_m_io4_out;
 wire s_m_io5_en;
 wire s_m_io5_opendrain;
 wire s_m_io5_out;
 wire s_m_io9_out;
 wire s_m_match_delayed1;
 wire s_m_packetdata_2_bit_16;
 wire s_m_packetdata_2_bit_17;
 wire \s_m_packetdata_2_rewired[0] ;
 wire \s_m_packetdata_2_rewired[10] ;
 wire \s_m_packetdata_2_rewired[11] ;
 wire \s_m_packetdata_2_rewired[12] ;
 wire \s_m_packetdata_2_rewired[13] ;
 wire \s_m_packetdata_2_rewired[14] ;
 wire \s_m_packetdata_2_rewired[15] ;
 wire \s_m_packetdata_2_rewired[18] ;
 wire \s_m_packetdata_2_rewired[19] ;
 wire \s_m_packetdata_2_rewired[1] ;
 wire \s_m_packetdata_2_rewired[20] ;
 wire \s_m_packetdata_2_rewired[21] ;
 wire \s_m_packetdata_2_rewired[22] ;
 wire \s_m_packetdata_2_rewired[23] ;
 wire \s_m_packetdata_2_rewired[2] ;
 wire \s_m_packetdata_2_rewired[3] ;
 wire \s_m_packetdata_2_rewired[4] ;
 wire \s_m_packetdata_2_rewired[5] ;
 wire \s_m_packetdata_2_rewired[6] ;
 wire \s_m_packetdata_2_rewired[7] ;
 wire \s_m_packetdata_2_rewired[8] ;
 wire \s_m_packetdata_2_rewired[9] ;
 wire \s_m_peekdata_data_2[0] ;
 wire \s_m_peekdata_data_2[1] ;
 wire \s_m_peekdata_data_2[2] ;
 wire \s_m_peekdata_data_2[3] ;
 wire \s_m_peekdata_data_2[4] ;
 wire \s_m_peekdata_data_2[5] ;
 wire \s_m_peekdata_data_2[6] ;
 wire \s_m_peekdata_data_2[7] ;
 wire s_m_phy_tx_valid_2;
 wire s_m_popempty;
 wire s_m_popempty_2;
 wire \s_m_pushdata_data[0] ;
 wire \s_m_pushdata_data[1] ;
 wire \s_m_pushdata_data[2] ;
 wire \s_m_pushdata_data[3] ;
 wire \s_m_pushdata_data[4] ;
 wire \s_m_pushdata_data[5] ;
 wire \s_m_pushdata_data[6] ;
 wire \s_m_pushdata_data[7] ;
 wire \s_m_pushdata_endpoint[0] ;
 wire \s_m_pushdata_endpoint[1] ;
 wire \s_m_pushdata_endpoint[2] ;
 wire \s_m_pushdata_endpoint[3] ;
 wire s_m_pushfull;
 wire s_m_pushfull_2;
 wire \s_m_status_linestate[0] ;
 wire \s_m_status_linestate[1] ;
 wire s_m_status_rxactive;
 wire \s_out_3[0] ;
 wire \s_out_3[1] ;
 wire \s_out_3[2] ;
 wire \s_out_3[3] ;
 wire \s_out_3[4] ;
 wire \s_out_3[5] ;
 wire \s_out_3[6] ;
 wire \s_out_3[7] ;
 wire s_out_valid_2;
 wire \scl_bitbangengine0.n3179_o ;
 wire \scl_bitbangengine0.n3198_o ;
 wire \scl_bitbangengine0.n3230_o ;
 wire \scl_bitbangengine0.n3241_o ;
 wire \scl_bitbangengine0.n3257_o ;
 wire \scl_bitbangengine0.n3258_o ;
 wire \scl_bitbangengine0.n3267_o ;
 wire \scl_bitbangengine0.n3336_o ;
 wire \scl_bitbangengine0.n3663_o[0] ;
 wire \scl_bitbangengine0.n3663_o[1] ;
 wire \scl_bitbangengine0.n3663_o[2] ;
 wire \scl_bitbangengine0.n3663_o[3] ;
 wire \scl_bitbangengine0.n3663_o[4] ;
 wire \scl_bitbangengine0.n3663_o[5] ;
 wire \scl_bitbangengine0.n3663_o[6] ;
 wire \scl_bitbangengine0.n3663_o[7] ;
 wire \scl_bitbangengine0.n3663_o[8] ;
 wire \scl_bitbangengine0.n3737_o ;
 wire \scl_bitbangengine0.n3740_o ;
 wire \scl_bitbangengine0.n3793_o ;
 wire \scl_bitbangengine0.n3817_o ;
 wire \scl_bitbangengine0.n3839_o ;
 wire \scl_bitbangengine0.n3865_o ;
 wire \scl_bitbangengine0.n3871_o ;
 wire \scl_bitbangengine0.n5401_o ;
 wire \scl_bitbangengine0.n5423_o[0] ;
 wire \scl_bitbangengine0.n5423_o[1] ;
 wire \scl_bitbangengine0.n5423_o[2] ;
 wire \scl_bitbangengine0.n5423_o[3] ;
 wire \scl_bitbangengine0.n5423_o[4] ;
 wire \scl_bitbangengine0.n5423_o[5] ;
 wire \scl_bitbangengine0.n5423_o[6] ;
 wire \scl_bitbangengine0.n5462_o[0] ;
 wire \scl_bitbangengine0.n5462_o[1] ;
 wire \scl_bitbangengine0.n5462_o[2] ;
 wire \scl_bitbangengine0.n5462_o[3] ;
 wire \scl_bitbangengine0.n5462_o[4] ;
 wire \scl_bitbangengine0.n5462_o[5] ;
 wire \scl_bitbangengine0.n5462_o[6] ;
 wire \scl_bitbangengine0.n5462_o[7] ;
 wire \scl_bitbangengine0.n5898_q[0] ;
 wire \scl_bitbangengine0.n5898_q[1] ;
 wire \scl_bitbangengine0.n5898_q[2] ;
 wire \scl_bitbangengine0.n5898_q[3] ;
 wire \scl_bitbangengine0.n5902_q ;
 wire \scl_bitbangengine0.n5903_q ;
 wire \scl_bitbangengine0.n5904_q ;
 wire \scl_bitbangengine0.n5905_q ;
 wire \scl_bitbangengine0.n5907_q ;
 wire \scl_bitbangengine0.n5909_q ;
 wire \scl_bitbangengine0.n5910_q ;
 wire \scl_bitbangengine0.n5911_q ;
 wire \scl_bitbangengine0.n5913_q ;
 wire \scl_bitbangengine0.n5915_q ;
 wire \scl_bitbangengine0.n5917_q ;
 wire \scl_bitbangengine0.n5918_q ;
 wire \scl_bitbangengine0.n5919_q ;
 wire \scl_bitbangengine0.n5920_q[0] ;
 wire \scl_bitbangengine0.n5920_q[10] ;
 wire \scl_bitbangengine0.n5920_q[11] ;
 wire \scl_bitbangengine0.n5920_q[12] ;
 wire \scl_bitbangengine0.n5920_q[13] ;
 wire \scl_bitbangengine0.n5920_q[14] ;
 wire \scl_bitbangengine0.n5920_q[15] ;
 wire \scl_bitbangengine0.n5920_q[16] ;
 wire \scl_bitbangengine0.n5920_q[17] ;
 wire \scl_bitbangengine0.n5920_q[18] ;
 wire \scl_bitbangengine0.n5920_q[19] ;
 wire \scl_bitbangengine0.n5920_q[1] ;
 wire \scl_bitbangengine0.n5920_q[2] ;
 wire \scl_bitbangengine0.n5920_q[3] ;
 wire \scl_bitbangengine0.n5920_q[4] ;
 wire \scl_bitbangengine0.n5920_q[5] ;
 wire \scl_bitbangengine0.n5920_q[6] ;
 wire \scl_bitbangengine0.n5920_q[7] ;
 wire \scl_bitbangengine0.n5920_q[8] ;
 wire \scl_bitbangengine0.n5920_q[9] ;
 wire \scl_bitbangengine0.n5921_q[0] ;
 wire \scl_bitbangengine0.n5921_q[1] ;
 wire \scl_bitbangengine0.n5921_q[2] ;
 wire \scl_bitbangengine0.n5921_q[3] ;
 wire \scl_bitbangengine0.n5921_q[4] ;
 wire \scl_bitbangengine0.n5921_q[5] ;
 wire \scl_bitbangengine0.n5921_q[6] ;
 wire \scl_bitbangengine0.n5921_q[7] ;
 wire \scl_bitbangengine0.n5923_q ;
 wire \scl_bitbangengine0.n5924_q[7] ;
 wire \scl_bitbangengine0.s_m_value[0] ;
 wire \scl_bitbangengine0.s_m_value[1] ;
 wire \scl_bitbangengine0.s_m_value[2] ;
 wire \scl_bitbangengine0.s_m_value_2[0] ;
 wire \scl_bitbangengine0.s_m_value_2[1] ;
 wire \scl_bitbangengine0.s_m_value_2[2] ;
 wire \scl_bitbangengine0.scl_counter0.n6954_o[0] ;
 wire \scl_bitbangengine0.scl_counter0.n6954_o[10] ;
 wire \scl_bitbangengine0.scl_counter0.n6954_o[11] ;
 wire \scl_bitbangengine0.scl_counter0.n6954_o[12] ;
 wire \scl_bitbangengine0.scl_counter0.n6954_o[13] ;
 wire \scl_bitbangengine0.scl_counter0.n6954_o[14] ;
 wire \scl_bitbangengine0.scl_counter0.n6954_o[15] ;
 wire \scl_bitbangengine0.scl_counter0.n6954_o[16] ;
 wire \scl_bitbangengine0.scl_counter0.n6954_o[1] ;
 wire \scl_bitbangengine0.scl_counter0.n6954_o[2] ;
 wire \scl_bitbangengine0.scl_counter0.n6954_o[3] ;
 wire \scl_bitbangengine0.scl_counter0.n6954_o[4] ;
 wire \scl_bitbangengine0.scl_counter0.n6954_o[5] ;
 wire \scl_bitbangengine0.scl_counter0.n6954_o[6] ;
 wire \scl_bitbangengine0.scl_counter0.n6954_o[7] ;
 wire \scl_bitbangengine0.scl_counter0.n6954_o[8] ;
 wire \scl_bitbangengine0.scl_counter0.n6954_o[9] ;
 wire \scl_bitbangengine0.scl_counter0.n6975_q[0] ;
 wire \scl_bitbangengine0.scl_counter0.n6975_q[10] ;
 wire \scl_bitbangengine0.scl_counter0.n6975_q[11] ;
 wire \scl_bitbangengine0.scl_counter0.n6975_q[12] ;
 wire \scl_bitbangengine0.scl_counter0.n6975_q[13] ;
 wire \scl_bitbangengine0.scl_counter0.n6975_q[14] ;
 wire \scl_bitbangengine0.scl_counter0.n6975_q[15] ;
 wire \scl_bitbangengine0.scl_counter0.n6975_q[16] ;
 wire \scl_bitbangengine0.scl_counter0.n6975_q[1] ;
 wire \scl_bitbangengine0.scl_counter0.n6975_q[2] ;
 wire \scl_bitbangengine0.scl_counter0.n6975_q[3] ;
 wire \scl_bitbangengine0.scl_counter0.n6975_q[4] ;
 wire \scl_bitbangengine0.scl_counter0.n6975_q[5] ;
 wire \scl_bitbangengine0.scl_counter0.n6975_q[6] ;
 wire \scl_bitbangengine0.scl_counter0.n6975_q[7] ;
 wire \scl_bitbangengine0.scl_counter0.n6975_q[8] ;
 wire \scl_bitbangengine0.scl_counter0.n6975_q[9] ;
 wire \scl_fifo0.n2689_o[0] ;
 wire \scl_fifo0.n2689_o[1] ;
 wire \scl_fifo0.n2689_o[2] ;
 wire \scl_fifo0.n2689_o[3] ;
 wire \scl_fifo0.n2694_o[0] ;
 wire \scl_fifo0.n2697_o[0] ;
 wire \scl_fifo0.n2697_o[1] ;
 wire \scl_fifo0.n2697_o[2] ;
 wire \scl_fifo0.n2697_o[3] ;
 wire \scl_fifo0.n2697_o[4] ;
 wire \scl_fifo0.n2700_o ;
 wire \scl_fifo0.n2711_o[0] ;
 wire \scl_fifo0.n2711_o[1] ;
 wire \scl_fifo0.n2711_o[2] ;
 wire \scl_fifo0.n2711_o[3] ;
 wire \scl_fifo0.n2722_o[1] ;
 wire \scl_fifo0.n2722_o[2] ;
 wire \scl_fifo0.n2722_o[3] ;
 wire \scl_fifo0.n2722_o[4] ;
 wire \scl_fifo0.n2726_o ;
 wire \scl_fifo0.n2737_o[0] ;
 wire \scl_fifo0.n2737_o[1] ;
 wire \scl_fifo0.n2737_o[2] ;
 wire \scl_fifo0.n2737_o[3] ;
 wire \scl_fifo0.n2746_o ;
 wire \scl_fifo0.n2781_q[4] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[0][0] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[0][1] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[0][2] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[0][3] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[0][4] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[0][5] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[0][6] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[0][7] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[10][0] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[10][1] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[10][2] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[10][3] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[10][4] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[10][5] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[10][6] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[10][7] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[11][0] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[11][1] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[11][2] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[11][3] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[11][4] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[11][5] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[11][6] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[11][7] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[12][0] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[12][1] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[12][2] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[12][3] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[12][4] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[12][5] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[12][6] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[12][7] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[13][0] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[13][1] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[13][2] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[13][3] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[13][4] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[13][5] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[13][6] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[13][7] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[14][0] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[14][1] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[14][2] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[14][3] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[14][4] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[14][5] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[14][6] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[14][7] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[15][0] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[15][1] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[15][2] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[15][3] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[15][4] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[15][5] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[15][6] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[15][7] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[1][0] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[1][1] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[1][2] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[1][3] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[1][4] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[1][5] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[1][6] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[1][7] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[2][0] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[2][1] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[2][2] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[2][3] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[2][4] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[2][5] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[2][6] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[2][7] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[3][0] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[3][1] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[3][2] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[3][3] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[3][4] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[3][5] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[3][6] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[3][7] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[4][0] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[4][1] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[4][2] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[4][3] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[4][4] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[4][5] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[4][6] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[4][7] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[5][0] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[5][1] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[5][2] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[5][3] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[5][4] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[5][5] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[5][6] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[5][7] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[6][0] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[6][1] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[6][2] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[6][3] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[6][4] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[6][5] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[6][6] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[6][7] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[7][0] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[7][1] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[7][2] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[7][3] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[7][4] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[7][5] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[7][6] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[7][7] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[8][0] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[8][1] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[8][2] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[8][3] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[8][4] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[8][5] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[8][6] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[8][7] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[9][0] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[9][1] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[9][2] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[9][3] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[9][4] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[9][5] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[9][6] ;
 wire \scl_fifo0.scl_memory0.physical_memory0.memory[9][7] ;
 wire \scl_fifo1.n6229_o[0] ;
 wire \scl_fifo1.n6229_o[1] ;
 wire \scl_fifo1.n6229_o[2] ;
 wire \scl_fifo1.n6229_o[3] ;
 wire \scl_fifo1.n6233_o[0] ;
 wire \scl_fifo1.n6233_o[1] ;
 wire \scl_fifo1.n6233_o[2] ;
 wire \scl_fifo1.n6233_o[3] ;
 wire \scl_fifo1.n6233_o[4] ;
 wire \scl_fifo1.n6238_o[0] ;
 wire \scl_fifo1.n6238_o[1] ;
 wire \scl_fifo1.n6238_o[2] ;
 wire \scl_fifo1.n6238_o[3] ;
 wire \scl_fifo1.n6238_o[4] ;
 wire \scl_fifo1.n6239_o[0] ;
 wire \scl_fifo1.n6239_o[1] ;
 wire \scl_fifo1.n6239_o[2] ;
 wire \scl_fifo1.n6239_o[3] ;
 wire \scl_fifo1.n6239_o[4] ;
 wire \scl_fifo1.n6242_o ;
 wire \scl_fifo1.n6267_o ;
 wire \scl_fifo1.n6278_o[0] ;
 wire \scl_fifo1.n6278_o[1] ;
 wire \scl_fifo1.n6278_o[2] ;
 wire \scl_fifo1.n6278_o[3] ;
 wire \scl_fifo1.n6287_o ;
 wire \scl_fifo1.n6321_q[0] ;
 wire \scl_fifo1.n6321_q[1] ;
 wire \scl_fifo1.n6321_q[2] ;
 wire \scl_fifo1.n6321_q[3] ;
 wire \scl_fifo1.n6321_q[4] ;
 wire \scl_fifo1.n6323_q[0] ;
 wire \scl_fifo1.n6323_q[1] ;
 wire \scl_fifo1.n6323_q[2] ;
 wire \scl_fifo1.n6323_q[3] ;
 wire \scl_fifo1.n6323_q[4] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[0][0] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[0][1] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[0][2] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[0][3] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[0][4] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[0][5] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[0][6] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[0][7] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[10][0] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[10][1] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[10][2] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[10][3] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[10][4] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[10][5] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[10][6] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[10][7] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[11][0] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[11][1] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[11][2] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[11][3] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[11][4] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[11][5] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[11][6] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[11][7] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[12][0] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[12][1] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[12][2] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[12][3] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[12][4] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[12][5] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[12][6] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[12][7] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[13][0] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[13][1] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[13][2] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[13][3] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[13][4] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[13][5] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[13][6] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[13][7] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[14][0] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[14][1] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[14][2] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[14][3] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[14][4] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[14][5] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[14][6] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[14][7] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[15][0] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[15][1] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[15][2] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[15][3] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[15][4] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[15][5] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[15][6] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[15][7] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[1][0] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[1][1] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[1][2] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[1][3] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[1][4] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[1][5] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[1][6] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[1][7] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[2][0] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[2][1] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[2][2] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[2][3] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[2][4] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[2][5] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[2][6] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[2][7] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[3][0] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[3][1] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[3][2] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[3][3] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[3][4] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[3][5] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[3][6] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[3][7] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[4][0] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[4][1] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[4][2] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[4][3] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[4][4] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[4][5] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[4][6] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[4][7] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[5][0] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[5][1] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[5][2] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[5][3] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[5][4] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[5][5] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[5][6] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[5][7] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[6][0] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[6][1] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[6][2] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[6][3] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[6][4] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[6][5] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[6][6] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[6][7] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[7][0] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[7][1] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[7][2] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[7][3] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[7][4] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[7][5] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[7][6] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[7][7] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[8][0] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[8][1] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[8][2] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[8][3] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[8][4] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[8][5] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[8][6] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[8][7] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[9][0] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[9][1] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[9][2] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[9][3] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[9][4] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[9][5] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[9][6] ;
 wire \scl_fifo1.scl_memory0.physical_memory0.memory[9][7] ;
 wire \scl_streamarbiter_2.n6146_o ;
 wire \scl_streamarbiter_2.n6171_o ;
 wire \scl_streamarbiter_2.n6192_q ;
 wire \scl_streamarbiter_2.n6194_q ;
 wire \scl_streamarbiter_2.n6195_q ;
 wire \scl_uartrx0.n5991_o ;
 wire \scl_uartrx0.n6047_o ;
 wire \scl_uartrx0.n6053_o ;
 wire \scl_uartrx0.n6074_o ;
 wire \scl_uartrx0.n6090_o ;
 wire \scl_uartrx0.n6119_q ;
 wire \scl_uartrx0.s_m_value[0] ;
 wire \scl_uartrx0.s_m_value[1] ;
 wire \scl_uartrx0.s_m_value[2] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7047_o[0] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7047_o[10] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7047_o[11] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7047_o[12] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7047_o[13] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7047_o[14] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7047_o[15] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7047_o[16] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7047_o[1] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7047_o[2] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7047_o[3] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7047_o[4] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7047_o[5] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7047_o[6] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7047_o[7] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7047_o[8] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7047_o[9] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7069_o[0] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7069_o[10] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7069_o[11] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7069_o[12] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7069_o[13] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7069_o[14] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7069_o[15] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7069_o[16] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7069_o[1] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7069_o[2] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7069_o[3] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7069_o[4] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7069_o[5] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7069_o[6] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7069_o[7] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7069_o[8] ;
 wire \scl_uartrx0.scl_baudrategenerator0.n7069_o[9] ;
 wire \scl_uarttx0.n2856_o[0] ;
 wire \scl_uarttx0.n2856_o[1] ;
 wire \scl_uarttx0.n2856_o[2] ;
 wire \scl_uarttx0.n2884_o ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6874_o[0] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6874_o[10] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6874_o[11] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6874_o[12] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6874_o[13] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6874_o[14] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6874_o[15] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6874_o[16] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6874_o[1] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6874_o[2] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6874_o[3] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6874_o[4] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6874_o[5] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6874_o[6] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6874_o[7] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6874_o[8] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6874_o[9] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6878_o[0] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6892_o[10] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6892_o[11] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6892_o[12] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6892_o[13] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6892_o[14] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6892_o[15] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6892_o[16] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6892_o[1] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6892_o[2] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6892_o[3] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6892_o[4] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6892_o[5] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6892_o[6] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6892_o[7] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6892_o[8] ;
 wire \scl_uarttx0.scl_baudrategenerator0.n6892_o[9] ;
 wire \scl_uarttx0.scl_counter0.n6919_o[0] ;
 wire \scl_uarttx0.scl_counter0.n6919_o[1] ;
 wire \scl_uarttx0.scl_counter0.n6919_o[3] ;
 wire \usbfunction0.functionreset0.in_unnamed[0] ;
 wire \usbfunction0.functionreset0.in_unnamed[1] ;
 wire \usbfunction0.functionreset0.in_unnamed[2] ;
 wire \usbfunction0.functionreset0.in_unnamed[3] ;
 wire \usbfunction0.functionreset0.in_unnamed[4] ;
 wire \usbfunction0.functionreset0.in_unnamed[5] ;
 wire \usbfunction0.functionreset0.in_unnamed[6] ;
 wire \usbfunction0.functionreset0.in_unnamed_2[0] ;
 wire \usbfunction0.functionreset0.in_unnamed_2[1] ;
 wire \usbfunction0.functionreset0.in_unnamed_2[2] ;
 wire \usbfunction0.functionreset0.in_unnamed_2[3] ;
 wire \usbfunction0.functionreset0.in_unnamed_3[0] ;
 wire \usbfunction0.functionreset0.in_unnamed_3[1] ;
 wire \usbfunction0.functionreset0.in_unnamed_3[2] ;
 wire \usbfunction0.functionreset0.in_unnamed_3[3] ;
 wire \usbfunction0.functionreset0.in_unnamed_3[4] ;
 wire \usbfunction0.functionreset0.in_unnamed_3[5] ;
 wire \usbfunction0.functionreset0.in_unnamed_3[6] ;
 wire \usbfunction0.functionreset0.in_unnamed_4[0] ;
 wire \usbfunction0.functionreset0.in_unnamed_4[1] ;
 wire \usbfunction0.functionreset0.n6674_o[0] ;
 wire \usbfunction0.functionreset0.n6674_o[1] ;
 wire \usbfunction0.functionreset0.n6674_o[2] ;
 wire \usbfunction0.functionreset0.n6674_o[3] ;
 wire \usbfunction0.functionreset0.n6674_o[4] ;
 wire \usbfunction0.functionreset0.n6674_o[5] ;
 wire \usbfunction0.functionreset0.n6674_o[6] ;
 wire \usbfunction0.functionreset0.n6674_o[7] ;
 wire \usbfunction0.functionreset0.n6674_o[8] ;
 wire \usbfunction0.functionreset0.n6674_o[9] ;
 wire \usbfunction0.functionreset0.n6683_o ;
 wire \usbfunction0.functionreset0.n6707_q[0] ;
 wire \usbfunction0.functionreset0.n6707_q[1] ;
 wire \usbfunction0.functionreset0.n6707_q[2] ;
 wire \usbfunction0.functionreset0.n6707_q[3] ;
 wire \usbfunction0.functionreset0.n6707_q[4] ;
 wire \usbfunction0.functionreset0.n6707_q[5] ;
 wire \usbfunction0.functionreset0.n6707_q[6] ;
 wire \usbfunction0.functionreset0.n6707_q[7] ;
 wire \usbfunction0.functionreset0.n6707_q[8] ;
 wire \usbfunction0.functionreset0.n6707_q[9] ;
 wire \usbfunction0.functionreset0.n6708_q ;
 wire \usbfunction0.n1083_o[0] ;
 wire \usbfunction0.n1083_o[1] ;
 wire \usbfunction0.n1083_o[2] ;
 wire \usbfunction0.n1083_o[3] ;
 wire \usbfunction0.n1083_o[4] ;
 wire \usbfunction0.n1083_o[5] ;
 wire \usbfunction0.n1083_o[6] ;
 wire \usbfunction0.n1101_o[0] ;
 wire \usbfunction0.n1101_o[1] ;
 wire \usbfunction0.n1101_o[2] ;
 wire \usbfunction0.n1101_o[3] ;
 wire \usbfunction0.n1101_o[4] ;
 wire \usbfunction0.n1101_o[5] ;
 wire \usbfunction0.n1101_o[6] ;
 wire \usbfunction0.n1101_o[7] ;
 wire \usbfunction0.n1189_o[0] ;
 wire \usbfunction0.n1189_o[1] ;
 wire \usbfunction0.n1189_o[2] ;
 wire \usbfunction0.n1189_o[3] ;
 wire \usbfunction0.n1359_o[0] ;
 wire \usbfunction0.n1359_o[1] ;
 wire \usbfunction0.n1360_o[0] ;
 wire \usbfunction0.n1360_o[1] ;
 wire \usbfunction0.n1360_o[2] ;
 wire \usbfunction0.n1360_o[3] ;
 wire \usbfunction0.n1581_o[0] ;
 wire \usbfunction0.n1581_o[1] ;
 wire \usbfunction0.n1583_o[0] ;
 wire \usbfunction0.n1583_o[1] ;
 wire \usbfunction0.n1583_o[2] ;
 wire \usbfunction0.n1583_o[3] ;
 wire \usbfunction0.n1583_o[4] ;
 wire \usbfunction0.n1583_o[5] ;
 wire \usbfunction0.n1583_o[6] ;
 wire \usbfunction0.n1630_o[0] ;
 wire \usbfunction0.n1630_o[10] ;
 wire \usbfunction0.n1630_o[11] ;
 wire \usbfunction0.n1630_o[12] ;
 wire \usbfunction0.n1630_o[13] ;
 wire \usbfunction0.n1630_o[14] ;
 wire \usbfunction0.n1630_o[15] ;
 wire \usbfunction0.n1630_o[1] ;
 wire \usbfunction0.n1630_o[2] ;
 wire \usbfunction0.n1630_o[3] ;
 wire \usbfunction0.n1630_o[4] ;
 wire \usbfunction0.n1630_o[5] ;
 wire \usbfunction0.n1630_o[6] ;
 wire \usbfunction0.n1630_o[7] ;
 wire \usbfunction0.n1630_o[8] ;
 wire \usbfunction0.n1630_o[9] ;
 wire \usbfunction0.n1687_o[0] ;
 wire \usbfunction0.n1687_o[10] ;
 wire \usbfunction0.n1687_o[11] ;
 wire \usbfunction0.n1687_o[12] ;
 wire \usbfunction0.n1687_o[13] ;
 wire \usbfunction0.n1687_o[14] ;
 wire \usbfunction0.n1687_o[1] ;
 wire \usbfunction0.n1687_o[2] ;
 wire \usbfunction0.n1687_o[3] ;
 wire \usbfunction0.n1687_o[4] ;
 wire \usbfunction0.n1687_o[5] ;
 wire \usbfunction0.n1687_o[6] ;
 wire \usbfunction0.n1687_o[7] ;
 wire \usbfunction0.n1687_o[8] ;
 wire \usbfunction0.n1687_o[9] ;
 wire \usbfunction0.n1974_o ;
 wire \usbfunction0.n2098_o ;
 wire \usbfunction0.n2254_o ;
 wire \usbfunction0.n2257_o[10] ;
 wire \usbfunction0.n2257_o[11] ;
 wire \usbfunction0.n2257_o[12] ;
 wire \usbfunction0.n2257_o[13] ;
 wire \usbfunction0.n2257_o[14] ;
 wire \usbfunction0.n2257_o[15] ;
 wire \usbfunction0.n2257_o[1] ;
 wire \usbfunction0.n2257_o[2] ;
 wire \usbfunction0.n2257_o[3] ;
 wire \usbfunction0.n2257_o[4] ;
 wire \usbfunction0.n2257_o[5] ;
 wire \usbfunction0.n2257_o[6] ;
 wire \usbfunction0.n2257_o[7] ;
 wire \usbfunction0.n2257_o[8] ;
 wire \usbfunction0.n2257_o[9] ;
 wire \usbfunction0.n2313_o[0] ;
 wire \usbfunction0.n2313_o[1] ;
 wire \usbfunction0.n2313_o[2] ;
 wire \usbfunction0.n2313_o[3] ;
 wire \usbfunction0.n2334_o[0] ;
 wire \usbfunction0.n2353_o[0] ;
 wire \usbfunction0.n2353_o[1] ;
 wire \usbfunction0.n2353_o[2] ;
 wire \usbfunction0.n2353_o[3] ;
 wire \usbfunction0.n2353_o[4] ;
 wire \usbfunction0.n2353_o[5] ;
 wire \usbfunction0.n2353_o[6] ;
 wire \usbfunction0.n2353_o[7] ;
 wire \usbfunction0.n2433_o[0] ;
 wire \usbfunction0.n2433_o[10] ;
 wire \usbfunction0.n2433_o[11] ;
 wire \usbfunction0.n2433_o[12] ;
 wire \usbfunction0.n2433_o[13] ;
 wire \usbfunction0.n2433_o[14] ;
 wire \usbfunction0.n2433_o[15] ;
 wire \usbfunction0.n2433_o[1] ;
 wire \usbfunction0.n2433_o[2] ;
 wire \usbfunction0.n2433_o[3] ;
 wire \usbfunction0.n2433_o[4] ;
 wire \usbfunction0.n2433_o[5] ;
 wire \usbfunction0.n2433_o[6] ;
 wire \usbfunction0.n2433_o[7] ;
 wire \usbfunction0.n2433_o[8] ;
 wire \usbfunction0.n2433_o[9] ;
 wire \usbfunction0.n2474_o[0] ;
 wire \usbfunction0.n2474_o[1] ;
 wire \usbfunction0.n2474_o[2] ;
 wire \usbfunction0.n2474_o[3] ;
 wire \usbfunction0.n2477_o[0] ;
 wire \usbfunction0.n2477_o[1] ;
 wire \usbfunction0.n2477_o[2] ;
 wire \usbfunction0.n2477_o[3] ;
 wire \usbfunction0.n2477_o[4] ;
 wire \usbfunction0.n2477_o[5] ;
 wire \usbfunction0.n2477_o[6] ;
 wire \usbfunction0.n2477_o[7] ;
 wire \usbfunction0.n2480_o[0] ;
 wire \usbfunction0.n2480_o[1] ;
 wire \usbfunction0.n2480_o[2] ;
 wire \usbfunction0.n2480_o[3] ;
 wire \usbfunction0.n2480_o[4] ;
 wire \usbfunction0.n2480_o[5] ;
 wire \usbfunction0.n2480_o[6] ;
 wire \usbfunction0.n2480_o[7] ;
 wire \usbfunction0.n2481_o[16] ;
 wire \usbfunction0.n2481_o[17] ;
 wire \usbfunction0.n2481_o[18] ;
 wire \usbfunction0.n2481_o[19] ;
 wire \usbfunction0.n2481_o[20] ;
 wire \usbfunction0.n2481_o[21] ;
 wire \usbfunction0.n2481_o[22] ;
 wire \usbfunction0.n2481_o[23] ;
 wire \usbfunction0.n2481_o[24] ;
 wire \usbfunction0.n2481_o[25] ;
 wire \usbfunction0.n2481_o[26] ;
 wire \usbfunction0.n2481_o[27] ;
 wire \usbfunction0.n2481_o[28] ;
 wire \usbfunction0.n2481_o[29] ;
 wire \usbfunction0.n2481_o[30] ;
 wire \usbfunction0.n2481_o[32] ;
 wire \usbfunction0.n2481_o[33] ;
 wire \usbfunction0.n2481_o[34] ;
 wire \usbfunction0.n2481_o[35] ;
 wire \usbfunction0.n2481_o[36] ;
 wire \usbfunction0.n2481_o[37] ;
 wire \usbfunction0.n2481_o[38] ;
 wire \usbfunction0.n2481_o[39] ;
 wire \usbfunction0.n2481_o[51] ;
 wire \usbfunction0.n2481_o[52] ;
 wire \usbfunction0.n2481_o[53] ;
 wire \usbfunction0.n2481_o[54] ;
 wire \usbfunction0.n2481_o[55] ;
 wire \usbfunction0.n2627_q ;
 wire \usbfunction0.n2628_q ;
 wire \usbfunction0.n2630_q ;
 wire \usbfunction0.n2631_q ;
 wire \usbfunction0.n2634_q[0] ;
 wire \usbfunction0.n2634_q[1] ;
 wire \usbfunction0.n2634_q[2] ;
 wire \usbfunction0.n2634_q[3] ;
 wire \usbfunction0.n2635_q[0] ;
 wire \usbfunction0.n2635_q[1] ;
 wire \usbfunction0.n2636_q ;
 wire \usbfunction0.n2637_q ;
 wire \usbfunction0.n2639_q ;
 wire \usbfunction0.n2640_q[0] ;
 wire \usbfunction0.n2640_q[1] ;
 wire \usbfunction0.n2640_q[2] ;
 wire \usbfunction0.n2640_q[3] ;
 wire \usbfunction0.n2642_q[0] ;
 wire \usbfunction0.n2642_q[1] ;
 wire \usbfunction0.n2642_q[2] ;
 wire \usbfunction0.n2642_q[3] ;
 wire \usbfunction0.n2644_q[0] ;
 wire \usbfunction0.n2644_q[10] ;
 wire \usbfunction0.n2644_q[11] ;
 wire \usbfunction0.n2644_q[12] ;
 wire \usbfunction0.n2644_q[13] ;
 wire \usbfunction0.n2644_q[14] ;
 wire \usbfunction0.n2644_q[15] ;
 wire \usbfunction0.n2644_q[1] ;
 wire \usbfunction0.n2644_q[2] ;
 wire \usbfunction0.n2644_q[3] ;
 wire \usbfunction0.n2644_q[4] ;
 wire \usbfunction0.n2644_q[5] ;
 wire \usbfunction0.n2644_q[6] ;
 wire \usbfunction0.n2644_q[7] ;
 wire \usbfunction0.n2644_q[8] ;
 wire \usbfunction0.n2644_q[9] ;
 wire \usbfunction0.n2645_q[2] ;
 wire \usbfunction0.n2648_q[0] ;
 wire \usbfunction0.n2648_q[10] ;
 wire \usbfunction0.n2648_q[11] ;
 wire \usbfunction0.n2648_q[12] ;
 wire \usbfunction0.n2648_q[13] ;
 wire \usbfunction0.n2648_q[14] ;
 wire \usbfunction0.n2648_q[15] ;
 wire \usbfunction0.n2648_q[1] ;
 wire \usbfunction0.n2648_q[2] ;
 wire \usbfunction0.n2648_q[3] ;
 wire \usbfunction0.n2648_q[4] ;
 wire \usbfunction0.n2648_q[5] ;
 wire \usbfunction0.n2648_q[6] ;
 wire \usbfunction0.n2648_q[7] ;
 wire \usbfunction0.n2648_q[8] ;
 wire \usbfunction0.n2648_q[9] ;
 wire \usbfunction0.n2649_q[0] ;
 wire \usbfunction0.n2649_q[1] ;
 wire \usbfunction0.n2649_q[2] ;
 wire \usbfunction0.n2649_q[3] ;
 wire \usbfunction0.n2649_q[4] ;
 wire \usbfunction0.n2649_q[5] ;
 wire \usbfunction0.n2649_q[6] ;
 wire \usbfunction0.n2649_q[7] ;
 wire \usbfunction0.n2650_q[0] ;
 wire \usbfunction0.n2650_q[1] ;
 wire \usbfunction0.n2650_q[2] ;
 wire \usbfunction0.n2650_q[3] ;
 wire \usbfunction0.n2650_q[4] ;
 wire \usbfunction0.n2650_q[5] ;
 wire \usbfunction0.n2650_q[6] ;
 wire \usbfunction0.n2650_q[7] ;
 wire \usbfunction0.n2651_q[0] ;
 wire \usbfunction0.n2651_q[1] ;
 wire \usbfunction0.n2651_q[2] ;
 wire \usbfunction0.n2651_q[3] ;
 wire \usbfunction0.n2651_q[4] ;
 wire \usbfunction0.n2651_q[5] ;
 wire \usbfunction0.n2651_q[6] ;
 wire \usbfunction0.n2651_q[7] ;
 wire \usbfunction0.n2652_q[0] ;
 wire \usbfunction0.n2652_q[1] ;
 wire \usbfunction0.n2652_q[2] ;
 wire \usbfunction0.n2652_q[3] ;
 wire \usbfunction0.n2652_q[4] ;
 wire \usbfunction0.n2652_q[5] ;
 wire \usbfunction0.n2652_q[6] ;
 wire \usbfunction0.n2652_q[7] ;
 wire \usbfunction0.n2653_q[0] ;
 wire \usbfunction0.n665_o[0] ;
 wire \usbfunction0.n665_o[1] ;
 wire \usbfunction0.n665_o[2] ;
 wire \usbfunction0.n665_o[3] ;
 wire \usbfunction0.n665_o[4] ;
 wire \usbfunction0.n665_o[5] ;
 wire \usbfunction0.n665_o[6] ;
 wire \usbfunction0.rxstream0.n6755_o ;
 wire \usbfunction0.s_m_descdata[0] ;
 wire \usbfunction0.s_m_descdata[1] ;
 wire \usbfunction0.s_m_descdata[2] ;
 wire \usbfunction0.s_m_descdata[3] ;
 wire \usbfunction0.s_m_descdata[4] ;
 wire \usbfunction0.s_m_descdata[5] ;
 wire \usbfunction0.s_m_descdata[6] ;
 wire \usbfunction0.s_m_descdata[7] ;
 wire \usbfunction0.s_m_rx_data[0] ;
 wire \usbfunction0.s_m_rx_data[1] ;
 wire \usbfunction0.s_m_rx_data[2] ;
 wire \usbfunction0.s_m_rx_data[3] ;
 wire \usbfunction0.s_m_rx_data[4] ;
 wire \usbfunction0.s_m_rx_data[5] ;
 wire \usbfunction0.s_m_rx_data[6] ;
 wire \usbfunction0.s_m_rx_data[7] ;
 wire \usbfunction0.s_m_rx_eop ;
 wire \usbfunction0.s_m_rx_error ;
 wire \usbfunction0.s_m_rx_sop ;
 wire \usbfunction0.s_m_rx_valid ;
 wire \usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8195_o[0] ;
 wire \usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8195_o[1] ;
 wire \usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8195_o[2] ;
 wire \usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8209_q[0] ;
 wire \usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8209_q[1] ;
 wire \usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8209_q[2] ;
 wire \usbfunction0.scl_usbgpiophy0.combinedbitcrc0.in_unnamed ;
 wire \usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[0] ;
 wire \usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[10] ;
 wire \usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[11] ;
 wire \usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[12] ;
 wire \usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[13] ;
 wire \usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[14] ;
 wire \usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[15] ;
 wire \usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[1] ;
 wire \usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[2] ;
 wire \usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[3] ;
 wire \usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[4] ;
 wire \usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[5] ;
 wire \usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[6] ;
 wire \usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[7] ;
 wire \usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[8] ;
 wire \usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[9] ;
 wire \usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.in_in_valid ;
 wire \usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7508_o ;
 wire \usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7634_o ;
 wire \usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7654_q[0] ;
 wire \usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7654_q[1] ;
 wire \usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7656_q ;
 wire \usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7657_q ;
 wire \usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.s_m_value[0] ;
 wire \usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.s_m_value[1] ;
 wire \usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.s_m_value[2] ;
 wire \usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.s_m_value[3] ;
 wire \usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.scl_counter0.n8128_o[0] ;
 wire \usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.scl_counter0.n8128_o[1] ;
 wire \usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.scl_counter0.n8128_o[2] ;
 wire \usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.scl_counter0.n8128_o[3] ;
 wire \usbfunction0.scl_usbgpiophy0.n6405_o ;
 wire \usbfunction0.scl_usbgpiophy0.n6411_o ;
 wire \usbfunction0.scl_usbgpiophy0.n6437_o ;
 wire \usbfunction0.scl_usbgpiophy0.n6449_o ;
 wire \usbfunction0.scl_usbgpiophy0.n6496_o ;
 wire \usbfunction0.scl_usbgpiophy0.n6500_o ;
 wire \usbfunction0.scl_usbgpiophy0.n6503_o ;
 wire \usbfunction0.scl_usbgpiophy0.n6529_o ;
 wire \usbfunction0.scl_usbgpiophy0.n6533_o ;
 wire \usbfunction0.scl_usbgpiophy0.n6553_o ;
 wire \usbfunction0.scl_usbgpiophy0.n6646_q ;
 wire \usbfunction0.scl_usbgpiophy0.n6649_q ;
 wire \usbfunction0.scl_usbgpiophy0.n6650_q ;
 wire \usbfunction0.scl_usbgpiophy0.n6651_q ;
 wire \usbfunction0.scl_usbgpiophy0.n6653_q ;
 wire \usbfunction0.scl_usbgpiophy0.n6654_q ;
 wire \usbfunction0.scl_usbgpiophy0.n6655_q ;
 wire \usbfunction0.scl_usbgpiophy0.nrzi0.n7721_q ;
 wire \usbfunction0.scl_usbgpiophy0.s_linein ;
 wire \usbfunction0.scl_usbgpiophy0.s_m_last ;
 wire \usbfunction0.scl_usbgpiophy0.s_out_2[0] ;
 wire \usbfunction0.scl_usbgpiophy0.s_out_2[1] ;
 wire \usbfunction0.scl_usbgpiophy0.s_out_2[2] ;
 wire \usbfunction0.scl_usbgpiophy0.s_out_2[3] ;
 wire \usbfunction0.scl_usbgpiophy0.s_out_2[4] ;
 wire \usbfunction0.scl_usbgpiophy0.s_out_2[5] ;
 wire \usbfunction0.scl_usbgpiophy0.s_out_2[6] ;
 wire \usbfunction0.scl_usbgpiophy0.s_out_2[7] ;
 wire \usbfunction0.scl_usbgpiophy0.s_ret_3 ;
 wire \usbfunction0.scl_usbgpiophy0.scl_addeopdeferred0.n7339_o ;
 wire \usbfunction0.scl_usbgpiophy0.scl_addeopdeferred0.n7349_q ;
 wire \usbfunction0.scl_usbgpiophy0.scl_addeopdeferred0.scl_eraselastbeat0.n8008_o ;
 wire \usbfunction0.scl_usbgpiophy0.scl_addeopdeferred0.scl_eraselastbeat0.n8041_q ;
 wire \usbfunction0.scl_usbgpiophy0.scl_addeopdeferred0.scl_eraselastbeat0.n8042_q ;
 wire \usbfunction0.scl_usbgpiophy0.scl_decodenrzi0.n7166_q ;
 wire \usbfunction0.scl_usbgpiophy0.scl_decodenrzi0.scl_counter0.n7944_q[0] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_decodenrzi0.scl_counter0.n7944_q[1] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_decodenrzi0.scl_counter0.n7944_q[2] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_extendwidth0.scl_counter0.n7961_o[0] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_extendwidth0.scl_counter0.n7961_o[1] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_extendwidth0.scl_counter0.n7961_o[2] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_extendwidth0.scl_counter0.n7984_q[0] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_extendwidth0.scl_counter0.n7984_q[1] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_extendwidth0.scl_counter0.n7984_q[2] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_insertbeat0.n7369_o ;
 wire \usbfunction0.scl_usbgpiophy0.scl_pulseextender0.n7741_o ;
 wire \usbfunction0.scl_usbgpiophy0.scl_pulseextender0.n7750_q ;
 wire \usbfunction0.scl_usbgpiophy0.scl_pulseextender0.scl_counter0.n8221_o[0] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_pulseextender0.scl_counter0.n8221_o[1] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_pulseextender0.scl_counter0.n8243_q[0] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_pulseextender0.scl_counter0.n8243_q[1] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_pulseextender1.n7766_o ;
 wire \usbfunction0.scl_usbgpiophy0.scl_pulseextender1.n7775_q ;
 wire \usbfunction0.scl_usbgpiophy0.scl_pulseextender1.scl_counter0.n8260_o[0] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_pulseextender1.scl_counter0.n8260_o[1] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_pulseextender1.scl_counter0.n8282_q[0] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_pulseextender1.scl_counter0.n8282_q[1] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_recoverdatadifferential0.scl_recoverdatadifferential_equalsampling_sky1300.detectsingleended0.n9022_q ;
 wire \usbfunction0.scl_usbgpiophy0.scl_recoverdatadifferential0.scl_recoverdatadifferential_equalsampling_sky1300.detectsingleended0.n9024_q ;
 wire \usbfunction0.scl_usbgpiophy0.scl_recoverdatadifferential0.scl_recoverdatadifferential_equalsampling_sky1300.detectsingleended0.n9025_q ;
 wire \usbfunction0.scl_usbgpiophy0.scl_recoverdatadifferential0.scl_recoverdatadifferential_equalsampling_sky1300.n7861_o ;
 wire \usbfunction0.scl_usbgpiophy0.scl_recoverdatadifferential0.scl_recoverdatadifferential_equalsampling_sky1300.n7883_q ;
 wire \usbfunction0.scl_usbgpiophy0.scl_reducewidth0.s_m_value[0] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_reducewidth0.s_m_value[1] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_reducewidth0.s_m_value[2] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_reducewidth0.scl_counter0.n8088_o[0] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_reducewidth0.scl_counter0.n8088_o[1] ;
 wire \usbfunction0.scl_usbgpiophy0.scl_reducewidth0.scl_counter0.n8088_o[2] ;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_leaf_0_clk_regs;
 wire clknet_leaf_1_clk_regs;
 wire clknet_leaf_2_clk_regs;
 wire clknet_leaf_3_clk_regs;
 wire clknet_leaf_4_clk_regs;
 wire clknet_leaf_5_clk_regs;
 wire clknet_leaf_6_clk_regs;
 wire clknet_leaf_7_clk_regs;
 wire clknet_leaf_8_clk_regs;
 wire clknet_leaf_9_clk_regs;
 wire clknet_leaf_10_clk_regs;
 wire clknet_leaf_11_clk_regs;
 wire clknet_leaf_12_clk_regs;
 wire clknet_leaf_13_clk_regs;
 wire clknet_leaf_14_clk_regs;
 wire clknet_leaf_15_clk_regs;
 wire clknet_leaf_16_clk_regs;
 wire clknet_leaf_17_clk_regs;
 wire clknet_leaf_18_clk_regs;
 wire clknet_leaf_19_clk_regs;
 wire clknet_leaf_20_clk_regs;
 wire clknet_leaf_21_clk_regs;
 wire clknet_leaf_22_clk_regs;
 wire clknet_leaf_23_clk_regs;
 wire clknet_leaf_24_clk_regs;
 wire clknet_leaf_25_clk_regs;
 wire clknet_leaf_26_clk_regs;
 wire clknet_leaf_27_clk_regs;
 wire clknet_leaf_28_clk_regs;
 wire clknet_leaf_29_clk_regs;
 wire clknet_leaf_30_clk_regs;
 wire clknet_leaf_31_clk_regs;
 wire clknet_leaf_32_clk_regs;
 wire clknet_leaf_33_clk_regs;
 wire clknet_leaf_34_clk_regs;
 wire clknet_leaf_35_clk_regs;
 wire clknet_leaf_36_clk_regs;
 wire clknet_leaf_37_clk_regs;
 wire clknet_leaf_38_clk_regs;
 wire clknet_leaf_39_clk_regs;
 wire clknet_leaf_40_clk_regs;
 wire clknet_leaf_41_clk_regs;
 wire clknet_leaf_42_clk_regs;
 wire clknet_leaf_43_clk_regs;
 wire clknet_leaf_44_clk_regs;
 wire clknet_leaf_45_clk_regs;
 wire clknet_leaf_46_clk_regs;
 wire clknet_leaf_47_clk_regs;
 wire clknet_leaf_48_clk_regs;
 wire clknet_leaf_49_clk_regs;
 wire clknet_leaf_50_clk_regs;
 wire clknet_leaf_51_clk_regs;
 wire clknet_leaf_52_clk_regs;
 wire clknet_leaf_53_clk_regs;
 wire clknet_leaf_54_clk_regs;
 wire clknet_leaf_55_clk_regs;
 wire clknet_leaf_56_clk_regs;
 wire clknet_leaf_57_clk_regs;
 wire clknet_leaf_58_clk_regs;
 wire clknet_leaf_59_clk_regs;
 wire clknet_leaf_60_clk_regs;
 wire clknet_leaf_61_clk_regs;
 wire clknet_leaf_62_clk_regs;
 wire clknet_leaf_63_clk_regs;
 wire clknet_leaf_64_clk_regs;
 wire clknet_leaf_65_clk_regs;
 wire clknet_leaf_66_clk_regs;
 wire clknet_leaf_67_clk_regs;
 wire clknet_leaf_68_clk_regs;
 wire clknet_leaf_69_clk_regs;
 wire clknet_leaf_70_clk_regs;
 wire clknet_leaf_71_clk_regs;
 wire clknet_leaf_72_clk_regs;
 wire clknet_leaf_73_clk_regs;
 wire clknet_leaf_74_clk_regs;
 wire clknet_leaf_75_clk_regs;
 wire clknet_leaf_76_clk_regs;
 wire clknet_leaf_77_clk_regs;
 wire clknet_leaf_78_clk_regs;
 wire clknet_leaf_79_clk_regs;
 wire clknet_leaf_80_clk_regs;
 wire clknet_leaf_81_clk_regs;
 wire clknet_leaf_82_clk_regs;
 wire clknet_leaf_83_clk_regs;
 wire clknet_leaf_84_clk_regs;
 wire clknet_leaf_85_clk_regs;
 wire clknet_leaf_86_clk_regs;
 wire clknet_leaf_87_clk_regs;
 wire clknet_leaf_88_clk_regs;
 wire clknet_leaf_89_clk_regs;
 wire clknet_leaf_90_clk_regs;
 wire clknet_leaf_91_clk_regs;
 wire clknet_leaf_92_clk_regs;
 wire clknet_leaf_93_clk_regs;
 wire clknet_leaf_94_clk_regs;
 wire clknet_leaf_95_clk_regs;
 wire clknet_leaf_96_clk_regs;
 wire clknet_leaf_97_clk_regs;
 wire clknet_leaf_98_clk_regs;
 wire clknet_leaf_99_clk_regs;
 wire clknet_leaf_100_clk_regs;
 wire clknet_leaf_101_clk_regs;
 wire clknet_leaf_102_clk_regs;
 wire clknet_leaf_103_clk_regs;
 wire clknet_leaf_104_clk_regs;
 wire clknet_leaf_105_clk_regs;
 wire clknet_leaf_106_clk_regs;
 wire clknet_leaf_107_clk_regs;
 wire clknet_leaf_108_clk_regs;
 wire clknet_leaf_109_clk_regs;
 wire clknet_leaf_110_clk_regs;
 wire clknet_leaf_111_clk_regs;
 wire clknet_leaf_112_clk_regs;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire clknet_5_0__leaf_clk_regs;
 wire clknet_5_1__leaf_clk_regs;
 wire clknet_5_2__leaf_clk_regs;
 wire clknet_5_3__leaf_clk_regs;
 wire clknet_5_4__leaf_clk_regs;
 wire clknet_5_5__leaf_clk_regs;
 wire clknet_5_6__leaf_clk_regs;
 wire clknet_5_7__leaf_clk_regs;
 wire clknet_5_8__leaf_clk_regs;
 wire clknet_5_9__leaf_clk_regs;
 wire clknet_5_10__leaf_clk_regs;
 wire clknet_5_11__leaf_clk_regs;
 wire clknet_5_12__leaf_clk_regs;
 wire clknet_5_13__leaf_clk_regs;
 wire clknet_5_14__leaf_clk_regs;
 wire clknet_5_15__leaf_clk_regs;
 wire clknet_5_16__leaf_clk_regs;
 wire clknet_5_17__leaf_clk_regs;
 wire clknet_5_18__leaf_clk_regs;
 wire clknet_5_19__leaf_clk_regs;
 wire clknet_5_20__leaf_clk_regs;
 wire clknet_5_21__leaf_clk_regs;
 wire clknet_5_22__leaf_clk_regs;
 wire clknet_5_23__leaf_clk_regs;
 wire clknet_5_24__leaf_clk_regs;
 wire clknet_5_25__leaf_clk_regs;
 wire clknet_5_26__leaf_clk_regs;
 wire clknet_5_27__leaf_clk_regs;
 wire clknet_5_28__leaf_clk_regs;
 wire clknet_5_29__leaf_clk_regs;
 wire clknet_5_30__leaf_clk_regs;
 wire clknet_5_31__leaf_clk_regs;
 wire delaynet_0_clk;
 wire delaynet_1_clk;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;

 sg13g2_inv_1 _4435_ (.Y(_0682_),
    .A(net1733));
 sg13g2_inv_1 _4436_ (.Y(_0683_),
    .A(\usbfunction0.n2313_o[1] ));
 sg13g2_inv_1 _4437_ (.Y(_0684_),
    .A(\usbfunction0.n2313_o[0] ));
 sg13g2_inv_1 _4438_ (.Y(_0685_),
    .A(net1124));
 sg13g2_inv_1 _4439_ (.Y(_0686_),
    .A(net1703));
 sg13g2_inv_1 _4440_ (.Y(_0687_),
    .A(net1872));
 sg13g2_inv_1 _4441_ (.Y(_0688_),
    .A(net1875));
 sg13g2_inv_1 _4442_ (.Y(_0689_),
    .A(net1735));
 sg13g2_inv_4 _4443_ (.A(net1504),
    .Y(_0690_));
 sg13g2_inv_1 _4444_ (.Y(_0691_),
    .A(net914));
 sg13g2_inv_4 _4445_ (.A(\scl_bitbangengine0.n3267_o ),
    .Y(_0692_));
 sg13g2_inv_1 _4446_ (.Y(_0693_),
    .A(net996));
 sg13g2_inv_2 _4447_ (.Y(_0694_),
    .A(\scl_bitbangengine0.n3258_o ));
 sg13g2_inv_2 _4448_ (.Y(_0695_),
    .A(net1798));
 sg13g2_inv_1 _4449_ (.Y(_0696_),
    .A(_0031_));
 sg13g2_inv_1 _4450_ (.Y(_0697_),
    .A(net1710));
 sg13g2_inv_1 _4451_ (.Y(_0698_),
    .A(_0032_));
 sg13g2_inv_1 _4452_ (.Y(_0699_),
    .A(\usbfunction0.n1583_o[4] ));
 sg13g2_inv_1 _4453_ (.Y(_0700_),
    .A(_0033_));
 sg13g2_inv_2 _4454_ (.Y(_0701_),
    .A(\usbfunction0.n2628_q ));
 sg13g2_inv_1 _4455_ (.Y(_0702_),
    .A(\usbfunction0.n2634_q[0] ));
 sg13g2_inv_2 _4456_ (.Y(_0703_),
    .A(net1649));
 sg13g2_inv_1 _4457_ (.Y(_0704_),
    .A(net1874));
 sg13g2_inv_2 _4458_ (.Y(_0705_),
    .A(net1477));
 sg13g2_inv_2 _4459_ (.Y(_0706_),
    .A(net1479));
 sg13g2_inv_1 _4460_ (.Y(_0707_),
    .A(n347_q));
 sg13g2_inv_1 _4461_ (.Y(_0708_),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[11] ));
 sg13g2_inv_1 _4462_ (.Y(_0709_),
    .A(net1588));
 sg13g2_inv_1 _4463_ (.Y(_0710_),
    .A(net687));
 sg13g2_inv_1 _4464_ (.Y(_0711_),
    .A(_0038_));
 sg13g2_inv_1 _4465_ (.Y(_0712_),
    .A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[1] ));
 sg13g2_inv_1 _4466_ (.Y(_0713_),
    .A(\usbfunction0.scl_usbgpiophy0.scl_insertbeat0.n7369_o ));
 sg13g2_inv_1 _4467_ (.Y(_0714_),
    .A(net832));
 sg13g2_inv_1 _4468_ (.Y(_0715_),
    .A(net1041));
 sg13g2_inv_1 _4469_ (.Y(_0716_),
    .A(net736));
 sg13g2_inv_1 _4470_ (.Y(_0717_),
    .A(net711));
 sg13g2_inv_1 _4471_ (.Y(_0718_),
    .A(s_m_popempty_2));
 sg13g2_inv_1 _4472_ (.Y(_0719_),
    .A(net1752));
 sg13g2_inv_1 _4473_ (.Y(_0720_),
    .A(\usbfunction0.n2650_q[7] ));
 sg13g2_inv_1 _4474_ (.Y(_0721_),
    .A(net984));
 sg13g2_inv_1 _4475_ (.Y(_0722_),
    .A(net1688));
 sg13g2_inv_2 _4476_ (.Y(_0723_),
    .A(\s_m_packetdata_2_rewired[0] ));
 sg13g2_inv_4 _4477_ (.A(n346_q),
    .Y(_0724_));
 sg13g2_inv_1 _4478_ (.Y(_0725_),
    .A(\scl_bitbangengine0.scl_counter0.n6975_q[0] ));
 sg13g2_inv_1 _4479_ (.Y(_0726_),
    .A(_0068_));
 sg13g2_inv_1 _4480_ (.Y(_0727_),
    .A(_0070_));
 sg13g2_inv_1 _4481_ (.Y(_0728_),
    .A(_0073_));
 sg13g2_inv_2 _4482_ (.Y(_0729_),
    .A(\scl_bitbangengine0.n3230_o ));
 sg13g2_inv_2 _4483_ (.Y(_0730_),
    .A(net1499));
 sg13g2_inv_2 _4484_ (.Y(_0731_),
    .A(net1498));
 sg13g2_inv_4 _4485_ (.A(net1492),
    .Y(_0732_));
 sg13g2_inv_1 _4486_ (.Y(_0733_),
    .A(net1801));
 sg13g2_inv_1 _4487_ (.Y(_0734_),
    .A(_0081_));
 sg13g2_inv_1 _4488_ (.Y(_0735_),
    .A(net1889));
 sg13g2_inv_1 _4489_ (.Y(_0736_),
    .A(net1774));
 sg13g2_inv_1 _4490_ (.Y(_0737_),
    .A(\scl_bitbangengine0.n5920_q[5] ));
 sg13g2_inv_1 _4491_ (.Y(_0738_),
    .A(net1151));
 sg13g2_inv_1 _4492_ (.Y(_0739_),
    .A(net1766));
 sg13g2_inv_1 _4493_ (.Y(_0740_),
    .A(net1584));
 sg13g2_inv_1 _4494_ (.Y(_0741_),
    .A(net881));
 sg13g2_inv_1 _4495_ (.Y(_0742_),
    .A(net1571));
 sg13g2_inv_1 _4496_ (.Y(_0743_),
    .A(net1577));
 sg13g2_inv_1 _4497_ (.Y(_0744_),
    .A(net1646));
 sg13g2_inv_1 _4498_ (.Y(_0745_),
    .A(net1054));
 sg13g2_inv_1 _4499_ (.Y(_0746_),
    .A(net734));
 sg13g2_inv_1 _4500_ (.Y(_0747_),
    .A(net683));
 sg13g2_inv_1 _4501_ (.Y(_0748_),
    .A(net878));
 sg13g2_inv_1 _4502_ (.Y(_0749_),
    .A(net896));
 sg13g2_inv_1 _4503_ (.Y(_0750_),
    .A(net1056));
 sg13g2_inv_1 _4504_ (.Y(_0751_),
    .A(net1003));
 sg13g2_inv_1 _4505_ (.Y(_0752_),
    .A(net1033));
 sg13g2_inv_1 _4506_ (.Y(_0753_),
    .A(net971));
 sg13g2_inv_1 _4507_ (.Y(_0754_),
    .A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[6] ));
 sg13g2_inv_1 _4508_ (.Y(_0755_),
    .A(net797));
 sg13g2_inv_1 _4509_ (.Y(_0756_),
    .A(net1163));
 sg13g2_inv_1 _4510_ (.Y(_0757_),
    .A(net1000));
 sg13g2_inv_1 _4511_ (.Y(_0758_),
    .A(net1060));
 sg13g2_inv_1 _4512_ (.Y(_0759_),
    .A(net870));
 sg13g2_inv_1 _4513_ (.Y(_0760_),
    .A(net1865));
 sg13g2_inv_1 _4514_ (.Y(_0761_),
    .A(\usbfunction0.n2652_q[6] ));
 sg13g2_inv_1 _4515_ (.Y(_0762_),
    .A(net1771));
 sg13g2_inv_1 _4516_ (.Y(_0763_),
    .A(net1709));
 sg13g2_inv_1 _4517_ (.Y(_0764_),
    .A(_0095_));
 sg13g2_inv_1 _4518_ (.Y(_0765_),
    .A(\usbfunction0.n2651_q[3] ));
 sg13g2_inv_1 _4519_ (.Y(_0766_),
    .A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[11] ));
 sg13g2_inv_1 _4520_ (.Y(_0767_),
    .A(net992));
 sg13g2_inv_1 _4521_ (.Y(_0768_),
    .A(net924));
 sg13g2_inv_1 _4522_ (.Y(_0769_),
    .A(net1058));
 sg13g2_inv_1 _4523_ (.Y(_0770_),
    .A(_0132_));
 sg13g2_inv_1 _4524_ (.Y(_0771_),
    .A(net1116));
 sg13g2_inv_2 _4525_ (.Y(_0772_),
    .A(\scl_bitbangengine0.n5915_q ));
 sg13g2_inv_1 _4526_ (.Y(_0773_),
    .A(\scl_bitbangengine0.n5423_o[6] ));
 sg13g2_inv_1 _4527_ (.Y(_0774_),
    .A(net1621));
 sg13g2_inv_1 _4528_ (.Y(_0775_),
    .A(net765));
 sg13g2_inv_1 _4529_ (.Y(_0776_),
    .A(net546));
 sg13g2_inv_1 _7831__2 (.Y(net529),
    .A(clknet_1_0__leaf_clk));
 sg13g2_nor4_1 _4531_ (.A(net1744),
    .B(net1090),
    .C(\usbfunction0.scl_usbgpiophy0.scl_recoverdatadifferential0.scl_recoverdatadifferential_equalsampling_sky1300.detectsingleended0.n9024_q ),
    .D(\usbfunction0.scl_usbgpiophy0.scl_recoverdatadifferential0.scl_recoverdatadifferential_equalsampling_sky1300.detectsingleended0.n9025_q ),
    .Y(\usbfunction0.scl_usbgpiophy0.scl_recoverdatadifferential0.scl_recoverdatadifferential_equalsampling_sky1300.n7861_o ));
 sg13g2_nor2_1 _4532_ (.A(net1006),
    .B(net1437),
    .Y(_0777_));
 sg13g2_nand2_1 _4533_ (.Y(_0778_),
    .A(\usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8209_q[1] ),
    .B(net588));
 sg13g2_or2_1 _4534_ (.X(_0779_),
    .B(_0778_),
    .A(\usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8209_q[0] ));
 sg13g2_nand2b_2 _4535_ (.Y(_0780_),
    .B(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7654_q[1] ),
    .A_N(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7654_q[0] ));
 sg13g2_nand3_1 _4536_ (.B(_0779_),
    .C(_0780_),
    .A(_0043_),
    .Y(_0781_));
 sg13g2_and2_2 _4537_ (.A(_0777_),
    .B(_0781_),
    .X(_0782_));
 sg13g2_nor2_1 _4538_ (.A(\usbfunction0.scl_usbgpiophy0.n6655_q ),
    .B(_0782_),
    .Y(_0783_));
 sg13g2_inv_2 _4539_ (.Y(\usbfunction0.scl_usbgpiophy0.n6496_o ),
    .A(_0783_));
 sg13g2_nand2_2 _4540_ (.Y(_0784_),
    .A(net1619),
    .B(_0783_));
 sg13g2_nand2b_1 _4541_ (.Y(_0785_),
    .B(\usbfunction0.scl_usbgpiophy0.scl_decodenrzi0.scl_counter0.n7944_q[1] ),
    .A_N(_0044_));
 sg13g2_nor2_1 _4542_ (.A(\usbfunction0.scl_usbgpiophy0.scl_decodenrzi0.scl_counter0.n7944_q[0] ),
    .B(_0785_),
    .Y(_0786_));
 sg13g2_nor2_1 _4543_ (.A(net1398),
    .B(_0786_),
    .Y(_0787_));
 sg13g2_nor2_1 _4544_ (.A(\usbfunction0.scl_usbgpiophy0.scl_decodenrzi0.n7166_q ),
    .B(_0784_),
    .Y(_0788_));
 sg13g2_xnor2_1 _4545_ (.Y(_0789_),
    .A(\usbfunction0.scl_usbgpiophy0.s_linein ),
    .B(_0788_));
 sg13g2_inv_1 _4546_ (.Y(\usbfunction0.s_m_rx_data[7] ),
    .A(_0789_));
 sg13g2_and2_1 _4547_ (.A(net1386),
    .B(_0789_),
    .X(_0790_));
 sg13g2_nand2_1 _4548_ (.Y(_0791_),
    .A(net559),
    .B(_0790_));
 sg13g2_nor2_1 _4549_ (.A(_0786_),
    .B(_0789_),
    .Y(_0792_));
 sg13g2_nor3_2 _4550_ (.A(net1398),
    .B(_0786_),
    .C(_0789_),
    .Y(_0793_));
 sg13g2_nand2_1 _4551_ (.Y(_0794_),
    .A(net1170),
    .B(_0793_));
 sg13g2_nand3_1 _4552_ (.B(net1670),
    .C(net1386),
    .A(net1023),
    .Y(_0795_));
 sg13g2_nor2_1 _4553_ (.A(\usbfunction0.scl_usbgpiophy0.n6437_o ),
    .B(net1436),
    .Y(_0796_));
 sg13g2_nand2b_1 _4554_ (.Y(_0797_),
    .B(net1386),
    .A_N(_0796_));
 sg13g2_nand3_1 _4555_ (.B(_0795_),
    .C(_0797_),
    .A(_0794_),
    .Y(_0798_));
 sg13g2_nor2b_1 _4556_ (.A(_0798_),
    .B_N(_0791_),
    .Y(_0799_));
 sg13g2_nand2_1 _4557_ (.Y(_0800_),
    .A(\usbfunction0.scl_usbgpiophy0.n6437_o ),
    .B(_0793_));
 sg13g2_nor2_1 _4558_ (.A(\usbfunction0.scl_usbgpiophy0.n6449_o ),
    .B(_0800_),
    .Y(_0801_));
 sg13g2_a221oi_1 _4559_ (.B2(net559),
    .C1(_0801_),
    .B1(_0799_),
    .A1(net1436),
    .Y(_0184_),
    .A2(net1386));
 sg13g2_nor2b_2 _4560_ (.A(net11),
    .B_N(net552),
    .Y(_0802_));
 sg13g2_and2_1 _4561_ (.A(net598),
    .B(_0802_),
    .X(_0803_));
 sg13g2_nand2_2 _4562_ (.Y(_0804_),
    .A(net598),
    .B(_0802_));
 sg13g2_nor2_1 _4563_ (.A(\usbfunction0.n2634_q[3] ),
    .B(\usbfunction0.n2634_q[2] ),
    .Y(_0805_));
 sg13g2_or2_1 _4564_ (.X(_0806_),
    .B(\usbfunction0.n2634_q[2] ),
    .A(\usbfunction0.n2634_q[3] ));
 sg13g2_nand3b_1 _4565_ (.B(\usbfunction0.n2634_q[0] ),
    .C(\usbfunction0.n2634_q[1] ),
    .Y(_0807_),
    .A_N(_0036_));
 sg13g2_nor2_1 _4566_ (.A(_0806_),
    .B(_0807_),
    .Y(_0808_));
 sg13g2_nand3_1 _4567_ (.B(\usbfunction0.n1581_o[0] ),
    .C(_0035_),
    .A(\usbfunction0.n1581_o[1] ),
    .Y(_0809_));
 sg13g2_nor3_1 _4568_ (.A(_0806_),
    .B(_0807_),
    .C(_0809_),
    .Y(_0810_));
 sg13g2_or4_2 _4569_ (.A(_0707_),
    .B(_0806_),
    .C(_0807_),
    .D(_0809_),
    .X(_0811_));
 sg13g2_inv_2 _4570_ (.Y(_0812_),
    .A(net1429));
 sg13g2_mux2_2 _4571_ (.A0(net1617),
    .A1(net1869),
    .S(net1429),
    .X(\n352_o[22] ));
 sg13g2_nor2_1 _4572_ (.A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[15] ),
    .B(\n352_o[22] ),
    .Y(_0813_));
 sg13g2_mux2_2 _4573_ (.A0(net1595),
    .A1(net1871),
    .S(net1429),
    .X(\n352_o[21] ));
 sg13g2_nand2_1 _4574_ (.Y(_0814_),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[14] ),
    .B(\n352_o[21] ));
 sg13g2_xor2_1 _4575_ (.B(\n352_o[21] ),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[14] ),
    .X(_0815_));
 sg13g2_mux2_2 _4576_ (.A0(\s_m_packetdata_2_rewired[18] ),
    .A1(net1804),
    .S(net1433),
    .X(\n352_o[18] ));
 sg13g2_inv_1 _4577_ (.Y(_0816_),
    .A(\n352_o[18] ));
 sg13g2_nor2_1 _4578_ (.A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[11] ),
    .B(\n352_o[18] ),
    .Y(_0817_));
 sg13g2_mux2_2 _4579_ (.A0(net1904),
    .A1(net1610),
    .S(net1429),
    .X(_0818_));
 sg13g2_inv_1 _4580_ (.Y(_0182_),
    .A(_0818_));
 sg13g2_nor2_1 _4581_ (.A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[9] ),
    .B(_0818_),
    .Y(_0819_));
 sg13g2_mux2_2 _4582_ (.A0(\s_m_packetdata_2_rewired[15] ),
    .A1(net1074),
    .S(net1433),
    .X(_0820_));
 sg13g2_inv_1 _4583_ (.Y(_0181_),
    .A(net1075));
 sg13g2_and2_1 _4584_ (.A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[8] ),
    .B(_0820_),
    .X(_0821_));
 sg13g2_mux2_2 _4585_ (.A0(net1161),
    .A1(net1660),
    .S(net1432),
    .X(_0822_));
 sg13g2_inv_1 _4586_ (.Y(_0180_),
    .A(_0822_));
 sg13g2_and2_1 _4587_ (.A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[7] ),
    .B(_0822_),
    .X(_0823_));
 sg13g2_mux2_2 _4588_ (.A0(net1696),
    .A1(net1816),
    .S(net1432),
    .X(\n352_o[13] ));
 sg13g2_nand2_1 _4589_ (.Y(_0824_),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[6] ),
    .B(\n352_o[13] ));
 sg13g2_mux2_2 _4590_ (.A0(net1739),
    .A1(net1852),
    .S(net1430),
    .X(\n352_o[12] ));
 sg13g2_and2_1 _4591_ (.A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[5] ),
    .B(\n352_o[12] ),
    .X(_0825_));
 sg13g2_mux2_2 _4592_ (.A0(\s_m_packetdata_2_rewired[11] ),
    .A1(net1859),
    .S(net1430),
    .X(\n352_o[11] ));
 sg13g2_nand2_1 _4593_ (.Y(_0826_),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[4] ),
    .B(\n352_o[11] ));
 sg13g2_mux2_2 _4594_ (.A0(net1794),
    .A1(net1835),
    .S(net1430),
    .X(\n352_o[10] ));
 sg13g2_and2_1 _4595_ (.A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[3] ),
    .B(\n352_o[10] ),
    .X(_0827_));
 sg13g2_mux2_2 _4596_ (.A0(\s_m_packetdata_2_rewired[9] ),
    .A1(net1137),
    .S(net1432),
    .X(_0828_));
 sg13g2_inv_1 _4597_ (.Y(_0179_),
    .A(net1138));
 sg13g2_and2_1 _4598_ (.A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[2] ),
    .B(_0828_),
    .X(_0829_));
 sg13g2_mux2_2 _4599_ (.A0(net1487),
    .A1(net1792),
    .S(net1432),
    .X(\n352_o[8] ));
 sg13g2_nand2_1 _4600_ (.Y(_0830_),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[1] ),
    .B(\n352_o[8] ));
 sg13g2_mux2_2 _4601_ (.A0(net1627),
    .A1(net1810),
    .S(net1431),
    .X(\n352_o[7] ));
 sg13g2_nand2_1 _4602_ (.Y(_0831_),
    .A(_0709_),
    .B(\n352_o[7] ));
 sg13g2_xnor2_1 _4603_ (.Y(_0832_),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[1] ),
    .B(\n352_o[8] ));
 sg13g2_o21ai_1 _4604_ (.B1(_0830_),
    .Y(_0833_),
    .A1(_0831_),
    .A2(_0832_));
 sg13g2_xor2_1 _4605_ (.B(_0828_),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[2] ),
    .X(_0834_));
 sg13g2_a21o_1 _4606_ (.A2(_0834_),
    .A1(_0833_),
    .B1(_0829_),
    .X(_0835_));
 sg13g2_xor2_1 _4607_ (.B(\n352_o[10] ),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[3] ),
    .X(_0836_));
 sg13g2_a21oi_1 _4608_ (.A1(_0835_),
    .A2(_0836_),
    .Y(_0837_),
    .B1(_0827_));
 sg13g2_nor2_1 _4609_ (.A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[4] ),
    .B(\n352_o[11] ),
    .Y(_0838_));
 sg13g2_xor2_1 _4610_ (.B(\n352_o[11] ),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[4] ),
    .X(_0839_));
 sg13g2_o21ai_1 _4611_ (.B1(_0826_),
    .Y(_0840_),
    .A1(_0837_),
    .A2(_0838_));
 sg13g2_xor2_1 _4612_ (.B(\n352_o[12] ),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[5] ),
    .X(_0841_));
 sg13g2_a21oi_1 _4613_ (.A1(_0840_),
    .A2(_0841_),
    .Y(_0842_),
    .B1(_0825_));
 sg13g2_nor2_1 _4614_ (.A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[6] ),
    .B(\n352_o[13] ),
    .Y(_0843_));
 sg13g2_xor2_1 _4615_ (.B(\n352_o[13] ),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[6] ),
    .X(_0844_));
 sg13g2_o21ai_1 _4616_ (.B1(_0824_),
    .Y(_0845_),
    .A1(_0842_),
    .A2(_0843_));
 sg13g2_xor2_1 _4617_ (.B(_0822_),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[7] ),
    .X(_0846_));
 sg13g2_a21o_1 _4618_ (.A2(_0846_),
    .A1(_0845_),
    .B1(_0823_),
    .X(_0847_));
 sg13g2_xor2_1 _4619_ (.B(_0820_),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[8] ),
    .X(_0848_));
 sg13g2_a21o_1 _4620_ (.A2(_0848_),
    .A1(_0847_),
    .B1(_0821_),
    .X(_0849_));
 sg13g2_a221oi_1 _4621_ (.B2(_0848_),
    .C1(_0821_),
    .B1(_0847_),
    .A1(\scl_uartrx0.scl_baudrategenerator0.n7047_o[9] ),
    .Y(_0850_),
    .A2(_0818_));
 sg13g2_mux2_2 _4622_ (.A0(s_m_packetdata_2_bit_17),
    .A1(net1775),
    .S(net1429),
    .X(\n352_o[17] ));
 sg13g2_nand2_1 _4623_ (.Y(_0851_),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[10] ),
    .B(\n352_o[17] ));
 sg13g2_inv_1 _4624_ (.Y(_0852_),
    .A(_0851_));
 sg13g2_xnor2_1 _4625_ (.Y(_0853_),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[10] ),
    .B(\n352_o[17] ));
 sg13g2_nor3_1 _4626_ (.A(_0819_),
    .B(_0850_),
    .C(_0853_),
    .Y(_0854_));
 sg13g2_or3_2 _4627_ (.A(_0819_),
    .B(_0850_),
    .C(_0853_),
    .X(_0855_));
 sg13g2_nand2_1 _4628_ (.Y(_0856_),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[11] ),
    .B(\n352_o[18] ));
 sg13g2_and2_1 _4629_ (.A(_0851_),
    .B(_0856_),
    .X(_0857_));
 sg13g2_nor2b_1 _4630_ (.A(_0817_),
    .B_N(_0856_),
    .Y(_0858_));
 sg13g2_a21oi_1 _4631_ (.A1(_0855_),
    .A2(_0857_),
    .Y(_0859_),
    .B1(_0817_));
 sg13g2_mux2_2 _4632_ (.A0(\s_m_packetdata_2_rewired[19] ),
    .A1(net1793),
    .S(net1429),
    .X(\n352_o[19] ));
 sg13g2_and2_1 _4633_ (.A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[12] ),
    .B(\n352_o[19] ),
    .X(_0860_));
 sg13g2_xor2_1 _4634_ (.B(\n352_o[19] ),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[12] ),
    .X(_0861_));
 sg13g2_inv_1 _4635_ (.Y(_0862_),
    .A(_0861_));
 sg13g2_mux2_2 _4636_ (.A0(net1759),
    .A1(net1829),
    .S(net1429),
    .X(\n352_o[20] ));
 sg13g2_nand2_1 _4637_ (.Y(_0863_),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[13] ),
    .B(\n352_o[20] ));
 sg13g2_xnor2_1 _4638_ (.Y(_0864_),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[13] ),
    .B(\n352_o[20] ));
 sg13g2_or2_1 _4639_ (.X(_0865_),
    .B(_0864_),
    .A(_0862_));
 sg13g2_a221oi_1 _4640_ (.B2(_0857_),
    .C1(_0865_),
    .B1(_0855_),
    .A1(_0708_),
    .Y(_0866_),
    .A2(_0816_));
 sg13g2_o21ai_1 _4641_ (.B1(_0860_),
    .Y(_0867_),
    .A1(\scl_uartrx0.scl_baudrategenerator0.n7047_o[13] ),
    .A2(\n352_o[20] ));
 sg13g2_nand2_1 _4642_ (.Y(_0868_),
    .A(_0863_),
    .B(_0867_));
 sg13g2_o21ai_1 _4643_ (.B1(_0815_),
    .Y(_0869_),
    .A1(_0866_),
    .A2(_0868_));
 sg13g2_a22oi_1 _4644_ (.Y(_0870_),
    .B1(\n352_o[21] ),
    .B2(\scl_uartrx0.scl_baudrategenerator0.n7047_o[14] ),
    .A2(\n352_o[22] ),
    .A1(\scl_uartrx0.scl_baudrategenerator0.n7047_o[15] ));
 sg13g2_a21oi_2 _4645_ (.B1(_0813_),
    .Y(_0871_),
    .A2(_0870_),
    .A1(_0869_));
 sg13g2_mux2_2 _4646_ (.A0(net1565),
    .A1(net1857),
    .S(net1429),
    .X(\n352_o[23] ));
 sg13g2_and2_1 _4647_ (.A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[16] ),
    .B(\n352_o[23] ),
    .X(_0872_));
 sg13g2_xor2_1 _4648_ (.B(\n352_o[23] ),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[16] ),
    .X(_0873_));
 sg13g2_xnor2_1 _4649_ (.Y(_0874_),
    .A(_0871_),
    .B(_0873_));
 sg13g2_inv_1 _4650_ (.Y(_0875_),
    .A(_0874_));
 sg13g2_or3_1 _4651_ (.A(_0815_),
    .B(_0866_),
    .C(_0868_),
    .X(_0876_));
 sg13g2_and2_1 _4652_ (.A(_0869_),
    .B(_0876_),
    .X(_0877_));
 sg13g2_a221oi_1 _4653_ (.B2(_0857_),
    .C1(_0862_),
    .B1(_0855_),
    .A1(_0708_),
    .Y(_0878_),
    .A2(_0816_));
 sg13g2_xnor2_1 _4654_ (.Y(_0879_),
    .A(_0859_),
    .B(_0861_));
 sg13g2_nor3_1 _4655_ (.A(_0852_),
    .B(_0854_),
    .C(_0858_),
    .Y(_0880_));
 sg13g2_o21ai_1 _4656_ (.B1(_0858_),
    .Y(_0881_),
    .A1(_0852_),
    .A2(_0854_));
 sg13g2_nand2b_1 _4657_ (.Y(_0882_),
    .B(_0881_),
    .A_N(_0880_));
 sg13g2_xor2_1 _4658_ (.B(_0848_),
    .A(_0847_),
    .X(_0883_));
 sg13g2_xnor2_1 _4659_ (.Y(_0884_),
    .A(_0845_),
    .B(_0846_));
 sg13g2_xnor2_1 _4660_ (.Y(_0885_),
    .A(_0840_),
    .B(_0841_));
 sg13g2_xnor2_1 _4661_ (.Y(_0886_),
    .A(_0837_),
    .B(_0839_));
 sg13g2_xnor2_1 _4662_ (.Y(_0887_),
    .A(_0833_),
    .B(_0834_));
 sg13g2_xnor2_1 _4663_ (.Y(_0888_),
    .A(_0831_),
    .B(_0832_));
 sg13g2_nor2_1 _4664_ (.A(_0887_),
    .B(_0888_),
    .Y(_0889_));
 sg13g2_xor2_1 _4665_ (.B(_0836_),
    .A(_0835_),
    .X(_0890_));
 sg13g2_nor2_1 _4666_ (.A(_0889_),
    .B(_0890_),
    .Y(_0891_));
 sg13g2_nor2b_1 _4667_ (.A(_0891_),
    .B_N(_0886_),
    .Y(_0892_));
 sg13g2_nor2b_1 _4668_ (.A(_0885_),
    .B_N(_0892_),
    .Y(_0893_));
 sg13g2_xnor2_1 _4669_ (.Y(_0894_),
    .A(_0842_),
    .B(_0844_));
 sg13g2_nor2_1 _4670_ (.A(_0893_),
    .B(_0894_),
    .Y(_0895_));
 sg13g2_and2_1 _4671_ (.A(_0884_),
    .B(_0895_),
    .X(_0896_));
 sg13g2_nand2b_1 _4672_ (.Y(_0897_),
    .B(_0896_),
    .A_N(_0883_));
 sg13g2_xnor2_1 _4673_ (.Y(_0898_),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[9] ),
    .B(_0818_));
 sg13g2_xnor2_1 _4674_ (.Y(_0899_),
    .A(_0849_),
    .B(_0898_));
 sg13g2_o21ai_1 _4675_ (.B1(_0853_),
    .Y(_0900_),
    .A1(_0819_),
    .A2(_0850_));
 sg13g2_and4_1 _4676_ (.A(_0855_),
    .B(_0897_),
    .C(_0899_),
    .D(_0900_),
    .X(_0901_));
 sg13g2_nor2b_1 _4677_ (.A(_0882_),
    .B_N(_0901_),
    .Y(_0902_));
 sg13g2_nand3b_1 _4678_ (.B(_0881_),
    .C(_0901_),
    .Y(_0903_),
    .A_N(_0880_));
 sg13g2_nand2_1 _4679_ (.Y(_0904_),
    .A(_0879_),
    .B(_0903_));
 sg13g2_o21ai_1 _4680_ (.B1(_0864_),
    .Y(_0905_),
    .A1(_0860_),
    .A2(_0878_));
 sg13g2_or3_1 _4681_ (.A(_0860_),
    .B(_0864_),
    .C(_0878_),
    .X(_0906_));
 sg13g2_nand2_1 _4682_ (.Y(_0907_),
    .A(_0905_),
    .B(_0906_));
 sg13g2_a22oi_1 _4683_ (.Y(_0908_),
    .B1(_0905_),
    .B2(_0906_),
    .A2(_0903_),
    .A1(_0879_));
 sg13g2_nand2_1 _4684_ (.Y(_0909_),
    .A(_0877_),
    .B(_0908_));
 sg13g2_xnor2_1 _4685_ (.Y(_0910_),
    .A(\scl_uartrx0.scl_baudrategenerator0.n7047_o[15] ),
    .B(\n352_o[22] ));
 sg13g2_nand3_1 _4686_ (.B(_0869_),
    .C(_0910_),
    .A(_0814_),
    .Y(_0911_));
 sg13g2_a21o_1 _4687_ (.A2(_0869_),
    .A1(_0814_),
    .B1(_0910_),
    .X(_0912_));
 sg13g2_nand2_1 _4688_ (.Y(_0913_),
    .A(_0911_),
    .B(_0912_));
 sg13g2_a22oi_1 _4689_ (.Y(_0914_),
    .B1(_0911_),
    .B2(_0912_),
    .A2(_0908_),
    .A1(_0877_));
 sg13g2_nand2_1 _4690_ (.Y(_0915_),
    .A(_0909_),
    .B(_0913_));
 sg13g2_nor2_1 _4691_ (.A(_0874_),
    .B(_0914_),
    .Y(_0916_));
 sg13g2_a21oi_1 _4692_ (.A1(_0871_),
    .A2(_0873_),
    .Y(_0917_),
    .B1(_0872_));
 sg13g2_a21o_1 _4693_ (.A2(_0873_),
    .A1(_0871_),
    .B1(_0872_),
    .X(_0918_));
 sg13g2_nor2_1 _4694_ (.A(_0916_),
    .B(_0918_),
    .Y(_0919_));
 sg13g2_o21ai_1 _4695_ (.B1(_0917_),
    .Y(_0920_),
    .A1(_0874_),
    .A2(_0914_));
 sg13g2_and3_1 _4696_ (.X(_0921_),
    .A(net11),
    .B(net938),
    .C(net1260));
 sg13g2_and2_2 _4697_ (.A(_0804_),
    .B(net1259),
    .X(_0922_));
 sg13g2_and2_1 _4698_ (.A(net878),
    .B(_0922_),
    .X(_0923_));
 sg13g2_nor3_1 _4699_ (.A(_0690_),
    .B(_0748_),
    .C(net1241),
    .Y(_0924_));
 sg13g2_and2_2 _4700_ (.A(net1842),
    .B(net1434),
    .X(_0925_));
 sg13g2_and2_2 _4701_ (.A(net1260),
    .B(_0925_),
    .X(_0926_));
 sg13g2_nand2_2 _4702_ (.Y(_0927_),
    .A(net1260),
    .B(_0925_));
 sg13g2_and2_1 _4703_ (.A(net1461),
    .B(\scl_uartrx0.s_m_value[0] ),
    .X(_0928_));
 sg13g2_nand3_1 _4704_ (.B(_0926_),
    .C(_0928_),
    .A(net1567),
    .Y(_0929_));
 sg13g2_inv_2 _4705_ (.Y(\scl_uartrx0.n6047_o ),
    .A(_0929_));
 sg13g2_or3_1 _4706_ (.A(_0921_),
    .B(_0923_),
    .C(\scl_uartrx0.n6047_o ),
    .X(_0930_));
 sg13g2_nor2_1 _4707_ (.A(net1435),
    .B(_0930_),
    .Y(_0931_));
 sg13g2_nor2_1 _4708_ (.A(_0921_),
    .B(_0929_),
    .Y(_0932_));
 sg13g2_a221oi_1 _4709_ (.B2(net552),
    .C1(_0921_),
    .B1(_0931_),
    .A1(_0924_),
    .Y(_0183_),
    .A2(_0929_));
 sg13g2_nand2b_1 _4710_ (.Y(_0933_),
    .B(net1473),
    .A_N(net1470));
 sg13g2_nand2_1 _4711_ (.Y(_0934_),
    .A(net1467),
    .B(net1464));
 sg13g2_nand2b_2 _4712_ (.Y(_0935_),
    .B(\s_m_pushdata_data[1] ),
    .A_N(net1476));
 sg13g2_or2_1 _4713_ (.X(_0936_),
    .B(\s_m_pushdata_data[0] ),
    .A(\s_m_pushdata_data[3] ));
 sg13g2_nor4_2 _4714_ (.A(_0933_),
    .B(_0934_),
    .C(_0935_),
    .Y(_0937_),
    .D(_0936_));
 sg13g2_or4_2 _4715_ (.A(_0933_),
    .B(_0934_),
    .C(_0935_),
    .D(_0936_),
    .X(_0938_));
 sg13g2_nand2_1 _4716_ (.Y(_0939_),
    .A(net912),
    .B(\usbfunction0.n2630_q ));
 sg13g2_nor2_2 _4717_ (.A(_0029_),
    .B(_0939_),
    .Y(_0940_));
 sg13g2_or2_1 _4718_ (.X(_0941_),
    .B(_0939_),
    .A(_0029_));
 sg13g2_nor2_1 _4719_ (.A(net1428),
    .B(net1426),
    .Y(_0942_));
 sg13g2_nand2_1 _4720_ (.Y(_0943_),
    .A(_0937_),
    .B(net1427));
 sg13g2_nor2b_1 _4721_ (.A(net1489),
    .B_N(net1883),
    .Y(_0944_));
 sg13g2_o21ai_1 _4722_ (.B1(_0944_),
    .Y(_0945_),
    .A1(_0938_),
    .A2(_0941_));
 sg13g2_nor2b_2 _4723_ (.A(net1490),
    .B_N(net1843),
    .Y(_0946_));
 sg13g2_nand3_1 _4724_ (.B(_0940_),
    .C(_0946_),
    .A(_0937_),
    .Y(_0947_));
 sg13g2_nand2_1 _4725_ (.Y(\usbfunction0.n665_o[3] ),
    .A(_0945_),
    .B(_0947_));
 sg13g2_nand3_1 _4726_ (.B(_0945_),
    .C(_0947_),
    .A(_0032_),
    .Y(_0948_));
 sg13g2_a21o_1 _4727_ (.A2(_0947_),
    .A1(_0945_),
    .B1(_0032_),
    .X(_0949_));
 sg13g2_nor2_1 _4728_ (.A(\usbfunction0.n2634_q[1] ),
    .B(\usbfunction0.n2634_q[0] ),
    .Y(_0950_));
 sg13g2_nor2b_1 _4729_ (.A(\usbfunction0.n2627_q ),
    .B_N(\usbfunction0.n1581_o[0] ),
    .Y(_0951_));
 sg13g2_o21ai_1 _4730_ (.B1(_0951_),
    .Y(_0952_),
    .A1(\usbfunction0.n1359_o[1] ),
    .A2(_0686_));
 sg13g2_nor4_1 _4731_ (.A(\usbfunction0.n1581_o[1] ),
    .B(\usbfunction0.n2634_q[1] ),
    .C(\usbfunction0.n2634_q[0] ),
    .D(_0952_),
    .Y(_0953_));
 sg13g2_nand3_1 _4732_ (.B(_0805_),
    .C(_0953_),
    .A(\usbfunction0.n2628_q ),
    .Y(_0954_));
 sg13g2_nor2b_1 _4733_ (.A(net1489),
    .B_N(net1885),
    .Y(_0955_));
 sg13g2_o21ai_1 _4734_ (.B1(_0955_),
    .Y(_0956_),
    .A1(net1428),
    .A2(net1426));
 sg13g2_nor2b_1 _4735_ (.A(net1490),
    .B_N(net1809),
    .Y(_0957_));
 sg13g2_nand3_1 _4736_ (.B(net1427),
    .C(_0957_),
    .A(_0937_),
    .Y(_0958_));
 sg13g2_nand2_1 _4737_ (.Y(\usbfunction0.n665_o[0] ),
    .A(_0956_),
    .B(_0958_));
 sg13g2_a221oi_1 _4738_ (.B2(_0695_),
    .C1(_0954_),
    .B1(\usbfunction0.n665_o[0] ),
    .A1(_0948_),
    .Y(_0959_),
    .A2(_0949_));
 sg13g2_nor2b_1 _4739_ (.A(net1489),
    .B_N(net1827),
    .Y(_0960_));
 sg13g2_o21ai_1 _4740_ (.B1(_0960_),
    .Y(_0961_),
    .A1(net1428),
    .A2(net1426));
 sg13g2_nor2b_1 _4741_ (.A(net1491),
    .B_N(net1789),
    .Y(_0962_));
 sg13g2_nand3_1 _4742_ (.B(net1427),
    .C(net1790),
    .A(_0937_),
    .Y(_0963_));
 sg13g2_nand2_1 _4743_ (.Y(\usbfunction0.n665_o[1] ),
    .A(_0961_),
    .B(_0963_));
 sg13g2_nand3_1 _4744_ (.B(_0961_),
    .C(_0963_),
    .A(_0030_),
    .Y(_0964_));
 sg13g2_a21o_1 _4745_ (.A2(_0963_),
    .A1(_0961_),
    .B1(_0030_),
    .X(_0965_));
 sg13g2_and2_1 _4746_ (.A(_0964_),
    .B(_0965_),
    .X(_0966_));
 sg13g2_nor2b_1 _4747_ (.A(net1489),
    .B_N(net1824),
    .Y(_0967_));
 sg13g2_o21ai_1 _4748_ (.B1(_0967_),
    .Y(_0968_),
    .A1(net1428),
    .A2(net1426));
 sg13g2_nor2b_1 _4749_ (.A(net1490),
    .B_N(net1687),
    .Y(_0969_));
 sg13g2_nand3_1 _4750_ (.B(net1427),
    .C(_0969_),
    .A(_0937_),
    .Y(_0970_));
 sg13g2_nand2_1 _4751_ (.Y(\usbfunction0.n665_o[6] ),
    .A(_0968_),
    .B(_0970_));
 sg13g2_nand3_1 _4752_ (.B(_0968_),
    .C(_0970_),
    .A(_0034_),
    .Y(_0971_));
 sg13g2_a21o_1 _4753_ (.A2(_0970_),
    .A1(_0968_),
    .B1(_0034_),
    .X(_0972_));
 sg13g2_a22oi_1 _4754_ (.Y(_0973_),
    .B1(_0971_),
    .B2(_0972_),
    .A2(_0965_),
    .A1(_0964_));
 sg13g2_nor2b_1 _4755_ (.A(net1489),
    .B_N(net1876),
    .Y(_0974_));
 sg13g2_o21ai_1 _4756_ (.B1(_0974_),
    .Y(_0975_),
    .A1(net1428),
    .A2(net1426));
 sg13g2_nor2b_1 _4757_ (.A(net1490),
    .B_N(net1788),
    .Y(_0976_));
 sg13g2_nand3_1 _4758_ (.B(net1427),
    .C(_0976_),
    .A(_0937_),
    .Y(_0977_));
 sg13g2_nand2_1 _4759_ (.Y(\usbfunction0.n665_o[2] ),
    .A(_0975_),
    .B(_0977_));
 sg13g2_nor2b_1 _4760_ (.A(net1490),
    .B_N(\usbfunction0.functionreset0.in_unnamed[4] ),
    .Y(_0978_));
 sg13g2_o21ai_1 _4761_ (.B1(_0978_),
    .Y(_0979_),
    .A1(net1428),
    .A2(net1426));
 sg13g2_nor2b_1 _4762_ (.A(net1490),
    .B_N(net1845),
    .Y(_0980_));
 sg13g2_nand3_1 _4763_ (.B(net1427),
    .C(_0980_),
    .A(_0937_),
    .Y(_0981_));
 sg13g2_nand2_1 _4764_ (.Y(\usbfunction0.n665_o[4] ),
    .A(_0979_),
    .B(net1846));
 sg13g2_a21oi_1 _4765_ (.A1(_0979_),
    .A2(_0981_),
    .Y(_0982_),
    .B1(\usbfunction0.n1583_o[4] ));
 sg13g2_nor2b_1 _4766_ (.A(net1490),
    .B_N(net1886),
    .Y(_0983_));
 sg13g2_o21ai_1 _4767_ (.B1(_0983_),
    .Y(_0984_),
    .A1(net1428),
    .A2(net1426));
 sg13g2_nor2b_1 _4768_ (.A(net1490),
    .B_N(\usbfunction0.functionreset0.in_unnamed_3[5] ),
    .Y(_0985_));
 sg13g2_nand3_1 _4769_ (.B(net1427),
    .C(_0985_),
    .A(_0937_),
    .Y(_0986_));
 sg13g2_nand2_1 _4770_ (.Y(\usbfunction0.n665_o[5] ),
    .A(_0984_),
    .B(_0986_));
 sg13g2_a221oi_1 _4771_ (.B2(_0033_),
    .C1(_0982_),
    .B1(\usbfunction0.n665_o[5] ),
    .A1(_0031_),
    .Y(_0987_),
    .A2(\usbfunction0.n665_o[2] ));
 sg13g2_and3_1 _4772_ (.X(_0988_),
    .A(_0700_),
    .B(_0984_),
    .C(_0986_));
 sg13g2_and3_1 _4773_ (.X(_0989_),
    .A(\usbfunction0.n1583_o[0] ),
    .B(_0956_),
    .C(_0958_));
 sg13g2_and3_1 _4774_ (.X(_0990_),
    .A(_0696_),
    .B(_0975_),
    .C(_0977_));
 sg13g2_and3_1 _4775_ (.X(_0991_),
    .A(\usbfunction0.n1583_o[4] ),
    .B(_0979_),
    .C(_0981_));
 sg13g2_nor4_1 _4776_ (.A(_0988_),
    .B(_0989_),
    .C(_0990_),
    .D(_0991_),
    .Y(_0992_));
 sg13g2_nand4_1 _4777_ (.B(_0973_),
    .C(_0987_),
    .A(_0959_),
    .Y(_0993_),
    .D(_0992_));
 sg13g2_xnor2_1 _4778_ (.Y(_0994_),
    .A(_0695_),
    .B(\usbfunction0.n665_o[0] ));
 sg13g2_xnor2_1 _4779_ (.Y(_0995_),
    .A(_0031_),
    .B(\usbfunction0.n665_o[2] ));
 sg13g2_nor2_1 _4780_ (.A(_0982_),
    .B(_0991_),
    .Y(_0996_));
 sg13g2_xnor2_1 _4781_ (.Y(_0997_),
    .A(_0700_),
    .B(\usbfunction0.n665_o[5] ));
 sg13g2_nand3_1 _4782_ (.B(_0945_),
    .C(_0947_),
    .A(_0698_),
    .Y(_0998_));
 sg13g2_a21o_1 _4783_ (.A2(_0972_),
    .A1(_0971_),
    .B1(_0994_),
    .X(_0999_));
 sg13g2_a21oi_1 _4784_ (.A1(_0032_),
    .A2(\usbfunction0.n665_o[3] ),
    .Y(_1000_),
    .B1(_0954_));
 sg13g2_nand4_1 _4785_ (.B(_0997_),
    .C(_0998_),
    .A(_0996_),
    .Y(_1001_),
    .D(_1000_));
 sg13g2_or4_1 _4786_ (.A(_0966_),
    .B(_0995_),
    .C(_0999_),
    .D(_1001_),
    .X(_1002_));
 sg13g2_mux2_2 _4787_ (.A0(_0703_),
    .A1(_0704_),
    .S(net1397),
    .X(_1003_));
 sg13g2_inv_2 _4788_ (.Y(\s_m_pushdata_endpoint[0] ),
    .A(_1003_));
 sg13g2_mux2_1 _4789_ (.A0(net1481),
    .A1(net1042),
    .S(net1396),
    .X(\s_m_pushdata_endpoint[1] ));
 sg13g2_or2_1 _4790_ (.X(_1004_),
    .B(net1381),
    .A(_1003_));
 sg13g2_mux2_2 _4791_ (.A0(net1478),
    .A1(net1765),
    .S(net1396),
    .X(\s_m_pushdata_endpoint[2] ));
 sg13g2_mux2_2 _4792_ (.A0(net1477),
    .A1(net1795),
    .S(net1396),
    .X(\s_m_pushdata_endpoint[3] ));
 sg13g2_nor2_1 _4793_ (.A(\s_m_pushdata_endpoint[2] ),
    .B(\s_m_pushdata_endpoint[3] ),
    .Y(_1005_));
 sg13g2_nor4_2 _4794_ (.A(_1003_),
    .B(net1381),
    .C(\s_m_pushdata_endpoint[2] ),
    .Y(_1006_),
    .D(\s_m_pushdata_endpoint[3] ));
 sg13g2_nand3_1 _4795_ (.B(net1427),
    .C(_1006_),
    .A(net1428),
    .Y(_1007_));
 sg13g2_xnor2_1 _4796_ (.Y(_1008_),
    .A(\usbfunction0.n2313_o[1] ),
    .B(\usbfunction0.n2640_q[1] ));
 sg13g2_xnor2_1 _4797_ (.Y(_1009_),
    .A(\usbfunction0.n2313_o[0] ),
    .B(\usbfunction0.n2640_q[0] ));
 sg13g2_xnor2_1 _4798_ (.Y(_1010_),
    .A(\usbfunction0.n2313_o[3] ),
    .B(\usbfunction0.n2640_q[3] ));
 sg13g2_xnor2_1 _4799_ (.Y(_1011_),
    .A(\usbfunction0.n2313_o[2] ),
    .B(\usbfunction0.n2640_q[2] ));
 sg13g2_nand4_1 _4800_ (.B(_1009_),
    .C(_1010_),
    .A(_1008_),
    .Y(_1012_),
    .D(_1011_));
 sg13g2_and2_1 _4801_ (.A(_0718_),
    .B(_1006_),
    .X(_1013_));
 sg13g2_and2_1 _4802_ (.A(_1012_),
    .B(_1013_),
    .X(_1014_));
 sg13g2_nor2b_1 _4803_ (.A(\usbfunction0.n2634_q[0] ),
    .B_N(\usbfunction0.n2634_q[1] ),
    .Y(_1015_));
 sg13g2_nor2b_1 _4804_ (.A(\usbfunction0.n2634_q[3] ),
    .B_N(\usbfunction0.n2634_q[2] ),
    .Y(_1016_));
 sg13g2_nand2_1 _4805_ (.Y(_1017_),
    .A(_1015_),
    .B(_1016_));
 sg13g2_inv_1 _4806_ (.Y(_1018_),
    .A(_1017_));
 sg13g2_nand4_1 _4807_ (.B(_1006_),
    .C(_1012_),
    .A(_0718_),
    .Y(_1019_),
    .D(_1018_));
 sg13g2_or4_1 _4808_ (.A(\usbfunction0.n2650_q[0] ),
    .B(\usbfunction0.n2650_q[1] ),
    .C(\usbfunction0.n2650_q[2] ),
    .D(\usbfunction0.n2650_q[3] ),
    .X(_1020_));
 sg13g2_nor2_1 _4809_ (.A(\usbfunction0.n2650_q[4] ),
    .B(_1020_),
    .Y(_1021_));
 sg13g2_nor3_1 _4810_ (.A(\usbfunction0.n2650_q[4] ),
    .B(\usbfunction0.n2650_q[5] ),
    .C(_1020_),
    .Y(_1022_));
 sg13g2_nand2b_1 _4811_ (.Y(_1023_),
    .B(_1021_),
    .A_N(\usbfunction0.n2650_q[5] ));
 sg13g2_nor2_1 _4812_ (.A(\usbfunction0.n2650_q[6] ),
    .B(_1023_),
    .Y(_1024_));
 sg13g2_nor3_2 _4813_ (.A(\usbfunction0.n2313_o[2] ),
    .B(\usbfunction0.n2313_o[1] ),
    .C(\usbfunction0.n2313_o[0] ),
    .Y(_1025_));
 sg13g2_a22oi_1 _4814_ (.Y(_1026_),
    .B1(_1025_),
    .B2(\usbfunction0.n2313_o[3] ),
    .A2(_1024_),
    .A1(_0720_));
 sg13g2_nand2_1 _4815_ (.Y(_1027_),
    .A(_0805_),
    .B(_1015_));
 sg13g2_and3_1 _4816_ (.X(_1028_),
    .A(_0805_),
    .B(_1015_),
    .C(_1026_));
 sg13g2_nand2_2 _4817_ (.Y(_1029_),
    .A(_0950_),
    .B(_1016_));
 sg13g2_nor2b_2 _4818_ (.A(net1394),
    .B_N(_1029_),
    .Y(_1030_));
 sg13g2_nand2b_1 _4819_ (.Y(_1031_),
    .B(_1029_),
    .A_N(net1394));
 sg13g2_nand3_1 _4820_ (.B(net1367),
    .C(_1030_),
    .A(_0719_),
    .Y(s_m_phy_tx_valid_2));
 sg13g2_nand4_1 _4821_ (.B(\usbfunction0.scl_usbgpiophy0.n6654_q ),
    .C(net1367),
    .A(_0719_),
    .Y(_1032_),
    .D(_1030_));
 sg13g2_and2_1 _4822_ (.A(_0721_),
    .B(_1032_),
    .X(_1033_));
 sg13g2_nand2_2 _4823_ (.Y(_1034_),
    .A(_0777_),
    .B(_0779_));
 sg13g2_nand2_1 _4824_ (.Y(_1035_),
    .A(net1488),
    .B(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.s_m_value[0] ));
 sg13g2_nand4_1 _4825_ (.B(net1132),
    .C(net1488),
    .A(net1878),
    .Y(_1036_),
    .D(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.s_m_value[0] ));
 sg13g2_nor2_1 _4826_ (.A(_1034_),
    .B(_1036_),
    .Y(_1037_));
 sg13g2_nor2_2 _4827_ (.A(_0043_),
    .B(_1037_),
    .Y(_1038_));
 sg13g2_or2_1 _4828_ (.X(_1039_),
    .B(_1037_),
    .A(_0043_));
 sg13g2_and2_2 _4829_ (.A(_1033_),
    .B(net1392),
    .X(_1040_));
 sg13g2_nor3_2 _4830_ (.A(\usbfunction0.scl_usbgpiophy0.scl_addeopdeferred0.n7349_q ),
    .B(net1365),
    .C(_1038_),
    .Y(_1041_));
 sg13g2_inv_1 _4831_ (.Y(_1042_),
    .A(_1041_));
 sg13g2_and3_1 _4832_ (.X(_1043_),
    .A(\scl_fifo1.n6321_q[0] ),
    .B(\scl_fifo1.n6321_q[1] ),
    .C(_1041_));
 sg13g2_nand3_1 _4833_ (.B(\scl_fifo1.n6321_q[3] ),
    .C(_1043_),
    .A(\scl_fifo1.n6321_q[2] ),
    .Y(_1044_));
 sg13g2_xnor2_1 _4834_ (.Y(_1045_),
    .A(net1164),
    .B(_1044_));
 sg13g2_mux2_1 _4835_ (.A0(net1105),
    .A1(net1165),
    .S(_1007_),
    .X(\scl_fifo1.n6238_o[4] ));
 sg13g2_xor2_1 _4836_ (.B(\scl_fifo1.n6238_o[4] ),
    .A(net1024),
    .X(_1046_));
 sg13g2_nor3_1 _4837_ (.A(\scl_fifo1.n6321_q[0] ),
    .B(\scl_fifo1.n6321_q[1] ),
    .C(_1042_),
    .Y(_1047_));
 sg13g2_nor2b_1 _4838_ (.A(_1041_),
    .B_N(net1153),
    .Y(_1048_));
 sg13g2_nor3_1 _4839_ (.A(_1043_),
    .B(_1047_),
    .C(_1048_),
    .Y(_1049_));
 sg13g2_mux2_2 _4840_ (.A0(\scl_fifo1.n6323_q[1] ),
    .A1(_1049_),
    .S(_1007_),
    .X(\scl_fifo1.n6238_o[1] ));
 sg13g2_xor2_1 _4841_ (.B(net1295),
    .A(\scl_fifo1.n6229_o[1] ),
    .X(_1050_));
 sg13g2_nor2_1 _4842_ (.A(\scl_fifo1.n6323_q[3] ),
    .B(_1007_),
    .Y(_1051_));
 sg13g2_nor2b_1 _4843_ (.A(net917),
    .B_N(_1043_),
    .Y(_1052_));
 sg13g2_xnor2_1 _4844_ (.Y(_1053_),
    .A(net1634),
    .B(_1052_));
 sg13g2_nand2b_1 _4845_ (.Y(_1054_),
    .B(_1007_),
    .A_N(_1053_));
 sg13g2_nand2b_2 _4846_ (.Y(_1055_),
    .B(_1054_),
    .A_N(_1051_));
 sg13g2_inv_2 _4847_ (.Y(\scl_fifo1.n6238_o[3] ),
    .A(net1274));
 sg13g2_xnor2_1 _4848_ (.Y(_1056_),
    .A(\scl_fifo1.n6229_o[3] ),
    .B(net1266));
 sg13g2_xor2_1 _4849_ (.B(_1041_),
    .A(net1618),
    .X(_1057_));
 sg13g2_nand2b_1 _4850_ (.Y(_1058_),
    .B(_1007_),
    .A_N(_1057_));
 sg13g2_o21ai_1 _4851_ (.B1(_1058_),
    .Y(_1059_),
    .A1(\scl_fifo1.n6323_q[0] ),
    .A2(_1007_));
 sg13g2_inv_1 _4852_ (.Y(\scl_fifo1.n6238_o[0] ),
    .A(net1322));
 sg13g2_xor2_1 _4853_ (.B(net1286),
    .A(\scl_fifo1.n6229_o[0] ),
    .X(_1060_));
 sg13g2_nor2_1 _4854_ (.A(\scl_fifo1.n6323_q[2] ),
    .B(_1007_),
    .Y(_1061_));
 sg13g2_xnor2_1 _4855_ (.Y(_1062_),
    .A(net917),
    .B(_1043_));
 sg13g2_inv_1 _4856_ (.Y(_1063_),
    .A(_1062_));
 sg13g2_a21o_2 _4857_ (.A2(_1063_),
    .A1(_1007_),
    .B1(_1061_),
    .X(_1064_));
 sg13g2_inv_1 _4858_ (.Y(\scl_fifo1.n6238_o[2] ),
    .A(_1064_));
 sg13g2_xor2_1 _4859_ (.B(net1273),
    .A(\scl_fifo1.n6229_o[2] ),
    .X(_1065_));
 sg13g2_nor3_1 _4860_ (.A(_1050_),
    .B(_1060_),
    .C(_1065_),
    .Y(_1066_));
 sg13g2_nand3_1 _4861_ (.B(_1056_),
    .C(_1066_),
    .A(_1046_),
    .Y(_0178_));
 sg13g2_nor2b_1 _4862_ (.A(\scl_streamarbiter_2.n6192_q ),
    .B_N(\scl_streamarbiter_2.n6195_q ),
    .Y(_1067_));
 sg13g2_nand2_1 _4863_ (.Y(_1068_),
    .A(_0724_),
    .B(_1067_));
 sg13g2_o21ai_1 _4864_ (.B1(_1068_),
    .Y(_1069_),
    .A1(\scl_streamarbiter_2.n6194_q ),
    .A2(_1067_));
 sg13g2_inv_1 _4865_ (.Y(\scl_streamarbiter_2.n6146_o ),
    .A(net1416));
 sg13g2_or2_2 _4866_ (.X(_1070_),
    .B(net1417),
    .A(s_m_pushfull_2));
 sg13g2_nor2_1 _4867_ (.A(\scl_bitbangengine0.n5898_q[3] ),
    .B(\scl_bitbangengine0.n5898_q[2] ),
    .Y(_1071_));
 sg13g2_nor2b_1 _4868_ (.A(_1070_),
    .B_N(_1071_),
    .Y(_1072_));
 sg13g2_nor2_1 _4869_ (.A(_0724_),
    .B(s_m_popempty),
    .Y(_1073_));
 sg13g2_nand2b_1 _4870_ (.Y(_1074_),
    .B(n346_q),
    .A_N(s_m_popempty));
 sg13g2_nor2_1 _4871_ (.A(net1503),
    .B(\scl_bitbangengine0.n5898_q[1] ),
    .Y(_1075_));
 sg13g2_nor2b_1 _4872_ (.A(_1074_),
    .B_N(_1075_),
    .Y(_1076_));
 sg13g2_and2_2 _4873_ (.A(_1072_),
    .B(_1076_),
    .X(_1077_));
 sg13g2_nand2_2 _4874_ (.Y(_1078_),
    .A(_1072_),
    .B(_1076_));
 sg13g2_nand2_2 _4875_ (.Y(_1079_),
    .A(\scl_bitbangengine0.n3179_o ),
    .B(_1077_));
 sg13g2_and3_1 _4876_ (.X(_1080_),
    .A(_0692_),
    .B(_0694_),
    .C(net1493));
 sg13g2_nor2_1 _4877_ (.A(net1500),
    .B(net1451),
    .Y(_1081_));
 sg13g2_and2_1 _4878_ (.A(_1080_),
    .B(_1081_),
    .X(_1082_));
 sg13g2_nand2_1 _4879_ (.Y(_1083_),
    .A(_1080_),
    .B(_1081_));
 sg13g2_a21o_1 _4880_ (.A2(_1082_),
    .A1(net1497),
    .B1(_1079_),
    .X(_1084_));
 sg13g2_nand2_1 _4881_ (.Y(_1085_),
    .A(net1495),
    .B(net1500));
 sg13g2_nor2_1 _4882_ (.A(\scl_bitbangengine0.n3230_o ),
    .B(net1451),
    .Y(_1086_));
 sg13g2_nand4_1 _4883_ (.B(net1500),
    .C(_1080_),
    .A(net1495),
    .Y(_1087_),
    .D(_1086_));
 sg13g2_nand2_2 _4884_ (.Y(_1088_),
    .A(_0692_),
    .B(\scl_bitbangengine0.n3258_o ));
 sg13g2_nor3_2 _4885_ (.A(\scl_bitbangengine0.n3267_o ),
    .B(\scl_bitbangengine0.n3258_o ),
    .C(net1493),
    .Y(_1089_));
 sg13g2_o21ai_1 _4886_ (.B1(_1089_),
    .Y(_1090_),
    .A1(net1498),
    .A2(_1085_));
 sg13g2_nand3_1 _4887_ (.B(_1088_),
    .C(_1090_),
    .A(_1087_),
    .Y(_1091_));
 sg13g2_nor3_2 _4888_ (.A(_1079_),
    .B(_1082_),
    .C(_1091_),
    .Y(_1092_));
 sg13g2_nand2b_1 _4889_ (.Y(_1093_),
    .B(net1503),
    .A_N(\scl_bitbangengine0.n5898_q[1] ));
 sg13g2_nor4_1 _4890_ (.A(\scl_bitbangengine0.n5898_q[3] ),
    .B(\scl_bitbangengine0.n5898_q[2] ),
    .C(_1070_),
    .D(_1093_),
    .Y(_1094_));
 sg13g2_nor2_2 _4891_ (.A(_1092_),
    .B(net1405),
    .Y(_1095_));
 sg13g2_nor2b_1 _4892_ (.A(_1079_),
    .B_N(_1089_),
    .Y(_1096_));
 sg13g2_nand3_1 _4893_ (.B(_1077_),
    .C(_1089_),
    .A(net1492),
    .Y(_1097_));
 sg13g2_nor2_1 _4894_ (.A(net1495),
    .B(_1097_),
    .Y(_1098_));
 sg13g2_nor4_2 _4895_ (.A(net1495),
    .B(_0729_),
    .C(net1498),
    .Y(_1099_),
    .D(_1097_));
 sg13g2_nor3_2 _4896_ (.A(net1495),
    .B(net1498),
    .C(_1097_),
    .Y(_1100_));
 sg13g2_and2_2 _4897_ (.A(net1502),
    .B(_1100_),
    .X(_1101_));
 sg13g2_nand3b_1 _4898_ (.B(_1095_),
    .C(\scl_streamarbiter_2.n6146_o ),
    .Y(_1102_),
    .A_N(_1101_));
 sg13g2_nor2_1 _4899_ (.A(_1079_),
    .B(_1088_),
    .Y(_1103_));
 sg13g2_nor2_1 _4900_ (.A(\scl_bitbangengine0.n5921_q[0] ),
    .B(\scl_bitbangengine0.n5921_q[1] ),
    .Y(_1104_));
 sg13g2_or4_2 _4901_ (.A(\scl_bitbangengine0.n5921_q[0] ),
    .B(\scl_bitbangengine0.n5921_q[1] ),
    .C(\scl_bitbangengine0.n5921_q[2] ),
    .D(\scl_bitbangengine0.n5921_q[3] ),
    .X(_1105_));
 sg13g2_or3_1 _4902_ (.A(\scl_bitbangengine0.n5921_q[4] ),
    .B(\scl_bitbangengine0.n5921_q[5] ),
    .C(_1105_),
    .X(_1106_));
 sg13g2_or2_1 _4903_ (.X(_1107_),
    .B(\scl_bitbangengine0.n5921_q[7] ),
    .A(\scl_bitbangengine0.n5921_q[6] ));
 sg13g2_or4_2 _4904_ (.A(\scl_bitbangengine0.n5921_q[4] ),
    .B(\scl_bitbangengine0.n5921_q[5] ),
    .C(_1105_),
    .D(_1107_),
    .X(_1108_));
 sg13g2_or3_1 _4905_ (.A(\scl_bitbangengine0.n3663_o[0] ),
    .B(\scl_bitbangengine0.n3663_o[1] ),
    .C(_1108_),
    .X(_1109_));
 sg13g2_or2_1 _4906_ (.X(_1110_),
    .B(\scl_bitbangengine0.n3663_o[3] ),
    .A(\scl_bitbangengine0.n3663_o[2] ));
 sg13g2_or4_2 _4907_ (.A(\scl_bitbangengine0.n3663_o[0] ),
    .B(\scl_bitbangengine0.n3663_o[1] ),
    .C(_1108_),
    .D(_1110_),
    .X(_1111_));
 sg13g2_nor3_2 _4908_ (.A(\scl_bitbangengine0.n3663_o[4] ),
    .B(\scl_bitbangengine0.n3663_o[5] ),
    .C(_1111_),
    .Y(_1112_));
 sg13g2_o21ai_1 _4909_ (.B1(\scl_bitbangengine0.n3663_o[5] ),
    .Y(_1113_),
    .A1(\scl_bitbangengine0.n3663_o[4] ),
    .A2(_1111_));
 sg13g2_nor2b_1 _4910_ (.A(_1112_),
    .B_N(_1113_),
    .Y(_1114_));
 sg13g2_xnor2_1 _4911_ (.Y(_1115_),
    .A(_0076_),
    .B(_1114_));
 sg13g2_nor2_1 _4912_ (.A(\scl_bitbangengine0.n3663_o[6] ),
    .B(\scl_bitbangengine0.n3663_o[7] ),
    .Y(_1116_));
 sg13g2_and2_1 _4913_ (.A(_1112_),
    .B(_1116_),
    .X(_1117_));
 sg13g2_xnor2_1 _4914_ (.Y(_1118_),
    .A(\scl_bitbangengine0.n3663_o[8] ),
    .B(_0080_));
 sg13g2_xnor2_1 _4915_ (.Y(_1119_),
    .A(_1117_),
    .B(_1118_));
 sg13g2_nand2_1 _4916_ (.Y(_1120_),
    .A(_1115_),
    .B(_1119_));
 sg13g2_and2_1 _4917_ (.A(_0078_),
    .B(_1112_),
    .X(_1121_));
 sg13g2_xor2_1 _4918_ (.B(_0079_),
    .A(\scl_bitbangengine0.n3663_o[7] ),
    .X(_1122_));
 sg13g2_xnor2_1 _4919_ (.Y(_1123_),
    .A(_1121_),
    .B(_1122_));
 sg13g2_xnor2_1 _4920_ (.Y(_1124_),
    .A(_0078_),
    .B(_1112_));
 sg13g2_xor2_1 _4921_ (.B(_1124_),
    .A(_0077_),
    .X(_1125_));
 sg13g2_xor2_1 _4922_ (.B(_1111_),
    .A(\scl_bitbangengine0.n3663_o[4] ),
    .X(_1126_));
 sg13g2_xnor2_1 _4923_ (.Y(_1127_),
    .A(_0075_),
    .B(_1126_));
 sg13g2_o21ai_1 _4924_ (.B1(\scl_bitbangengine0.n3663_o[1] ),
    .Y(_1128_),
    .A1(\scl_bitbangengine0.n3663_o[0] ),
    .A2(_1108_));
 sg13g2_a21oi_1 _4925_ (.A1(_1109_),
    .A2(_1128_),
    .Y(_1129_),
    .B1(_0071_));
 sg13g2_and3_1 _4926_ (.X(_1130_),
    .A(_0071_),
    .B(_1109_),
    .C(_1128_));
 sg13g2_nor4_1 _4927_ (.A(\scl_bitbangengine0.n3663_o[0] ),
    .B(\scl_bitbangengine0.n3663_o[1] ),
    .C(_0728_),
    .D(_1108_),
    .Y(_1131_));
 sg13g2_xnor2_1 _4928_ (.Y(_1132_),
    .A(\scl_bitbangengine0.n3663_o[3] ),
    .B(_0074_));
 sg13g2_xnor2_1 _4929_ (.Y(_1133_),
    .A(_1131_),
    .B(_1132_));
 sg13g2_o21ai_1 _4930_ (.B1(_1133_),
    .Y(_1134_),
    .A1(_1129_),
    .A2(_1130_));
 sg13g2_xnor2_1 _4931_ (.Y(_1135_),
    .A(_0728_),
    .B(_1109_));
 sg13g2_nor2_1 _4932_ (.A(_0072_),
    .B(_1135_),
    .Y(_1136_));
 sg13g2_and2_1 _4933_ (.A(_0072_),
    .B(_1135_),
    .X(_1137_));
 sg13g2_xor2_1 _4934_ (.B(_1108_),
    .A(\scl_bitbangengine0.n3663_o[0] ),
    .X(_1138_));
 sg13g2_nand2b_1 _4935_ (.Y(_1139_),
    .B(_0070_),
    .A_N(_1138_));
 sg13g2_xnor2_1 _4936_ (.Y(_1140_),
    .A(_0070_),
    .B(_1138_));
 sg13g2_xnor2_1 _4937_ (.Y(_1141_),
    .A(\scl_bitbangengine0.n5921_q[7] ),
    .B(_0069_));
 sg13g2_nand2b_1 _4938_ (.Y(_1142_),
    .B(_0068_),
    .A_N(_0067_));
 sg13g2_o21ai_1 _4939_ (.B1(_1142_),
    .Y(_1143_),
    .A1(_1106_),
    .A2(_1141_));
 sg13g2_a21oi_1 _4940_ (.A1(_0726_),
    .A2(_0067_),
    .Y(_1144_),
    .B1(_1141_));
 sg13g2_nor2_1 _4941_ (.A(_1106_),
    .B(_1144_),
    .Y(_1145_));
 sg13g2_mux2_1 _4942_ (.A0(_1144_),
    .A1(_1145_),
    .S(_1143_),
    .X(_1146_));
 sg13g2_o21ai_1 _4943_ (.B1(\scl_bitbangengine0.n5921_q[5] ),
    .Y(_1147_),
    .A1(\scl_bitbangengine0.n5921_q[4] ),
    .A2(_1105_));
 sg13g2_nand2_1 _4944_ (.Y(_1148_),
    .A(_1106_),
    .B(_1147_));
 sg13g2_xor2_1 _4945_ (.B(_1148_),
    .A(_0066_),
    .X(_1149_));
 sg13g2_xnor2_1 _4946_ (.Y(_1150_),
    .A(\scl_bitbangengine0.n5921_q[4] ),
    .B(_1105_));
 sg13g2_xnor2_1 _4947_ (.Y(_1151_),
    .A(_0065_),
    .B(_1150_));
 sg13g2_xor2_1 _4948_ (.B(\scl_bitbangengine0.scl_counter0.n6975_q[1] ),
    .A(\scl_bitbangengine0.n5921_q[1] ),
    .X(_1152_));
 sg13g2_a21oi_1 _4949_ (.A1(_0725_),
    .A2(\scl_bitbangengine0.n5921_q[0] ),
    .Y(_1153_),
    .B1(_1152_));
 sg13g2_o21ai_1 _4950_ (.B1(_1152_),
    .Y(_1154_),
    .A1(_0725_),
    .A2(\scl_bitbangengine0.n5921_q[0] ));
 sg13g2_nand2b_1 _4951_ (.Y(_1155_),
    .B(_1154_),
    .A_N(_1153_));
 sg13g2_nand2_1 _4952_ (.Y(_1156_),
    .A(_0063_),
    .B(_1104_));
 sg13g2_xnor2_1 _4953_ (.Y(_1157_),
    .A(\scl_bitbangengine0.n5921_q[3] ),
    .B(_0064_));
 sg13g2_xnor2_1 _4954_ (.Y(_1158_),
    .A(_1156_),
    .B(_1157_));
 sg13g2_xnor2_1 _4955_ (.Y(_1159_),
    .A(_0063_),
    .B(_1104_));
 sg13g2_xnor2_1 _4956_ (.Y(_1160_),
    .A(_0062_),
    .B(_1159_));
 sg13g2_nor4_2 _4957_ (.A(_1151_),
    .B(_1155_),
    .C(_1158_),
    .Y(_1161_),
    .D(_1160_));
 sg13g2_nand4_1 _4958_ (.B(_1146_),
    .C(_1149_),
    .A(_1140_),
    .Y(_1162_),
    .D(_1161_));
 sg13g2_nor4_1 _4959_ (.A(_1134_),
    .B(_1136_),
    .C(_1137_),
    .D(_1162_),
    .Y(_1163_));
 sg13g2_nand3_1 _4960_ (.B(_1127_),
    .C(_1163_),
    .A(_1125_),
    .Y(_1164_));
 sg13g2_nor3_1 _4961_ (.A(_1120_),
    .B(_1123_),
    .C(_1164_),
    .Y(_1165_));
 sg13g2_and2_2 _4962_ (.A(_1103_),
    .B(net1371),
    .X(_1166_));
 sg13g2_xnor2_1 _4963_ (.Y(_1167_),
    .A(\scl_bitbangengine0.n3663_o[7] ),
    .B(_1121_));
 sg13g2_nor2b_1 _4964_ (.A(_0079_),
    .B_N(_1167_),
    .Y(_1168_));
 sg13g2_nand2b_1 _4965_ (.Y(_1169_),
    .B(_0075_),
    .A_N(_1126_));
 sg13g2_nand2b_1 _4966_ (.Y(_1170_),
    .B(_1126_),
    .A_N(_0075_));
 sg13g2_nor2b_1 _4967_ (.A(_1167_),
    .B_N(_0079_),
    .Y(_1171_));
 sg13g2_nand3_1 _4968_ (.B(_1149_),
    .C(_1161_),
    .A(_1139_),
    .Y(_1172_));
 sg13g2_a21oi_1 _4969_ (.A1(_0727_),
    .A2(_1138_),
    .Y(_1173_),
    .B1(_1172_));
 sg13g2_nand4_1 _4970_ (.B(_1169_),
    .C(_1170_),
    .A(_1146_),
    .Y(_1174_),
    .D(_1173_));
 sg13g2_or3_1 _4971_ (.A(_1134_),
    .B(_1136_),
    .C(_1137_),
    .X(_1175_));
 sg13g2_nor4_1 _4972_ (.A(_1168_),
    .B(_1171_),
    .C(_1174_),
    .D(_1175_),
    .Y(_1176_));
 sg13g2_nand4_1 _4973_ (.B(_1119_),
    .C(_1125_),
    .A(_1115_),
    .Y(_1177_),
    .D(_1176_));
 sg13g2_nor3_2 _4974_ (.A(_1079_),
    .B(_1088_),
    .C(_1177_),
    .Y(_1178_));
 sg13g2_a21oi_1 _4975_ (.A1(net1493),
    .A2(_1166_),
    .Y(_1179_),
    .B1(_1102_));
 sg13g2_xnor2_1 _4976_ (.Y(_1180_),
    .A(\scl_bitbangengine0.n5902_q ),
    .B(net14));
 sg13g2_nor4_1 _4977_ (.A(\scl_bitbangengine0.n5920_q[1] ),
    .B(\scl_bitbangengine0.n5920_q[2] ),
    .C(\scl_bitbangengine0.n5920_q[3] ),
    .D(\scl_bitbangengine0.n5920_q[16] ),
    .Y(_1181_));
 sg13g2_nand3_1 _4978_ (.B(\scl_bitbangengine0.n5920_q[0] ),
    .C(_1181_),
    .A(\scl_bitbangengine0.n5904_q ),
    .Y(_1182_));
 sg13g2_nor4_2 _4979_ (.A(\scl_bitbangengine0.n5920_q[4] ),
    .B(\scl_bitbangengine0.n5920_q[5] ),
    .C(\scl_bitbangengine0.n5920_q[6] ),
    .Y(_1183_),
    .D(\scl_bitbangengine0.n5920_q[7] ));
 sg13g2_nor3_1 _4980_ (.A(\scl_bitbangengine0.n5920_q[17] ),
    .B(\scl_bitbangengine0.n5920_q[19] ),
    .C(\scl_bitbangengine0.n5920_q[18] ),
    .Y(_1184_));
 sg13g2_nor4_2 _4981_ (.A(\scl_bitbangengine0.n5920_q[9] ),
    .B(\scl_bitbangengine0.n5920_q[8] ),
    .C(\scl_bitbangengine0.n5920_q[11] ),
    .Y(_1185_),
    .D(\scl_bitbangengine0.n5920_q[10] ));
 sg13g2_nand4_1 _4982_ (.B(_0740_),
    .C(_0741_),
    .A(_0739_),
    .Y(_1186_),
    .D(_0742_));
 sg13g2_nand3_1 _4983_ (.B(_1184_),
    .C(_1185_),
    .A(_1183_),
    .Y(_1187_));
 sg13g2_nor3_2 _4984_ (.A(_1182_),
    .B(_1186_),
    .C(_1187_),
    .Y(_1188_));
 sg13g2_a21o_2 _4985_ (.A2(_1180_),
    .A1(\scl_bitbangengine0.n5903_q ),
    .B1(_1188_),
    .X(_1189_));
 sg13g2_nor2b_1 _4986_ (.A(_0133_),
    .B_N(\scl_bitbangengine0.s_m_value_2[2] ),
    .Y(_1190_));
 sg13g2_xor2_1 _4987_ (.B(\scl_bitbangengine0.s_m_value_2[0] ),
    .A(\scl_bitbangengine0.n5905_q ),
    .X(_1191_));
 sg13g2_a21oi_1 _4988_ (.A1(_1190_),
    .A2(_1191_),
    .Y(_1192_),
    .B1(_1189_));
 sg13g2_nand2b_2 _4989_ (.Y(_1193_),
    .B(\scl_bitbangengine0.n5898_q[1] ),
    .A_N(net1503));
 sg13g2_nand2b_1 _4990_ (.Y(_1194_),
    .B(\scl_bitbangengine0.n5898_q[3] ),
    .A_N(\scl_bitbangengine0.n5898_q[2] ));
 sg13g2_a21oi_2 _4991_ (.B1(_1194_),
    .Y(_1195_),
    .A2(_1070_),
    .A1(\scl_bitbangengine0.n5910_q ));
 sg13g2_nand2_2 _4992_ (.Y(_1196_),
    .A(net1371),
    .B(_1195_));
 sg13g2_nor2_2 _4993_ (.A(_1193_),
    .B(_1196_),
    .Y(_1197_));
 sg13g2_xnor2_1 _4994_ (.Y(_1198_),
    .A(\scl_bitbangengine0.n5917_q ),
    .B(_1197_));
 sg13g2_nand2_1 _4995_ (.Y(_1199_),
    .A(\scl_bitbangengine0.n5910_q ),
    .B(_1198_));
 sg13g2_nand3_1 _4996_ (.B(_1071_),
    .C(_1073_),
    .A(\scl_bitbangengine0.n5898_q[1] ),
    .Y(_1200_));
 sg13g2_nor2_1 _4997_ (.A(\scl_bitbangengine0.n5898_q[0] ),
    .B(_1200_),
    .Y(_1201_));
 sg13g2_nor3_2 _4998_ (.A(net1503),
    .B(\scl_bitbangengine0.n3336_o ),
    .C(_1200_),
    .Y(_1202_));
 sg13g2_nor2_2 _4999_ (.A(_1166_),
    .B(_1202_),
    .Y(_1203_));
 sg13g2_mux2_1 _5000_ (.A0(net1496),
    .A1(net1877),
    .S(_1203_),
    .X(_1204_));
 sg13g2_nand4_1 _5001_ (.B(\scl_bitbangengine0.n5898_q[1] ),
    .C(_1071_),
    .A(net1503),
    .Y(_1205_),
    .D(_1073_));
 sg13g2_nor2_2 _5002_ (.A(\scl_bitbangengine0.n3336_o ),
    .B(_1205_),
    .Y(_1206_));
 sg13g2_mux2_1 _5003_ (.A0(net1669),
    .A1(net1496),
    .S(net1414),
    .X(\scl_bitbangengine0.n3793_o ));
 sg13g2_xor2_1 _5004_ (.B(_1204_),
    .A(net12),
    .X(_1207_));
 sg13g2_a21oi_1 _5005_ (.A1(\scl_bitbangengine0.n5911_q ),
    .A2(_1074_),
    .Y(_1208_),
    .B1(_1093_));
 sg13g2_nand3_1 _5006_ (.B(_1195_),
    .C(_1208_),
    .A(net1371),
    .Y(_1209_));
 sg13g2_a21oi_2 _5007_ (.B1(_1209_),
    .Y(_1210_),
    .A2(_1207_),
    .A1(\scl_bitbangengine0.n3793_o ));
 sg13g2_inv_2 _5008_ (.Y(_1211_),
    .A(_1210_));
 sg13g2_or2_2 _5009_ (.X(_1212_),
    .B(_1210_),
    .A(_1197_));
 sg13g2_nor2b_1 _5010_ (.A(_1199_),
    .B_N(_1212_),
    .Y(_1213_));
 sg13g2_nand2b_2 _5011_ (.Y(_1214_),
    .B(_1212_),
    .A_N(_1199_));
 sg13g2_nand2b_2 _5012_ (.Y(_1215_),
    .B(net1270),
    .A_N(_1192_));
 sg13g2_a22oi_1 _5013_ (.Y(_1216_),
    .B1(_1179_),
    .B2(_1215_),
    .A2(net1417),
    .A1(_0151_));
 sg13g2_nor2b_1 _5014_ (.A(net556),
    .B_N(_1216_),
    .Y(_0177_));
 sg13g2_and2_1 _5015_ (.A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[10] ),
    .B(\n352_o[17] ),
    .X(_1217_));
 sg13g2_xor2_1 _5016_ (.B(\n352_o[17] ),
    .A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[10] ),
    .X(_1218_));
 sg13g2_xnor2_1 _5017_ (.Y(_1219_),
    .A(_0766_),
    .B(\n352_o[18] ));
 sg13g2_and2_1 _5018_ (.A(_1218_),
    .B(_1219_),
    .X(_1220_));
 sg13g2_and2_1 _5019_ (.A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[8] ),
    .B(_0820_),
    .X(_1221_));
 sg13g2_nand2_1 _5020_ (.Y(_1222_),
    .A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[8] ),
    .B(_0820_));
 sg13g2_o21ai_1 _5021_ (.B1(_1221_),
    .Y(_1223_),
    .A1(\scl_uarttx0.scl_baudrategenerator0.n6874_o[9] ),
    .A2(_0818_));
 sg13g2_inv_1 _5022_ (.Y(_1224_),
    .A(_1223_));
 sg13g2_a21oi_1 _5023_ (.A1(\scl_uarttx0.scl_baudrategenerator0.n6874_o[9] ),
    .A2(_0818_),
    .Y(_1225_),
    .B1(_1224_));
 sg13g2_and2_1 _5024_ (.A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[7] ),
    .B(_0822_),
    .X(_1226_));
 sg13g2_nand2_1 _5025_ (.Y(_1227_),
    .A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[6] ),
    .B(\n352_o[13] ));
 sg13g2_xnor2_1 _5026_ (.Y(_1228_),
    .A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[6] ),
    .B(\n352_o[13] ));
 sg13g2_nor2_1 _5027_ (.A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[5] ),
    .B(\n352_o[12] ),
    .Y(_1229_));
 sg13g2_nand2_1 _5028_ (.Y(_1230_),
    .A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[3] ),
    .B(\n352_o[10] ));
 sg13g2_and2_1 _5029_ (.A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[2] ),
    .B(_0828_),
    .X(_1231_));
 sg13g2_nand2_1 _5030_ (.Y(_1232_),
    .A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[1] ),
    .B(\n352_o[8] ));
 sg13g2_nand2_1 _5031_ (.Y(_1233_),
    .A(net611),
    .B(\n352_o[7] ));
 sg13g2_xnor2_1 _5032_ (.Y(_1234_),
    .A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[1] ),
    .B(\n352_o[8] ));
 sg13g2_o21ai_1 _5033_ (.B1(_1232_),
    .Y(_1235_),
    .A1(_1233_),
    .A2(_1234_));
 sg13g2_xor2_1 _5034_ (.B(_0828_),
    .A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[2] ),
    .X(_1236_));
 sg13g2_a21oi_1 _5035_ (.A1(_1235_),
    .A2(_1236_),
    .Y(_1237_),
    .B1(_1231_));
 sg13g2_nor2_1 _5036_ (.A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[3] ),
    .B(\n352_o[10] ),
    .Y(_1238_));
 sg13g2_xor2_1 _5037_ (.B(\n352_o[10] ),
    .A(net1901),
    .X(_1239_));
 sg13g2_o21ai_1 _5038_ (.B1(_1230_),
    .Y(_1240_),
    .A1(_1237_),
    .A2(_1238_));
 sg13g2_and2_1 _5039_ (.A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[4] ),
    .B(\n352_o[11] ),
    .X(_1241_));
 sg13g2_xor2_1 _5040_ (.B(\n352_o[11] ),
    .A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[4] ),
    .X(_1242_));
 sg13g2_xor2_1 _5041_ (.B(\n352_o[12] ),
    .A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[5] ),
    .X(_1243_));
 sg13g2_and2_1 _5042_ (.A(_1242_),
    .B(_1243_),
    .X(_1244_));
 sg13g2_nor2b_1 _5043_ (.A(_1229_),
    .B_N(_1241_),
    .Y(_1245_));
 sg13g2_a221oi_1 _5044_ (.B2(_1244_),
    .C1(_1245_),
    .B1(_1240_),
    .A1(\scl_uarttx0.scl_baudrategenerator0.n6874_o[5] ),
    .Y(_1246_),
    .A2(\n352_o[12] ));
 sg13g2_o21ai_1 _5045_ (.B1(_1227_),
    .Y(_1247_),
    .A1(_1228_),
    .A2(_1246_));
 sg13g2_xor2_1 _5046_ (.B(_0822_),
    .A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[7] ),
    .X(_1248_));
 sg13g2_a21oi_2 _5047_ (.B1(_1226_),
    .Y(_1249_),
    .A2(_1248_),
    .A1(_1247_));
 sg13g2_xor2_1 _5048_ (.B(_0818_),
    .A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[9] ),
    .X(_1250_));
 sg13g2_nor2_1 _5049_ (.A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[8] ),
    .B(_0820_),
    .Y(_1251_));
 sg13g2_nor2_1 _5050_ (.A(_1221_),
    .B(_1251_),
    .Y(_1252_));
 sg13g2_nand2_1 _5051_ (.Y(_1253_),
    .A(_1250_),
    .B(_1252_));
 sg13g2_o21ai_1 _5052_ (.B1(_1225_),
    .Y(_1254_),
    .A1(_1249_),
    .A2(_1253_));
 sg13g2_o21ai_1 _5053_ (.B1(_1217_),
    .Y(_1255_),
    .A1(\scl_uarttx0.scl_baudrategenerator0.n6874_o[11] ),
    .A2(\n352_o[18] ));
 sg13g2_o21ai_1 _5054_ (.B1(_1255_),
    .Y(_1256_),
    .A1(_0766_),
    .A2(_0816_));
 sg13g2_a21o_1 _5055_ (.A2(_1254_),
    .A1(_1220_),
    .B1(_1256_),
    .X(_1257_));
 sg13g2_and2_1 _5056_ (.A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[12] ),
    .B(\n352_o[19] ),
    .X(_1258_));
 sg13g2_xor2_1 _5057_ (.B(\n352_o[19] ),
    .A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[12] ),
    .X(_1259_));
 sg13g2_inv_1 _5058_ (.Y(_1260_),
    .A(_1259_));
 sg13g2_xnor2_1 _5059_ (.Y(_1261_),
    .A(_1257_),
    .B(_1259_));
 sg13g2_inv_1 _5060_ (.Y(_1262_),
    .A(_1261_));
 sg13g2_o21ai_1 _5061_ (.B1(_1222_),
    .Y(_1263_),
    .A1(_1249_),
    .A2(_1251_));
 sg13g2_xor2_1 _5062_ (.B(_1263_),
    .A(_1250_),
    .X(_1264_));
 sg13g2_xor2_1 _5063_ (.B(_1254_),
    .A(_1218_),
    .X(_1265_));
 sg13g2_xnor2_1 _5064_ (.Y(_1266_),
    .A(_1249_),
    .B(_1252_));
 sg13g2_xnor2_1 _5065_ (.Y(_1267_),
    .A(_1247_),
    .B(_1248_));
 sg13g2_xnor2_1 _5066_ (.Y(_1268_),
    .A(_1228_),
    .B(_1246_));
 sg13g2_xnor2_1 _5067_ (.Y(_1269_),
    .A(_1233_),
    .B(_1234_));
 sg13g2_xnor2_1 _5068_ (.Y(_1270_),
    .A(_1235_),
    .B(_1236_));
 sg13g2_nor2_1 _5069_ (.A(_1269_),
    .B(_1270_),
    .Y(_1271_));
 sg13g2_xnor2_1 _5070_ (.Y(_1272_),
    .A(_1237_),
    .B(_1239_));
 sg13g2_nor2_1 _5071_ (.A(_1271_),
    .B(_1272_),
    .Y(_1273_));
 sg13g2_xnor2_1 _5072_ (.Y(_1274_),
    .A(_1240_),
    .B(_1242_));
 sg13g2_a21oi_1 _5073_ (.A1(_1240_),
    .A2(_1242_),
    .Y(_1275_),
    .B1(_1241_));
 sg13g2_xor2_1 _5074_ (.B(_1275_),
    .A(_1243_),
    .X(_1276_));
 sg13g2_nor2_1 _5075_ (.A(_1274_),
    .B(_1276_),
    .Y(_1277_));
 sg13g2_nor3_2 _5076_ (.A(_1273_),
    .B(_1274_),
    .C(_1276_),
    .Y(_1278_));
 sg13g2_nand2_1 _5077_ (.Y(_1279_),
    .A(_1267_),
    .B(_1268_));
 sg13g2_nor3_1 _5078_ (.A(_1266_),
    .B(_1278_),
    .C(_1279_),
    .Y(_1280_));
 sg13g2_or3_1 _5079_ (.A(_1266_),
    .B(_1278_),
    .C(_1279_),
    .X(_1281_));
 sg13g2_nand3_1 _5080_ (.B(_1265_),
    .C(_1281_),
    .A(_1264_),
    .Y(_1282_));
 sg13g2_a21oi_1 _5081_ (.A1(_1218_),
    .A2(_1254_),
    .Y(_1283_),
    .B1(_1217_));
 sg13g2_xor2_1 _5082_ (.B(_1283_),
    .A(_1219_),
    .X(_1284_));
 sg13g2_nor2_1 _5083_ (.A(_1282_),
    .B(_1284_),
    .Y(_1285_));
 sg13g2_nor2_1 _5084_ (.A(_1262_),
    .B(_1285_),
    .Y(_1286_));
 sg13g2_o21ai_1 _5085_ (.B1(_1261_),
    .Y(_1287_),
    .A1(_1282_),
    .A2(_1284_));
 sg13g2_and2_1 _5086_ (.A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[13] ),
    .B(\n352_o[20] ),
    .X(_1288_));
 sg13g2_or2_1 _5087_ (.X(_1289_),
    .B(\n352_o[20] ),
    .A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[13] ));
 sg13g2_nand2b_1 _5088_ (.Y(_1290_),
    .B(_1289_),
    .A_N(_1288_));
 sg13g2_a21oi_1 _5089_ (.A1(_1257_),
    .A2(_1259_),
    .Y(_1291_),
    .B1(_1258_));
 sg13g2_xnor2_1 _5090_ (.Y(_1292_),
    .A(_1290_),
    .B(_1291_));
 sg13g2_nand2_1 _5091_ (.Y(_1293_),
    .A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[14] ),
    .B(\n352_o[21] ));
 sg13g2_xor2_1 _5092_ (.B(\n352_o[21] ),
    .A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[14] ),
    .X(_1294_));
 sg13g2_inv_1 _5093_ (.Y(_1295_),
    .A(_1294_));
 sg13g2_nor2_1 _5094_ (.A(_1260_),
    .B(_1290_),
    .Y(_1296_));
 sg13g2_a221oi_1 _5095_ (.B2(_1257_),
    .C1(_1288_),
    .B1(_1296_),
    .A1(_1258_),
    .Y(_1297_),
    .A2(_1289_));
 sg13g2_xnor2_1 _5096_ (.Y(_1298_),
    .A(_1294_),
    .B(_1297_));
 sg13g2_nor2b_1 _5097_ (.A(_1292_),
    .B_N(_1298_),
    .Y(_1299_));
 sg13g2_nand3b_1 _5098_ (.B(_1298_),
    .C(_1287_),
    .Y(_1300_),
    .A_N(_1292_));
 sg13g2_nor2_1 _5099_ (.A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[15] ),
    .B(\n352_o[22] ),
    .Y(_1301_));
 sg13g2_inv_1 _5100_ (.Y(_1302_),
    .A(_1301_));
 sg13g2_xor2_1 _5101_ (.B(\n352_o[22] ),
    .A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[15] ),
    .X(_1303_));
 sg13g2_o21ai_1 _5102_ (.B1(_1293_),
    .Y(_1304_),
    .A1(_1295_),
    .A2(_1297_));
 sg13g2_xnor2_1 _5103_ (.Y(_1305_),
    .A(_1303_),
    .B(_1304_));
 sg13g2_and2_1 _5104_ (.A(_1300_),
    .B(_1305_),
    .X(_1306_));
 sg13g2_a22oi_1 _5105_ (.Y(_1307_),
    .B1(\n352_o[21] ),
    .B2(\scl_uarttx0.scl_baudrategenerator0.n6874_o[14] ),
    .A2(\n352_o[22] ),
    .A1(\scl_uarttx0.scl_baudrategenerator0.n6874_o[15] ));
 sg13g2_o21ai_1 _5106_ (.B1(_1307_),
    .Y(_1308_),
    .A1(_1295_),
    .A2(_1297_));
 sg13g2_xnor2_1 _5107_ (.Y(_1309_),
    .A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[16] ),
    .B(\n352_o[23] ));
 sg13g2_inv_1 _5108_ (.Y(_1310_),
    .A(_1309_));
 sg13g2_and3_1 _5109_ (.X(_1311_),
    .A(_1302_),
    .B(_1308_),
    .C(_1310_));
 sg13g2_nand3_1 _5110_ (.B(_1308_),
    .C(_1309_),
    .A(_1302_),
    .Y(_1312_));
 sg13g2_a21o_1 _5111_ (.A2(_1308_),
    .A1(_1302_),
    .B1(_1309_),
    .X(_1313_));
 sg13g2_and2_1 _5112_ (.A(_1312_),
    .B(_1313_),
    .X(_1314_));
 sg13g2_a22oi_1 _5113_ (.Y(_1315_),
    .B1(_1312_),
    .B2(_1313_),
    .A2(_1305_),
    .A1(_1300_));
 sg13g2_a21o_2 _5114_ (.A2(\n352_o[23] ),
    .A1(\scl_uarttx0.scl_baudrategenerator0.n6874_o[16] ),
    .B1(_1311_),
    .X(_1316_));
 sg13g2_nor2_2 _5115_ (.A(_1315_),
    .B(_1316_),
    .Y(_1317_));
 sg13g2_nor3_2 _5116_ (.A(n346_q),
    .B(s_m_popempty),
    .C(_1317_),
    .Y(_1318_));
 sg13g2_and2_1 _5117_ (.A(net1737),
    .B(_1318_),
    .X(_1319_));
 sg13g2_nand3_1 _5118_ (.B(\scl_uarttx0.n2856_o[1] ),
    .C(\scl_uarttx0.n2856_o[2] ),
    .A(\scl_uarttx0.n2856_o[0] ),
    .Y(_1320_));
 sg13g2_nand3_1 _5119_ (.B(net1642),
    .C(_1319_),
    .A(\scl_uarttx0.n2856_o[1] ),
    .Y(_1321_));
 sg13g2_nor2b_1 _5120_ (.A(\scl_uarttx0.n2856_o[1] ),
    .B_N(\scl_uarttx0.n2856_o[0] ),
    .Y(_1322_));
 sg13g2_o21ai_1 _5121_ (.B1(\scl_uarttx0.n2856_o[0] ),
    .Y(_1323_),
    .A1(\scl_uarttx0.n2856_o[1] ),
    .A2(_0767_));
 sg13g2_nor2b_1 _5122_ (.A(_1323_),
    .B_N(_1318_),
    .Y(_1324_));
 sg13g2_o21ai_1 _5123_ (.B1(_1321_),
    .Y(_0176_),
    .A1(net1642),
    .A2(_1324_));
 sg13g2_nor2_1 _5124_ (.A(_0767_),
    .B(_1320_),
    .Y(_1325_));
 sg13g2_o21ai_1 _5125_ (.B1(_1325_),
    .Y(_1326_),
    .A1(_1315_),
    .A2(_1316_));
 sg13g2_nand3b_1 _5126_ (.B(_1076_),
    .C(\scl_bitbangengine0.n5898_q[3] ),
    .Y(_1327_),
    .A_N(\scl_bitbangengine0.n5898_q[2] ));
 sg13g2_nand3b_1 _5127_ (.B(\scl_bitbangengine0.n5898_q[2] ),
    .C(_1073_),
    .Y(_1328_),
    .A_N(\scl_bitbangengine0.n5898_q[3] ));
 sg13g2_nand4_1 _5128_ (.B(_1200_),
    .C(_1327_),
    .A(n346_q),
    .Y(_1329_),
    .D(_1328_));
 sg13g2_nand2b_1 _5129_ (.Y(_1330_),
    .B(_1077_),
    .A_N(_1092_));
 sg13g2_a21oi_1 _5130_ (.A1(_1103_),
    .A2(_1177_),
    .Y(_1331_),
    .B1(_1330_));
 sg13g2_nor3_1 _5131_ (.A(net1406),
    .B(_1329_),
    .C(_1331_),
    .Y(_1332_));
 sg13g2_xnor2_1 _5132_ (.Y(_1333_),
    .A(\scl_bitbangengine0.n5905_q ),
    .B(\scl_bitbangengine0.s_m_value[0] ));
 sg13g2_nor3_1 _5133_ (.A(_0120_),
    .B(_0768_),
    .C(_1333_),
    .Y(_1334_));
 sg13g2_or2_1 _5134_ (.X(_1335_),
    .B(_1334_),
    .A(_1189_));
 sg13g2_nor2_2 _5135_ (.A(_0733_),
    .B(_1211_),
    .Y(_1336_));
 sg13g2_nand2_2 _5136_ (.Y(_1337_),
    .A(\scl_bitbangengine0.n5911_q ),
    .B(_1210_));
 sg13g2_nand2_1 _5137_ (.Y(_1338_),
    .A(_1335_),
    .B(_1336_));
 sg13g2_a221oi_1 _5138_ (.B2(_1338_),
    .C1(s_m_popempty),
    .B1(_1332_),
    .A1(_0724_),
    .Y(_1339_),
    .A2(_1326_));
 sg13g2_xnor2_1 _5139_ (.Y(_1340_),
    .A(\scl_fifo0.n2737_o[1] ),
    .B(\scl_fifo0.n2737_o[0] ));
 sg13g2_mux2_2 _5140_ (.A0(_0118_),
    .A1(_1340_),
    .S(_1339_),
    .X(_1341_));
 sg13g2_inv_1 _5141_ (.Y(\scl_fifo0.n2697_o[1] ),
    .A(net1235));
 sg13g2_xnor2_1 _5142_ (.Y(_1342_),
    .A(\scl_fifo0.n2737_o[0] ),
    .B(_1339_));
 sg13g2_inv_2 _5143_ (.Y(\scl_fifo0.n2697_o[0] ),
    .A(net1228));
 sg13g2_xnor2_1 _5144_ (.Y(_1343_),
    .A(_0711_),
    .B(net1237));
 sg13g2_xnor2_1 _5145_ (.Y(_1344_),
    .A(net1641),
    .B(\scl_fifo0.n2697_o[0] ));
 sg13g2_nand3_1 _5146_ (.B(\scl_fifo0.n2737_o[0] ),
    .C(_1339_),
    .A(\scl_fifo0.n2737_o[1] ),
    .Y(_1345_));
 sg13g2_nor2_1 _5147_ (.A(_0127_),
    .B(_1345_),
    .Y(_1346_));
 sg13g2_xnor2_1 _5148_ (.Y(_1347_),
    .A(_0127_),
    .B(_1345_));
 sg13g2_inv_1 _5149_ (.Y(\scl_fifo0.n2697_o[2] ),
    .A(net1189));
 sg13g2_xnor2_1 _5150_ (.Y(_1348_),
    .A(_0121_),
    .B(net1180));
 sg13g2_nor3_1 _5151_ (.A(_1343_),
    .B(_1344_),
    .C(_1348_),
    .Y(_1349_));
 sg13g2_xor2_1 _5152_ (.B(_1346_),
    .A(_0128_),
    .X(_1350_));
 sg13g2_inv_1 _5153_ (.Y(\scl_fifo0.n2697_o[3] ),
    .A(_1350_));
 sg13g2_xnor2_1 _5154_ (.Y(_1351_),
    .A(net1836),
    .B(_1350_));
 sg13g2_nand2_1 _5155_ (.Y(_1352_),
    .A(\scl_fifo0.n2737_o[2] ),
    .B(\scl_fifo0.n2737_o[3] ));
 sg13g2_nor2_1 _5156_ (.A(_1345_),
    .B(_1352_),
    .Y(_1353_));
 sg13g2_xnor2_1 _5157_ (.Y(\scl_fifo0.n2697_o[4] ),
    .A(net1026),
    .B(_1353_));
 sg13g2_xnor2_1 _5158_ (.Y(_1354_),
    .A(net1058),
    .B(\scl_fifo0.n2697_o[4] ));
 sg13g2_nand3_1 _5159_ (.B(_1351_),
    .C(_1354_),
    .A(_1349_),
    .Y(_0175_));
 sg13g2_nor2_2 _5160_ (.A(net1764),
    .B(_0787_),
    .Y(_1355_));
 sg13g2_inv_1 _5161_ (.Y(s_m_status_rxactive),
    .A(_1355_));
 sg13g2_nand2_1 _5162_ (.Y(_1356_),
    .A(\usbfunction0.n2634_q[3] ),
    .B(_0950_));
 sg13g2_nor3_1 _5163_ (.A(_0701_),
    .B(\usbfunction0.n2634_q[2] ),
    .C(_1356_),
    .Y(_1357_));
 sg13g2_and3_1 _5164_ (.X(_1358_),
    .A(\usbfunction0.n2634_q[1] ),
    .B(\usbfunction0.n2634_q[0] ),
    .C(_1016_));
 sg13g2_and2_2 _5165_ (.A(\usbfunction0.n2628_q ),
    .B(_1358_),
    .X(_1359_));
 sg13g2_or3_1 _5166_ (.A(_0808_),
    .B(_1357_),
    .C(_1359_),
    .X(_1360_));
 sg13g2_nor2_2 _5167_ (.A(_1014_),
    .B(_1017_),
    .Y(_1361_));
 sg13g2_nand2b_1 _5168_ (.Y(_1362_),
    .B(_1018_),
    .A_N(_1014_));
 sg13g2_o21ai_1 _5169_ (.B1(_1362_),
    .Y(_1363_),
    .A1(_1026_),
    .A2(_1027_));
 sg13g2_nor2_1 _5170_ (.A(_1360_),
    .B(_1363_),
    .Y(_1364_));
 sg13g2_and2_2 _5171_ (.A(\usbfunction0.n2631_q ),
    .B(\usbfunction0.n2630_q ),
    .X(_1365_));
 sg13g2_nand2_2 _5172_ (.Y(_1366_),
    .A(net1570),
    .B(\usbfunction0.n2630_q ));
 sg13g2_nand2_1 _5173_ (.Y(_1367_),
    .A(_1358_),
    .B(_1365_));
 sg13g2_nand2_1 _5174_ (.Y(_1368_),
    .A(\s_m_pushdata_endpoint[0] ),
    .B(net1381));
 sg13g2_nor4_1 _5175_ (.A(_0701_),
    .B(\usbfunction0.n2634_q[1] ),
    .C(_0702_),
    .D(_0806_),
    .Y(_1369_));
 sg13g2_nor2_1 _5176_ (.A(\usbfunction0.n1359_o[1] ),
    .B(\usbfunction0.n1359_o[0] ),
    .Y(_1370_));
 sg13g2_nand4_1 _5177_ (.B(_0951_),
    .C(_1369_),
    .A(\usbfunction0.n1581_o[1] ),
    .Y(_1371_),
    .D(_1370_));
 sg13g2_inv_2 _5178_ (.Y(_1372_),
    .A(net1415));
 sg13g2_nor3_1 _5179_ (.A(\s_m_packetdata_2_rewired[6] ),
    .B(\s_m_packetdata_2_rewired[5] ),
    .C(_1371_),
    .Y(_1373_));
 sg13g2_nor4_2 _5180_ (.A(\s_m_packetdata_2_rewired[1] ),
    .B(\s_m_packetdata_2_rewired[3] ),
    .C(\s_m_packetdata_2_rewired[2] ),
    .Y(_1374_),
    .D(\s_m_packetdata_2_rewired[4] ));
 sg13g2_nand3_1 _5181_ (.B(_1373_),
    .C(_1374_),
    .A(_0723_),
    .Y(_1375_));
 sg13g2_nor3_1 _5182_ (.A(\s_m_packetdata_2_rewired[15] ),
    .B(\s_m_packetdata_2_rewired[14] ),
    .C(\s_m_packetdata_2_rewired[12] ),
    .Y(_1376_));
 sg13g2_nor2b_2 _5183_ (.A(\s_m_packetdata_2_rewired[13] ),
    .B_N(_1376_),
    .Y(_1377_));
 sg13g2_nand3b_1 _5184_ (.B(_1377_),
    .C(\s_m_packetdata_2_rewired[11] ),
    .Y(_1378_),
    .A_N(\s_m_packetdata_2_rewired[10] ));
 sg13g2_or2_1 _5185_ (.X(_1379_),
    .B(_1378_),
    .A(_1375_));
 sg13g2_nor4_1 _5186_ (.A(\s_m_packetdata_2_rewired[23] ),
    .B(\s_m_packetdata_2_rewired[22] ),
    .C(\s_m_packetdata_2_rewired[21] ),
    .D(\s_m_packetdata_2_rewired[20] ),
    .Y(_1380_));
 sg13g2_nor2_1 _5187_ (.A(\s_m_packetdata_2_rewired[19] ),
    .B(\s_m_packetdata_2_rewired[18] ),
    .Y(_1381_));
 sg13g2_nor3_1 _5188_ (.A(\s_m_packetdata_2_rewired[19] ),
    .B(\s_m_packetdata_2_rewired[18] ),
    .C(s_m_packetdata_2_bit_17),
    .Y(_1382_));
 sg13g2_nand3_1 _5189_ (.B(_1380_),
    .C(_1382_),
    .A(s_m_packetdata_2_bit_16),
    .Y(_1383_));
 sg13g2_nand2b_2 _5190_ (.Y(_1384_),
    .B(net1487),
    .A_N(net1486));
 sg13g2_nor3_2 _5191_ (.A(\usbfunction0.n2481_o[17] ),
    .B(\usbfunction0.n2481_o[19] ),
    .C(\usbfunction0.n2481_o[18] ),
    .Y(_1385_));
 sg13g2_nor2b_1 _5192_ (.A(\usbfunction0.n2481_o[16] ),
    .B_N(_1385_),
    .Y(_1386_));
 sg13g2_nor4_2 _5193_ (.A(\usbfunction0.n2481_o[21] ),
    .B(\usbfunction0.n2481_o[20] ),
    .C(\usbfunction0.n2481_o[23] ),
    .Y(_1387_),
    .D(\usbfunction0.n2481_o[22] ));
 sg13g2_inv_1 _5194_ (.Y(_1388_),
    .A(_1387_));
 sg13g2_nand2_1 _5195_ (.Y(_1389_),
    .A(_1386_),
    .B(_1387_));
 sg13g2_nor4_1 _5196_ (.A(_1379_),
    .B(_1383_),
    .C(_1384_),
    .D(_1389_),
    .Y(_1390_));
 sg13g2_nor2_1 _5197_ (.A(_0053_),
    .B(net1380),
    .Y(_1391_));
 sg13g2_nor2_1 _5198_ (.A(\s_m_packetdata_2_rewired[11] ),
    .B(\s_m_packetdata_2_rewired[10] ),
    .Y(_1392_));
 sg13g2_nand3_1 _5199_ (.B(_1377_),
    .C(_1392_),
    .A(_1373_),
    .Y(_1393_));
 sg13g2_nor2b_1 _5200_ (.A(s_m_packetdata_2_bit_16),
    .B_N(_1380_),
    .Y(_1394_));
 sg13g2_and2_2 _5201_ (.A(_1382_),
    .B(_1394_),
    .X(_1395_));
 sg13g2_nand2_1 _5202_ (.Y(_1396_),
    .A(_1387_),
    .B(_1395_));
 sg13g2_nand2b_1 _5203_ (.Y(_1397_),
    .B(_1395_),
    .A_N(_1389_));
 sg13g2_nor3_1 _5204_ (.A(_1384_),
    .B(_1393_),
    .C(_1397_),
    .Y(_1398_));
 sg13g2_nand2_1 _5205_ (.Y(_1399_),
    .A(\usbfunction0.n2098_o ),
    .B(_1398_));
 sg13g2_inv_1 _5206_ (.Y(_1400_),
    .A(net1376));
 sg13g2_nor2b_2 _5207_ (.A(net1482),
    .B_N(net1483),
    .Y(_1401_));
 sg13g2_nand3_1 _5208_ (.B(net1484),
    .C(_1401_),
    .A(net1485),
    .Y(_1402_));
 sg13g2_nand3b_1 _5209_ (.B(_1386_),
    .C(_1387_),
    .Y(_1403_),
    .A_N(_1384_));
 sg13g2_nor3_1 _5210_ (.A(\s_m_packetdata_2_rewired[6] ),
    .B(\s_m_packetdata_2_rewired[5] ),
    .C(_1371_),
    .Y(_1404_));
 sg13g2_nand3_1 _5211_ (.B(_1374_),
    .C(_1404_),
    .A(_0723_),
    .Y(_1405_));
 sg13g2_nor4_1 _5212_ (.A(_1378_),
    .B(_1383_),
    .C(_1403_),
    .D(_1405_),
    .Y(_1406_));
 sg13g2_nand4_1 _5213_ (.B(_1392_),
    .C(_1395_),
    .A(_1377_),
    .Y(_1407_),
    .D(_1404_));
 sg13g2_o21ai_1 _5214_ (.B1(_1391_),
    .Y(_1408_),
    .A1(net1377),
    .A2(_1402_));
 sg13g2_nor2_2 _5215_ (.A(\s_m_pushdata_endpoint[0] ),
    .B(net1381),
    .Y(_1409_));
 sg13g2_or2_1 _5216_ (.X(_1410_),
    .B(net1381),
    .A(\s_m_pushdata_endpoint[0] ));
 sg13g2_nor2_1 _5217_ (.A(_0050_),
    .B(net1378),
    .Y(_1411_));
 sg13g2_nor2_2 _5218_ (.A(net1485),
    .B(net1484),
    .Y(_1412_));
 sg13g2_nand2_1 _5219_ (.Y(_1413_),
    .A(_1401_),
    .B(_1412_));
 sg13g2_o21ai_1 _5220_ (.B1(_1411_),
    .Y(_1414_),
    .A1(net1375),
    .A2(_1413_));
 sg13g2_nor2_1 _5221_ (.A(_0051_),
    .B(net1378),
    .Y(_1415_));
 sg13g2_nor2b_2 _5222_ (.A(net1484),
    .B_N(net1485),
    .Y(_1416_));
 sg13g2_nand2_1 _5223_ (.Y(_1417_),
    .A(_1401_),
    .B(_1416_));
 sg13g2_o21ai_1 _5224_ (.B1(_1415_),
    .Y(_1418_),
    .A1(net1375),
    .A2(_1417_));
 sg13g2_nand2_1 _5225_ (.Y(_1419_),
    .A(_1003_),
    .B(net1381));
 sg13g2_nor2_1 _5226_ (.A(_0052_),
    .B(net1378),
    .Y(_1420_));
 sg13g2_nor2b_2 _5227_ (.A(net1485),
    .B_N(net1484),
    .Y(_1421_));
 sg13g2_nand2_1 _5228_ (.Y(_1422_),
    .A(_1401_),
    .B(_1421_));
 sg13g2_o21ai_1 _5229_ (.B1(_1420_),
    .Y(_1423_),
    .A1(net1375),
    .A2(_1422_));
 sg13g2_mux4_1 _5230_ (.S0(\s_m_pushdata_endpoint[0] ),
    .A0(_1414_),
    .A1(_1418_),
    .A2(_1423_),
    .A3(_1408_),
    .S1(net1381),
    .X(_1424_));
 sg13g2_nor2_1 _5231_ (.A(\s_m_pushdata_endpoint[3] ),
    .B(_1424_),
    .Y(_1425_));
 sg13g2_nor2_1 _5232_ (.A(_0060_),
    .B(net1378),
    .Y(_1426_));
 sg13g2_nand3_1 _5233_ (.B(net1482),
    .C(_1421_),
    .A(net1483),
    .Y(_1427_));
 sg13g2_o21ai_1 _5234_ (.B1(_1426_),
    .Y(_1428_),
    .A1(net1375),
    .A2(_1427_));
 sg13g2_nor2_1 _5235_ (.A(_1419_),
    .B(_1428_),
    .Y(_1429_));
 sg13g2_nand3_1 _5236_ (.B(net1482),
    .C(_1416_),
    .A(net1483),
    .Y(_1430_));
 sg13g2_nor2_1 _5237_ (.A(net1375),
    .B(_1430_),
    .Y(_1431_));
 sg13g2_nor3_2 _5238_ (.A(_0059_),
    .B(net1378),
    .C(_1431_),
    .Y(_1432_));
 sg13g2_o21ai_1 _5239_ (.B1(\s_m_pushdata_endpoint[0] ),
    .Y(_1433_),
    .A1(net1381),
    .A2(_1432_));
 sg13g2_nor2_1 _5240_ (.A(_0058_),
    .B(net1380),
    .Y(_1434_));
 sg13g2_nand3_1 _5241_ (.B(net1482),
    .C(_1412_),
    .A(net1483),
    .Y(_1435_));
 sg13g2_o21ai_1 _5242_ (.B1(_1434_),
    .Y(_1436_),
    .A1(net1377),
    .A2(_1435_));
 sg13g2_nor2_1 _5243_ (.A(_1410_),
    .B(_1436_),
    .Y(_1437_));
 sg13g2_nor2_1 _5244_ (.A(_1429_),
    .B(_1437_),
    .Y(_1438_));
 sg13g2_nor2_2 _5245_ (.A(net1483),
    .B(net1482),
    .Y(_1439_));
 sg13g2_and2_1 _5246_ (.A(_1412_),
    .B(_1439_),
    .X(_1440_));
 sg13g2_nand2_2 _5247_ (.Y(_1441_),
    .A(_1412_),
    .B(_1439_));
 sg13g2_nand4_1 _5248_ (.B(net1484),
    .C(net1483),
    .A(net1485),
    .Y(_1442_),
    .D(net1482));
 sg13g2_nor2b_1 _5249_ (.A(_0046_),
    .B_N(_1442_),
    .Y(_1443_));
 sg13g2_nor3_1 _5250_ (.A(net1376),
    .B(_1440_),
    .C(_1443_),
    .Y(_1444_));
 sg13g2_a21oi_1 _5251_ (.A1(_1400_),
    .A2(_1441_),
    .Y(_1445_),
    .B1(\usbfunction0.n1687_o[14] ));
 sg13g2_nor3_2 _5252_ (.A(net1378),
    .B(_1444_),
    .C(_1445_),
    .Y(_1446_));
 sg13g2_o21ai_1 _5253_ (.B1(\s_m_pushdata_endpoint[3] ),
    .Y(_1447_),
    .A1(_1368_),
    .A2(_1446_));
 sg13g2_a21oi_1 _5254_ (.A1(_1433_),
    .A2(_1438_),
    .Y(_1448_),
    .B1(_1447_));
 sg13g2_o21ai_1 _5255_ (.B1(\s_m_pushdata_endpoint[2] ),
    .Y(_1449_),
    .A1(_1425_),
    .A2(_1448_));
 sg13g2_o21ai_1 _5256_ (.B1(net1841),
    .Y(_1450_),
    .A1(net1376),
    .A2(_1441_));
 sg13g2_nand2_1 _5257_ (.Y(_1451_),
    .A(_1005_),
    .B(_1409_));
 sg13g2_nor2_2 _5258_ (.A(net1384),
    .B(_1451_),
    .Y(_1452_));
 sg13g2_nand2_1 _5259_ (.Y(_1453_),
    .A(net1703),
    .B(_1452_));
 sg13g2_a21oi_1 _5260_ (.A1(net1703),
    .A2(_1452_),
    .Y(_1454_),
    .B1(_1450_));
 sg13g2_and2_1 _5261_ (.A(_1409_),
    .B(_1454_),
    .X(_1455_));
 sg13g2_nor2_1 _5262_ (.A(_0047_),
    .B(net1379),
    .Y(_1456_));
 sg13g2_nand2_1 _5263_ (.Y(_1457_),
    .A(_1416_),
    .B(_1439_));
 sg13g2_o21ai_1 _5264_ (.B1(_1456_),
    .Y(_1458_),
    .A1(net1375),
    .A2(_1457_));
 sg13g2_nor2_1 _5265_ (.A(_1004_),
    .B(_1458_),
    .Y(_1459_));
 sg13g2_nor2_1 _5266_ (.A(_0048_),
    .B(net1379),
    .Y(_1460_));
 sg13g2_nand2_1 _5267_ (.Y(_1461_),
    .A(_1421_),
    .B(_1439_));
 sg13g2_o21ai_1 _5268_ (.B1(_1460_),
    .Y(_1462_),
    .A1(net1377),
    .A2(_1461_));
 sg13g2_or2_1 _5269_ (.X(_1463_),
    .B(_1462_),
    .A(_1419_));
 sg13g2_nor2_1 _5270_ (.A(_0049_),
    .B(net1380),
    .Y(_1464_));
 sg13g2_nand3_1 _5271_ (.B(net1484),
    .C(_1439_),
    .A(net1485),
    .Y(_1465_));
 sg13g2_o21ai_1 _5272_ (.B1(_1464_),
    .Y(_1466_),
    .A1(net1377),
    .A2(_1465_));
 sg13g2_o21ai_1 _5273_ (.B1(_1463_),
    .Y(_1467_),
    .A1(_1368_),
    .A2(_1466_));
 sg13g2_nor4_1 _5274_ (.A(\s_m_pushdata_endpoint[3] ),
    .B(_1455_),
    .C(_1459_),
    .D(_1467_),
    .Y(_1468_));
 sg13g2_nor2_1 _5275_ (.A(_0057_),
    .B(net1378),
    .Y(_1469_));
 sg13g2_nor2b_2 _5276_ (.A(net1483),
    .B_N(net1482),
    .Y(_1470_));
 sg13g2_nand3_1 _5277_ (.B(net1484),
    .C(_1470_),
    .A(net1485),
    .Y(_1471_));
 sg13g2_o21ai_1 _5278_ (.B1(_1469_),
    .Y(_1472_),
    .A1(net1375),
    .A2(_1471_));
 sg13g2_nor2_1 _5279_ (.A(_1368_),
    .B(_1472_),
    .Y(_1473_));
 sg13g2_nor2_1 _5280_ (.A(_0055_),
    .B(net1379),
    .Y(_1474_));
 sg13g2_nand2_1 _5281_ (.Y(_1475_),
    .A(_1416_),
    .B(_1470_));
 sg13g2_o21ai_1 _5282_ (.B1(_1474_),
    .Y(_1476_),
    .A1(net1376),
    .A2(_1475_));
 sg13g2_nor2_1 _5283_ (.A(_1004_),
    .B(_1476_),
    .Y(_1477_));
 sg13g2_nor2_1 _5284_ (.A(_0056_),
    .B(net1378),
    .Y(_1478_));
 sg13g2_nand2_1 _5285_ (.Y(_1479_),
    .A(_1421_),
    .B(_1470_));
 sg13g2_o21ai_1 _5286_ (.B1(_1478_),
    .Y(_1480_),
    .A1(net1375),
    .A2(_1479_));
 sg13g2_nor2_1 _5287_ (.A(_1419_),
    .B(_1480_),
    .Y(_1481_));
 sg13g2_nor2_1 _5288_ (.A(_0054_),
    .B(net1380),
    .Y(_1482_));
 sg13g2_nand2_1 _5289_ (.Y(_1483_),
    .A(_1412_),
    .B(_1470_));
 sg13g2_o21ai_1 _5290_ (.B1(_1482_),
    .Y(_1484_),
    .A1(net1377),
    .A2(_1483_));
 sg13g2_o21ai_1 _5291_ (.B1(\s_m_pushdata_endpoint[3] ),
    .Y(_1485_),
    .A1(_1410_),
    .A2(_1484_));
 sg13g2_nor4_1 _5292_ (.A(_1473_),
    .B(_1477_),
    .C(_1481_),
    .D(_1485_),
    .Y(_1486_));
 sg13g2_or2_1 _5293_ (.X(_1487_),
    .B(_1486_),
    .A(\s_m_pushdata_endpoint[2] ));
 sg13g2_o21ai_1 _5294_ (.B1(_1449_),
    .Y(_1488_),
    .A1(_1468_),
    .A2(_1487_));
 sg13g2_xnor2_1 _5295_ (.Y(_1489_),
    .A(net1460),
    .B(_1488_));
 sg13g2_xor2_1 _5296_ (.B(_1488_),
    .A(net1464),
    .X(_1490_));
 sg13g2_inv_1 _5297_ (.Y(_1491_),
    .A(_1490_));
 sg13g2_nor4_1 _5298_ (.A(net1454),
    .B(net1470),
    .C(net1473),
    .D(net1853),
    .Y(_1492_));
 sg13g2_nand2b_1 _5299_ (.Y(_1493_),
    .B(_1492_),
    .A_N(_0935_));
 sg13g2_nor2_1 _5300_ (.A(_1490_),
    .B(_1493_),
    .Y(_1494_));
 sg13g2_a21oi_1 _5301_ (.A1(_1489_),
    .A2(_1494_),
    .Y(_1495_),
    .B1(_1367_));
 sg13g2_nor2b_1 _5302_ (.A(_1495_),
    .B_N(_1364_),
    .Y(_1496_));
 sg13g2_nor2b_1 _5303_ (.A(net1902),
    .B_N(\usbfunction0.n1359_o[1] ),
    .Y(_1497_));
 sg13g2_nor2b_1 _5304_ (.A(net1384),
    .B_N(_1370_),
    .Y(_1498_));
 sg13g2_and2_1 _5305_ (.A(_1452_),
    .B(_1497_),
    .X(_1499_));
 sg13g2_a221oi_1 _5306_ (.B2(_1451_),
    .C1(\usbfunction0.n2634_q[2] ),
    .B1(_1498_),
    .A1(_1452_),
    .Y(_1500_),
    .A2(_1497_));
 sg13g2_or2_1 _5307_ (.X(_1501_),
    .B(_1013_),
    .A(net622));
 sg13g2_nand3b_1 _5308_ (.B(_1451_),
    .C(_1497_),
    .Y(_1502_),
    .A_N(net1384));
 sg13g2_nand2b_1 _5309_ (.Y(_1503_),
    .B(_1501_),
    .A_N(_1502_));
 sg13g2_nor2b_1 _5310_ (.A(_1029_),
    .B_N(_1040_),
    .Y(_1504_));
 sg13g2_a22oi_1 _5311_ (.Y(_1505_),
    .B1(_1504_),
    .B2(_0693_),
    .A2(_1503_),
    .A1(_1500_));
 sg13g2_and2_1 _5312_ (.A(_1496_),
    .B(_1505_),
    .X(\usbfunction0.n2474_o[2] ));
 sg13g2_nor2_1 _5313_ (.A(\usbfunction0.n2634_q[0] ),
    .B(_1498_),
    .Y(_1506_));
 sg13g2_a21oi_1 _5314_ (.A1(_1453_),
    .A2(_1506_),
    .Y(_1507_),
    .B1(_1369_));
 sg13g2_nand2_1 _5315_ (.Y(_1508_),
    .A(_1364_),
    .B(_1507_));
 sg13g2_nor2_1 _5316_ (.A(_1495_),
    .B(_1508_),
    .Y(\usbfunction0.n2474_o[0] ));
 sg13g2_nor3_1 _5317_ (.A(net1888),
    .B(_1498_),
    .C(_1504_),
    .Y(_1509_));
 sg13g2_nor2b_1 _5318_ (.A(_1509_),
    .B_N(_1496_),
    .Y(\usbfunction0.n2474_o[1] ));
 sg13g2_nor4_1 _5319_ (.A(_1367_),
    .B(_1489_),
    .C(_1491_),
    .D(_1493_),
    .Y(_1510_));
 sg13g2_nor2_1 _5320_ (.A(net1870),
    .B(_1510_),
    .Y(_1511_));
 sg13g2_or2_1 _5321_ (.X(_1512_),
    .B(_1511_),
    .A(_1360_));
 sg13g2_inv_1 _5322_ (.Y(\usbfunction0.n2474_o[3] ),
    .A(_1512_));
 sg13g2_nand2_1 _5323_ (.Y(_1513_),
    .A(net876),
    .B(net1431));
 sg13g2_o21ai_1 _5324_ (.B1(_1513_),
    .Y(\n352_o[0] ),
    .A1(_0723_),
    .A2(net1430));
 sg13g2_mux2_1 _5325_ (.A0(\s_m_packetdata_2_rewired[1] ),
    .A1(net1070),
    .S(net1430),
    .X(\n352_o[1] ));
 sg13g2_mux2_1 _5326_ (.A0(\s_m_packetdata_2_rewired[2] ),
    .A1(net1573),
    .S(net1430),
    .X(\n352_o[2] ));
 sg13g2_mux2_1 _5327_ (.A0(\s_m_packetdata_2_rewired[3] ),
    .A1(net1100),
    .S(net1430),
    .X(\n352_o[3] ));
 sg13g2_mux2_1 _5328_ (.A0(\s_m_packetdata_2_rewired[4] ),
    .A1(net1149),
    .S(net1430),
    .X(\n352_o[4] ));
 sg13g2_mux2_1 _5329_ (.A0(\s_m_packetdata_2_rewired[5] ),
    .A1(net1082),
    .S(net1431),
    .X(\n352_o[5] ));
 sg13g2_mux2_1 _5330_ (.A0(\s_m_packetdata_2_rewired[6] ),
    .A1(net1112),
    .S(net1431),
    .X(\n352_o[6] ));
 sg13g2_a21oi_1 _5331_ (.A1(_0748_),
    .A2(net1434),
    .Y(_0024_),
    .B1(_0930_));
 sg13g2_a21oi_1 _5332_ (.A1(_0690_),
    .A2(_0923_),
    .Y(_1514_),
    .B1(_0925_));
 sg13g2_nor4_1 _5333_ (.A(_0921_),
    .B(_0924_),
    .C(\scl_uartrx0.n6047_o ),
    .D(_1514_),
    .Y(_0023_));
 sg13g2_nor3_1 _5334_ (.A(net559),
    .B(\usbfunction0.scl_usbgpiophy0.n6449_o ),
    .C(\usbfunction0.scl_usbgpiophy0.n6411_o ),
    .Y(_1515_));
 sg13g2_nand3_1 _5335_ (.B(_0796_),
    .C(_1515_),
    .A(net1386),
    .Y(_1516_));
 sg13g2_inv_1 _5336_ (.Y(_1517_),
    .A(net1368));
 sg13g2_nand4_1 _5337_ (.B(net537),
    .C(\usbfunction0.scl_usbgpiophy0.scl_extendwidth0.scl_counter0.n7984_q[2] ),
    .A(\usbfunction0.scl_usbgpiophy0.scl_extendwidth0.scl_counter0.n7984_q[1] ),
    .Y(_1518_),
    .D(_1517_));
 sg13g2_inv_1 _5338_ (.Y(\usbfunction0.s_m_rx_valid ),
    .A(net538));
 sg13g2_nor2_1 _5339_ (.A(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7654_q[1] ),
    .B(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7654_q[0] ),
    .Y(_1519_));
 sg13g2_nor3_1 _5340_ (.A(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.s_m_value[1] ),
    .B(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.s_m_value[0] ),
    .C(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.s_m_value[2] ),
    .Y(_1520_));
 sg13g2_nand3_1 _5341_ (.B(_1519_),
    .C(_1520_),
    .A(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.s_m_value[3] ),
    .Y(_1521_));
 sg13g2_nor2b_1 _5342_ (.A(_0045_),
    .B_N(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.s_m_value[2] ),
    .Y(_1522_));
 sg13g2_nor2_1 _5343_ (.A(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.s_m_value[1] ),
    .B(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.s_m_value[0] ),
    .Y(_1523_));
 sg13g2_nand3b_1 _5344_ (.B(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.s_m_value[0] ),
    .C(\usbfunction0.scl_usbgpiophy0.s_out_2[5] ),
    .Y(_1524_),
    .A_N(net1488));
 sg13g2_nor2b_1 _5345_ (.A(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.s_m_value[0] ),
    .B_N(net1488),
    .Y(_1525_));
 sg13g2_a22oi_1 _5346_ (.Y(_1526_),
    .B1(_1525_),
    .B2(\usbfunction0.scl_usbgpiophy0.s_out_2[6] ),
    .A2(_1523_),
    .A1(\usbfunction0.scl_usbgpiophy0.s_out_2[4] ));
 sg13g2_nand2_1 _5347_ (.Y(_1527_),
    .A(_1524_),
    .B(_1526_));
 sg13g2_nor2b_1 _5348_ (.A(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.s_m_value[2] ),
    .B_N(_0045_),
    .Y(_1528_));
 sg13g2_mux4_1 _5349_ (.S0(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.s_m_value[0] ),
    .A0(\usbfunction0.scl_usbgpiophy0.s_out_2[0] ),
    .A1(\usbfunction0.scl_usbgpiophy0.s_out_2[1] ),
    .A2(\usbfunction0.scl_usbgpiophy0.s_out_2[2] ),
    .A3(\usbfunction0.scl_usbgpiophy0.s_out_2[3] ),
    .S1(net1488),
    .X(_1529_));
 sg13g2_a22oi_1 _5350_ (.Y(_1530_),
    .B1(_1528_),
    .B2(_1529_),
    .A2(_1527_),
    .A1(_1522_));
 sg13g2_a21oi_1 _5351_ (.A1(_1035_),
    .A2(_1522_),
    .Y(_1531_),
    .B1(_1528_));
 sg13g2_o21ai_1 _5352_ (.B1(_1531_),
    .Y(_1532_),
    .A1(_0713_),
    .A2(\usbfunction0.scl_usbgpiophy0.s_out_2[7] ));
 sg13g2_o21ai_1 _5353_ (.B1(_1532_),
    .Y(_1533_),
    .A1(_0713_),
    .A2(_1530_));
 sg13g2_mux2_1 _5354_ (.A0(_1533_),
    .A1(net1629),
    .S(_1521_),
    .X(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7508_o ));
 sg13g2_nand2_1 _5355_ (.Y(_1534_),
    .A(net1170),
    .B(_0799_));
 sg13g2_nand2_1 _5356_ (.Y(_1535_),
    .A(net1640),
    .B(_0790_));
 sg13g2_o21ai_1 _5357_ (.B1(_1534_),
    .Y(_0028_),
    .A1(net1436),
    .A2(_1535_));
 sg13g2_o21ai_1 _5358_ (.B1(_0793_),
    .Y(_1536_),
    .A1(net1640),
    .A2(net1170));
 sg13g2_a22oi_1 _5359_ (.Y(_1537_),
    .B1(_0790_),
    .B2(\usbfunction0.scl_usbgpiophy0.n6437_o ),
    .A2(net1386),
    .A1(net1436));
 sg13g2_nand4_1 _5360_ (.B(_0795_),
    .C(_1536_),
    .A(net1023),
    .Y(_1538_),
    .D(_1537_));
 sg13g2_o21ai_1 _5361_ (.B1(_1538_),
    .Y(_0027_),
    .A1(_0791_),
    .A2(_0798_));
 sg13g2_nand2_1 _5362_ (.Y(_1539_),
    .A(net1640),
    .B(_0799_));
 sg13g2_nand3b_1 _5363_ (.B(_1535_),
    .C(_1536_),
    .Y(_1540_),
    .A_N(net1436));
 sg13g2_o21ai_1 _5364_ (.B1(_1539_),
    .Y(_0026_),
    .A1(_0795_),
    .A2(_1540_));
 sg13g2_a21o_1 _5365_ (.A2(_0931_),
    .A1(net938),
    .B1(_0932_),
    .X(_0025_));
 sg13g2_nor4_1 _5366_ (.A(net1700),
    .B(net1683),
    .C(net603),
    .D(net1671),
    .Y(_1541_));
 sg13g2_nor2_1 _5367_ (.A(net1677),
    .B(net583),
    .Y(_1542_));
 sg13g2_nor4_1 _5368_ (.A(net794),
    .B(net1754),
    .C(net1679),
    .D(net1647),
    .Y(_1543_));
 sg13g2_and3_2 _5369_ (.X(\usbfunction0.functionreset0.n6683_o ),
    .A(_1541_),
    .B(_1542_),
    .C(_1543_));
 sg13g2_and4_2 _5370_ (.A(_0721_),
    .B(net1394),
    .C(_1032_),
    .D(net1392),
    .X(_1544_));
 sg13g2_nand4_1 _5371_ (.B(net1394),
    .C(_1032_),
    .A(_0721_),
    .Y(_1545_),
    .D(net1392));
 sg13g2_xnor2_1 _5372_ (.Y(_1546_),
    .A(net1897),
    .B(net1350));
 sg13g2_nand2_1 _5373_ (.Y(_1547_),
    .A(_0085_),
    .B(net1418));
 sg13g2_o21ai_1 _5374_ (.B1(_1547_),
    .Y(_1548_),
    .A1(net1418),
    .A2(_1546_));
 sg13g2_nor2_1 _5375_ (.A(_1372_),
    .B(_1548_),
    .Y(_1549_));
 sg13g2_nand3b_1 _5376_ (.B(\s_m_packetdata_2_rewired[10] ),
    .C(_1377_),
    .Y(_1550_),
    .A_N(\s_m_packetdata_2_rewired[11] ));
 sg13g2_or2_1 _5377_ (.X(_1551_),
    .B(_1550_),
    .A(_1375_));
 sg13g2_nand2b_1 _5378_ (.Y(_1552_),
    .B(net1486),
    .A_N(net1487));
 sg13g2_nor3_1 _5379_ (.A(_1388_),
    .B(_1551_),
    .C(_1552_),
    .Y(_1553_));
 sg13g2_nor3_2 _5380_ (.A(_0722_),
    .B(\usbfunction0.n2481_o[19] ),
    .C(\usbfunction0.n2481_o[18] ),
    .Y(_1554_));
 sg13g2_nor3_2 _5381_ (.A(net1486),
    .B(net1487),
    .C(_1379_),
    .Y(_1555_));
 sg13g2_inv_1 _5382_ (.Y(_1556_),
    .A(_1555_));
 sg13g2_nor3_2 _5383_ (.A(net1486),
    .B(net1487),
    .C(_1379_),
    .Y(_1557_));
 sg13g2_or2_1 _5384_ (.X(_1558_),
    .B(_1552_),
    .A(_1551_));
 sg13g2_nor2_1 _5385_ (.A(_1396_),
    .B(_1558_),
    .Y(_1559_));
 sg13g2_and2_2 _5386_ (.A(_1554_),
    .B(_1559_),
    .X(_1560_));
 sg13g2_nor2b_2 _5387_ (.A(\usbfunction0.n2481_o[16] ),
    .B_N(_1560_),
    .Y(_1561_));
 sg13g2_nor3_1 _5388_ (.A(_1549_),
    .B(_1557_),
    .C(_1561_),
    .Y(_1562_));
 sg13g2_inv_1 _5389_ (.Y(_1563_),
    .A(_1562_));
 sg13g2_nor3_1 _5390_ (.A(\usbfunction0.n2650_q[0] ),
    .B(\usbfunction0.n2650_q[1] ),
    .C(net1350),
    .Y(_1564_));
 sg13g2_nor4_1 _5391_ (.A(\usbfunction0.n2650_q[0] ),
    .B(\usbfunction0.n2650_q[1] ),
    .C(\usbfunction0.n2650_q[2] ),
    .D(net1350),
    .Y(_1565_));
 sg13g2_nor2_1 _5392_ (.A(_1020_),
    .B(net1350),
    .Y(_1566_));
 sg13g2_xor2_1 _5393_ (.B(_1566_),
    .A(_0090_),
    .X(_1567_));
 sg13g2_xnor2_1 _5394_ (.Y(_1568_),
    .A(net1840),
    .B(_1566_));
 sg13g2_o21ai_1 _5395_ (.B1(net1415),
    .Y(_1569_),
    .A1(\usbfunction0.n2652_q[4] ),
    .A2(net1423));
 sg13g2_a21oi_1 _5396_ (.A1(net1423),
    .A2(_1567_),
    .Y(_1570_),
    .B1(_1569_));
 sg13g2_nand4_1 _5397_ (.B(_1385_),
    .C(_1395_),
    .A(\usbfunction0.n2481_o[16] ),
    .Y(_1571_),
    .D(_1553_));
 sg13g2_nand3_1 _5398_ (.B(_1387_),
    .C(_1554_),
    .A(\usbfunction0.n2481_o[16] ),
    .Y(_1572_));
 sg13g2_nor3_2 _5399_ (.A(_1383_),
    .B(_1558_),
    .C(_1572_),
    .Y(_1573_));
 sg13g2_and3_2 _5400_ (.X(_1574_),
    .A(\usbfunction0.n2481_o[16] ),
    .B(_1385_),
    .C(_1559_));
 sg13g2_or3_2 _5401_ (.A(_1570_),
    .B(_1573_),
    .C(_1574_),
    .X(_1575_));
 sg13g2_inv_1 _5402_ (.Y(_1576_),
    .A(_1575_));
 sg13g2_xnor2_1 _5403_ (.Y(_1577_),
    .A(_0699_),
    .B(_1575_));
 sg13g2_a21oi_1 _5404_ (.A1(_1022_),
    .A2(_1544_),
    .Y(_1578_),
    .B1(_0760_));
 sg13g2_nor3_1 _5405_ (.A(net1865),
    .B(_1023_),
    .C(net1350),
    .Y(_1579_));
 sg13g2_nor2_1 _5406_ (.A(_1578_),
    .B(_1579_),
    .Y(_1580_));
 sg13g2_o21ai_1 _5407_ (.B1(net1422),
    .Y(_1581_),
    .A1(_1578_),
    .A2(_1579_));
 sg13g2_a21oi_1 _5408_ (.A1(_0761_),
    .A2(net1420),
    .Y(_1582_),
    .B1(_1372_));
 sg13g2_a21o_1 _5409_ (.A2(_1582_),
    .A1(_1581_),
    .B1(_1561_),
    .X(_1583_));
 sg13g2_xor2_1 _5410_ (.B(_1583_),
    .A(\usbfunction0.n1583_o[6] ),
    .X(_1584_));
 sg13g2_nand2_1 _5411_ (.Y(_1585_),
    .A(_1024_),
    .B(_1544_));
 sg13g2_xor2_1 _5412_ (.B(_1585_),
    .A(net1812),
    .X(_1586_));
 sg13g2_xnor2_1 _5413_ (.Y(_1587_),
    .A(net1812),
    .B(_1585_));
 sg13g2_o21ai_1 _5414_ (.B1(net1415),
    .Y(_1588_),
    .A1(net1881),
    .A2(net1422));
 sg13g2_a21oi_1 _5415_ (.A1(net1422),
    .A2(_1587_),
    .Y(_1589_),
    .B1(_1588_));
 sg13g2_inv_1 _5416_ (.Y(_1590_),
    .A(_1589_));
 sg13g2_and2_1 _5417_ (.A(_0086_),
    .B(_1589_),
    .X(_1591_));
 sg13g2_nor2_1 _5418_ (.A(_0086_),
    .B(_1589_),
    .Y(_1592_));
 sg13g2_or3_1 _5419_ (.A(_1584_),
    .B(_1591_),
    .C(_1592_),
    .X(_1593_));
 sg13g2_nand2_1 _5420_ (.Y(_1594_),
    .A(_1021_),
    .B(_1544_));
 sg13g2_xor2_1 _5421_ (.B(_1594_),
    .A(net1838),
    .X(_1595_));
 sg13g2_xnor2_1 _5422_ (.Y(_1596_),
    .A(_0089_),
    .B(_1594_));
 sg13g2_o21ai_1 _5423_ (.B1(net1415),
    .Y(_1597_),
    .A1(\usbfunction0.n2652_q[5] ),
    .A2(net1422));
 sg13g2_a21oi_1 _5424_ (.A1(net1423),
    .A2(_1596_),
    .Y(_1598_),
    .B1(_1597_));
 sg13g2_nand3_1 _5425_ (.B(_1381_),
    .C(_1394_),
    .A(s_m_packetdata_2_bit_17),
    .Y(_1599_));
 sg13g2_nor3_2 _5426_ (.A(_1558_),
    .B(_1572_),
    .C(_1599_),
    .Y(_1600_));
 sg13g2_or2_1 _5427_ (.X(_1601_),
    .B(_1600_),
    .A(_1598_));
 sg13g2_xor2_1 _5428_ (.B(_1601_),
    .A(\usbfunction0.n1583_o[5] ),
    .X(_1602_));
 sg13g2_xnor2_1 _5429_ (.Y(_1603_),
    .A(net1822),
    .B(_1565_));
 sg13g2_o21ai_1 _5430_ (.B1(net1415),
    .Y(_1604_),
    .A1(net1418),
    .A2(_1603_));
 sg13g2_a21oi_1 _5431_ (.A1(_0762_),
    .A2(net1418),
    .Y(_1605_),
    .B1(_1604_));
 sg13g2_inv_1 _5432_ (.Y(_1606_),
    .A(_1605_));
 sg13g2_nand2_1 _5433_ (.Y(_1607_),
    .A(_0698_),
    .B(_1606_));
 sg13g2_xnor2_1 _5434_ (.Y(_1608_),
    .A(net1799),
    .B(_1564_));
 sg13g2_nor2_1 _5435_ (.A(net1418),
    .B(_1608_),
    .Y(_1609_));
 sg13g2_o21ai_1 _5436_ (.B1(net1415),
    .Y(_1610_),
    .A1(\usbfunction0.n2652_q[2] ),
    .A2(net1423));
 sg13g2_nor2_1 _5437_ (.A(_1609_),
    .B(_1610_),
    .Y(_1611_));
 sg13g2_nand2_1 _5438_ (.Y(_1612_),
    .A(\usbfunction0.n2481_o[16] ),
    .B(_1560_));
 sg13g2_inv_1 _5439_ (.Y(_1613_),
    .A(_1612_));
 sg13g2_nor2_2 _5440_ (.A(_1611_),
    .B(_1613_),
    .Y(_1614_));
 sg13g2_inv_1 _5441_ (.Y(_1615_),
    .A(_1614_));
 sg13g2_xor2_1 _5442_ (.B(_1614_),
    .A(\usbfunction0.n1583_o[2] ),
    .X(_1616_));
 sg13g2_nand2_1 _5443_ (.Y(_1617_),
    .A(_0032_),
    .B(_1605_));
 sg13g2_nor3_1 _5444_ (.A(_1577_),
    .B(_1593_),
    .C(_1602_),
    .Y(_1618_));
 sg13g2_nand4_1 _5445_ (.B(_1616_),
    .C(_1617_),
    .A(_1607_),
    .Y(_1619_),
    .D(_1618_));
 sg13g2_xnor2_1 _5446_ (.Y(_1620_),
    .A(\usbfunction0.n2650_q[0] ),
    .B(\usbfunction0.n2650_q[1] ));
 sg13g2_nand2_1 _5447_ (.Y(_1621_),
    .A(_1544_),
    .B(_1620_));
 sg13g2_o21ai_1 _5448_ (.B1(_1621_),
    .Y(_1622_),
    .A1(net1777),
    .A2(_1544_));
 sg13g2_nand2_1 _5449_ (.Y(_1623_),
    .A(_0093_),
    .B(net1418));
 sg13g2_o21ai_1 _5450_ (.B1(_1623_),
    .Y(_1624_),
    .A1(net1418),
    .A2(_1622_));
 sg13g2_nor2_1 _5451_ (.A(_1372_),
    .B(_1624_),
    .Y(_1625_));
 sg13g2_or3_2 _5452_ (.A(net1486),
    .B(net1487),
    .C(_1393_),
    .X(_1626_));
 sg13g2_and2_1 _5453_ (.A(_1571_),
    .B(_1626_),
    .X(_1627_));
 sg13g2_or2_1 _5454_ (.X(_1628_),
    .B(_1600_),
    .A(_1573_));
 sg13g2_nor2_2 _5455_ (.A(_1561_),
    .B(_1574_),
    .Y(_1629_));
 sg13g2_inv_1 _5456_ (.Y(_1630_),
    .A(_1629_));
 sg13g2_nand2_2 _5457_ (.Y(_1631_),
    .A(_1626_),
    .B(_1629_));
 sg13g2_or3_2 _5458_ (.A(_1625_),
    .B(_1628_),
    .C(_1631_),
    .X(_1632_));
 sg13g2_xnor2_1 _5459_ (.Y(_1633_),
    .A(\usbfunction0.n1583_o[1] ),
    .B(_1632_));
 sg13g2_o21ai_1 _5460_ (.B1(_1633_),
    .Y(_1634_),
    .A1(_0695_),
    .A2(_1563_));
 sg13g2_nand2_1 _5461_ (.Y(_1635_),
    .A(_0030_),
    .B(_1632_));
 sg13g2_a21o_1 _5462_ (.A2(_1635_),
    .A1(_1634_),
    .B1(_1619_),
    .X(_1636_));
 sg13g2_o21ai_1 _5463_ (.B1(_1617_),
    .Y(_1637_),
    .A1(_0696_),
    .A2(_1614_));
 sg13g2_nand3_1 _5464_ (.B(_1618_),
    .C(_1637_),
    .A(_1607_),
    .Y(_1638_));
 sg13g2_a21oi_1 _5465_ (.A1(_0034_),
    .A2(_1583_),
    .Y(_1639_),
    .B1(_1591_));
 sg13g2_o21ai_1 _5466_ (.B1(_1638_),
    .Y(_1640_),
    .A1(_1592_),
    .A2(_1639_));
 sg13g2_nor3_1 _5467_ (.A(\usbfunction0.n1583_o[4] ),
    .B(_1576_),
    .C(_1602_),
    .Y(_1641_));
 sg13g2_a21oi_1 _5468_ (.A1(_0033_),
    .A2(_1601_),
    .Y(_1642_),
    .B1(_1641_));
 sg13g2_o21ai_1 _5469_ (.B1(_1636_),
    .Y(_1643_),
    .A1(_1593_),
    .A2(_1642_));
 sg13g2_nor2_1 _5470_ (.A(\usbfunction0.n1583_o[0] ),
    .B(_1562_),
    .Y(_1644_));
 sg13g2_nor3_1 _5471_ (.A(_1619_),
    .B(_1634_),
    .C(_1644_),
    .Y(_1645_));
 sg13g2_nor2_1 _5472_ (.A(net1594),
    .B(net1479),
    .Y(_1646_));
 sg13g2_nor4_1 _5473_ (.A(\usbfunction0.n2481_o[53] ),
    .B(\usbfunction0.n2481_o[52] ),
    .C(\usbfunction0.n2481_o[55] ),
    .D(\usbfunction0.n2481_o[54] ),
    .Y(_1647_));
 sg13g2_nor4_1 _5474_ (.A(net1477),
    .B(net1478),
    .C(net1480),
    .D(\usbfunction0.n2481_o[51] ),
    .Y(_1648_));
 sg13g2_nand2_1 _5475_ (.Y(_1649_),
    .A(_1647_),
    .B(_1648_));
 sg13g2_nor3_1 _5476_ (.A(net1415),
    .B(_1645_),
    .C(_1649_),
    .Y(_1650_));
 sg13g2_o21ai_1 _5477_ (.B1(_1650_),
    .Y(_1651_),
    .A1(_1640_),
    .A2(_1643_));
 sg13g2_mux2_1 _5478_ (.A0(net1798),
    .A1(_1563_),
    .S(_1651_),
    .X(\usbfunction0.n2353_o[0] ));
 sg13g2_nand4_1 _5479_ (.B(_1508_),
    .C(_1509_),
    .A(\usbfunction0.n2474_o[2] ),
    .Y(_1652_),
    .D(_1512_));
 sg13g2_mux2_1 _5480_ (.A0(\usbfunction0.n2353_o[0] ),
    .A1(_1546_),
    .S(net1178),
    .X(\usbfunction0.n2480_o[0] ));
 sg13g2_mux2_1 _5481_ (.A0(net1667),
    .A1(_1632_),
    .S(_1651_),
    .X(\usbfunction0.n2353_o[1] ));
 sg13g2_mux2_1 _5482_ (.A0(\usbfunction0.n2353_o[1] ),
    .A1(_1622_),
    .S(net1178),
    .X(\usbfunction0.n2480_o[1] ));
 sg13g2_mux2_1 _5483_ (.A0(net1656),
    .A1(_1615_),
    .S(_1651_),
    .X(\usbfunction0.n2353_o[2] ));
 sg13g2_mux2_1 _5484_ (.A0(\usbfunction0.n2353_o[2] ),
    .A1(_1608_),
    .S(net1178),
    .X(\usbfunction0.n2480_o[2] ));
 sg13g2_o21ai_1 _5485_ (.B1(_1606_),
    .Y(\usbfunction0.n2353_o[3] ),
    .A1(_0697_),
    .A2(_1651_));
 sg13g2_mux2_1 _5486_ (.A0(\usbfunction0.n2353_o[3] ),
    .A1(net1823),
    .S(net1179),
    .X(\usbfunction0.n2480_o[3] ));
 sg13g2_mux2_1 _5487_ (.A0(net1768),
    .A1(_1575_),
    .S(_1651_),
    .X(\usbfunction0.n2353_o[4] ));
 sg13g2_mux2_1 _5488_ (.A0(\usbfunction0.n2353_o[4] ),
    .A1(_1568_),
    .S(net1179),
    .X(\usbfunction0.n2480_o[4] ));
 sg13g2_mux2_1 _5489_ (.A0(net1753),
    .A1(_1601_),
    .S(_1651_),
    .X(\usbfunction0.n2353_o[5] ));
 sg13g2_mux2_1 _5490_ (.A0(\usbfunction0.n2353_o[5] ),
    .A1(_1595_),
    .S(net1179),
    .X(\usbfunction0.n2480_o[5] ));
 sg13g2_mux2_1 _5491_ (.A0(net1776),
    .A1(_1583_),
    .S(_1651_),
    .X(\usbfunction0.n2353_o[6] ));
 sg13g2_mux2_1 _5492_ (.A0(\usbfunction0.n2353_o[6] ),
    .A1(_1580_),
    .S(net1179),
    .X(\usbfunction0.n2480_o[6] ));
 sg13g2_o21ai_1 _5493_ (.B1(_1590_),
    .Y(\usbfunction0.n2353_o[7] ),
    .A1(_0703_),
    .A2(_1651_));
 sg13g2_mux2_1 _5494_ (.A0(\usbfunction0.n2353_o[7] ),
    .A1(_1586_),
    .S(net1179),
    .X(\usbfunction0.n2480_o[7] ));
 sg13g2_xnor2_1 _5495_ (.Y(_1653_),
    .A(\usbfunction0.n2649_q[0] ),
    .B(_1544_));
 sg13g2_xnor2_1 _5496_ (.Y(_1654_),
    .A(\usbfunction0.n2649_q[0] ),
    .B(_1545_));
 sg13g2_nand2_1 _5497_ (.Y(_1655_),
    .A(net1423),
    .B(_1653_));
 sg13g2_a21oi_1 _5498_ (.A1(_0763_),
    .A2(net1419),
    .Y(_1656_),
    .B1(_1631_));
 sg13g2_nor3_2 _5499_ (.A(_1557_),
    .B(_1573_),
    .C(_1600_),
    .Y(_1657_));
 sg13g2_nand2_1 _5500_ (.Y(_1658_),
    .A(_1612_),
    .B(_1657_));
 sg13g2_a21oi_1 _5501_ (.A1(_1655_),
    .A2(_1656_),
    .Y(_1659_),
    .B1(_1658_));
 sg13g2_nand2b_1 _5502_ (.Y(_1660_),
    .B(net1575),
    .A_N(net1491));
 sg13g2_a21oi_1 _5503_ (.A1(_1555_),
    .A2(net1576),
    .Y(\usbfunction0.n1101_o[0] ),
    .B1(_1659_));
 sg13g2_nor2_1 _5504_ (.A(net1179),
    .B(\usbfunction0.n1101_o[0] ),
    .Y(_1661_));
 sg13g2_a21oi_1 _5505_ (.A1(net1179),
    .A2(_1653_),
    .Y(\usbfunction0.n2477_o[0] ),
    .B1(_1661_));
 sg13g2_nand2_1 _5506_ (.Y(_1662_),
    .A(net1863),
    .B(_1545_));
 sg13g2_nand2_1 _5507_ (.Y(_1663_),
    .A(\usbfunction0.n2649_q[0] ),
    .B(\usbfunction0.n2649_q[1] ));
 sg13g2_xor2_1 _5508_ (.B(\usbfunction0.n2649_q[1] ),
    .A(\usbfunction0.n2649_q[0] ),
    .X(_1664_));
 sg13g2_mux2_2 _5509_ (.A0(_0764_),
    .A1(_1664_),
    .S(_1544_),
    .X(_1665_));
 sg13g2_o21ai_1 _5510_ (.B1(_1662_),
    .Y(_1666_),
    .A1(net1350),
    .A2(_1664_));
 sg13g2_nand2_1 _5511_ (.Y(_1667_),
    .A(net1424),
    .B(_1665_));
 sg13g2_nand2_1 _5512_ (.Y(_1668_),
    .A(\usbfunction0.n2651_q[1] ),
    .B(net1419));
 sg13g2_nand3_1 _5513_ (.B(_1667_),
    .C(_1668_),
    .A(_1626_),
    .Y(_1669_));
 sg13g2_a21oi_1 _5514_ (.A1(_1571_),
    .A2(_1669_),
    .Y(_1670_),
    .B1(_1560_));
 sg13g2_nor3_1 _5515_ (.A(_1573_),
    .B(_1613_),
    .C(_1670_),
    .Y(_1671_));
 sg13g2_nor3_1 _5516_ (.A(_1557_),
    .B(_1600_),
    .C(_1671_),
    .Y(_1672_));
 sg13g2_nand2b_1 _5517_ (.Y(_1673_),
    .B(net809),
    .A_N(net1489));
 sg13g2_a21oi_1 _5518_ (.A1(_1555_),
    .A2(_1673_),
    .Y(\usbfunction0.n1101_o[1] ),
    .B1(_1672_));
 sg13g2_nor2_1 _5519_ (.A(net1176),
    .B(\usbfunction0.n1101_o[1] ),
    .Y(_1674_));
 sg13g2_a21oi_1 _5520_ (.A1(net1176),
    .A2(_1666_),
    .Y(\usbfunction0.n2477_o[1] ),
    .B1(_1674_));
 sg13g2_nor2_1 _5521_ (.A(net1350),
    .B(_1663_),
    .Y(_1675_));
 sg13g2_nor3_2 _5522_ (.A(_0096_),
    .B(net1350),
    .C(_1663_),
    .Y(_1676_));
 sg13g2_xnor2_1 _5523_ (.Y(_1677_),
    .A(_0096_),
    .B(_1675_));
 sg13g2_xor2_1 _5524_ (.B(_1675_),
    .A(net1882),
    .X(_1678_));
 sg13g2_nor2_1 _5525_ (.A(net1419),
    .B(net1313),
    .Y(_1679_));
 sg13g2_a21oi_1 _5526_ (.A1(\usbfunction0.n2651_q[2] ),
    .A2(net1419),
    .Y(_1680_),
    .B1(_1679_));
 sg13g2_a21oi_1 _5527_ (.A1(_1626_),
    .A2(_1680_),
    .Y(_1681_),
    .B1(_1630_));
 sg13g2_o21ai_1 _5528_ (.B1(_1657_),
    .Y(_1682_),
    .A1(_1613_),
    .A2(_1681_));
 sg13g2_nand2b_1 _5529_ (.Y(_1683_),
    .B(net958),
    .A_N(net1489));
 sg13g2_o21ai_1 _5530_ (.B1(_1682_),
    .Y(\usbfunction0.n1101_o[2] ),
    .A1(_1556_),
    .A2(_1683_));
 sg13g2_nor2_1 _5531_ (.A(net1176),
    .B(\usbfunction0.n1101_o[2] ),
    .Y(_1684_));
 sg13g2_a21oi_1 _5532_ (.A1(net1176),
    .A2(net1313),
    .Y(\usbfunction0.n2477_o[2] ),
    .B1(_1684_));
 sg13g2_xnor2_1 _5533_ (.Y(_1685_),
    .A(_0097_),
    .B(_1676_));
 sg13g2_xor2_1 _5534_ (.B(_1676_),
    .A(_0097_),
    .X(_1686_));
 sg13g2_o21ai_1 _5535_ (.B1(_1626_),
    .Y(_1687_),
    .A1(_0765_),
    .A2(net1424));
 sg13g2_a21oi_1 _5536_ (.A1(net1424),
    .A2(_1685_),
    .Y(_1688_),
    .B1(_1687_));
 sg13g2_or3_1 _5537_ (.A(_1560_),
    .B(_1574_),
    .C(_1688_),
    .X(_1689_));
 sg13g2_nand2b_1 _5538_ (.Y(_1690_),
    .B(net934),
    .A_N(net1489));
 sg13g2_a22oi_1 _5539_ (.Y(\usbfunction0.n1101_o[3] ),
    .B1(_1690_),
    .B2(_1555_),
    .A2(_1689_),
    .A1(_1657_));
 sg13g2_nor2_1 _5540_ (.A(net1176),
    .B(\usbfunction0.n1101_o[3] ),
    .Y(_1691_));
 sg13g2_a21oi_1 _5541_ (.A1(net1176),
    .A2(net1307),
    .Y(\usbfunction0.n2477_o[3] ),
    .B1(_1691_));
 sg13g2_and3_2 _5542_ (.X(_1692_),
    .A(\usbfunction0.n2649_q[2] ),
    .B(\usbfunction0.n2649_q[3] ),
    .C(_1675_));
 sg13g2_nor2b_1 _5543_ (.A(_0098_),
    .B_N(_1692_),
    .Y(_1693_));
 sg13g2_xnor2_1 _5544_ (.Y(_1694_),
    .A(_0098_),
    .B(_1692_));
 sg13g2_xor2_1 _5545_ (.B(_1692_),
    .A(net1900),
    .X(_1695_));
 sg13g2_nor2_1 _5546_ (.A(net1418),
    .B(_1694_),
    .Y(_1696_));
 sg13g2_o21ai_1 _5547_ (.B1(_1626_),
    .Y(_1697_),
    .A1(net1899),
    .A2(net1424));
 sg13g2_o21ai_1 _5548_ (.B1(_1571_),
    .Y(_1698_),
    .A1(_1696_),
    .A2(_1697_));
 sg13g2_nor2_1 _5549_ (.A(_1560_),
    .B(_1573_),
    .Y(_1699_));
 sg13g2_a21oi_1 _5550_ (.A1(_1698_),
    .A2(_1699_),
    .Y(_1700_),
    .B1(_1600_));
 sg13g2_nor2_1 _5551_ (.A(_1555_),
    .B(_1700_),
    .Y(\usbfunction0.n1101_o[4] ));
 sg13g2_nor2_1 _5552_ (.A(net1177),
    .B(\usbfunction0.n1101_o[4] ),
    .Y(_1701_));
 sg13g2_a21oi_1 _5553_ (.A1(net1177),
    .A2(net1277),
    .Y(\usbfunction0.n2477_o[4] ),
    .B1(_1701_));
 sg13g2_xor2_1 _5554_ (.B(_1693_),
    .A(_0099_),
    .X(_1702_));
 sg13g2_xnor2_1 _5555_ (.Y(_1703_),
    .A(_0099_),
    .B(_1693_));
 sg13g2_o21ai_1 _5556_ (.B1(_1627_),
    .Y(_1704_),
    .A1(net1894),
    .A2(net1424));
 sg13g2_a21oi_1 _5557_ (.A1(net1424),
    .A2(net1268),
    .Y(_1705_),
    .B1(_1704_));
 sg13g2_nor3_1 _5558_ (.A(_1560_),
    .B(_1628_),
    .C(_1705_),
    .Y(_1706_));
 sg13g2_nor2_1 _5559_ (.A(_1555_),
    .B(_1706_),
    .Y(\usbfunction0.n1101_o[5] ));
 sg13g2_nor2_1 _5560_ (.A(net1177),
    .B(\usbfunction0.n1101_o[5] ),
    .Y(_1707_));
 sg13g2_a21oi_1 _5561_ (.A1(net1177),
    .A2(net1268),
    .Y(\usbfunction0.n2477_o[5] ),
    .B1(_1707_));
 sg13g2_nand3_1 _5562_ (.B(\usbfunction0.n2649_q[5] ),
    .C(_1692_),
    .A(\usbfunction0.n2649_q[4] ),
    .Y(_1708_));
 sg13g2_nor2_1 _5563_ (.A(_0100_),
    .B(_1708_),
    .Y(_1709_));
 sg13g2_xor2_1 _5564_ (.B(_1708_),
    .A(_0100_),
    .X(_1710_));
 sg13g2_xnor2_1 _5565_ (.Y(_1711_),
    .A(_0100_),
    .B(_1708_));
 sg13g2_nor2_1 _5566_ (.A(net1419),
    .B(_1710_),
    .Y(_1712_));
 sg13g2_nor2_1 _5567_ (.A(net1873),
    .B(net1423),
    .Y(_1713_));
 sg13g2_nor3_1 _5568_ (.A(_1631_),
    .B(_1712_),
    .C(_1713_),
    .Y(_1714_));
 sg13g2_nand2b_1 _5569_ (.Y(_1715_),
    .B(_1612_),
    .A_N(_1628_));
 sg13g2_nor2_1 _5570_ (.A(_1714_),
    .B(_1715_),
    .Y(_1716_));
 sg13g2_nor2_1 _5571_ (.A(_1555_),
    .B(_1716_),
    .Y(\usbfunction0.n1101_o[6] ));
 sg13g2_nor2_1 _5572_ (.A(net1177),
    .B(\usbfunction0.n1101_o[6] ),
    .Y(_1717_));
 sg13g2_a21oi_1 _5573_ (.A1(net1176),
    .A2(net1267),
    .Y(\usbfunction0.n2477_o[6] ),
    .B1(_1717_));
 sg13g2_xnor2_1 _5574_ (.Y(_1718_),
    .A(net1896),
    .B(_1709_));
 sg13g2_xor2_1 _5575_ (.B(_1709_),
    .A(net1850),
    .X(_1719_));
 sg13g2_nor2_1 _5576_ (.A(net1419),
    .B(net1264),
    .Y(_1720_));
 sg13g2_nor2_1 _5577_ (.A(net919),
    .B(net1423),
    .Y(_1721_));
 sg13g2_nor4_1 _5578_ (.A(_1631_),
    .B(_1658_),
    .C(_1720_),
    .D(_1721_),
    .Y(\usbfunction0.n1101_o[7] ));
 sg13g2_nor2_1 _5579_ (.A(net1177),
    .B(\usbfunction0.n1101_o[7] ),
    .Y(_1722_));
 sg13g2_a21oi_1 _5580_ (.A1(net1176),
    .A2(_1719_),
    .Y(\usbfunction0.n2477_o[7] ),
    .B1(_1722_));
 sg13g2_a21o_1 _5581_ (.A2(net1384),
    .A1(net1602),
    .B1(_1452_),
    .X(\usbfunction0.n1630_o[0] ));
 sg13g2_and2_1 _5582_ (.A(_0035_),
    .B(_1357_),
    .X(_1723_));
 sg13g2_and2_1 _5583_ (.A(net548),
    .B(_1723_),
    .X(_1724_));
 sg13g2_nand2_1 _5584_ (.Y(_1725_),
    .A(\usbfunction0.n1630_o[0] ),
    .B(net1404));
 sg13g2_xnor2_1 _5585_ (.Y(\usbfunction0.n2433_o[0] ),
    .A(_1454_),
    .B(_1725_));
 sg13g2_nor4_2 _5586_ (.A(_0703_),
    .B(net1477),
    .C(net1479),
    .Y(_1726_),
    .D(net1481));
 sg13g2_mux2_1 _5587_ (.A0(_1726_),
    .A1(net897),
    .S(net1385),
    .X(\usbfunction0.n1630_o[1] ));
 sg13g2_nand2_1 _5588_ (.Y(_1727_),
    .A(net897),
    .B(net1403));
 sg13g2_xor2_1 _5589_ (.B(_1727_),
    .A(_1458_),
    .X(\usbfunction0.n2433_o[1] ));
 sg13g2_nand2_1 _5590_ (.Y(_1728_),
    .A(net1028),
    .B(net1397));
 sg13g2_nor2b_2 _5591_ (.A(\usbfunction0.n1360_o[0] ),
    .B_N(net1481),
    .Y(_1729_));
 sg13g2_nand2_1 _5592_ (.Y(_1730_),
    .A(_1646_),
    .B(_1729_));
 sg13g2_o21ai_1 _5593_ (.B1(_1728_),
    .Y(\usbfunction0.n1630_o[2] ),
    .A1(net1385),
    .A2(_1730_));
 sg13g2_nand2_1 _5594_ (.Y(_1731_),
    .A(net1028),
    .B(net1403));
 sg13g2_xor2_1 _5595_ (.B(_1731_),
    .A(_1462_),
    .X(\usbfunction0.n2433_o[2] ));
 sg13g2_nand2_1 _5596_ (.Y(_1732_),
    .A(net1127),
    .B(net1397));
 sg13g2_nand3_1 _5597_ (.B(net1480),
    .C(_1646_),
    .A(net1625),
    .Y(_1733_));
 sg13g2_o21ai_1 _5598_ (.B1(_1732_),
    .Y(\usbfunction0.n1630_o[3] ),
    .A1(net1385),
    .A2(_1733_));
 sg13g2_nand2_1 _5599_ (.Y(_1734_),
    .A(net1127),
    .B(net1403));
 sg13g2_xor2_1 _5600_ (.B(_1734_),
    .A(_1466_),
    .X(\usbfunction0.n2433_o[3] ));
 sg13g2_nor4_1 _5601_ (.A(\usbfunction0.n1360_o[0] ),
    .B(net1477),
    .C(_0706_),
    .D(net1480),
    .Y(_1735_));
 sg13g2_mux2_1 _5602_ (.A0(_1735_),
    .A1(net926),
    .S(net1382),
    .X(\usbfunction0.n1630_o[4] ));
 sg13g2_nand2_1 _5603_ (.Y(_1736_),
    .A(net926),
    .B(net1402));
 sg13g2_xor2_1 _5604_ (.B(_1736_),
    .A(_1414_),
    .X(\usbfunction0.n2433_o[4] ));
 sg13g2_nand2_1 _5605_ (.Y(_1737_),
    .A(net900),
    .B(net1396));
 sg13g2_nor2_1 _5606_ (.A(_0703_),
    .B(net1480),
    .Y(_1738_));
 sg13g2_nand3_1 _5607_ (.B(net1478),
    .C(_1738_),
    .A(_0705_),
    .Y(_1739_));
 sg13g2_o21ai_1 _5608_ (.B1(_1737_),
    .Y(\usbfunction0.n1630_o[5] ),
    .A1(net1382),
    .A2(_1739_));
 sg13g2_nand2_1 _5609_ (.Y(_1740_),
    .A(net900),
    .B(net1402));
 sg13g2_xor2_1 _5610_ (.B(_1740_),
    .A(_1418_),
    .X(\usbfunction0.n2433_o[5] ));
 sg13g2_nand2_1 _5611_ (.Y(_1741_),
    .A(net776),
    .B(net1396));
 sg13g2_nand3_1 _5612_ (.B(net1479),
    .C(_1729_),
    .A(_0705_),
    .Y(_1742_));
 sg13g2_o21ai_1 _5613_ (.B1(_1741_),
    .Y(\usbfunction0.n1630_o[6] ),
    .A1(net1383),
    .A2(_1742_));
 sg13g2_nand2_1 _5614_ (.Y(_1743_),
    .A(net776),
    .B(net1402));
 sg13g2_xor2_1 _5615_ (.B(_1743_),
    .A(_1423_),
    .X(\usbfunction0.n2433_o[6] ));
 sg13g2_nand2_1 _5616_ (.Y(_1744_),
    .A(net761),
    .B(net1397));
 sg13g2_nand4_1 _5617_ (.B(_0705_),
    .C(net1478),
    .A(net1625),
    .Y(_1745_),
    .D(net1481));
 sg13g2_o21ai_1 _5618_ (.B1(_1744_),
    .Y(\usbfunction0.n1630_o[7] ),
    .A1(net1385),
    .A2(net1626));
 sg13g2_nand2_1 _5619_ (.Y(_1746_),
    .A(net761),
    .B(net1403));
 sg13g2_xor2_1 _5620_ (.B(_1746_),
    .A(_1408_),
    .X(\usbfunction0.n2433_o[7] ));
 sg13g2_or3_1 _5621_ (.A(\usbfunction0.n1360_o[0] ),
    .B(_0705_),
    .C(net1480),
    .X(_1747_));
 sg13g2_nor3_1 _5622_ (.A(net1479),
    .B(net1385),
    .C(_1747_),
    .Y(_1748_));
 sg13g2_a21o_1 _5623_ (.A2(net1385),
    .A1(net774),
    .B1(_1748_),
    .X(\usbfunction0.n1630_o[8] ));
 sg13g2_nand2_1 _5624_ (.Y(_1749_),
    .A(net774),
    .B(net1403));
 sg13g2_xor2_1 _5625_ (.B(_1749_),
    .A(_1484_),
    .X(\usbfunction0.n2433_o[8] ));
 sg13g2_nand2_1 _5626_ (.Y(_1750_),
    .A(net1477),
    .B(_1738_));
 sg13g2_nor3_1 _5627_ (.A(net1478),
    .B(net1383),
    .C(_1750_),
    .Y(_1751_));
 sg13g2_a21o_1 _5628_ (.A2(net1383),
    .A1(net631),
    .B1(_1751_),
    .X(\usbfunction0.n1630_o[9] ));
 sg13g2_nand2_1 _5629_ (.Y(_1752_),
    .A(net631),
    .B(net1402));
 sg13g2_xor2_1 _5630_ (.B(_1752_),
    .A(_1476_),
    .X(\usbfunction0.n2433_o[9] ));
 sg13g2_nand2_1 _5631_ (.Y(_1753_),
    .A(net1477),
    .B(_1729_));
 sg13g2_nor3_1 _5632_ (.A(net1478),
    .B(net1382),
    .C(_1753_),
    .Y(_1754_));
 sg13g2_a21o_1 _5633_ (.A2(net1382),
    .A1(net771),
    .B1(_1754_),
    .X(\usbfunction0.n1630_o[10] ));
 sg13g2_nand2_1 _5634_ (.Y(_1755_),
    .A(net771),
    .B(net1402));
 sg13g2_xor2_1 _5635_ (.B(_1755_),
    .A(_1480_),
    .X(\usbfunction0.n2433_o[10] ));
 sg13g2_nand3_1 _5636_ (.B(net1477),
    .C(net1480),
    .A(\usbfunction0.n1360_o[0] ),
    .Y(_1756_));
 sg13g2_nor3_1 _5637_ (.A(net1478),
    .B(net1383),
    .C(_1756_),
    .Y(_1757_));
 sg13g2_a21o_1 _5638_ (.A2(net1382),
    .A1(net909),
    .B1(_1757_),
    .X(\usbfunction0.n1630_o[11] ));
 sg13g2_nand2_1 _5639_ (.Y(_1758_),
    .A(net909),
    .B(net1402));
 sg13g2_xor2_1 _5640_ (.B(_1758_),
    .A(_1472_),
    .X(\usbfunction0.n2433_o[11] ));
 sg13g2_nor3_1 _5641_ (.A(_0706_),
    .B(net1397),
    .C(_1747_),
    .Y(_1759_));
 sg13g2_a21o_1 _5642_ (.A2(net1385),
    .A1(net939),
    .B1(_1759_),
    .X(\usbfunction0.n1630_o[12] ));
 sg13g2_nand2_1 _5643_ (.Y(_1760_),
    .A(net939),
    .B(net1403));
 sg13g2_xor2_1 _5644_ (.B(_1760_),
    .A(_1436_),
    .X(\usbfunction0.n2433_o[12] ));
 sg13g2_nor3_1 _5645_ (.A(_0706_),
    .B(net1396),
    .C(_1750_),
    .Y(_1761_));
 sg13g2_a21o_1 _5646_ (.A2(net1382),
    .A1(net692),
    .B1(_1761_),
    .X(\usbfunction0.n1630_o[13] ));
 sg13g2_nand2_1 _5647_ (.Y(_1762_),
    .A(net692),
    .B(net1402));
 sg13g2_xnor2_1 _5648_ (.Y(\usbfunction0.n2433_o[13] ),
    .A(_1432_),
    .B(_1762_));
 sg13g2_nor3_1 _5649_ (.A(_0706_),
    .B(net1396),
    .C(_1753_),
    .Y(_1763_));
 sg13g2_a21o_1 _5650_ (.A2(net1382),
    .A1(net817),
    .B1(_1763_),
    .X(\usbfunction0.n1630_o[14] ));
 sg13g2_nand2_1 _5651_ (.Y(_1764_),
    .A(net817),
    .B(net1402));
 sg13g2_xor2_1 _5652_ (.B(_1764_),
    .A(_1428_),
    .X(\usbfunction0.n2433_o[14] ));
 sg13g2_nor3_1 _5653_ (.A(_0706_),
    .B(net1396),
    .C(_1756_),
    .Y(_1765_));
 sg13g2_a21o_1 _5654_ (.A2(net1382),
    .A1(net624),
    .B1(_1765_),
    .X(\usbfunction0.n1630_o[15] ));
 sg13g2_nand2_1 _5655_ (.Y(_1766_),
    .A(net624),
    .B(net1403));
 sg13g2_xnor2_1 _5656_ (.Y(\usbfunction0.n2433_o[15] ),
    .A(_1446_),
    .B(_1766_));
 sg13g2_nand2_1 _5657_ (.Y(_1767_),
    .A(net1421),
    .B(\usbfunction0.n1630_o[1] ));
 sg13g2_and2_1 _5658_ (.A(net843),
    .B(_1767_),
    .X(_1768_));
 sg13g2_nor2_1 _5659_ (.A(net843),
    .B(_1767_),
    .Y(_1769_));
 sg13g2_or3_2 _5660_ (.A(\usbfunction0.n2098_o ),
    .B(_1403_),
    .C(_1407_),
    .X(_1770_));
 sg13g2_nor2_1 _5661_ (.A(_1457_),
    .B(_1770_),
    .Y(_1771_));
 sg13g2_nor4_1 _5662_ (.A(net1390),
    .B(_1768_),
    .C(_1769_),
    .D(_1771_),
    .Y(\usbfunction0.n2257_o[1] ));
 sg13g2_nand2_1 _5663_ (.Y(_1772_),
    .A(net1425),
    .B(\usbfunction0.n1630_o[2] ));
 sg13g2_and2_1 _5664_ (.A(net841),
    .B(_1772_),
    .X(_1773_));
 sg13g2_nor2_1 _5665_ (.A(net841),
    .B(_1772_),
    .Y(_1774_));
 sg13g2_nor2_1 _5666_ (.A(_1461_),
    .B(net1388),
    .Y(_1775_));
 sg13g2_nor4_1 _5667_ (.A(net1390),
    .B(_1773_),
    .C(_1774_),
    .D(_1775_),
    .Y(\usbfunction0.n2257_o[2] ));
 sg13g2_nand2_1 _5668_ (.Y(_1776_),
    .A(net1425),
    .B(\usbfunction0.n1630_o[3] ));
 sg13g2_xnor2_1 _5669_ (.Y(_1777_),
    .A(net840),
    .B(_1776_));
 sg13g2_nor2_1 _5670_ (.A(_1465_),
    .B(net1388),
    .Y(_1778_));
 sg13g2_nor3_1 _5671_ (.A(net1390),
    .B(_1777_),
    .C(_1778_),
    .Y(\usbfunction0.n2257_o[3] ));
 sg13g2_nand2_1 _5672_ (.Y(_1779_),
    .A(net1421),
    .B(\usbfunction0.n1630_o[4] ));
 sg13g2_and2_1 _5673_ (.A(net700),
    .B(_1779_),
    .X(_1780_));
 sg13g2_nor2_1 _5674_ (.A(net700),
    .B(_1779_),
    .Y(_1781_));
 sg13g2_nor2_1 _5675_ (.A(_1413_),
    .B(net1387),
    .Y(_1782_));
 sg13g2_nor4_1 _5676_ (.A(net1389),
    .B(_1780_),
    .C(_1781_),
    .D(_1782_),
    .Y(\usbfunction0.n2257_o[4] ));
 sg13g2_nand2_1 _5677_ (.Y(_1783_),
    .A(net1421),
    .B(\usbfunction0.n1630_o[5] ));
 sg13g2_and2_1 _5678_ (.A(net879),
    .B(_1783_),
    .X(_1784_));
 sg13g2_nor2_1 _5679_ (.A(net879),
    .B(_1783_),
    .Y(_1785_));
 sg13g2_nor2_1 _5680_ (.A(_1417_),
    .B(net1387),
    .Y(_1786_));
 sg13g2_nor4_1 _5681_ (.A(net1389),
    .B(_1784_),
    .C(_1785_),
    .D(_1786_),
    .Y(\usbfunction0.n2257_o[5] ));
 sg13g2_nand2_1 _5682_ (.Y(_1787_),
    .A(net1422),
    .B(\usbfunction0.n1630_o[6] ));
 sg13g2_and2_1 _5683_ (.A(net678),
    .B(_1787_),
    .X(_1788_));
 sg13g2_nor2_1 _5684_ (.A(net678),
    .B(_1787_),
    .Y(_1789_));
 sg13g2_nor2_1 _5685_ (.A(_1422_),
    .B(net1387),
    .Y(_1790_));
 sg13g2_nor4_1 _5686_ (.A(net1390),
    .B(_1788_),
    .C(_1789_),
    .D(_1790_),
    .Y(\usbfunction0.n2257_o[6] ));
 sg13g2_nand2_1 _5687_ (.Y(_1791_),
    .A(net1425),
    .B(\usbfunction0.n1630_o[7] ));
 sg13g2_and2_1 _5688_ (.A(net727),
    .B(_1791_),
    .X(_1792_));
 sg13g2_nor2_1 _5689_ (.A(net727),
    .B(_1791_),
    .Y(_1793_));
 sg13g2_nor2_1 _5690_ (.A(_1402_),
    .B(net1388),
    .Y(_1794_));
 sg13g2_nor4_1 _5691_ (.A(net1390),
    .B(_1792_),
    .C(_1793_),
    .D(_1794_),
    .Y(\usbfunction0.n2257_o[7] ));
 sg13g2_nand2_1 _5692_ (.Y(_1795_),
    .A(net1425),
    .B(\usbfunction0.n1630_o[8] ));
 sg13g2_and2_1 _5693_ (.A(net714),
    .B(_1795_),
    .X(_1796_));
 sg13g2_nor2_1 _5694_ (.A(net714),
    .B(_1795_),
    .Y(_1797_));
 sg13g2_nor2_1 _5695_ (.A(_1483_),
    .B(net1388),
    .Y(_1798_));
 sg13g2_nor4_1 _5696_ (.A(net1390),
    .B(_1796_),
    .C(_1797_),
    .D(_1798_),
    .Y(\usbfunction0.n2257_o[8] ));
 sg13g2_nand2_1 _5697_ (.Y(_1799_),
    .A(net1422),
    .B(\usbfunction0.n1630_o[9] ));
 sg13g2_and2_1 _5698_ (.A(net751),
    .B(_1799_),
    .X(_1800_));
 sg13g2_nor2_1 _5699_ (.A(net751),
    .B(_1799_),
    .Y(_1801_));
 sg13g2_nor2_1 _5700_ (.A(_1475_),
    .B(net1388),
    .Y(_1802_));
 sg13g2_nor4_1 _5701_ (.A(net1390),
    .B(_1800_),
    .C(_1801_),
    .D(_1802_),
    .Y(\usbfunction0.n2257_o[9] ));
 sg13g2_nand2_1 _5702_ (.Y(_1803_),
    .A(net1421),
    .B(\usbfunction0.n1630_o[10] ));
 sg13g2_and2_1 _5703_ (.A(net661),
    .B(_1803_),
    .X(_1804_));
 sg13g2_nor2_1 _5704_ (.A(net661),
    .B(_1803_),
    .Y(_1805_));
 sg13g2_nor2_1 _5705_ (.A(_1479_),
    .B(net1387),
    .Y(_1806_));
 sg13g2_nor4_1 _5706_ (.A(net1389),
    .B(_1804_),
    .C(_1805_),
    .D(_1806_),
    .Y(\usbfunction0.n2257_o[10] ));
 sg13g2_nand2_1 _5707_ (.Y(_1807_),
    .A(net1421),
    .B(\usbfunction0.n1630_o[11] ));
 sg13g2_and2_1 _5708_ (.A(net827),
    .B(_1807_),
    .X(_1808_));
 sg13g2_nor2_1 _5709_ (.A(net827),
    .B(_1807_),
    .Y(_1809_));
 sg13g2_nor2_1 _5710_ (.A(_1471_),
    .B(net1387),
    .Y(_1810_));
 sg13g2_nor4_2 _5711_ (.A(net1389),
    .B(_1808_),
    .C(_1809_),
    .Y(\usbfunction0.n2257_o[11] ),
    .D(_1810_));
 sg13g2_nand2_1 _5712_ (.Y(_1811_),
    .A(net1425),
    .B(\usbfunction0.n1630_o[12] ));
 sg13g2_xnor2_1 _5713_ (.Y(_1812_),
    .A(net866),
    .B(_1811_));
 sg13g2_nor2_1 _5714_ (.A(_1435_),
    .B(net1388),
    .Y(_1813_));
 sg13g2_nor3_1 _5715_ (.A(net1389),
    .B(_1812_),
    .C(_1813_),
    .Y(\usbfunction0.n2257_o[12] ));
 sg13g2_nand2_1 _5716_ (.Y(_1814_),
    .A(net1421),
    .B(\usbfunction0.n1630_o[13] ));
 sg13g2_and2_1 _5717_ (.A(net821),
    .B(_1814_),
    .X(_1815_));
 sg13g2_nor2_1 _5718_ (.A(net821),
    .B(_1814_),
    .Y(_1816_));
 sg13g2_nor2_1 _5719_ (.A(_1430_),
    .B(net1387),
    .Y(_1817_));
 sg13g2_nor4_1 _5720_ (.A(net1389),
    .B(_1815_),
    .C(_1816_),
    .D(_1817_),
    .Y(\usbfunction0.n2257_o[13] ));
 sg13g2_nand2_1 _5721_ (.Y(_1818_),
    .A(net1421),
    .B(\usbfunction0.n1630_o[14] ));
 sg13g2_and2_1 _5722_ (.A(net911),
    .B(_1818_),
    .X(_1819_));
 sg13g2_nor2_1 _5723_ (.A(net911),
    .B(_1818_),
    .Y(_1820_));
 sg13g2_nor2_1 _5724_ (.A(_1427_),
    .B(net1387),
    .Y(_1821_));
 sg13g2_nor4_2 _5725_ (.A(net1389),
    .B(_1819_),
    .C(_1820_),
    .Y(\usbfunction0.n2257_o[14] ),
    .D(_1821_));
 sg13g2_nand2_1 _5726_ (.Y(_1822_),
    .A(net1421),
    .B(\usbfunction0.n1630_o[15] ));
 sg13g2_xnor2_1 _5727_ (.Y(_1823_),
    .A(net705),
    .B(_1822_));
 sg13g2_nor2_1 _5728_ (.A(_1442_),
    .B(net1388),
    .Y(_1824_));
 sg13g2_nor3_1 _5729_ (.A(net1389),
    .B(_1823_),
    .C(_1824_),
    .Y(\usbfunction0.n2257_o[15] ));
 sg13g2_nand2_1 _5730_ (.Y(_1825_),
    .A(net1422),
    .B(\usbfunction0.n1630_o[0] ));
 sg13g2_xor2_1 _5731_ (.B(_1825_),
    .A(net1839),
    .X(_1826_));
 sg13g2_nor2_1 _5732_ (.A(_1441_),
    .B(net1387),
    .Y(_1827_));
 sg13g2_a21oi_1 _5733_ (.A1(_1453_),
    .A2(_1826_),
    .Y(\usbfunction0.n2254_o ),
    .B1(_1827_));
 sg13g2_xor2_1 _5734_ (.B(\n352_o[7] ),
    .A(net611),
    .X(\scl_uarttx0.scl_baudrategenerator0.n6878_o[0] ));
 sg13g2_nand2b_1 _5735_ (.Y(_1828_),
    .B(\s_m_packetdata_2_rewired[5] ),
    .A_N(\s_m_packetdata_2_rewired[6] ));
 sg13g2_or2_1 _5736_ (.X(_1829_),
    .B(_1828_),
    .A(_1371_));
 sg13g2_nor4_1 _5737_ (.A(\usbfunction0.n2481_o[37] ),
    .B(\usbfunction0.n2481_o[36] ),
    .C(\usbfunction0.n2481_o[39] ),
    .D(\usbfunction0.n2481_o[38] ),
    .Y(_1830_));
 sg13g2_nor4_1 _5738_ (.A(\usbfunction0.n2481_o[28] ),
    .B(\usbfunction0.n2481_o[30] ),
    .C(\usbfunction0.n2481_o[32] ),
    .D(\usbfunction0.n2481_o[33] ),
    .Y(_1831_));
 sg13g2_nand3_1 _5739_ (.B(_1376_),
    .C(_1392_),
    .A(\s_m_packetdata_2_rewired[13] ),
    .Y(_1832_));
 sg13g2_nor4_1 _5740_ (.A(\usbfunction0.n2098_o ),
    .B(\usbfunction0.n2481_o[29] ),
    .C(\usbfunction0.n2481_o[35] ),
    .D(\usbfunction0.n2481_o[34] ),
    .Y(_1833_));
 sg13g2_nand4_1 _5741_ (.B(_1830_),
    .C(_1831_),
    .A(_1440_),
    .Y(_1834_),
    .D(_1833_));
 sg13g2_nor3_1 _5742_ (.A(\s_m_packetdata_2_rewired[7] ),
    .B(_0723_),
    .C(_1828_),
    .Y(_1835_));
 sg13g2_nand2_1 _5743_ (.Y(_1836_),
    .A(_1374_),
    .B(_1835_));
 sg13g2_nor4_1 _5744_ (.A(_1552_),
    .B(_1832_),
    .C(_1834_),
    .D(_1836_),
    .Y(_1837_));
 sg13g2_nand2b_2 _5745_ (.Y(_1838_),
    .B(_1837_),
    .A_N(_1829_));
 sg13g2_inv_1 _5746_ (.Y(_1839_),
    .A(_1838_));
 sg13g2_mux2_2 _5747_ (.A0(s_m_packetdata_2_bit_17),
    .A1(net1834),
    .S(_1838_),
    .X(n350_o));
 sg13g2_mux2_2 _5748_ (.A0(net1803),
    .A1(net1811),
    .S(_1838_),
    .X(n183_o));
 sg13g2_nand2b_1 _5749_ (.Y(\usbfunction0.n1189_o[0] ),
    .B(net1576),
    .A_N(net1391));
 sg13g2_nor2_1 _5750_ (.A(net1391),
    .B(_1673_),
    .Y(\usbfunction0.n1189_o[1] ));
 sg13g2_nor2_1 _5751_ (.A(net1391),
    .B(_1683_),
    .Y(\usbfunction0.n1189_o[2] ));
 sg13g2_nor2_1 _5752_ (.A(net1391),
    .B(_1690_),
    .Y(\usbfunction0.n1189_o[3] ));
 sg13g2_nor2_2 _5753_ (.A(_1384_),
    .B(_1551_),
    .Y(_1840_));
 sg13g2_mux2_1 _5754_ (.A0(_0957_),
    .A1(net1803),
    .S(_1840_),
    .X(\usbfunction0.n1083_o[0] ));
 sg13g2_mux2_1 _5755_ (.A0(net1790),
    .A1(s_m_packetdata_2_bit_17),
    .S(_1840_),
    .X(\usbfunction0.n1083_o[1] ));
 sg13g2_mux2_1 _5756_ (.A0(_0976_),
    .A1(net1767),
    .S(_1840_),
    .X(\usbfunction0.n1083_o[2] ));
 sg13g2_mux2_1 _5757_ (.A0(_0946_),
    .A1(\s_m_packetdata_2_rewired[19] ),
    .S(_1840_),
    .X(\usbfunction0.n1083_o[3] ));
 sg13g2_mux2_1 _5758_ (.A0(_0980_),
    .A1(net1759),
    .S(_1840_),
    .X(\usbfunction0.n1083_o[4] ));
 sg13g2_mux2_1 _5759_ (.A0(_0985_),
    .A1(net1595),
    .S(_1840_),
    .X(\usbfunction0.n1083_o[5] ));
 sg13g2_mux2_1 _5760_ (.A0(_0969_),
    .A1(net1617),
    .S(_1840_),
    .X(\usbfunction0.n1083_o[6] ));
 sg13g2_nor2_1 _5761_ (.A(\usbfunction0.n2627_q ),
    .B(\usbfunction0.n1974_o ),
    .Y(_1841_));
 sg13g2_nor4_2 _5762_ (.A(\usbfunction0.functionreset0.in_unnamed_2[1] ),
    .B(\usbfunction0.functionreset0.in_unnamed_2[0] ),
    .C(\usbfunction0.functionreset0.in_unnamed_2[3] ),
    .Y(_1842_),
    .D(\usbfunction0.functionreset0.in_unnamed_2[2] ));
 sg13g2_nor3_1 _5763_ (.A(\usbfunction0.n2634_q[2] ),
    .B(_1356_),
    .C(_1842_),
    .Y(_1843_));
 sg13g2_nor2b_1 _5764_ (.A(_0036_),
    .B_N(_1843_),
    .Y(_1844_));
 sg13g2_nand2_1 _5765_ (.Y(_1845_),
    .A(_1006_),
    .B(_1844_));
 sg13g2_or2_1 _5766_ (.X(_1846_),
    .B(_1845_),
    .A(_1841_));
 sg13g2_and2_1 _5767_ (.A(\usbfunction0.n2631_q ),
    .B(_1843_),
    .X(_1847_));
 sg13g2_and4_1 _5768_ (.A(_0041_),
    .B(_0040_),
    .C(_1006_),
    .D(_1847_),
    .X(_1848_));
 sg13g2_inv_1 _5769_ (.Y(_1849_),
    .A(net1364));
 sg13g2_nor2b_2 _5770_ (.A(\scl_fifo0.n2689_o[1] ),
    .B_N(\scl_fifo0.n2689_o[0] ),
    .Y(_1850_));
 sg13g2_nor2b_2 _5771_ (.A(\scl_fifo0.n2689_o[0] ),
    .B_N(\scl_fifo0.n2689_o[1] ),
    .Y(_1851_));
 sg13g2_o21ai_1 _5772_ (.B1(_1848_),
    .Y(_1852_),
    .A1(_1850_),
    .A2(_1851_));
 sg13g2_or2_1 _5773_ (.X(_1853_),
    .B(_1848_),
    .A(_0039_));
 sg13g2_nand3_1 _5774_ (.B(_1852_),
    .C(_1853_),
    .A(net1362),
    .Y(_1854_));
 sg13g2_o21ai_1 _5775_ (.B1(_1854_),
    .Y(_1855_),
    .A1(_0711_),
    .A2(net1362));
 sg13g2_nor3_1 _5776_ (.A(\usbfunction0.n2627_q ),
    .B(\usbfunction0.n1974_o ),
    .C(_1845_),
    .Y(_1856_));
 sg13g2_nand3_1 _5777_ (.B(_1841_),
    .C(_1844_),
    .A(_1006_),
    .Y(_1857_));
 sg13g2_nand2b_1 _5778_ (.Y(_1858_),
    .B(_1855_),
    .A_N(_1857_));
 sg13g2_xnor2_1 _5779_ (.Y(\scl_fifo0.n2722_o[1] ),
    .A(_1855_),
    .B(net1361));
 sg13g2_nand3_1 _5780_ (.B(\scl_fifo0.n2689_o[0] ),
    .C(net1364),
    .A(\scl_fifo0.n2689_o[1] ),
    .Y(_1859_));
 sg13g2_nor2_1 _5781_ (.A(_0122_),
    .B(_1859_),
    .Y(_1860_));
 sg13g2_o21ai_1 _5782_ (.B1(net1362),
    .Y(_1861_),
    .A1(_0122_),
    .A2(_1859_));
 sg13g2_a21o_1 _5783_ (.A2(_1859_),
    .A1(_0122_),
    .B1(_1861_),
    .X(_1862_));
 sg13g2_o21ai_1 _5784_ (.B1(_1862_),
    .Y(_1863_),
    .A1(_0121_),
    .A2(net1362));
 sg13g2_inv_1 _5785_ (.Y(_1864_),
    .A(_1863_));
 sg13g2_or2_1 _5786_ (.X(_1865_),
    .B(_1863_),
    .A(_1858_));
 sg13g2_xnor2_1 _5787_ (.Y(\scl_fifo0.n2722_o[2] ),
    .A(_1858_),
    .B(_1863_));
 sg13g2_nor2_1 _5788_ (.A(net1836),
    .B(_1846_),
    .Y(_1866_));
 sg13g2_xnor2_1 _5789_ (.Y(_1867_),
    .A(_0124_),
    .B(_1860_));
 sg13g2_a21oi_1 _5790_ (.A1(_1846_),
    .A2(_1867_),
    .Y(_1868_),
    .B1(_1866_));
 sg13g2_nand4_1 _5791_ (.B(net1361),
    .C(_1864_),
    .A(_1855_),
    .Y(_1869_),
    .D(_1868_));
 sg13g2_xnor2_1 _5792_ (.Y(_1870_),
    .A(_1865_),
    .B(_1868_));
 sg13g2_inv_1 _5793_ (.Y(\scl_fifo0.n2722_o[3] ),
    .A(_1870_));
 sg13g2_nor2_1 _5794_ (.A(net1858),
    .B(net1362),
    .Y(_1871_));
 sg13g2_nand2_1 _5795_ (.Y(_1872_),
    .A(\scl_fifo0.n2689_o[2] ),
    .B(\scl_fifo0.n2689_o[3] ));
 sg13g2_nor2_1 _5796_ (.A(_1859_),
    .B(_1872_),
    .Y(_1873_));
 sg13g2_xnor2_1 _5797_ (.Y(_1874_),
    .A(_0126_),
    .B(net1349));
 sg13g2_a21oi_1 _5798_ (.A1(net1362),
    .A2(_1874_),
    .Y(_1875_),
    .B1(_1871_));
 sg13g2_o21ai_1 _5799_ (.B1(net1361),
    .Y(_1876_),
    .A1(_1869_),
    .A2(_1875_));
 sg13g2_a21o_1 _5800_ (.A2(_1875_),
    .A1(_1869_),
    .B1(_1876_),
    .X(_1877_));
 sg13g2_o21ai_1 _5801_ (.B1(_1877_),
    .Y(\scl_fifo0.n2722_o[4] ),
    .A1(net1361),
    .A2(_1875_));
 sg13g2_xor2_1 _5802_ (.B(net1364),
    .A(\scl_fifo0.n2689_o[0] ),
    .X(_1878_));
 sg13g2_nor2_1 _5803_ (.A(net1641),
    .B(net1362),
    .Y(_1879_));
 sg13g2_a21oi_2 _5804_ (.B1(_1879_),
    .Y(_1880_),
    .A2(_1878_),
    .A1(net1362));
 sg13g2_inv_1 _5805_ (.Y(\scl_fifo0.n2694_o[0] ),
    .A(_1880_));
 sg13g2_xor2_1 _5806_ (.B(_1318_),
    .A(net1737),
    .X(\scl_uarttx0.scl_counter0.n6919_o[0] ));
 sg13g2_xor2_1 _5807_ (.B(_1319_),
    .A(net1848),
    .X(\scl_uarttx0.scl_counter0.n6919_o[1] ));
 sg13g2_xnor2_1 _5808_ (.Y(\scl_uarttx0.scl_counter0.n6919_o[3] ),
    .A(net992),
    .B(_1321_));
 sg13g2_nor2_1 _5809_ (.A(_1269_),
    .B(net1262),
    .Y(_1881_));
 sg13g2_xor2_1 _5810_ (.B(net1262),
    .A(_1269_),
    .X(\scl_uarttx0.scl_baudrategenerator0.n6892_o[1] ));
 sg13g2_xnor2_1 _5811_ (.Y(\scl_uarttx0.scl_baudrategenerator0.n6892_o[2] ),
    .A(_1270_),
    .B(_1881_));
 sg13g2_nor2_1 _5812_ (.A(_1271_),
    .B(net1262),
    .Y(_1882_));
 sg13g2_xor2_1 _5813_ (.B(_1882_),
    .A(_1272_),
    .X(\scl_uarttx0.scl_baudrategenerator0.n6892_o[3] ));
 sg13g2_nor2_1 _5814_ (.A(_1273_),
    .B(net1261),
    .Y(_1883_));
 sg13g2_nand2b_1 _5815_ (.Y(_1884_),
    .B(_1883_),
    .A_N(_1274_));
 sg13g2_xnor2_1 _5816_ (.Y(\scl_uarttx0.scl_baudrategenerator0.n6892_o[4] ),
    .A(_1274_),
    .B(_1883_));
 sg13g2_a22oi_1 _5817_ (.Y(\scl_uarttx0.scl_baudrategenerator0.n6892_o[5] ),
    .B1(_1884_),
    .B2(_1276_),
    .A2(_1883_),
    .A1(_1277_));
 sg13g2_nor2_1 _5818_ (.A(_1278_),
    .B(net1261),
    .Y(_1885_));
 sg13g2_xnor2_1 _5819_ (.Y(\scl_uarttx0.scl_baudrategenerator0.n6892_o[6] ),
    .A(_1268_),
    .B(_1885_));
 sg13g2_nand2b_1 _5820_ (.Y(_1886_),
    .B(_1885_),
    .A_N(_1279_));
 sg13g2_a21o_1 _5821_ (.A2(_1885_),
    .A1(_1268_),
    .B1(_1267_),
    .X(_1887_));
 sg13g2_nand2_1 _5822_ (.Y(\scl_uarttx0.scl_baudrategenerator0.n6892_o[7] ),
    .A(_1886_),
    .B(_1887_));
 sg13g2_xnor2_1 _5823_ (.Y(\scl_uarttx0.scl_baudrategenerator0.n6892_o[8] ),
    .A(_1266_),
    .B(_1886_));
 sg13g2_nor2_1 _5824_ (.A(_1280_),
    .B(net1261),
    .Y(_1888_));
 sg13g2_xor2_1 _5825_ (.B(_1888_),
    .A(_1264_),
    .X(\scl_uarttx0.scl_baudrategenerator0.n6892_o[9] ));
 sg13g2_nor2_1 _5826_ (.A(_1282_),
    .B(net1262),
    .Y(_1889_));
 sg13g2_a21oi_1 _5827_ (.A1(_1264_),
    .A2(_1888_),
    .Y(_1890_),
    .B1(_1265_));
 sg13g2_nor2_1 _5828_ (.A(_1889_),
    .B(_1890_),
    .Y(\scl_uarttx0.scl_baudrategenerator0.n6892_o[10] ));
 sg13g2_xnor2_1 _5829_ (.Y(\scl_uarttx0.scl_baudrategenerator0.n6892_o[11] ),
    .A(_1284_),
    .B(_1889_));
 sg13g2_nor2_1 _5830_ (.A(_1285_),
    .B(net1261),
    .Y(_1891_));
 sg13g2_xnor2_1 _5831_ (.Y(\scl_uarttx0.scl_baudrategenerator0.n6892_o[12] ),
    .A(_1261_),
    .B(_1891_));
 sg13g2_nor3_1 _5832_ (.A(_1286_),
    .B(_1292_),
    .C(net1261),
    .Y(_1892_));
 sg13g2_o21ai_1 _5833_ (.B1(_1292_),
    .Y(_1893_),
    .A1(_1286_),
    .A2(net1261));
 sg13g2_nor2b_1 _5834_ (.A(_1892_),
    .B_N(_1893_),
    .Y(\scl_uarttx0.scl_baudrategenerator0.n6892_o[13] ));
 sg13g2_xor2_1 _5835_ (.B(_1892_),
    .A(_1298_),
    .X(\scl_uarttx0.scl_baudrategenerator0.n6892_o[14] ));
 sg13g2_a21oi_1 _5836_ (.A1(_1287_),
    .A2(_1299_),
    .Y(_1894_),
    .B1(net1261));
 sg13g2_xnor2_1 _5837_ (.Y(\scl_uarttx0.scl_baudrategenerator0.n6892_o[15] ),
    .A(_1305_),
    .B(_1894_));
 sg13g2_nor2_1 _5838_ (.A(_1306_),
    .B(net1261),
    .Y(_1895_));
 sg13g2_mux2_1 _5839_ (.A0(_1306_),
    .A1(_1895_),
    .S(_1314_),
    .X(\scl_uarttx0.scl_baudrategenerator0.n6892_o[16] ));
 sg13g2_nor2_1 _5840_ (.A(net721),
    .B(net1370),
    .Y(\scl_bitbangengine0.scl_counter0.n6954_o[0] ));
 sg13g2_nand2_1 _5841_ (.Y(_1896_),
    .A(net721),
    .B(net1868));
 sg13g2_or2_1 _5842_ (.X(_1897_),
    .B(net1868),
    .A(net721));
 sg13g2_and3_1 _5843_ (.X(\scl_bitbangengine0.scl_counter0.n6954_o[1] ),
    .A(_1177_),
    .B(_1896_),
    .C(_1897_));
 sg13g2_and2_1 _5844_ (.A(net1657),
    .B(_1896_),
    .X(_1898_));
 sg13g2_nor2_1 _5845_ (.A(net1657),
    .B(_1896_),
    .Y(_1899_));
 sg13g2_nor3_1 _5846_ (.A(net1370),
    .B(net1658),
    .C(_1899_),
    .Y(\scl_bitbangengine0.scl_counter0.n6954_o[2] ));
 sg13g2_xor2_1 _5847_ (.B(_1899_),
    .A(net1600),
    .X(_1900_));
 sg13g2_nor2_1 _5848_ (.A(net1370),
    .B(net1601),
    .Y(\scl_bitbangengine0.scl_counter0.n6954_o[3] ));
 sg13g2_nand4_1 _5849_ (.B(\scl_bitbangengine0.scl_counter0.n6975_q[1] ),
    .C(\scl_bitbangengine0.scl_counter0.n6975_q[2] ),
    .A(\scl_bitbangengine0.scl_counter0.n6975_q[0] ),
    .Y(_1901_),
    .D(\scl_bitbangengine0.scl_counter0.n6975_q[3] ));
 sg13g2_and2_1 _5850_ (.A(net1705),
    .B(_1901_),
    .X(_1902_));
 sg13g2_nor2_1 _5851_ (.A(net1705),
    .B(_1901_),
    .Y(_1903_));
 sg13g2_nor3_1 _5852_ (.A(net1369),
    .B(net1706),
    .C(_1903_),
    .Y(\scl_bitbangengine0.scl_counter0.n6954_o[4] ));
 sg13g2_xor2_1 _5853_ (.B(_1903_),
    .A(net1079),
    .X(_1904_));
 sg13g2_nor2_1 _5854_ (.A(net1369),
    .B(net1080),
    .Y(\scl_bitbangengine0.scl_counter0.n6954_o[5] ));
 sg13g2_nand2_1 _5855_ (.Y(_1905_),
    .A(\scl_bitbangengine0.scl_counter0.n6975_q[4] ),
    .B(\scl_bitbangengine0.scl_counter0.n6975_q[5] ));
 sg13g2_nor2_1 _5856_ (.A(_1901_),
    .B(_1905_),
    .Y(_1906_));
 sg13g2_nor2b_1 _5857_ (.A(_1906_),
    .B_N(net1728),
    .Y(_1907_));
 sg13g2_nor3_1 _5858_ (.A(net1728),
    .B(_1901_),
    .C(_1905_),
    .Y(_1908_));
 sg13g2_nor3_1 _5859_ (.A(net1369),
    .B(net1729),
    .C(_1908_),
    .Y(\scl_bitbangengine0.scl_counter0.n6954_o[6] ));
 sg13g2_xnor2_1 _5860_ (.Y(_1909_),
    .A(net1749),
    .B(_1908_));
 sg13g2_nor2b_1 _5861_ (.A(net1369),
    .B_N(net1750),
    .Y(\scl_bitbangengine0.scl_counter0.n6954_o[7] ));
 sg13g2_nand3_1 _5862_ (.B(\scl_bitbangengine0.scl_counter0.n6975_q[7] ),
    .C(_1906_),
    .A(\scl_bitbangengine0.scl_counter0.n6975_q[6] ),
    .Y(_1910_));
 sg13g2_and2_1 _5863_ (.A(net1813),
    .B(_1910_),
    .X(_1911_));
 sg13g2_nor2_1 _5864_ (.A(net1813),
    .B(_1910_),
    .Y(_1912_));
 sg13g2_nor3_1 _5865_ (.A(net1369),
    .B(net1814),
    .C(_1912_),
    .Y(\scl_bitbangengine0.scl_counter0.n6954_o[8] ));
 sg13g2_xor2_1 _5866_ (.B(_1912_),
    .A(net1661),
    .X(_1913_));
 sg13g2_nor2_1 _5867_ (.A(net1370),
    .B(net1662),
    .Y(\scl_bitbangengine0.scl_counter0.n6954_o[9] ));
 sg13g2_nand2_1 _5868_ (.Y(_1914_),
    .A(\scl_bitbangengine0.scl_counter0.n6975_q[8] ),
    .B(\scl_bitbangengine0.scl_counter0.n6975_q[9] ));
 sg13g2_nor2_1 _5869_ (.A(_1910_),
    .B(_1914_),
    .Y(_1915_));
 sg13g2_nor2b_1 _5870_ (.A(_1915_),
    .B_N(net1746),
    .Y(_1916_));
 sg13g2_nor3_1 _5871_ (.A(net1746),
    .B(_1910_),
    .C(_1914_),
    .Y(_1917_));
 sg13g2_nor3_1 _5872_ (.A(net1369),
    .B(net1747),
    .C(_1917_),
    .Y(\scl_bitbangengine0.scl_counter0.n6954_o[10] ));
 sg13g2_xor2_1 _5873_ (.B(_1917_),
    .A(net1585),
    .X(_1918_));
 sg13g2_nor2_1 _5874_ (.A(net1370),
    .B(net1586),
    .Y(\scl_bitbangengine0.scl_counter0.n6954_o[11] ));
 sg13g2_and2_1 _5875_ (.A(\scl_bitbangengine0.scl_counter0.n6975_q[10] ),
    .B(\scl_bitbangengine0.scl_counter0.n6975_q[11] ),
    .X(_1919_));
 sg13g2_nand2_1 _5876_ (.Y(_1920_),
    .A(_1915_),
    .B(_1919_));
 sg13g2_and2_1 _5877_ (.A(net1796),
    .B(_1920_),
    .X(_1921_));
 sg13g2_nor2_1 _5878_ (.A(net1796),
    .B(_1920_),
    .Y(_1922_));
 sg13g2_nor3_1 _5879_ (.A(net1369),
    .B(net1797),
    .C(_1922_),
    .Y(\scl_bitbangengine0.scl_counter0.n6954_o[12] ));
 sg13g2_xor2_1 _5880_ (.B(_1922_),
    .A(net1039),
    .X(_1923_));
 sg13g2_nor2_1 _5881_ (.A(net1369),
    .B(net1040),
    .Y(\scl_bitbangengine0.scl_counter0.n6954_o[13] ));
 sg13g2_nand4_1 _5882_ (.B(\scl_bitbangengine0.scl_counter0.n6975_q[13] ),
    .C(_1915_),
    .A(\scl_bitbangengine0.scl_counter0.n6975_q[12] ),
    .Y(_1924_),
    .D(_1919_));
 sg13g2_inv_1 _5883_ (.Y(_1925_),
    .A(_1924_));
 sg13g2_and2_1 _5884_ (.A(net1607),
    .B(_1924_),
    .X(_1926_));
 sg13g2_nor2_1 _5885_ (.A(net1607),
    .B(_1924_),
    .Y(_1927_));
 sg13g2_nor3_1 _5886_ (.A(net1371),
    .B(net1608),
    .C(_1927_),
    .Y(\scl_bitbangengine0.scl_counter0.n6954_o[14] ));
 sg13g2_xor2_1 _5887_ (.B(_1927_),
    .A(net1781),
    .X(_1928_));
 sg13g2_nor2_1 _5888_ (.A(net1370),
    .B(net1782),
    .Y(\scl_bitbangengine0.scl_counter0.n6954_o[15] ));
 sg13g2_nand3_1 _5889_ (.B(\scl_bitbangengine0.scl_counter0.n6975_q[15] ),
    .C(_1925_),
    .A(\scl_bitbangengine0.scl_counter0.n6975_q[14] ),
    .Y(_1929_));
 sg13g2_xnor2_1 _5890_ (.Y(_1930_),
    .A(net985),
    .B(_1929_));
 sg13g2_nor2_1 _5891_ (.A(net1370),
    .B(net986),
    .Y(\scl_bitbangengine0.scl_counter0.n6954_o[16] ));
 sg13g2_nand2_1 _5892_ (.Y(_1931_),
    .A(net931),
    .B(_1214_));
 sg13g2_nor2_2 _5893_ (.A(\scl_bitbangengine0.n5915_q ),
    .B(_1214_),
    .Y(_1932_));
 sg13g2_nor2_1 _5894_ (.A(_0690_),
    .B(\scl_bitbangengine0.n5909_q ),
    .Y(_1933_));
 sg13g2_a21oi_1 _5895_ (.A1(net10),
    .A2(\scl_bitbangengine0.n5909_q ),
    .Y(_1934_),
    .B1(_1933_));
 sg13g2_nor2_2 _5896_ (.A(_0772_),
    .B(net1269),
    .Y(_1935_));
 sg13g2_a22oi_1 _5897_ (.Y(_1936_),
    .B1(_1934_),
    .B2(_1935_),
    .A2(_1932_),
    .A1(_0135_));
 sg13g2_and3_1 _5898_ (.X(\scl_bitbangengine0.n5462_o[0] ),
    .A(_1215_),
    .B(_1931_),
    .C(_1936_));
 sg13g2_nand2_1 _5899_ (.Y(_1937_),
    .A(net1146),
    .B(_1214_));
 sg13g2_a22oi_1 _5900_ (.Y(_1938_),
    .B1(_1935_),
    .B2(net931),
    .A2(_1932_),
    .A1(_0136_));
 sg13g2_and3_1 _5901_ (.X(\scl_bitbangengine0.n5462_o[1] ),
    .A(net1265),
    .B(_1937_),
    .C(_1938_));
 sg13g2_nand2_1 _5902_ (.Y(_1939_),
    .A(net1563),
    .B(net1269));
 sg13g2_a22oi_1 _5903_ (.Y(_1940_),
    .B1(_1935_),
    .B2(net1146),
    .A2(_1932_),
    .A1(_0137_));
 sg13g2_and3_1 _5904_ (.X(\scl_bitbangengine0.n5462_o[2] ),
    .A(net1265),
    .B(_1939_),
    .C(_1940_));
 sg13g2_nand2_1 _5905_ (.Y(_1941_),
    .A(net1663),
    .B(net1269));
 sg13g2_a22oi_1 _5906_ (.Y(_1942_),
    .B1(_1935_),
    .B2(net1563),
    .A2(_1932_),
    .A1(net1590));
 sg13g2_and3_1 _5907_ (.X(\scl_bitbangengine0.n5462_o[3] ),
    .A(net1265),
    .B(_1941_),
    .C(_1942_));
 sg13g2_nand2_1 _5908_ (.Y(_1943_),
    .A(net1590),
    .B(net1269));
 sg13g2_a22oi_1 _5909_ (.Y(_1944_),
    .B1(_1935_),
    .B2(_0137_),
    .A2(_1932_),
    .A1(net1135));
 sg13g2_and3_1 _5910_ (.X(\scl_bitbangengine0.n5462_o[4] ),
    .A(net1265),
    .B(_1943_),
    .C(_1944_));
 sg13g2_nand2_1 _5911_ (.Y(_1945_),
    .A(net1135),
    .B(net1269));
 sg13g2_a22oi_1 _5912_ (.Y(_1946_),
    .B1(_1935_),
    .B2(_0138_),
    .A2(_1932_),
    .A1(_0140_));
 sg13g2_and3_1 _5913_ (.X(\scl_bitbangengine0.n5462_o[5] ),
    .A(net1265),
    .B(_1945_),
    .C(_1946_));
 sg13g2_o21ai_1 _5914_ (.B1(net1265),
    .Y(_1947_),
    .A1(_0774_),
    .A2(net1271));
 sg13g2_nor3_1 _5915_ (.A(\scl_bitbangengine0.n5915_q ),
    .B(\scl_bitbangengine0.n5924_q[7] ),
    .C(net1269),
    .Y(_1948_));
 sg13g2_a21o_1 _5916_ (.A2(_1935_),
    .A1(net1135),
    .B1(_1948_),
    .X(_1949_));
 sg13g2_nor2_1 _5917_ (.A(_1947_),
    .B(_1949_),
    .Y(\scl_bitbangengine0.n5462_o[6] ));
 sg13g2_o21ai_1 _5918_ (.B1(net1265),
    .Y(_1950_),
    .A1(net1651),
    .A2(net1271));
 sg13g2_a22oi_1 _5919_ (.Y(_1951_),
    .B1(_1935_),
    .B2(_0773_),
    .A2(_1934_),
    .A1(_1932_));
 sg13g2_nor2b_1 _5920_ (.A(_1950_),
    .B_N(_1951_),
    .Y(\scl_bitbangengine0.n5462_o[7] ));
 sg13g2_nand2_2 _5921_ (.Y(_1952_),
    .A(net1503),
    .B(\scl_bitbangengine0.n5898_q[1] ));
 sg13g2_nor2_1 _5922_ (.A(_1194_),
    .B(_1952_),
    .Y(_1953_));
 sg13g2_nand2_1 _5923_ (.Y(_1954_),
    .A(net1371),
    .B(_1953_));
 sg13g2_nor2b_1 _5924_ (.A(_1197_),
    .B_N(_1954_),
    .Y(_1955_));
 sg13g2_o21ai_1 _5925_ (.B1(_1955_),
    .Y(_1956_),
    .A1(\scl_bitbangengine0.n5913_q ),
    .A2(_1211_));
 sg13g2_nand2b_1 _5926_ (.Y(_1957_),
    .B(net1088),
    .A_N(net859));
 sg13g2_o21ai_1 _5927_ (.B1(_1957_),
    .Y(_1958_),
    .A1(net1088),
    .A2(_1956_));
 sg13g2_nor2_1 _5928_ (.A(_1177_),
    .B(_1958_),
    .Y(_1959_));
 sg13g2_xor2_1 _5929_ (.B(_1959_),
    .A(_1204_),
    .X(\scl_bitbangengine0.n5401_o ));
 sg13g2_nor2_1 _5930_ (.A(net1692),
    .B(_1100_),
    .Y(_1960_));
 sg13g2_a21oi_1 _5931_ (.A1(_0730_),
    .A2(_1100_),
    .Y(\scl_bitbangengine0.n3871_o ),
    .B1(_1960_));
 sg13g2_mux2_1 _5932_ (.A0(net1066),
    .A1(net1496),
    .S(_1202_),
    .X(\scl_bitbangengine0.n3839_o ));
 sg13g2_xnor2_1 _5933_ (.Y(_1961_),
    .A(_0709_),
    .B(\n352_o[7] ));
 sg13g2_nand2_1 _5934_ (.Y(\scl_uartrx0.scl_baudrategenerator0.n7069_o[0] ),
    .A(net1434),
    .B(net1589));
 sg13g2_nand2b_1 _5935_ (.Y(_1962_),
    .B(_0922_),
    .A_N(_0888_));
 sg13g2_o21ai_1 _5936_ (.B1(_0888_),
    .Y(_1963_),
    .A1(net1435),
    .A2(net1241));
 sg13g2_a21o_1 _5937_ (.A2(_1963_),
    .A1(_1962_),
    .B1(net1435),
    .X(\scl_uartrx0.scl_baudrategenerator0.n7069_o[1] ));
 sg13g2_a221oi_1 _5938_ (.B2(_0887_),
    .C1(net1435),
    .B1(_1962_),
    .A1(_0889_),
    .Y(\scl_uartrx0.scl_baudrategenerator0.n7069_o[2] ),
    .A2(net1259));
 sg13g2_o21ai_1 _5939_ (.B1(_0890_),
    .Y(_1964_),
    .A1(_0889_),
    .A2(net1241));
 sg13g2_or3_1 _5940_ (.A(_0889_),
    .B(_0890_),
    .C(net1241),
    .X(_1965_));
 sg13g2_nand3_1 _5941_ (.B(_1964_),
    .C(_1965_),
    .A(net1434),
    .Y(\scl_uartrx0.scl_baudrategenerator0.n7069_o[3] ));
 sg13g2_nor2_1 _5942_ (.A(_0891_),
    .B(net1241),
    .Y(_1966_));
 sg13g2_nand2_1 _5943_ (.Y(_1967_),
    .A(_0892_),
    .B(net1259));
 sg13g2_xnor2_1 _5944_ (.Y(_1968_),
    .A(_0886_),
    .B(_1966_));
 sg13g2_nand2_1 _5945_ (.Y(\scl_uartrx0.scl_baudrategenerator0.n7069_o[4] ),
    .A(net1434),
    .B(_1968_));
 sg13g2_o21ai_1 _5946_ (.B1(net1434),
    .Y(_1969_),
    .A1(_0885_),
    .A2(_1967_));
 sg13g2_a21oi_1 _5947_ (.A1(_0885_),
    .A2(_1967_),
    .Y(\scl_uartrx0.scl_baudrategenerator0.n7069_o[5] ),
    .B1(_1969_));
 sg13g2_nor2_1 _5948_ (.A(_0893_),
    .B(net1241),
    .Y(_1970_));
 sg13g2_o21ai_1 _5949_ (.B1(net1434),
    .Y(_1971_),
    .A1(_0894_),
    .A2(_1970_));
 sg13g2_a21oi_1 _5950_ (.A1(_0894_),
    .A2(_1970_),
    .Y(\scl_uartrx0.scl_baudrategenerator0.n7069_o[6] ),
    .B1(_1971_));
 sg13g2_nand2_1 _5951_ (.Y(_1972_),
    .A(_0896_),
    .B(_0922_));
 sg13g2_a21o_1 _5952_ (.A2(_0922_),
    .A1(_0895_),
    .B1(_0884_),
    .X(_1973_));
 sg13g2_a21oi_1 _5953_ (.A1(_1972_),
    .A2(_1973_),
    .Y(\scl_uartrx0.scl_baudrategenerator0.n7069_o[7] ),
    .B1(net1435));
 sg13g2_a21oi_1 _5954_ (.A1(_0883_),
    .A2(_1972_),
    .Y(_1974_),
    .B1(net1435));
 sg13g2_o21ai_1 _5955_ (.B1(_1974_),
    .Y(\scl_uartrx0.scl_baudrategenerator0.n7069_o[8] ),
    .A1(_0897_),
    .A2(net1241));
 sg13g2_a21oi_1 _5956_ (.A1(_0897_),
    .A2(net1259),
    .Y(_1975_),
    .B1(_0899_));
 sg13g2_and3_1 _5957_ (.X(_1976_),
    .A(_0897_),
    .B(_0899_),
    .C(net1259));
 sg13g2_o21ai_1 _5958_ (.B1(net1434),
    .Y(\scl_uartrx0.scl_baudrategenerator0.n7069_o[9] ),
    .A1(_1975_),
    .A2(_1976_));
 sg13g2_nand2_1 _5959_ (.Y(_1977_),
    .A(_0901_),
    .B(_0922_));
 sg13g2_a221oi_1 _5960_ (.B2(_0900_),
    .C1(_1976_),
    .B1(_0855_),
    .A1(net598),
    .Y(_1978_),
    .A2(_0802_));
 sg13g2_a21oi_1 _5961_ (.A1(_0901_),
    .A2(_0922_),
    .Y(\scl_uartrx0.scl_baudrategenerator0.n7069_o[10] ),
    .B1(_1978_));
 sg13g2_a221oi_1 _5962_ (.B2(_0882_),
    .C1(net1435),
    .B1(_1977_),
    .A1(_0902_),
    .Y(\scl_uartrx0.scl_baudrategenerator0.n7069_o[11] ),
    .A2(net1259));
 sg13g2_nor2_1 _5963_ (.A(_0902_),
    .B(net1241),
    .Y(_1979_));
 sg13g2_a21oi_1 _5964_ (.A1(_0879_),
    .A2(_1979_),
    .Y(_1980_),
    .B1(net1435));
 sg13g2_o21ai_1 _5965_ (.B1(_1980_),
    .Y(\scl_uartrx0.scl_baudrategenerator0.n7069_o[12] ),
    .A1(_0879_),
    .A2(_1979_));
 sg13g2_a21oi_1 _5966_ (.A1(_0904_),
    .A2(net1259),
    .Y(_1981_),
    .B1(_0907_));
 sg13g2_a22oi_1 _5967_ (.Y(\scl_uartrx0.scl_baudrategenerator0.n7069_o[13] ),
    .B1(_1981_),
    .B2(_0804_),
    .A2(_0922_),
    .A1(_0908_));
 sg13g2_a21oi_1 _5968_ (.A1(_0908_),
    .A2(_0922_),
    .Y(_1982_),
    .B1(_0877_));
 sg13g2_o21ai_1 _5969_ (.B1(_0804_),
    .Y(_1983_),
    .A1(_0909_),
    .A2(_0919_));
 sg13g2_nor2_1 _5970_ (.A(_1982_),
    .B(_1983_),
    .Y(\scl_uartrx0.scl_baudrategenerator0.n7069_o[14] ));
 sg13g2_a21oi_1 _5971_ (.A1(_0909_),
    .A2(net1259),
    .Y(_1984_),
    .B1(_0913_));
 sg13g2_nor2_1 _5972_ (.A(_0915_),
    .B(_0917_),
    .Y(_1985_));
 sg13g2_or3_1 _5973_ (.A(_0803_),
    .B(_1984_),
    .C(_1985_),
    .X(\scl_uartrx0.scl_baudrategenerator0.n7069_o[15] ));
 sg13g2_a21oi_1 _5974_ (.A1(_0915_),
    .A2(_0918_),
    .Y(_1986_),
    .B1(_0875_));
 sg13g2_nor3_1 _5975_ (.A(_0803_),
    .B(_0916_),
    .C(_1986_),
    .Y(\scl_uartrx0.scl_baudrategenerator0.n7069_o[16] ));
 sg13g2_nand2_2 _5976_ (.Y(_1987_),
    .A(net1423),
    .B(_1006_));
 sg13g2_mux2_1 _5977_ (.A0(_1057_),
    .A1(net1611),
    .S(net1363),
    .X(\scl_fifo1.n6239_o[0] ));
 sg13g2_mux2_1 _5978_ (.A0(_1049_),
    .A1(net1144),
    .S(net1363),
    .X(\scl_fifo1.n6239_o[1] ));
 sg13g2_nand2_1 _5979_ (.Y(_1988_),
    .A(net892),
    .B(net1363));
 sg13g2_o21ai_1 _5980_ (.B1(_1988_),
    .Y(\scl_fifo1.n6239_o[2] ),
    .A1(_1063_),
    .A2(net1363));
 sg13g2_mux2_1 _5981_ (.A0(_1053_),
    .A1(net1603),
    .S(_1987_),
    .X(\scl_fifo1.n6239_o[3] ));
 sg13g2_mux2_1 _5982_ (.A0(_1045_),
    .A1(net1105),
    .S(_1987_),
    .X(\scl_fifo1.n6239_o[4] ));
 sg13g2_nand2_1 _5983_ (.Y(_1989_),
    .A(_0150_),
    .B(_1216_));
 sg13g2_xor2_1 _5984_ (.B(net1257),
    .A(net561),
    .X(\scl_fifo1.n6233_o[0] ));
 sg13g2_nand4_1 _5985_ (.B(_0150_),
    .C(\scl_fifo1.n6229_o[1] ),
    .A(\scl_fifo1.n6229_o[0] ),
    .Y(_1990_),
    .D(_1216_));
 sg13g2_or3_2 _5986_ (.A(\scl_fifo1.n6229_o[0] ),
    .B(\scl_fifo1.n6229_o[1] ),
    .C(net1257),
    .X(_1991_));
 sg13g2_nand2_1 _5987_ (.Y(_1992_),
    .A(_1990_),
    .B(_1991_));
 sg13g2_a21oi_1 _5988_ (.A1(net541),
    .A2(net1257),
    .Y(\scl_fifo1.n6233_o[1] ),
    .B1(_1992_));
 sg13g2_nor2_1 _5989_ (.A(_0153_),
    .B(_1990_),
    .Y(_1993_));
 sg13g2_xor2_1 _5990_ (.B(_1990_),
    .A(net651),
    .X(\scl_fifo1.n6233_o[2] ));
 sg13g2_xnor2_1 _5991_ (.Y(\scl_fifo1.n6233_o[3] ),
    .A(net581),
    .B(_1993_));
 sg13g2_nand2_2 _5992_ (.Y(_1994_),
    .A(\scl_fifo1.n6229_o[2] ),
    .B(\scl_fifo1.n6229_o[3] ));
 sg13g2_nor2_1 _5993_ (.A(_1990_),
    .B(_1994_),
    .Y(_1995_));
 sg13g2_xnor2_1 _5994_ (.Y(\scl_fifo1.n6233_o[4] ),
    .A(net1024),
    .B(net1224));
 sg13g2_nor2b_1 _5995_ (.A(s_m_io0_opendrain),
    .B_N(s_m_io0_out),
    .Y(n106_o));
 sg13g2_nor2b_1 _5996_ (.A(s_m_io2_opendrain),
    .B_N(s_m_io2_out),
    .Y(n118_o));
 sg13g2_nor2b_1 _5997_ (.A(s_m_io3_opendrain),
    .B_N(s_m_io3_out),
    .Y(n124_o));
 sg13g2_nor2b_1 _5998_ (.A(s_m_io4_opendrain),
    .B_N(s_m_io4_out),
    .Y(n130_o));
 sg13g2_nor2b_1 _5999_ (.A(s_m_io5_opendrain),
    .B_N(s_m_io5_out),
    .Y(n136_o));
 sg13g2_mux2_2 _6000_ (.A0(n153_o),
    .A1(n183_o),
    .S(_0724_),
    .X(uo_out[0]));
 sg13g2_mux2_2 _6001_ (.A0(s_m_io9_out),
    .A1(n350_o),
    .S(_0724_),
    .X(uo_out[1]));
 sg13g2_nand2b_1 _6002_ (.Y(_1996_),
    .B(s_m_io0_en),
    .A_N(_0119_));
 sg13g2_a21oi_2 _6003_ (.B1(_1996_),
    .Y(uio_oe[0]),
    .A2(s_m_io0_opendrain),
    .A1(s_m_io0_out));
 sg13g2_nand2_1 _6004_ (.Y(_1997_),
    .A(s_m_io1_out),
    .B(s_m_io1_opendrain));
 sg13g2_a21o_1 _6005_ (.A2(_1997_),
    .A1(s_m_io1_en),
    .B1(_0119_),
    .X(uio_oe[1]));
 sg13g2_nand2b_1 _6006_ (.Y(_1998_),
    .B(s_m_io2_en),
    .A_N(_0119_));
 sg13g2_a21oi_2 _6007_ (.B1(_1998_),
    .Y(uio_oe[2]),
    .A2(s_m_io2_opendrain),
    .A1(s_m_io2_out));
 sg13g2_nand2b_1 _6008_ (.Y(_1999_),
    .B(s_m_io3_en),
    .A_N(_0119_));
 sg13g2_a21oi_2 _6009_ (.B1(_1999_),
    .Y(uio_oe[3]),
    .A2(s_m_io3_opendrain),
    .A1(s_m_io3_out));
 sg13g2_nand2b_1 _6010_ (.Y(_2000_),
    .B(s_m_io4_en),
    .A_N(_0119_));
 sg13g2_a21oi_2 _6011_ (.B1(_2000_),
    .Y(uio_oe[4]),
    .A2(s_m_io4_opendrain),
    .A1(s_m_io4_out));
 sg13g2_nand2b_1 _6012_ (.Y(_2001_),
    .B(s_m_io5_en),
    .A_N(_0119_));
 sg13g2_a21oi_2 _6013_ (.B1(_2001_),
    .Y(uio_oe[5]),
    .A2(s_m_io5_opendrain),
    .A1(s_m_io5_out));
 sg13g2_mux4_1 _6014_ (.S0(\scl_uarttx0.n2856_o[1] ),
    .A0(net1502),
    .A1(net1498),
    .A2(net1493),
    .A3(\scl_bitbangengine0.n3258_o ),
    .S1(\scl_uarttx0.n2856_o[2] ),
    .X(_2002_));
 sg13g2_nand2b_1 _6015_ (.Y(_2003_),
    .B(_2002_),
    .A_N(\scl_uarttx0.n2856_o[0] ));
 sg13g2_nand2_1 _6016_ (.Y(_2004_),
    .A(\scl_bitbangengine0.n3267_o ),
    .B(_1322_));
 sg13g2_nand3_1 _6017_ (.B(\scl_uarttx0.n2856_o[0] ),
    .C(\scl_uarttx0.n2856_o[1] ),
    .A(net1497),
    .Y(_2005_));
 sg13g2_o21ai_1 _6018_ (.B1(_1322_),
    .Y(_2006_),
    .A1(net1501),
    .A2(\scl_uarttx0.n2856_o[2] ));
 sg13g2_a22oi_1 _6019_ (.Y(_2007_),
    .B1(_2005_),
    .B2(_2006_),
    .A2(_2004_),
    .A1(\scl_uarttx0.n2856_o[2] ));
 sg13g2_nand3b_1 _6020_ (.B(\scl_uarttx0.n2884_o ),
    .C(_2003_),
    .Y(_2008_),
    .A_N(_2007_));
 sg13g2_a22oi_1 _6021_ (.Y(_2009_),
    .B1(_2008_),
    .B2(_1320_),
    .A2(_1325_),
    .A1(net1492));
 sg13g2_nand3b_1 _6022_ (.B(s_m_io1_out),
    .C(n346_q),
    .Y(_2010_),
    .A_N(s_m_io1_opendrain));
 sg13g2_o21ai_1 _6023_ (.B1(_2010_),
    .Y(uio_out[1]),
    .A1(n346_q),
    .A2(_2009_));
 sg13g2_mux2_1 _6024_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[9][0] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[8][0] ),
    .S(net1229),
    .X(_2011_));
 sg13g2_nand2_1 _6025_ (.Y(_2012_),
    .A(net1235),
    .B(_2011_));
 sg13g2_mux2_1 _6026_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[11][0] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[10][0] ),
    .S(net1229),
    .X(_2013_));
 sg13g2_a21oi_1 _6027_ (.A1(net1191),
    .A2(_2013_),
    .Y(_2014_),
    .B1(net1180));
 sg13g2_mux2_1 _6028_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[13][0] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[12][0] ),
    .S(net1226),
    .X(_2015_));
 sg13g2_mux2_1 _6029_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[15][0] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[14][0] ),
    .S(net1228),
    .X(_2016_));
 sg13g2_nand2_1 _6030_ (.Y(_2017_),
    .A(net1191),
    .B(_2016_));
 sg13g2_a21oi_1 _6031_ (.A1(net1235),
    .A2(_2015_),
    .Y(_2018_),
    .B1(net1189));
 sg13g2_a22oi_1 _6032_ (.Y(_2019_),
    .B1(_2017_),
    .B2(_2018_),
    .A2(_2014_),
    .A1(_2012_));
 sg13g2_mux2_1 _6033_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[1][0] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[0][0] ),
    .S(net1230),
    .X(_2020_));
 sg13g2_nand2_1 _6034_ (.Y(_2021_),
    .A(net1239),
    .B(_2020_));
 sg13g2_mux2_1 _6035_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[3][0] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[2][0] ),
    .S(net1231),
    .X(_2022_));
 sg13g2_a21oi_1 _6036_ (.A1(net1193),
    .A2(_2022_),
    .Y(_2023_),
    .B1(net1181));
 sg13g2_mux2_1 _6037_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[5][0] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[4][0] ),
    .S(net1231),
    .X(_2024_));
 sg13g2_nand2_1 _6038_ (.Y(_2025_),
    .A(net1239),
    .B(_2024_));
 sg13g2_mux2_1 _6039_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[7][0] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[6][0] ),
    .S(net1231),
    .X(_2026_));
 sg13g2_a21oi_1 _6040_ (.A1(net1193),
    .A2(_2026_),
    .Y(_2027_),
    .B1(_1347_));
 sg13g2_a221oi_1 _6041_ (.B2(_2027_),
    .C1(net1174),
    .B1(_2025_),
    .A1(_2021_),
    .Y(_2028_),
    .A2(_2023_));
 sg13g2_a21o_2 _6042_ (.A2(_2019_),
    .A1(net1173),
    .B1(_2028_),
    .X(_0000_));
 sg13g2_mux2_1 _6043_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[9][1] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[8][1] ),
    .S(net1225),
    .X(_2029_));
 sg13g2_nand2_1 _6044_ (.Y(_2030_),
    .A(net1235),
    .B(_2029_));
 sg13g2_mux2_1 _6045_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[11][1] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[10][1] ),
    .S(net1225),
    .X(_2031_));
 sg13g2_a21oi_1 _6046_ (.A1(net1191),
    .A2(_2031_),
    .Y(_2032_),
    .B1(net1180));
 sg13g2_mux2_1 _6047_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[13][1] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[12][1] ),
    .S(net1227),
    .X(_2033_));
 sg13g2_mux2_1 _6048_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[15][1] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[14][1] ),
    .S(net1228),
    .X(_2034_));
 sg13g2_nand2_1 _6049_ (.Y(_2035_),
    .A(net1191),
    .B(_2034_));
 sg13g2_a21oi_1 _6050_ (.A1(net1235),
    .A2(_2033_),
    .Y(_2036_),
    .B1(net1189));
 sg13g2_a22oi_1 _6051_ (.Y(_2037_),
    .B1(_2035_),
    .B2(_2036_),
    .A2(_2032_),
    .A1(_2030_));
 sg13g2_mux2_1 _6052_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[1][1] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[0][1] ),
    .S(net1226),
    .X(_2038_));
 sg13g2_nand2_1 _6053_ (.Y(_2039_),
    .A(net1238),
    .B(_2038_));
 sg13g2_mux2_1 _6054_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[3][1] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[2][1] ),
    .S(net1233),
    .X(_2040_));
 sg13g2_a21oi_1 _6055_ (.A1(net1195),
    .A2(_2040_),
    .Y(_2041_),
    .B1(net1181));
 sg13g2_mux2_1 _6056_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[5][1] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[4][1] ),
    .S(net1230),
    .X(_2042_));
 sg13g2_nand2_1 _6057_ (.Y(_2043_),
    .A(net1238),
    .B(_2042_));
 sg13g2_mux2_1 _6058_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[7][1] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[6][1] ),
    .S(net1230),
    .X(_2044_));
 sg13g2_a21oi_1 _6059_ (.A1(net1193),
    .A2(_2044_),
    .Y(_2045_),
    .B1(_1347_));
 sg13g2_a221oi_1 _6060_ (.B2(_2045_),
    .C1(net1173),
    .B1(_2043_),
    .A1(_2039_),
    .Y(_2046_),
    .A2(_2041_));
 sg13g2_a21o_1 _6061_ (.A2(_2037_),
    .A1(net1173),
    .B1(_2046_),
    .X(_0001_));
 sg13g2_mux2_1 _6062_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[9][2] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[8][2] ),
    .S(net1227),
    .X(_2047_));
 sg13g2_nand2_1 _6063_ (.Y(_2048_),
    .A(_1341_),
    .B(_2047_));
 sg13g2_mux2_1 _6064_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[11][2] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[10][2] ),
    .S(net1227),
    .X(_2049_));
 sg13g2_a21oi_1 _6065_ (.A1(net1192),
    .A2(_2049_),
    .Y(_2050_),
    .B1(net1180));
 sg13g2_mux2_1 _6066_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[13][2] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[12][2] ),
    .S(net1227),
    .X(_2051_));
 sg13g2_mux2_1 _6067_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[15][2] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[14][2] ),
    .S(net1227),
    .X(_2052_));
 sg13g2_nand2_1 _6068_ (.Y(_2053_),
    .A(net1192),
    .B(_2052_));
 sg13g2_a21oi_1 _6069_ (.A1(net1237),
    .A2(_2051_),
    .Y(_2054_),
    .B1(net1189));
 sg13g2_a22oi_1 _6070_ (.Y(_2055_),
    .B1(_2053_),
    .B2(_2054_),
    .A2(_2050_),
    .A1(_2048_));
 sg13g2_mux2_1 _6071_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[1][2] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[0][2] ),
    .S(net1232),
    .X(_2056_));
 sg13g2_nand2_1 _6072_ (.Y(_2057_),
    .A(net1240),
    .B(_2056_));
 sg13g2_mux2_1 _6073_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[3][2] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[2][2] ),
    .S(net1233),
    .X(_2058_));
 sg13g2_a21oi_1 _6074_ (.A1(net1194),
    .A2(_2058_),
    .Y(_2059_),
    .B1(net1182));
 sg13g2_mux2_1 _6075_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[5][2] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[4][2] ),
    .S(net1233),
    .X(_2060_));
 sg13g2_nand2_1 _6076_ (.Y(_2061_),
    .A(net1240),
    .B(_2060_));
 sg13g2_mux2_1 _6077_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[7][2] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[6][2] ),
    .S(net1232),
    .X(_2062_));
 sg13g2_a21oi_1 _6078_ (.A1(net1194),
    .A2(_2062_),
    .Y(_2063_),
    .B1(net1190));
 sg13g2_a221oi_1 _6079_ (.B2(_2063_),
    .C1(net1175),
    .B1(_2061_),
    .A1(_2057_),
    .Y(_2064_),
    .A2(_2059_));
 sg13g2_a21o_1 _6080_ (.A2(_2055_),
    .A1(net1175),
    .B1(_2064_),
    .X(_0002_));
 sg13g2_mux2_1 _6081_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[9][3] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[8][3] ),
    .S(net1225),
    .X(_2065_));
 sg13g2_nand2_1 _6082_ (.Y(_2066_),
    .A(net1235),
    .B(_2065_));
 sg13g2_mux2_1 _6083_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[11][3] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[10][3] ),
    .S(net1226),
    .X(_2067_));
 sg13g2_a21oi_1 _6084_ (.A1(net1192),
    .A2(_2067_),
    .Y(_2068_),
    .B1(net1180));
 sg13g2_mux2_1 _6085_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[13][3] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[12][3] ),
    .S(net1227),
    .X(_2069_));
 sg13g2_mux2_1 _6086_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[15][3] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[14][3] ),
    .S(net1228),
    .X(_2070_));
 sg13g2_nand2_1 _6087_ (.Y(_2071_),
    .A(net1192),
    .B(_2070_));
 sg13g2_a21oi_1 _6088_ (.A1(net1237),
    .A2(_2069_),
    .Y(_2072_),
    .B1(net1189));
 sg13g2_a22oi_1 _6089_ (.Y(_2073_),
    .B1(_2071_),
    .B2(_2072_),
    .A2(_2068_),
    .A1(_2066_));
 sg13g2_mux2_1 _6090_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[1][3] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[0][3] ),
    .S(net1230),
    .X(_2074_));
 sg13g2_nand2_1 _6091_ (.Y(_2075_),
    .A(net1238),
    .B(_2074_));
 sg13g2_mux2_1 _6092_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[3][3] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[2][3] ),
    .S(net1233),
    .X(_2076_));
 sg13g2_a21oi_1 _6093_ (.A1(net1193),
    .A2(_2076_),
    .Y(_2077_),
    .B1(net1181));
 sg13g2_mux2_1 _6094_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[5][3] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[4][3] ),
    .S(net1231),
    .X(_2078_));
 sg13g2_nand2_1 _6095_ (.Y(_2079_),
    .A(net1239),
    .B(_2078_));
 sg13g2_mux2_1 _6096_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[7][3] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[6][3] ),
    .S(net1231),
    .X(_2080_));
 sg13g2_a21oi_1 _6097_ (.A1(net1194),
    .A2(_2080_),
    .Y(_2081_),
    .B1(net1190));
 sg13g2_a221oi_1 _6098_ (.B2(_2081_),
    .C1(net1173),
    .B1(_2079_),
    .A1(_2075_),
    .Y(_2082_),
    .A2(_2077_));
 sg13g2_a21o_1 _6099_ (.A2(_2073_),
    .A1(net1175),
    .B1(_2082_),
    .X(_0003_));
 sg13g2_mux2_1 _6100_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[9][4] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[8][4] ),
    .S(net1225),
    .X(_2083_));
 sg13g2_nand2_1 _6101_ (.Y(_2084_),
    .A(net1235),
    .B(_2083_));
 sg13g2_mux2_1 _6102_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[11][4] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[10][4] ),
    .S(net1225),
    .X(_2085_));
 sg13g2_a21oi_1 _6103_ (.A1(net1191),
    .A2(_2085_),
    .Y(_2086_),
    .B1(net1180));
 sg13g2_mux2_1 _6104_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[13][4] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[12][4] ),
    .S(net1225),
    .X(_2087_));
 sg13g2_mux2_1 _6105_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[15][4] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[14][4] ),
    .S(net1227),
    .X(_2088_));
 sg13g2_nand2_1 _6106_ (.Y(_2089_),
    .A(net1192),
    .B(_2088_));
 sg13g2_a21oi_1 _6107_ (.A1(net1236),
    .A2(_2087_),
    .Y(_2090_),
    .B1(net1189));
 sg13g2_a22oi_1 _6108_ (.Y(_2091_),
    .B1(_2089_),
    .B2(_2090_),
    .A2(_2086_),
    .A1(_2084_));
 sg13g2_mux2_1 _6109_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[1][4] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[0][4] ),
    .S(net1226),
    .X(_2092_));
 sg13g2_nand2_1 _6110_ (.Y(_2093_),
    .A(net1238),
    .B(_2092_));
 sg13g2_mux2_1 _6111_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[3][4] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[2][4] ),
    .S(net1233),
    .X(_2094_));
 sg13g2_a21oi_1 _6112_ (.A1(net1193),
    .A2(_2094_),
    .Y(_2095_),
    .B1(net1181));
 sg13g2_mux2_1 _6113_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[5][4] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[4][4] ),
    .S(net1230),
    .X(_2096_));
 sg13g2_nand2_1 _6114_ (.Y(_2097_),
    .A(net1238),
    .B(_2096_));
 sg13g2_mux2_1 _6115_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[7][4] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[6][4] ),
    .S(net1230),
    .X(_2098_));
 sg13g2_a21oi_1 _6116_ (.A1(net1193),
    .A2(_2098_),
    .Y(_2099_),
    .B1(net1190));
 sg13g2_a221oi_1 _6117_ (.B2(_2099_),
    .C1(net1173),
    .B1(_2097_),
    .A1(_2093_),
    .Y(_2100_),
    .A2(_2095_));
 sg13g2_a21o_1 _6118_ (.A2(_2091_),
    .A1(net1173),
    .B1(_2100_),
    .X(_0004_));
 sg13g2_mux2_1 _6119_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[9][5] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[8][5] ),
    .S(net1226),
    .X(_2101_));
 sg13g2_nand2_1 _6120_ (.Y(_2102_),
    .A(net1236),
    .B(_2101_));
 sg13g2_mux2_1 _6121_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[11][5] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[10][5] ),
    .S(net1226),
    .X(_2103_));
 sg13g2_a21oi_1 _6122_ (.A1(net1191),
    .A2(_2103_),
    .Y(_2104_),
    .B1(net1180));
 sg13g2_mux2_1 _6123_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[13][5] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[12][5] ),
    .S(net1226),
    .X(_2105_));
 sg13g2_mux2_1 _6124_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[15][5] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[14][5] ),
    .S(net1228),
    .X(_2106_));
 sg13g2_nand2_1 _6125_ (.Y(_2107_),
    .A(net1191),
    .B(_2106_));
 sg13g2_a21oi_1 _6126_ (.A1(net1236),
    .A2(_2105_),
    .Y(_2108_),
    .B1(net1189));
 sg13g2_a22oi_1 _6127_ (.Y(_2109_),
    .B1(_2107_),
    .B2(_2108_),
    .A2(_2104_),
    .A1(_2102_));
 sg13g2_mux2_1 _6128_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[1][5] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[0][5] ),
    .S(net1230),
    .X(_2110_));
 sg13g2_nand2_1 _6129_ (.Y(_2111_),
    .A(net1238),
    .B(_2110_));
 sg13g2_mux2_1 _6130_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[3][5] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[2][5] ),
    .S(net1233),
    .X(_2112_));
 sg13g2_a21oi_1 _6131_ (.A1(net1193),
    .A2(_2112_),
    .Y(_2113_),
    .B1(net1181));
 sg13g2_mux2_1 _6132_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[5][5] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[4][5] ),
    .S(net1231),
    .X(_2114_));
 sg13g2_nand2_1 _6133_ (.Y(_2115_),
    .A(net1239),
    .B(_2114_));
 sg13g2_mux2_1 _6134_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[7][5] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[6][5] ),
    .S(net1231),
    .X(_2116_));
 sg13g2_a21oi_1 _6135_ (.A1(net1194),
    .A2(_2116_),
    .Y(_2117_),
    .B1(net1190));
 sg13g2_a221oi_1 _6136_ (.B2(_2117_),
    .C1(net1174),
    .B1(_2115_),
    .A1(_2111_),
    .Y(_2118_),
    .A2(_2113_));
 sg13g2_a21o_1 _6137_ (.A2(_2109_),
    .A1(net1173),
    .B1(_2118_),
    .X(_0005_));
 sg13g2_mux4_1 _6138_ (.S0(\scl_fifo0.n2697_o[0] ),
    .A0(\scl_fifo0.scl_memory0.physical_memory0.memory[10][6] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[11][6] ),
    .A2(\scl_fifo0.scl_memory0.physical_memory0.memory[8][6] ),
    .A3(\scl_fifo0.scl_memory0.physical_memory0.memory[9][6] ),
    .S1(net1237),
    .X(_2119_));
 sg13g2_nor2_1 _6139_ (.A(net1182),
    .B(_2119_),
    .Y(_2120_));
 sg13g2_mux2_1 _6140_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[13][6] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[12][6] ),
    .S(net1229),
    .X(_2121_));
 sg13g2_nand2b_1 _6141_ (.Y(_2122_),
    .B(\scl_fifo0.n2697_o[0] ),
    .A_N(\scl_fifo0.scl_memory0.physical_memory0.memory[15][6] ));
 sg13g2_a21oi_1 _6142_ (.A1(_0775_),
    .A2(net1228),
    .Y(_2123_),
    .B1(net1237));
 sg13g2_a221oi_1 _6143_ (.B2(_2123_),
    .C1(net1190),
    .B1(_2122_),
    .A1(net1237),
    .Y(_2124_),
    .A2(_2121_));
 sg13g2_nor3_2 _6144_ (.A(_1350_),
    .B(_2120_),
    .C(_2124_),
    .Y(_2125_));
 sg13g2_mux2_1 _6145_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[1][6] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[0][6] ),
    .S(net1230),
    .X(_2126_));
 sg13g2_nand2_1 _6146_ (.Y(_2127_),
    .A(net1240),
    .B(_2126_));
 sg13g2_mux2_1 _6147_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[3][6] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[2][6] ),
    .S(net1233),
    .X(_2128_));
 sg13g2_a21oi_1 _6148_ (.A1(net1194),
    .A2(_2128_),
    .Y(_2129_),
    .B1(net1181));
 sg13g2_mux2_1 _6149_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[5][6] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[4][6] ),
    .S(net1234),
    .X(_2130_));
 sg13g2_nand2_1 _6150_ (.Y(_2131_),
    .A(net1240),
    .B(_2130_));
 sg13g2_mux2_1 _6151_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[7][6] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[6][6] ),
    .S(net1232),
    .X(_2132_));
 sg13g2_a21oi_1 _6152_ (.A1(net1195),
    .A2(_2132_),
    .Y(_2133_),
    .B1(net1190));
 sg13g2_a221oi_1 _6153_ (.B2(_2133_),
    .C1(net1175),
    .B1(_2131_),
    .A1(_2127_),
    .Y(_2134_),
    .A2(_2129_));
 sg13g2_or2_1 _6154_ (.X(_0006_),
    .B(_2134_),
    .A(_2125_));
 sg13g2_mux2_1 _6155_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[9][7] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[8][7] ),
    .S(net1225),
    .X(_2135_));
 sg13g2_nand2_1 _6156_ (.Y(_2136_),
    .A(net1235),
    .B(_2135_));
 sg13g2_mux2_1 _6157_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[11][7] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[10][7] ),
    .S(net1225),
    .X(_2137_));
 sg13g2_a21oi_1 _6158_ (.A1(net1191),
    .A2(_2137_),
    .Y(_2138_),
    .B1(net1180));
 sg13g2_mux2_1 _6159_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[13][7] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[12][7] ),
    .S(net1227),
    .X(_2139_));
 sg13g2_mux2_1 _6160_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[15][7] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[14][7] ),
    .S(net1228),
    .X(_2140_));
 sg13g2_nand2_1 _6161_ (.Y(_2141_),
    .A(net1192),
    .B(_2140_));
 sg13g2_a21oi_1 _6162_ (.A1(net1237),
    .A2(_2139_),
    .Y(_2142_),
    .B1(net1189));
 sg13g2_a22oi_1 _6163_ (.Y(_2143_),
    .B1(_2141_),
    .B2(_2142_),
    .A2(_2138_),
    .A1(_2136_));
 sg13g2_mux2_1 _6164_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[1][7] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[0][7] ),
    .S(net1232),
    .X(_2144_));
 sg13g2_nand2_1 _6165_ (.Y(_2145_),
    .A(net1238),
    .B(_2144_));
 sg13g2_mux2_1 _6166_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[3][7] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[2][7] ),
    .S(net1233),
    .X(_2146_));
 sg13g2_a21oi_1 _6167_ (.A1(net1194),
    .A2(_2146_),
    .Y(_2147_),
    .B1(net1181));
 sg13g2_mux2_1 _6168_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[5][7] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[4][7] ),
    .S(net1231),
    .X(_2148_));
 sg13g2_nand2_1 _6169_ (.Y(_2149_),
    .A(net1238),
    .B(_2148_));
 sg13g2_mux2_1 _6170_ (.A0(\scl_fifo0.scl_memory0.physical_memory0.memory[7][7] ),
    .A1(\scl_fifo0.scl_memory0.physical_memory0.memory[6][7] ),
    .S(net1232),
    .X(_2150_));
 sg13g2_a21oi_1 _6171_ (.A1(net1193),
    .A2(_2150_),
    .Y(_2151_),
    .B1(net1190));
 sg13g2_a221oi_1 _6172_ (.B2(_2151_),
    .C1(net1173),
    .B1(_2149_),
    .A1(_2145_),
    .Y(_2152_),
    .A2(_2147_));
 sg13g2_a21o_1 _6173_ (.A2(_2143_),
    .A1(net1174),
    .B1(_2152_),
    .X(_0007_));
 sg13g2_nor2_2 _6174_ (.A(\usbfunction0.functionreset0.in_unnamed_4[1] ),
    .B(\usbfunction0.functionreset0.in_unnamed_4[0] ),
    .Y(_2153_));
 sg13g2_or2_1 _6175_ (.X(_2154_),
    .B(\usbfunction0.functionreset0.in_unnamed_4[0] ),
    .A(\usbfunction0.functionreset0.in_unnamed_4[1] ));
 sg13g2_nand2_1 _6176_ (.Y(\usbfunction0.functionreset0.n6674_o[0] ),
    .A(net583),
    .B(_2153_));
 sg13g2_and2_1 _6177_ (.A(net1677),
    .B(net583),
    .X(_2155_));
 sg13g2_nor3_1 _6178_ (.A(_1542_),
    .B(_2154_),
    .C(_2155_),
    .Y(\usbfunction0.functionreset0.n6674_o[1] ));
 sg13g2_a21oi_1 _6179_ (.A1(net1754),
    .A2(_2155_),
    .Y(_2156_),
    .B1(_2154_));
 sg13g2_o21ai_1 _6180_ (.B1(_2156_),
    .Y(_2157_),
    .A1(net1754),
    .A2(_2155_));
 sg13g2_inv_1 _6181_ (.Y(\usbfunction0.functionreset0.n6674_o[2] ),
    .A(net1755));
 sg13g2_a21oi_1 _6182_ (.A1(\usbfunction0.functionreset0.n6707_q[2] ),
    .A2(_2155_),
    .Y(_2158_),
    .B1(net794));
 sg13g2_and3_1 _6183_ (.X(_2159_),
    .A(net794),
    .B(\usbfunction0.functionreset0.n6707_q[2] ),
    .C(_2155_));
 sg13g2_nor3_1 _6184_ (.A(_2154_),
    .B(net795),
    .C(_2159_),
    .Y(\usbfunction0.functionreset0.n6674_o[3] ));
 sg13g2_and2_1 _6185_ (.A(net1647),
    .B(_2159_),
    .X(_2160_));
 sg13g2_o21ai_1 _6186_ (.B1(_2153_),
    .Y(_2161_),
    .A1(net1647),
    .A2(_2159_));
 sg13g2_nor2_1 _6187_ (.A(_2160_),
    .B(net1648),
    .Y(\usbfunction0.functionreset0.n6674_o[4] ));
 sg13g2_and2_1 _6188_ (.A(net1679),
    .B(_2160_),
    .X(_2162_));
 sg13g2_o21ai_1 _6189_ (.B1(_2153_),
    .Y(_2163_),
    .A1(net1679),
    .A2(_2160_));
 sg13g2_nor2_1 _6190_ (.A(_2162_),
    .B(net1680),
    .Y(\usbfunction0.functionreset0.n6674_o[5] ));
 sg13g2_and2_1 _6191_ (.A(net1683),
    .B(_2162_),
    .X(_2164_));
 sg13g2_o21ai_1 _6192_ (.B1(_2153_),
    .Y(_2165_),
    .A1(net1683),
    .A2(_2162_));
 sg13g2_nor2_1 _6193_ (.A(_2164_),
    .B(net1684),
    .Y(\usbfunction0.functionreset0.n6674_o[6] ));
 sg13g2_and2_1 _6194_ (.A(net1700),
    .B(_2164_),
    .X(_2166_));
 sg13g2_o21ai_1 _6195_ (.B1(_2153_),
    .Y(_2167_),
    .A1(net1700),
    .A2(_2164_));
 sg13g2_nor2_1 _6196_ (.A(_2166_),
    .B(net1701),
    .Y(\usbfunction0.functionreset0.n6674_o[7] ));
 sg13g2_and2_1 _6197_ (.A(net1671),
    .B(_2166_),
    .X(_2168_));
 sg13g2_o21ai_1 _6198_ (.B1(_2153_),
    .Y(_2169_),
    .A1(net1671),
    .A2(_2166_));
 sg13g2_nor2_1 _6199_ (.A(_2168_),
    .B(net1672),
    .Y(\usbfunction0.functionreset0.n6674_o[8] ));
 sg13g2_o21ai_1 _6200_ (.B1(_2153_),
    .Y(_2170_),
    .A1(net603),
    .A2(_2168_));
 sg13g2_a21oi_1 _6201_ (.A1(net603),
    .A2(_2168_),
    .Y(\usbfunction0.functionreset0.n6674_o[9] ),
    .B1(_2170_));
 sg13g2_nor2b_2 _6202_ (.A(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7654_q[1] ),
    .B_N(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7654_q[0] ),
    .Y(_2171_));
 sg13g2_xnor2_1 _6203_ (.Y(_2172_),
    .A(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7654_q[1] ),
    .B(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7654_q[0] ));
 sg13g2_xor2_1 _6204_ (.B(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7654_q[0] ),
    .A(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7654_q[1] ),
    .X(_2173_));
 sg13g2_nand2_1 _6205_ (.Y(_2174_),
    .A(\usbfunction0.scl_usbgpiophy0.n6653_q ),
    .B(_2172_));
 sg13g2_nand2_1 _6206_ (.Y(_2175_),
    .A(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7657_q ),
    .B(_2173_));
 sg13g2_o21ai_1 _6207_ (.B1(_2175_),
    .Y(_2176_),
    .A1(_1355_),
    .A2(_2174_));
 sg13g2_nand2_1 _6208_ (.Y(_2177_),
    .A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.in_unnamed ),
    .B(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[0] ));
 sg13g2_o21ai_1 _6209_ (.B1(_2177_),
    .Y(_2178_),
    .A1(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.in_unnamed ),
    .A2(_0715_));
 sg13g2_nor2_1 _6210_ (.A(_2176_),
    .B(_2178_),
    .Y(_2179_));
 sg13g2_mux2_1 _6211_ (.A0(_2179_),
    .A1(_1533_),
    .S(_0780_),
    .X(_2180_));
 sg13g2_nand2_1 _6212_ (.Y(_2181_),
    .A(_0779_),
    .B(_2180_));
 sg13g2_xor2_1 _6213_ (.B(_2181_),
    .A(\usbfunction0.scl_usbgpiophy0.nrzi0.n7721_q ),
    .X(_2182_));
 sg13g2_nor2b_1 _6214_ (.A(\usbfunction0.scl_usbgpiophy0.n6655_q ),
    .B_N(_2182_),
    .Y(\usbfunction0.scl_usbgpiophy0.n6500_o ));
 sg13g2_nor2_1 _6215_ (.A(\usbfunction0.scl_usbgpiophy0.n6655_q ),
    .B(_2182_),
    .Y(\usbfunction0.scl_usbgpiophy0.n6503_o ));
 sg13g2_mux2_1 _6216_ (.A0(\scl_fifo1.scl_memory0.physical_memory0.memory[0][0] ),
    .A1(\scl_fifo1.scl_memory0.physical_memory0.memory[1][0] ),
    .S(net1288),
    .X(_2183_));
 sg13g2_and2_1 _6217_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[3][0] ),
    .B(net1288),
    .X(_2184_));
 sg13g2_a21oi_1 _6218_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[2][0] ),
    .A2(net1321),
    .Y(_2185_),
    .B1(_2184_));
 sg13g2_a21oi_1 _6219_ (.A1(net1300),
    .A2(_2185_),
    .Y(_2186_),
    .B1(net1273));
 sg13g2_o21ai_1 _6220_ (.B1(_2186_),
    .Y(_2187_),
    .A1(net1300),
    .A2(_2183_));
 sg13g2_nand2_1 _6221_ (.Y(_2188_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[4][0] ),
    .B(net1325));
 sg13g2_a21oi_1 _6222_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[5][0] ),
    .A2(net1288),
    .Y(_2189_),
    .B1(net1303));
 sg13g2_and2_1 _6223_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[7][0] ),
    .B(net1289),
    .X(_2190_));
 sg13g2_a21oi_1 _6224_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[6][0] ),
    .A2(net1321),
    .Y(_2191_),
    .B1(_2190_));
 sg13g2_a221oi_1 _6225_ (.B2(net1303),
    .C1(net1280),
    .B1(_2191_),
    .A1(_2188_),
    .Y(_2192_),
    .A2(_2189_));
 sg13g2_nor2_1 _6226_ (.A(net1266),
    .B(_2192_),
    .Y(_2193_));
 sg13g2_nand2_1 _6227_ (.Y(_2194_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[12][0] ),
    .B(net1319));
 sg13g2_a21oi_1 _6228_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[13][0] ),
    .A2(net1285),
    .Y(_2195_),
    .B1(net1298));
 sg13g2_and2_1 _6229_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[15][0] ),
    .B(net1285),
    .X(_2196_));
 sg13g2_a21oi_1 _6230_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[14][0] ),
    .A2(net1319),
    .Y(_2197_),
    .B1(_2196_));
 sg13g2_a221oi_1 _6231_ (.B2(net1298),
    .C1(net1281),
    .B1(_2197_),
    .A1(_2194_),
    .Y(_2198_),
    .A2(_2195_));
 sg13g2_mux2_1 _6232_ (.A0(\scl_fifo1.scl_memory0.physical_memory0.memory[8][0] ),
    .A1(\scl_fifo1.scl_memory0.physical_memory0.memory[9][0] ),
    .S(net1283),
    .X(_2199_));
 sg13g2_and2_1 _6233_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[11][0] ),
    .B(net1282),
    .X(_2200_));
 sg13g2_a21oi_1 _6234_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[10][0] ),
    .A2(net1317),
    .Y(_2201_),
    .B1(_2200_));
 sg13g2_a21oi_1 _6235_ (.A1(net1294),
    .A2(_2201_),
    .Y(_2202_),
    .B1(net1272));
 sg13g2_o21ai_1 _6236_ (.B1(_2202_),
    .Y(_2203_),
    .A1(net1294),
    .A2(_2199_));
 sg13g2_nor2_1 _6237_ (.A(net1274),
    .B(_2198_),
    .Y(_2204_));
 sg13g2_a22oi_1 _6238_ (.Y(_0008_),
    .B1(_2203_),
    .B2(_2204_),
    .A2(_2193_),
    .A1(_2187_));
 sg13g2_and2_1 _6239_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[3][1] ),
    .B(net1292),
    .X(_2205_));
 sg13g2_a21oi_1 _6240_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[2][1] ),
    .A2(net1324),
    .Y(_2206_),
    .B1(_2205_));
 sg13g2_nand2_1 _6241_ (.Y(_2207_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[0][1] ),
    .B(net1322));
 sg13g2_a21oi_1 _6242_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[1][1] ),
    .A2(net1290),
    .Y(_2208_),
    .B1(net1300));
 sg13g2_a221oi_1 _6243_ (.B2(_2208_),
    .C1(\scl_fifo1.n6238_o[2] ),
    .B1(_2207_),
    .A1(net1300),
    .Y(_2209_),
    .A2(_2206_));
 sg13g2_nand2_1 _6244_ (.Y(_2210_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[4][1] ),
    .B(net1324));
 sg13g2_a21oi_1 _6245_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[5][1] ),
    .A2(net1292),
    .Y(_2211_),
    .B1(net1301));
 sg13g2_and2_1 _6246_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[7][1] ),
    .B(net1291),
    .X(_2212_));
 sg13g2_a21oi_1 _6247_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[6][1] ),
    .A2(net1324),
    .Y(_2213_),
    .B1(_2212_));
 sg13g2_a221oi_1 _6248_ (.B2(net1301),
    .C1(net1280),
    .B1(_2213_),
    .A1(_2210_),
    .Y(_2214_),
    .A2(_2211_));
 sg13g2_nor3_2 _6249_ (.A(\scl_fifo1.n6238_o[3] ),
    .B(_2209_),
    .C(_2214_),
    .Y(_2215_));
 sg13g2_nand2_1 _6250_ (.Y(_2216_),
    .A(net1895),
    .B(net1318));
 sg13g2_a21oi_1 _6251_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[13][1] ),
    .A2(net1284),
    .Y(_2217_),
    .B1(net1296));
 sg13g2_and2_1 _6252_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[15][1] ),
    .B(net1283),
    .X(_2218_));
 sg13g2_a21oi_1 _6253_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[14][1] ),
    .A2(net1318),
    .Y(_2219_),
    .B1(_2218_));
 sg13g2_a221oi_1 _6254_ (.B2(net1296),
    .C1(net1281),
    .B1(_2219_),
    .A1(_2216_),
    .Y(_2220_),
    .A2(_2217_));
 sg13g2_mux2_1 _6255_ (.A0(\scl_fifo1.scl_memory0.physical_memory0.memory[8][1] ),
    .A1(\scl_fifo1.scl_memory0.physical_memory0.memory[9][1] ),
    .S(net1282),
    .X(_2221_));
 sg13g2_and2_1 _6256_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[11][1] ),
    .B(net1282),
    .X(_2222_));
 sg13g2_a21oi_1 _6257_ (.A1(net949),
    .A2(net1317),
    .Y(_2223_),
    .B1(_2222_));
 sg13g2_a21oi_1 _6258_ (.A1(net1294),
    .A2(_2223_),
    .Y(_2224_),
    .B1(net1272));
 sg13g2_o21ai_1 _6259_ (.B1(_2224_),
    .Y(_2225_),
    .A1(net1294),
    .A2(_2221_));
 sg13g2_nor2_1 _6260_ (.A(net1274),
    .B(_2220_),
    .Y(_2226_));
 sg13g2_a21oi_1 _6261_ (.A1(_2225_),
    .A2(_2226_),
    .Y(_0009_),
    .B1(_2215_));
 sg13g2_mux2_1 _6262_ (.A0(\scl_fifo1.scl_memory0.physical_memory0.memory[0][2] ),
    .A1(\scl_fifo1.scl_memory0.physical_memory0.memory[1][2] ),
    .S(net1292),
    .X(_2227_));
 sg13g2_and2_1 _6263_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[3][2] ),
    .B(net1290),
    .X(_2228_));
 sg13g2_a21oi_1 _6264_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[2][2] ),
    .A2(net1322),
    .Y(_2229_),
    .B1(_2228_));
 sg13g2_a21oi_1 _6265_ (.A1(net1301),
    .A2(_2229_),
    .Y(_2230_),
    .B1(net1273));
 sg13g2_o21ai_1 _6266_ (.B1(_2230_),
    .Y(_2231_),
    .A1(net1301),
    .A2(_2227_));
 sg13g2_nand2_1 _6267_ (.Y(_2232_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[4][2] ),
    .B(net1323));
 sg13g2_a21oi_1 _6268_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[5][2] ),
    .A2(net1291),
    .Y(_2233_),
    .B1(net1302));
 sg13g2_and2_1 _6269_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[7][2] ),
    .B(net1291),
    .X(_2234_));
 sg13g2_a21oi_1 _6270_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[6][2] ),
    .A2(net1323),
    .Y(_2235_),
    .B1(_2234_));
 sg13g2_a221oi_1 _6271_ (.B2(net1301),
    .C1(net1280),
    .B1(_2235_),
    .A1(_2232_),
    .Y(_2236_),
    .A2(_2233_));
 sg13g2_nor2_1 _6272_ (.A(\scl_fifo1.n6238_o[3] ),
    .B(_2236_),
    .Y(_2237_));
 sg13g2_nand2_1 _6273_ (.Y(_2238_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[8][2] ),
    .B(net1319));
 sg13g2_a21oi_1 _6274_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[9][2] ),
    .A2(net1286),
    .Y(_2239_),
    .B1(net1298));
 sg13g2_and2_1 _6275_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[11][2] ),
    .B(net1284),
    .X(_2240_));
 sg13g2_a21oi_1 _6276_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[10][2] ),
    .A2(net1319),
    .Y(_2241_),
    .B1(_2240_));
 sg13g2_a221oi_1 _6277_ (.B2(net1298),
    .C1(net1272),
    .B1(_2241_),
    .A1(_2238_),
    .Y(_2242_),
    .A2(_2239_));
 sg13g2_mux2_1 _6278_ (.A0(\scl_fifo1.scl_memory0.physical_memory0.memory[12][2] ),
    .A1(\scl_fifo1.scl_memory0.physical_memory0.memory[13][2] ),
    .S(net1284),
    .X(_2243_));
 sg13g2_and2_1 _6279_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[15][2] ),
    .B(net1285),
    .X(_2244_));
 sg13g2_a21oi_1 _6280_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[14][2] ),
    .A2(net1320),
    .Y(_2245_),
    .B1(_2244_));
 sg13g2_a21oi_1 _6281_ (.A1(net1299),
    .A2(_2245_),
    .Y(_2246_),
    .B1(net1281));
 sg13g2_o21ai_1 _6282_ (.B1(_2246_),
    .Y(_2247_),
    .A1(net1298),
    .A2(_2243_));
 sg13g2_nor2_1 _6283_ (.A(net1274),
    .B(_2242_),
    .Y(_2248_));
 sg13g2_a22oi_1 _6284_ (.Y(_0010_),
    .B1(_2247_),
    .B2(_2248_),
    .A2(_2237_),
    .A1(_2231_));
 sg13g2_and2_1 _6285_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[3][3] ),
    .B(net1290),
    .X(_2249_));
 sg13g2_a21oi_1 _6286_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[2][3] ),
    .A2(net1324),
    .Y(_2250_),
    .B1(_2249_));
 sg13g2_nand2_1 _6287_ (.Y(_2251_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[0][3] ),
    .B(net1322));
 sg13g2_a21oi_1 _6288_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[1][3] ),
    .A2(net1290),
    .Y(_2252_),
    .B1(net1300));
 sg13g2_a221oi_1 _6289_ (.B2(_2252_),
    .C1(\scl_fifo1.n6238_o[2] ),
    .B1(_2251_),
    .A1(net1300),
    .Y(_2253_),
    .A2(_2250_));
 sg13g2_nand2_1 _6290_ (.Y(_2254_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[4][3] ),
    .B(net1323));
 sg13g2_a21oi_1 _6291_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[5][3] ),
    .A2(net1291),
    .Y(_2255_),
    .B1(net1302));
 sg13g2_and2_1 _6292_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[7][3] ),
    .B(net1291),
    .X(_2256_));
 sg13g2_a21oi_1 _6293_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[6][3] ),
    .A2(net1323),
    .Y(_2257_),
    .B1(_2256_));
 sg13g2_a221oi_1 _6294_ (.B2(net1302),
    .C1(net1280),
    .B1(_2257_),
    .A1(_2254_),
    .Y(_2258_),
    .A2(_2255_));
 sg13g2_nor3_2 _6295_ (.A(net1266),
    .B(_2253_),
    .C(_2258_),
    .Y(_2259_));
 sg13g2_nand2_1 _6296_ (.Y(_2260_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[12][3] ),
    .B(net1318));
 sg13g2_a21oi_1 _6297_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[13][3] ),
    .A2(net1283),
    .Y(_2261_),
    .B1(net1296));
 sg13g2_and2_1 _6298_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[15][3] ),
    .B(net1283),
    .X(_2262_));
 sg13g2_a21oi_1 _6299_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[14][3] ),
    .A2(net1318),
    .Y(_2263_),
    .B1(_2262_));
 sg13g2_a221oi_1 _6300_ (.B2(net1297),
    .C1(net1281),
    .B1(_2263_),
    .A1(_2260_),
    .Y(_2264_),
    .A2(_2261_));
 sg13g2_mux2_1 _6301_ (.A0(net682),
    .A1(\scl_fifo1.scl_memory0.physical_memory0.memory[9][3] ),
    .S(net1282),
    .X(_2265_));
 sg13g2_and2_1 _6302_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[11][3] ),
    .B(net1282),
    .X(_2266_));
 sg13g2_a21oi_1 _6303_ (.A1(net1017),
    .A2(net1317),
    .Y(_2267_),
    .B1(_2266_));
 sg13g2_a21oi_1 _6304_ (.A1(net1294),
    .A2(_2267_),
    .Y(_2268_),
    .B1(net1272));
 sg13g2_o21ai_1 _6305_ (.B1(_2268_),
    .Y(_2269_),
    .A1(net1294),
    .A2(_2265_));
 sg13g2_nor2_1 _6306_ (.A(net1274),
    .B(_2264_),
    .Y(_2270_));
 sg13g2_a21oi_1 _6307_ (.A1(_2269_),
    .A2(_2270_),
    .Y(_0011_),
    .B1(_2259_));
 sg13g2_mux2_1 _6308_ (.A0(\scl_fifo1.scl_memory0.physical_memory0.memory[0][4] ),
    .A1(\scl_fifo1.scl_memory0.physical_memory0.memory[1][4] ),
    .S(net1288),
    .X(_2271_));
 sg13g2_and2_1 _6309_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[3][4] ),
    .B(net1288),
    .X(_2272_));
 sg13g2_a21oi_1 _6310_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[2][4] ),
    .A2(net1321),
    .Y(_2273_),
    .B1(_2272_));
 sg13g2_a21oi_1 _6311_ (.A1(net1300),
    .A2(_2273_),
    .Y(_2274_),
    .B1(net1273));
 sg13g2_o21ai_1 _6312_ (.B1(_2274_),
    .Y(_2275_),
    .A1(net1300),
    .A2(_2271_));
 sg13g2_nand2_1 _6313_ (.Y(_2276_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[4][4] ),
    .B(net1321));
 sg13g2_a21oi_1 _6314_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[5][4] ),
    .A2(net1288),
    .Y(_2277_),
    .B1(net1303));
 sg13g2_and2_1 _6315_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[7][4] ),
    .B(net1289),
    .X(_2278_));
 sg13g2_a21oi_1 _6316_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[6][4] ),
    .A2(net1321),
    .Y(_2279_),
    .B1(_2278_));
 sg13g2_a221oi_1 _6317_ (.B2(net1303),
    .C1(net1280),
    .B1(_2279_),
    .A1(_2276_),
    .Y(_2280_),
    .A2(_2277_));
 sg13g2_nor2_1 _6318_ (.A(net1266),
    .B(_2280_),
    .Y(_2281_));
 sg13g2_nand2_1 _6319_ (.Y(_2282_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[12][4] ),
    .B(net1319));
 sg13g2_a21oi_1 _6320_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[13][4] ),
    .A2(net1284),
    .Y(_2283_),
    .B1(net1298));
 sg13g2_and2_1 _6321_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[15][4] ),
    .B(net1285),
    .X(_2284_));
 sg13g2_a21oi_1 _6322_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[14][4] ),
    .A2(net1319),
    .Y(_2285_),
    .B1(_2284_));
 sg13g2_a221oi_1 _6323_ (.B2(net1298),
    .C1(net1281),
    .B1(_2285_),
    .A1(_2282_),
    .Y(_2286_),
    .A2(_2283_));
 sg13g2_mux2_1 _6324_ (.A0(\scl_fifo1.scl_memory0.physical_memory0.memory[8][4] ),
    .A1(\scl_fifo1.scl_memory0.physical_memory0.memory[9][4] ),
    .S(net1286),
    .X(_2287_));
 sg13g2_and2_1 _6325_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[11][4] ),
    .B(net1282),
    .X(_2288_));
 sg13g2_a21oi_1 _6326_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[10][4] ),
    .A2(net1317),
    .Y(_2289_),
    .B1(_2288_));
 sg13g2_a21oi_1 _6327_ (.A1(net1295),
    .A2(_2289_),
    .Y(_2290_),
    .B1(net1272));
 sg13g2_o21ai_1 _6328_ (.B1(_2290_),
    .Y(_2291_),
    .A1(net1295),
    .A2(_2287_));
 sg13g2_nor2_1 _6329_ (.A(net1274),
    .B(_2286_),
    .Y(_2292_));
 sg13g2_a22oi_1 _6330_ (.Y(_0012_),
    .B1(_2291_),
    .B2(_2292_),
    .A2(_2281_),
    .A1(_2275_));
 sg13g2_and2_1 _6331_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[3][5] ),
    .B(net1290),
    .X(_2293_));
 sg13g2_a21oi_1 _6332_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[2][5] ),
    .A2(net1322),
    .Y(_2294_),
    .B1(_2293_));
 sg13g2_nand2_1 _6333_ (.Y(_2295_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[0][5] ),
    .B(net1322));
 sg13g2_a21oi_1 _6334_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[1][5] ),
    .A2(net1290),
    .Y(_2296_),
    .B1(net1301));
 sg13g2_a221oi_1 _6335_ (.B2(_2296_),
    .C1(\scl_fifo1.n6238_o[2] ),
    .B1(_2295_),
    .A1(net1301),
    .Y(_2297_),
    .A2(_2294_));
 sg13g2_nand2_1 _6336_ (.Y(_2298_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[4][5] ),
    .B(net1323));
 sg13g2_a21oi_1 _6337_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[5][5] ),
    .A2(net1291),
    .Y(_2299_),
    .B1(net1302));
 sg13g2_and2_1 _6338_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[7][5] ),
    .B(net1291),
    .X(_2300_));
 sg13g2_a21oi_1 _6339_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[6][5] ),
    .A2(net1323),
    .Y(_2301_),
    .B1(_2300_));
 sg13g2_a221oi_1 _6340_ (.B2(net1301),
    .C1(net1280),
    .B1(_2301_),
    .A1(_2298_),
    .Y(_2302_),
    .A2(_2299_));
 sg13g2_nor3_2 _6341_ (.A(net1266),
    .B(_2297_),
    .C(_2302_),
    .Y(_2303_));
 sg13g2_nand2_1 _6342_ (.Y(_2304_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[12][5] ),
    .B(net1318));
 sg13g2_a21oi_1 _6343_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[13][5] ),
    .A2(net1284),
    .Y(_2305_),
    .B1(net1297));
 sg13g2_and2_1 _6344_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[15][5] ),
    .B(net1283),
    .X(_2306_));
 sg13g2_a21oi_1 _6345_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[14][5] ),
    .A2(net1318),
    .Y(_2307_),
    .B1(_2306_));
 sg13g2_a221oi_1 _6346_ (.B2(net1296),
    .C1(net1281),
    .B1(_2307_),
    .A1(_2304_),
    .Y(_2308_),
    .A2(_2305_));
 sg13g2_mux2_1 _6347_ (.A0(\scl_fifo1.scl_memory0.physical_memory0.memory[8][5] ),
    .A1(\scl_fifo1.scl_memory0.physical_memory0.memory[9][5] ),
    .S(net1282),
    .X(_2309_));
 sg13g2_and2_1 _6348_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[11][5] ),
    .B(net1287),
    .X(_2310_));
 sg13g2_a21oi_1 _6349_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[10][5] ),
    .A2(net1317),
    .Y(_2311_),
    .B1(_2310_));
 sg13g2_a21oi_1 _6350_ (.A1(net1296),
    .A2(_2311_),
    .Y(_2312_),
    .B1(net1272));
 sg13g2_o21ai_1 _6351_ (.B1(_2312_),
    .Y(_2313_),
    .A1(net1296),
    .A2(_2309_));
 sg13g2_nor2_1 _6352_ (.A(net1274),
    .B(_2308_),
    .Y(_2314_));
 sg13g2_a21oi_2 _6353_ (.B1(_2303_),
    .Y(_0013_),
    .A2(_2314_),
    .A1(_2313_));
 sg13g2_and2_1 _6354_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[3][6] ),
    .B(net1290),
    .X(_2315_));
 sg13g2_a21oi_1 _6355_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[2][6] ),
    .A2(net1322),
    .Y(_2316_),
    .B1(_2315_));
 sg13g2_nand2_1 _6356_ (.Y(_2317_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[0][6] ),
    .B(net1322));
 sg13g2_a21oi_1 _6357_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[1][6] ),
    .A2(net1290),
    .Y(_2318_),
    .B1(net1304));
 sg13g2_a221oi_1 _6358_ (.B2(_2318_),
    .C1(net1273),
    .B1(_2317_),
    .A1(net1304),
    .Y(_2319_),
    .A2(_2316_));
 sg13g2_nand2_1 _6359_ (.Y(_2320_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[4][6] ),
    .B(net1323));
 sg13g2_a21oi_1 _6360_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[5][6] ),
    .A2(net1292),
    .Y(_2321_),
    .B1(net1302));
 sg13g2_and2_1 _6361_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[7][6] ),
    .B(net1291),
    .X(_2322_));
 sg13g2_a21oi_1 _6362_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[6][6] ),
    .A2(net1323),
    .Y(_2323_),
    .B1(_2322_));
 sg13g2_a221oi_1 _6363_ (.B2(net1302),
    .C1(net1280),
    .B1(_2323_),
    .A1(_2320_),
    .Y(_2324_),
    .A2(_2321_));
 sg13g2_nor3_2 _6364_ (.A(net1266),
    .B(_2319_),
    .C(_2324_),
    .Y(_2325_));
 sg13g2_nand2_1 _6365_ (.Y(_2326_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[12][6] ),
    .B(net1318));
 sg13g2_a21oi_1 _6366_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[13][6] ),
    .A2(net1284),
    .Y(_2327_),
    .B1(net1297));
 sg13g2_and2_1 _6367_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[15][6] ),
    .B(net1287),
    .X(_2328_));
 sg13g2_a21oi_1 _6368_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[14][6] ),
    .A2(net1318),
    .Y(_2329_),
    .B1(_2328_));
 sg13g2_a221oi_1 _6369_ (.B2(net1297),
    .C1(net1281),
    .B1(_2329_),
    .A1(_2326_),
    .Y(_2330_),
    .A2(_2327_));
 sg13g2_and2_1 _6370_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[11][6] ),
    .B(net1282),
    .X(_2331_));
 sg13g2_a21oi_1 _6371_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[10][6] ),
    .A2(net1317),
    .Y(_2332_),
    .B1(_2331_));
 sg13g2_nand2_1 _6372_ (.Y(_2333_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[8][6] ),
    .B(net1317));
 sg13g2_a21oi_1 _6373_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[9][6] ),
    .A2(net1283),
    .Y(_2334_),
    .B1(net1294));
 sg13g2_a221oi_1 _6374_ (.B2(_2334_),
    .C1(net1272),
    .B1(_2333_),
    .A1(net1295),
    .Y(_2335_),
    .A2(_2332_));
 sg13g2_nor3_1 _6375_ (.A(net1274),
    .B(_2330_),
    .C(_2335_),
    .Y(_2336_));
 sg13g2_nor2_1 _6376_ (.A(_2325_),
    .B(_2336_),
    .Y(_0014_));
 sg13g2_mux2_1 _6377_ (.A0(\scl_fifo1.scl_memory0.physical_memory0.memory[4][7] ),
    .A1(\scl_fifo1.scl_memory0.physical_memory0.memory[5][7] ),
    .S(net1288),
    .X(_2337_));
 sg13g2_and2_1 _6378_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[7][7] ),
    .B(net1289),
    .X(_2338_));
 sg13g2_a21oi_1 _6379_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[6][7] ),
    .A2(net1321),
    .Y(_2339_),
    .B1(_2338_));
 sg13g2_a21oi_1 _6380_ (.A1(net1303),
    .A2(_2339_),
    .Y(_2340_),
    .B1(net1280));
 sg13g2_o21ai_1 _6381_ (.B1(_2340_),
    .Y(_2341_),
    .A1(net1303),
    .A2(_2337_));
 sg13g2_nand2_1 _6382_ (.Y(_2342_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[0][7] ),
    .B(net1321));
 sg13g2_a21oi_1 _6383_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[1][7] ),
    .A2(net1289),
    .Y(_2343_),
    .B1(net1303));
 sg13g2_and2_1 _6384_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[3][7] ),
    .B(net1288),
    .X(_2344_));
 sg13g2_a21oi_1 _6385_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[2][7] ),
    .A2(net1321),
    .Y(_2345_),
    .B1(_2344_));
 sg13g2_a221oi_1 _6386_ (.B2(net1303),
    .C1(net1273),
    .B1(_2345_),
    .A1(_2342_),
    .Y(_2346_),
    .A2(_2343_));
 sg13g2_nor2_1 _6387_ (.A(net1266),
    .B(_2346_),
    .Y(_2347_));
 sg13g2_nand2_1 _6388_ (.Y(_2348_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[12][7] ),
    .B(net1319));
 sg13g2_a21oi_1 _6389_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[13][7] ),
    .A2(net1284),
    .Y(_2349_),
    .B1(net1298));
 sg13g2_and2_1 _6390_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[15][7] ),
    .B(net1284),
    .X(_2350_));
 sg13g2_a21oi_1 _6391_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[14][7] ),
    .A2(net1320),
    .Y(_2351_),
    .B1(_2350_));
 sg13g2_a221oi_1 _6392_ (.B2(net1299),
    .C1(net1281),
    .B1(_2351_),
    .A1(_2348_),
    .Y(_2352_),
    .A2(_2349_));
 sg13g2_and2_1 _6393_ (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[11][7] ),
    .B(net1287),
    .X(_2353_));
 sg13g2_a21oi_1 _6394_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[10][7] ),
    .A2(net1317),
    .Y(_2354_),
    .B1(_2353_));
 sg13g2_nand2_1 _6395_ (.Y(_2355_),
    .A(\scl_fifo1.scl_memory0.physical_memory0.memory[8][7] ),
    .B(net1319));
 sg13g2_a21oi_1 _6396_ (.A1(\scl_fifo1.scl_memory0.physical_memory0.memory[9][7] ),
    .A2(net1286),
    .Y(_2356_),
    .B1(net1296));
 sg13g2_a221oi_1 _6397_ (.B2(_2356_),
    .C1(net1272),
    .B1(_2355_),
    .A1(net1296),
    .Y(_2357_),
    .A2(_2354_));
 sg13g2_nor3_1 _6398_ (.A(_1055_),
    .B(_2352_),
    .C(_2357_),
    .Y(_2358_));
 sg13g2_a21oi_2 _6399_ (.B1(_2358_),
    .Y(_0015_),
    .A2(_2347_),
    .A1(_2341_));
 sg13g2_nand2_1 _6400_ (.Y(_2359_),
    .A(_1703_),
    .B(_1710_));
 sg13g2_nor2_2 _6401_ (.A(_1665_),
    .B(net1312),
    .Y(_2360_));
 sg13g2_nand2_1 _6402_ (.Y(_2361_),
    .A(net1316),
    .B(net1314));
 sg13g2_nor2_1 _6403_ (.A(net1330),
    .B(_1665_),
    .Y(_2362_));
 sg13g2_nand2_2 _6404_ (.Y(_2363_),
    .A(_1653_),
    .B(net1316));
 sg13g2_nand2_2 _6405_ (.Y(_2364_),
    .A(net1315),
    .B(_2362_));
 sg13g2_nand2_1 _6406_ (.Y(_2365_),
    .A(net1329),
    .B(net1314));
 sg13g2_nand2_2 _6407_ (.Y(_2366_),
    .A(_1665_),
    .B(net1314));
 sg13g2_nor2_2 _6408_ (.A(_1653_),
    .B(net1316),
    .Y(_2367_));
 sg13g2_nand2_2 _6409_ (.Y(_2368_),
    .A(net1330),
    .B(_1665_));
 sg13g2_nand2_2 _6410_ (.Y(_2369_),
    .A(net1315),
    .B(_2367_));
 sg13g2_nand2_1 _6411_ (.Y(_2370_),
    .A(_2364_),
    .B(_2369_));
 sg13g2_nand2_1 _6412_ (.Y(_2371_),
    .A(net1308),
    .B(_2370_));
 sg13g2_nand2_2 _6413_ (.Y(_2372_),
    .A(net1329),
    .B(net1305));
 sg13g2_nand2b_1 _6414_ (.Y(_2373_),
    .B(_2366_),
    .A_N(_2372_));
 sg13g2_nand2_1 _6415_ (.Y(_2374_),
    .A(_2371_),
    .B(_2373_));
 sg13g2_nand2_1 _6416_ (.Y(_2375_),
    .A(net1329),
    .B(net1312));
 sg13g2_nor2_1 _6417_ (.A(net1305),
    .B(_2375_),
    .Y(_2376_));
 sg13g2_nand2_2 _6418_ (.Y(_2377_),
    .A(_1666_),
    .B(_2376_));
 sg13g2_nor2_2 _6419_ (.A(net1276),
    .B(_2377_),
    .Y(_2378_));
 sg13g2_nand2_1 _6420_ (.Y(_2379_),
    .A(_2363_),
    .B(_2366_));
 sg13g2_nor2_2 _6421_ (.A(net1307),
    .B(net1278),
    .Y(_2380_));
 sg13g2_nand2_1 _6422_ (.Y(_2381_),
    .A(net1309),
    .B(net1275));
 sg13g2_nand2_1 _6423_ (.Y(_2382_),
    .A(net1316),
    .B(net1312));
 sg13g2_inv_1 _6424_ (.Y(_2383_),
    .A(_2382_));
 sg13g2_nand4_1 _6425_ (.B(_2366_),
    .C(_2380_),
    .A(_2363_),
    .Y(_2384_),
    .D(_2382_));
 sg13g2_nor2_2 _6426_ (.A(net1308),
    .B(net1278),
    .Y(_2385_));
 sg13g2_o21ai_1 _6427_ (.B1(_2384_),
    .Y(_2386_),
    .A1(net1276),
    .A2(_2377_));
 sg13g2_a221oi_1 _6428_ (.B2(_2385_),
    .C1(_2386_),
    .B1(_2379_),
    .A1(net1279),
    .Y(_2387_),
    .A2(_2374_));
 sg13g2_nor2_1 _6429_ (.A(net1314),
    .B(_2372_),
    .Y(_2388_));
 sg13g2_nor2_1 _6430_ (.A(net1276),
    .B(_2388_),
    .Y(_2389_));
 sg13g2_nor2_1 _6431_ (.A(net1316),
    .B(net1314),
    .Y(_2390_));
 sg13g2_nand2_2 _6432_ (.Y(_2391_),
    .A(_1665_),
    .B(net1312));
 sg13g2_nand4_1 _6433_ (.B(_2363_),
    .C(_2368_),
    .A(net1308),
    .Y(_2392_),
    .D(_2391_));
 sg13g2_a21oi_1 _6434_ (.A1(net1329),
    .A2(_2366_),
    .Y(_2393_),
    .B1(net1279));
 sg13g2_a22oi_1 _6435_ (.Y(_2394_),
    .B1(_2393_),
    .B2(_2372_),
    .A2(_2392_),
    .A1(_2389_));
 sg13g2_nand2b_1 _6436_ (.Y(_2395_),
    .B(_1702_),
    .A_N(_2394_));
 sg13g2_nand2_1 _6437_ (.Y(_2396_),
    .A(net1311),
    .B(_2363_));
 sg13g2_nor2_1 _6438_ (.A(_2367_),
    .B(_2396_),
    .Y(_2397_));
 sg13g2_inv_1 _6439_ (.Y(_2398_),
    .A(_2397_));
 sg13g2_o21ai_1 _6440_ (.B1(net1306),
    .Y(_2399_),
    .A1(_2370_),
    .A2(_2397_));
 sg13g2_nor2_1 _6441_ (.A(net1279),
    .B(_1702_),
    .Y(_2400_));
 sg13g2_nand2_1 _6442_ (.Y(_2401_),
    .A(_1665_),
    .B(net1310));
 sg13g2_nand2_1 _6443_ (.Y(_2402_),
    .A(net1309),
    .B(_2367_));
 sg13g2_nand3_1 _6444_ (.B(_2400_),
    .C(_2402_),
    .A(_2399_),
    .Y(_2403_));
 sg13g2_nand2_1 _6445_ (.Y(_2404_),
    .A(net1316),
    .B(net1305));
 sg13g2_nor2_1 _6446_ (.A(net1309),
    .B(_2364_),
    .Y(_2405_));
 sg13g2_nand2_2 _6447_ (.Y(_2406_),
    .A(_1653_),
    .B(net1312));
 sg13g2_nor2_2 _6448_ (.A(net1329),
    .B(net1316),
    .Y(_2407_));
 sg13g2_nand2_1 _6449_ (.Y(_2408_),
    .A(net1312),
    .B(_2407_));
 sg13g2_nand2_2 _6450_ (.Y(_2409_),
    .A(_1665_),
    .B(net1305));
 sg13g2_nor3_1 _6451_ (.A(net1315),
    .B(net1305),
    .C(_2407_),
    .Y(_2410_));
 sg13g2_nor4_1 _6452_ (.A(net1275),
    .B(net1268),
    .C(_2405_),
    .D(_2410_),
    .Y(_2411_));
 sg13g2_o21ai_1 _6453_ (.B1(_2411_),
    .Y(_2412_),
    .A1(_2406_),
    .A2(_2409_));
 sg13g2_nand4_1 _6454_ (.B(_2395_),
    .C(_2403_),
    .A(net1267),
    .Y(_2413_),
    .D(_2412_));
 sg13g2_nor2_2 _6455_ (.A(_1703_),
    .B(net1267),
    .Y(_2414_));
 sg13g2_nand4_1 _6456_ (.B(_2371_),
    .C(_2375_),
    .A(net1276),
    .Y(_2415_),
    .D(_2404_));
 sg13g2_o21ai_1 _6457_ (.B1(_2369_),
    .Y(_2416_),
    .A1(net1314),
    .A2(_2363_));
 sg13g2_nand2_2 _6458_ (.Y(_2417_),
    .A(net1306),
    .B(net1279));
 sg13g2_nand2b_1 _6459_ (.Y(_2418_),
    .B(_2416_),
    .A_N(_2417_));
 sg13g2_nand2_2 _6460_ (.Y(_2419_),
    .A(net1308),
    .B(net1279));
 sg13g2_nand4_1 _6461_ (.B(net1278),
    .C(_2364_),
    .A(net1308),
    .Y(_2420_),
    .D(_2391_));
 sg13g2_nand3_1 _6462_ (.B(_2418_),
    .C(_2420_),
    .A(_2415_),
    .Y(_2421_));
 sg13g2_o21ai_1 _6463_ (.B1(_2413_),
    .Y(_2422_),
    .A1(_2359_),
    .A2(_2387_));
 sg13g2_a21oi_1 _6464_ (.A1(_2414_),
    .A2(_2421_),
    .Y(_2423_),
    .B1(_2422_));
 sg13g2_nor2_1 _6465_ (.A(net1276),
    .B(_2376_),
    .Y(_2424_));
 sg13g2_o21ai_1 _6466_ (.B1(_2424_),
    .Y(_2425_),
    .A1(_2372_),
    .A2(_2383_));
 sg13g2_nand2_2 _6467_ (.Y(_2426_),
    .A(net1329),
    .B(_2391_));
 sg13g2_o21ai_1 _6468_ (.B1(net1276),
    .Y(_2427_),
    .A1(net1305),
    .A2(_2426_));
 sg13g2_nand3_1 _6469_ (.B(_2425_),
    .C(_2427_),
    .A(net1263),
    .Y(_2428_));
 sg13g2_o21ai_1 _6470_ (.B1(_2428_),
    .Y(_0016_),
    .A1(net1263),
    .A2(_2423_));
 sg13g2_nand2_1 _6471_ (.Y(_2429_),
    .A(net1316),
    .B(_2388_));
 sg13g2_nor2_1 _6472_ (.A(_2365_),
    .B(_2417_),
    .Y(_2430_));
 sg13g2_nor2_1 _6473_ (.A(_1719_),
    .B(_2430_),
    .Y(_2431_));
 sg13g2_nand3_1 _6474_ (.B(net1309),
    .C(_2367_),
    .A(net1313),
    .Y(_2432_));
 sg13g2_a21oi_1 _6475_ (.A1(net1308),
    .A2(_2360_),
    .Y(_2433_),
    .B1(_2388_));
 sg13g2_a21oi_1 _6476_ (.A1(_2432_),
    .A2(_2433_),
    .Y(_2434_),
    .B1(net1275));
 sg13g2_nand2_1 _6477_ (.Y(_2435_),
    .A(_2368_),
    .B(_2396_));
 sg13g2_xnor2_1 _6478_ (.Y(_2436_),
    .A(_2409_),
    .B(_2435_));
 sg13g2_a21oi_1 _6479_ (.A1(net1275),
    .A2(_2436_),
    .Y(_2437_),
    .B1(_2434_));
 sg13g2_o21ai_1 _6480_ (.B1(net1267),
    .Y(_2438_),
    .A1(_2381_),
    .A2(_2408_));
 sg13g2_nand3_1 _6481_ (.B(_2406_),
    .C(_2426_),
    .A(_2385_),
    .Y(_2439_));
 sg13g2_o21ai_1 _6482_ (.B1(_2439_),
    .Y(_2440_),
    .A1(_2382_),
    .A2(_2417_));
 sg13g2_a21oi_1 _6483_ (.A1(_1710_),
    .A2(_2437_),
    .Y(_2441_),
    .B1(net1268));
 sg13g2_o21ai_1 _6484_ (.B1(_2441_),
    .Y(_2442_),
    .A1(_2438_),
    .A2(_2440_));
 sg13g2_nand2_1 _6485_ (.Y(_2443_),
    .A(_2363_),
    .B(_2369_));
 sg13g2_a21oi_1 _6486_ (.A1(_0097_),
    .A2(net1314),
    .Y(_2444_),
    .B1(net1277));
 sg13g2_nor2_1 _6487_ (.A(_2368_),
    .B(_2417_),
    .Y(_2445_));
 sg13g2_a21o_1 _6488_ (.A2(_2444_),
    .A1(_2407_),
    .B1(_2445_),
    .X(_2446_));
 sg13g2_a221oi_1 _6489_ (.B2(_2385_),
    .C1(_2446_),
    .B1(_2443_),
    .A1(_2380_),
    .Y(_2447_),
    .A2(_2397_));
 sg13g2_nor2b_1 _6490_ (.A(_2447_),
    .B_N(_2414_),
    .Y(_2448_));
 sg13g2_o21ai_1 _6491_ (.B1(net1278),
    .Y(_2449_),
    .A1(net1306),
    .A2(_2369_));
 sg13g2_a21oi_1 _6492_ (.A1(net1306),
    .A2(_2362_),
    .Y(_2450_),
    .B1(_2449_));
 sg13g2_and3_1 _6493_ (.X(_2451_),
    .A(net1275),
    .B(_2391_),
    .C(_2409_));
 sg13g2_nor4_1 _6494_ (.A(_1703_),
    .B(_1710_),
    .C(_2450_),
    .D(_2451_),
    .Y(_2452_));
 sg13g2_nor3_1 _6495_ (.A(net1264),
    .B(_2448_),
    .C(_2452_),
    .Y(_2453_));
 sg13g2_a22oi_1 _6496_ (.Y(_0017_),
    .B1(_2442_),
    .B2(_2453_),
    .A2(_2431_),
    .A1(_2429_));
 sg13g2_nor2_1 _6497_ (.A(net1311),
    .B(net1279),
    .Y(_2454_));
 sg13g2_a21oi_1 _6498_ (.A1(_2401_),
    .A2(_2454_),
    .Y(_2455_),
    .B1(_2378_));
 sg13g2_nor2_1 _6499_ (.A(_2364_),
    .B(_2381_),
    .Y(_2456_));
 sg13g2_nand2_2 _6500_ (.Y(_2457_),
    .A(_0097_),
    .B(_2360_));
 sg13g2_a21oi_1 _6501_ (.A1(_2366_),
    .A2(_2398_),
    .Y(_2458_),
    .B1(_2419_));
 sg13g2_o21ai_1 _6502_ (.B1(_1703_),
    .Y(_2459_),
    .A1(net1275),
    .A2(_2457_));
 sg13g2_nor3_1 _6503_ (.A(_2456_),
    .B(_2458_),
    .C(_2459_),
    .Y(_2460_));
 sg13g2_a21oi_1 _6504_ (.A1(net1268),
    .A2(_2455_),
    .Y(_2461_),
    .B1(_2460_));
 sg13g2_nand2_1 _6505_ (.Y(_2462_),
    .A(net1315),
    .B(_2445_));
 sg13g2_nand4_1 _6506_ (.B(net1278),
    .C(_2361_),
    .A(net1310),
    .Y(_2463_),
    .D(_2396_));
 sg13g2_o21ai_1 _6507_ (.B1(_2385_),
    .Y(_2464_),
    .A1(_2370_),
    .A2(_2390_));
 sg13g2_nand4_1 _6508_ (.B(net1278),
    .C(_2401_),
    .A(net1330),
    .Y(_2465_),
    .D(_2457_));
 sg13g2_nand4_1 _6509_ (.B(net1329),
    .C(net1277),
    .A(_0097_),
    .Y(_2466_),
    .D(_2360_));
 sg13g2_nand4_1 _6510_ (.B(_2462_),
    .C(_2463_),
    .A(net1268),
    .Y(_2467_),
    .D(_2464_));
 sg13g2_nand3_1 _6511_ (.B(_2465_),
    .C(_2466_),
    .A(_1703_),
    .Y(_2468_));
 sg13g2_a22oi_1 _6512_ (.Y(_2469_),
    .B1(_2467_),
    .B2(_2468_),
    .A2(_2416_),
    .A1(_2380_));
 sg13g2_nor2_1 _6513_ (.A(net1267),
    .B(_2469_),
    .Y(_2470_));
 sg13g2_a21oi_1 _6514_ (.A1(net1267),
    .A2(_2461_),
    .Y(_2471_),
    .B1(_2470_));
 sg13g2_nand3_1 _6515_ (.B(net1310),
    .C(_2361_),
    .A(net1330),
    .Y(_2472_));
 sg13g2_a21oi_1 _6516_ (.A1(_2373_),
    .A2(_2472_),
    .Y(_2473_),
    .B1(net1278));
 sg13g2_nand4_1 _6517_ (.B(net1311),
    .C(net1279),
    .A(net1329),
    .Y(_2474_),
    .D(_2409_));
 sg13g2_nor2_1 _6518_ (.A(_1719_),
    .B(_2473_),
    .Y(_2475_));
 sg13g2_a22oi_1 _6519_ (.Y(_0018_),
    .B1(_2474_),
    .B2(_2475_),
    .A2(_2471_),
    .A1(_1719_));
 sg13g2_nand3_1 _6520_ (.B(_2369_),
    .C(_2429_),
    .A(net1276),
    .Y(_2476_));
 sg13g2_nand2_1 _6521_ (.Y(_2477_),
    .A(net1263),
    .B(_2476_));
 sg13g2_a221oi_1 _6522_ (.B2(net1314),
    .C1(_2378_),
    .B1(_2445_),
    .A1(_2366_),
    .Y(_2478_),
    .A2(_2380_));
 sg13g2_o21ai_1 _6523_ (.B1(_2432_),
    .Y(_2479_),
    .A1(_2406_),
    .A2(_2409_));
 sg13g2_a21oi_1 _6524_ (.A1(_2400_),
    .A2(_2479_),
    .Y(_2480_),
    .B1(_1710_));
 sg13g2_o21ai_1 _6525_ (.B1(_2480_),
    .Y(_2481_),
    .A1(_1703_),
    .A2(_2478_));
 sg13g2_nand2b_1 _6526_ (.Y(_2482_),
    .B(_2429_),
    .A_N(_2449_));
 sg13g2_a21oi_1 _6527_ (.A1(_2369_),
    .A2(_2408_),
    .Y(_2483_),
    .B1(net1308));
 sg13g2_o21ai_1 _6528_ (.B1(net1275),
    .Y(_2484_),
    .A1(net1305),
    .A2(_2365_));
 sg13g2_o21ai_1 _6529_ (.B1(_2482_),
    .Y(_2485_),
    .A1(_2483_),
    .A2(_2484_));
 sg13g2_nand2b_1 _6530_ (.Y(_2486_),
    .B(_2485_),
    .A_N(_2359_));
 sg13g2_a22oi_1 _6531_ (.Y(_2487_),
    .B1(_2407_),
    .B2(_2454_),
    .A2(_2367_),
    .A1(net1311));
 sg13g2_o21ai_1 _6532_ (.B1(_2414_),
    .Y(_2488_),
    .A1(_2385_),
    .A2(_2487_));
 sg13g2_nand4_1 _6533_ (.B(_2481_),
    .C(_2486_),
    .A(_1719_),
    .Y(_2489_),
    .D(_2488_));
 sg13g2_o21ai_1 _6534_ (.B1(_2489_),
    .Y(_0019_),
    .A1(_2389_),
    .A2(_2477_));
 sg13g2_nand4_1 _6535_ (.B(_1703_),
    .C(_2380_),
    .A(net1311),
    .Y(_2490_),
    .D(_2407_));
 sg13g2_and2_1 _6536_ (.A(net1278),
    .B(_2372_),
    .X(_2491_));
 sg13g2_nand4_1 _6537_ (.B(net1311),
    .C(_2401_),
    .A(_0099_),
    .Y(_2492_),
    .D(_2491_));
 sg13g2_a21oi_1 _6538_ (.A1(_2490_),
    .A2(_2492_),
    .Y(_2493_),
    .B1(_1710_));
 sg13g2_nand4_1 _6539_ (.B(_1710_),
    .C(_2366_),
    .A(net1330),
    .Y(_2494_),
    .D(_2380_));
 sg13g2_a21oi_1 _6540_ (.A1(_2462_),
    .A2(_2494_),
    .Y(_2495_),
    .B1(net1268));
 sg13g2_nor3_1 _6541_ (.A(net1264),
    .B(_2493_),
    .C(_2495_),
    .Y(_2496_));
 sg13g2_nor2b_1 _6542_ (.A(_2378_),
    .B_N(_2466_),
    .Y(_2497_));
 sg13g2_a21oi_1 _6543_ (.A1(_2431_),
    .A2(_2497_),
    .Y(_0020_),
    .B1(_2496_));
 sg13g2_nor2_1 _6544_ (.A(_2360_),
    .B(_2372_),
    .Y(_2498_));
 sg13g2_o21ai_1 _6545_ (.B1(_2424_),
    .Y(_2499_),
    .A1(net1308),
    .A2(_2426_));
 sg13g2_o21ai_1 _6546_ (.B1(_2499_),
    .Y(_2500_),
    .A1(_2427_),
    .A2(_2498_));
 sg13g2_nand2_1 _6547_ (.Y(_2501_),
    .A(_2472_),
    .B(_2491_));
 sg13g2_a21oi_1 _6548_ (.A1(_2484_),
    .A2(_2501_),
    .Y(_2502_),
    .B1(_1711_));
 sg13g2_a21oi_1 _6549_ (.A1(_2369_),
    .A2(_2408_),
    .Y(_2503_),
    .B1(_2419_));
 sg13g2_nor3_1 _6550_ (.A(_1653_),
    .B(net1275),
    .C(_2457_),
    .Y(_2504_));
 sg13g2_nor3_1 _6551_ (.A(_2438_),
    .B(_2503_),
    .C(_2504_),
    .Y(_2505_));
 sg13g2_nor3_1 _6552_ (.A(net1268),
    .B(_2502_),
    .C(_2505_),
    .Y(_2506_));
 sg13g2_nand4_1 _6553_ (.B(_2367_),
    .C(_2385_),
    .A(net1312),
    .Y(_2507_),
    .D(_2414_));
 sg13g2_nor2_1 _6554_ (.A(net1263),
    .B(_2506_),
    .Y(_2508_));
 sg13g2_a22oi_1 _6555_ (.Y(_0021_),
    .B1(_2507_),
    .B2(_2508_),
    .A2(_2500_),
    .A1(net1263));
 sg13g2_o21ai_1 _6556_ (.B1(_2491_),
    .Y(_2509_),
    .A1(net1305),
    .A2(_2426_));
 sg13g2_nand3_1 _6557_ (.B(_2365_),
    .C(_2368_),
    .A(net1277),
    .Y(_2510_));
 sg13g2_nor2_1 _6558_ (.A(_2359_),
    .B(_2385_),
    .Y(_2511_));
 sg13g2_nand3_1 _6559_ (.B(_2510_),
    .C(_2511_),
    .A(_2509_),
    .Y(_2512_));
 sg13g2_and3_1 _6560_ (.X(_2513_),
    .A(_1711_),
    .B(_2400_),
    .C(_2405_));
 sg13g2_nand3_1 _6561_ (.B(net1267),
    .C(_2362_),
    .A(net1311),
    .Y(_2514_));
 sg13g2_nor3_1 _6562_ (.A(_1703_),
    .B(_2419_),
    .C(_2514_),
    .Y(_2515_));
 sg13g2_o21ai_1 _6563_ (.B1(net1330),
    .Y(_2516_),
    .A1(net1311),
    .A2(_2419_));
 sg13g2_nor3_1 _6564_ (.A(net1263),
    .B(_2513_),
    .C(_2515_),
    .Y(_2517_));
 sg13g2_a22oi_1 _6565_ (.Y(_0022_),
    .B1(_2517_),
    .B2(_2512_),
    .A2(_2516_),
    .A1(net1263));
 sg13g2_nor2_1 _6566_ (.A(net785),
    .B(_1516_),
    .Y(_2518_));
 sg13g2_a21oi_1 _6567_ (.A1(net785),
    .A2(_1516_),
    .Y(_2519_),
    .B1(_1355_));
 sg13g2_nor2b_1 _6568_ (.A(_2518_),
    .B_N(net786),
    .Y(\usbfunction0.scl_usbgpiophy0.scl_extendwidth0.scl_counter0.n7961_o[0] ));
 sg13g2_nor2_1 _6569_ (.A(net1142),
    .B(_2518_),
    .Y(_2520_));
 sg13g2_and2_1 _6570_ (.A(net1142),
    .B(_2518_),
    .X(_2521_));
 sg13g2_nor3_1 _6571_ (.A(_1355_),
    .B(_2520_),
    .C(_2521_),
    .Y(\usbfunction0.scl_usbgpiophy0.scl_extendwidth0.scl_counter0.n7961_o[1] ));
 sg13g2_o21ai_1 _6572_ (.B1(s_m_status_rxactive),
    .Y(_2522_),
    .A1(net608),
    .A2(_2521_));
 sg13g2_a21oi_1 _6573_ (.A1(net608),
    .A2(_2521_),
    .Y(\usbfunction0.scl_usbgpiophy0.scl_extendwidth0.scl_counter0.n7961_o[2] ),
    .B1(_2522_));
 sg13g2_nor2_1 _6574_ (.A(_0043_),
    .B(_1034_),
    .Y(_2523_));
 sg13g2_or2_2 _6575_ (.X(_2524_),
    .B(_1034_),
    .A(_0043_));
 sg13g2_nor2_1 _6576_ (.A(net543),
    .B(_2524_),
    .Y(_2525_));
 sg13g2_o21ai_1 _6577_ (.B1(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.in_in_valid ),
    .Y(_2526_),
    .A1(net543),
    .A2(_2524_));
 sg13g2_a21oi_1 _6578_ (.A1(net543),
    .A2(_2524_),
    .Y(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.scl_counter0.n8088_o[0] ),
    .B1(_2526_));
 sg13g2_nand2_1 _6579_ (.Y(_2527_),
    .A(net1488),
    .B(_2525_));
 sg13g2_o21ai_1 _6580_ (.B1(net835),
    .Y(_2528_),
    .A1(net1488),
    .A2(_2525_));
 sg13g2_nor2b_1 _6581_ (.A(net836),
    .B_N(_2527_),
    .Y(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.scl_counter0.n8088_o[1] ));
 sg13g2_o21ai_1 _6582_ (.B1(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.in_in_valid ),
    .Y(_2529_),
    .A1(net554),
    .A2(_2527_));
 sg13g2_a21oi_1 _6583_ (.A1(net554),
    .A2(_2527_),
    .Y(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.scl_counter0.n8088_o[2] ),
    .B1(_2529_));
 sg13g2_a21o_2 _6584_ (.A2(_0780_),
    .A1(_0043_),
    .B1(_1034_),
    .X(_2530_));
 sg13g2_nor2_1 _6585_ (.A(net1682),
    .B(_2530_),
    .Y(_2531_));
 sg13g2_a21oi_1 _6586_ (.A1(net1682),
    .A2(_2530_),
    .Y(_2532_),
    .B1(_2171_));
 sg13g2_nor2b_1 _6587_ (.A(_2531_),
    .B_N(_2532_),
    .Y(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.scl_counter0.n8128_o[0] ));
 sg13g2_nor2b_1 _6588_ (.A(_2531_),
    .B_N(net1581),
    .Y(_2533_));
 sg13g2_nor3_2 _6589_ (.A(net1682),
    .B(net1581),
    .C(_2530_),
    .Y(_2534_));
 sg13g2_nor3_1 _6590_ (.A(_2171_),
    .B(net1582),
    .C(_2534_),
    .Y(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.scl_counter0.n8128_o[1] ));
 sg13g2_nand2_1 _6591_ (.Y(_2535_),
    .A(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.s_m_value[2] ),
    .B(_2534_));
 sg13g2_a21oi_1 _6592_ (.A1(net1727),
    .A2(_2534_),
    .Y(_2536_),
    .B1(_2171_));
 sg13g2_o21ai_1 _6593_ (.B1(_2536_),
    .Y(_2537_),
    .A1(net1727),
    .A2(_2534_));
 sg13g2_inv_1 _6594_ (.Y(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.scl_counter0.n8128_o[2] ),
    .A(_2537_));
 sg13g2_xor2_1 _6595_ (.B(_2535_),
    .A(net1719),
    .X(_2538_));
 sg13g2_nor2_1 _6596_ (.A(_2171_),
    .B(net1720),
    .Y(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.scl_counter0.n8128_o[3] ));
 sg13g2_and2_1 _6597_ (.A(_0782_),
    .B(_2181_),
    .X(_2539_));
 sg13g2_and3_1 _6598_ (.X(_2540_),
    .A(net1015),
    .B(_0782_),
    .C(_2180_));
 sg13g2_nor2_1 _6599_ (.A(net1015),
    .B(_0782_),
    .Y(_2541_));
 sg13g2_nor3_1 _6600_ (.A(_2539_),
    .B(_2540_),
    .C(_2541_),
    .Y(\usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8195_o[0] ));
 sg13g2_xnor2_1 _6601_ (.Y(_2542_),
    .A(net1637),
    .B(_2540_));
 sg13g2_nor2_1 _6602_ (.A(_2539_),
    .B(_2542_),
    .Y(\usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8195_o[1] ));
 sg13g2_a21oi_1 _6603_ (.A1(\usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8209_q[1] ),
    .A2(_2540_),
    .Y(_2543_),
    .B1(net588));
 sg13g2_nand2_1 _6604_ (.Y(_2544_),
    .A(_0778_),
    .B(_2180_));
 sg13g2_a21oi_1 _6605_ (.A1(_0782_),
    .A2(_2544_),
    .Y(\usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8195_o[2] ),
    .B1(net589));
 sg13g2_nor2_1 _6606_ (.A(net562),
    .B(net1436),
    .Y(\usbfunction0.scl_usbgpiophy0.scl_pulseextender0.scl_counter0.n8221_o[0] ));
 sg13g2_nand2_1 _6607_ (.Y(_2545_),
    .A(net562),
    .B(\usbfunction0.scl_usbgpiophy0.scl_pulseextender0.scl_counter0.n8243_q[1] ));
 sg13g2_xnor2_1 _6608_ (.Y(_2546_),
    .A(net562),
    .B(net1035));
 sg13g2_nor2_1 _6609_ (.A(net1436),
    .B(_2546_),
    .Y(\usbfunction0.scl_usbgpiophy0.scl_pulseextender0.scl_counter0.n8221_o[1] ));
 sg13g2_nand4_1 _6610_ (.B(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.s_m_value[0] ),
    .C(net1727),
    .A(net1757),
    .Y(_2547_),
    .D(net1719));
 sg13g2_nor2b_1 _6611_ (.A(net1713),
    .B_N(_1033_),
    .Y(_2548_));
 sg13g2_a21oi_2 _6612_ (.B1(_1036_),
    .Y(_2549_),
    .A2(_2548_),
    .A1(_0749_));
 sg13g2_nand2b_1 _6613_ (.Y(_2550_),
    .B(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7508_o ),
    .A_N(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7654_q[1] ));
 sg13g2_nand3_1 _6614_ (.B(_2549_),
    .C(_2550_),
    .A(_2172_),
    .Y(_2551_));
 sg13g2_o21ai_1 _6615_ (.B1(_2551_),
    .Y(_2552_),
    .A1(_0780_),
    .A2(_2547_));
 sg13g2_nand2b_1 _6616_ (.Y(_2553_),
    .B(_2552_),
    .A_N(_2530_));
 sg13g2_inv_1 _6617_ (.Y(_2554_),
    .A(_2553_));
 sg13g2_nor3_1 _6618_ (.A(net546),
    .B(\usbfunction0.scl_usbgpiophy0.scl_pulseextender1.scl_counter0.n8282_q[1] ),
    .C(_2554_),
    .Y(\usbfunction0.scl_usbgpiophy0.scl_pulseextender1.scl_counter0.n8260_o[0] ));
 sg13g2_nor3_1 _6619_ (.A(_0776_),
    .B(net558),
    .C(_2554_),
    .Y(\usbfunction0.scl_usbgpiophy0.scl_pulseextender1.scl_counter0.n8260_o[1] ));
 sg13g2_and3_1 _6620_ (.X(\usbfunction0.s_m_rx_eop ),
    .A(net1096),
    .B(\usbfunction0.scl_usbgpiophy0.n6650_q ),
    .C(_1355_));
 sg13g2_xor2_1 _6621_ (.B(_1870_),
    .A(net1168),
    .X(_2555_));
 sg13g2_xor2_1 _6622_ (.B(_1880_),
    .A(\scl_fifo0.n2737_o[0] ),
    .X(_2556_));
 sg13g2_xor2_1 _6623_ (.B(\scl_fifo0.n2722_o[1] ),
    .A(_0118_),
    .X(_2557_));
 sg13g2_xor2_1 _6624_ (.B(\scl_fifo0.n2722_o[2] ),
    .A(_0127_),
    .X(_2558_));
 sg13g2_nand3_1 _6625_ (.B(_2557_),
    .C(_2558_),
    .A(_2556_),
    .Y(_2559_));
 sg13g2_xor2_1 _6626_ (.B(\scl_fifo0.n2722_o[4] ),
    .A(net1026),
    .X(_2560_));
 sg13g2_nor3_1 _6627_ (.A(_2555_),
    .B(_2559_),
    .C(_2560_),
    .Y(\scl_fifo0.n2746_o ));
 sg13g2_nor2b_1 _6628_ (.A(_1216_),
    .B_N(net564),
    .Y(\scl_streamarbiter_2.n6171_o ));
 sg13g2_xnor2_1 _6629_ (.Y(_2561_),
    .A(\scl_fifo1.n6278_o[0] ),
    .B(\scl_fifo1.n6233_o[0] ));
 sg13g2_xor2_1 _6630_ (.B(\scl_fifo1.n6233_o[1] ),
    .A(\scl_fifo1.n6278_o[1] ),
    .X(_2562_));
 sg13g2_nand2b_1 _6631_ (.Y(_2563_),
    .B(\scl_fifo1.n6233_o[2] ),
    .A_N(\scl_fifo1.n6278_o[2] ));
 sg13g2_nand2b_1 _6632_ (.Y(_2564_),
    .B(\scl_fifo1.n6278_o[2] ),
    .A_N(\scl_fifo1.n6233_o[2] ));
 sg13g2_xnor2_1 _6633_ (.Y(_2565_),
    .A(net1769),
    .B(\scl_fifo1.n6233_o[4] ));
 sg13g2_xor2_1 _6634_ (.B(\scl_fifo1.n6233_o[3] ),
    .A(\scl_fifo1.n6278_o[3] ),
    .X(_2566_));
 sg13g2_nand3_1 _6635_ (.B(_2563_),
    .C(_2564_),
    .A(_2561_),
    .Y(_2567_));
 sg13g2_nor4_2 _6636_ (.A(_2562_),
    .B(_2565_),
    .C(_2566_),
    .Y(\scl_fifo1.n6287_o ),
    .D(_2567_));
 sg13g2_nand3b_1 _6637_ (.B(_1006_),
    .C(_1847_),
    .Y(_2568_),
    .A_N(_0040_));
 sg13g2_a21oi_1 _6638_ (.A1(net548),
    .A2(_2568_),
    .Y(\usbfunction0.rxstream0.n6755_o ),
    .B1(_1844_));
 sg13g2_nor2b_1 _6639_ (.A(net749),
    .B_N(net570),
    .Y(_2569_));
 sg13g2_and2_1 _6640_ (.A(net1097),
    .B(_2569_),
    .X(\usbfunction0.s_m_rx_error ));
 sg13g2_a21oi_1 _6641_ (.A1(net1437),
    .A2(net1386),
    .Y(\usbfunction0.scl_usbgpiophy0.n6529_o ),
    .B1(_1355_));
 sg13g2_a21oi_1 _6642_ (.A1(net530),
    .A2(net538),
    .Y(\usbfunction0.scl_usbgpiophy0.n6533_o ),
    .B1(_1355_));
 sg13g2_nor2_2 _6643_ (.A(net1096),
    .B(net538),
    .Y(_2570_));
 sg13g2_nand2b_1 _6644_ (.Y(_2571_),
    .B(net540),
    .A_N(net536));
 sg13g2_a21oi_1 _6645_ (.A1(_2570_),
    .A2(_2571_),
    .Y(_2572_),
    .B1(net570));
 sg13g2_nor2_1 _6646_ (.A(\usbfunction0.s_m_rx_eop ),
    .B(net571),
    .Y(\usbfunction0.scl_usbgpiophy0.n6553_o ));
 sg13g2_nor2_1 _6647_ (.A(_1036_),
    .B(_2524_),
    .Y(_2573_));
 sg13g2_nor2_1 _6648_ (.A(_2548_),
    .B(_2573_),
    .Y(\usbfunction0.scl_usbgpiophy0.scl_addeopdeferred0.scl_eraselastbeat0.n8008_o ));
 sg13g2_nor2_1 _6649_ (.A(_1033_),
    .B(_2573_),
    .Y(\usbfunction0.scl_usbgpiophy0.scl_addeopdeferred0.n7339_o ));
 sg13g2_a21o_1 _6650_ (.A2(_2524_),
    .A1(net1020),
    .B1(_1519_),
    .X(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7634_o ));
 sg13g2_a21o_1 _6651_ (.A2(_2545_),
    .A1(net1006),
    .B1(net1436),
    .X(\usbfunction0.scl_usbgpiophy0.scl_pulseextender0.n7741_o ));
 sg13g2_nand2b_1 _6652_ (.Y(\usbfunction0.scl_usbgpiophy0.s_ret_3 ),
    .B(_2553_),
    .A_N(net627));
 sg13g2_nand3_1 _6653_ (.B(net558),
    .C(_2553_),
    .A(_0776_),
    .Y(_2574_));
 sg13g2_and2_1 _6654_ (.A(\usbfunction0.scl_usbgpiophy0.s_ret_3 ),
    .B(_2574_),
    .X(\usbfunction0.scl_usbgpiophy0.scl_pulseextender1.n7766_o ));
 sg13g2_a21oi_1 _6655_ (.A1(_1005_),
    .A2(_1409_),
    .Y(_2575_),
    .B1(net1420));
 sg13g2_inv_1 _6656_ (.Y(_2576_),
    .A(_2575_));
 sg13g2_o21ai_1 _6657_ (.B1(_2576_),
    .Y(_2577_),
    .A1(net1694),
    .A2(_1361_));
 sg13g2_a21oi_1 _6658_ (.A1(_0684_),
    .A2(_1361_),
    .Y(_0187_),
    .B1(_2577_));
 sg13g2_o21ai_1 _6659_ (.B1(_2576_),
    .Y(_2578_),
    .A1(net1654),
    .A2(_1361_));
 sg13g2_a21oi_1 _6660_ (.A1(_0683_),
    .A2(_1361_),
    .Y(_0188_),
    .B1(_2578_));
 sg13g2_o21ai_1 _6661_ (.B1(_2576_),
    .Y(_2579_),
    .A1(net1613),
    .A2(_1361_));
 sg13g2_a21oi_1 _6662_ (.A1(_0682_),
    .A2(_1361_),
    .Y(_0189_),
    .B1(_2579_));
 sg13g2_o21ai_1 _6663_ (.B1(_2576_),
    .Y(_2580_),
    .A1(net1561),
    .A2(_1361_));
 sg13g2_a21oi_1 _6664_ (.A1(\usbfunction0.n2313_o[3] ),
    .A2(_1361_),
    .Y(_0190_),
    .B1(_2580_));
 sg13g2_nand2_1 _6665_ (.Y(_2581_),
    .A(net622),
    .B(_1362_));
 sg13g2_o21ai_1 _6666_ (.B1(_2581_),
    .Y(_0191_),
    .A1(_1012_),
    .A2(_1017_));
 sg13g2_a21o_1 _6667_ (.A2(net1426),
    .A1(net912),
    .B1(_1363_),
    .X(_0192_));
 sg13g2_a21oi_1 _6668_ (.A1(_1192_),
    .A2(net1271),
    .Y(_2582_),
    .B1(net1673));
 sg13g2_a21oi_1 _6669_ (.A1(net1673),
    .A2(net1270),
    .Y(_0193_),
    .B1(net1674));
 sg13g2_xnor2_1 _6670_ (.Y(_2583_),
    .A(\scl_bitbangengine0.s_m_value_2[0] ),
    .B(_0133_));
 sg13g2_nand3_1 _6671_ (.B(net1270),
    .C(_2583_),
    .A(_1192_),
    .Y(_2584_));
 sg13g2_o21ai_1 _6672_ (.B1(_2584_),
    .Y(_0194_),
    .A1(_0771_),
    .A2(net1270));
 sg13g2_nand3_1 _6673_ (.B(net1116),
    .C(net1270),
    .A(net1673),
    .Y(_2585_));
 sg13g2_nand2b_1 _6674_ (.Y(_2586_),
    .B(_2585_),
    .A_N(net1785));
 sg13g2_nand4_1 _6675_ (.B(net1116),
    .C(net1785),
    .A(net1673),
    .Y(_2587_),
    .D(net1270));
 sg13g2_and3_1 _6676_ (.X(_0195_),
    .A(net1265),
    .B(_2586_),
    .C(_2587_));
 sg13g2_nor2_1 _6677_ (.A(net745),
    .B(net1349),
    .Y(_2588_));
 sg13g2_a21oi_1 _6678_ (.A1(net1454),
    .A2(net1349),
    .Y(_0196_),
    .B1(_2588_));
 sg13g2_nor2_1 _6679_ (.A(net642),
    .B(net1348),
    .Y(_2589_));
 sg13g2_a21oi_1 _6680_ (.A1(net1457),
    .A2(net1348),
    .Y(_0197_),
    .B1(_2589_));
 sg13g2_mux2_1 _6681_ (.A0(net737),
    .A1(net1474),
    .S(net1348),
    .X(_0198_));
 sg13g2_nor2_1 _6682_ (.A(net810),
    .B(net1348),
    .Y(_2590_));
 sg13g2_a21oi_1 _6683_ (.A1(net1460),
    .A2(net1348),
    .Y(_0199_),
    .B1(_2590_));
 sg13g2_mux2_1 _6684_ (.A0(net697),
    .A1(net1473),
    .S(net1348),
    .X(_0200_));
 sg13g2_mux2_1 _6685_ (.A0(net702),
    .A1(net1470),
    .S(net1348),
    .X(_0201_));
 sg13g2_mux2_1 _6686_ (.A0(net1011),
    .A1(net1467),
    .S(net1349),
    .X(_0202_));
 sg13g2_mux2_1 _6687_ (.A0(net675),
    .A1(net1464),
    .S(net1348),
    .X(_0203_));
 sg13g2_nor2_1 _6688_ (.A(_1193_),
    .B(_1328_),
    .Y(_2591_));
 sg13g2_nor2_1 _6689_ (.A(_1328_),
    .B(_1952_),
    .Y(_2592_));
 sg13g2_nor3_1 _6690_ (.A(_0084_),
    .B(_1328_),
    .C(_1952_),
    .Y(_2593_));
 sg13g2_nor2_1 _6691_ (.A(_1077_),
    .B(net1412),
    .Y(_2594_));
 sg13g2_o21ai_1 _6692_ (.B1(_2594_),
    .Y(_2595_),
    .A1(_1193_),
    .A2(_1196_));
 sg13g2_nor2_1 _6693_ (.A(_1077_),
    .B(net1413),
    .Y(_2596_));
 sg13g2_o21ai_1 _6694_ (.B1(net1374),
    .Y(_2597_),
    .A1(_1193_),
    .A2(_1196_));
 sg13g2_or2_2 _6695_ (.X(_2598_),
    .B(net1359),
    .A(net1412));
 sg13g2_nor3_2 _6696_ (.A(\scl_bitbangengine0.n5920_q[0] ),
    .B(\scl_bitbangengine0.n5920_q[1] ),
    .C(\scl_bitbangengine0.n5920_q[2] ),
    .Y(_2599_));
 sg13g2_nor2b_2 _6697_ (.A(\scl_bitbangengine0.n5920_q[3] ),
    .B_N(_2599_),
    .Y(_2600_));
 sg13g2_xor2_1 _6698_ (.B(_2599_),
    .A(net1778),
    .X(_2601_));
 sg13g2_nand2_2 _6699_ (.Y(_2602_),
    .A(net1502),
    .B(\scl_bitbangengine0.n5919_q ));
 sg13g2_nor2_1 _6700_ (.A(_0083_),
    .B(_2602_),
    .Y(_2603_));
 sg13g2_nor3_2 _6701_ (.A(net1451),
    .B(_0083_),
    .C(_2602_),
    .Y(_2604_));
 sg13g2_and2_1 _6702_ (.A(net1497),
    .B(_2604_),
    .X(_2605_));
 sg13g2_xor2_1 _6703_ (.B(_2604_),
    .A(net1497),
    .X(_2606_));
 sg13g2_xnor2_1 _6704_ (.Y(_2607_),
    .A(net1497),
    .B(_2604_));
 sg13g2_a22oi_1 _6705_ (.Y(_2608_),
    .B1(_2606_),
    .B2(net1413),
    .A2(_2601_),
    .A1(net1374));
 sg13g2_xor2_1 _6706_ (.B(\scl_bitbangengine0.n5919_q ),
    .A(net1502),
    .X(_2609_));
 sg13g2_nand2b_1 _6707_ (.Y(_2610_),
    .B(net1411),
    .A_N(_2609_));
 sg13g2_o21ai_1 _6708_ (.B1(_2610_),
    .Y(_2611_),
    .A1(net1778),
    .A2(_2598_));
 sg13g2_a21oi_1 _6709_ (.A1(net1359),
    .A2(_2608_),
    .Y(_0204_),
    .B1(_2611_));
 sg13g2_xnor2_1 _6710_ (.Y(_2612_),
    .A(_0736_),
    .B(_2600_));
 sg13g2_and2_1 _6711_ (.A(net1494),
    .B(_2605_),
    .X(_2613_));
 sg13g2_xor2_1 _6712_ (.B(_2605_),
    .A(net1494),
    .X(_2614_));
 sg13g2_a22oi_1 _6713_ (.Y(_2615_),
    .B1(_2614_),
    .B2(net1413),
    .A2(_2612_),
    .A1(net1374));
 sg13g2_nor2_1 _6714_ (.A(net1411),
    .B(_2615_),
    .Y(_2616_));
 sg13g2_xnor2_1 _6715_ (.Y(_2617_),
    .A(net1501),
    .B(_2602_));
 sg13g2_a22oi_1 _6716_ (.Y(_2618_),
    .B1(_2617_),
    .B2(net1411),
    .A2(_2616_),
    .A1(net1359));
 sg13g2_o21ai_1 _6717_ (.B1(_2618_),
    .Y(_0205_),
    .A1(_0736_),
    .A2(_2598_));
 sg13g2_and3_1 _6718_ (.X(_2619_),
    .A(_0736_),
    .B(_0737_),
    .C(_2600_));
 sg13g2_a21oi_1 _6719_ (.A1(_0736_),
    .A2(_2600_),
    .Y(_2620_),
    .B1(_0737_));
 sg13g2_or2_1 _6720_ (.X(_2621_),
    .B(_2620_),
    .A(_2619_));
 sg13g2_and2_1 _6721_ (.A(\scl_bitbangengine0.n3267_o ),
    .B(_2613_),
    .X(_2622_));
 sg13g2_xnor2_1 _6722_ (.Y(_2623_),
    .A(_0692_),
    .B(_2613_));
 sg13g2_a22oi_1 _6723_ (.Y(_2624_),
    .B1(_2623_),
    .B2(net1413),
    .A2(_2621_),
    .A1(net1374));
 sg13g2_xnor2_1 _6724_ (.Y(_2625_),
    .A(net1451),
    .B(_2603_));
 sg13g2_nand2b_1 _6725_ (.Y(_2626_),
    .B(net1411),
    .A_N(_2625_));
 sg13g2_o21ai_1 _6726_ (.B1(_2626_),
    .Y(_2627_),
    .A1(net1716),
    .A2(_2598_));
 sg13g2_a21oi_1 _6727_ (.A1(net1359),
    .A2(_2624_),
    .Y(_0206_),
    .B1(_2627_));
 sg13g2_nor2_1 _6728_ (.A(net1037),
    .B(_2598_),
    .Y(_2628_));
 sg13g2_nand2_2 _6729_ (.Y(_2629_),
    .A(\scl_bitbangengine0.n3258_o ),
    .B(_2622_));
 sg13g2_xnor2_1 _6730_ (.Y(_2630_),
    .A(_0694_),
    .B(_2622_));
 sg13g2_nand2_1 _6731_ (.Y(_2631_),
    .A(_0145_),
    .B(_2619_));
 sg13g2_xnor2_1 _6732_ (.Y(_2632_),
    .A(_0145_),
    .B(_2619_));
 sg13g2_a221oi_1 _6733_ (.B2(net1374),
    .C1(net1411),
    .B1(_2632_),
    .A1(net1413),
    .Y(_2633_),
    .A2(_2630_));
 sg13g2_a221oi_1 _6734_ (.B2(net1359),
    .C1(_2628_),
    .B1(_2633_),
    .A1(net1411),
    .Y(_0207_),
    .A2(_2607_));
 sg13g2_nor2_2 _6735_ (.A(_0732_),
    .B(_2629_),
    .Y(_2634_));
 sg13g2_xnor2_1 _6736_ (.Y(_2635_),
    .A(net1492),
    .B(_2629_));
 sg13g2_xnor2_1 _6737_ (.Y(_2636_),
    .A(_0732_),
    .B(_2629_));
 sg13g2_xnor2_1 _6738_ (.Y(_2637_),
    .A(net1786),
    .B(_2631_));
 sg13g2_a22oi_1 _6739_ (.Y(_2638_),
    .B1(_2637_),
    .B2(net1374),
    .A2(_2635_),
    .A1(net1413));
 sg13g2_nand2b_1 _6740_ (.Y(_2639_),
    .B(net1411),
    .A_N(_2614_));
 sg13g2_o21ai_1 _6741_ (.B1(_2639_),
    .Y(_2640_),
    .A1(net1786),
    .A2(_2598_));
 sg13g2_a21oi_1 _6742_ (.A1(net1359),
    .A2(_2638_),
    .Y(_0208_),
    .B1(_2640_));
 sg13g2_nand2_2 _6743_ (.Y(_2641_),
    .A(_1183_),
    .B(_2600_));
 sg13g2_xnor2_1 _6744_ (.Y(_2642_),
    .A(\scl_bitbangengine0.n5920_q[8] ),
    .B(_2641_));
 sg13g2_a221oi_1 _6745_ (.B2(net1374),
    .C1(net1412),
    .B1(_2642_),
    .A1(_2591_),
    .Y(_2643_),
    .A2(_2634_));
 sg13g2_nand2b_1 _6746_ (.Y(_2644_),
    .B(net1411),
    .A_N(_2623_));
 sg13g2_o21ai_1 _6747_ (.B1(_2644_),
    .Y(_2645_),
    .A1(net1867),
    .A2(_2598_));
 sg13g2_a21oi_1 _6748_ (.A1(net1360),
    .A2(_2643_),
    .Y(_0209_),
    .B1(_2645_));
 sg13g2_nor2_1 _6749_ (.A(_1079_),
    .B(_1087_),
    .Y(_2646_));
 sg13g2_o21ai_1 _6750_ (.B1(_1327_),
    .Y(_2647_),
    .A1(_1193_),
    .A2(_1328_));
 sg13g2_nand4_1 _6751_ (.B(\scl_bitbangengine0.n5898_q[2] ),
    .C(_1075_),
    .A(\scl_bitbangengine0.n5898_q[3] ),
    .Y(_2648_),
    .D(_1180_));
 sg13g2_nor2_1 _6752_ (.A(_2592_),
    .B(_2647_),
    .Y(_2649_));
 sg13g2_nand3_1 _6753_ (.B(_2648_),
    .C(_2649_),
    .A(_1205_),
    .Y(_2650_));
 sg13g2_nor3_1 _6754_ (.A(net1406),
    .B(_2646_),
    .C(_2650_),
    .Y(_2651_));
 sg13g2_nor2b_1 _6755_ (.A(_1092_),
    .B_N(_2651_),
    .Y(_2652_));
 sg13g2_nand3_1 _6756_ (.B(_1086_),
    .C(_1098_),
    .A(net1500),
    .Y(_2653_));
 sg13g2_nor2_1 _6757_ (.A(_1079_),
    .B(_1083_),
    .Y(_2654_));
 sg13g2_nor2_1 _6758_ (.A(net1492),
    .B(_1078_),
    .Y(_2655_));
 sg13g2_nor2_2 _6759_ (.A(\scl_bitbangengine0.n5898_q[1] ),
    .B(_1328_),
    .Y(_2656_));
 sg13g2_nor4_1 _6760_ (.A(_1201_),
    .B(_2654_),
    .C(net1373),
    .D(_2656_),
    .Y(_2657_));
 sg13g2_and3_1 _6761_ (.X(_2658_),
    .A(_2652_),
    .B(_2653_),
    .C(_2657_));
 sg13g2_and2_1 _6762_ (.A(net683),
    .B(_1100_),
    .X(_2659_));
 sg13g2_nor3_2 _6763_ (.A(net1451),
    .B(_1085_),
    .C(_1097_),
    .Y(_2660_));
 sg13g2_nand2_1 _6764_ (.Y(_2661_),
    .A(net1495),
    .B(_1096_));
 sg13g2_nor3_1 _6765_ (.A(net1501),
    .B(net1498),
    .C(_2661_),
    .Y(_2662_));
 sg13g2_nor3_1 _6766_ (.A(net1501),
    .B(net1498),
    .C(_2661_),
    .Y(_2663_));
 sg13g2_nor3_1 _6767_ (.A(_2659_),
    .B(_2660_),
    .C(_2663_),
    .Y(_2664_));
 sg13g2_nand3_1 _6768_ (.B(_2658_),
    .C(_2664_),
    .A(_1955_),
    .Y(_2665_));
 sg13g2_nor2_1 _6769_ (.A(_1210_),
    .B(_2665_),
    .Y(_2666_));
 sg13g2_nand2_1 _6770_ (.Y(_2667_),
    .A(net1503),
    .B(_2656_));
 sg13g2_nor2_1 _6771_ (.A(net1866),
    .B(_2667_),
    .Y(_2668_));
 sg13g2_nand2b_1 _6772_ (.Y(_2669_),
    .B(net1373),
    .A_N(_0083_));
 sg13g2_a22oi_1 _6773_ (.Y(_2670_),
    .B1(_2664_),
    .B2(_2669_),
    .A2(_2660_),
    .A1(net1502));
 sg13g2_nor2b_1 _6774_ (.A(_2670_),
    .B_N(_2651_),
    .Y(_2671_));
 sg13g2_nor2b_1 _6775_ (.A(_0084_),
    .B_N(_2647_),
    .Y(_2672_));
 sg13g2_o21ai_1 _6776_ (.B1(_1954_),
    .Y(_2673_),
    .A1(_2671_),
    .A2(_2672_));
 sg13g2_a21oi_1 _6777_ (.A1(_1189_),
    .A2(_1197_),
    .Y(_2674_),
    .B1(_2673_));
 sg13g2_o21ai_1 _6778_ (.B1(_0141_),
    .Y(_2675_),
    .A1(_1193_),
    .A2(_1196_));
 sg13g2_o21ai_1 _6779_ (.B1(_2674_),
    .Y(_2676_),
    .A1(_1211_),
    .A2(_2675_));
 sg13g2_nor3_1 _6780_ (.A(_2666_),
    .B(_2668_),
    .C(_2676_),
    .Y(_2677_));
 sg13g2_a21o_1 _6781_ (.A2(_2666_),
    .A1(net1503),
    .B1(_2677_),
    .X(_0210_));
 sg13g2_nor3_1 _6782_ (.A(net1898),
    .B(_1210_),
    .C(_2665_),
    .Y(_2678_));
 sg13g2_nor3_2 _6783_ (.A(net1497),
    .B(_1079_),
    .C(_1083_),
    .Y(_2679_));
 sg13g2_or2_1 _6784_ (.X(_2680_),
    .B(_2679_),
    .A(_2662_));
 sg13g2_nand2b_1 _6785_ (.Y(_2681_),
    .B(_2652_),
    .A_N(_2656_));
 sg13g2_nor4_1 _6786_ (.A(_1197_),
    .B(_2678_),
    .C(_2680_),
    .D(_2681_),
    .Y(_0211_));
 sg13g2_nand4_1 _6787_ (.B(_2648_),
    .C(_2649_),
    .A(_1200_),
    .Y(_2682_),
    .D(_2667_));
 sg13g2_nor4_1 _6788_ (.A(_1092_),
    .B(net1406),
    .C(_2679_),
    .D(_2682_),
    .Y(_2683_));
 sg13g2_nand3b_1 _6789_ (.B(_2683_),
    .C(_1955_),
    .Y(_2684_),
    .A_N(_2659_));
 sg13g2_nor2_1 _6790_ (.A(net1751),
    .B(_2665_),
    .Y(_2685_));
 sg13g2_nor2_1 _6791_ (.A(_2684_),
    .B(_2685_),
    .Y(_0212_));
 sg13g2_a21o_1 _6792_ (.A2(_2647_),
    .A1(\scl_bitbangengine0.n3817_o ),
    .B1(_2592_),
    .X(_2686_));
 sg13g2_nor3_1 _6793_ (.A(_1212_),
    .B(_2680_),
    .C(_2686_),
    .Y(_2687_));
 sg13g2_a21oi_1 _6794_ (.A1(_1189_),
    .A2(_1197_),
    .Y(_2688_),
    .B1(_2687_));
 sg13g2_nand2_1 _6795_ (.Y(_2689_),
    .A(_1954_),
    .B(_2667_));
 sg13g2_nor2_1 _6796_ (.A(_2688_),
    .B(_2689_),
    .Y(_2690_));
 sg13g2_nor3_1 _6797_ (.A(_2666_),
    .B(_2668_),
    .C(_2690_),
    .Y(_2691_));
 sg13g2_a21o_1 _6798_ (.A2(_2666_),
    .A1(net1800),
    .B1(_2691_),
    .X(_0213_));
 sg13g2_nor2_1 _6799_ (.A(_1335_),
    .B(_1337_),
    .Y(_2692_));
 sg13g2_nor2_1 _6800_ (.A(net752),
    .B(_2692_),
    .Y(_2693_));
 sg13g2_a21oi_1 _6801_ (.A1(net752),
    .A2(_1336_),
    .Y(_0214_),
    .B1(_2693_));
 sg13g2_nand2_1 _6802_ (.Y(_2694_),
    .A(net566),
    .B(_1337_));
 sg13g2_nor3_1 _6803_ (.A(_0120_),
    .B(_0131_),
    .C(_1337_),
    .Y(_2695_));
 sg13g2_nand2_1 _6804_ (.Y(_2696_),
    .A(_0120_),
    .B(_0131_));
 sg13g2_nand2_1 _6805_ (.Y(_2697_),
    .A(_2692_),
    .B(_2696_));
 sg13g2_o21ai_1 _6806_ (.B1(net567),
    .Y(_0215_),
    .A1(_2695_),
    .A2(_2697_));
 sg13g2_o21ai_1 _6807_ (.B1(_2692_),
    .Y(_2698_),
    .A1(_0770_),
    .A2(_2695_));
 sg13g2_a21o_1 _6808_ (.A2(_2695_),
    .A1(_0770_),
    .B1(_2698_),
    .X(_2699_));
 sg13g2_o21ai_1 _6809_ (.B1(_2699_),
    .Y(_0216_),
    .A1(_0768_),
    .A2(_1336_));
 sg13g2_a22oi_1 _6810_ (.Y(_2700_),
    .B1(net1373),
    .B2(net1861),
    .A2(_1078_),
    .A1(\scl_bitbangengine0.n5905_q ));
 sg13g2_inv_1 _6811_ (.Y(_0217_),
    .A(net1862));
 sg13g2_nor2_2 _6812_ (.A(\scl_uartrx0.s_m_value[2] ),
    .B(_0734_),
    .Y(_2701_));
 sg13g2_nor2_1 _6813_ (.A(net1461),
    .B(\scl_uartrx0.s_m_value[0] ),
    .Y(_2702_));
 sg13g2_nor2b_2 _6814_ (.A(_0081_),
    .B_N(\scl_uartrx0.s_m_value[2] ),
    .Y(_2703_));
 sg13g2_nand2_1 _6815_ (.Y(_2704_),
    .A(\scl_uartrx0.s_m_value[2] ),
    .B(_0734_));
 sg13g2_nand2_1 _6816_ (.Y(_2705_),
    .A(_2702_),
    .B(_2703_));
 sg13g2_nor2_1 _6817_ (.A(\scl_uartrx0.s_m_value[1] ),
    .B(_0082_),
    .Y(_2706_));
 sg13g2_a21oi_1 _6818_ (.A1(net1461),
    .A2(_0734_),
    .Y(_2707_),
    .B1(_2706_));
 sg13g2_nand2_1 _6819_ (.Y(_2708_),
    .A(_2705_),
    .B(_2707_));
 sg13g2_a21oi_1 _6820_ (.A1(_0928_),
    .A2(_2701_),
    .Y(_2709_),
    .B1(_2708_));
 sg13g2_and2_1 _6821_ (.A(_2701_),
    .B(_2702_),
    .X(_2710_));
 sg13g2_nand3b_1 _6822_ (.B(_2709_),
    .C(_0926_),
    .Y(_2711_),
    .A_N(_2710_));
 sg13g2_nand2b_1 _6823_ (.Y(_2712_),
    .B(net1461),
    .A_N(\scl_uartrx0.s_m_value[0] ));
 sg13g2_nor3_1 _6824_ (.A(\scl_uartrx0.s_m_value[2] ),
    .B(_0734_),
    .C(_2712_),
    .Y(_2713_));
 sg13g2_nand2_1 _6825_ (.Y(_2714_),
    .A(net1504),
    .B(_2713_));
 sg13g2_nand2_1 _6826_ (.Y(_2715_),
    .A(net788),
    .B(_2711_));
 sg13g2_o21ai_1 _6827_ (.B1(_2715_),
    .Y(_0218_),
    .A1(_2711_),
    .A2(_2714_));
 sg13g2_nor2b_1 _6828_ (.A(net1461),
    .B_N(\scl_uartrx0.s_m_value[0] ),
    .Y(_2716_));
 sg13g2_nand2b_1 _6829_ (.Y(_2717_),
    .B(\scl_uartrx0.s_m_value[0] ),
    .A_N(net1461));
 sg13g2_nor2_2 _6830_ (.A(_0927_),
    .B(_2701_),
    .Y(_2718_));
 sg13g2_o21ai_1 _6831_ (.B1(_2718_),
    .Y(_2719_),
    .A1(_2704_),
    .A2(_2716_));
 sg13g2_nand2_1 _6832_ (.Y(_2720_),
    .A(net1504),
    .B(_2703_));
 sg13g2_nand2_1 _6833_ (.Y(_2721_),
    .A(net868),
    .B(_2719_));
 sg13g2_nand2_1 _6834_ (.Y(_2722_),
    .A(_2716_),
    .B(_2718_));
 sg13g2_o21ai_1 _6835_ (.B1(_2721_),
    .Y(_0219_),
    .A1(_2720_),
    .A2(_2722_));
 sg13g2_o21ai_1 _6836_ (.B1(_1084_),
    .Y(_2723_),
    .A1(net1866),
    .A2(_1077_));
 sg13g2_nand2b_1 _6837_ (.Y(_0220_),
    .B(_2723_),
    .A_N(_2660_));
 sg13g2_nor3_2 _6838_ (.A(\scl_fifo1.n6229_o[2] ),
    .B(\scl_fifo1.n6229_o[3] ),
    .C(_1991_),
    .Y(_2724_));
 sg13g2_mux2_1 _6839_ (.A0(net9),
    .A1(net1),
    .S(net1499),
    .X(_2725_));
 sg13g2_nand2_1 _6840_ (.Y(_2726_),
    .A(net1502),
    .B(net1406));
 sg13g2_a22oi_1 _6841_ (.Y(_2727_),
    .B1(_2725_),
    .B2(_1101_),
    .A2(_1178_),
    .A1(net9));
 sg13g2_nand3_1 _6842_ (.B(_2726_),
    .C(_2727_),
    .A(net1269),
    .Y(_2728_));
 sg13g2_a22oi_1 _6843_ (.Y(_2729_),
    .B1(_1936_),
    .B2(_2728_),
    .A2(net1416),
    .A1(net674));
 sg13g2_nor2_1 _6844_ (.A(net654),
    .B(net1187),
    .Y(_2730_));
 sg13g2_a21oi_1 _6845_ (.A1(net1187),
    .A2(net1255),
    .Y(_0221_),
    .B1(_2730_));
 sg13g2_mux2_1 _6846_ (.A0(net10),
    .A1(net2),
    .S(net1499),
    .X(_2731_));
 sg13g2_a22oi_1 _6847_ (.Y(_2732_),
    .B1(_2731_),
    .B2(_1101_),
    .A2(_1178_),
    .A1(net10));
 sg13g2_a22oi_1 _6848_ (.Y(_2733_),
    .B1(_1095_),
    .B2(_2732_),
    .A2(net1405),
    .A1(_0730_));
 sg13g2_or2_1 _6849_ (.X(_2734_),
    .B(_2733_),
    .A(net1271));
 sg13g2_a22oi_1 _6850_ (.Y(_2735_),
    .B1(_1938_),
    .B2(_2734_),
    .A2(net1416),
    .A1(\s_out_3[1] ));
 sg13g2_nor2_1 _6851_ (.A(net956),
    .B(net1188),
    .Y(_2736_));
 sg13g2_a21oi_1 _6852_ (.A1(net1188),
    .A2(net1254),
    .Y(_0222_),
    .B1(_2736_));
 sg13g2_and2_1 _6853_ (.A(\s_out_3[2] ),
    .B(net1417),
    .X(_2737_));
 sg13g2_nand2_1 _6854_ (.Y(_2738_),
    .A(net1504),
    .B(_1166_));
 sg13g2_nand2_1 _6855_ (.Y(_2739_),
    .A(net1499),
    .B(net3));
 sg13g2_o21ai_1 _6856_ (.B1(_2739_),
    .Y(_2740_),
    .A1(_0690_),
    .A2(net1500));
 sg13g2_a22oi_1 _6857_ (.Y(_2741_),
    .B1(_1099_),
    .B2(_2740_),
    .A2(net1405),
    .A1(\scl_bitbangengine0.n3737_o ));
 sg13g2_nand3_1 _6858_ (.B(_2738_),
    .C(_2741_),
    .A(net1269),
    .Y(_2742_));
 sg13g2_a21o_2 _6859_ (.A2(_2742_),
    .A1(_1940_),
    .B1(_2737_),
    .X(_2743_));
 sg13g2_mux2_1 _6860_ (.A0(net743),
    .A1(net1252),
    .S(net1188),
    .X(_0223_));
 sg13g2_nor2_1 _6861_ (.A(_1092_),
    .B(net1270),
    .Y(_2744_));
 sg13g2_mux2_1 _6862_ (.A0(net12),
    .A1(net4),
    .S(net1499),
    .X(_2745_));
 sg13g2_a22oi_1 _6863_ (.Y(_2746_),
    .B1(_1099_),
    .B2(_2745_),
    .A2(net1405),
    .A1(net1495));
 sg13g2_nand2_1 _6864_ (.Y(_2747_),
    .A(net12),
    .B(_1166_));
 sg13g2_nand3_1 _6865_ (.B(_2746_),
    .C(_2747_),
    .A(_2744_),
    .Y(_2748_));
 sg13g2_a22oi_1 _6866_ (.Y(_2749_),
    .B1(_1942_),
    .B2(_2748_),
    .A2(net1416),
    .A1(\s_out_3[3] ));
 sg13g2_nor2_1 _6867_ (.A(net837),
    .B(net1188),
    .Y(_2750_));
 sg13g2_a21oi_1 _6868_ (.A1(net1187),
    .A2(net1250),
    .Y(_0224_),
    .B1(_2750_));
 sg13g2_nand2_1 _6869_ (.Y(_2751_),
    .A(net13),
    .B(_1166_));
 sg13g2_mux2_1 _6870_ (.A0(net13),
    .A1(net5),
    .S(net1500),
    .X(_2752_));
 sg13g2_a22oi_1 _6871_ (.Y(_2753_),
    .B1(_1099_),
    .B2(_2752_),
    .A2(net1405),
    .A1(net1493));
 sg13g2_nand3_1 _6872_ (.B(_2751_),
    .C(_2753_),
    .A(_2744_),
    .Y(_2754_));
 sg13g2_a22oi_1 _6873_ (.Y(_2755_),
    .B1(_1944_),
    .B2(_2754_),
    .A2(net1416),
    .A1(net716));
 sg13g2_nor2_1 _6874_ (.A(net805),
    .B(net1187),
    .Y(_2756_));
 sg13g2_a21oi_1 _6875_ (.A1(net1187),
    .A2(net1247),
    .Y(_0225_),
    .B1(_2756_));
 sg13g2_mux2_1 _6876_ (.A0(net14),
    .A1(net6),
    .S(net1499),
    .X(_2757_));
 sg13g2_a22oi_1 _6877_ (.Y(_2758_),
    .B1(_2757_),
    .B2(_1101_),
    .A2(_1178_),
    .A1(net14));
 sg13g2_a22oi_1 _6878_ (.Y(_2759_),
    .B1(_1095_),
    .B2(_2758_),
    .A2(net1405),
    .A1(_0692_));
 sg13g2_or2_1 _6879_ (.X(_2760_),
    .B(_2759_),
    .A(net1270));
 sg13g2_a22oi_1 _6880_ (.Y(_2761_),
    .B1(_1946_),
    .B2(_2760_),
    .A2(net1416),
    .A1(\s_out_3[5] ));
 sg13g2_nor2_1 _6881_ (.A(net845),
    .B(net1188),
    .Y(_2762_));
 sg13g2_a21oi_1 _6882_ (.A1(net1187),
    .A2(net1245),
    .Y(_0226_),
    .B1(_2762_));
 sg13g2_nand3_1 _6883_ (.B(net7),
    .C(_1101_),
    .A(net1499),
    .Y(_2763_));
 sg13g2_a22oi_1 _6884_ (.Y(_2764_),
    .B1(_1095_),
    .B2(_2763_),
    .A2(net1405),
    .A1(_0694_));
 sg13g2_nor2_1 _6885_ (.A(net1271),
    .B(_2764_),
    .Y(_2765_));
 sg13g2_nor2_1 _6886_ (.A(_1949_),
    .B(_2765_),
    .Y(_2766_));
 sg13g2_a21oi_2 _6887_ (.B1(_2766_),
    .Y(_2767_),
    .A2(net1416),
    .A1(\s_out_3[6] ));
 sg13g2_nor2_1 _6888_ (.A(net894),
    .B(net1188),
    .Y(_2768_));
 sg13g2_a21oi_1 _6889_ (.A1(net1188),
    .A2(net1222),
    .Y(_0227_),
    .B1(_2768_));
 sg13g2_nand3_1 _6890_ (.B(net8),
    .C(_1101_),
    .A(net1499),
    .Y(_2769_));
 sg13g2_a22oi_1 _6891_ (.Y(_2770_),
    .B1(_1095_),
    .B2(_2769_),
    .A2(net1405),
    .A1(_0732_));
 sg13g2_or2_1 _6892_ (.X(_2771_),
    .B(_2770_),
    .A(net1271));
 sg13g2_a22oi_1 _6893_ (.Y(_2772_),
    .B1(_1951_),
    .B2(_2771_),
    .A2(net1416),
    .A1(net686));
 sg13g2_nor2_1 _6894_ (.A(net928),
    .B(net1187),
    .Y(_2773_));
 sg13g2_a21oi_1 _6895_ (.A1(net1187),
    .A2(net1242),
    .Y(_0228_),
    .B1(_2773_));
 sg13g2_o21ai_1 _6896_ (.B1(_1503_),
    .Y(_0229_),
    .A1(_0693_),
    .A2(_1499_));
 sg13g2_a21o_1 _6897_ (.A2(_1177_),
    .A1(net859),
    .B1(_1956_),
    .X(_0230_));
 sg13g2_nand2_1 _6898_ (.Y(_2774_),
    .A(\scl_bitbangengine0.n3336_o ),
    .B(_1201_));
 sg13g2_nand2_1 _6899_ (.Y(_2775_),
    .A(net595),
    .B(net1400));
 sg13g2_o21ai_1 _6900_ (.B1(_2775_),
    .Y(_0231_),
    .A1(_0732_),
    .A2(net1400));
 sg13g2_nor2_1 _6901_ (.A(_2654_),
    .B(_2663_),
    .Y(_2776_));
 sg13g2_nand2_1 _6902_ (.Y(_2777_),
    .A(net747),
    .B(_2776_));
 sg13g2_o21ai_1 _6903_ (.B1(_2777_),
    .Y(_0232_),
    .A1(_0747_),
    .A2(_2776_));
 sg13g2_nand2_1 _6904_ (.Y(_2778_),
    .A(net594),
    .B(net1400));
 sg13g2_o21ai_1 _6905_ (.B1(_2778_),
    .Y(_0233_),
    .A1(_0694_),
    .A2(net1400));
 sg13g2_nor2_1 _6906_ (.A(_0730_),
    .B(_1203_),
    .Y(_2779_));
 sg13g2_a221oi_1 _6907_ (.B2(net1801),
    .C1(_2779_),
    .B1(_1210_),
    .A1(net1890),
    .Y(_2780_),
    .A2(_1203_));
 sg13g2_nand2_1 _6908_ (.Y(_2781_),
    .A(\scl_bitbangengine0.n5905_q ),
    .B(\scl_bitbangengine0.n5915_q ));
 sg13g2_o21ai_1 _6909_ (.B1(\scl_bitbangengine0.n5915_q ),
    .Y(_2782_),
    .A1(_0131_),
    .A2(_2781_));
 sg13g2_a21oi_1 _6910_ (.A1(_0131_),
    .A2(_2781_),
    .Y(_2783_),
    .B1(_2782_));
 sg13g2_a21oi_2 _6911_ (.B1(_2783_),
    .Y(_2784_),
    .A2(_0772_),
    .A1(_0131_));
 sg13g2_xor2_1 _6912_ (.B(_2782_),
    .A(_0120_),
    .X(_2785_));
 sg13g2_nor3_1 _6913_ (.A(_0120_),
    .B(_0131_),
    .C(_2781_),
    .Y(_2786_));
 sg13g2_xor2_1 _6914_ (.B(\scl_bitbangengine0.n5915_q ),
    .A(_0132_),
    .X(_2787_));
 sg13g2_xnor2_1 _6915_ (.Y(_2788_),
    .A(_2786_),
    .B(_2787_));
 sg13g2_mux4_1 _6916_ (.S0(_2785_),
    .A0(net1493),
    .A1(\scl_bitbangengine0.n3258_o ),
    .A2(\scl_bitbangengine0.n3267_o ),
    .A3(net1492),
    .S1(_2784_),
    .X(_2789_));
 sg13g2_inv_1 _6917_ (.Y(_2790_),
    .A(_2789_));
 sg13g2_nor2_1 _6918_ (.A(\scl_bitbangengine0.n3737_o ),
    .B(_2784_),
    .Y(_2791_));
 sg13g2_a21oi_1 _6919_ (.A1(\scl_bitbangengine0.n3865_o ),
    .A2(_2784_),
    .Y(_2792_),
    .B1(_2791_));
 sg13g2_nor2_1 _6920_ (.A(net1502),
    .B(_2784_),
    .Y(_2793_));
 sg13g2_a21oi_1 _6921_ (.A1(_0083_),
    .A2(_2784_),
    .Y(_2794_),
    .B1(_2793_));
 sg13g2_nand2b_1 _6922_ (.Y(_2795_),
    .B(_2794_),
    .A_N(_2785_));
 sg13g2_a21oi_1 _6923_ (.A1(_2785_),
    .A2(_2792_),
    .Y(_2796_),
    .B1(_2788_));
 sg13g2_a22oi_1 _6924_ (.Y(_2797_),
    .B1(_2795_),
    .B2(_2796_),
    .A2(_2790_),
    .A1(_2788_));
 sg13g2_nor3_1 _6925_ (.A(\scl_bitbangengine0.n5905_q ),
    .B(_1337_),
    .C(_2797_),
    .Y(_2798_));
 sg13g2_nor2_1 _6926_ (.A(_2780_),
    .B(_2798_),
    .Y(_2799_));
 sg13g2_nand2_2 _6927_ (.Y(_2800_),
    .A(\scl_bitbangengine0.n5905_q ),
    .B(_1336_));
 sg13g2_o21ai_1 _6928_ (.B1(_2799_),
    .Y(_2801_),
    .A1(net1492),
    .A2(_2800_));
 sg13g2_inv_1 _6929_ (.Y(_0234_),
    .A(net1891));
 sg13g2_nand2_1 _6930_ (.Y(_2802_),
    .A(net597),
    .B(net1400));
 sg13g2_o21ai_1 _6931_ (.B1(_2802_),
    .Y(_0235_),
    .A1(_0692_),
    .A2(net1400));
 sg13g2_mux2_1 _6932_ (.A0(net1493),
    .A1(net1013),
    .S(net1401),
    .X(_0236_));
 sg13g2_a22oi_1 _6933_ (.Y(_2803_),
    .B1(net1373),
    .B2(\scl_bitbangengine0.n3267_o ),
    .A2(_1078_),
    .A1(net1166));
 sg13g2_inv_1 _6934_ (.Y(_0237_),
    .A(net1167));
 sg13g2_mux2_1 _6935_ (.A0(net1496),
    .A1(net1016),
    .S(net1400),
    .X(_0238_));
 sg13g2_a21o_1 _6936_ (.A2(_1078_),
    .A1(net1014),
    .B1(_2654_),
    .X(_0239_));
 sg13g2_nand2_1 _6937_ (.Y(_2804_),
    .A(net635),
    .B(net1401));
 sg13g2_o21ai_1 _6938_ (.B1(_2804_),
    .Y(_0240_),
    .A1(net1451),
    .A2(net1400));
 sg13g2_a21oi_1 _6939_ (.A1(_0691_),
    .A2(_1078_),
    .Y(_0241_),
    .B1(_2679_));
 sg13g2_nand2_1 _6940_ (.Y(_2805_),
    .A(net706),
    .B(net1401));
 sg13g2_o21ai_1 _6941_ (.B1(_2805_),
    .Y(_0242_),
    .A1(_0730_),
    .A2(net1401));
 sg13g2_nand2_1 _6942_ (.Y(_2806_),
    .A(_1081_),
    .B(_1098_));
 sg13g2_nand2_1 _6943_ (.Y(_2807_),
    .A(net1022),
    .B(_2806_));
 sg13g2_o21ai_1 _6944_ (.B1(_2807_),
    .Y(_0243_),
    .A1(_0747_),
    .A2(_2806_));
 sg13g2_nand2_1 _6945_ (.Y(_2808_),
    .A(net945),
    .B(net1401));
 sg13g2_o21ai_1 _6946_ (.B1(_2808_),
    .Y(_0244_),
    .A1(_0729_),
    .A2(net1401));
 sg13g2_nand2b_2 _6947_ (.Y(_2809_),
    .B(_2656_),
    .A_N(\scl_bitbangengine0.n5898_q[0] ));
 sg13g2_nand2_1 _6948_ (.Y(_2810_),
    .A(net994),
    .B(net1399));
 sg13g2_o21ai_1 _6949_ (.B1(_2810_),
    .Y(_0245_),
    .A1(_0692_),
    .A2(net1399));
 sg13g2_nor4_1 _6950_ (.A(_0927_),
    .B(_2708_),
    .C(_2710_),
    .D(_2713_),
    .Y(_2811_));
 sg13g2_and3_1 _6951_ (.X(_2812_),
    .A(net1504),
    .B(_0928_),
    .C(_2701_));
 sg13g2_mux2_1 _6952_ (.A0(net1098),
    .A1(_2812_),
    .S(_2811_),
    .X(_0246_));
 sg13g2_nor2_1 _6953_ (.A(net981),
    .B(net1414),
    .Y(_2813_));
 sg13g2_a21oi_1 _6954_ (.A1(_0692_),
    .A2(net1414),
    .Y(_0247_),
    .B1(_2813_));
 sg13g2_and2_1 _6955_ (.A(_0747_),
    .B(\scl_bitbangengine0.n3839_o ),
    .X(_2814_));
 sg13g2_o21ai_1 _6956_ (.B1(_0141_),
    .Y(_2815_),
    .A1(_0747_),
    .A2(\scl_bitbangengine0.n3839_o ));
 sg13g2_nor4_1 _6957_ (.A(net1492),
    .B(_1078_),
    .C(_2814_),
    .D(_2815_),
    .Y(_2816_));
 sg13g2_a21o_1 _6958_ (.A2(_1078_),
    .A1(net1088),
    .B1(_2816_),
    .X(_0248_));
 sg13g2_nor2_1 _6959_ (.A(net1129),
    .B(_1202_),
    .Y(_2817_));
 sg13g2_a21oi_1 _6960_ (.A1(_0692_),
    .A2(_1202_),
    .Y(_0249_),
    .B1(net1130));
 sg13g2_nand2_1 _6961_ (.Y(_2818_),
    .A(net888),
    .B(_2809_));
 sg13g2_o21ai_1 _6962_ (.B1(net889),
    .Y(_0250_),
    .A1(_0729_),
    .A2(_2809_));
 sg13g2_mux2_1 _6963_ (.A0(net1494),
    .A1(net1665),
    .S(net1399),
    .X(_0251_));
 sg13g2_mux2_1 _6964_ (.A0(net825),
    .A1(net1494),
    .S(net1414),
    .X(_0252_));
 sg13g2_nand3_1 _6965_ (.B(_1081_),
    .C(_1096_),
    .A(net1495),
    .Y(_2819_));
 sg13g2_mux2_1 _6966_ (.A0(net683),
    .A1(\scl_bitbangengine0.n5913_q ),
    .S(_2819_),
    .X(_0253_));
 sg13g2_nand2b_1 _6967_ (.Y(_2820_),
    .B(_1202_),
    .A_N(net1494));
 sg13g2_o21ai_1 _6968_ (.B1(_2820_),
    .Y(_2821_),
    .A1(net1832),
    .A2(_1202_));
 sg13g2_nor2_1 _6969_ (.A(_2797_),
    .B(_2800_),
    .Y(_2822_));
 sg13g2_a21oi_1 _6970_ (.A1(_2800_),
    .A2(_2821_),
    .Y(_0254_),
    .B1(_2822_));
 sg13g2_nand2_1 _6971_ (.Y(_2823_),
    .A(net576),
    .B(net1373));
 sg13g2_o21ai_1 _6972_ (.B1(_2823_),
    .Y(_0255_),
    .A1(_0772_),
    .A2(net1373));
 sg13g2_nand2_1 _6973_ (.Y(_2824_),
    .A(net885),
    .B(_1203_));
 sg13g2_o21ai_1 _6974_ (.B1(_2824_),
    .Y(_0256_),
    .A1(_0729_),
    .A2(_1203_));
 sg13g2_nor2_1 _6975_ (.A(net987),
    .B(_2655_),
    .Y(_2825_));
 sg13g2_xnor2_1 _6976_ (.Y(_2826_),
    .A(net1502),
    .B(net1498));
 sg13g2_a21oi_1 _6977_ (.A1(net1373),
    .A2(_2826_),
    .Y(_0257_),
    .B1(_2825_));
 sg13g2_mux2_1 _6978_ (.A0(net1496),
    .A1(net1690),
    .S(net1399),
    .X(_0258_));
 sg13g2_o21ai_1 _6979_ (.B1(net1373),
    .Y(_2827_),
    .A1(\scl_bitbangengine0.n3258_o ),
    .A2(net1493));
 sg13g2_o21ai_1 _6980_ (.B1(_2827_),
    .Y(_0259_),
    .A1(_0733_),
    .A2(_1077_));
 sg13g2_nand2_1 _6981_ (.Y(_2828_),
    .A(_2703_),
    .B(_2712_));
 sg13g2_nand2_1 _6982_ (.Y(_2829_),
    .A(_2701_),
    .B(_2717_));
 sg13g2_nand2_1 _6983_ (.Y(_2830_),
    .A(_2718_),
    .B(_2828_));
 sg13g2_nor2_1 _6984_ (.A(_2712_),
    .B(_2720_),
    .Y(_2831_));
 sg13g2_mux2_1 _6985_ (.A0(_2831_),
    .A1(net1638),
    .S(_2830_),
    .X(_0260_));
 sg13g2_nand2_1 _6986_ (.Y(_2832_),
    .A(net1031),
    .B(net1399));
 sg13g2_o21ai_1 _6987_ (.B1(_2832_),
    .Y(_0261_),
    .A1(_0731_),
    .A2(net1399));
 sg13g2_nand3_1 _6988_ (.B(_2707_),
    .C(_2829_),
    .A(_0926_),
    .Y(_2833_));
 sg13g2_nand3_1 _6989_ (.B(_2702_),
    .C(_2703_),
    .A(net1504),
    .Y(_2834_));
 sg13g2_nand2_1 _6990_ (.Y(_2835_),
    .A(net716),
    .B(_2833_));
 sg13g2_o21ai_1 _6991_ (.B1(net717),
    .Y(_0262_),
    .A1(_2833_),
    .A2(_2834_));
 sg13g2_a21oi_1 _6992_ (.A1(net828),
    .A2(_1327_),
    .Y(_2836_),
    .B1(_2592_));
 sg13g2_a21oi_1 _6993_ (.A1(_2592_),
    .A2(_2634_),
    .Y(_0263_),
    .B1(_2836_));
 sg13g2_nor2_1 _6994_ (.A(net738),
    .B(net1414),
    .Y(_2837_));
 sg13g2_a21oi_1 _6995_ (.A1(net1451),
    .A2(net1414),
    .Y(_0264_),
    .B1(_2837_));
 sg13g2_nor2_2 _6996_ (.A(net1903),
    .B(_1327_),
    .Y(_2838_));
 sg13g2_mux2_1 _6997_ (.A0(net1851),
    .A1(_2609_),
    .S(net1410),
    .X(_0265_));
 sg13g2_mux2_1 _6998_ (.A0(net1773),
    .A1(_2617_),
    .S(net1410),
    .X(_0266_));
 sg13g2_mux2_1 _6999_ (.A0(net823),
    .A1(_2625_),
    .S(net1410),
    .X(_0267_));
 sg13g2_nor2_1 _7000_ (.A(net1708),
    .B(net1410),
    .Y(_2839_));
 sg13g2_a21oi_1 _7001_ (.A1(_2607_),
    .A2(net1410),
    .Y(_0268_),
    .B1(_2839_));
 sg13g2_mux2_1 _7002_ (.A0(net1779),
    .A1(_2614_),
    .S(_2838_),
    .X(_0269_));
 sg13g2_mux2_1 _7003_ (.A0(net1668),
    .A1(_2623_),
    .S(_2838_),
    .X(_0270_));
 sg13g2_mux2_1 _7004_ (.A0(net856),
    .A1(_2630_),
    .S(_2838_),
    .X(_0271_));
 sg13g2_nor2_1 _7005_ (.A(net1745),
    .B(net1410),
    .Y(_2840_));
 sg13g2_a21oi_1 _7006_ (.A1(_2636_),
    .A2(net1410),
    .Y(_0272_),
    .B1(_2840_));
 sg13g2_mux2_1 _7007_ (.A0(net1693),
    .A1(_2634_),
    .S(net1410),
    .X(_0273_));
 sg13g2_nand2_1 _7008_ (.Y(_2841_),
    .A(net820),
    .B(_1203_));
 sg13g2_o21ai_1 _7009_ (.B1(_2841_),
    .Y(_0274_),
    .A1(net1451),
    .A2(_1203_));
 sg13g2_nor2_1 _7010_ (.A(net850),
    .B(_1206_),
    .Y(_2842_));
 sg13g2_a21oi_1 _7011_ (.A1(_0729_),
    .A2(_1206_),
    .Y(_0275_),
    .B1(net851));
 sg13g2_nand2_1 _7012_ (.Y(_2843_),
    .A(net861),
    .B(net1399));
 sg13g2_o21ai_1 _7013_ (.B1(_2843_),
    .Y(_0276_),
    .A1(_0730_),
    .A2(net1399));
 sg13g2_nor2_1 _7014_ (.A(net760),
    .B(net1414),
    .Y(_2844_));
 sg13g2_a21oi_1 _7015_ (.A1(_0730_),
    .A2(net1414),
    .Y(_0277_),
    .B1(_2844_));
 sg13g2_nor2_1 _7016_ (.A(net598),
    .B(net552),
    .Y(_2845_));
 sg13g2_nor2_1 _7017_ (.A(_0802_),
    .B(_2845_),
    .Y(_0278_));
 sg13g2_nand3b_1 _7018_ (.B(_2709_),
    .C(_0926_),
    .Y(_2846_),
    .A_N(_2713_));
 sg13g2_nand2_1 _7019_ (.Y(_2847_),
    .A(net1504),
    .B(_2710_));
 sg13g2_nand2_1 _7020_ (.Y(_2848_),
    .A(net674),
    .B(_2846_));
 sg13g2_o21ai_1 _7021_ (.B1(_2848_),
    .Y(_0284_),
    .A1(_2846_),
    .A2(_2847_));
 sg13g2_nor2_1 _7022_ (.A(net670),
    .B(net1361),
    .Y(_2849_));
 sg13g2_a21oi_1 _7023_ (.A1(net1361),
    .A2(_1880_),
    .Y(_0285_),
    .B1(_2849_));
 sg13g2_o21ai_1 _7024_ (.B1(_1858_),
    .Y(_0286_),
    .A1(_0710_),
    .A2(net1361));
 sg13g2_mux2_1 _7025_ (.A0(net658),
    .A1(\scl_fifo0.n2722_o[2] ),
    .S(net1361),
    .X(_0287_));
 sg13g2_nand2_1 _7026_ (.Y(_2850_),
    .A(net578),
    .B(_1857_));
 sg13g2_o21ai_1 _7027_ (.B1(net579),
    .Y(_0288_),
    .A1(_1857_),
    .A2(_1870_));
 sg13g2_o21ai_1 _7028_ (.B1(_1877_),
    .Y(_0289_),
    .A1(_0769_),
    .A2(_1856_));
 sg13g2_o21ai_1 _7029_ (.B1(_2718_),
    .Y(_2851_),
    .A1(_0928_),
    .A2(_2704_));
 sg13g2_nand2_1 _7030_ (.Y(_2852_),
    .A(net686),
    .B(_2851_));
 sg13g2_o21ai_1 _7031_ (.B1(_2852_),
    .Y(_0290_),
    .A1(_0690_),
    .A2(_2851_));
 sg13g2_nand4_1 _7032_ (.B(net1488),
    .C(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.s_m_value[0] ),
    .A(net1132),
    .Y(_2853_),
    .D(_2523_));
 sg13g2_a22oi_1 _7033_ (.Y(_0291_),
    .B1(net1133),
    .B2(_0713_),
    .A2(_2549_),
    .A1(_2523_));
 sg13g2_mux2_1 _7034_ (.A0(net540),
    .A1(net536),
    .S(_1516_),
    .X(_0292_));
 sg13g2_mux2_1 _7035_ (.A0(net532),
    .A1(net540),
    .S(net1368),
    .X(_0293_));
 sg13g2_mux2_1 _7036_ (.A0(net534),
    .A1(net532),
    .S(net1368),
    .X(_0294_));
 sg13g2_mux2_1 _7037_ (.A0(net533),
    .A1(net534),
    .S(net1368),
    .X(_0295_));
 sg13g2_mux2_1 _7038_ (.A0(net531),
    .A1(net533),
    .S(net1368),
    .X(_0296_));
 sg13g2_mux2_1 _7039_ (.A0(net535),
    .A1(net531),
    .S(net1368),
    .X(_0297_));
 sg13g2_nand2_1 _7040_ (.Y(_2854_),
    .A(net535),
    .B(net1368));
 sg13g2_o21ai_1 _7041_ (.B1(_2854_),
    .Y(_0298_),
    .A1(_0789_),
    .A2(net1368));
 sg13g2_nor4_2 _7042_ (.A(net1486),
    .B(net1487),
    .C(_1829_),
    .Y(_2855_),
    .D(_1832_));
 sg13g2_nor2_1 _7043_ (.A(_1834_),
    .B(_1836_),
    .Y(_2856_));
 sg13g2_a22oi_1 _7044_ (.Y(_2857_),
    .B1(_2855_),
    .B2(_2856_),
    .A2(_1829_),
    .A1(net755));
 sg13g2_inv_1 _7045_ (.Y(_0299_),
    .A(net756));
 sg13g2_nand3_1 _7046_ (.B(_2704_),
    .C(_2829_),
    .A(_0926_),
    .Y(_2858_));
 sg13g2_nand2_1 _7047_ (.Y(_2859_),
    .A(net689),
    .B(_2858_));
 sg13g2_nand3_1 _7048_ (.B(_2701_),
    .C(_2716_),
    .A(net1504),
    .Y(_2860_));
 sg13g2_o21ai_1 _7049_ (.B1(_2859_),
    .Y(_0300_),
    .A1(_2858_),
    .A2(_2860_));
 sg13g2_nand4_1 _7050_ (.B(\scl_fifo0.n2689_o[3] ),
    .C(net1364),
    .A(\scl_fifo0.n2689_o[2] ),
    .Y(_2861_),
    .D(_1851_));
 sg13g2_nand2_1 _7051_ (.Y(_2862_),
    .A(net672),
    .B(net1358));
 sg13g2_o21ai_1 _7052_ (.B1(_2862_),
    .Y(_0301_),
    .A1(net1454),
    .A2(net1357));
 sg13g2_nand2_1 _7053_ (.Y(_2863_),
    .A(net615),
    .B(net1357));
 sg13g2_o21ai_1 _7054_ (.B1(_2863_),
    .Y(_0302_),
    .A1(net1457),
    .A2(net1357));
 sg13g2_mux2_1 _7055_ (.A0(net1474),
    .A1(net1120),
    .S(net1357),
    .X(_0303_));
 sg13g2_nand2_1 _7056_ (.Y(_2864_),
    .A(net652),
    .B(net1358));
 sg13g2_o21ai_1 _7057_ (.B1(_2864_),
    .Y(_0304_),
    .A1(net1460),
    .A2(net1358));
 sg13g2_mux2_1 _7058_ (.A0(net1473),
    .A1(net1125),
    .S(net1357),
    .X(_0305_));
 sg13g2_mux2_1 _7059_ (.A0(net1470),
    .A1(net1122),
    .S(net1357),
    .X(_0306_));
 sg13g2_nor2_1 _7060_ (.A(net1465),
    .B(net1358),
    .Y(_2865_));
 sg13g2_a21oi_1 _7061_ (.A1(_0775_),
    .A2(net1357),
    .Y(_0307_),
    .B1(_2865_));
 sg13g2_mux2_1 _7062_ (.A0(net1464),
    .A1(net1061),
    .S(net1357),
    .X(_0308_));
 sg13g2_nand4_1 _7063_ (.B(\scl_fifo0.n2689_o[3] ),
    .C(net1364),
    .A(\scl_fifo0.n2689_o[2] ),
    .Y(_2866_),
    .D(_1850_));
 sg13g2_nand2_1 _7064_ (.Y(_2867_),
    .A(net585),
    .B(net1356));
 sg13g2_o21ai_1 _7065_ (.B1(_2867_),
    .Y(_0309_),
    .A1(net1452),
    .A2(net1356));
 sg13g2_nand2_1 _7066_ (.Y(_2868_),
    .A(net586),
    .B(net1356));
 sg13g2_o21ai_1 _7067_ (.B1(_2868_),
    .Y(_0310_),
    .A1(net1456),
    .A2(net1356));
 sg13g2_mux2_1 _7068_ (.A0(net1474),
    .A1(net964),
    .S(net1356),
    .X(_0311_));
 sg13g2_nand2_1 _7069_ (.Y(_2869_),
    .A(net587),
    .B(_2866_));
 sg13g2_o21ai_1 _7070_ (.B1(_2869_),
    .Y(_0312_),
    .A1(net1459),
    .A2(_2866_));
 sg13g2_mux2_1 _7071_ (.A0(net1471),
    .A1(net954),
    .S(net1356),
    .X(_0313_));
 sg13g2_mux2_1 _7072_ (.A0(net1468),
    .A1(net959),
    .S(net1356),
    .X(_0314_));
 sg13g2_mux2_1 _7073_ (.A0(net1466),
    .A1(net990),
    .S(_2866_),
    .X(_0315_));
 sg13g2_mux2_1 _7074_ (.A0(net1462),
    .A1(net907),
    .S(net1356),
    .X(_0316_));
 sg13g2_nor2_2 _7075_ (.A(\scl_fifo0.n2689_o[1] ),
    .B(\scl_fifo0.n2689_o[0] ),
    .Y(_2870_));
 sg13g2_nand4_1 _7076_ (.B(\scl_fifo0.n2689_o[3] ),
    .C(net1364),
    .A(\scl_fifo0.n2689_o[2] ),
    .Y(_2871_),
    .D(_2870_));
 sg13g2_nand2_1 _7077_ (.Y(_2872_),
    .A(net701),
    .B(net1355));
 sg13g2_o21ai_1 _7078_ (.B1(_2872_),
    .Y(_0317_),
    .A1(net1452),
    .A2(_2871_));
 sg13g2_nand2_1 _7079_ (.Y(_2873_),
    .A(net726),
    .B(net1355));
 sg13g2_o21ai_1 _7080_ (.B1(_2873_),
    .Y(_0318_),
    .A1(net1456),
    .A2(net1355));
 sg13g2_mux2_1 _7081_ (.A0(net1474),
    .A1(net1107),
    .S(net1355),
    .X(_0319_));
 sg13g2_nand2_1 _7082_ (.Y(_2874_),
    .A(net619),
    .B(_2871_));
 sg13g2_o21ai_1 _7083_ (.B1(_2874_),
    .Y(_0320_),
    .A1(net1459),
    .A2(_2871_));
 sg13g2_mux2_1 _7084_ (.A0(net1471),
    .A1(net1072),
    .S(net1355),
    .X(_0321_));
 sg13g2_mux2_1 _7085_ (.A0(net1468),
    .A1(net1095),
    .S(net1355),
    .X(_0322_));
 sg13g2_mux2_1 _7086_ (.A0(net1465),
    .A1(net1119),
    .S(net1355),
    .X(_0323_));
 sg13g2_mux2_1 _7087_ (.A0(net1462),
    .A1(net1064),
    .S(net1355),
    .X(_0324_));
 sg13g2_nor2b_1 _7088_ (.A(\scl_fifo0.n2689_o[2] ),
    .B_N(\scl_fifo0.n2689_o[3] ),
    .Y(_2875_));
 sg13g2_nor2b_2 _7089_ (.A(_1859_),
    .B_N(_2875_),
    .Y(_2876_));
 sg13g2_nor2_1 _7090_ (.A(net694),
    .B(_2876_),
    .Y(_2877_));
 sg13g2_a21oi_1 _7091_ (.A1(net1452),
    .A2(_2876_),
    .Y(_0325_),
    .B1(_2877_));
 sg13g2_nor2_1 _7092_ (.A(net637),
    .B(net1347),
    .Y(_2878_));
 sg13g2_a21oi_1 _7093_ (.A1(net1455),
    .A2(net1347),
    .Y(_0326_),
    .B1(_2878_));
 sg13g2_mux2_1 _7094_ (.A0(net773),
    .A1(net1474),
    .S(net1347),
    .X(_0327_));
 sg13g2_nor2_1 _7095_ (.A(net646),
    .B(net1347),
    .Y(_2879_));
 sg13g2_a21oi_1 _7096_ (.A1(net1459),
    .A2(net1347),
    .Y(_0328_),
    .B1(_2879_));
 sg13g2_mux2_1 _7097_ (.A0(net644),
    .A1(net1471),
    .S(net1347),
    .X(_0329_));
 sg13g2_mux2_1 _7098_ (.A0(net725),
    .A1(net1468),
    .S(net1347),
    .X(_0330_));
 sg13g2_mux2_1 _7099_ (.A0(net918),
    .A1(net1465),
    .S(_2876_),
    .X(_0331_));
 sg13g2_mux2_1 _7100_ (.A0(net677),
    .A1(net1462),
    .S(net1347),
    .X(_0332_));
 sg13g2_and2_1 _7101_ (.A(net1364),
    .B(_2875_),
    .X(_2880_));
 sg13g2_nand2_2 _7102_ (.Y(_2881_),
    .A(_1851_),
    .B(_2880_));
 sg13g2_nand2_1 _7103_ (.Y(_2882_),
    .A(net648),
    .B(_2881_));
 sg13g2_o21ai_1 _7104_ (.B1(_2882_),
    .Y(_0333_),
    .A1(net1452),
    .A2(_2881_));
 sg13g2_nand2_1 _7105_ (.Y(_2883_),
    .A(net636),
    .B(net1346));
 sg13g2_o21ai_1 _7106_ (.B1(_2883_),
    .Y(_0334_),
    .A1(net1455),
    .A2(net1346));
 sg13g2_mux2_1 _7107_ (.A0(net1474),
    .A1(net1063),
    .S(net1346),
    .X(_0335_));
 sg13g2_nand2_1 _7108_ (.Y(_2884_),
    .A(net707),
    .B(net1346));
 sg13g2_o21ai_1 _7109_ (.B1(_2884_),
    .Y(_0336_),
    .A1(net1458),
    .A2(net1346));
 sg13g2_mux2_1 _7110_ (.A0(net1471),
    .A1(net1065),
    .S(net1346),
    .X(_0337_));
 sg13g2_mux2_1 _7111_ (.A0(net1468),
    .A1(net1069),
    .S(net1346),
    .X(_0338_));
 sg13g2_mux2_1 _7112_ (.A0(net1465),
    .A1(net1036),
    .S(_2881_),
    .X(_0339_));
 sg13g2_mux2_1 _7113_ (.A0(net1462),
    .A1(net1047),
    .S(net1346),
    .X(_0340_));
 sg13g2_nor3_2 _7114_ (.A(\scl_fifo0.n2689_o[2] ),
    .B(\scl_fifo0.n2689_o[3] ),
    .C(_1849_),
    .Y(_2885_));
 sg13g2_nand2_2 _7115_ (.Y(_2886_),
    .A(_2870_),
    .B(_2885_));
 sg13g2_nand2_1 _7116_ (.Y(_2887_),
    .A(net655),
    .B(net1328));
 sg13g2_o21ai_1 _7117_ (.B1(_2887_),
    .Y(_0341_),
    .A1(net1452),
    .A2(net1328));
 sg13g2_nand2_1 _7118_ (.Y(_2888_),
    .A(net638),
    .B(net1328));
 sg13g2_o21ai_1 _7119_ (.B1(_2888_),
    .Y(_0342_),
    .A1(net1455),
    .A2(_2886_));
 sg13g2_mux2_1 _7120_ (.A0(net1475),
    .A1(net1099),
    .S(net1328),
    .X(_0343_));
 sg13g2_nand2_1 _7121_ (.Y(_2889_),
    .A(net656),
    .B(net1328));
 sg13g2_o21ai_1 _7122_ (.B1(_2889_),
    .Y(_0344_),
    .A1(net1458),
    .A2(net1328));
 sg13g2_mux2_1 _7123_ (.A0(net1471),
    .A1(net1569),
    .S(net1328),
    .X(_0345_));
 sg13g2_mux2_1 _7124_ (.A0(net1468),
    .A1(net1086),
    .S(net1328),
    .X(_0346_));
 sg13g2_mux2_1 _7125_ (.A0(net1465),
    .A1(net1091),
    .S(_2886_),
    .X(_0347_));
 sg13g2_mux2_1 _7126_ (.A0(net1462),
    .A1(net1141),
    .S(_2886_),
    .X(_0348_));
 sg13g2_nand2_1 _7127_ (.Y(_2890_),
    .A(_2870_),
    .B(_2880_));
 sg13g2_nand2_1 _7128_ (.Y(_2891_),
    .A(net645),
    .B(net1344));
 sg13g2_o21ai_1 _7129_ (.B1(_2891_),
    .Y(_0349_),
    .A1(net1452),
    .A2(net1345));
 sg13g2_nand2_1 _7130_ (.Y(_2892_),
    .A(net630),
    .B(net1344));
 sg13g2_o21ai_1 _7131_ (.B1(_2892_),
    .Y(_0350_),
    .A1(net1455),
    .A2(net1344));
 sg13g2_mux2_1 _7132_ (.A0(net1474),
    .A1(net1067),
    .S(net1345),
    .X(_0351_));
 sg13g2_nand2_1 _7133_ (.Y(_2893_),
    .A(net650),
    .B(net1344));
 sg13g2_o21ai_1 _7134_ (.B1(_2893_),
    .Y(_0352_),
    .A1(net1458),
    .A2(net1344));
 sg13g2_mux2_1 _7135_ (.A0(net1471),
    .A1(net1081),
    .S(net1344),
    .X(_0353_));
 sg13g2_mux2_1 _7136_ (.A0(net1468),
    .A1(net1121),
    .S(net1344),
    .X(_0354_));
 sg13g2_mux2_1 _7137_ (.A0(net1465),
    .A1(net1092),
    .S(net1345),
    .X(_0355_));
 sg13g2_mux2_1 _7138_ (.A0(net1462),
    .A1(net1111),
    .S(net1344),
    .X(_0356_));
 sg13g2_nor2b_1 _7139_ (.A(\scl_fifo0.n2689_o[3] ),
    .B_N(\scl_fifo0.n2689_o[2] ),
    .Y(_2894_));
 sg13g2_nor2b_2 _7140_ (.A(_1859_),
    .B_N(_2894_),
    .Y(_2895_));
 sg13g2_nor2_1 _7141_ (.A(net704),
    .B(_2895_),
    .Y(_2896_));
 sg13g2_a21oi_1 _7142_ (.A1(net1453),
    .A2(_2895_),
    .Y(_0357_),
    .B1(_2896_));
 sg13g2_nor2_1 _7143_ (.A(net842),
    .B(net1343),
    .Y(_2897_));
 sg13g2_a21oi_1 _7144_ (.A1(net1456),
    .A2(net1343),
    .Y(_0358_),
    .B1(_2897_));
 sg13g2_mux2_1 _7145_ (.A0(net664),
    .A1(net1475),
    .S(net1343),
    .X(_0359_));
 sg13g2_nor2_1 _7146_ (.A(net647),
    .B(net1343),
    .Y(_2898_));
 sg13g2_a21oi_1 _7147_ (.A1(net1459),
    .A2(_2895_),
    .Y(_0360_),
    .B1(_2898_));
 sg13g2_mux2_1 _7148_ (.A0(net657),
    .A1(net1472),
    .S(net1343),
    .X(_0361_));
 sg13g2_mux2_1 _7149_ (.A0(net793),
    .A1(net1469),
    .S(net1343),
    .X(_0362_));
 sg13g2_mux2_1 _7150_ (.A0(net732),
    .A1(net1466),
    .S(net1343),
    .X(_0363_));
 sg13g2_mux2_1 _7151_ (.A0(net715),
    .A1(net1463),
    .S(net1343),
    .X(_0364_));
 sg13g2_and2_1 _7152_ (.A(net1364),
    .B(_2894_),
    .X(_2899_));
 sg13g2_nand2_2 _7153_ (.Y(_2900_),
    .A(_1851_),
    .B(_2899_));
 sg13g2_nand2_1 _7154_ (.Y(_2901_),
    .A(net719),
    .B(_2900_));
 sg13g2_o21ai_1 _7155_ (.B1(_2901_),
    .Y(_0365_),
    .A1(net1453),
    .A2(_2900_));
 sg13g2_nand2_1 _7156_ (.Y(_2902_),
    .A(net663),
    .B(net1342));
 sg13g2_o21ai_1 _7157_ (.B1(_2902_),
    .Y(_0366_),
    .A1(net1456),
    .A2(net1342));
 sg13g2_mux2_1 _7158_ (.A0(net1475),
    .A1(net1045),
    .S(net1342),
    .X(_0367_));
 sg13g2_nand2_1 _7159_ (.Y(_2903_),
    .A(net691),
    .B(net1342));
 sg13g2_o21ai_1 _7160_ (.B1(_2903_),
    .Y(_0368_),
    .A1(net1458),
    .A2(net1342));
 sg13g2_mux2_1 _7161_ (.A0(net1472),
    .A1(net1087),
    .S(net1342),
    .X(_0369_));
 sg13g2_mux2_1 _7162_ (.A0(net1469),
    .A1(net1115),
    .S(_2900_),
    .X(_0370_));
 sg13g2_mux2_1 _7163_ (.A0(net1466),
    .A1(net1048),
    .S(net1342),
    .X(_0371_));
 sg13g2_mux2_1 _7164_ (.A0(net1463),
    .A1(net1073),
    .S(net1342),
    .X(_0372_));
 sg13g2_nand2_1 _7165_ (.Y(_2904_),
    .A(_1850_),
    .B(_2899_));
 sg13g2_nand2_1 _7166_ (.Y(_2905_),
    .A(net569),
    .B(net1341));
 sg13g2_o21ai_1 _7167_ (.B1(_2905_),
    .Y(_0373_),
    .A1(net1453),
    .A2(net1340));
 sg13g2_nand2_1 _7168_ (.Y(_2906_),
    .A(net592),
    .B(net1340));
 sg13g2_o21ai_1 _7169_ (.B1(_2906_),
    .Y(_0374_),
    .A1(net1455),
    .A2(net1340));
 sg13g2_mux2_1 _7170_ (.A0(net1475),
    .A1(net950),
    .S(net1341),
    .X(_0375_));
 sg13g2_nand2_1 _7171_ (.Y(_2907_),
    .A(net563),
    .B(net1340));
 sg13g2_o21ai_1 _7172_ (.B1(_2907_),
    .Y(_0376_),
    .A1(net1458),
    .A2(net1340));
 sg13g2_mux2_1 _7173_ (.A0(net1472),
    .A1(net973),
    .S(net1340),
    .X(_0377_));
 sg13g2_mux2_1 _7174_ (.A0(net1469),
    .A1(net998),
    .S(net1340),
    .X(_0378_));
 sg13g2_mux2_1 _7175_ (.A0(net1466),
    .A1(net970),
    .S(net1341),
    .X(_0379_));
 sg13g2_mux2_1 _7176_ (.A0(net1463),
    .A1(net1002),
    .S(net1340),
    .X(_0380_));
 sg13g2_nand2_1 _7177_ (.Y(_2908_),
    .A(_2870_),
    .B(_2899_));
 sg13g2_nand2_1 _7178_ (.Y(_2909_),
    .A(net662),
    .B(net1339));
 sg13g2_o21ai_1 _7179_ (.B1(_2909_),
    .Y(_0381_),
    .A1(net1453),
    .A2(net1338));
 sg13g2_nand2_1 _7180_ (.Y(_2910_),
    .A(net722),
    .B(net1338));
 sg13g2_o21ai_1 _7181_ (.B1(_2910_),
    .Y(_0382_),
    .A1(net1455),
    .A2(net1338));
 sg13g2_mux2_1 _7182_ (.A0(net1475),
    .A1(net1110),
    .S(net1339),
    .X(_0383_));
 sg13g2_nand2_1 _7183_ (.Y(_2911_),
    .A(net626),
    .B(net1338));
 sg13g2_o21ai_1 _7184_ (.B1(_2911_),
    .Y(_0384_),
    .A1(net1458),
    .A2(net1338));
 sg13g2_mux2_1 _7185_ (.A0(net1472),
    .A1(net1046),
    .S(net1338),
    .X(_0385_));
 sg13g2_mux2_1 _7186_ (.A0(net1469),
    .A1(net1108),
    .S(net1338),
    .X(_0386_));
 sg13g2_mux2_1 _7187_ (.A0(net1466),
    .A1(net1078),
    .S(net1339),
    .X(_0387_));
 sg13g2_mux2_1 _7188_ (.A0(net1463),
    .A1(net1118),
    .S(net1338),
    .X(_0388_));
 sg13g2_nor3_2 _7189_ (.A(\scl_fifo0.n2689_o[2] ),
    .B(\scl_fifo0.n2689_o[3] ),
    .C(_1859_),
    .Y(_2912_));
 sg13g2_nor2_1 _7190_ (.A(net699),
    .B(_2912_),
    .Y(_2913_));
 sg13g2_a21oi_1 _7191_ (.A1(net1453),
    .A2(net1337),
    .Y(_0389_),
    .B1(_2913_));
 sg13g2_nor2_1 _7192_ (.A(net665),
    .B(net1337),
    .Y(_2914_));
 sg13g2_a21oi_1 _7193_ (.A1(net1457),
    .A2(net1337),
    .Y(_0390_),
    .B1(_2914_));
 sg13g2_mux2_1 _7194_ (.A0(net709),
    .A1(net1475),
    .S(net1337),
    .X(_0391_));
 sg13g2_nor2_1 _7195_ (.A(net728),
    .B(net1337),
    .Y(_2915_));
 sg13g2_a21oi_1 _7196_ (.A1(net1459),
    .A2(net1337),
    .Y(_0392_),
    .B1(_2915_));
 sg13g2_mux2_1 _7197_ (.A0(net667),
    .A1(net1472),
    .S(net1337),
    .X(_0393_));
 sg13g2_mux2_1 _7198_ (.A0(net695),
    .A1(\s_m_pushdata_data[5] ),
    .S(_2912_),
    .X(_0394_));
 sg13g2_mux2_1 _7199_ (.A0(net660),
    .A1(net1466),
    .S(net1337),
    .X(_0395_));
 sg13g2_mux2_1 _7200_ (.A0(net680),
    .A1(net1464),
    .S(_2912_),
    .X(_0396_));
 sg13g2_nand2_2 _7201_ (.Y(_2916_),
    .A(_1850_),
    .B(_2885_));
 sg13g2_nand2_1 _7202_ (.Y(_2917_),
    .A(net573),
    .B(net1327));
 sg13g2_o21ai_1 _7203_ (.B1(_2917_),
    .Y(_0397_),
    .A1(net1452),
    .A2(net1327));
 sg13g2_nand2_1 _7204_ (.Y(_2918_),
    .A(net613),
    .B(_2916_));
 sg13g2_o21ai_1 _7205_ (.B1(_2918_),
    .Y(_0398_),
    .A1(net1455),
    .A2(_2916_));
 sg13g2_mux2_1 _7206_ (.A0(net1475),
    .A1(net979),
    .S(net1327),
    .X(_0399_));
 sg13g2_nand2_1 _7207_ (.Y(_2919_),
    .A(net593),
    .B(net1327));
 sg13g2_o21ai_1 _7208_ (.B1(_2919_),
    .Y(_0400_),
    .A1(net1458),
    .A2(net1327));
 sg13g2_mux2_1 _7209_ (.A0(net1471),
    .A1(net941),
    .S(net1327),
    .X(_0401_));
 sg13g2_mux2_1 _7210_ (.A0(net1468),
    .A1(net935),
    .S(net1327),
    .X(_0402_));
 sg13g2_mux2_1 _7211_ (.A0(net1465),
    .A1(net1025),
    .S(_2916_),
    .X(_0403_));
 sg13g2_mux2_1 _7212_ (.A0(net1462),
    .A1(net1005),
    .S(net1327),
    .X(_0404_));
 sg13g2_nand2_2 _7213_ (.Y(_2920_),
    .A(_1851_),
    .B(_2885_));
 sg13g2_nand2_1 _7214_ (.Y(_2921_),
    .A(net659),
    .B(net1326));
 sg13g2_o21ai_1 _7215_ (.B1(_2921_),
    .Y(_0405_),
    .A1(net1453),
    .A2(net1326));
 sg13g2_nand2_1 _7216_ (.Y(_2922_),
    .A(net712),
    .B(_2920_));
 sg13g2_o21ai_1 _7217_ (.B1(_2922_),
    .Y(_0406_),
    .A1(net1457),
    .A2(_2920_));
 sg13g2_mux2_1 _7218_ (.A0(net1475),
    .A1(net1114),
    .S(_2920_),
    .X(_0407_));
 sg13g2_nand2_1 _7219_ (.Y(_2923_),
    .A(net679),
    .B(net1326));
 sg13g2_o21ai_1 _7220_ (.B1(_2923_),
    .Y(_0408_),
    .A1(net1459),
    .A2(net1326));
 sg13g2_mux2_1 _7221_ (.A0(net1472),
    .A1(net1102),
    .S(net1326),
    .X(_0409_));
 sg13g2_mux2_1 _7222_ (.A0(net1470),
    .A1(net1139),
    .S(net1326),
    .X(_0410_));
 sg13g2_mux2_1 _7223_ (.A0(net1466),
    .A1(net1068),
    .S(net1326),
    .X(_0411_));
 sg13g2_mux2_1 _7224_ (.A0(net1463),
    .A1(net1148),
    .S(net1326),
    .X(_0412_));
 sg13g2_nor3_1 _7225_ (.A(\n352_o[11] ),
    .B(\n352_o[10] ),
    .C(_0828_),
    .Y(_2924_));
 sg13g2_nand2_1 _7226_ (.Y(_2925_),
    .A(\n352_o[8] ),
    .B(_2924_));
 sg13g2_nor3_1 _7227_ (.A(\usbfunction0.n2481_o[32] ),
    .B(\usbfunction0.n2481_o[35] ),
    .C(\usbfunction0.n2481_o[34] ),
    .Y(_2926_));
 sg13g2_and4_2 _7228_ (.A(\usbfunction0.n2481_o[33] ),
    .B(_1395_),
    .C(_1830_),
    .D(_2926_),
    .X(_2927_));
 sg13g2_nand4_1 _7229_ (.B(\s_m_packetdata_2_rewired[13] ),
    .C(_0812_),
    .A(\s_m_packetdata_2_rewired[15] ),
    .Y(_2928_),
    .D(_2927_));
 sg13g2_nor4_1 _7230_ (.A(_0180_),
    .B(\n352_o[12] ),
    .C(_2925_),
    .D(_2928_),
    .Y(_2929_));
 sg13g2_nor4_1 _7231_ (.A(\n352_o[3] ),
    .B(\n352_o[4] ),
    .C(\n352_o[5] ),
    .D(\n352_o[6] ),
    .Y(_2930_));
 sg13g2_nor4_1 _7232_ (.A(\n352_o[7] ),
    .B(\n352_o[0] ),
    .C(\n352_o[1] ),
    .D(\n352_o[2] ),
    .Y(_2931_));
 sg13g2_nand3_1 _7233_ (.B(_2930_),
    .C(_2931_),
    .A(_2929_),
    .Y(_2932_));
 sg13g2_o21ai_1 _7234_ (.B1(_2932_),
    .Y(_0413_),
    .A1(_0724_),
    .A2(_0812_));
 sg13g2_a21oi_1 _7235_ (.A1(net1267),
    .A2(_2400_),
    .Y(_2933_),
    .B1(_2414_));
 sg13g2_nor3_1 _7236_ (.A(net1263),
    .B(_2377_),
    .C(_2933_),
    .Y(_0414_));
 sg13g2_a22oi_1 _7237_ (.Y(_2934_),
    .B1(_2609_),
    .B2(_2591_),
    .A2(_2596_),
    .A1(_0735_));
 sg13g2_xor2_1 _7238_ (.B(_2934_),
    .A(net1360),
    .X(_0415_));
 sg13g2_nor2_1 _7239_ (.A(net1722),
    .B(net1360),
    .Y(_2935_));
 sg13g2_xnor2_1 _7240_ (.Y(_2936_),
    .A(\scl_bitbangengine0.n5920_q[0] ),
    .B(net1722));
 sg13g2_a22oi_1 _7241_ (.Y(_2937_),
    .B1(_2936_),
    .B2(_2596_),
    .A2(_2617_),
    .A1(net1413));
 sg13g2_a21oi_1 _7242_ (.A1(net1360),
    .A2(_2937_),
    .Y(_0416_),
    .B1(_2935_));
 sg13g2_o21ai_1 _7243_ (.B1(net1605),
    .Y(_2938_),
    .A1(\scl_bitbangengine0.n5920_q[0] ),
    .A2(\scl_bitbangengine0.n5920_q[1] ));
 sg13g2_nand2b_1 _7244_ (.Y(_2939_),
    .B(_2938_),
    .A_N(_2599_));
 sg13g2_a22oi_1 _7245_ (.Y(_2940_),
    .B1(_2939_),
    .B2(net1374),
    .A2(_2625_),
    .A1(net1413));
 sg13g2_nor2_1 _7246_ (.A(net1605),
    .B(net1359),
    .Y(_2941_));
 sg13g2_a21oi_1 _7247_ (.A1(net1359),
    .A2(_2940_),
    .Y(_0417_),
    .B1(_2941_));
 sg13g2_or4_1 _7248_ (.A(_0810_),
    .B(_1359_),
    .C(_1372_),
    .D(net1404),
    .X(_2942_));
 sg13g2_a21oi_1 _7249_ (.A1(\usbfunction0.n1974_o ),
    .A2(_1723_),
    .Y(_2943_),
    .B1(_2942_));
 sg13g2_o21ai_1 _7250_ (.B1(_2943_),
    .Y(_2944_),
    .A1(_1501_),
    .A2(_1502_));
 sg13g2_a21oi_2 _7251_ (.B1(_2944_),
    .Y(_2945_),
    .A2(_1040_),
    .A1(\usbfunction0.n2636_q ));
 sg13g2_a21o_1 _7252_ (.A2(_2945_),
    .A1(net1741),
    .B1(_2942_),
    .X(_0418_));
 sg13g2_nor3_1 _7253_ (.A(_1359_),
    .B(_1839_),
    .C(_2855_),
    .Y(_2946_));
 sg13g2_nand2b_1 _7254_ (.Y(_2947_),
    .B(_1552_),
    .A_N(_1393_));
 sg13g2_a21oi_1 _7255_ (.A1(net1486),
    .A2(_1397_),
    .Y(_2948_),
    .B1(_2947_));
 sg13g2_nor4_1 _7256_ (.A(net1380),
    .B(_1555_),
    .C(_1840_),
    .D(_2948_),
    .Y(_2949_));
 sg13g2_nand3_1 _7257_ (.B(_2946_),
    .C(_2949_),
    .A(_1629_),
    .Y(_2950_));
 sg13g2_nor2_1 _7258_ (.A(_1715_),
    .B(_2950_),
    .Y(_2951_));
 sg13g2_o21ai_1 _7259_ (.B1(net1415),
    .Y(_2952_),
    .A1(_1501_),
    .A2(_1502_));
 sg13g2_a21oi_1 _7260_ (.A1(_2951_),
    .A2(_2952_),
    .Y(_2953_),
    .B1(_1723_));
 sg13g2_nor4_1 _7261_ (.A(_0810_),
    .B(net1404),
    .C(_2945_),
    .D(_2953_),
    .Y(_2954_));
 sg13g2_a21o_1 _7262_ (.A2(_2945_),
    .A1(net1724),
    .B1(_2954_),
    .X(_0419_));
 sg13g2_nor2_1 _7263_ (.A(net599),
    .B(_2570_),
    .Y(_2955_));
 sg13g2_a21oi_1 _7264_ (.A1(net599),
    .A2(_1517_),
    .Y(_0420_),
    .B1(_2955_));
 sg13g2_nand2_1 _7265_ (.Y(_2956_),
    .A(_2173_),
    .B(_2530_));
 sg13g2_o21ai_1 _7266_ (.B1(_2956_),
    .Y(_2957_),
    .A1(_1517_),
    .A2(_2173_));
 sg13g2_nand2_1 _7267_ (.Y(_2958_),
    .A(net749),
    .B(net1352));
 sg13g2_nand2_1 _7268_ (.Y(_2959_),
    .A(_1533_),
    .B(_2171_));
 sg13g2_o21ai_1 _7269_ (.B1(_2959_),
    .Y(_2960_),
    .A1(_0789_),
    .A2(_2171_));
 sg13g2_xnor2_1 _7270_ (.Y(_2961_),
    .A(_2179_),
    .B(_2960_));
 sg13g2_nand2_2 _7271_ (.Y(_2962_),
    .A(_0780_),
    .B(_2961_));
 sg13g2_nand2_1 _7272_ (.Y(_2963_),
    .A(_0689_),
    .B(_2962_));
 sg13g2_nor2_1 _7273_ (.A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[1] ),
    .B(_2176_),
    .Y(_2964_));
 sg13g2_nor4_1 _7274_ (.A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[7] ),
    .B(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[8] ),
    .C(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[9] ),
    .D(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[10] ),
    .Y(_2965_));
 sg13g2_nor4_1 _7275_ (.A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[2] ),
    .B(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[3] ),
    .C(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[4] ),
    .D(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[5] ),
    .Y(_2966_));
 sg13g2_nand4_1 _7276_ (.B(_0715_),
    .C(_2965_),
    .A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.in_unnamed ),
    .Y(_2967_),
    .D(_2966_));
 sg13g2_or4_1 _7277_ (.A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[1] ),
    .B(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[6] ),
    .C(_2176_),
    .D(_2962_),
    .X(_2968_));
 sg13g2_o21ai_1 _7278_ (.B1(_2963_),
    .Y(_2969_),
    .A1(_2967_),
    .A2(_2968_));
 sg13g2_nor2_1 _7279_ (.A(net711),
    .B(_2176_),
    .Y(_2970_));
 sg13g2_xnor2_1 _7280_ (.Y(_2971_),
    .A(_2962_),
    .B(_2970_));
 sg13g2_nor2_2 _7281_ (.A(_2176_),
    .B(net1353),
    .Y(_2972_));
 sg13g2_nor3_1 _7282_ (.A(net610),
    .B(_2176_),
    .C(net1353),
    .Y(_2973_));
 sg13g2_nand4_1 _7283_ (.B(_0759_),
    .C(_2969_),
    .A(net736),
    .Y(_2974_),
    .D(_2973_));
 sg13g2_o21ai_1 _7284_ (.B1(_2958_),
    .Y(_0421_),
    .A1(_2971_),
    .A2(_2974_));
 sg13g2_nor3_1 _7285_ (.A(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7654_q[1] ),
    .B(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7654_q[0] ),
    .C(_0043_),
    .Y(_2975_));
 sg13g2_a21oi_1 _7286_ (.A1(net540),
    .A2(_2570_),
    .Y(_2976_),
    .B1(_2975_));
 sg13g2_o21ai_1 _7287_ (.B1(_2976_),
    .Y(_0422_),
    .A1(_0689_),
    .A2(_2570_));
 sg13g2_nor2_1 _7288_ (.A(net849),
    .B(net1224),
    .Y(_2977_));
 sg13g2_a21oi_1 _7289_ (.A1(net1224),
    .A2(net1255),
    .Y(_0423_),
    .B1(_2977_));
 sg13g2_nor2_1 _7290_ (.A(net813),
    .B(net1223),
    .Y(_2978_));
 sg13g2_a21oi_1 _7291_ (.A1(net1223),
    .A2(net1253),
    .Y(_0424_),
    .B1(_2978_));
 sg13g2_mux2_1 _7292_ (.A0(net880),
    .A1(net1251),
    .S(net1224),
    .X(_0425_));
 sg13g2_nor2_1 _7293_ (.A(net803),
    .B(net1223),
    .Y(_2979_));
 sg13g2_a21oi_1 _7294_ (.A1(net1223),
    .A2(net1249),
    .Y(_0426_),
    .B1(_2979_));
 sg13g2_nor2_1 _7295_ (.A(net730),
    .B(net1224),
    .Y(_2980_));
 sg13g2_a21oi_1 _7296_ (.A1(net1224),
    .A2(net1246),
    .Y(_0427_),
    .B1(_2980_));
 sg13g2_nor2_1 _7297_ (.A(net848),
    .B(net1223),
    .Y(_2981_));
 sg13g2_a21oi_1 _7298_ (.A1(net1223),
    .A2(net1244),
    .Y(_0428_),
    .B1(_2981_));
 sg13g2_nor2_1 _7299_ (.A(net944),
    .B(net1223),
    .Y(_2982_));
 sg13g2_a21oi_1 _7300_ (.A1(net1223),
    .A2(net1221),
    .Y(_0429_),
    .B1(_2982_));
 sg13g2_nor2_1 _7301_ (.A(net800),
    .B(net1224),
    .Y(_2983_));
 sg13g2_a21oi_1 _7302_ (.A1(net1224),
    .A2(net1242),
    .Y(_0430_),
    .B1(_2983_));
 sg13g2_nand2b_2 _7303_ (.Y(_2984_),
    .B(\scl_fifo1.n6229_o[1] ),
    .A_N(\scl_fifo1.n6229_o[0] ));
 sg13g2_nor3_2 _7304_ (.A(net1257),
    .B(_1994_),
    .C(_2984_),
    .Y(_2985_));
 sg13g2_nor2_1 _7305_ (.A(net763),
    .B(net1220),
    .Y(_2986_));
 sg13g2_a21oi_1 _7306_ (.A1(net1255),
    .A2(net1220),
    .Y(_0431_),
    .B1(_2986_));
 sg13g2_nor2_1 _7307_ (.A(net865),
    .B(net1219),
    .Y(_2987_));
 sg13g2_a21oi_1 _7308_ (.A1(net1253),
    .A2(net1219),
    .Y(_0432_),
    .B1(_2987_));
 sg13g2_mux2_1 _7309_ (.A0(net923),
    .A1(net1251),
    .S(net1220),
    .X(_0433_));
 sg13g2_nor2_1 _7310_ (.A(net830),
    .B(net1219),
    .Y(_2988_));
 sg13g2_a21oi_1 _7311_ (.A1(net1249),
    .A2(net1219),
    .Y(_0434_),
    .B1(_2988_));
 sg13g2_nor2_1 _7312_ (.A(net916),
    .B(net1220),
    .Y(_2989_));
 sg13g2_a21oi_1 _7313_ (.A1(net1246),
    .A2(net1220),
    .Y(_0435_),
    .B1(_2989_));
 sg13g2_nor2_1 _7314_ (.A(net960),
    .B(net1219),
    .Y(_2990_));
 sg13g2_a21oi_1 _7315_ (.A1(net1244),
    .A2(net1219),
    .Y(_0436_),
    .B1(_2990_));
 sg13g2_nor2_1 _7316_ (.A(net754),
    .B(net1219),
    .Y(_2991_));
 sg13g2_a21oi_1 _7317_ (.A1(net1221),
    .A2(net1219),
    .Y(_0437_),
    .B1(_2991_));
 sg13g2_nor2_1 _7318_ (.A(net783),
    .B(net1220),
    .Y(_2992_));
 sg13g2_a21oi_1 _7319_ (.A1(net1243),
    .A2(net1220),
    .Y(_0438_),
    .B1(_2992_));
 sg13g2_nand2b_2 _7320_ (.Y(_2993_),
    .B(\scl_fifo1.n6229_o[0] ),
    .A_N(\scl_fifo1.n6229_o[1] ));
 sg13g2_nor3_1 _7321_ (.A(net1257),
    .B(_1994_),
    .C(_2993_),
    .Y(_2994_));
 sg13g2_nor2_1 _7322_ (.A(net816),
    .B(net1218),
    .Y(_2995_));
 sg13g2_a21oi_1 _7323_ (.A1(net1256),
    .A2(net1218),
    .Y(_0439_),
    .B1(_2995_));
 sg13g2_nor2_1 _7324_ (.A(net806),
    .B(net1217),
    .Y(_2996_));
 sg13g2_a21oi_1 _7325_ (.A1(net1253),
    .A2(net1217),
    .Y(_0440_),
    .B1(_2996_));
 sg13g2_mux2_1 _7326_ (.A0(net968),
    .A1(net1251),
    .S(net1218),
    .X(_0441_));
 sg13g2_nor2_1 _7327_ (.A(net834),
    .B(net1218),
    .Y(_2997_));
 sg13g2_a21oi_1 _7328_ (.A1(net1249),
    .A2(net1218),
    .Y(_0442_),
    .B1(_2997_));
 sg13g2_nor2_1 _7329_ (.A(net780),
    .B(net1218),
    .Y(_2998_));
 sg13g2_a21oi_1 _7330_ (.A1(net1246),
    .A2(net1218),
    .Y(_0443_),
    .B1(_2998_));
 sg13g2_nor2_1 _7331_ (.A(net899),
    .B(net1217),
    .Y(_2999_));
 sg13g2_a21oi_1 _7332_ (.A1(net1244),
    .A2(net1217),
    .Y(_0444_),
    .B1(_2999_));
 sg13g2_nor2_1 _7333_ (.A(net943),
    .B(net1217),
    .Y(_3000_));
 sg13g2_a21oi_1 _7334_ (.A1(net1221),
    .A2(net1217),
    .Y(_0445_),
    .B1(_3000_));
 sg13g2_nor2_1 _7335_ (.A(net983),
    .B(net1217),
    .Y(_3001_));
 sg13g2_a21oi_1 _7336_ (.A1(net1243),
    .A2(net1217),
    .Y(_0446_),
    .B1(_3001_));
 sg13g2_nor2_1 _7337_ (.A(_1991_),
    .B(_1994_),
    .Y(_3002_));
 sg13g2_nor2_1 _7338_ (.A(net955),
    .B(net1186),
    .Y(_3003_));
 sg13g2_a21oi_1 _7339_ (.A1(net1256),
    .A2(net1186),
    .Y(_0447_),
    .B1(_3003_));
 sg13g2_nor2_1 _7340_ (.A(net742),
    .B(net1185),
    .Y(_3004_));
 sg13g2_a21oi_1 _7341_ (.A1(net1253),
    .A2(net1185),
    .Y(_0448_),
    .B1(_3004_));
 sg13g2_mux2_1 _7342_ (.A0(net733),
    .A1(net1251),
    .S(net1186),
    .X(_0449_));
 sg13g2_nor2_1 _7343_ (.A(net784),
    .B(net1185),
    .Y(_3005_));
 sg13g2_a21oi_1 _7344_ (.A1(net1249),
    .A2(net1185),
    .Y(_0450_),
    .B1(_3005_));
 sg13g2_nor2_1 _7345_ (.A(net822),
    .B(net1186),
    .Y(_3006_));
 sg13g2_a21oi_1 _7346_ (.A1(net1246),
    .A2(net1186),
    .Y(_0451_),
    .B1(_3006_));
 sg13g2_nor2_1 _7347_ (.A(net801),
    .B(net1185),
    .Y(_3007_));
 sg13g2_a21oi_1 _7348_ (.A1(net1244),
    .A2(net1185),
    .Y(_0452_),
    .B1(_3007_));
 sg13g2_nor2_1 _7349_ (.A(net905),
    .B(net1185),
    .Y(_3008_));
 sg13g2_a21oi_1 _7350_ (.A1(net1221),
    .A2(net1185),
    .Y(_0453_),
    .B1(_3008_));
 sg13g2_nor2_1 _7351_ (.A(net847),
    .B(net1186),
    .Y(_3009_));
 sg13g2_a21oi_1 _7352_ (.A1(net1243),
    .A2(net1186),
    .Y(_0454_),
    .B1(_3009_));
 sg13g2_nand2b_2 _7353_ (.Y(_3010_),
    .B(\scl_fifo1.n6229_o[3] ),
    .A_N(\scl_fifo1.n6229_o[2] ));
 sg13g2_nor2_1 _7354_ (.A(_1990_),
    .B(_3010_),
    .Y(_3011_));
 sg13g2_nor2_1 _7355_ (.A(net855),
    .B(net1216),
    .Y(_3012_));
 sg13g2_a21oi_1 _7356_ (.A1(net1256),
    .A2(net1216),
    .Y(_0455_),
    .B1(_3012_));
 sg13g2_nor2_1 _7357_ (.A(net708),
    .B(net1215),
    .Y(_3013_));
 sg13g2_a21oi_1 _7358_ (.A1(net1253),
    .A2(net1215),
    .Y(_0456_),
    .B1(_3013_));
 sg13g2_mux2_1 _7359_ (.A0(net957),
    .A1(net1251),
    .S(net1216),
    .X(_0457_));
 sg13g2_nor2_1 _7360_ (.A(net953),
    .B(net1215),
    .Y(_3014_));
 sg13g2_a21oi_1 _7361_ (.A1(net1249),
    .A2(net1215),
    .Y(_0458_),
    .B1(_3014_));
 sg13g2_nor2_1 _7362_ (.A(net952),
    .B(net1215),
    .Y(_3015_));
 sg13g2_a21oi_1 _7363_ (.A1(net1248),
    .A2(net1215),
    .Y(_0459_),
    .B1(_3015_));
 sg13g2_nor2_1 _7364_ (.A(net814),
    .B(net1216),
    .Y(_3016_));
 sg13g2_a21oi_1 _7365_ (.A1(net1244),
    .A2(net1216),
    .Y(_0460_),
    .B1(_3016_));
 sg13g2_nor2_1 _7366_ (.A(net729),
    .B(net1215),
    .Y(_3017_));
 sg13g2_a21oi_1 _7367_ (.A1(net1221),
    .A2(net1215),
    .Y(_0461_),
    .B1(_3017_));
 sg13g2_nor2_1 _7368_ (.A(net770),
    .B(net1216),
    .Y(_3018_));
 sg13g2_a21oi_1 _7369_ (.A1(net1243),
    .A2(net1216),
    .Y(_0462_),
    .B1(_3018_));
 sg13g2_nor3_1 _7370_ (.A(net1257),
    .B(_2984_),
    .C(_3010_),
    .Y(_3019_));
 sg13g2_nor2_1 _7371_ (.A(net839),
    .B(net1214),
    .Y(_3020_));
 sg13g2_a21oi_1 _7372_ (.A1(net1256),
    .A2(net1214),
    .Y(_0463_),
    .B1(_3020_));
 sg13g2_nor2_1 _7373_ (.A(net949),
    .B(net1212),
    .Y(_3021_));
 sg13g2_a21oi_1 _7374_ (.A1(net1253),
    .A2(net1212),
    .Y(_0464_),
    .B1(_3021_));
 sg13g2_mux2_1 _7375_ (.A0(net824),
    .A1(net1251),
    .S(net1214),
    .X(_0465_));
 sg13g2_nor2_1 _7376_ (.A(net1017),
    .B(net1212),
    .Y(_3022_));
 sg13g2_a21oi_1 _7377_ (.A1(net1249),
    .A2(net1212),
    .Y(_0466_),
    .B1(_3022_));
 sg13g2_nor2_1 _7378_ (.A(net883),
    .B(net1212),
    .Y(_3023_));
 sg13g2_a21oi_1 _7379_ (.A1(net1248),
    .A2(net1212),
    .Y(_0467_),
    .B1(_3023_));
 sg13g2_nor2_1 _7380_ (.A(net792),
    .B(net1213),
    .Y(_3024_));
 sg13g2_a21oi_1 _7381_ (.A1(net1244),
    .A2(net1213),
    .Y(_0468_),
    .B1(_3024_));
 sg13g2_nor2_1 _7382_ (.A(net980),
    .B(net1213),
    .Y(_3025_));
 sg13g2_a21oi_1 _7383_ (.A1(net1221),
    .A2(net1213),
    .Y(_0469_),
    .B1(_3025_));
 sg13g2_nor2_1 _7384_ (.A(net858),
    .B(net1212),
    .Y(_3026_));
 sg13g2_a21oi_1 _7385_ (.A1(net1243),
    .A2(net1212),
    .Y(_0470_),
    .B1(_3026_));
 sg13g2_nor3_1 _7386_ (.A(net1257),
    .B(_2993_),
    .C(_3010_),
    .Y(_3027_));
 sg13g2_nor2_1 _7387_ (.A(net867),
    .B(net1211),
    .Y(_3028_));
 sg13g2_a21oi_1 _7388_ (.A1(net1256),
    .A2(net1211),
    .Y(_0471_),
    .B1(_3028_));
 sg13g2_nor2_1 _7389_ (.A(net844),
    .B(net1210),
    .Y(_3029_));
 sg13g2_a21oi_1 _7390_ (.A1(net1253),
    .A2(net1210),
    .Y(_0472_),
    .B1(_3029_));
 sg13g2_mux2_1 _7391_ (.A0(net863),
    .A1(net1251),
    .S(net1211),
    .X(_0473_));
 sg13g2_nor2_1 _7392_ (.A(net951),
    .B(net1210),
    .Y(_3030_));
 sg13g2_a21oi_1 _7393_ (.A1(net1249),
    .A2(net1210),
    .Y(_0474_),
    .B1(_3030_));
 sg13g2_nor2_1 _7394_ (.A(net804),
    .B(net1211),
    .Y(_3031_));
 sg13g2_a21oi_1 _7395_ (.A1(net1246),
    .A2(net1211),
    .Y(_0475_),
    .B1(_3031_));
 sg13g2_nor2_1 _7396_ (.A(net982),
    .B(net1210),
    .Y(_3032_));
 sg13g2_a21oi_1 _7397_ (.A1(net1244),
    .A2(net1210),
    .Y(_0476_),
    .B1(_3032_));
 sg13g2_nor2_1 _7398_ (.A(net748),
    .B(net1210),
    .Y(_3033_));
 sg13g2_a21oi_1 _7399_ (.A1(net1221),
    .A2(net1210),
    .Y(_0477_),
    .B1(_3033_));
 sg13g2_nor2_1 _7400_ (.A(net891),
    .B(net1211),
    .Y(_3034_));
 sg13g2_a21oi_1 _7401_ (.A1(net1243),
    .A2(net1211),
    .Y(_0478_),
    .B1(_3034_));
 sg13g2_nor4_2 _7402_ (.A(\scl_fifo1.n6229_o[0] ),
    .B(\scl_fifo1.n6229_o[1] ),
    .C(net1257),
    .Y(_3035_),
    .D(_3010_));
 sg13g2_nor2_1 _7403_ (.A(net731),
    .B(net1209),
    .Y(_3036_));
 sg13g2_a21oi_1 _7404_ (.A1(net1256),
    .A2(net1209),
    .Y(_0479_),
    .B1(_3036_));
 sg13g2_nor2_1 _7405_ (.A(net607),
    .B(net1208),
    .Y(_3037_));
 sg13g2_a21oi_1 _7406_ (.A1(net1253),
    .A2(net1208),
    .Y(_0480_),
    .B1(_3037_));
 sg13g2_mux2_1 _7407_ (.A0(net854),
    .A1(net1251),
    .S(net1209),
    .X(_0481_));
 sg13g2_nor2_1 _7408_ (.A(net682),
    .B(net1208),
    .Y(_3038_));
 sg13g2_a21oi_1 _7409_ (.A1(net1249),
    .A2(net1208),
    .Y(_0482_),
    .B1(_3038_));
 sg13g2_nor2_1 _7410_ (.A(net769),
    .B(net1209),
    .Y(_3039_));
 sg13g2_a21oi_1 _7411_ (.A1(net1246),
    .A2(net1209),
    .Y(_0483_),
    .B1(_3039_));
 sg13g2_nor2_1 _7412_ (.A(net685),
    .B(net1208),
    .Y(_3040_));
 sg13g2_a21oi_1 _7413_ (.A1(net1244),
    .A2(net1208),
    .Y(_0484_),
    .B1(_3040_));
 sg13g2_nor2_1 _7414_ (.A(net757),
    .B(net1208),
    .Y(_3041_));
 sg13g2_a21oi_1 _7415_ (.A1(net1221),
    .A2(net1208),
    .Y(_0485_),
    .B1(_3041_));
 sg13g2_nor2_1 _7416_ (.A(net744),
    .B(net1209),
    .Y(_3042_));
 sg13g2_a21oi_1 _7417_ (.A1(net1243),
    .A2(net1209),
    .Y(_0486_),
    .B1(_3042_));
 sg13g2_nand2b_2 _7418_ (.Y(_3043_),
    .B(\scl_fifo1.n6229_o[2] ),
    .A_N(\scl_fifo1.n6229_o[3] ));
 sg13g2_nor2_1 _7419_ (.A(_1990_),
    .B(_3043_),
    .Y(_3044_));
 sg13g2_nor2_1 _7420_ (.A(net991),
    .B(net1207),
    .Y(_3045_));
 sg13g2_a21oi_1 _7421_ (.A1(net1256),
    .A2(net1207),
    .Y(_0487_),
    .B1(_3045_));
 sg13g2_nor2_1 _7422_ (.A(net720),
    .B(net1206),
    .Y(_3046_));
 sg13g2_a21oi_1 _7423_ (.A1(net1254),
    .A2(net1206),
    .Y(_0488_),
    .B1(_3046_));
 sg13g2_mux2_1 _7424_ (.A0(net922),
    .A1(net1252),
    .S(net1206),
    .X(_0489_));
 sg13g2_nor2_1 _7425_ (.A(net739),
    .B(net1206),
    .Y(_3047_));
 sg13g2_a21oi_1 _7426_ (.A1(net1250),
    .A2(net1206),
    .Y(_0490_),
    .B1(_3047_));
 sg13g2_nor2_1 _7427_ (.A(net872),
    .B(net1207),
    .Y(_3048_));
 sg13g2_a21oi_1 _7428_ (.A1(net1247),
    .A2(net1207),
    .Y(_0491_),
    .B1(_3048_));
 sg13g2_nor2_1 _7429_ (.A(net741),
    .B(net1207),
    .Y(_3049_));
 sg13g2_a21oi_1 _7430_ (.A1(net1245),
    .A2(net1206),
    .Y(_0492_),
    .B1(_3049_));
 sg13g2_nor2_1 _7431_ (.A(net799),
    .B(net1206),
    .Y(_3050_));
 sg13g2_a21oi_1 _7432_ (.A1(net1222),
    .A2(net1206),
    .Y(_0493_),
    .B1(_3050_));
 sg13g2_nor2_1 _7433_ (.A(net875),
    .B(net1207),
    .Y(_3051_));
 sg13g2_a21oi_1 _7434_ (.A1(net1242),
    .A2(net1207),
    .Y(_0494_),
    .B1(_3051_));
 sg13g2_nor3_2 _7435_ (.A(net1258),
    .B(_2984_),
    .C(_3043_),
    .Y(_3052_));
 sg13g2_nor2_1 _7436_ (.A(net838),
    .B(net1204),
    .Y(_3053_));
 sg13g2_a21oi_1 _7437_ (.A1(_2729_),
    .A2(net1204),
    .Y(_0495_),
    .B1(_3053_));
 sg13g2_nor2_1 _7438_ (.A(net853),
    .B(net1205),
    .Y(_3054_));
 sg13g2_a21oi_1 _7439_ (.A1(net1254),
    .A2(net1205),
    .Y(_0496_),
    .B1(_3054_));
 sg13g2_mux2_1 _7440_ (.A0(net937),
    .A1(net1252),
    .S(net1204),
    .X(_0497_));
 sg13g2_nor2_1 _7441_ (.A(net906),
    .B(net1205),
    .Y(_3055_));
 sg13g2_a21oi_1 _7442_ (.A1(net1250),
    .A2(net1205),
    .Y(_0498_),
    .B1(_3055_));
 sg13g2_nor2_1 _7443_ (.A(net961),
    .B(net1204),
    .Y(_3056_));
 sg13g2_a21oi_1 _7444_ (.A1(net1247),
    .A2(net1204),
    .Y(_0499_),
    .B1(_3056_));
 sg13g2_nor2_1 _7445_ (.A(net759),
    .B(net1205),
    .Y(_3057_));
 sg13g2_a21oi_1 _7446_ (.A1(net1245),
    .A2(net1204),
    .Y(_0500_),
    .B1(_3057_));
 sg13g2_nor2_1 _7447_ (.A(net965),
    .B(net1205),
    .Y(_3058_));
 sg13g2_a21oi_1 _7448_ (.A1(net1222),
    .A2(net1205),
    .Y(_0501_),
    .B1(_3058_));
 sg13g2_nor2_1 _7449_ (.A(net929),
    .B(net1204),
    .Y(_3059_));
 sg13g2_a21oi_1 _7450_ (.A1(net1242),
    .A2(net1204),
    .Y(_0502_),
    .B1(_3059_));
 sg13g2_nor3_2 _7451_ (.A(net1258),
    .B(_2993_),
    .C(_3043_),
    .Y(_3060_));
 sg13g2_nor2_1 _7452_ (.A(net904),
    .B(net1202),
    .Y(_3061_));
 sg13g2_a21oi_1 _7453_ (.A1(net1255),
    .A2(net1202),
    .Y(_0503_),
    .B1(_3061_));
 sg13g2_nor2_1 _7454_ (.A(net930),
    .B(net1203),
    .Y(_3062_));
 sg13g2_a21oi_1 _7455_ (.A1(net1254),
    .A2(net1203),
    .Y(_0504_),
    .B1(_3062_));
 sg13g2_mux2_1 _7456_ (.A0(net978),
    .A1(net1252),
    .S(net1203),
    .X(_0505_));
 sg13g2_nor2_1 _7457_ (.A(net740),
    .B(net1203),
    .Y(_3063_));
 sg13g2_a21oi_1 _7458_ (.A1(net1250),
    .A2(net1203),
    .Y(_0506_),
    .B1(_3063_));
 sg13g2_nor2_1 _7459_ (.A(net1034),
    .B(net1202),
    .Y(_3064_));
 sg13g2_a21oi_1 _7460_ (.A1(net1246),
    .A2(net1202),
    .Y(_0507_),
    .B1(_3064_));
 sg13g2_nor2_1 _7461_ (.A(net807),
    .B(net1202),
    .Y(_3065_));
 sg13g2_a21oi_1 _7462_ (.A1(net1245),
    .A2(net1202),
    .Y(_0508_),
    .B1(_3065_));
 sg13g2_nor2_1 _7463_ (.A(net829),
    .B(net1203),
    .Y(_3066_));
 sg13g2_a21oi_1 _7464_ (.A1(net1222),
    .A2(net1203),
    .Y(_0509_),
    .B1(_3066_));
 sg13g2_nor2_1 _7465_ (.A(net921),
    .B(net1202),
    .Y(_3067_));
 sg13g2_a21oi_1 _7466_ (.A1(_2772_),
    .A2(net1202),
    .Y(_0510_),
    .B1(_3067_));
 sg13g2_nor2_1 _7467_ (.A(_1991_),
    .B(_3043_),
    .Y(_3068_));
 sg13g2_nor2_1 _7468_ (.A(net920),
    .B(net1183),
    .Y(_3069_));
 sg13g2_a21oi_1 _7469_ (.A1(net1255),
    .A2(net1183),
    .Y(_0511_),
    .B1(_3069_));
 sg13g2_nor2_1 _7470_ (.A(net862),
    .B(net1184),
    .Y(_3070_));
 sg13g2_a21oi_1 _7471_ (.A1(net1254),
    .A2(net1184),
    .Y(_0512_),
    .B1(_3070_));
 sg13g2_mux2_1 _7472_ (.A0(net884),
    .A1(net1252),
    .S(net1184),
    .X(_0513_));
 sg13g2_nor2_1 _7473_ (.A(net815),
    .B(net1184),
    .Y(_3071_));
 sg13g2_a21oi_1 _7474_ (.A1(net1250),
    .A2(net1184),
    .Y(_0514_),
    .B1(_3071_));
 sg13g2_nor2_1 _7475_ (.A(net781),
    .B(net1183),
    .Y(_3072_));
 sg13g2_a21oi_1 _7476_ (.A1(net1246),
    .A2(net1183),
    .Y(_0515_),
    .B1(_3072_));
 sg13g2_nor2_1 _7477_ (.A(net989),
    .B(net1183),
    .Y(_3073_));
 sg13g2_a21oi_1 _7478_ (.A1(net1245),
    .A2(net1183),
    .Y(_0516_),
    .B1(_3073_));
 sg13g2_nor2_1 _7479_ (.A(net962),
    .B(net1184),
    .Y(_3074_));
 sg13g2_a21oi_1 _7480_ (.A1(net1222),
    .A2(net1184),
    .Y(_0517_),
    .B1(_3074_));
 sg13g2_nor2_1 _7481_ (.A(net710),
    .B(net1183),
    .Y(_3075_));
 sg13g2_a21oi_1 _7482_ (.A1(net1242),
    .A2(net1183),
    .Y(_0518_),
    .B1(_3075_));
 sg13g2_nor3_2 _7483_ (.A(\scl_fifo1.n6229_o[2] ),
    .B(\scl_fifo1.n6229_o[3] ),
    .C(_1990_),
    .Y(_3076_));
 sg13g2_nor2_1 _7484_ (.A(net997),
    .B(net1200),
    .Y(_3077_));
 sg13g2_a21oi_1 _7485_ (.A1(net1255),
    .A2(net1200),
    .Y(_0519_),
    .B1(_3077_));
 sg13g2_nor2_1 _7486_ (.A(net766),
    .B(net1201),
    .Y(_3078_));
 sg13g2_a21oi_1 _7487_ (.A1(net1254),
    .A2(net1201),
    .Y(_0520_),
    .B1(_3078_));
 sg13g2_mux2_1 _7488_ (.A0(net812),
    .A1(net1252),
    .S(net1201),
    .X(_0521_));
 sg13g2_nor2_1 _7489_ (.A(net758),
    .B(net1201),
    .Y(_3079_));
 sg13g2_a21oi_1 _7490_ (.A1(net1250),
    .A2(net1201),
    .Y(_0522_),
    .B1(_3079_));
 sg13g2_nor2_1 _7491_ (.A(net764),
    .B(net1200),
    .Y(_3080_));
 sg13g2_a21oi_1 _7492_ (.A1(net1247),
    .A2(net1200),
    .Y(_0523_),
    .B1(_3080_));
 sg13g2_nor2_1 _7493_ (.A(net1008),
    .B(net1200),
    .Y(_3081_));
 sg13g2_a21oi_1 _7494_ (.A1(net1245),
    .A2(net1200),
    .Y(_0524_),
    .B1(_3081_));
 sg13g2_nor2_1 _7495_ (.A(net948),
    .B(net1201),
    .Y(_3082_));
 sg13g2_a21oi_1 _7496_ (.A1(net1222),
    .A2(net1201),
    .Y(_0525_),
    .B1(_3082_));
 sg13g2_nor2_1 _7497_ (.A(net913),
    .B(net1200),
    .Y(_3083_));
 sg13g2_a21oi_1 _7498_ (.A1(net1242),
    .A2(net1200),
    .Y(_0526_),
    .B1(_3083_));
 sg13g2_nor4_2 _7499_ (.A(\scl_fifo1.n6229_o[2] ),
    .B(\scl_fifo1.n6229_o[3] ),
    .C(net1258),
    .Y(_3084_),
    .D(_2984_));
 sg13g2_nor2_1 _7500_ (.A(net778),
    .B(net1198),
    .Y(_3085_));
 sg13g2_a21oi_1 _7501_ (.A1(net1255),
    .A2(net1198),
    .Y(_0527_),
    .B1(_3085_));
 sg13g2_nor2_1 _7502_ (.A(net808),
    .B(net1199),
    .Y(_3086_));
 sg13g2_a21oi_1 _7503_ (.A1(net1254),
    .A2(net1199),
    .Y(_0528_),
    .B1(_3086_));
 sg13g2_mux2_1 _7504_ (.A0(net864),
    .A1(net1252),
    .S(net1199),
    .X(_0529_));
 sg13g2_nor2_1 _7505_ (.A(net908),
    .B(net1199),
    .Y(_3087_));
 sg13g2_a21oi_1 _7506_ (.A1(net1250),
    .A2(net1199),
    .Y(_0530_),
    .B1(_3087_));
 sg13g2_nor2_1 _7507_ (.A(net977),
    .B(net1198),
    .Y(_3088_));
 sg13g2_a21oi_1 _7508_ (.A1(net1247),
    .A2(net1198),
    .Y(_0531_),
    .B1(_3088_));
 sg13g2_nor2_1 _7509_ (.A(net787),
    .B(net1198),
    .Y(_3089_));
 sg13g2_a21oi_1 _7510_ (.A1(net1245),
    .A2(net1198),
    .Y(_0532_),
    .B1(_3089_));
 sg13g2_nor2_1 _7511_ (.A(net969),
    .B(net1199),
    .Y(_3090_));
 sg13g2_a21oi_1 _7512_ (.A1(net1222),
    .A2(net1199),
    .Y(_0533_),
    .B1(_3090_));
 sg13g2_nor2_1 _7513_ (.A(net933),
    .B(net1198),
    .Y(_3091_));
 sg13g2_a21oi_1 _7514_ (.A1(net1242),
    .A2(net1198),
    .Y(_0534_),
    .B1(_3091_));
 sg13g2_nor4_2 _7515_ (.A(\scl_fifo1.n6229_o[2] ),
    .B(\scl_fifo1.n6229_o[3] ),
    .C(net1258),
    .Y(_3092_),
    .D(_2993_));
 sg13g2_nor2_1 _7516_ (.A(net846),
    .B(net1196),
    .Y(_3093_));
 sg13g2_a21oi_1 _7517_ (.A1(net1255),
    .A2(net1196),
    .Y(_0535_),
    .B1(_3093_));
 sg13g2_nor2_1 _7518_ (.A(net802),
    .B(net1197),
    .Y(_3094_));
 sg13g2_a21oi_1 _7519_ (.A1(net1254),
    .A2(net1197),
    .Y(_0536_),
    .B1(_3094_));
 sg13g2_mux2_1 _7520_ (.A0(net895),
    .A1(net1252),
    .S(net1197),
    .X(_0537_));
 sg13g2_nor2_1 _7521_ (.A(net871),
    .B(net1197),
    .Y(_3095_));
 sg13g2_a21oi_1 _7522_ (.A1(net1250),
    .A2(net1196),
    .Y(_0538_),
    .B1(_3095_));
 sg13g2_nor2_1 _7523_ (.A(net999),
    .B(net1196),
    .Y(_3096_));
 sg13g2_a21oi_1 _7524_ (.A1(net1247),
    .A2(net1196),
    .Y(_0539_),
    .B1(_3096_));
 sg13g2_nor2_1 _7525_ (.A(net887),
    .B(net1197),
    .Y(_3097_));
 sg13g2_a21oi_1 _7526_ (.A1(net1245),
    .A2(net1196),
    .Y(_0540_),
    .B1(_3097_));
 sg13g2_nor2_1 _7527_ (.A(net782),
    .B(net1197),
    .Y(_3098_));
 sg13g2_a21oi_1 _7528_ (.A1(net1222),
    .A2(net1197),
    .Y(_0541_),
    .B1(_3098_));
 sg13g2_nor2_1 _7529_ (.A(net942),
    .B(net1196),
    .Y(_3099_));
 sg13g2_a21oi_1 _7530_ (.A1(net1242),
    .A2(net1196),
    .Y(_0542_),
    .B1(_3099_));
 sg13g2_nand2_1 _7531_ (.Y(_3100_),
    .A(_1850_),
    .B(_2880_));
 sg13g2_nand2_1 _7532_ (.Y(_3101_),
    .A(net574),
    .B(net1334));
 sg13g2_o21ai_1 _7533_ (.B1(_3101_),
    .Y(_0543_),
    .A1(net1452),
    .A2(net1335));
 sg13g2_nand2_1 _7534_ (.Y(_3102_),
    .A(net575),
    .B(net1334));
 sg13g2_o21ai_1 _7535_ (.B1(_3102_),
    .Y(_0544_),
    .A1(net1455),
    .A2(net1334));
 sg13g2_mux2_1 _7536_ (.A0(net1474),
    .A1(net936),
    .S(net1335),
    .X(_0545_));
 sg13g2_nand2_1 _7537_ (.Y(_3103_),
    .A(net591),
    .B(net1334));
 sg13g2_o21ai_1 _7538_ (.B1(_3103_),
    .Y(_0546_),
    .A1(net1458),
    .A2(net1334));
 sg13g2_mux2_1 _7539_ (.A0(net1471),
    .A1(net976),
    .S(net1334),
    .X(_0547_));
 sg13g2_mux2_1 _7540_ (.A0(net1468),
    .A1(net963),
    .S(net1334),
    .X(_0548_));
 sg13g2_mux2_1 _7541_ (.A0(net1465),
    .A1(net1049),
    .S(net1335),
    .X(_0549_));
 sg13g2_mux2_1 _7542_ (.A0(net1462),
    .A1(net947),
    .S(net1334),
    .X(_0550_));
 sg13g2_mux2_1 _7543_ (.A0(net1090),
    .A1(net779),
    .S(net1398),
    .X(_0551_));
 sg13g2_a21o_1 _7544_ (.A2(net1386),
    .A1(net1023),
    .B1(net1670),
    .X(_3104_));
 sg13g2_and2_1 _7545_ (.A(_0795_),
    .B(_3104_),
    .X(_0552_));
 sg13g2_mux2_1 _7546_ (.A0(net1090),
    .A1(net545),
    .S(net1620),
    .X(_0553_));
 sg13g2_nor3_1 _7547_ (.A(net1090),
    .B(net1437),
    .C(net1398),
    .Y(_3105_));
 sg13g2_a21o_1 _7548_ (.A2(_0784_),
    .A1(net542),
    .B1(_3105_),
    .X(_0554_));
 sg13g2_nand2_2 _7549_ (.Y(_3106_),
    .A(s_m_phy_tx_valid_2),
    .B(net1392));
 sg13g2_nand2_1 _7550_ (.Y(_3107_),
    .A(net835),
    .B(net1393));
 sg13g2_o21ai_1 _7551_ (.B1(_3107_),
    .Y(_0555_),
    .A1(net984),
    .A2(_3106_));
 sg13g2_a22oi_1 _7552_ (.Y(_3108_),
    .B1(_0793_),
    .B2(net628),
    .A2(net1398),
    .A1(\usbfunction0.scl_usbgpiophy0.scl_decodenrzi0.scl_counter0.n7944_q[0] ));
 sg13g2_inv_1 _7553_ (.Y(_0556_),
    .A(net629));
 sg13g2_nor2_1 _7554_ (.A(net628),
    .B(net1398),
    .Y(_3109_));
 sg13g2_nor2_1 _7555_ (.A(net1030),
    .B(_3109_),
    .Y(_3110_));
 sg13g2_nand2_1 _7556_ (.Y(_3111_),
    .A(net1030),
    .B(_3109_));
 sg13g2_o21ai_1 _7557_ (.B1(_3111_),
    .Y(_3112_),
    .A1(net1398),
    .A2(_0792_));
 sg13g2_nor2_1 _7558_ (.A(_3110_),
    .B(_3112_),
    .Y(_0557_));
 sg13g2_nor2_1 _7559_ (.A(_0156_),
    .B(_0785_),
    .Y(_3113_));
 sg13g2_a21oi_1 _7560_ (.A1(_0044_),
    .A2(_3111_),
    .Y(_3114_),
    .B1(_3113_));
 sg13g2_a22oi_1 _7561_ (.Y(_3115_),
    .B1(_0793_),
    .B2(_3114_),
    .A2(net1398),
    .A1(net601));
 sg13g2_inv_1 _7562_ (.Y(_0558_),
    .A(net602));
 sg13g2_nand2_1 _7563_ (.Y(_3116_),
    .A(net723),
    .B(_1038_));
 sg13g2_nand2_1 _7564_ (.Y(_3117_),
    .A(\usbfunction0.s_m_descdata[0] ),
    .B(net1395));
 sg13g2_nand3_1 _7565_ (.B(_1029_),
    .C(_3117_),
    .A(net1367),
    .Y(_3118_));
 sg13g2_o21ai_1 _7566_ (.B1(_3118_),
    .Y(_3119_),
    .A1(\s_m_peekdata_data_2[0] ),
    .A2(net1366));
 sg13g2_o21ai_1 _7567_ (.B1(_3116_),
    .Y(_0559_),
    .A1(net1393),
    .A2(_3119_));
 sg13g2_nand2_1 _7568_ (.Y(_3120_),
    .A(net620),
    .B(net1393));
 sg13g2_nand2b_1 _7569_ (.Y(_3121_),
    .B(net1395),
    .A_N(\usbfunction0.s_m_descdata[1] ));
 sg13g2_o21ai_1 _7570_ (.B1(_3121_),
    .Y(_3122_),
    .A1(\s_m_peekdata_data_2[1] ),
    .A2(net1366));
 sg13g2_o21ai_1 _7571_ (.B1(_3120_),
    .Y(_0560_),
    .A1(_3106_),
    .A2(_3122_));
 sg13g2_nand2_1 _7572_ (.Y(_3123_),
    .A(net633),
    .B(net1393));
 sg13g2_nand3_1 _7573_ (.B(\usbfunction0.n2635_q[0] ),
    .C(\usbfunction0.n2635_q[1] ),
    .A(\usbfunction0.n2636_q ),
    .Y(_3124_));
 sg13g2_o21ai_1 _7574_ (.B1(net1367),
    .Y(_3125_),
    .A1(_1031_),
    .A2(_3124_));
 sg13g2_a21oi_1 _7575_ (.A1(\usbfunction0.s_m_descdata[2] ),
    .A2(net1395),
    .Y(_3126_),
    .B1(_3125_));
 sg13g2_o21ai_1 _7576_ (.B1(_1039_),
    .Y(_3127_),
    .A1(\s_m_peekdata_data_2[2] ),
    .A2(net1366));
 sg13g2_o21ai_1 _7577_ (.B1(_3123_),
    .Y(_0561_),
    .A1(_3126_),
    .A2(_3127_));
 sg13g2_nand2_1 _7578_ (.Y(_3128_),
    .A(\usbfunction0.n1630_o[15] ),
    .B(\usbfunction0.n2257_o[15] ));
 sg13g2_a22oi_1 _7579_ (.Y(_3129_),
    .B1(\usbfunction0.n2257_o[8] ),
    .B2(\usbfunction0.n1630_o[8] ),
    .A2(\usbfunction0.n2257_o[2] ),
    .A1(\usbfunction0.n1630_o[2] ));
 sg13g2_a22oi_1 _7580_ (.Y(_3130_),
    .B1(\usbfunction0.n2257_o[12] ),
    .B2(\usbfunction0.n1630_o[12] ),
    .A2(\usbfunction0.n2257_o[3] ),
    .A1(\usbfunction0.n1630_o[3] ));
 sg13g2_a22oi_1 _7581_ (.Y(_3131_),
    .B1(\usbfunction0.n2257_o[6] ),
    .B2(\usbfunction0.n1630_o[6] ),
    .A2(\usbfunction0.n2257_o[1] ),
    .A1(\usbfunction0.n1630_o[1] ));
 sg13g2_nand3_1 _7582_ (.B(_3130_),
    .C(_3131_),
    .A(_3129_),
    .Y(_3132_));
 sg13g2_a221oi_1 _7583_ (.B2(\usbfunction0.n1630_o[9] ),
    .C1(_3132_),
    .B1(\usbfunction0.n2257_o[9] ),
    .A1(\usbfunction0.n1630_o[7] ),
    .Y(_3133_),
    .A2(\usbfunction0.n2257_o[7] ));
 sg13g2_a22oi_1 _7584_ (.Y(_3134_),
    .B1(\usbfunction0.n2257_o[14] ),
    .B2(\usbfunction0.n1630_o[14] ),
    .A2(\usbfunction0.n2257_o[13] ),
    .A1(\usbfunction0.n1630_o[13] ));
 sg13g2_a22oi_1 _7585_ (.Y(_3135_),
    .B1(\usbfunction0.n2257_o[11] ),
    .B2(\usbfunction0.n1630_o[11] ),
    .A2(\usbfunction0.n2257_o[4] ),
    .A1(\usbfunction0.n1630_o[4] ));
 sg13g2_a22oi_1 _7586_ (.Y(_3136_),
    .B1(\usbfunction0.n2257_o[10] ),
    .B2(\usbfunction0.n1630_o[10] ),
    .A2(\usbfunction0.n2257_o[5] ),
    .A1(\usbfunction0.n1630_o[5] ));
 sg13g2_nand4_1 _7587_ (.B(_3134_),
    .C(_3135_),
    .A(_3128_),
    .Y(_3137_),
    .D(_3136_));
 sg13g2_a21oi_1 _7588_ (.A1(\usbfunction0.n1630_o[0] ),
    .A2(\usbfunction0.n2254_o ),
    .Y(_3138_),
    .B1(_3137_));
 sg13g2_a21o_2 _7589_ (.A2(_3138_),
    .A1(_3133_),
    .B1(_1029_),
    .X(_3139_));
 sg13g2_nand2b_1 _7590_ (.Y(_3140_),
    .B(\usbfunction0.n2635_q[1] ),
    .A_N(\usbfunction0.n2635_q[0] ));
 sg13g2_nor2_1 _7591_ (.A(_0117_),
    .B(_3140_),
    .Y(_3141_));
 sg13g2_a221oi_1 _7592_ (.B2(_3141_),
    .C1(_3125_),
    .B1(_1030_),
    .A1(\usbfunction0.s_m_descdata[3] ),
    .Y(_3142_),
    .A2(net1394));
 sg13g2_o21ai_1 _7593_ (.B1(_1039_),
    .Y(_3143_),
    .A1(\s_m_peekdata_data_2[3] ),
    .A2(net1365));
 sg13g2_a21oi_1 _7594_ (.A1(_3139_),
    .A2(_3142_),
    .Y(_3144_),
    .B1(_3143_));
 sg13g2_a21o_1 _7595_ (.A2(_1038_),
    .A1(net1009),
    .B1(_3144_),
    .X(_0562_));
 sg13g2_a22oi_1 _7596_ (.Y(_3145_),
    .B1(_1030_),
    .B2(\usbfunction0.n2636_q ),
    .A2(net1394),
    .A1(\usbfunction0.s_m_descdata[4] ));
 sg13g2_o21ai_1 _7597_ (.B1(net1392),
    .Y(_3146_),
    .A1(\s_m_peekdata_data_2[4] ),
    .A2(net1365));
 sg13g2_a21oi_1 _7598_ (.A1(net1365),
    .A2(_3145_),
    .Y(_3147_),
    .B1(_3146_));
 sg13g2_a21o_1 _7599_ (.A2(net1393),
    .A1(net902),
    .B1(_3147_),
    .X(_0563_));
 sg13g2_nand2_1 _7600_ (.Y(_3148_),
    .A(\usbfunction0.s_m_descdata[5] ),
    .B(net1395));
 sg13g2_o21ai_1 _7601_ (.B1(net1392),
    .Y(_3149_),
    .A1(\s_m_peekdata_data_2[5] ),
    .A2(net1365));
 sg13g2_a21oi_1 _7602_ (.A1(net1366),
    .A2(_3148_),
    .Y(_3150_),
    .B1(_3149_));
 sg13g2_a21o_1 _7603_ (.A2(net1393),
    .A1(net1076),
    .B1(_3150_),
    .X(_0564_));
 sg13g2_nand2_1 _7604_ (.Y(_3151_),
    .A(net617),
    .B(net1393));
 sg13g2_nand4_1 _7605_ (.B(\usbfunction0.n2635_q[1] ),
    .C(net1367),
    .A(\usbfunction0.n2635_q[0] ),
    .Y(_3152_),
    .D(_1030_));
 sg13g2_nand2b_1 _7606_ (.Y(_3153_),
    .B(net1395),
    .A_N(\usbfunction0.s_m_descdata[6] ));
 sg13g2_o21ai_1 _7607_ (.B1(_3153_),
    .Y(_3154_),
    .A1(\s_m_peekdata_data_2[6] ),
    .A2(net1365));
 sg13g2_nand2b_1 _7608_ (.Y(_3155_),
    .B(_3152_),
    .A_N(_3154_));
 sg13g2_o21ai_1 _7609_ (.B1(_3151_),
    .Y(_0565_),
    .A1(_3106_),
    .A2(_3155_));
 sg13g2_nand3b_1 _7610_ (.B(_3124_),
    .C(_3140_),
    .Y(_3156_),
    .A_N(_0117_));
 sg13g2_a21oi_1 _7611_ (.A1(_1029_),
    .A2(_3156_),
    .Y(_3157_),
    .B1(net1394));
 sg13g2_a22oi_1 _7612_ (.Y(_3158_),
    .B1(_3139_),
    .B2(_3157_),
    .A2(net1394),
    .A1(\usbfunction0.s_m_descdata[7] ));
 sg13g2_o21ai_1 _7613_ (.B1(net1392),
    .Y(_3159_),
    .A1(\s_m_peekdata_data_2[7] ),
    .A2(net1365));
 sg13g2_a21o_1 _7614_ (.A2(_3158_),
    .A1(net1365),
    .B1(_3159_),
    .X(_3160_));
 sg13g2_o21ai_1 _7615_ (.B1(_3160_),
    .Y(_0566_),
    .A1(_0714_),
    .A2(net1392));
 sg13g2_nand2b_1 _7616_ (.Y(_3161_),
    .B(net668),
    .A_N(_0782_));
 sg13g2_nand2b_1 _7617_ (.Y(_3162_),
    .B(_0782_),
    .A_N(_2182_));
 sg13g2_a21oi_1 _7618_ (.A1(_3161_),
    .A2(_3162_),
    .Y(_0567_),
    .B1(_2554_));
 sg13g2_a21oi_1 _7619_ (.A1(_0749_),
    .A2(net1393),
    .Y(_0568_),
    .B1(_1040_));
 sg13g2_nor3_2 _7620_ (.A(\scl_bitbangengine0.n5920_q[9] ),
    .B(\scl_bitbangengine0.n5920_q[8] ),
    .C(_2641_),
    .Y(_3163_));
 sg13g2_o21ai_1 _7621_ (.B1(net1726),
    .Y(_3164_),
    .A1(\scl_bitbangengine0.n5920_q[8] ),
    .A2(_2641_));
 sg13g2_nand2b_1 _7622_ (.Y(_3165_),
    .B(_3164_),
    .A_N(_3163_));
 sg13g2_a22oi_1 _7623_ (.Y(_3166_),
    .B1(_3165_),
    .B2(_2594_),
    .A2(_2630_),
    .A1(net1412));
 sg13g2_nor2_1 _7624_ (.A(net1726),
    .B(_2595_),
    .Y(_3167_));
 sg13g2_a21oi_1 _7625_ (.A1(_2595_),
    .A2(_3166_),
    .Y(_0569_),
    .B1(_3167_));
 sg13g2_nor2_1 _7626_ (.A(net1103),
    .B(_2595_),
    .Y(_3168_));
 sg13g2_nand2_1 _7627_ (.Y(_3169_),
    .A(_0142_),
    .B(_3163_));
 sg13g2_xnor2_1 _7628_ (.Y(_3170_),
    .A(_0142_),
    .B(_3163_));
 sg13g2_a22oi_1 _7629_ (.Y(_3171_),
    .B1(_3170_),
    .B2(_2594_),
    .A2(_2635_),
    .A1(net1412));
 sg13g2_a21oi_1 _7630_ (.A1(_2595_),
    .A2(_3171_),
    .Y(_0570_),
    .B1(_3168_));
 sg13g2_nand2_1 _7631_ (.Y(_3172_),
    .A(net605),
    .B(net1353));
 sg13g2_xnor2_1 _7632_ (.Y(_3173_),
    .A(_2962_),
    .B(_2964_));
 sg13g2_o21ai_1 _7633_ (.B1(_3172_),
    .Y(_0571_),
    .A1(net1352),
    .A2(_3173_));
 sg13g2_a22oi_1 _7634_ (.Y(_0572_),
    .B1(_2972_),
    .B2(_0750_),
    .A2(net1351),
    .A1(_0712_));
 sg13g2_a22oi_1 _7635_ (.Y(_0573_),
    .B1(net1336),
    .B2(_0751_),
    .A2(net1354),
    .A1(_0750_));
 sg13g2_a22oi_1 _7636_ (.Y(_0574_),
    .B1(net1336),
    .B2(_0752_),
    .A2(net1354),
    .A1(_0751_));
 sg13g2_a22oi_1 _7637_ (.Y(_0575_),
    .B1(net1336),
    .B2(_0753_),
    .A2(net1354),
    .A1(_0752_));
 sg13g2_nor3_1 _7638_ (.A(net1044),
    .B(_2176_),
    .C(net1353),
    .Y(_3174_));
 sg13g2_a21oi_1 _7639_ (.A1(_0753_),
    .A2(net1351),
    .Y(_0576_),
    .B1(_3174_));
 sg13g2_a22oi_1 _7640_ (.Y(_0577_),
    .B1(net1336),
    .B2(_0755_),
    .A2(net1351),
    .A1(_0754_));
 sg13g2_a22oi_1 _7641_ (.Y(_0578_),
    .B1(net1336),
    .B2(_0756_),
    .A2(net1351),
    .A1(_0755_));
 sg13g2_a22oi_1 _7642_ (.Y(_0579_),
    .B1(net1336),
    .B2(_0757_),
    .A2(net1351),
    .A1(_0756_));
 sg13g2_a22oi_1 _7643_ (.Y(_0580_),
    .B1(net1336),
    .B2(_0758_),
    .A2(net1351),
    .A1(_0757_));
 sg13g2_a22oi_1 _7644_ (.Y(_0581_),
    .B1(net1336),
    .B2(_0715_),
    .A2(net1351),
    .A1(_0758_));
 sg13g2_a22oi_1 _7645_ (.Y(_0582_),
    .B1(_2972_),
    .B2(_0759_),
    .A2(net1351),
    .A1(_0715_));
 sg13g2_a22oi_1 _7646_ (.Y(_0583_),
    .B1(_2972_),
    .B2(_0716_),
    .A2(net1352),
    .A1(_0759_));
 sg13g2_nand2_1 _7647_ (.Y(_3175_),
    .A(net736),
    .B(net1352));
 sg13g2_o21ai_1 _7648_ (.B1(_3175_),
    .Y(_0584_),
    .A1(net1352),
    .A2(_2971_));
 sg13g2_a21oi_1 _7649_ (.A1(_0717_),
    .A2(net1352),
    .Y(_0585_),
    .B1(_2973_));
 sg13g2_nand2_1 _7650_ (.Y(_3176_),
    .A(net610),
    .B(net1352));
 sg13g2_o21ai_1 _7651_ (.B1(_3176_),
    .Y(_0586_),
    .A1(net1352),
    .A2(_2962_));
 sg13g2_nor3_1 _7652_ (.A(net1903),
    .B(_1328_),
    .C(_1952_),
    .Y(_3177_));
 sg13g2_nor2_1 _7653_ (.A(net640),
    .B(net1408),
    .Y(_3178_));
 sg13g2_a21oi_1 _7654_ (.A1(_2609_),
    .A2(net1409),
    .Y(_0587_),
    .B1(_3178_));
 sg13g2_mux2_1 _7655_ (.A0(net1711),
    .A1(_2617_),
    .S(net1408),
    .X(_0588_));
 sg13g2_mux2_1 _7656_ (.A0(net831),
    .A1(_2625_),
    .S(net1408),
    .X(_0589_));
 sg13g2_nor2_1 _7657_ (.A(net1580),
    .B(net1408),
    .Y(_3179_));
 sg13g2_a21oi_1 _7658_ (.A1(_2607_),
    .A2(net1408),
    .Y(_0590_),
    .B1(_3179_));
 sg13g2_mux2_1 _7659_ (.A0(net1761),
    .A1(_2614_),
    .S(net1408),
    .X(_0591_));
 sg13g2_mux2_1 _7660_ (.A0(net1587),
    .A1(_2623_),
    .S(net1408),
    .X(_0592_));
 sg13g2_mux2_1 _7661_ (.A0(net819),
    .A1(_2630_),
    .S(net1408),
    .X(_0593_));
 sg13g2_nor2_1 _7662_ (.A(net1653),
    .B(net1409),
    .Y(_3180_));
 sg13g2_a21oi_1 _7663_ (.A1(_2636_),
    .A2(net1409),
    .Y(_0594_),
    .B1(_3180_));
 sg13g2_nor2_2 _7664_ (.A(_0084_),
    .B(_1327_),
    .Y(_3181_));
 sg13g2_nor2_1 _7665_ (.A(_1077_),
    .B(net1407),
    .Y(_3182_));
 sg13g2_nor2b_1 _7666_ (.A(_1197_),
    .B_N(net1372),
    .Y(_3183_));
 sg13g2_xnor2_1 _7667_ (.Y(_3184_),
    .A(net1151),
    .B(_3169_));
 sg13g2_a221oi_1 _7668_ (.B2(_3184_),
    .C1(net1333),
    .B1(_3182_),
    .A1(_2609_),
    .Y(_3185_),
    .A2(net1407));
 sg13g2_a21oi_1 _7669_ (.A1(_0738_),
    .A2(net1333),
    .Y(_0595_),
    .B1(_3185_));
 sg13g2_nand3_1 _7670_ (.B(_1185_),
    .C(_2600_),
    .A(_1183_),
    .Y(_3186_));
 sg13g2_xnor2_1 _7671_ (.Y(_3187_),
    .A(net1766),
    .B(_3186_));
 sg13g2_a221oi_1 _7672_ (.B2(_3187_),
    .C1(net1332),
    .B1(net1372),
    .A1(_2617_),
    .Y(_3188_),
    .A2(net1407));
 sg13g2_a21oi_1 _7673_ (.A1(_0739_),
    .A2(net1331),
    .Y(_0596_),
    .B1(_3188_));
 sg13g2_nor3_2 _7674_ (.A(\scl_bitbangengine0.n5920_q[12] ),
    .B(\scl_bitbangengine0.n5920_q[13] ),
    .C(_3186_),
    .Y(_3189_));
 sg13g2_o21ai_1 _7675_ (.B1(net1584),
    .Y(_3190_),
    .A1(\scl_bitbangengine0.n5920_q[12] ),
    .A2(_3186_));
 sg13g2_nand2b_1 _7676_ (.Y(_3191_),
    .B(_3190_),
    .A_N(_3189_));
 sg13g2_a221oi_1 _7677_ (.B2(_3191_),
    .C1(net1332),
    .B1(net1372),
    .A1(_2625_),
    .Y(_3192_),
    .A2(net1407));
 sg13g2_a21oi_1 _7678_ (.A1(_0740_),
    .A2(net1331),
    .Y(_0597_),
    .B1(_3192_));
 sg13g2_nand2_1 _7679_ (.Y(_3193_),
    .A(_0143_),
    .B(_3189_));
 sg13g2_xnor2_1 _7680_ (.Y(_3194_),
    .A(_0143_),
    .B(_3189_));
 sg13g2_a221oi_1 _7681_ (.B2(_3194_),
    .C1(net1331),
    .B1(net1372),
    .A1(_2606_),
    .Y(_3195_),
    .A2(net1407));
 sg13g2_a21oi_1 _7682_ (.A1(_0741_),
    .A2(net1331),
    .Y(_0598_),
    .B1(_3195_));
 sg13g2_xnor2_1 _7683_ (.Y(_3196_),
    .A(net1571),
    .B(_3193_));
 sg13g2_a221oi_1 _7684_ (.B2(_3196_),
    .C1(net1332),
    .B1(net1372),
    .A1(_2614_),
    .Y(_3197_),
    .A2(net1407));
 sg13g2_a21oi_1 _7685_ (.A1(_0742_),
    .A2(net1331),
    .Y(_0599_),
    .B1(_3197_));
 sg13g2_nor3_2 _7686_ (.A(\scl_bitbangengine0.n5920_q[16] ),
    .B(_1186_),
    .C(_3186_),
    .Y(_3198_));
 sg13g2_o21ai_1 _7687_ (.B1(net1577),
    .Y(_3199_),
    .A1(_1186_),
    .A2(_3186_));
 sg13g2_nand2b_1 _7688_ (.Y(_3200_),
    .B(_3199_),
    .A_N(_3198_));
 sg13g2_a221oi_1 _7689_ (.B2(_3200_),
    .C1(net1331),
    .B1(net1372),
    .A1(_2623_),
    .Y(_3201_),
    .A2(net1407));
 sg13g2_a21oi_1 _7690_ (.A1(_0743_),
    .A2(net1331),
    .Y(_0600_),
    .B1(_3201_));
 sg13g2_and2_1 _7691_ (.A(_0744_),
    .B(_3198_),
    .X(_3202_));
 sg13g2_xnor2_1 _7692_ (.Y(_3203_),
    .A(_0744_),
    .B(_3198_));
 sg13g2_a221oi_1 _7693_ (.B2(_3203_),
    .C1(net1331),
    .B1(net1372),
    .A1(_2630_),
    .Y(_3204_),
    .A2(net1407));
 sg13g2_a21oi_1 _7694_ (.A1(_0744_),
    .A2(net1332),
    .Y(_0601_),
    .B1(_3204_));
 sg13g2_nand2_1 _7695_ (.Y(_3205_),
    .A(_0144_),
    .B(_3202_));
 sg13g2_xnor2_1 _7696_ (.Y(_3206_),
    .A(_0144_),
    .B(_3202_));
 sg13g2_a221oi_1 _7697_ (.B2(_3206_),
    .C1(net1332),
    .B1(net1372),
    .A1(_2635_),
    .Y(_3207_),
    .A2(_3181_));
 sg13g2_a21oi_1 _7698_ (.A1(_0746_),
    .A2(net1333),
    .Y(_0602_),
    .B1(_3207_));
 sg13g2_xnor2_1 _7699_ (.Y(_3208_),
    .A(net1054),
    .B(_3205_));
 sg13g2_a221oi_1 _7700_ (.B2(_3208_),
    .C1(net1333),
    .B1(_3182_),
    .A1(_2634_),
    .Y(_3209_),
    .A2(_3181_));
 sg13g2_a21oi_1 _7701_ (.A1(_0745_),
    .A2(net1333),
    .Y(_0603_),
    .B1(_3209_));
 sg13g2_nor2b_1 _7702_ (.A(net1758),
    .B_N(_2975_),
    .Y(_3210_));
 sg13g2_nand4_1 _7703_ (.B(_0779_),
    .C(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7508_o ),
    .A(_0777_),
    .Y(_3211_),
    .D(_3210_));
 sg13g2_nand3_1 _7704_ (.B(_2523_),
    .C(_2549_),
    .A(_2171_),
    .Y(_3212_));
 sg13g2_nand2_1 _7705_ (.Y(_3213_),
    .A(_3211_),
    .B(_3212_));
 sg13g2_nand3_1 _7706_ (.B(_3211_),
    .C(_3212_),
    .A(net1762),
    .Y(_3214_));
 sg13g2_o21ai_1 _7707_ (.B1(_3214_),
    .Y(_0604_),
    .A1(_2549_),
    .A2(_3211_));
 sg13g2_a21oi_1 _7708_ (.A1(_2549_),
    .A2(_3213_),
    .Y(_3215_),
    .B1(net1820));
 sg13g2_nor3_1 _7709_ (.A(_0780_),
    .B(_1034_),
    .C(net1758),
    .Y(_3216_));
 sg13g2_nor2_1 _7710_ (.A(net1821),
    .B(_3216_),
    .Y(_0605_));
 sg13g2_nor2b_1 _7711_ (.A(\usbfunction0.n2313_o[3] ),
    .B_N(\usbfunction0.n2631_q ),
    .Y(_3217_));
 sg13g2_nand2b_1 _7712_ (.Y(_3218_),
    .B(\usbfunction0.n2631_q ),
    .A_N(\usbfunction0.n2313_o[3] ));
 sg13g2_nor2_1 _7713_ (.A(net767),
    .B(net1441),
    .Y(_3219_));
 sg13g2_a21oi_1 _7714_ (.A1(_0723_),
    .A2(net1441),
    .Y(_0606_),
    .B1(_3219_));
 sg13g2_mux2_1 _7715_ (.A0(net1172),
    .A1(\s_m_packetdata_2_rewired[1] ),
    .S(net1441),
    .X(_0607_));
 sg13g2_mux2_1 _7716_ (.A0(\s_m_packetdata_2_rewired[10] ),
    .A1(net1578),
    .S(net1441),
    .X(_0608_));
 sg13g2_mux2_1 _7717_ (.A0(\s_m_packetdata_2_rewired[11] ),
    .A1(net1675),
    .S(net1442),
    .X(_0609_));
 sg13g2_mux2_1 _7718_ (.A0(\s_m_packetdata_2_rewired[12] ),
    .A1(net1632),
    .S(net1442),
    .X(_0610_));
 sg13g2_mux2_1 _7719_ (.A0(net1696),
    .A1(net1702),
    .S(net1440),
    .X(_0611_));
 sg13g2_mux2_1 _7720_ (.A0(net1161),
    .A1(\s_m_packetdata_2_rewired[6] ),
    .S(net1440),
    .X(_0612_));
 sg13g2_mux2_1 _7721_ (.A0(\s_m_packetdata_2_rewired[15] ),
    .A1(net1627),
    .S(net1440),
    .X(_0613_));
 sg13g2_mux2_1 _7722_ (.A0(net1803),
    .A1(net1487),
    .S(net1441),
    .X(_0614_));
 sg13g2_mux2_1 _7723_ (.A0(net1880),
    .A1(net1486),
    .S(net1440),
    .X(_0615_));
 sg13g2_mux2_1 _7724_ (.A0(net1767),
    .A1(net1794),
    .S(net1440),
    .X(_0616_));
 sg13g2_mux2_1 _7725_ (.A0(\s_m_packetdata_2_rewired[19] ),
    .A1(net1830),
    .S(net1442),
    .X(_0617_));
 sg13g2_mux2_1 _7726_ (.A0(\s_m_packetdata_2_rewired[20] ),
    .A1(net1739),
    .S(net1442),
    .X(_0618_));
 sg13g2_mux2_1 _7727_ (.A0(net1595),
    .A1(net1696),
    .S(net1440),
    .X(_0619_));
 sg13g2_mux2_1 _7728_ (.A0(net1617),
    .A1(net1161),
    .S(net1440),
    .X(_0620_));
 sg13g2_mux2_1 _7729_ (.A0(net1565),
    .A1(\s_m_packetdata_2_rewired[15] ),
    .S(net1440),
    .X(_0621_));
 sg13g2_mux2_1 _7730_ (.A0(net1803),
    .A1(net1826),
    .S(net1449),
    .X(_0622_));
 sg13g2_nor2_1 _7731_ (.A(s_m_packetdata_2_bit_17),
    .B(net1446),
    .Y(_3220_));
 sg13g2_a21oi_1 _7732_ (.A1(_0722_),
    .A2(net1446),
    .Y(_0623_),
    .B1(_3220_));
 sg13g2_mux2_1 _7733_ (.A0(net1767),
    .A1(net1756),
    .S(net1447),
    .X(_0624_));
 sg13g2_mux2_1 _7734_ (.A0(\s_m_packetdata_2_rewired[19] ),
    .A1(net1783),
    .S(net1446),
    .X(_0625_));
 sg13g2_mux2_1 _7735_ (.A0(net1759),
    .A1(net1772),
    .S(net1446),
    .X(_0626_));
 sg13g2_mux2_1 _7736_ (.A0(net1595),
    .A1(net1644),
    .S(net1446),
    .X(_0627_));
 sg13g2_mux2_1 _7737_ (.A0(net1617),
    .A1(net1597),
    .S(net1446),
    .X(_0628_));
 sg13g2_mux2_1 _7738_ (.A0(net1565),
    .A1(net1599),
    .S(net1449),
    .X(_0629_));
 sg13g2_mux2_1 _7739_ (.A0(\usbfunction0.n2481_o[16] ),
    .A1(net974),
    .S(net1445),
    .X(_0630_));
 sg13g2_nor2_1 _7740_ (.A(net966),
    .B(net1443),
    .Y(_3221_));
 sg13g2_a21oi_1 _7741_ (.A1(_0722_),
    .A2(net1443),
    .Y(_0631_),
    .B1(_3221_));
 sg13g2_mux2_1 _7742_ (.A0(net1756),
    .A1(net1483),
    .S(net1447),
    .X(_0632_));
 sg13g2_mux2_1 _7743_ (.A0(\usbfunction0.n2481_o[19] ),
    .A1(net1052),
    .S(net1447),
    .X(_0633_));
 sg13g2_mux2_1 _7744_ (.A0(\usbfunction0.n2481_o[20] ),
    .A1(net1155),
    .S(net1447),
    .X(_0634_));
 sg13g2_mux2_1 _7745_ (.A0(net1644),
    .A1(net1093),
    .S(net1447),
    .X(_0635_));
 sg13g2_mux2_1 _7746_ (.A0(net1597),
    .A1(\usbfunction0.n2481_o[30] ),
    .S(net1446),
    .X(_0636_));
 sg13g2_mux2_1 _7747_ (.A0(net1599),
    .A1(net1154),
    .S(net1446),
    .X(_0637_));
 sg13g2_mux2_1 _7748_ (.A0(net1485),
    .A1(net1615),
    .S(net1445),
    .X(_0638_));
 sg13g2_mux2_1 _7749_ (.A0(net1484),
    .A1(net1650),
    .S(net1448),
    .X(_0639_));
 sg13g2_mux2_1 _7750_ (.A0(net790),
    .A1(\usbfunction0.n2481_o[34] ),
    .S(net1448),
    .X(_0640_));
 sg13g2_mux2_1 _7751_ (.A0(net1482),
    .A1(net1691),
    .S(net1448),
    .X(_0641_));
 sg13g2_mux2_1 _7752_ (.A0(net1155),
    .A1(net1084),
    .S(net1448),
    .X(_0642_));
 sg13g2_mux2_1 _7753_ (.A0(net1093),
    .A1(\usbfunction0.n2481_o[37] ),
    .S(net1448),
    .X(_0643_));
 sg13g2_mux2_1 _7754_ (.A0(net1623),
    .A1(\usbfunction0.n2481_o[38] ),
    .S(net1448),
    .X(_0644_));
 sg13g2_mux2_1 _7755_ (.A0(net1154),
    .A1(net1109),
    .S(net1448),
    .X(_0645_));
 sg13g2_nor2_1 _7756_ (.A(net1615),
    .B(net1445),
    .Y(_3222_));
 sg13g2_a21oi_1 _7757_ (.A1(_0695_),
    .A2(net1445),
    .Y(_0646_),
    .B1(_3222_));
 sg13g2_mux2_1 _7758_ (.A0(net1667),
    .A1(net1650),
    .S(net1443),
    .X(_0647_));
 sg13g2_mux2_1 _7759_ (.A0(net1656),
    .A1(net1721),
    .S(net1443),
    .X(_0648_));
 sg13g2_nor2_1 _7760_ (.A(net1691),
    .B(net1445),
    .Y(_3223_));
 sg13g2_a21oi_1 _7761_ (.A1(_0697_),
    .A2(net1444),
    .Y(_0649_),
    .B1(_3223_));
 sg13g2_nor2_1 _7762_ (.A(net1084),
    .B(net1444),
    .Y(_3224_));
 sg13g2_a21oi_1 _7763_ (.A1(_0699_),
    .A2(net1445),
    .Y(_0650_),
    .B1(_3224_));
 sg13g2_mux2_1 _7764_ (.A0(\usbfunction0.n1583_o[5] ),
    .A1(net1635),
    .S(net1443),
    .X(_0651_));
 sg13g2_mux2_1 _7765_ (.A0(\usbfunction0.n1583_o[6] ),
    .A1(net1685),
    .S(net1443),
    .X(_0652_));
 sg13g2_nor2_1 _7766_ (.A(net1109),
    .B(net1444),
    .Y(_3225_));
 sg13g2_a21oi_1 _7767_ (.A1(_0703_),
    .A2(net1444),
    .Y(_0653_),
    .B1(_3225_));
 sg13g2_nor2_1 _7768_ (.A(net1480),
    .B(net1439),
    .Y(_3226_));
 sg13g2_a21oi_1 _7769_ (.A1(_0695_),
    .A2(net1439),
    .Y(_0654_),
    .B1(_3226_));
 sg13g2_nor2_1 _7770_ (.A(net1667),
    .B(net1444),
    .Y(_3227_));
 sg13g2_a21oi_1 _7771_ (.A1(_0706_),
    .A2(net1444),
    .Y(_0655_),
    .B1(_3227_));
 sg13g2_nor2_1 _7772_ (.A(net1656),
    .B(net1444),
    .Y(_3228_));
 sg13g2_a21oi_1 _7773_ (.A1(_0705_),
    .A2(net1444),
    .Y(_0656_),
    .B1(_3228_));
 sg13g2_nor2_1 _7774_ (.A(net1018),
    .B(net1439),
    .Y(_3229_));
 sg13g2_a21oi_1 _7775_ (.A1(_0697_),
    .A2(net1439),
    .Y(_0657_),
    .B1(_3229_));
 sg13g2_nor2_1 _7776_ (.A(net1050),
    .B(net1439),
    .Y(_3230_));
 sg13g2_a21oi_1 _7777_ (.A1(_0699_),
    .A2(net1439),
    .Y(_0658_),
    .B1(_3230_));
 sg13g2_mux2_1 _7778_ (.A0(\usbfunction0.n1583_o[5] ),
    .A1(net1592),
    .S(net1450),
    .X(_0659_));
 sg13g2_mux2_1 _7779_ (.A0(\usbfunction0.n1583_o[6] ),
    .A1(net1159),
    .S(net1450),
    .X(_0660_));
 sg13g2_nor2_1 _7780_ (.A(net873),
    .B(net1438),
    .Y(_3231_));
 sg13g2_a21oi_1 _7781_ (.A1(_0703_),
    .A2(net1438),
    .Y(_0661_),
    .B1(_3231_));
 sg13g2_nor2_1 _7782_ (.A(net1480),
    .B(net1450),
    .Y(_3232_));
 sg13g2_a21oi_1 _7783_ (.A1(net1454),
    .A2(net1450),
    .Y(_0662_),
    .B1(_3232_));
 sg13g2_nor2_1 _7784_ (.A(net1478),
    .B(net1450),
    .Y(_3233_));
 sg13g2_a21oi_1 _7785_ (.A1(net1457),
    .A2(net1450),
    .Y(_0663_),
    .B1(_3233_));
 sg13g2_nor2_1 _7786_ (.A(net1476),
    .B(net1438),
    .Y(_3234_));
 sg13g2_a21oi_1 _7787_ (.A1(_0705_),
    .A2(net1438),
    .Y(_0664_),
    .B1(_3234_));
 sg13g2_nor2_1 _7788_ (.A(net1018),
    .B(net1450),
    .Y(_3235_));
 sg13g2_a21oi_1 _7789_ (.A1(net1460),
    .A2(net1450),
    .Y(_0665_),
    .B1(_3235_));
 sg13g2_mux2_1 _7790_ (.A0(net1473),
    .A1(net1050),
    .S(net1438),
    .X(_0666_));
 sg13g2_mux2_1 _7791_ (.A0(net1470),
    .A1(net1592),
    .S(net1438),
    .X(_0667_));
 sg13g2_mux2_1 _7792_ (.A0(net1467),
    .A1(net1159),
    .S(net1438),
    .X(_0668_));
 sg13g2_mux2_1 _7793_ (.A0(net1464),
    .A1(net873),
    .S(net1438),
    .X(_0669_));
 sg13g2_nor3_1 _7794_ (.A(\usbfunction0.n2636_q ),
    .B(net1741),
    .C(net1724),
    .Y(_3236_));
 sg13g2_a21oi_1 _7795_ (.A1(\usbfunction0.n2636_q ),
    .A2(_1040_),
    .Y(_0670_),
    .B1(net1742));
 sg13g2_o21ai_1 _7796_ (.B1(_0701_),
    .Y(_3237_),
    .A1(net1697),
    .A2(_1365_));
 sg13g2_a21oi_1 _7797_ (.A1(net1454),
    .A2(_1365_),
    .Y(_0671_),
    .B1(net1698));
 sg13g2_o21ai_1 _7798_ (.B1(_0701_),
    .Y(_3238_),
    .A1(net1806),
    .A2(_1365_));
 sg13g2_a21oi_1 _7799_ (.A1(net1457),
    .A2(_1365_),
    .Y(_0672_),
    .B1(net1807));
 sg13g2_o21ai_1 _7800_ (.B1(_0701_),
    .Y(_3239_),
    .A1(net1476),
    .A2(_1366_));
 sg13g2_a21oi_1 _7801_ (.A1(_0686_),
    .A2(_1366_),
    .Y(_0673_),
    .B1(_3239_));
 sg13g2_o21ai_1 _7802_ (.B1(_0701_),
    .Y(_3240_),
    .A1(net1731),
    .A2(_1365_));
 sg13g2_a21oi_1 _7803_ (.A1(net1460),
    .A2(_1365_),
    .Y(_0674_),
    .B1(net1732));
 sg13g2_o21ai_1 _7804_ (.B1(_0029_),
    .Y(_3241_),
    .A1(\usbfunction0.scl_usbgpiophy0.scl_addeopdeferred0.n7349_q ),
    .A2(_3106_));
 sg13g2_nor2_1 _7805_ (.A(_0683_),
    .B(_0684_),
    .Y(_3242_));
 sg13g2_nand3_1 _7806_ (.B(\usbfunction0.n2313_o[2] ),
    .C(_3242_),
    .A(\usbfunction0.n2313_o[3] ),
    .Y(_3243_));
 sg13g2_nand2_1 _7807_ (.Y(_3244_),
    .A(_3241_),
    .B(_3243_));
 sg13g2_nor2_1 _7808_ (.A(net550),
    .B(_3244_),
    .Y(_3245_));
 sg13g2_nor2_1 _7809_ (.A(\usbfunction0.n2313_o[0] ),
    .B(_3241_),
    .Y(_3246_));
 sg13g2_nand2_2 _7810_ (.Y(_3247_),
    .A(_1029_),
    .B(_1366_));
 sg13g2_nor3_1 _7811_ (.A(_3245_),
    .B(_3246_),
    .C(_3247_),
    .Y(_0675_));
 sg13g2_xor2_1 _7812_ (.B(\usbfunction0.n2313_o[0] ),
    .A(net1817),
    .X(_3248_));
 sg13g2_nor2_1 _7813_ (.A(_3244_),
    .B(_3248_),
    .Y(_3249_));
 sg13g2_nor2_1 _7814_ (.A(net1817),
    .B(_3241_),
    .Y(_3250_));
 sg13g2_nor3_1 _7815_ (.A(_3247_),
    .B(_3249_),
    .C(net1818),
    .Y(_0676_));
 sg13g2_a21oi_1 _7816_ (.A1(_3241_),
    .A2(_3242_),
    .Y(_3251_),
    .B1(net1733));
 sg13g2_nor4_1 _7817_ (.A(_0682_),
    .B(_0683_),
    .C(_0684_),
    .D(_3244_),
    .Y(_3252_));
 sg13g2_nor3_1 _7818_ (.A(_3247_),
    .B(_3251_),
    .C(_3252_),
    .Y(_0677_));
 sg13g2_nor2_1 _7819_ (.A(net1854),
    .B(_3252_),
    .Y(_3253_));
 sg13g2_nor2_1 _7820_ (.A(_3247_),
    .B(net1855),
    .Y(_0678_));
 sg13g2_xnor2_1 _7821_ (.Y(_0679_),
    .A(net1717),
    .B(_0927_));
 sg13g2_nor2_1 _7822_ (.A(net1157),
    .B(_0927_),
    .Y(_3254_));
 sg13g2_nand2_1 _7823_ (.Y(_3255_),
    .A(net1461),
    .B(_3254_));
 sg13g2_xor2_1 _7824_ (.B(_3254_),
    .A(net1461),
    .X(_0680_));
 sg13g2_xnor2_1 _7825_ (.Y(_0681_),
    .A(net1567),
    .B(_3255_));
 sg13g2_mux2_1 _7826_ (.A0(_1057_),
    .A1(net1611),
    .S(net1363),
    .X(_0279_));
 sg13g2_mux2_1 _7827_ (.A0(_1049_),
    .A1(net1144),
    .S(net1363),
    .X(_0280_));
 sg13g2_o21ai_1 _7828_ (.B1(_1988_),
    .Y(_0281_),
    .A1(_1063_),
    .A2(net1363));
 sg13g2_mux2_1 _7829_ (.A0(_1053_),
    .A1(net1603),
    .S(net1363),
    .X(_0282_));
 sg13g2_mux2_1 _7830_ (.A0(net1165),
    .A1(net1105),
    .S(_1987_),
    .X(_0283_));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_dfrbp_1 _7832_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net18),
    .D(_0008_),
    .Q_N(_3722_),
    .Q(\s_m_peekdata_data_2[0] ));
 sg13g2_dfrbp_1 _7833_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net19),
    .D(_0009_),
    .Q_N(_3723_),
    .Q(\s_m_peekdata_data_2[1] ));
 sg13g2_dfrbp_1 _7834_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net20),
    .D(_0010_),
    .Q_N(_3724_),
    .Q(\s_m_peekdata_data_2[2] ));
 sg13g2_dfrbp_1 _7835_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net21),
    .D(_0011_),
    .Q_N(_3725_),
    .Q(\s_m_peekdata_data_2[3] ));
 sg13g2_dfrbp_1 _7836_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net22),
    .D(_0012_),
    .Q_N(_3726_),
    .Q(\s_m_peekdata_data_2[4] ));
 sg13g2_dfrbp_1 _7837_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net23),
    .D(_0013_),
    .Q_N(_3727_),
    .Q(\s_m_peekdata_data_2[5] ));
 sg13g2_dfrbp_1 _7838_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net24),
    .D(_0014_),
    .Q_N(_3728_),
    .Q(\s_m_peekdata_data_2[6] ));
 sg13g2_dfrbp_1 _7839_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net27),
    .D(_0015_),
    .Q_N(_3729_),
    .Q(\s_m_peekdata_data_2[7] ));
 sg13g2_dfrbp_1 _7840_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net1507),
    .D(\usbfunction0.s_m_rx_valid ),
    .Q_N(_0029_),
    .Q(\usbfunction0.n2631_q ));
 sg13g2_dfrbp_1 _7841_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net1538),
    .D(net1695),
    .Q_N(_3721_),
    .Q(\usbfunction0.n2640_q[0] ));
 sg13g2_dfrbp_1 _7842_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net1538),
    .D(net1655),
    .Q_N(_3720_),
    .Q(\usbfunction0.n2640_q[1] ));
 sg13g2_dfrbp_1 _7843_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net1508),
    .D(net1614),
    .Q_N(_3719_),
    .Q(\usbfunction0.n2640_q[2] ));
 sg13g2_dfrbp_1 _7844_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net1507),
    .D(net1562),
    .Q_N(\usbfunction0.n2640_q[3] ),
    .Q(_0161_));
 sg13g2_dfrbp_1 _7845_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net1508),
    .D(\usbfunction0.n2474_o[0] ),
    .Q_N(_3730_),
    .Q(\usbfunction0.n2634_q[0] ));
 sg13g2_dfrbp_1 _7846_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net1508),
    .D(\usbfunction0.n2474_o[1] ),
    .Q_N(_3731_),
    .Q(\usbfunction0.n2634_q[1] ));
 sg13g2_dfrbp_1 _7847_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net1508),
    .D(\usbfunction0.n2474_o[2] ),
    .Q_N(_3732_),
    .Q(\usbfunction0.n2634_q[2] ));
 sg13g2_dfrbp_1 _7848_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net1508),
    .D(\usbfunction0.n2474_o[3] ),
    .Q_N(_3718_),
    .Q(\usbfunction0.n2634_q[3] ));
 sg13g2_dfrbp_1 _7849_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net1538),
    .D(net623),
    .Q_N(_3717_),
    .Q(\usbfunction0.n2639_q ));
 sg13g2_dfrbp_1 _7850_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net1508),
    .D(_0192_),
    .Q_N(_3733_),
    .Q(\usbfunction0.n2637_q ));
 sg13g2_dfrbp_1 _7851_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net29),
    .D(net545),
    .Q_N(_3734_),
    .Q(\usbfunction0.functionreset0.in_unnamed_4[0] ));
 sg13g2_dfrbp_1 _7852_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net31),
    .D(net542),
    .Q_N(_3735_),
    .Q(\usbfunction0.functionreset0.in_unnamed_4[1] ));
 sg13g2_dfrbp_1 _7853_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net1509),
    .D(net1169),
    .Q_N(_0040_),
    .Q(s_m_pushfull));
 sg13g2_dfrbp_1 _7854_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net1526),
    .D(net1837),
    .Q_N(s_m_popempty),
    .Q(_0162_));
 sg13g2_dfrbp_1 _7855_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net1510),
    .D(\scl_fifo0.n2697_o[0] ),
    .Q_N(_3736_),
    .Q(\scl_fifo0.n2737_o[0] ));
 sg13g2_dfrbp_1 _7856_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net1510),
    .D(net1194),
    .Q_N(_0118_),
    .Q(\scl_fifo0.n2737_o[1] ));
 sg13g2_dfrbp_1 _7857_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net1509),
    .D(net1181),
    .Q_N(_0127_),
    .Q(\scl_fifo0.n2737_o[2] ));
 sg13g2_dfrbp_1 _7858_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net1509),
    .D(net1175),
    .Q_N(_0128_),
    .Q(\scl_fifo0.n2737_o[3] ));
 sg13g2_dfrbp_1 _7859_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net1509),
    .D(net1027),
    .Q_N(_0129_),
    .Q(\scl_fifo0.n2726_o ));
 sg13g2_dfrbp_1 _7860_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net1530),
    .D(_0193_),
    .Q_N(_3716_),
    .Q(\scl_bitbangengine0.s_m_value_2[0] ));
 sg13g2_dfrbp_1 _7861_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net1530),
    .D(net1117),
    .Q_N(_0133_),
    .Q(\scl_bitbangengine0.s_m_value_2[1] ));
 sg13g2_dfrbp_1 _7862_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net1530),
    .D(_0195_),
    .Q_N(_3737_),
    .Q(\scl_bitbangengine0.s_m_value_2[2] ));
 sg13g2_dfrbp_1 _7863_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net1510),
    .D(\scl_fifo0.n2694_o[0] ),
    .Q_N(_3738_),
    .Q(\scl_fifo0.n2689_o[0] ));
 sg13g2_dfrbp_1 _7864_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net1510),
    .D(\scl_fifo0.n2722_o[1] ),
    .Q_N(_0039_),
    .Q(\scl_fifo0.n2689_o[1] ));
 sg13g2_dfrbp_1 _7865_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net1505),
    .D(\scl_fifo0.n2722_o[2] ),
    .Q_N(_0122_),
    .Q(\scl_fifo0.n2689_o[2] ));
 sg13g2_dfrbp_1 _7866_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net1505),
    .D(\scl_fifo0.n2722_o[3] ),
    .Q_N(_0124_),
    .Q(\scl_fifo0.n2689_o[3] ));
 sg13g2_dfrbp_1 _7867_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net1505),
    .D(\scl_fifo0.n2722_o[4] ),
    .Q_N(_0126_),
    .Q(\scl_fifo0.n2781_q[4] ));
 sg13g2_dfrbp_1 _7868_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net1514),
    .D(net1738),
    .Q_N(_3739_),
    .Q(\scl_uarttx0.n2856_o[0] ));
 sg13g2_dfrbp_1 _7869_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net1514),
    .D(net1849),
    .Q_N(_3715_),
    .Q(\scl_uarttx0.n2856_o[1] ));
 sg13g2_dfrbp_1 _7870_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net1513),
    .D(net1643),
    .Q_N(\scl_uarttx0.n2856_o[2] ),
    .Q(_0163_));
 sg13g2_dfrbp_1 _7871_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net1513),
    .D(net993),
    .Q_N(_3740_),
    .Q(\scl_uarttx0.n2884_o ));
 sg13g2_dfrbp_1 _7872_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net1545),
    .D(net612),
    .Q_N(_3741_),
    .Q(\scl_uarttx0.scl_baudrategenerator0.n6874_o[0] ));
 sg13g2_dfrbp_1 _7873_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net1545),
    .D(\scl_uarttx0.scl_baudrategenerator0.n6892_o[1] ),
    .Q_N(_3742_),
    .Q(\scl_uarttx0.scl_baudrategenerator0.n6874_o[1] ));
 sg13g2_dfrbp_1 _7874_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net1545),
    .D(\scl_uarttx0.scl_baudrategenerator0.n6892_o[2] ),
    .Q_N(_3743_),
    .Q(\scl_uarttx0.scl_baudrategenerator0.n6874_o[2] ));
 sg13g2_dfrbp_1 _7875_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net1545),
    .D(\scl_uarttx0.scl_baudrategenerator0.n6892_o[3] ),
    .Q_N(_3744_),
    .Q(\scl_uarttx0.scl_baudrategenerator0.n6874_o[3] ));
 sg13g2_dfrbp_1 _7876_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net1545),
    .D(\scl_uarttx0.scl_baudrategenerator0.n6892_o[4] ),
    .Q_N(_3745_),
    .Q(\scl_uarttx0.scl_baudrategenerator0.n6874_o[4] ));
 sg13g2_dfrbp_1 _7877_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net1545),
    .D(\scl_uarttx0.scl_baudrategenerator0.n6892_o[5] ),
    .Q_N(_3746_),
    .Q(\scl_uarttx0.scl_baudrategenerator0.n6874_o[5] ));
 sg13g2_dfrbp_1 _7878_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net1546),
    .D(\scl_uarttx0.scl_baudrategenerator0.n6892_o[6] ),
    .Q_N(_3747_),
    .Q(\scl_uarttx0.scl_baudrategenerator0.n6874_o[6] ));
 sg13g2_dfrbp_1 _7879_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net1546),
    .D(\scl_uarttx0.scl_baudrategenerator0.n6892_o[7] ),
    .Q_N(_3748_),
    .Q(\scl_uarttx0.scl_baudrategenerator0.n6874_o[7] ));
 sg13g2_dfrbp_1 _7880_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net1541),
    .D(\scl_uarttx0.scl_baudrategenerator0.n6892_o[8] ),
    .Q_N(_3749_),
    .Q(\scl_uarttx0.scl_baudrategenerator0.n6874_o[8] ));
 sg13g2_dfrbp_1 _7881_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net1555),
    .D(\scl_uarttx0.scl_baudrategenerator0.n6892_o[9] ),
    .Q_N(_3750_),
    .Q(\scl_uarttx0.scl_baudrategenerator0.n6874_o[9] ));
 sg13g2_dfrbp_1 _7882_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net1555),
    .D(\scl_uarttx0.scl_baudrategenerator0.n6892_o[10] ),
    .Q_N(_3751_),
    .Q(\scl_uarttx0.scl_baudrategenerator0.n6874_o[10] ));
 sg13g2_dfrbp_1 _7883_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net1555),
    .D(\scl_uarttx0.scl_baudrategenerator0.n6892_o[11] ),
    .Q_N(_3752_),
    .Q(\scl_uarttx0.scl_baudrategenerator0.n6874_o[11] ));
 sg13g2_dfrbp_1 _7884_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net1555),
    .D(\scl_uarttx0.scl_baudrategenerator0.n6892_o[12] ),
    .Q_N(_3753_),
    .Q(\scl_uarttx0.scl_baudrategenerator0.n6874_o[12] ));
 sg13g2_dfrbp_1 _7885_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net1555),
    .D(\scl_uarttx0.scl_baudrategenerator0.n6892_o[13] ),
    .Q_N(_3754_),
    .Q(\scl_uarttx0.scl_baudrategenerator0.n6874_o[13] ));
 sg13g2_dfrbp_1 _7886_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net1555),
    .D(\scl_uarttx0.scl_baudrategenerator0.n6892_o[14] ),
    .Q_N(_3755_),
    .Q(\scl_uarttx0.scl_baudrategenerator0.n6874_o[14] ));
 sg13g2_dfrbp_1 _7887_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net1556),
    .D(\scl_uarttx0.scl_baudrategenerator0.n6892_o[15] ),
    .Q_N(_3756_),
    .Q(\scl_uarttx0.scl_baudrategenerator0.n6874_o[15] ));
 sg13g2_dfrbp_1 _7888_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net1556),
    .D(\scl_uarttx0.scl_baudrategenerator0.n6892_o[16] ),
    .Q_N(_3714_),
    .Q(\scl_uarttx0.scl_baudrategenerator0.n6874_o[16] ));
 sg13g2_dfrbp_1 _7889_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net222),
    .D(net746),
    .Q_N(_3713_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[15][0] ));
 sg13g2_dfrbp_1 _7890_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net221),
    .D(net643),
    .Q_N(_3712_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[15][1] ));
 sg13g2_dfrbp_1 _7891_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net220),
    .D(_0198_),
    .Q_N(_3711_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[15][2] ));
 sg13g2_dfrbp_1 _7892_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net219),
    .D(net811),
    .Q_N(_3710_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[15][3] ));
 sg13g2_dfrbp_1 _7893_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net218),
    .D(net698),
    .Q_N(_3709_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[15][4] ));
 sg13g2_dfrbp_1 _7894_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net217),
    .D(net703),
    .Q_N(_3708_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[15][5] ));
 sg13g2_dfrbp_1 _7895_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net216),
    .D(net1012),
    .Q_N(_3707_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[15][6] ));
 sg13g2_dfrbp_1 _7896_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net215),
    .D(net676),
    .Q_N(_3706_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[15][7] ));
 sg13g2_dfrbp_1 _7897_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net213),
    .D(_0204_),
    .Q_N(_3705_),
    .Q(\scl_bitbangengine0.n5920_q[3] ));
 sg13g2_dfrbp_1 _7898_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net212),
    .D(_0205_),
    .Q_N(_3704_),
    .Q(\scl_bitbangengine0.n5920_q[4] ));
 sg13g2_dfrbp_1 _7899_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net210),
    .D(_0206_),
    .Q_N(_3703_),
    .Q(\scl_bitbangengine0.n5920_q[5] ));
 sg13g2_dfrbp_1 _7900_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net209),
    .D(net1038),
    .Q_N(_0145_),
    .Q(\scl_bitbangengine0.n5920_q[6] ));
 sg13g2_dfrbp_1 _7901_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net208),
    .D(net1787),
    .Q_N(_3702_),
    .Q(\scl_bitbangengine0.n5920_q[7] ));
 sg13g2_dfrbp_1 _7902_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net207),
    .D(_0209_),
    .Q_N(_3701_),
    .Q(\scl_bitbangengine0.n5920_q[8] ));
 sg13g2_dfrbp_1 _7903_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net1522),
    .D(net1893),
    .Q_N(_3700_),
    .Q(\scl_bitbangengine0.n5898_q[0] ));
 sg13g2_dfrbp_1 _7904_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net1522),
    .D(_0211_),
    .Q_N(_3699_),
    .Q(\scl_bitbangengine0.n5898_q[1] ));
 sg13g2_dfrbp_1 _7905_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net1513),
    .D(_0212_),
    .Q_N(_3698_),
    .Q(\scl_bitbangengine0.n5898_q[2] ));
 sg13g2_dfrbp_1 _7906_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net1513),
    .D(_0213_),
    .Q_N(_3697_),
    .Q(\scl_bitbangengine0.n5898_q[3] ));
 sg13g2_dfrbp_1 _7907_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net1530),
    .D(net753),
    .Q_N(_0131_),
    .Q(\scl_bitbangengine0.s_m_value[0] ));
 sg13g2_dfrbp_1 _7908_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net1530),
    .D(net568),
    .Q_N(_0120_),
    .Q(\scl_bitbangengine0.s_m_value[1] ));
 sg13g2_dfrbp_1 _7909_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net1530),
    .D(net925),
    .Q_N(_0132_),
    .Q(\scl_bitbangengine0.s_m_value[2] ));
 sg13g2_dfrbp_1 _7910_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net1519),
    .D(\scl_bitbangengine0.scl_counter0.n6954_o[0] ),
    .Q_N(_3757_),
    .Q(\scl_bitbangengine0.scl_counter0.n6975_q[0] ));
 sg13g2_dfrbp_1 _7911_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net1515),
    .D(\scl_bitbangengine0.scl_counter0.n6954_o[1] ),
    .Q_N(_3758_),
    .Q(\scl_bitbangengine0.scl_counter0.n6975_q[1] ));
 sg13g2_dfrbp_1 _7912_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net1519),
    .D(net1659),
    .Q_N(_0062_),
    .Q(\scl_bitbangengine0.scl_counter0.n6975_q[2] ));
 sg13g2_dfrbp_1 _7913_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net1515),
    .D(\scl_bitbangengine0.scl_counter0.n6954_o[3] ),
    .Q_N(_0064_),
    .Q(\scl_bitbangengine0.scl_counter0.n6975_q[3] ));
 sg13g2_dfrbp_1 _7914_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net1515),
    .D(net1707),
    .Q_N(_0065_),
    .Q(\scl_bitbangengine0.scl_counter0.n6975_q[4] ));
 sg13g2_dfrbp_1 _7915_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net1515),
    .D(\scl_bitbangengine0.scl_counter0.n6954_o[5] ),
    .Q_N(_0066_),
    .Q(\scl_bitbangengine0.scl_counter0.n6975_q[5] ));
 sg13g2_dfrbp_1 _7916_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net1515),
    .D(net1730),
    .Q_N(_0067_),
    .Q(\scl_bitbangengine0.scl_counter0.n6975_q[6] ));
 sg13g2_dfrbp_1 _7917_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net1515),
    .D(\scl_bitbangengine0.scl_counter0.n6954_o[7] ),
    .Q_N(_0069_),
    .Q(\scl_bitbangengine0.scl_counter0.n6975_q[7] ));
 sg13g2_dfrbp_1 _7918_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net1516),
    .D(net1815),
    .Q_N(_0070_),
    .Q(\scl_bitbangengine0.scl_counter0.n6975_q[8] ));
 sg13g2_dfrbp_1 _7919_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net1515),
    .D(\scl_bitbangengine0.scl_counter0.n6954_o[9] ),
    .Q_N(_0071_),
    .Q(\scl_bitbangengine0.scl_counter0.n6975_q[9] ));
 sg13g2_dfrbp_1 _7920_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net1516),
    .D(net1748),
    .Q_N(_0072_),
    .Q(\scl_bitbangengine0.scl_counter0.n6975_q[10] ));
 sg13g2_dfrbp_1 _7921_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net1516),
    .D(\scl_bitbangengine0.scl_counter0.n6954_o[11] ),
    .Q_N(_0074_),
    .Q(\scl_bitbangengine0.scl_counter0.n6975_q[11] ));
 sg13g2_dfrbp_1 _7922_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net1516),
    .D(\scl_bitbangengine0.scl_counter0.n6954_o[12] ),
    .Q_N(_0075_),
    .Q(\scl_bitbangengine0.scl_counter0.n6975_q[12] ));
 sg13g2_dfrbp_1 _7923_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net1516),
    .D(\scl_bitbangengine0.scl_counter0.n6954_o[13] ),
    .Q_N(_0076_),
    .Q(\scl_bitbangengine0.scl_counter0.n6975_q[13] ));
 sg13g2_dfrbp_1 _7924_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net1517),
    .D(net1609),
    .Q_N(_0077_),
    .Q(\scl_bitbangengine0.scl_counter0.n6975_q[14] ));
 sg13g2_dfrbp_1 _7925_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net1517),
    .D(\scl_bitbangengine0.scl_counter0.n6954_o[15] ),
    .Q_N(_0079_),
    .Q(\scl_bitbangengine0.scl_counter0.n6975_q[15] ));
 sg13g2_dfrbp_1 _7926_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net1517),
    .D(\scl_bitbangengine0.scl_counter0.n6954_o[16] ),
    .Q_N(_0080_),
    .Q(\scl_bitbangengine0.scl_counter0.n6975_q[16] ));
 sg13g2_dfrbp_1 _7927_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net206),
    .D(_0217_),
    .Q_N(_3696_),
    .Q(\scl_bitbangengine0.n5905_q ));
 sg13g2_dfrbp_1 _7928_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net204),
    .D(net789),
    .Q_N(_3695_),
    .Q(\s_out_3[2] ));
 sg13g2_dfrbp_1 _7929_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net203),
    .D(net869),
    .Q_N(_3694_),
    .Q(\s_out_3[5] ));
 sg13g2_dfrbp_1 _7930_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net1513),
    .D(_0220_),
    .Q_N(_0084_),
    .Q(\scl_bitbangengine0.n3817_o ));
 sg13g2_dfrbp_1 _7931_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net202),
    .D(_0221_),
    .Q_N(_3693_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[0][0] ));
 sg13g2_dfrbp_1 _7932_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net201),
    .D(_0222_),
    .Q_N(_3692_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[0][1] ));
 sg13g2_dfrbp_1 _7933_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net200),
    .D(_0223_),
    .Q_N(_3691_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[0][2] ));
 sg13g2_dfrbp_1 _7934_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net199),
    .D(_0224_),
    .Q_N(_3690_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[0][3] ));
 sg13g2_dfrbp_1 _7935_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net198),
    .D(_0225_),
    .Q_N(_3689_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[0][4] ));
 sg13g2_dfrbp_1 _7936_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net197),
    .D(_0226_),
    .Q_N(_3688_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[0][5] ));
 sg13g2_dfrbp_1 _7937_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net196),
    .D(_0227_),
    .Q_N(_3687_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[0][6] ));
 sg13g2_dfrbp_1 _7938_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net195),
    .D(_0228_),
    .Q_N(_3686_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[0][7] ));
 sg13g2_dfrbp_1 _7939_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net194),
    .D(_0229_),
    .Q_N(_3685_),
    .Q(\usbfunction0.n2645_q[2] ));
 sg13g2_dfrbp_1 _7940_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net1522),
    .D(net860),
    .Q_N(_3684_),
    .Q(\scl_bitbangengine0.n5923_q ));
 sg13g2_dfrbp_1 _7941_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net1520),
    .D(net596),
    .Q_N(_3683_),
    .Q(s_m_io15_out));
 sg13g2_dfrbp_1 _7942_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net192),
    .D(_0232_),
    .Q_N(_3682_),
    .Q(\scl_bitbangengine0.n5902_q ));
 sg13g2_dfrbp_1 _7943_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net1520),
    .D(_0233_),
    .Q_N(_3681_),
    .Q(s_m_io14_out));
 sg13g2_dfrbp_1 _7944_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net1521),
    .D(_0234_),
    .Q_N(_3680_),
    .Q(s_m_io1_out));
 sg13g2_dfrbp_1 _7945_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net1521),
    .D(_0235_),
    .Q_N(_3759_),
    .Q(s_m_io13_out));
 sg13g2_dfrbp_1 _7946_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net191),
    .D(\scl_bitbangengine0.n3871_o ),
    .Q_N(_3679_),
    .Q(\scl_bitbangengine0.n3336_o ));
 sg13g2_dfrbp_1 _7947_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net1521),
    .D(_0236_),
    .Q_N(_3678_),
    .Q(s_m_io12_out));
 sg13g2_dfrbp_1 _7948_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net190),
    .D(_0237_),
    .Q_N(_3677_),
    .Q(\scl_bitbangengine0.n5910_q ));
 sg13g2_dfrbp_1 _7949_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net1531),
    .D(_0238_),
    .Q_N(_3676_),
    .Q(s_m_io11_out));
 sg13g2_dfrbp_1 _7950_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net188),
    .D(_0239_),
    .Q_N(_3675_),
    .Q(\scl_bitbangengine0.n5903_q ));
 sg13g2_dfrbp_1 _7951_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net1521),
    .D(_0240_),
    .Q_N(_3674_),
    .Q(s_m_io10_out));
 sg13g2_dfrbp_1 _7952_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net186),
    .D(net915),
    .Q_N(_3673_),
    .Q(\scl_bitbangengine0.n5904_q ));
 sg13g2_dfrbp_1 _7953_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net1521),
    .D(_0242_),
    .Q_N(_3672_),
    .Q(s_m_io9_out));
 sg13g2_dfrbp_1 _7954_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net1520),
    .D(_0243_),
    .Q_N(_3671_),
    .Q(\scl_bitbangengine0.n5909_q ));
 sg13g2_dfrbp_1 _7955_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net1521),
    .D(net946),
    .Q_N(_3760_),
    .Q(n153_o));
 sg13g2_dfrbp_1 _7956_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net1520),
    .D(\scl_bitbangengine0.n3839_o ),
    .Q_N(_3670_),
    .Q(\scl_bitbangengine0.n5907_q ));
 sg13g2_dfrbp_1 _7957_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net1518),
    .D(net995),
    .Q_N(_3761_),
    .Q(s_m_io5_opendrain));
 sg13g2_dfrbp_1 _7958_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net1532),
    .D(net932),
    .Q_N(_0134_),
    .Q(\scl_bitbangengine0.n5423_o[0] ));
 sg13g2_dfrbp_1 _7959_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net1532),
    .D(net1147),
    .Q_N(_0135_),
    .Q(\scl_bitbangengine0.n5423_o[1] ));
 sg13g2_dfrbp_1 _7960_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net1532),
    .D(net1564),
    .Q_N(_0136_),
    .Q(\scl_bitbangengine0.n5423_o[2] ));
 sg13g2_dfrbp_1 _7961_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net1532),
    .D(\scl_bitbangengine0.n5462_o[3] ),
    .Q_N(_0137_),
    .Q(\scl_bitbangengine0.n5423_o[3] ));
 sg13g2_dfrbp_1 _7962_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net1532),
    .D(net1591),
    .Q_N(_0138_),
    .Q(\scl_bitbangengine0.n5423_o[4] ));
 sg13g2_dfrbp_1 _7963_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net1532),
    .D(net1136),
    .Q_N(_0139_),
    .Q(\scl_bitbangengine0.n5423_o[5] ));
 sg13g2_dfrbp_1 _7964_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net1531),
    .D(net1622),
    .Q_N(_0140_),
    .Q(\scl_bitbangengine0.n5423_o[6] ));
 sg13g2_dfrbp_1 _7965_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net1531),
    .D(net1652),
    .Q_N(_3669_),
    .Q(\scl_bitbangengine0.n5924_q[7] ));
 sg13g2_dfrbp_1 _7966_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net184),
    .D(_0246_),
    .Q_N(_3668_),
    .Q(\s_out_3[3] ));
 sg13g2_dfrbp_1 _7967_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net1518),
    .D(_0247_),
    .Q_N(_3667_),
    .Q(s_m_io5_en));
 sg13g2_dfrbp_1 _7968_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net183),
    .D(net1089),
    .Q_N(_3666_),
    .Q(\scl_bitbangengine0.n5918_q ));
 sg13g2_dfrbp_1 _7969_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net1516),
    .D(net1131),
    .Q_N(_3665_),
    .Q(s_m_io5_out));
 sg13g2_dfrbp_1 _7970_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net1517),
    .D(net890),
    .Q_N(_3664_),
    .Q(s_m_io0_opendrain));
 sg13g2_dfrbp_1 _7971_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net1516),
    .D(net1666),
    .Q_N(_3663_),
    .Q(s_m_io4_opendrain));
 sg13g2_dfrbp_1 _7972_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net1518),
    .D(net826),
    .Q_N(_3662_),
    .Q(s_m_io4_en));
 sg13g2_dfrbp_1 _7973_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net1522),
    .D(net684),
    .Q_N(_0141_),
    .Q(\scl_bitbangengine0.n5913_q ));
 sg13g2_dfrbp_1 _7974_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net1520),
    .D(net1833),
    .Q_N(_3661_),
    .Q(s_m_io4_out));
 sg13g2_dfrbp_1 _7975_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net97),
    .D(net577),
    .Q_N(_3762_),
    .Q(\scl_bitbangengine0.n5915_q ));
 sg13g2_dfrbp_1 _7976_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net1517),
    .D(\scl_bitbangengine0.n3793_o ),
    .Q_N(_3660_),
    .Q(s_m_io3_en));
 sg13g2_dfrbp_1 _7977_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net1517),
    .D(net886),
    .Q_N(_3763_),
    .Q(s_m_io0_out));
 sg13g2_dfrbp_1 _7978_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net1520),
    .D(\scl_bitbangengine0.n5401_o ),
    .Q_N(_3659_),
    .Q(s_m_io3_out));
 sg13g2_dfrbp_1 _7979_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net181),
    .D(net988),
    .Q_N(_3658_),
    .Q(\scl_bitbangengine0.n5917_q ));
 sg13g2_dfrbp_1 _7980_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net1517),
    .D(_0258_),
    .Q_N(_3657_),
    .Q(s_m_io3_opendrain));
 sg13g2_dfrbp_1 _7981_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net101),
    .D(net1802),
    .Q_N(_3764_),
    .Q(\scl_bitbangengine0.n5911_q ));
 sg13g2_dfrbp_1 _7982_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net102),
    .D(_0016_),
    .Q_N(_3765_),
    .Q(\usbfunction0.s_m_descdata[0] ));
 sg13g2_dfrbp_1 _7983_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net103),
    .D(_0017_),
    .Q_N(_3766_),
    .Q(\usbfunction0.s_m_descdata[1] ));
 sg13g2_dfrbp_1 _7984_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net104),
    .D(_0018_),
    .Q_N(_3767_),
    .Q(\usbfunction0.s_m_descdata[2] ));
 sg13g2_dfrbp_1 _7985_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net105),
    .D(_0019_),
    .Q_N(_3768_),
    .Q(\usbfunction0.s_m_descdata[3] ));
 sg13g2_dfrbp_1 _7986_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net106),
    .D(_0020_),
    .Q_N(_3769_),
    .Q(\usbfunction0.s_m_descdata[4] ));
 sg13g2_dfrbp_1 _7987_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net126),
    .D(_0021_),
    .Q_N(_3770_),
    .Q(\usbfunction0.s_m_descdata[5] ));
 sg13g2_dfrbp_1 _7988_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net180),
    .D(_0022_),
    .Q_N(_3656_),
    .Q(\usbfunction0.s_m_descdata[6] ));
 sg13g2_dfrbp_1 _7989_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net178),
    .D(net1639),
    .Q_N(_3655_),
    .Q(\s_out_3[6] ));
 sg13g2_dfrbp_1 _7990_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net1518),
    .D(net1032),
    .Q_N(_3654_),
    .Q(s_m_io2_opendrain));
 sg13g2_dfrbp_1 _7991_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net177),
    .D(net718),
    .Q_N(_3653_),
    .Q(\s_out_3[4] ));
 sg13g2_dfrbp_1 _7992_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net1513),
    .D(_0263_),
    .Q_N(\scl_bitbangengine0.n5919_q ),
    .Q(_0164_));
 sg13g2_dfrbp_1 _7993_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net1516),
    .D(_0264_),
    .Q_N(_3652_),
    .Q(s_m_io2_en));
 sg13g2_dfrbp_1 _7994_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net1511),
    .D(_0265_),
    .Q_N(_3651_),
    .Q(\scl_bitbangengine0.n3663_o[0] ));
 sg13g2_dfrbp_1 _7995_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net1512),
    .D(_0266_),
    .Q_N(_3650_),
    .Q(\scl_bitbangengine0.n3663_o[1] ));
 sg13g2_dfrbp_1 _7996_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net1511),
    .D(_0267_),
    .Q_N(_0073_),
    .Q(\scl_bitbangengine0.n3663_o[2] ));
 sg13g2_dfrbp_1 _7997_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net1511),
    .D(_0268_),
    .Q_N(_3649_),
    .Q(\scl_bitbangengine0.n3663_o[3] ));
 sg13g2_dfrbp_1 _7998_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net1512),
    .D(net1780),
    .Q_N(_3648_),
    .Q(\scl_bitbangengine0.n3663_o[4] ));
 sg13g2_dfrbp_1 _7999_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net1512),
    .D(_0270_),
    .Q_N(_3647_),
    .Q(\scl_bitbangengine0.n3663_o[5] ));
 sg13g2_dfrbp_1 _8000_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net1519),
    .D(net857),
    .Q_N(_0078_),
    .Q(\scl_bitbangengine0.n3663_o[6] ));
 sg13g2_dfrbp_1 _8001_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net1522),
    .D(_0272_),
    .Q_N(_3646_),
    .Q(\scl_bitbangengine0.n3663_o[7] ));
 sg13g2_dfrbp_1 _8002_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net1513),
    .D(_0273_),
    .Q_N(_3645_),
    .Q(\scl_bitbangengine0.n3663_o[8] ));
 sg13g2_dfrbp_1 _8003_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net1518),
    .D(_0274_),
    .Q_N(_3644_),
    .Q(s_m_io2_out));
 sg13g2_dfrbp_1 _8004_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net1517),
    .D(net852),
    .Q_N(_3643_),
    .Q(s_m_io0_en));
 sg13g2_dfrbp_1 _8005_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net1520),
    .D(_0276_),
    .Q_N(_3642_),
    .Q(s_m_io1_opendrain));
 sg13g2_dfrbp_1 _8006_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net1520),
    .D(_0277_),
    .Q_N(_3641_),
    .Q(s_m_io1_en));
 sg13g2_dfrbp_1 _8007_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net1558),
    .D(_0278_),
    .Q_N(_3771_),
    .Q(\scl_uartrx0.n6119_q ));
 sg13g2_dfrbp_1 _8008_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net1546),
    .D(\scl_uartrx0.scl_baudrategenerator0.n7069_o[0] ),
    .Q_N(_0037_),
    .Q(\scl_uartrx0.scl_baudrategenerator0.n7047_o[0] ));
 sg13g2_dfrbp_1 _8009_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net1545),
    .D(\scl_uartrx0.scl_baudrategenerator0.n7069_o[1] ),
    .Q_N(_3772_),
    .Q(\scl_uartrx0.scl_baudrategenerator0.n7047_o[1] ));
 sg13g2_dfrbp_1 _8010_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net1558),
    .D(\scl_uartrx0.scl_baudrategenerator0.n7069_o[2] ),
    .Q_N(_3773_),
    .Q(\scl_uartrx0.scl_baudrategenerator0.n7047_o[2] ));
 sg13g2_dfrbp_1 _8011_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net1545),
    .D(\scl_uartrx0.scl_baudrategenerator0.n7069_o[3] ),
    .Q_N(_3774_),
    .Q(\scl_uartrx0.scl_baudrategenerator0.n7047_o[3] ));
 sg13g2_dfrbp_1 _8012_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net1557),
    .D(\scl_uartrx0.scl_baudrategenerator0.n7069_o[4] ),
    .Q_N(_3775_),
    .Q(\scl_uartrx0.scl_baudrategenerator0.n7047_o[4] ));
 sg13g2_dfrbp_1 _8013_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net1557),
    .D(\scl_uartrx0.scl_baudrategenerator0.n7069_o[5] ),
    .Q_N(_3776_),
    .Q(\scl_uartrx0.scl_baudrategenerator0.n7047_o[5] ));
 sg13g2_dfrbp_1 _8014_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net1557),
    .D(\scl_uartrx0.scl_baudrategenerator0.n7069_o[6] ),
    .Q_N(_3777_),
    .Q(\scl_uartrx0.scl_baudrategenerator0.n7047_o[6] ));
 sg13g2_dfrbp_1 _8015_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net1557),
    .D(\scl_uartrx0.scl_baudrategenerator0.n7069_o[7] ),
    .Q_N(_3778_),
    .Q(\scl_uartrx0.scl_baudrategenerator0.n7047_o[7] ));
 sg13g2_dfrbp_1 _8016_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net1557),
    .D(\scl_uartrx0.scl_baudrategenerator0.n7069_o[8] ),
    .Q_N(_3779_),
    .Q(\scl_uartrx0.scl_baudrategenerator0.n7047_o[8] ));
 sg13g2_dfrbp_1 _8017_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net1557),
    .D(\scl_uartrx0.scl_baudrategenerator0.n7069_o[9] ),
    .Q_N(_3780_),
    .Q(\scl_uartrx0.scl_baudrategenerator0.n7047_o[9] ));
 sg13g2_dfrbp_1 _8018_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net1557),
    .D(\scl_uartrx0.scl_baudrategenerator0.n7069_o[10] ),
    .Q_N(_3781_),
    .Q(\scl_uartrx0.scl_baudrategenerator0.n7047_o[10] ));
 sg13g2_dfrbp_1 _8019_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net1557),
    .D(\scl_uartrx0.scl_baudrategenerator0.n7069_o[11] ),
    .Q_N(_3782_),
    .Q(\scl_uartrx0.scl_baudrategenerator0.n7047_o[11] ));
 sg13g2_dfrbp_1 _8020_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net1555),
    .D(\scl_uartrx0.scl_baudrategenerator0.n7069_o[12] ),
    .Q_N(_3783_),
    .Q(\scl_uartrx0.scl_baudrategenerator0.n7047_o[12] ));
 sg13g2_dfrbp_1 _8021_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net1555),
    .D(\scl_uartrx0.scl_baudrategenerator0.n7069_o[13] ),
    .Q_N(_3784_),
    .Q(\scl_uartrx0.scl_baudrategenerator0.n7047_o[13] ));
 sg13g2_dfrbp_1 _8022_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net1558),
    .D(\scl_uartrx0.scl_baudrategenerator0.n7069_o[14] ),
    .Q_N(_3785_),
    .Q(\scl_uartrx0.scl_baudrategenerator0.n7047_o[14] ));
 sg13g2_dfrbp_1 _8023_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net1558),
    .D(\scl_uartrx0.scl_baudrategenerator0.n7069_o[15] ),
    .Q_N(_3786_),
    .Q(\scl_uartrx0.scl_baudrategenerator0.n7047_o[15] ));
 sg13g2_dfrbp_1 _8024_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net1556),
    .D(\scl_uartrx0.scl_baudrategenerator0.n7069_o[16] ),
    .Q_N(_3787_),
    .Q(\scl_uartrx0.scl_baudrategenerator0.n7047_o[16] ));
 sg13g2_dfrbp_1 _8025_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net174),
    .D(\scl_uartrx0.n6047_o ),
    .Q_N(_0151_),
    .Q(s_out_valid_2));
 sg13g2_dfrbp_1 _8026_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net1550),
    .D(_0279_),
    .Q_N(_3640_),
    .Q(\scl_fifo1.n6323_q[0] ));
 sg13g2_dfrbp_1 _8027_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net1550),
    .D(net1145),
    .Q_N(_3639_),
    .Q(\scl_fifo1.n6323_q[1] ));
 sg13g2_dfrbp_1 _8028_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net1550),
    .D(_0281_),
    .Q_N(_3638_),
    .Q(\scl_fifo1.n6323_q[2] ));
 sg13g2_dfrbp_1 _8029_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net1550),
    .D(_0282_),
    .Q_N(_3637_),
    .Q(\scl_fifo1.n6323_q[3] ));
 sg13g2_dfrbp_1 _8030_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net1551),
    .D(_0283_),
    .Q_N(_3636_),
    .Q(\scl_fifo1.n6323_q[4] ));
 sg13g2_dfrbp_1 _8031_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net134),
    .D(_0284_),
    .Q_N(_3788_),
    .Q(\s_out_3[0] ));
 sg13g2_dfrbp_1 _8032_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net1553),
    .D(net565),
    .Q_N(_3635_),
    .Q(\scl_streamarbiter_2.n6192_q ));
 sg13g2_dfrbp_1 _8033_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net1533),
    .D(net557),
    .Q_N(\scl_streamarbiter_2.n6195_q ),
    .Q(_0165_));
 sg13g2_dfrbp_1 _8034_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net1532),
    .D(\scl_streamarbiter_2.n6146_o ),
    .Q_N(_3789_),
    .Q(\scl_streamarbiter_2.n6194_q ));
 sg13g2_dfrbp_1 _8035_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net1552),
    .D(net1283),
    .Q_N(_3790_),
    .Q(\scl_fifo1.n6321_q[0] ));
 sg13g2_dfrbp_1 _8036_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net1552),
    .D(net1294),
    .Q_N(_0146_),
    .Q(\scl_fifo1.n6321_q[1] ));
 sg13g2_dfrbp_1 _8037_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net1550),
    .D(net1273),
    .Q_N(_0147_),
    .Q(\scl_fifo1.n6321_q[2] ));
 sg13g2_dfrbp_1 _8038_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net1550),
    .D(net1266),
    .Q_N(_0148_),
    .Q(\scl_fifo1.n6321_q[3] ));
 sg13g2_dfrbp_1 _8039_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net1551),
    .D(\scl_fifo1.n6238_o[4] ),
    .Q_N(_3634_),
    .Q(\scl_fifo1.n6321_q[4] ));
 sg13g2_dfrbp_1 _8040_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net1552),
    .D(_0178_),
    .Q_N(s_m_popempty_2),
    .Q(_0166_));
 sg13g2_dfrbp_1 _8041_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net1533),
    .D(net1770),
    .Q_N(_0150_),
    .Q(s_m_pushfull_2));
 sg13g2_dfrbp_1 _8042_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net1550),
    .D(net1612),
    .Q_N(_3791_),
    .Q(\scl_fifo1.n6278_o[0] ));
 sg13g2_dfrbp_1 _8043_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net1550),
    .D(\scl_fifo1.n6239_o[1] ),
    .Q_N(_3792_),
    .Q(\scl_fifo1.n6278_o[1] ));
 sg13g2_dfrbp_1 _8044_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net1551),
    .D(net893),
    .Q_N(_3793_),
    .Q(\scl_fifo1.n6278_o[2] ));
 sg13g2_dfrbp_1 _8045_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net1551),
    .D(net1604),
    .Q_N(_3794_),
    .Q(\scl_fifo1.n6278_o[3] ));
 sg13g2_dfrbp_1 _8046_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net1551),
    .D(net1106),
    .Q_N(_3633_),
    .Q(\scl_fifo1.n6267_o ));
 sg13g2_dfrbp_1 _8047_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net1510),
    .D(net671),
    .Q_N(_0130_),
    .Q(\scl_fifo0.n2711_o[0] ));
 sg13g2_dfrbp_1 _8048_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net1505),
    .D(net688),
    .Q_N(_0038_),
    .Q(\scl_fifo0.n2711_o[1] ));
 sg13g2_dfrbp_1 _8049_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net1505),
    .D(_0287_),
    .Q_N(_0121_),
    .Q(\scl_fifo0.n2711_o[2] ));
 sg13g2_dfrbp_1 _8050_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net1509),
    .D(net580),
    .Q_N(_0123_),
    .Q(\scl_fifo0.n2711_o[3] ));
 sg13g2_dfrbp_1 _8051_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net1509),
    .D(net1059),
    .Q_N(_0125_),
    .Q(\scl_fifo0.n2700_o ));
 sg13g2_dfrbp_1 _8052_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net1553),
    .D(\scl_fifo1.n6233_o[0] ),
    .Q_N(_0149_),
    .Q(\scl_fifo1.n6229_o[0] ));
 sg13g2_dfrbp_1 _8053_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net1554),
    .D(\scl_fifo1.n6233_o[1] ),
    .Q_N(_0152_),
    .Q(\scl_fifo1.n6229_o[1] ));
 sg13g2_dfrbp_1 _8054_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net1554),
    .D(\scl_fifo1.n6233_o[2] ),
    .Q_N(_0153_),
    .Q(\scl_fifo1.n6229_o[2] ));
 sg13g2_dfrbp_1 _8055_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net1554),
    .D(net582),
    .Q_N(_0154_),
    .Q(\scl_fifo1.n6229_o[3] ));
 sg13g2_dfrbp_1 _8056_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net1551),
    .D(\scl_fifo1.n6233_o[4] ),
    .Q_N(_0155_),
    .Q(\scl_fifo1.n6242_o ));
 sg13g2_dfrbp_1 _8057_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net172),
    .D(_0290_),
    .Q_N(_3632_),
    .Q(\s_out_3[7] ));
 sg13g2_dfrbp_1 _8058_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net1528),
    .D(net1134),
    .Q_N(_3795_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_insertbeat0.n7369_o ));
 sg13g2_dfrbp_1 _8059_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net1543),
    .D(net877),
    .Q_N(_3796_),
    .Q(\n353_q[0] ));
 sg13g2_dfrbp_1 _8060_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net1543),
    .D(net1071),
    .Q_N(_3797_),
    .Q(\n353_q[1] ));
 sg13g2_dfrbp_1 _8061_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net1543),
    .D(net1574),
    .Q_N(_3798_),
    .Q(\n353_q[2] ));
 sg13g2_dfrbp_1 _8062_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net1548),
    .D(net1101),
    .Q_N(_3799_),
    .Q(\n353_q[3] ));
 sg13g2_dfrbp_1 _8063_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net1543),
    .D(net1150),
    .Q_N(_3800_),
    .Q(\n353_q[4] ));
 sg13g2_dfrbp_1 _8064_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net1543),
    .D(net1083),
    .Q_N(_3801_),
    .Q(\n353_q[5] ));
 sg13g2_dfrbp_1 _8065_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net1543),
    .D(net1113),
    .Q_N(_3802_),
    .Q(\n353_q[6] ));
 sg13g2_dfrbp_1 _8066_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net1544),
    .D(\n352_o[7] ),
    .Q_N(_3803_),
    .Q(\n353_q[7] ));
 sg13g2_dfrbp_1 _8067_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net1544),
    .D(\n352_o[8] ),
    .Q_N(_3631_),
    .Q(\n353_q[8] ));
 sg13g2_dfrbp_1 _8068_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net1544),
    .D(_0179_),
    .Q_N(\n353_q[9] ),
    .Q(_0167_));
 sg13g2_dfrbp_1 _8069_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net1544),
    .D(\n352_o[10] ),
    .Q_N(_3804_),
    .Q(\n353_q[10] ));
 sg13g2_dfrbp_1 _8070_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net1543),
    .D(net1860),
    .Q_N(_3805_),
    .Q(\n353_q[11] ));
 sg13g2_dfrbp_1 _8071_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net1543),
    .D(\n352_o[12] ),
    .Q_N(_3806_),
    .Q(\n353_q[12] ));
 sg13g2_dfrbp_1 _8072_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net1546),
    .D(\n352_o[13] ),
    .Q_N(_3630_),
    .Q(\n353_q[13] ));
 sg13g2_dfrbp_1 _8073_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net1547),
    .D(_0180_),
    .Q_N(\n353_q[14] ),
    .Q(_0168_));
 sg13g2_dfrbp_1 _8074_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net1546),
    .D(_0181_),
    .Q_N(\n353_q[15] ),
    .Q(_0169_));
 sg13g2_dfrbp_1 _8075_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net1541),
    .D(_0182_),
    .Q_N(\n353_q[16] ),
    .Q(_0170_));
 sg13g2_dfrbp_1 _8076_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net1541),
    .D(\n352_o[17] ),
    .Q_N(_3807_),
    .Q(\n353_q[17] ));
 sg13g2_dfrbp_1 _8077_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net1546),
    .D(net1805),
    .Q_N(_3808_),
    .Q(\n353_q[18] ));
 sg13g2_dfrbp_1 _8078_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net1541),
    .D(\n352_o[19] ),
    .Q_N(_3809_),
    .Q(\n353_q[19] ));
 sg13g2_dfrbp_1 _8079_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net1541),
    .D(\n352_o[20] ),
    .Q_N(_3810_),
    .Q(\n353_q[20] ));
 sg13g2_dfrbp_1 _8080_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net1542),
    .D(\n352_o[21] ),
    .Q_N(_3811_),
    .Q(\n353_q[21] ));
 sg13g2_dfrbp_1 _8081_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net1542),
    .D(\n352_o[22] ),
    .Q_N(_3812_),
    .Q(\n353_q[22] ));
 sg13g2_dfrbp_1 _8082_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net1541),
    .D(\n352_o[23] ),
    .Q_N(_3813_),
    .Q(\n353_q[23] ));
 sg13g2_dfrbp_1 _8083_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net1541),
    .D(n350_o),
    .Q_N(_3814_),
    .Q(n351_q));
 sg13g2_dfrbp_1 _8084_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net1541),
    .D(n183_o),
    .Q_N(_3629_),
    .Q(n349_q));
 sg13g2_dfrbp_1 _8085_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net166),
    .D(_0292_),
    .Q_N(_3628_),
    .Q(\usbfunction0.s_m_rx_data[0] ));
 sg13g2_dfrbp_1 _8086_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net165),
    .D(_0293_),
    .Q_N(_3627_),
    .Q(\usbfunction0.s_m_rx_data[1] ));
 sg13g2_dfrbp_1 _8087_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net164),
    .D(_0294_),
    .Q_N(_3626_),
    .Q(\usbfunction0.s_m_rx_data[2] ));
 sg13g2_dfrbp_1 _8088_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net163),
    .D(_0295_),
    .Q_N(_3625_),
    .Q(\usbfunction0.s_m_rx_data[3] ));
 sg13g2_dfrbp_1 _8089_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net162),
    .D(_0296_),
    .Q_N(_3624_),
    .Q(\usbfunction0.s_m_rx_data[4] ));
 sg13g2_dfrbp_1 _8090_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net154),
    .D(_0297_),
    .Q_N(_3623_),
    .Q(\usbfunction0.s_m_rx_data[5] ));
 sg13g2_dfrbp_1 _8091_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net153),
    .D(_0298_),
    .Q_N(_3622_),
    .Q(\usbfunction0.s_m_rx_data[6] ));
 sg13g2_dfrbp_1 _8092_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net1542),
    .D(_0299_),
    .Q_N(_3621_),
    .Q(n347_q));
 sg13g2_dfrbp_1 _8093_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net155),
    .D(net690),
    .Q_N(_3815_),
    .Q(\s_out_3[1] ));
 sg13g2_dfrbp_1 _8094_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net156),
    .D(_0000_),
    .Q_N(\scl_bitbangengine0.n3241_o ),
    .Q(\scl_bitbangengine0.n3230_o ));
 sg13g2_dfrbp_1 _8095_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net157),
    .D(_0001_),
    .Q_N(_0083_),
    .Q(\scl_bitbangengine0.n3198_o ));
 sg13g2_dfrbp_1 _8096_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net158),
    .D(_0002_),
    .Q_N(_3816_),
    .Q(\scl_bitbangengine0.n3737_o ));
 sg13g2_dfrbp_1 _8097_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net159),
    .D(_0003_),
    .Q_N(\scl_bitbangengine0.n3865_o ),
    .Q(\scl_bitbangengine0.n3740_o ));
 sg13g2_dfrbp_1 _8098_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net160),
    .D(_0004_),
    .Q_N(_3817_),
    .Q(\scl_bitbangengine0.n3257_o ));
 sg13g2_dfrbp_1 _8099_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net161),
    .D(_0005_),
    .Q_N(_3818_),
    .Q(\scl_bitbangengine0.n3267_o ));
 sg13g2_dfrbp_1 _8100_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net211),
    .D(_0006_),
    .Q_N(_3819_),
    .Q(\scl_bitbangengine0.n3258_o ));
 sg13g2_dfrbp_1 _8101_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net152),
    .D(_0007_),
    .Q_N(_3620_),
    .Q(\scl_bitbangengine0.n3179_o ));
 sg13g2_dfrbp_1 _8102_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net151),
    .D(net673),
    .Q_N(_3619_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[14][0] ));
 sg13g2_dfrbp_1 _8103_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net150),
    .D(net616),
    .Q_N(_3618_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[14][1] ));
 sg13g2_dfrbp_1 _8104_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net149),
    .D(_0303_),
    .Q_N(_3617_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[14][2] ));
 sg13g2_dfrbp_1 _8105_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net148),
    .D(net653),
    .Q_N(_3616_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[14][3] ));
 sg13g2_dfrbp_1 _8106_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net147),
    .D(net1126),
    .Q_N(_3615_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[14][4] ));
 sg13g2_dfrbp_1 _8107_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net146),
    .D(net1123),
    .Q_N(_3614_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[14][5] ));
 sg13g2_dfrbp_1 _8108_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net145),
    .D(_0307_),
    .Q_N(_3613_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[14][6] ));
 sg13g2_dfrbp_1 _8109_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net144),
    .D(net1062),
    .Q_N(_3612_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[14][7] ));
 sg13g2_dfrbp_1 _8110_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net143),
    .D(_0309_),
    .Q_N(_3611_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[13][0] ));
 sg13g2_dfrbp_1 _8111_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net142),
    .D(_0310_),
    .Q_N(_3610_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[13][1] ));
 sg13g2_dfrbp_1 _8112_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net141),
    .D(_0311_),
    .Q_N(_3609_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[13][2] ));
 sg13g2_dfrbp_1 _8113_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net140),
    .D(_0312_),
    .Q_N(_3608_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[13][3] ));
 sg13g2_dfrbp_1 _8114_ (.CLK(clknet_leaf_112_clk_regs),
    .RESET_B(net139),
    .D(_0313_),
    .Q_N(_3607_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[13][4] ));
 sg13g2_dfrbp_1 _8115_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net138),
    .D(_0314_),
    .Q_N(_3606_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[13][5] ));
 sg13g2_dfrbp_1 _8116_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net137),
    .D(_0315_),
    .Q_N(_3605_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[13][6] ));
 sg13g2_dfrbp_1 _8117_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net136),
    .D(_0316_),
    .Q_N(_3604_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[13][7] ));
 sg13g2_dfrbp_1 _8118_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net135),
    .D(_0317_),
    .Q_N(_3603_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[12][0] ));
 sg13g2_dfrbp_1 _8119_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net133),
    .D(_0318_),
    .Q_N(_3602_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[12][1] ));
 sg13g2_dfrbp_1 _8120_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net132),
    .D(_0319_),
    .Q_N(_3601_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[12][2] ));
 sg13g2_dfrbp_1 _8121_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net131),
    .D(_0320_),
    .Q_N(_3600_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[12][3] ));
 sg13g2_dfrbp_1 _8122_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net130),
    .D(_0321_),
    .Q_N(_3599_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[12][4] ));
 sg13g2_dfrbp_1 _8123_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net129),
    .D(_0322_),
    .Q_N(_3598_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[12][5] ));
 sg13g2_dfrbp_1 _8124_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net128),
    .D(_0323_),
    .Q_N(_3597_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[12][6] ));
 sg13g2_dfrbp_1 _8125_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net127),
    .D(_0324_),
    .Q_N(_3596_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[12][7] ));
 sg13g2_dfrbp_1 _8126_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net125),
    .D(_0325_),
    .Q_N(_3595_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[11][0] ));
 sg13g2_dfrbp_1 _8127_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net124),
    .D(_0326_),
    .Q_N(_3594_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[11][1] ));
 sg13g2_dfrbp_1 _8128_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net123),
    .D(_0327_),
    .Q_N(_3593_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[11][2] ));
 sg13g2_dfrbp_1 _8129_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net122),
    .D(_0328_),
    .Q_N(_3592_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[11][3] ));
 sg13g2_dfrbp_1 _8130_ (.CLK(clknet_leaf_112_clk_regs),
    .RESET_B(net121),
    .D(_0329_),
    .Q_N(_3591_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[11][4] ));
 sg13g2_dfrbp_1 _8131_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net120),
    .D(_0330_),
    .Q_N(_3590_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[11][5] ));
 sg13g2_dfrbp_1 _8132_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net119),
    .D(_0331_),
    .Q_N(_3589_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[11][6] ));
 sg13g2_dfrbp_1 _8133_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net118),
    .D(_0332_),
    .Q_N(_3588_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[11][7] ));
 sg13g2_dfrbp_1 _8134_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net117),
    .D(net649),
    .Q_N(_3587_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[10][0] ));
 sg13g2_dfrbp_1 _8135_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net116),
    .D(_0334_),
    .Q_N(_3586_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[10][1] ));
 sg13g2_dfrbp_1 _8136_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net115),
    .D(_0335_),
    .Q_N(_3585_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[10][2] ));
 sg13g2_dfrbp_1 _8137_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net114),
    .D(_0336_),
    .Q_N(_3584_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[10][3] ));
 sg13g2_dfrbp_1 _8138_ (.CLK(clknet_leaf_112_clk_regs),
    .RESET_B(net113),
    .D(_0337_),
    .Q_N(_3583_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[10][4] ));
 sg13g2_dfrbp_1 _8139_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net112),
    .D(_0338_),
    .Q_N(_3582_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[10][5] ));
 sg13g2_dfrbp_1 _8140_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net111),
    .D(_0339_),
    .Q_N(_3581_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[10][6] ));
 sg13g2_dfrbp_1 _8141_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net110),
    .D(_0340_),
    .Q_N(_3580_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[10][7] ));
 sg13g2_dfrbp_1 _8142_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net109),
    .D(_0341_),
    .Q_N(_3579_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[0][0] ));
 sg13g2_dfrbp_1 _8143_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net108),
    .D(net639),
    .Q_N(_3578_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[0][1] ));
 sg13g2_dfrbp_1 _8144_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net107),
    .D(_0343_),
    .Q_N(_3577_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[0][2] ));
 sg13g2_dfrbp_1 _8145_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net100),
    .D(_0344_),
    .Q_N(_3576_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[0][3] ));
 sg13g2_dfrbp_1 _8146_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net99),
    .D(_0345_),
    .Q_N(_3575_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[0][4] ));
 sg13g2_dfrbp_1 _8147_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net98),
    .D(_0346_),
    .Q_N(_3574_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[0][5] ));
 sg13g2_dfrbp_1 _8148_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net96),
    .D(_0347_),
    .Q_N(_3573_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[0][6] ));
 sg13g2_dfrbp_1 _8149_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net95),
    .D(_0348_),
    .Q_N(_3572_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[0][7] ));
 sg13g2_dfrbp_1 _8150_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net94),
    .D(_0349_),
    .Q_N(_3571_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[8][0] ));
 sg13g2_dfrbp_1 _8151_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net93),
    .D(_0350_),
    .Q_N(_3570_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[8][1] ));
 sg13g2_dfrbp_1 _8152_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net92),
    .D(_0351_),
    .Q_N(_3569_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[8][2] ));
 sg13g2_dfrbp_1 _8153_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net91),
    .D(_0352_),
    .Q_N(_3568_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[8][3] ));
 sg13g2_dfrbp_1 _8154_ (.CLK(clknet_leaf_112_clk_regs),
    .RESET_B(net90),
    .D(_0353_),
    .Q_N(_3567_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[8][4] ));
 sg13g2_dfrbp_1 _8155_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net89),
    .D(_0354_),
    .Q_N(_3566_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[8][5] ));
 sg13g2_dfrbp_1 _8156_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net88),
    .D(_0355_),
    .Q_N(_3565_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[8][6] ));
 sg13g2_dfrbp_1 _8157_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net87),
    .D(_0356_),
    .Q_N(_3564_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[8][7] ));
 sg13g2_dfrbp_1 _8158_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net86),
    .D(_0357_),
    .Q_N(_3563_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[7][0] ));
 sg13g2_dfrbp_1 _8159_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net85),
    .D(_0358_),
    .Q_N(_3562_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[7][1] ));
 sg13g2_dfrbp_1 _8160_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net84),
    .D(_0359_),
    .Q_N(_3561_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[7][2] ));
 sg13g2_dfrbp_1 _8161_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net83),
    .D(_0360_),
    .Q_N(_3560_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[7][3] ));
 sg13g2_dfrbp_1 _8162_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net82),
    .D(_0361_),
    .Q_N(_3559_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[7][4] ));
 sg13g2_dfrbp_1 _8163_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net81),
    .D(_0362_),
    .Q_N(_3558_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[7][5] ));
 sg13g2_dfrbp_1 _8164_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net80),
    .D(_0363_),
    .Q_N(_3557_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[7][6] ));
 sg13g2_dfrbp_1 _8165_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net79),
    .D(_0364_),
    .Q_N(_3556_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[7][7] ));
 sg13g2_dfrbp_1 _8166_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net78),
    .D(_0365_),
    .Q_N(_3555_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[6][0] ));
 sg13g2_dfrbp_1 _8167_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net77),
    .D(_0366_),
    .Q_N(_3554_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[6][1] ));
 sg13g2_dfrbp_1 _8168_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net76),
    .D(_0367_),
    .Q_N(_3553_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[6][2] ));
 sg13g2_dfrbp_1 _8169_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net75),
    .D(_0368_),
    .Q_N(_3552_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[6][3] ));
 sg13g2_dfrbp_1 _8170_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net74),
    .D(_0369_),
    .Q_N(_3551_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[6][4] ));
 sg13g2_dfrbp_1 _8171_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net73),
    .D(_0370_),
    .Q_N(_3550_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[6][5] ));
 sg13g2_dfrbp_1 _8172_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net72),
    .D(_0371_),
    .Q_N(_3549_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[6][6] ));
 sg13g2_dfrbp_1 _8173_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net71),
    .D(_0372_),
    .Q_N(_3548_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[6][7] ));
 sg13g2_dfrbp_1 _8174_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net70),
    .D(_0373_),
    .Q_N(_3547_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[5][0] ));
 sg13g2_dfrbp_1 _8175_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net69),
    .D(_0374_),
    .Q_N(_3546_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[5][1] ));
 sg13g2_dfrbp_1 _8176_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net68),
    .D(_0375_),
    .Q_N(_3545_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[5][2] ));
 sg13g2_dfrbp_1 _8177_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net67),
    .D(_0376_),
    .Q_N(_3544_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[5][3] ));
 sg13g2_dfrbp_1 _8178_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net66),
    .D(_0377_),
    .Q_N(_3543_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[5][4] ));
 sg13g2_dfrbp_1 _8179_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net65),
    .D(_0378_),
    .Q_N(_3542_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[5][5] ));
 sg13g2_dfrbp_1 _8180_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net64),
    .D(_0379_),
    .Q_N(_3541_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[5][6] ));
 sg13g2_dfrbp_1 _8181_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net63),
    .D(_0380_),
    .Q_N(_3540_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[5][7] ));
 sg13g2_dfrbp_1 _8182_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net62),
    .D(_0381_),
    .Q_N(_3539_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[4][0] ));
 sg13g2_dfrbp_1 _8183_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net61),
    .D(_0382_),
    .Q_N(_3538_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[4][1] ));
 sg13g2_dfrbp_1 _8184_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net60),
    .D(_0383_),
    .Q_N(_3537_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[4][2] ));
 sg13g2_dfrbp_1 _8185_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net59),
    .D(_0384_),
    .Q_N(_3536_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[4][3] ));
 sg13g2_dfrbp_1 _8186_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net58),
    .D(_0385_),
    .Q_N(_3535_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[4][4] ));
 sg13g2_dfrbp_1 _8187_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net57),
    .D(_0386_),
    .Q_N(_3534_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[4][5] ));
 sg13g2_dfrbp_1 _8188_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net56),
    .D(_0387_),
    .Q_N(_3533_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[4][6] ));
 sg13g2_dfrbp_1 _8189_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net55),
    .D(_0388_),
    .Q_N(_3532_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[4][7] ));
 sg13g2_dfrbp_1 _8190_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net54),
    .D(_0389_),
    .Q_N(_3531_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[3][0] ));
 sg13g2_dfrbp_1 _8191_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net53),
    .D(net666),
    .Q_N(_3530_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[3][1] ));
 sg13g2_dfrbp_1 _8192_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net52),
    .D(_0391_),
    .Q_N(_3529_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[3][2] ));
 sg13g2_dfrbp_1 _8193_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net51),
    .D(_0392_),
    .Q_N(_3528_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[3][3] ));
 sg13g2_dfrbp_1 _8194_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net50),
    .D(_0393_),
    .Q_N(_3527_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[3][4] ));
 sg13g2_dfrbp_1 _8195_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net49),
    .D(net696),
    .Q_N(_3526_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[3][5] ));
 sg13g2_dfrbp_1 _8196_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net48),
    .D(_0395_),
    .Q_N(_3525_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[3][6] ));
 sg13g2_dfrbp_1 _8197_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net47),
    .D(net681),
    .Q_N(_3524_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[3][7] ));
 sg13g2_dfrbp_1 _8198_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net46),
    .D(_0397_),
    .Q_N(_3523_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[1][0] ));
 sg13g2_dfrbp_1 _8199_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net45),
    .D(net614),
    .Q_N(_3522_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[1][1] ));
 sg13g2_dfrbp_1 _8200_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net44),
    .D(_0399_),
    .Q_N(_3521_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[1][2] ));
 sg13g2_dfrbp_1 _8201_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net43),
    .D(_0400_),
    .Q_N(_3520_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[1][3] ));
 sg13g2_dfrbp_1 _8202_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net42),
    .D(_0401_),
    .Q_N(_3519_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[1][4] ));
 sg13g2_dfrbp_1 _8203_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net41),
    .D(_0402_),
    .Q_N(_3518_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[1][5] ));
 sg13g2_dfrbp_1 _8204_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net40),
    .D(_0403_),
    .Q_N(_3517_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[1][6] ));
 sg13g2_dfrbp_1 _8205_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net39),
    .D(_0404_),
    .Q_N(_3516_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[1][7] ));
 sg13g2_dfrbp_1 _8206_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net38),
    .D(_0405_),
    .Q_N(_3515_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[2][0] ));
 sg13g2_dfrbp_1 _8207_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net37),
    .D(net713),
    .Q_N(_3514_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[2][1] ));
 sg13g2_dfrbp_1 _8208_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net36),
    .D(_0407_),
    .Q_N(_3513_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[2][2] ));
 sg13g2_dfrbp_1 _8209_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net35),
    .D(_0408_),
    .Q_N(_3512_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[2][3] ));
 sg13g2_dfrbp_1 _8210_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net34),
    .D(_0409_),
    .Q_N(_3511_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[2][4] ));
 sg13g2_dfrbp_1 _8211_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net33),
    .D(net1140),
    .Q_N(_3510_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[2][5] ));
 sg13g2_dfrbp_1 _8212_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net32),
    .D(_0411_),
    .Q_N(_3509_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[2][6] ));
 sg13g2_dfrbp_1 _8213_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net30),
    .D(_0412_),
    .Q_N(_3508_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[2][7] ));
 sg13g2_dfrbp_1 _8214_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net1558),
    .D(net553),
    .Q_N(\scl_uartrx0.n6053_o ),
    .Q(_0171_));
 sg13g2_dfrbp_1 _8215_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net1556),
    .D(_0023_),
    .Q_N(_3820_),
    .Q(\scl_uartrx0.n5991_o ));
 sg13g2_dfrbp_1 _8216_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net1556),
    .D(_0024_),
    .Q_N(_3821_),
    .Q(\scl_uartrx0.n6074_o ));
 sg13g2_dfrbp_1 _8217_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net1556),
    .D(_0025_),
    .Q_N(_3507_),
    .Q(\scl_uartrx0.n6090_o ));
 sg13g2_dfrbp_1 _8218_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net1514),
    .D(_0413_),
    .Q_N(_0119_),
    .Q(n346_q));
 sg13g2_dfrbp_1 _8219_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net214),
    .D(_0414_),
    .Q_N(_3822_),
    .Q(\usbfunction0.s_m_descdata[7] ));
 sg13g2_dfrbp_1 _8220_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net1509),
    .D(net549),
    .Q_N(_0041_),
    .Q(\usbfunction0.n1974_o ));
 sg13g2_dfrbp_1 _8221_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net1553),
    .D(net584),
    .Q_N(_3823_),
    .Q(\usbfunction0.functionreset0.n6707_q[0] ));
 sg13g2_dfrbp_1 _8222_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net1553),
    .D(net1678),
    .Q_N(_3824_),
    .Q(\usbfunction0.functionreset0.n6707_q[1] ));
 sg13g2_dfrbp_1 _8223_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net1553),
    .D(\usbfunction0.functionreset0.n6674_o[2] ),
    .Q_N(_3825_),
    .Q(\usbfunction0.functionreset0.n6707_q[2] ));
 sg13g2_dfrbp_1 _8224_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net1532),
    .D(net796),
    .Q_N(_3826_),
    .Q(\usbfunction0.functionreset0.n6707_q[3] ));
 sg13g2_dfrbp_1 _8225_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net1533),
    .D(\usbfunction0.functionreset0.n6674_o[4] ),
    .Q_N(_3827_),
    .Q(\usbfunction0.functionreset0.n6707_q[4] ));
 sg13g2_dfrbp_1 _8226_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net1534),
    .D(\usbfunction0.functionreset0.n6674_o[5] ),
    .Q_N(_3828_),
    .Q(\usbfunction0.functionreset0.n6707_q[5] ));
 sg13g2_dfrbp_1 _8227_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net1534),
    .D(\usbfunction0.functionreset0.n6674_o[6] ),
    .Q_N(_3829_),
    .Q(\usbfunction0.functionreset0.n6707_q[6] ));
 sg13g2_dfrbp_1 _8228_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net1553),
    .D(\usbfunction0.functionreset0.n6674_o[7] ),
    .Q_N(_3830_),
    .Q(\usbfunction0.functionreset0.n6707_q[7] ));
 sg13g2_dfrbp_1 _8229_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net1553),
    .D(\usbfunction0.functionreset0.n6674_o[8] ),
    .Q_N(_3831_),
    .Q(\usbfunction0.functionreset0.n6707_q[8] ));
 sg13g2_dfrbp_1 _8230_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net1553),
    .D(net604),
    .Q_N(_3832_),
    .Q(\usbfunction0.functionreset0.n6707_q[9] ));
 sg13g2_dfrbp_1 _8231_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net1539),
    .D(\usbfunction0.functionreset0.n6683_o ),
    .Q_N(_3506_),
    .Q(\usbfunction0.functionreset0.n6708_q ));
 sg13g2_dfrbp_1 _8232_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net26),
    .D(_0415_),
    .Q_N(_3505_),
    .Q(\scl_bitbangengine0.n5920_q[0] ));
 sg13g2_dfrbp_1 _8233_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net25),
    .D(net1723),
    .Q_N(_3504_),
    .Q(\scl_bitbangengine0.n5920_q[1] ));
 sg13g2_dfrbp_1 _8234_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net17),
    .D(net1606),
    .Q_N(_3503_),
    .Q(\scl_bitbangengine0.n5920_q[2] ));
 sg13g2_dfrbp_1 _8235_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net1528),
    .D(net560),
    .Q_N(\usbfunction0.scl_usbgpiophy0.n6405_o ),
    .Q(_0172_));
 sg13g2_dfrbp_1 _8236_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net1528),
    .D(_0026_),
    .Q_N(_3833_),
    .Q(\usbfunction0.scl_usbgpiophy0.n6437_o ));
 sg13g2_dfrbp_1 _8237_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net1528),
    .D(net1171),
    .Q_N(_3834_),
    .Q(\usbfunction0.scl_usbgpiophy0.n6411_o ));
 sg13g2_dfrbp_1 _8238_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net1528),
    .D(_0028_),
    .Q_N(_3835_),
    .Q(\usbfunction0.scl_usbgpiophy0.n6449_o ));
 sg13g2_dfrbp_1 _8239_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net1507),
    .D(s_m_status_rxactive),
    .Q_N(_3502_),
    .Q(\usbfunction0.scl_usbgpiophy0.n6650_q ));
 sg13g2_dfrbp_1 _8240_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net1538),
    .D(_0418_),
    .Q_N(_3501_),
    .Q(\usbfunction0.n2635_q[0] ));
 sg13g2_dfrbp_1 _8241_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net1538),
    .D(net1725),
    .Q_N(_3500_),
    .Q(\usbfunction0.n2635_q[1] ));
 sg13g2_dfrbp_1 _8242_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net1527),
    .D(net600),
    .Q_N(_3836_),
    .Q(\usbfunction0.scl_usbgpiophy0.n6653_q ));
 sg13g2_dfrbp_1 _8243_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net1524),
    .D(\usbfunction0.scl_usbgpiophy0.s_ret_3 ),
    .Q_N(_3837_),
    .Q(\usbfunction0.scl_usbgpiophy0.n6655_q ));
 sg13g2_dfrbp_1 _8244_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net1529),
    .D(\usbfunction0.scl_usbgpiophy0.n6529_o ),
    .Q_N(_3838_),
    .Q(\usbfunction0.scl_usbgpiophy0.n6646_q ));
 sg13g2_dfrbp_1 _8245_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net1538),
    .D(s_m_phy_tx_valid_2),
    .Q_N(_3839_),
    .Q(\usbfunction0.scl_usbgpiophy0.n6654_q ));
 sg13g2_dfrbp_1 _8246_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net1507),
    .D(net539),
    .Q_N(\usbfunction0.s_m_rx_sop ),
    .Q(\usbfunction0.scl_usbgpiophy0.n6649_q ));
 sg13g2_dfrbp_1 _8247_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net525),
    .D(net750),
    .Q_N(_3499_),
    .Q(s_m_match_delayed1));
 sg13g2_dfrbp_1 _8248_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net224),
    .D(net1736),
    .Q_N(_3840_),
    .Q(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.in_unnamed ));
 sg13g2_dfrbp_1 _8249_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net1507),
    .D(net572),
    .Q_N(_3841_),
    .Q(\usbfunction0.scl_usbgpiophy0.n6651_q ));
 sg13g2_dfrbp_1 _8250_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net1531),
    .D(net15),
    .Q_N(_3842_),
    .Q(\usbfunction0.scl_usbgpiophy0.s_linein ));
 sg13g2_dfrbp_1 _8251_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net1530),
    .D(net1437),
    .Q_N(_0042_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_recoverdatadifferential0.scl_recoverdatadifferential_equalsampling_sky1300.n7883_q ));
 sg13g2_dfrbp_1 _8252_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net524),
    .D(_0423_),
    .Q_N(_3498_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[15][0] ));
 sg13g2_dfrbp_1 _8253_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net523),
    .D(_0424_),
    .Q_N(_3497_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[15][1] ));
 sg13g2_dfrbp_1 _8254_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net522),
    .D(_0425_),
    .Q_N(_3496_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[15][2] ));
 sg13g2_dfrbp_1 _8255_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net475),
    .D(_0426_),
    .Q_N(_3495_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[15][3] ));
 sg13g2_dfrbp_1 _8256_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net444),
    .D(_0427_),
    .Q_N(_3494_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[15][4] ));
 sg13g2_dfrbp_1 _8257_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net443),
    .D(_0428_),
    .Q_N(_3493_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[15][5] ));
 sg13g2_dfrbp_1 _8258_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net442),
    .D(_0429_),
    .Q_N(_3492_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[15][6] ));
 sg13g2_dfrbp_1 _8259_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net441),
    .D(_0430_),
    .Q_N(_3491_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[15][7] ));
 sg13g2_dfrbp_1 _8260_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net440),
    .D(_0431_),
    .Q_N(_3490_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[14][0] ));
 sg13g2_dfrbp_1 _8261_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net439),
    .D(_0432_),
    .Q_N(_3489_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[14][1] ));
 sg13g2_dfrbp_1 _8262_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net438),
    .D(_0433_),
    .Q_N(_3488_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[14][2] ));
 sg13g2_dfrbp_1 _8263_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net437),
    .D(_0434_),
    .Q_N(_3487_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[14][3] ));
 sg13g2_dfrbp_1 _8264_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net436),
    .D(_0435_),
    .Q_N(_3486_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[14][4] ));
 sg13g2_dfrbp_1 _8265_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net435),
    .D(_0436_),
    .Q_N(_3485_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[14][5] ));
 sg13g2_dfrbp_1 _8266_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net434),
    .D(_0437_),
    .Q_N(_3484_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[14][6] ));
 sg13g2_dfrbp_1 _8267_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net433),
    .D(_0438_),
    .Q_N(_3483_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[14][7] ));
 sg13g2_dfrbp_1 _8268_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net432),
    .D(_0439_),
    .Q_N(_3482_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[13][0] ));
 sg13g2_dfrbp_1 _8269_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net431),
    .D(_0440_),
    .Q_N(_3481_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[13][1] ));
 sg13g2_dfrbp_1 _8270_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net430),
    .D(_0441_),
    .Q_N(_3480_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[13][2] ));
 sg13g2_dfrbp_1 _8271_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net429),
    .D(_0442_),
    .Q_N(_3479_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[13][3] ));
 sg13g2_dfrbp_1 _8272_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net428),
    .D(_0443_),
    .Q_N(_3478_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[13][4] ));
 sg13g2_dfrbp_1 _8273_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net427),
    .D(_0444_),
    .Q_N(_3477_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[13][5] ));
 sg13g2_dfrbp_1 _8274_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net426),
    .D(_0445_),
    .Q_N(_3476_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[13][6] ));
 sg13g2_dfrbp_1 _8275_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net425),
    .D(_0446_),
    .Q_N(_3475_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[13][7] ));
 sg13g2_dfrbp_1 _8276_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net424),
    .D(_0447_),
    .Q_N(_3474_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[12][0] ));
 sg13g2_dfrbp_1 _8277_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net423),
    .D(_0448_),
    .Q_N(_3473_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[12][1] ));
 sg13g2_dfrbp_1 _8278_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net422),
    .D(_0449_),
    .Q_N(_3472_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[12][2] ));
 sg13g2_dfrbp_1 _8279_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net421),
    .D(_0450_),
    .Q_N(_3471_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[12][3] ));
 sg13g2_dfrbp_1 _8280_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net420),
    .D(_0451_),
    .Q_N(_3470_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[12][4] ));
 sg13g2_dfrbp_1 _8281_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net419),
    .D(_0452_),
    .Q_N(_3469_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[12][5] ));
 sg13g2_dfrbp_1 _8282_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net418),
    .D(_0453_),
    .Q_N(_3468_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[12][6] ));
 sg13g2_dfrbp_1 _8283_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net417),
    .D(_0454_),
    .Q_N(_3467_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[12][7] ));
 sg13g2_dfrbp_1 _8284_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net416),
    .D(_0455_),
    .Q_N(_3466_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[11][0] ));
 sg13g2_dfrbp_1 _8285_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net415),
    .D(_0456_),
    .Q_N(_3465_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[11][1] ));
 sg13g2_dfrbp_1 _8286_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net414),
    .D(_0457_),
    .Q_N(_3464_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[11][2] ));
 sg13g2_dfrbp_1 _8287_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net413),
    .D(_0458_),
    .Q_N(_3463_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[11][3] ));
 sg13g2_dfrbp_1 _8288_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net412),
    .D(_0459_),
    .Q_N(_3462_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[11][4] ));
 sg13g2_dfrbp_1 _8289_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net411),
    .D(_0460_),
    .Q_N(_3461_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[11][5] ));
 sg13g2_dfrbp_1 _8290_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net410),
    .D(_0461_),
    .Q_N(_3460_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[11][6] ));
 sg13g2_dfrbp_1 _8291_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net409),
    .D(_0462_),
    .Q_N(_3459_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[11][7] ));
 sg13g2_dfrbp_1 _8292_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net408),
    .D(_0463_),
    .Q_N(_3458_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[10][0] ));
 sg13g2_dfrbp_1 _8293_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net407),
    .D(_0464_),
    .Q_N(_3457_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[10][1] ));
 sg13g2_dfrbp_1 _8294_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net406),
    .D(_0465_),
    .Q_N(_3456_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[10][2] ));
 sg13g2_dfrbp_1 _8295_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net405),
    .D(_0466_),
    .Q_N(_3455_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[10][3] ));
 sg13g2_dfrbp_1 _8296_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net404),
    .D(_0467_),
    .Q_N(_3454_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[10][4] ));
 sg13g2_dfrbp_1 _8297_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net403),
    .D(_0468_),
    .Q_N(_3453_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[10][5] ));
 sg13g2_dfrbp_1 _8298_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net402),
    .D(_0469_),
    .Q_N(_3452_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[10][6] ));
 sg13g2_dfrbp_1 _8299_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net401),
    .D(_0470_),
    .Q_N(_3451_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[10][7] ));
 sg13g2_dfrbp_1 _8300_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net400),
    .D(_0471_),
    .Q_N(_3450_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[9][0] ));
 sg13g2_dfrbp_1 _8301_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net399),
    .D(_0472_),
    .Q_N(_3449_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[9][1] ));
 sg13g2_dfrbp_1 _8302_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net398),
    .D(_0473_),
    .Q_N(_3448_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[9][2] ));
 sg13g2_dfrbp_1 _8303_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net397),
    .D(_0474_),
    .Q_N(_3447_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[9][3] ));
 sg13g2_dfrbp_1 _8304_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net396),
    .D(_0475_),
    .Q_N(_3446_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[9][4] ));
 sg13g2_dfrbp_1 _8305_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net395),
    .D(_0476_),
    .Q_N(_3445_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[9][5] ));
 sg13g2_dfrbp_1 _8306_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net394),
    .D(_0477_),
    .Q_N(_3444_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[9][6] ));
 sg13g2_dfrbp_1 _8307_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net393),
    .D(_0478_),
    .Q_N(_3443_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[9][7] ));
 sg13g2_dfrbp_1 _8308_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net392),
    .D(_0479_),
    .Q_N(_3442_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[8][0] ));
 sg13g2_dfrbp_1 _8309_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net391),
    .D(_0480_),
    .Q_N(_3441_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[8][1] ));
 sg13g2_dfrbp_1 _8310_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net390),
    .D(_0481_),
    .Q_N(_3440_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[8][2] ));
 sg13g2_dfrbp_1 _8311_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net389),
    .D(_0482_),
    .Q_N(_3439_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[8][3] ));
 sg13g2_dfrbp_1 _8312_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net388),
    .D(_0483_),
    .Q_N(_3438_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[8][4] ));
 sg13g2_dfrbp_1 _8313_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net387),
    .D(_0484_),
    .Q_N(_3437_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[8][5] ));
 sg13g2_dfrbp_1 _8314_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net386),
    .D(_0485_),
    .Q_N(_3436_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[8][6] ));
 sg13g2_dfrbp_1 _8315_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net385),
    .D(_0486_),
    .Q_N(_3435_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[8][7] ));
 sg13g2_dfrbp_1 _8316_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net384),
    .D(_0487_),
    .Q_N(_3434_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[7][0] ));
 sg13g2_dfrbp_1 _8317_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net383),
    .D(_0488_),
    .Q_N(_3433_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[7][1] ));
 sg13g2_dfrbp_1 _8318_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net382),
    .D(_0489_),
    .Q_N(_3432_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[7][2] ));
 sg13g2_dfrbp_1 _8319_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net381),
    .D(_0490_),
    .Q_N(_3431_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[7][3] ));
 sg13g2_dfrbp_1 _8320_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net380),
    .D(_0491_),
    .Q_N(_3430_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[7][4] ));
 sg13g2_dfrbp_1 _8321_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net379),
    .D(_0492_),
    .Q_N(_3429_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[7][5] ));
 sg13g2_dfrbp_1 _8322_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net376),
    .D(_0493_),
    .Q_N(_3428_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[7][6] ));
 sg13g2_dfrbp_1 _8323_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net375),
    .D(_0494_),
    .Q_N(_3427_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[7][7] ));
 sg13g2_dfrbp_1 _8324_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net374),
    .D(_0495_),
    .Q_N(_3426_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[6][0] ));
 sg13g2_dfrbp_1 _8325_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net373),
    .D(_0496_),
    .Q_N(_3425_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[6][1] ));
 sg13g2_dfrbp_1 _8326_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net372),
    .D(_0497_),
    .Q_N(_3424_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[6][2] ));
 sg13g2_dfrbp_1 _8327_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net371),
    .D(_0498_),
    .Q_N(_3423_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[6][3] ));
 sg13g2_dfrbp_1 _8328_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net370),
    .D(_0499_),
    .Q_N(_3422_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[6][4] ));
 sg13g2_dfrbp_1 _8329_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net369),
    .D(_0500_),
    .Q_N(_3421_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[6][5] ));
 sg13g2_dfrbp_1 _8330_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net368),
    .D(_0501_),
    .Q_N(_3420_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[6][6] ));
 sg13g2_dfrbp_1 _8331_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net367),
    .D(_0502_),
    .Q_N(_3419_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[6][7] ));
 sg13g2_dfrbp_1 _8332_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net366),
    .D(_0503_),
    .Q_N(_3418_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[5][0] ));
 sg13g2_dfrbp_1 _8333_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net365),
    .D(_0504_),
    .Q_N(_3417_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[5][1] ));
 sg13g2_dfrbp_1 _8334_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net364),
    .D(_0505_),
    .Q_N(_3416_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[5][2] ));
 sg13g2_dfrbp_1 _8335_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net363),
    .D(_0506_),
    .Q_N(_3415_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[5][3] ));
 sg13g2_dfrbp_1 _8336_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net362),
    .D(_0507_),
    .Q_N(_3414_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[5][4] ));
 sg13g2_dfrbp_1 _8337_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net361),
    .D(_0508_),
    .Q_N(_3413_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[5][5] ));
 sg13g2_dfrbp_1 _8338_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net360),
    .D(_0509_),
    .Q_N(_3412_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[5][6] ));
 sg13g2_dfrbp_1 _8339_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net326),
    .D(_0510_),
    .Q_N(_3843_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[5][7] ));
 sg13g2_dfrbp_1 _8340_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net1531),
    .D(net16),
    .Q_N(_3411_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_recoverdatadifferential0.scl_recoverdatadifferential_equalsampling_sky1300.detectsingleended0.n9022_q ));
 sg13g2_dfrbp_1 _8341_ (.CLK(net528),
    .RESET_B(net359),
    .D(net16),
    .Q_N(_3410_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_recoverdatadifferential0.scl_recoverdatadifferential_equalsampling_sky1300.detectsingleended0.n9024_q ));
 sg13g2_dfrbp_1 _8342_ (.CLK(net529),
    .RESET_B(net358),
    .D(net15),
    .Q_N(_3409_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_recoverdatadifferential0.scl_recoverdatadifferential_equalsampling_sky1300.detectsingleended0.n9025_q ));
 sg13g2_dfrbp_1 _8343_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net357),
    .D(_0511_),
    .Q_N(_3408_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[4][0] ));
 sg13g2_dfrbp_1 _8344_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net356),
    .D(_0512_),
    .Q_N(_3407_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[4][1] ));
 sg13g2_dfrbp_1 _8345_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net355),
    .D(_0513_),
    .Q_N(_3406_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[4][2] ));
 sg13g2_dfrbp_1 _8346_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net354),
    .D(_0514_),
    .Q_N(_3405_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[4][3] ));
 sg13g2_dfrbp_1 _8347_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net353),
    .D(_0515_),
    .Q_N(_3404_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[4][4] ));
 sg13g2_dfrbp_1 _8348_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net352),
    .D(_0516_),
    .Q_N(_3403_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[4][5] ));
 sg13g2_dfrbp_1 _8349_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net351),
    .D(_0517_),
    .Q_N(_3402_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[4][6] ));
 sg13g2_dfrbp_1 _8350_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net350),
    .D(_0518_),
    .Q_N(_3401_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[4][7] ));
 sg13g2_dfrbp_1 _8351_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net349),
    .D(_0519_),
    .Q_N(_3400_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[3][0] ));
 sg13g2_dfrbp_1 _8352_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net348),
    .D(_0520_),
    .Q_N(_3399_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[3][1] ));
 sg13g2_dfrbp_1 _8353_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net347),
    .D(_0521_),
    .Q_N(_3398_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[3][2] ));
 sg13g2_dfrbp_1 _8354_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net346),
    .D(_0522_),
    .Q_N(_3397_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[3][3] ));
 sg13g2_dfrbp_1 _8355_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net345),
    .D(_0523_),
    .Q_N(_3396_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[3][4] ));
 sg13g2_dfrbp_1 _8356_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net342),
    .D(_0524_),
    .Q_N(_3395_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[3][5] ));
 sg13g2_dfrbp_1 _8357_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net341),
    .D(_0525_),
    .Q_N(_3394_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[3][6] ));
 sg13g2_dfrbp_1 _8358_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net339),
    .D(_0526_),
    .Q_N(_3393_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[3][7] ));
 sg13g2_dfrbp_1 _8359_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net338),
    .D(_0527_),
    .Q_N(_3392_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[2][0] ));
 sg13g2_dfrbp_1 _8360_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net337),
    .D(_0528_),
    .Q_N(_3391_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[2][1] ));
 sg13g2_dfrbp_1 _8361_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net336),
    .D(_0529_),
    .Q_N(_3390_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[2][2] ));
 sg13g2_dfrbp_1 _8362_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net335),
    .D(_0530_),
    .Q_N(_3389_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[2][3] ));
 sg13g2_dfrbp_1 _8363_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net334),
    .D(_0531_),
    .Q_N(_3388_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[2][4] ));
 sg13g2_dfrbp_1 _8364_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net333),
    .D(_0532_),
    .Q_N(_3387_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[2][5] ));
 sg13g2_dfrbp_1 _8365_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net332),
    .D(_0533_),
    .Q_N(_3386_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[2][6] ));
 sg13g2_dfrbp_1 _8366_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net331),
    .D(_0534_),
    .Q_N(_3385_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[2][7] ));
 sg13g2_dfrbp_1 _8367_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net330),
    .D(_0535_),
    .Q_N(_3384_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[1][0] ));
 sg13g2_dfrbp_1 _8368_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net329),
    .D(_0536_),
    .Q_N(_3383_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[1][1] ));
 sg13g2_dfrbp_1 _8369_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net328),
    .D(_0537_),
    .Q_N(_3382_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[1][2] ));
 sg13g2_dfrbp_1 _8370_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net327),
    .D(_0538_),
    .Q_N(_3381_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[1][3] ));
 sg13g2_dfrbp_1 _8371_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net325),
    .D(_0539_),
    .Q_N(_3380_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[1][4] ));
 sg13g2_dfrbp_1 _8372_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net324),
    .D(_0540_),
    .Q_N(_3379_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[1][5] ));
 sg13g2_dfrbp_1 _8373_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net323),
    .D(_0541_),
    .Q_N(_3378_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[1][6] ));
 sg13g2_dfrbp_1 _8374_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net322),
    .D(_0542_),
    .Q_N(_3377_),
    .Q(\scl_fifo1.scl_memory0.physical_memory0.memory[1][7] ));
 sg13g2_dfrbp_1 _8375_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net321),
    .D(_0543_),
    .Q_N(_3376_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[9][0] ));
 sg13g2_dfrbp_1 _8376_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net320),
    .D(_0544_),
    .Q_N(_3375_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[9][1] ));
 sg13g2_dfrbp_1 _8377_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net319),
    .D(_0545_),
    .Q_N(_3374_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[9][2] ));
 sg13g2_dfrbp_1 _8378_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net318),
    .D(_0546_),
    .Q_N(_3373_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[9][3] ));
 sg13g2_dfrbp_1 _8379_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net317),
    .D(_0547_),
    .Q_N(_3372_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[9][4] ));
 sg13g2_dfrbp_1 _8380_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net316),
    .D(_0548_),
    .Q_N(_3371_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[9][5] ));
 sg13g2_dfrbp_1 _8381_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net315),
    .D(_0549_),
    .Q_N(_3370_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[9][6] ));
 sg13g2_dfrbp_1 _8382_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net314),
    .D(_0550_),
    .Q_N(_3369_),
    .Q(\scl_fifo0.scl_memory0.physical_memory0.memory[9][7] ));
 sg13g2_dfrbp_1 _8383_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net1530),
    .D(_0551_),
    .Q_N(_3368_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_decodenrzi0.n7166_q ));
 sg13g2_dfrbp_1 _8384_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net1529),
    .D(_0552_),
    .Q_N(_3367_),
    .Q(\usbfunction0.scl_usbgpiophy0.s_m_last ));
 sg13g2_dfrbp_1 _8385_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net313),
    .D(_0553_),
    .Q_N(_3366_),
    .Q(\s_m_status_linestate[0] ));
 sg13g2_dfrbp_1 _8386_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net312),
    .D(_0554_),
    .Q_N(_3365_),
    .Q(\s_m_status_linestate[1] ));
 sg13g2_dfrbp_1 _8387_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net1528),
    .D(_0555_),
    .Q_N(_0043_),
    .Q(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.in_in_valid ));
 sg13g2_dfrbp_1 _8388_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net1507),
    .D(\usbfunction0.scl_usbgpiophy0.scl_extendwidth0.scl_counter0.n7961_o[0] ),
    .Q_N(_0157_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_extendwidth0.scl_counter0.n7984_q[0] ));
 sg13g2_dfrbp_1 _8389_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net1507),
    .D(net1143),
    .Q_N(_3844_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_extendwidth0.scl_counter0.n7984_q[1] ));
 sg13g2_dfrbp_1 _8390_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net1507),
    .D(net609),
    .Q_N(_3364_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_extendwidth0.scl_counter0.n7984_q[2] ));
 sg13g2_dfrbp_1 _8391_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net1524),
    .D(_0556_),
    .Q_N(_0156_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_decodenrzi0.scl_counter0.n7944_q[0] ));
 sg13g2_dfrbp_1 _8392_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net1533),
    .D(_0557_),
    .Q_N(_3363_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_decodenrzi0.scl_counter0.n7944_q[1] ));
 sg13g2_dfrbp_1 _8393_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net1524),
    .D(_0558_),
    .Q_N(_0044_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_decodenrzi0.scl_counter0.n7944_q[2] ));
 sg13g2_dfrbp_1 _8394_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net311),
    .D(net724),
    .Q_N(_3362_),
    .Q(\usbfunction0.scl_usbgpiophy0.s_out_2[0] ));
 sg13g2_dfrbp_1 _8395_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net310),
    .D(net621),
    .Q_N(_3361_),
    .Q(\usbfunction0.scl_usbgpiophy0.s_out_2[1] ));
 sg13g2_dfrbp_1 _8396_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net309),
    .D(net634),
    .Q_N(_3360_),
    .Q(\usbfunction0.scl_usbgpiophy0.s_out_2[2] ));
 sg13g2_dfrbp_1 _8397_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net308),
    .D(net1010),
    .Q_N(_3359_),
    .Q(\usbfunction0.scl_usbgpiophy0.s_out_2[3] ));
 sg13g2_dfrbp_1 _8398_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net307),
    .D(net903),
    .Q_N(_3358_),
    .Q(\usbfunction0.scl_usbgpiophy0.s_out_2[4] ));
 sg13g2_dfrbp_1 _8399_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net306),
    .D(net1077),
    .Q_N(_3357_),
    .Q(\usbfunction0.scl_usbgpiophy0.s_out_2[5] ));
 sg13g2_dfrbp_1 _8400_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net305),
    .D(net618),
    .Q_N(_3356_),
    .Q(\usbfunction0.scl_usbgpiophy0.s_out_2[6] ));
 sg13g2_dfrbp_1 _8401_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net340),
    .D(net833),
    .Q_N(_3845_),
    .Q(\usbfunction0.scl_usbgpiophy0.s_out_2[7] ));
 sg13g2_dfrbp_1 _8402_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net1527),
    .D(net1714),
    .Q_N(_3355_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_addeopdeferred0.scl_eraselastbeat0.n8042_q ));
 sg13g2_dfrbp_1 _8403_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net1524),
    .D(net669),
    .Q_N(\usbfunction0.scl_usbgpiophy0.nrzi0.n7721_q ),
    .Q(_0173_));
 sg13g2_dfrbp_1 _8404_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net343),
    .D(_0568_),
    .Q_N(_3846_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_addeopdeferred0.scl_eraselastbeat0.n8041_q ));
 sg13g2_dfrbp_1 _8405_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net1528),
    .D(net1879),
    .Q_N(_3354_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_addeopdeferred0.n7349_q ));
 sg13g2_dfrbp_1 _8406_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net303),
    .D(_0569_),
    .Q_N(_3353_),
    .Q(\scl_bitbangengine0.n5920_q[9] ));
 sg13g2_dfrbp_1 _8407_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net344),
    .D(net1104),
    .Q_N(_0142_),
    .Q(\scl_bitbangengine0.n5920_q[10] ));
 sg13g2_dfrbp_1 _8408_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net1527),
    .D(net544),
    .Q_N(_0158_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.s_m_value[0] ));
 sg13g2_dfrbp_1 _8409_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net1527),
    .D(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.scl_counter0.n8088_o[1] ),
    .Q_N(_3847_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.s_m_value[1] ));
 sg13g2_dfrbp_1 _8410_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net1527),
    .D(net555),
    .Q_N(_0045_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.s_m_value[2] ));
 sg13g2_dfrbp_1 _8411_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net1526),
    .D(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.scl_counter0.n8128_o[0] ),
    .Q_N(_0159_),
    .Q(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.s_m_value[0] ));
 sg13g2_dfrbp_1 _8412_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net1526),
    .D(net1583),
    .Q_N(_0160_),
    .Q(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.s_m_value[1] ));
 sg13g2_dfrbp_1 _8413_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net1526),
    .D(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.scl_counter0.n8128_o[2] ),
    .Q_N(_3848_),
    .Q(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.s_m_value[2] ));
 sg13g2_dfrbp_1 _8414_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net1526),
    .D(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.scl_counter0.n8128_o[3] ),
    .Q_N(_3849_),
    .Q(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.s_m_value[3] ));
 sg13g2_dfrbp_1 _8415_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net377),
    .D(net1630),
    .Q_N(_3850_),
    .Q(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7656_q ));
 sg13g2_dfrbp_1 _8416_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net1527),
    .D(net1021),
    .Q_N(_3352_),
    .Q(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7657_q ));
 sg13g2_dfrbp_1 _8417_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net302),
    .D(net606),
    .Q_N(_3351_),
    .Q(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[0] ));
 sg13g2_dfrbp_1 _8418_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net301),
    .D(net1057),
    .Q_N(_3350_),
    .Q(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[1] ));
 sg13g2_dfrbp_1 _8419_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net300),
    .D(net1004),
    .Q_N(_3349_),
    .Q(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[2] ));
 sg13g2_dfrbp_1 _8420_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net299),
    .D(_0574_),
    .Q_N(_3348_),
    .Q(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[3] ));
 sg13g2_dfrbp_1 _8421_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net298),
    .D(net972),
    .Q_N(_3347_),
    .Q(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[4] ));
 sg13g2_dfrbp_1 _8422_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net297),
    .D(_0576_),
    .Q_N(_3346_),
    .Q(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[5] ));
 sg13g2_dfrbp_1 _8423_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net296),
    .D(net798),
    .Q_N(_3345_),
    .Q(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[6] ));
 sg13g2_dfrbp_1 _8424_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net295),
    .D(_0578_),
    .Q_N(_3344_),
    .Q(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[7] ));
 sg13g2_dfrbp_1 _8425_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net294),
    .D(net1001),
    .Q_N(_3343_),
    .Q(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[8] ));
 sg13g2_dfrbp_1 _8426_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net293),
    .D(_0580_),
    .Q_N(_3342_),
    .Q(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[9] ));
 sg13g2_dfrbp_1 _8427_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net292),
    .D(_0581_),
    .Q_N(_3341_),
    .Q(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[10] ));
 sg13g2_dfrbp_1 _8428_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net291),
    .D(_0582_),
    .Q_N(_3340_),
    .Q(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[11] ));
 sg13g2_dfrbp_1 _8429_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net290),
    .D(_0583_),
    .Q_N(_3339_),
    .Q(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[12] ));
 sg13g2_dfrbp_1 _8430_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net289),
    .D(_0584_),
    .Q_N(_3338_),
    .Q(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[13] ));
 sg13g2_dfrbp_1 _8431_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net288),
    .D(_0585_),
    .Q_N(_3337_),
    .Q(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[14] ));
 sg13g2_dfrbp_1 _8432_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net287),
    .D(_0586_),
    .Q_N(_3336_),
    .Q(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[15] ));
 sg13g2_dfrbp_1 _8433_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net1511),
    .D(net641),
    .Q_N(\scl_bitbangengine0.n5921_q[0] ),
    .Q(_0174_));
 sg13g2_dfrbp_1 _8434_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net1512),
    .D(_0588_),
    .Q_N(_3335_),
    .Q(\scl_bitbangengine0.n5921_q[1] ));
 sg13g2_dfrbp_1 _8435_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net1511),
    .D(_0589_),
    .Q_N(_0063_),
    .Q(\scl_bitbangengine0.n5921_q[2] ));
 sg13g2_dfrbp_1 _8436_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net1511),
    .D(_0590_),
    .Q_N(_3334_),
    .Q(\scl_bitbangengine0.n5921_q[3] ));
 sg13g2_dfrbp_1 _8437_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net1511),
    .D(_0591_),
    .Q_N(_3333_),
    .Q(\scl_bitbangengine0.n5921_q[4] ));
 sg13g2_dfrbp_1 _8438_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net1511),
    .D(_0592_),
    .Q_N(_3332_),
    .Q(\scl_bitbangengine0.n5921_q[5] ));
 sg13g2_dfrbp_1 _8439_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net1515),
    .D(_0593_),
    .Q_N(_0068_),
    .Q(\scl_bitbangengine0.n5921_q[6] ));
 sg13g2_dfrbp_1 _8440_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net1513),
    .D(_0594_),
    .Q_N(_3331_),
    .Q(\scl_bitbangengine0.n5921_q[7] ));
 sg13g2_dfrbp_1 _8441_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net285),
    .D(net1152),
    .Q_N(_3330_),
    .Q(\scl_bitbangengine0.n5920_q[11] ));
 sg13g2_dfrbp_1 _8442_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net284),
    .D(_0596_),
    .Q_N(_3329_),
    .Q(\scl_bitbangengine0.n5920_q[12] ));
 sg13g2_dfrbp_1 _8443_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net283),
    .D(_0597_),
    .Q_N(_3328_),
    .Q(\scl_bitbangengine0.n5920_q[13] ));
 sg13g2_dfrbp_1 _8444_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net282),
    .D(net882),
    .Q_N(_0143_),
    .Q(\scl_bitbangengine0.n5920_q[14] ));
 sg13g2_dfrbp_1 _8445_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net281),
    .D(net1572),
    .Q_N(_3327_),
    .Q(\scl_bitbangengine0.n5920_q[15] ));
 sg13g2_dfrbp_1 _8446_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net280),
    .D(_0600_),
    .Q_N(_3326_),
    .Q(\scl_bitbangengine0.n5920_q[16] ));
 sg13g2_dfrbp_1 _8447_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net279),
    .D(_0601_),
    .Q_N(_3325_),
    .Q(\scl_bitbangengine0.n5920_q[17] ));
 sg13g2_dfrbp_1 _8448_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net278),
    .D(net735),
    .Q_N(_0144_),
    .Q(\scl_bitbangengine0.n5920_q[18] ));
 sg13g2_dfrbp_1 _8449_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net378),
    .D(net1055),
    .Q_N(_3851_),
    .Q(\scl_bitbangengine0.n5920_q[19] ));
 sg13g2_dfrbp_1 _8450_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net1525),
    .D(\usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8195_o[0] ),
    .Q_N(_3852_),
    .Q(\usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8209_q[0] ));
 sg13g2_dfrbp_1 _8451_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net1525),
    .D(\usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8195_o[1] ),
    .Q_N(_3853_),
    .Q(\usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8209_q[1] ));
 sg13g2_dfrbp_1 _8452_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net1525),
    .D(net590),
    .Q_N(_3324_),
    .Q(\usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8209_q[2] ));
 sg13g2_dfrbp_1 _8453_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net1527),
    .D(net1763),
    .Q_N(_3323_),
    .Q(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7654_q[0] ));
 sg13g2_dfrbp_1 _8454_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net1527),
    .D(_0605_),
    .Q_N(_3854_),
    .Q(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7654_q[1] ));
 sg13g2_dfrbp_1 _8455_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net1525),
    .D(\usbfunction0.scl_usbgpiophy0.scl_pulseextender0.scl_counter0.n8221_o[0] ),
    .Q_N(_3855_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_pulseextender0.scl_counter0.n8243_q[0] ));
 sg13g2_dfrbp_1 _8456_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net1524),
    .D(\usbfunction0.scl_usbgpiophy0.scl_pulseextender0.scl_counter0.n8221_o[1] ),
    .Q_N(_3856_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_pulseextender0.scl_counter0.n8243_q[1] ));
 sg13g2_dfrbp_1 _8457_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net1525),
    .D(net1007),
    .Q_N(_3857_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_pulseextender0.n7750_q ));
 sg13g2_dfrbp_1 _8458_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net1524),
    .D(net547),
    .Q_N(_3858_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_pulseextender1.scl_counter0.n8282_q[0] ));
 sg13g2_dfrbp_1 _8459_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net1524),
    .D(\usbfunction0.scl_usbgpiophy0.scl_pulseextender1.scl_counter0.n8260_o[1] ),
    .Q_N(_3859_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_pulseextender1.scl_counter0.n8282_q[1] ));
 sg13g2_dfrbp_1 _8460_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net1524),
    .D(\usbfunction0.scl_usbgpiophy0.scl_pulseextender1.n7766_o ),
    .Q_N(_3322_),
    .Q(\usbfunction0.scl_usbgpiophy0.scl_pulseextender1.n7775_q ));
 sg13g2_dfrbp_1 _8461_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net277),
    .D(net768),
    .Q_N(_3321_),
    .Q(\s_m_packetdata_2_rewired[0] ));
 sg13g2_dfrbp_1 _8462_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net276),
    .D(net1560),
    .Q_N(_3320_),
    .Q(\s_m_packetdata_2_rewired[1] ));
 sg13g2_dfrbp_1 _8463_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net275),
    .D(net1579),
    .Q_N(_3319_),
    .Q(\s_m_packetdata_2_rewired[2] ));
 sg13g2_dfrbp_1 _8464_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net274),
    .D(net1676),
    .Q_N(_3318_),
    .Q(\s_m_packetdata_2_rewired[3] ));
 sg13g2_dfrbp_1 _8465_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net273),
    .D(net1633),
    .Q_N(_3317_),
    .Q(\s_m_packetdata_2_rewired[4] ));
 sg13g2_dfrbp_1 _8466_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net272),
    .D(_0611_),
    .Q_N(_3316_),
    .Q(\s_m_packetdata_2_rewired[5] ));
 sg13g2_dfrbp_1 _8467_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net271),
    .D(net1162),
    .Q_N(_3315_),
    .Q(\s_m_packetdata_2_rewired[6] ));
 sg13g2_dfrbp_1 _8468_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net270),
    .D(net1628),
    .Q_N(_3314_),
    .Q(\s_m_packetdata_2_rewired[7] ));
 sg13g2_dfrbp_1 _8469_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net269),
    .D(_0614_),
    .Q_N(_3313_),
    .Q(\s_m_packetdata_2_rewired[8] ));
 sg13g2_dfrbp_1 _8470_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net268),
    .D(_0615_),
    .Q_N(_3312_),
    .Q(\s_m_packetdata_2_rewired[9] ));
 sg13g2_dfrbp_1 _8471_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net267),
    .D(_0616_),
    .Q_N(_3311_),
    .Q(\s_m_packetdata_2_rewired[10] ));
 sg13g2_dfrbp_1 _8472_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net266),
    .D(net1831),
    .Q_N(_3310_),
    .Q(\s_m_packetdata_2_rewired[11] ));
 sg13g2_dfrbp_1 _8473_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net265),
    .D(net1740),
    .Q_N(_3309_),
    .Q(\s_m_packetdata_2_rewired[12] ));
 sg13g2_dfrbp_1 _8474_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net264),
    .D(_0619_),
    .Q_N(_3308_),
    .Q(\s_m_packetdata_2_rewired[13] ));
 sg13g2_dfrbp_1 _8475_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net263),
    .D(_0620_),
    .Q_N(_3307_),
    .Q(\s_m_packetdata_2_rewired[14] ));
 sg13g2_dfrbp_1 _8476_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net262),
    .D(net1566),
    .Q_N(_3306_),
    .Q(\s_m_packetdata_2_rewired[15] ));
 sg13g2_dfrbp_1 _8477_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net261),
    .D(_0622_),
    .Q_N(_3305_),
    .Q(s_m_packetdata_2_bit_16));
 sg13g2_dfrbp_1 _8478_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net260),
    .D(net1689),
    .Q_N(_3304_),
    .Q(s_m_packetdata_2_bit_17));
 sg13g2_dfrbp_1 _8479_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net259),
    .D(_0624_),
    .Q_N(_3303_),
    .Q(\s_m_packetdata_2_rewired[18] ));
 sg13g2_dfrbp_1 _8480_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net258),
    .D(net1784),
    .Q_N(_3302_),
    .Q(\s_m_packetdata_2_rewired[19] ));
 sg13g2_dfrbp_1 _8481_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net257),
    .D(_0626_),
    .Q_N(_3301_),
    .Q(\s_m_packetdata_2_rewired[20] ));
 sg13g2_dfrbp_1 _8482_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net256),
    .D(_0627_),
    .Q_N(_3300_),
    .Q(\s_m_packetdata_2_rewired[21] ));
 sg13g2_dfrbp_1 _8483_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net255),
    .D(_0628_),
    .Q_N(_3299_),
    .Q(\s_m_packetdata_2_rewired[22] ));
 sg13g2_dfrbp_1 _8484_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net254),
    .D(_0629_),
    .Q_N(_3298_),
    .Q(\s_m_packetdata_2_rewired[23] ));
 sg13g2_dfrbp_1 _8485_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net253),
    .D(net975),
    .Q_N(_3297_),
    .Q(\usbfunction0.n2481_o[16] ));
 sg13g2_dfrbp_1 _8486_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net252),
    .D(net967),
    .Q_N(_3296_),
    .Q(\usbfunction0.n2481_o[17] ));
 sg13g2_dfrbp_1 _8487_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net251),
    .D(_0632_),
    .Q_N(_3295_),
    .Q(\usbfunction0.n2481_o[18] ));
 sg13g2_dfrbp_1 _8488_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net250),
    .D(net1053),
    .Q_N(_3294_),
    .Q(\usbfunction0.n2481_o[19] ));
 sg13g2_dfrbp_1 _8489_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net249),
    .D(net1156),
    .Q_N(_3293_),
    .Q(\usbfunction0.n2481_o[20] ));
 sg13g2_dfrbp_1 _8490_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net248),
    .D(_0635_),
    .Q_N(_3292_),
    .Q(\usbfunction0.n2481_o[21] ));
 sg13g2_dfrbp_1 _8491_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net247),
    .D(net1598),
    .Q_N(_3291_),
    .Q(\usbfunction0.n2481_o[22] ));
 sg13g2_dfrbp_1 _8492_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net246),
    .D(_0637_),
    .Q_N(_3290_),
    .Q(\usbfunction0.n2481_o[23] ));
 sg13g2_dfrbp_1 _8493_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net245),
    .D(_0638_),
    .Q_N(_3289_),
    .Q(\usbfunction0.n2481_o[24] ));
 sg13g2_dfrbp_1 _8494_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net244),
    .D(_0639_),
    .Q_N(_3288_),
    .Q(\usbfunction0.n2481_o[25] ));
 sg13g2_dfrbp_1 _8495_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net243),
    .D(net791),
    .Q_N(_3287_),
    .Q(\usbfunction0.n2481_o[26] ));
 sg13g2_dfrbp_1 _8496_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net242),
    .D(_0641_),
    .Q_N(_3286_),
    .Q(\usbfunction0.n2481_o[27] ));
 sg13g2_dfrbp_1 _8497_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net241),
    .D(_0642_),
    .Q_N(_3285_),
    .Q(\usbfunction0.n2481_o[28] ));
 sg13g2_dfrbp_1 _8498_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net240),
    .D(net1094),
    .Q_N(_3284_),
    .Q(\usbfunction0.n2481_o[29] ));
 sg13g2_dfrbp_1 _8499_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net239),
    .D(net1624),
    .Q_N(_3283_),
    .Q(\usbfunction0.n2481_o[30] ));
 sg13g2_dfrbp_1 _8500_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net238),
    .D(_0645_),
    .Q_N(_3282_),
    .Q(\usbfunction0.n2098_o ));
 sg13g2_dfrbp_1 _8501_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net237),
    .D(net1616),
    .Q_N(_3281_),
    .Q(\usbfunction0.n2481_o[32] ));
 sg13g2_dfrbp_1 _8502_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net236),
    .D(_0647_),
    .Q_N(_3280_),
    .Q(\usbfunction0.n2481_o[33] ));
 sg13g2_dfrbp_1 _8503_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net235),
    .D(_0648_),
    .Q_N(_3279_),
    .Q(\usbfunction0.n2481_o[34] ));
 sg13g2_dfrbp_1 _8504_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net234),
    .D(_0649_),
    .Q_N(_3278_),
    .Q(\usbfunction0.n2481_o[35] ));
 sg13g2_dfrbp_1 _8505_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net233),
    .D(net1085),
    .Q_N(_3277_),
    .Q(\usbfunction0.n2481_o[36] ));
 sg13g2_dfrbp_1 _8506_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net232),
    .D(net1636),
    .Q_N(_3276_),
    .Q(\usbfunction0.n2481_o[37] ));
 sg13g2_dfrbp_1 _8507_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net231),
    .D(net1686),
    .Q_N(_3275_),
    .Q(\usbfunction0.n2481_o[38] ));
 sg13g2_dfrbp_1 _8508_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net230),
    .D(_0653_),
    .Q_N(_3274_),
    .Q(\usbfunction0.n2481_o[39] ));
 sg13g2_dfrbp_1 _8509_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net229),
    .D(_0654_),
    .Q_N(_3273_),
    .Q(\usbfunction0.n1583_o[0] ));
 sg13g2_dfrbp_1 _8510_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net228),
    .D(_0655_),
    .Q_N(_0030_),
    .Q(\usbfunction0.n1583_o[1] ));
 sg13g2_dfrbp_1 _8511_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net227),
    .D(_0656_),
    .Q_N(_0031_),
    .Q(\usbfunction0.n1583_o[2] ));
 sg13g2_dfrbp_1 _8512_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net226),
    .D(net1019),
    .Q_N(_0032_),
    .Q(\usbfunction0.n1583_o[3] ));
 sg13g2_dfrbp_1 _8513_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net225),
    .D(net1051),
    .Q_N(_3272_),
    .Q(\usbfunction0.n1583_o[4] ));
 sg13g2_dfrbp_1 _8514_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net223),
    .D(net1593),
    .Q_N(_0033_),
    .Q(\usbfunction0.n1583_o[5] ));
 sg13g2_dfrbp_1 _8515_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net205),
    .D(net1160),
    .Q_N(_0034_),
    .Q(\usbfunction0.n1583_o[6] ));
 sg13g2_dfrbp_1 _8516_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net193),
    .D(net874),
    .Q_N(_0086_),
    .Q(\usbfunction0.n1360_o[0] ));
 sg13g2_dfrbp_1 _8517_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net189),
    .D(_0662_),
    .Q_N(_3271_),
    .Q(\usbfunction0.n1360_o[1] ));
 sg13g2_dfrbp_1 _8518_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net187),
    .D(_0663_),
    .Q_N(_3270_),
    .Q(\usbfunction0.n1360_o[2] ));
 sg13g2_dfrbp_1 _8519_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net185),
    .D(_0664_),
    .Q_N(_3269_),
    .Q(\usbfunction0.n1360_o[3] ));
 sg13g2_dfrbp_1 _8520_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net182),
    .D(_0665_),
    .Q_N(_3268_),
    .Q(\usbfunction0.n2481_o[51] ));
 sg13g2_dfrbp_1 _8521_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net179),
    .D(_0666_),
    .Q_N(_3267_),
    .Q(\usbfunction0.n2481_o[52] ));
 sg13g2_dfrbp_1 _8522_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net176),
    .D(_0667_),
    .Q_N(_3266_),
    .Q(\usbfunction0.n2481_o[53] ));
 sg13g2_dfrbp_1 _8523_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net175),
    .D(_0668_),
    .Q_N(_3265_),
    .Q(\usbfunction0.n2481_o[54] ));
 sg13g2_dfrbp_1 _8524_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net445),
    .D(_0669_),
    .Q_N(_3860_),
    .Q(\usbfunction0.n2481_o[55] ));
 sg13g2_dfrbp_1 _8525_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net446),
    .D(net530),
    .Q_N(_3861_),
    .Q(\usbfunction0.n2630_q ));
 sg13g2_dfrbp_1 _8526_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net447),
    .D(\s_m_pushdata_endpoint[0] ),
    .Q_N(_3862_),
    .Q(\usbfunction0.n2642_q[0] ));
 sg13g2_dfrbp_1 _8527_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net448),
    .D(net1043),
    .Q_N(_3863_),
    .Q(\usbfunction0.n2642_q[1] ));
 sg13g2_dfrbp_1 _8528_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net449),
    .D(\s_m_pushdata_endpoint[2] ),
    .Q_N(_3864_),
    .Q(\usbfunction0.n2642_q[2] ));
 sg13g2_dfrbp_1 _8529_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net450),
    .D(\s_m_pushdata_endpoint[3] ),
    .Q_N(_3865_),
    .Q(\usbfunction0.n2642_q[3] ));
 sg13g2_dfrbp_1 _8530_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net451),
    .D(\usbfunction0.n1630_o[0] ),
    .Q_N(_3866_),
    .Q(\usbfunction0.n2644_q[0] ));
 sg13g2_dfrbp_1 _8531_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net452),
    .D(\usbfunction0.n1630_o[1] ),
    .Q_N(_3867_),
    .Q(\usbfunction0.n2644_q[1] ));
 sg13g2_dfrbp_1 _8532_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net453),
    .D(\usbfunction0.n1630_o[2] ),
    .Q_N(_3868_),
    .Q(\usbfunction0.n2644_q[2] ));
 sg13g2_dfrbp_1 _8533_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net454),
    .D(\usbfunction0.n1630_o[3] ),
    .Q_N(_3869_),
    .Q(\usbfunction0.n2644_q[3] ));
 sg13g2_dfrbp_1 _8534_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net455),
    .D(\usbfunction0.n1630_o[4] ),
    .Q_N(_3870_),
    .Q(\usbfunction0.n2644_q[4] ));
 sg13g2_dfrbp_1 _8535_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net456),
    .D(\usbfunction0.n1630_o[5] ),
    .Q_N(_3871_),
    .Q(\usbfunction0.n2644_q[5] ));
 sg13g2_dfrbp_1 _8536_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net457),
    .D(\usbfunction0.n1630_o[6] ),
    .Q_N(_3872_),
    .Q(\usbfunction0.n2644_q[6] ));
 sg13g2_dfrbp_1 _8537_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net458),
    .D(\usbfunction0.n1630_o[7] ),
    .Q_N(_3873_),
    .Q(\usbfunction0.n2644_q[7] ));
 sg13g2_dfrbp_1 _8538_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net459),
    .D(\usbfunction0.n1630_o[8] ),
    .Q_N(_3874_),
    .Q(\usbfunction0.n2644_q[8] ));
 sg13g2_dfrbp_1 _8539_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net460),
    .D(\usbfunction0.n1630_o[9] ),
    .Q_N(_3875_),
    .Q(\usbfunction0.n2644_q[9] ));
 sg13g2_dfrbp_1 _8540_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net461),
    .D(\usbfunction0.n1630_o[10] ),
    .Q_N(_3876_),
    .Q(\usbfunction0.n2644_q[10] ));
 sg13g2_dfrbp_1 _8541_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net462),
    .D(\usbfunction0.n1630_o[11] ),
    .Q_N(_3877_),
    .Q(\usbfunction0.n2644_q[11] ));
 sg13g2_dfrbp_1 _8542_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net463),
    .D(\usbfunction0.n1630_o[12] ),
    .Q_N(_3878_),
    .Q(\usbfunction0.n2644_q[12] ));
 sg13g2_dfrbp_1 _8543_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net464),
    .D(\usbfunction0.n1630_o[13] ),
    .Q_N(_3879_),
    .Q(\usbfunction0.n2644_q[13] ));
 sg13g2_dfrbp_1 _8544_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net465),
    .D(\usbfunction0.n1630_o[14] ),
    .Q_N(_3880_),
    .Q(\usbfunction0.n2644_q[14] ));
 sg13g2_dfrbp_1 _8545_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net466),
    .D(\usbfunction0.n1630_o[15] ),
    .Q_N(_3881_),
    .Q(\usbfunction0.n2644_q[15] ));
 sg13g2_dfrbp_1 _8546_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net1542),
    .D(\usbfunction0.n1083_o[0] ),
    .Q_N(_3882_),
    .Q(\usbfunction0.functionreset0.in_unnamed_3[0] ));
 sg13g2_dfrbp_1 _8547_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net1548),
    .D(net1791),
    .Q_N(_3883_),
    .Q(\usbfunction0.functionreset0.in_unnamed_3[1] ));
 sg13g2_dfrbp_1 _8548_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net1548),
    .D(\usbfunction0.n1083_o[2] ),
    .Q_N(_3884_),
    .Q(\usbfunction0.functionreset0.in_unnamed_3[2] ));
 sg13g2_dfrbp_1 _8549_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net1548),
    .D(net1844),
    .Q_N(_3885_),
    .Q(\usbfunction0.functionreset0.in_unnamed_3[3] ));
 sg13g2_dfrbp_1 _8550_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net1542),
    .D(net1760),
    .Q_N(_3886_),
    .Q(\usbfunction0.functionreset0.in_unnamed_3[4] ));
 sg13g2_dfrbp_1 _8551_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net1548),
    .D(net1596),
    .Q_N(_3887_),
    .Q(\usbfunction0.functionreset0.in_unnamed_3[5] ));
 sg13g2_dfrbp_1 _8552_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net1548),
    .D(\usbfunction0.n1083_o[6] ),
    .Q_N(_3888_),
    .Q(\usbfunction0.functionreset0.in_unnamed_3[6] ));
 sg13g2_dfrbp_1 _8553_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net467),
    .D(net536),
    .Q_N(_3889_),
    .Q(\s_m_pushdata_data[0] ));
 sg13g2_dfrbp_1 _8554_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net468),
    .D(net540),
    .Q_N(_3890_),
    .Q(\s_m_pushdata_data[1] ));
 sg13g2_dfrbp_1 _8555_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net469),
    .D(net532),
    .Q_N(_3891_),
    .Q(\s_m_pushdata_data[2] ));
 sg13g2_dfrbp_1 _8556_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net470),
    .D(net534),
    .Q_N(_3892_),
    .Q(\s_m_pushdata_data[3] ));
 sg13g2_dfrbp_1 _8557_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net471),
    .D(net533),
    .Q_N(_3893_),
    .Q(\s_m_pushdata_data[4] ));
 sg13g2_dfrbp_1 _8558_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net472),
    .D(net531),
    .Q_N(_3894_),
    .Q(\s_m_pushdata_data[5] ));
 sg13g2_dfrbp_1 _8559_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net473),
    .D(net535),
    .Q_N(_0061_),
    .Q(\s_m_pushdata_data[6] ));
 sg13g2_dfrbp_1 _8560_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net474),
    .D(\usbfunction0.s_m_rx_data[7] ),
    .Q_N(_3895_),
    .Q(\s_m_pushdata_data[7] ));
 sg13g2_dfrbp_1 _8561_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net1539),
    .D(\usbfunction0.n1189_o[0] ),
    .Q_N(_3896_),
    .Q(\usbfunction0.functionreset0.in_unnamed_2[0] ));
 sg13g2_dfrbp_1 _8562_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net1539),
    .D(\usbfunction0.n1189_o[1] ),
    .Q_N(_3897_),
    .Q(\usbfunction0.functionreset0.in_unnamed_2[1] ));
 sg13g2_dfrbp_1 _8563_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net1538),
    .D(\usbfunction0.n1189_o[2] ),
    .Q_N(_3898_),
    .Q(\usbfunction0.functionreset0.in_unnamed_2[2] ));
 sg13g2_dfrbp_1 _8564_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net1540),
    .D(\usbfunction0.n1189_o[3] ),
    .Q_N(_3264_),
    .Q(\usbfunction0.functionreset0.in_unnamed_2[3] ));
 sg13g2_dfrbp_1 _8565_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net1538),
    .D(net1743),
    .Q_N(_0117_),
    .Q(\usbfunction0.n2636_q ));
 sg13g2_dfrbp_1 _8566_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net1506),
    .D(\usbfunction0.n2254_o ),
    .Q_N(_3899_),
    .Q(\usbfunction0.n2648_q[0] ));
 sg13g2_dfrbp_1 _8567_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net1536),
    .D(\usbfunction0.n2257_o[1] ),
    .Q_N(_0102_),
    .Q(\usbfunction0.n2648_q[1] ));
 sg13g2_dfrbp_1 _8568_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net1536),
    .D(\usbfunction0.n2257_o[2] ),
    .Q_N(_0103_),
    .Q(\usbfunction0.n2648_q[2] ));
 sg13g2_dfrbp_1 _8569_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net1537),
    .D(\usbfunction0.n2257_o[3] ),
    .Q_N(_0104_),
    .Q(\usbfunction0.n2648_q[3] ));
 sg13g2_dfrbp_1 _8570_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net1506),
    .D(\usbfunction0.n2257_o[4] ),
    .Q_N(_0105_),
    .Q(\usbfunction0.n2648_q[4] ));
 sg13g2_dfrbp_1 _8571_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net1506),
    .D(\usbfunction0.n2257_o[5] ),
    .Q_N(_0106_),
    .Q(\usbfunction0.n2648_q[5] ));
 sg13g2_dfrbp_1 _8572_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net1536),
    .D(\usbfunction0.n2257_o[6] ),
    .Q_N(_0107_),
    .Q(\usbfunction0.n2648_q[6] ));
 sg13g2_dfrbp_1 _8573_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net1536),
    .D(\usbfunction0.n2257_o[7] ),
    .Q_N(_0108_),
    .Q(\usbfunction0.n2648_q[7] ));
 sg13g2_dfrbp_1 _8574_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net1536),
    .D(\usbfunction0.n2257_o[8] ),
    .Q_N(_0109_),
    .Q(\usbfunction0.n2648_q[8] ));
 sg13g2_dfrbp_1 _8575_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net1536),
    .D(\usbfunction0.n2257_o[9] ),
    .Q_N(_0110_),
    .Q(\usbfunction0.n2648_q[9] ));
 sg13g2_dfrbp_1 _8576_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net1506),
    .D(\usbfunction0.n2257_o[10] ),
    .Q_N(_0111_),
    .Q(\usbfunction0.n2648_q[10] ));
 sg13g2_dfrbp_1 _8577_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net1506),
    .D(\usbfunction0.n2257_o[11] ),
    .Q_N(_0112_),
    .Q(\usbfunction0.n2648_q[11] ));
 sg13g2_dfrbp_1 _8578_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net1537),
    .D(\usbfunction0.n2257_o[12] ),
    .Q_N(_0113_),
    .Q(\usbfunction0.n2648_q[12] ));
 sg13g2_dfrbp_1 _8579_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net1505),
    .D(\usbfunction0.n2257_o[13] ),
    .Q_N(_0114_),
    .Q(\usbfunction0.n2648_q[13] ));
 sg13g2_dfrbp_1 _8580_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net1505),
    .D(\usbfunction0.n2257_o[14] ),
    .Q_N(_0115_),
    .Q(\usbfunction0.n2648_q[14] ));
 sg13g2_dfrbp_1 _8581_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net1505),
    .D(\usbfunction0.n2257_o[15] ),
    .Q_N(_0116_),
    .Q(\usbfunction0.n2648_q[15] ));
 sg13g2_dfrbp_1 _8582_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net1508),
    .D(net1097),
    .Q_N(_0036_),
    .Q(\usbfunction0.n2628_q ));
 sg13g2_dfrbp_1 _8583_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net476),
    .D(\usbfunction0.n2477_o[0] ),
    .Q_N(_3900_),
    .Q(\usbfunction0.n2649_q[0] ));
 sg13g2_dfrbp_1 _8584_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net477),
    .D(\usbfunction0.n2477_o[1] ),
    .Q_N(_0095_),
    .Q(\usbfunction0.n2649_q[1] ));
 sg13g2_dfrbp_1 _8585_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net478),
    .D(\usbfunction0.n2477_o[2] ),
    .Q_N(_0096_),
    .Q(\usbfunction0.n2649_q[2] ));
 sg13g2_dfrbp_1 _8586_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net479),
    .D(\usbfunction0.n2477_o[3] ),
    .Q_N(_0097_),
    .Q(\usbfunction0.n2649_q[3] ));
 sg13g2_dfrbp_1 _8587_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net480),
    .D(\usbfunction0.n2477_o[4] ),
    .Q_N(_0098_),
    .Q(\usbfunction0.n2649_q[4] ));
 sg13g2_dfrbp_1 _8588_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net481),
    .D(\usbfunction0.n2477_o[5] ),
    .Q_N(_0099_),
    .Q(\usbfunction0.n2649_q[5] ));
 sg13g2_dfrbp_1 _8589_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net482),
    .D(\usbfunction0.n2477_o[6] ),
    .Q_N(_0100_),
    .Q(\usbfunction0.n2649_q[6] ));
 sg13g2_dfrbp_1 _8590_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net483),
    .D(\usbfunction0.n2477_o[7] ),
    .Q_N(_0101_),
    .Q(\usbfunction0.n2649_q[7] ));
 sg13g2_dfrbp_1 _8591_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net484),
    .D(\usbfunction0.n2480_o[0] ),
    .Q_N(_3901_),
    .Q(\usbfunction0.n2650_q[0] ));
 sg13g2_dfrbp_1 _8592_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net485),
    .D(\usbfunction0.n2480_o[1] ),
    .Q_N(_0094_),
    .Q(\usbfunction0.n2650_q[1] ));
 sg13g2_dfrbp_1 _8593_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net486),
    .D(\usbfunction0.n2480_o[2] ),
    .Q_N(_0092_),
    .Q(\usbfunction0.n2650_q[2] ));
 sg13g2_dfrbp_1 _8594_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net487),
    .D(\usbfunction0.n2480_o[3] ),
    .Q_N(_0091_),
    .Q(\usbfunction0.n2650_q[3] ));
 sg13g2_dfrbp_1 _8595_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net488),
    .D(\usbfunction0.n2480_o[4] ),
    .Q_N(_0090_),
    .Q(\usbfunction0.n2650_q[4] ));
 sg13g2_dfrbp_1 _8596_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net489),
    .D(\usbfunction0.n2480_o[5] ),
    .Q_N(_0089_),
    .Q(\usbfunction0.n2650_q[5] ));
 sg13g2_dfrbp_1 _8597_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net490),
    .D(\usbfunction0.n2480_o[6] ),
    .Q_N(_0088_),
    .Q(\usbfunction0.n2650_q[6] ));
 sg13g2_dfrbp_1 _8598_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net491),
    .D(\usbfunction0.n2480_o[7] ),
    .Q_N(_0087_),
    .Q(\usbfunction0.n2650_q[7] ));
 sg13g2_dfrbp_1 _8599_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net492),
    .D(\usbfunction0.n1101_o[0] ),
    .Q_N(_3902_),
    .Q(\usbfunction0.n2651_q[0] ));
 sg13g2_dfrbp_1 _8600_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net493),
    .D(\usbfunction0.n1101_o[1] ),
    .Q_N(_3903_),
    .Q(\usbfunction0.n2651_q[1] ));
 sg13g2_dfrbp_1 _8601_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net494),
    .D(\usbfunction0.n1101_o[2] ),
    .Q_N(_3904_),
    .Q(\usbfunction0.n2651_q[2] ));
 sg13g2_dfrbp_1 _8602_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net495),
    .D(\usbfunction0.n1101_o[3] ),
    .Q_N(_3905_),
    .Q(\usbfunction0.n2651_q[3] ));
 sg13g2_dfrbp_1 _8603_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net496),
    .D(\usbfunction0.n1101_o[4] ),
    .Q_N(_3906_),
    .Q(\usbfunction0.n2651_q[4] ));
 sg13g2_dfrbp_1 _8604_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net497),
    .D(\usbfunction0.n1101_o[5] ),
    .Q_N(_3907_),
    .Q(\usbfunction0.n2651_q[5] ));
 sg13g2_dfrbp_1 _8605_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net498),
    .D(\usbfunction0.n1101_o[6] ),
    .Q_N(_3908_),
    .Q(\usbfunction0.n2651_q[6] ));
 sg13g2_dfrbp_1 _8606_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net499),
    .D(\usbfunction0.n1101_o[7] ),
    .Q_N(_3909_),
    .Q(\usbfunction0.n2651_q[7] ));
 sg13g2_dfrbp_1 _8607_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net500),
    .D(\usbfunction0.n2353_o[0] ),
    .Q_N(_0085_),
    .Q(\usbfunction0.n2652_q[0] ));
 sg13g2_dfrbp_1 _8608_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net501),
    .D(\usbfunction0.n2353_o[1] ),
    .Q_N(_0093_),
    .Q(\usbfunction0.n2652_q[1] ));
 sg13g2_dfrbp_1 _8609_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net502),
    .D(\usbfunction0.n2353_o[2] ),
    .Q_N(_3910_),
    .Q(\usbfunction0.n2652_q[2] ));
 sg13g2_dfrbp_1 _8610_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net503),
    .D(\usbfunction0.n2353_o[3] ),
    .Q_N(_3911_),
    .Q(\usbfunction0.n2652_q[3] ));
 sg13g2_dfrbp_1 _8611_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net504),
    .D(\usbfunction0.n2353_o[4] ),
    .Q_N(_3912_),
    .Q(\usbfunction0.n2652_q[4] ));
 sg13g2_dfrbp_1 _8612_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net505),
    .D(\usbfunction0.n2353_o[5] ),
    .Q_N(_3913_),
    .Q(\usbfunction0.n2652_q[5] ));
 sg13g2_dfrbp_1 _8613_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net506),
    .D(\usbfunction0.n2353_o[6] ),
    .Q_N(_3914_),
    .Q(\usbfunction0.n2652_q[6] ));
 sg13g2_dfrbp_1 _8614_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net507),
    .D(\usbfunction0.n2353_o[7] ),
    .Q_N(_3915_),
    .Q(\usbfunction0.n2652_q[7] ));
 sg13g2_dfrbp_1 _8615_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net508),
    .D(\usbfunction0.n2433_o[0] ),
    .Q_N(_3916_),
    .Q(\usbfunction0.n2653_q[0] ));
 sg13g2_dfrbp_1 _8616_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net509),
    .D(net898),
    .Q_N(_0047_),
    .Q(\usbfunction0.n1687_o[0] ));
 sg13g2_dfrbp_1 _8617_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net510),
    .D(net1029),
    .Q_N(_0048_),
    .Q(\usbfunction0.n1687_o[1] ));
 sg13g2_dfrbp_1 _8618_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net511),
    .D(net1128),
    .Q_N(_0049_),
    .Q(\usbfunction0.n1687_o[2] ));
 sg13g2_dfrbp_1 _8619_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net512),
    .D(net927),
    .Q_N(_0050_),
    .Q(\usbfunction0.n1687_o[3] ));
 sg13g2_dfrbp_1 _8620_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net513),
    .D(net901),
    .Q_N(_0051_),
    .Q(\usbfunction0.n1687_o[4] ));
 sg13g2_dfrbp_1 _8621_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net514),
    .D(net777),
    .Q_N(_0052_),
    .Q(\usbfunction0.n1687_o[5] ));
 sg13g2_dfrbp_1 _8622_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net515),
    .D(net762),
    .Q_N(_0053_),
    .Q(\usbfunction0.n1687_o[6] ));
 sg13g2_dfrbp_1 _8623_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net516),
    .D(net775),
    .Q_N(_0054_),
    .Q(\usbfunction0.n1687_o[7] ));
 sg13g2_dfrbp_1 _8624_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net517),
    .D(net632),
    .Q_N(_0055_),
    .Q(\usbfunction0.n1687_o[8] ));
 sg13g2_dfrbp_1 _8625_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net518),
    .D(net772),
    .Q_N(_0056_),
    .Q(\usbfunction0.n1687_o[9] ));
 sg13g2_dfrbp_1 _8626_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net519),
    .D(net910),
    .Q_N(_0057_),
    .Q(\usbfunction0.n1687_o[10] ));
 sg13g2_dfrbp_1 _8627_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net520),
    .D(net940),
    .Q_N(_0058_),
    .Q(\usbfunction0.n1687_o[11] ));
 sg13g2_dfrbp_1 _8628_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net521),
    .D(net693),
    .Q_N(_0059_),
    .Q(\usbfunction0.n1687_o[12] ));
 sg13g2_dfrbp_1 _8629_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net527),
    .D(net818),
    .Q_N(_0060_),
    .Q(\usbfunction0.n1687_o[13] ));
 sg13g2_dfrbp_1 _8630_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net173),
    .D(net625),
    .Q_N(_0046_),
    .Q(\usbfunction0.n1687_o[14] ));
 sg13g2_dfrbp_1 _8631_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net171),
    .D(net1699),
    .Q_N(_3263_),
    .Q(\usbfunction0.n1581_o[0] ));
 sg13g2_dfrbp_1 _8632_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net169),
    .D(net1808),
    .Q_N(_3262_),
    .Q(\usbfunction0.n1581_o[1] ));
 sg13g2_dfrbp_1 _8633_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net167),
    .D(net1704),
    .Q_N(_3261_),
    .Q(\usbfunction0.n1359_o[0] ));
 sg13g2_dfrbp_1 _8634_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net526),
    .D(_0674_),
    .Q_N(_3260_),
    .Q(\usbfunction0.n1359_o[1] ));
 sg13g2_dfrbp_1 _8635_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net304),
    .D(net551),
    .Q_N(\usbfunction0.n2334_o[0] ),
    .Q(\usbfunction0.n2313_o[0] ));
 sg13g2_dfrbp_1 _8636_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net286),
    .D(net1819),
    .Q_N(_3259_),
    .Q(\usbfunction0.n2313_o[1] ));
 sg13g2_dfrbp_1 _8637_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net170),
    .D(net1734),
    .Q_N(_3258_),
    .Q(\usbfunction0.n2313_o[2] ));
 sg13g2_dfrbp_1 _8638_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net28),
    .D(net1856),
    .Q_N(_3257_),
    .Q(\usbfunction0.n2313_o[3] ));
 sg13g2_dfrbp_1 _8639_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net1533),
    .D(net1718),
    .Q_N(_0082_),
    .Q(\scl_uartrx0.s_m_value[0] ));
 sg13g2_dfrbp_1 _8640_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net1533),
    .D(net1158),
    .Q_N(_3256_),
    .Q(\scl_uartrx0.s_m_value[1] ));
 sg13g2_dfrbp_1 _8641_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net1533),
    .D(net1568),
    .Q_N(_0081_),
    .Q(\scl_uartrx0.s_m_value[2] ));
 sg13g2_dfrbp_1 _8642_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net1540),
    .D(\usbfunction0.n665_o[0] ),
    .Q_N(_3917_),
    .Q(\usbfunction0.functionreset0.in_unnamed[0] ));
 sg13g2_dfrbp_1 _8643_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net1537),
    .D(net1828),
    .Q_N(_3918_),
    .Q(\usbfunction0.functionreset0.in_unnamed[1] ));
 sg13g2_dfrbp_1 _8644_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net1537),
    .D(\usbfunction0.n665_o[2] ),
    .Q_N(_3919_),
    .Q(\usbfunction0.functionreset0.in_unnamed[2] ));
 sg13g2_dfrbp_1 _8645_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net1540),
    .D(net1884),
    .Q_N(_3920_),
    .Q(\usbfunction0.functionreset0.in_unnamed[3] ));
 sg13g2_dfrbp_1 _8646_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net1537),
    .D(net1847),
    .Q_N(_3921_),
    .Q(\usbfunction0.functionreset0.in_unnamed[4] ));
 sg13g2_dfrbp_1 _8647_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net1536),
    .D(net1887),
    .Q_N(_3922_),
    .Q(\usbfunction0.functionreset0.in_unnamed[5] ));
 sg13g2_dfrbp_1 _8648_ (.CLK(clknet_leaf_89_clk_regs),
    .RESET_B(net1536),
    .D(net1825),
    .Q_N(_3923_),
    .Q(\usbfunction0.functionreset0.in_unnamed[6] ));
 sg13g2_dfrbp_1 _8649_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net168),
    .D(\usbfunction0.s_m_rx_error ),
    .Q_N(_0035_),
    .Q(\usbfunction0.n2627_q ));
 sg13g2_tiehi _7832__18 (.L_HI(net18));
 sg13g2_tiehi _7833__19 (.L_HI(net19));
 sg13g2_tiehi _7834__20 (.L_HI(net20));
 sg13g2_tiehi _7835__21 (.L_HI(net21));
 sg13g2_tiehi _7836__22 (.L_HI(net22));
 sg13g2_tiehi _7837__23 (.L_HI(net23));
 sg13g2_tiehi _7838__24 (.L_HI(net24));
 sg13g2_tiehi _8233__25 (.L_HI(net25));
 sg13g2_tiehi _8232__26 (.L_HI(net26));
 sg13g2_tiehi _7839__27 (.L_HI(net27));
 sg13g2_tiehi _8638__28 (.L_HI(net28));
 sg13g2_tiehi _7851__29 (.L_HI(net29));
 sg13g2_tiehi _8213__30 (.L_HI(net30));
 sg13g2_tiehi _7852__31 (.L_HI(net31));
 sg13g2_tiehi _8212__32 (.L_HI(net32));
 sg13g2_tiehi _8211__33 (.L_HI(net33));
 sg13g2_tiehi _8210__34 (.L_HI(net34));
 sg13g2_tiehi _8209__35 (.L_HI(net35));
 sg13g2_tiehi _8208__36 (.L_HI(net36));
 sg13g2_tiehi _8207__37 (.L_HI(net37));
 sg13g2_tiehi _8206__38 (.L_HI(net38));
 sg13g2_tiehi _8205__39 (.L_HI(net39));
 sg13g2_tiehi _8204__40 (.L_HI(net40));
 sg13g2_tiehi _8203__41 (.L_HI(net41));
 sg13g2_tiehi _8202__42 (.L_HI(net42));
 sg13g2_tiehi _8201__43 (.L_HI(net43));
 sg13g2_tiehi _8200__44 (.L_HI(net44));
 sg13g2_tiehi _8199__45 (.L_HI(net45));
 sg13g2_tiehi _8198__46 (.L_HI(net46));
 sg13g2_tiehi _8197__47 (.L_HI(net47));
 sg13g2_tiehi _8196__48 (.L_HI(net48));
 sg13g2_tiehi _8195__49 (.L_HI(net49));
 sg13g2_tiehi _8194__50 (.L_HI(net50));
 sg13g2_tiehi _8193__51 (.L_HI(net51));
 sg13g2_tiehi _8192__52 (.L_HI(net52));
 sg13g2_tiehi _8191__53 (.L_HI(net53));
 sg13g2_tiehi _8190__54 (.L_HI(net54));
 sg13g2_tiehi _8189__55 (.L_HI(net55));
 sg13g2_tiehi _8188__56 (.L_HI(net56));
 sg13g2_tiehi _8187__57 (.L_HI(net57));
 sg13g2_tiehi _8186__58 (.L_HI(net58));
 sg13g2_tiehi _8185__59 (.L_HI(net59));
 sg13g2_tiehi _8184__60 (.L_HI(net60));
 sg13g2_tiehi _8183__61 (.L_HI(net61));
 sg13g2_tiehi _8182__62 (.L_HI(net62));
 sg13g2_tiehi _8181__63 (.L_HI(net63));
 sg13g2_tiehi _8180__64 (.L_HI(net64));
 sg13g2_tiehi _8179__65 (.L_HI(net65));
 sg13g2_tiehi _8178__66 (.L_HI(net66));
 sg13g2_tiehi _8177__67 (.L_HI(net67));
 sg13g2_tiehi _8176__68 (.L_HI(net68));
 sg13g2_tiehi _8175__69 (.L_HI(net69));
 sg13g2_tiehi _8174__70 (.L_HI(net70));
 sg13g2_tiehi _8173__71 (.L_HI(net71));
 sg13g2_tiehi _8172__72 (.L_HI(net72));
 sg13g2_tiehi _8171__73 (.L_HI(net73));
 sg13g2_tiehi _8170__74 (.L_HI(net74));
 sg13g2_tiehi _8169__75 (.L_HI(net75));
 sg13g2_tiehi _8168__76 (.L_HI(net76));
 sg13g2_tiehi _8167__77 (.L_HI(net77));
 sg13g2_tiehi _8166__78 (.L_HI(net78));
 sg13g2_tiehi _8165__79 (.L_HI(net79));
 sg13g2_tiehi _8164__80 (.L_HI(net80));
 sg13g2_tiehi _8163__81 (.L_HI(net81));
 sg13g2_tiehi _8162__82 (.L_HI(net82));
 sg13g2_tiehi _8161__83 (.L_HI(net83));
 sg13g2_tiehi _8160__84 (.L_HI(net84));
 sg13g2_tiehi _8159__85 (.L_HI(net85));
 sg13g2_tiehi _8158__86 (.L_HI(net86));
 sg13g2_tiehi _8157__87 (.L_HI(net87));
 sg13g2_tiehi _8156__88 (.L_HI(net88));
 sg13g2_tiehi _8155__89 (.L_HI(net89));
 sg13g2_tiehi _8154__90 (.L_HI(net90));
 sg13g2_tiehi _8153__91 (.L_HI(net91));
 sg13g2_tiehi _8152__92 (.L_HI(net92));
 sg13g2_tiehi _8151__93 (.L_HI(net93));
 sg13g2_tiehi _8150__94 (.L_HI(net94));
 sg13g2_tiehi _8149__95 (.L_HI(net95));
 sg13g2_tiehi _8148__96 (.L_HI(net96));
 sg13g2_tiehi _7975__97 (.L_HI(net97));
 sg13g2_tiehi _8147__98 (.L_HI(net98));
 sg13g2_tiehi _8146__99 (.L_HI(net99));
 sg13g2_tiehi _8145__100 (.L_HI(net100));
 sg13g2_tiehi _7981__101 (.L_HI(net101));
 sg13g2_tiehi _7982__102 (.L_HI(net102));
 sg13g2_tiehi _7983__103 (.L_HI(net103));
 sg13g2_tiehi _7984__104 (.L_HI(net104));
 sg13g2_tiehi _7985__105 (.L_HI(net105));
 sg13g2_tiehi _7986__106 (.L_HI(net106));
 sg13g2_tiehi _8144__107 (.L_HI(net107));
 sg13g2_tiehi _8143__108 (.L_HI(net108));
 sg13g2_tiehi _8142__109 (.L_HI(net109));
 sg13g2_tiehi _8141__110 (.L_HI(net110));
 sg13g2_tiehi _8140__111 (.L_HI(net111));
 sg13g2_tiehi _8139__112 (.L_HI(net112));
 sg13g2_tiehi _8138__113 (.L_HI(net113));
 sg13g2_tiehi _8137__114 (.L_HI(net114));
 sg13g2_tiehi _8136__115 (.L_HI(net115));
 sg13g2_tiehi _8135__116 (.L_HI(net116));
 sg13g2_tiehi _8134__117 (.L_HI(net117));
 sg13g2_tiehi _8133__118 (.L_HI(net118));
 sg13g2_tiehi _8132__119 (.L_HI(net119));
 sg13g2_tiehi _8131__120 (.L_HI(net120));
 sg13g2_tiehi _8130__121 (.L_HI(net121));
 sg13g2_tiehi _8129__122 (.L_HI(net122));
 sg13g2_tiehi _8128__123 (.L_HI(net123));
 sg13g2_tiehi _8127__124 (.L_HI(net124));
 sg13g2_tiehi _8126__125 (.L_HI(net125));
 sg13g2_tiehi _7987__126 (.L_HI(net126));
 sg13g2_tiehi _8125__127 (.L_HI(net127));
 sg13g2_tiehi _8124__128 (.L_HI(net128));
 sg13g2_tiehi _8123__129 (.L_HI(net129));
 sg13g2_tiehi _8122__130 (.L_HI(net130));
 sg13g2_tiehi _8121__131 (.L_HI(net131));
 sg13g2_tiehi _8120__132 (.L_HI(net132));
 sg13g2_tiehi _8119__133 (.L_HI(net133));
 sg13g2_tiehi _8031__134 (.L_HI(net134));
 sg13g2_tiehi _8118__135 (.L_HI(net135));
 sg13g2_tiehi _8117__136 (.L_HI(net136));
 sg13g2_tiehi _8116__137 (.L_HI(net137));
 sg13g2_tiehi _8115__138 (.L_HI(net138));
 sg13g2_tiehi _8114__139 (.L_HI(net139));
 sg13g2_tiehi _8113__140 (.L_HI(net140));
 sg13g2_tiehi _8112__141 (.L_HI(net141));
 sg13g2_tiehi _8111__142 (.L_HI(net142));
 sg13g2_tiehi _8110__143 (.L_HI(net143));
 sg13g2_tiehi _8109__144 (.L_HI(net144));
 sg13g2_tiehi _8108__145 (.L_HI(net145));
 sg13g2_tiehi _8107__146 (.L_HI(net146));
 sg13g2_tiehi _8106__147 (.L_HI(net147));
 sg13g2_tiehi _8105__148 (.L_HI(net148));
 sg13g2_tiehi _8104__149 (.L_HI(net149));
 sg13g2_tiehi _8103__150 (.L_HI(net150));
 sg13g2_tiehi _8102__151 (.L_HI(net151));
 sg13g2_tiehi _8101__152 (.L_HI(net152));
 sg13g2_tiehi _8091__153 (.L_HI(net153));
 sg13g2_tiehi _8090__154 (.L_HI(net154));
 sg13g2_tiehi _8093__155 (.L_HI(net155));
 sg13g2_tiehi _8094__156 (.L_HI(net156));
 sg13g2_tiehi _8095__157 (.L_HI(net157));
 sg13g2_tiehi _8096__158 (.L_HI(net158));
 sg13g2_tiehi _8097__159 (.L_HI(net159));
 sg13g2_tiehi _8098__160 (.L_HI(net160));
 sg13g2_tiehi _8099__161 (.L_HI(net161));
 sg13g2_tiehi _8089__162 (.L_HI(net162));
 sg13g2_tiehi _8088__163 (.L_HI(net163));
 sg13g2_tiehi _8087__164 (.L_HI(net164));
 sg13g2_tiehi _8086__165 (.L_HI(net165));
 sg13g2_tiehi _8085__166 (.L_HI(net166));
 sg13g2_tiehi _8633__167 (.L_HI(net167));
 sg13g2_tiehi _8649__168 (.L_HI(net168));
 sg13g2_tiehi _8632__169 (.L_HI(net169));
 sg13g2_tiehi _8637__170 (.L_HI(net170));
 sg13g2_tiehi _8631__171 (.L_HI(net171));
 sg13g2_tiehi _8057__172 (.L_HI(net172));
 sg13g2_tiehi _8630__173 (.L_HI(net173));
 sg13g2_tiehi _8025__174 (.L_HI(net174));
 sg13g2_tiehi _8523__175 (.L_HI(net175));
 sg13g2_tiehi _8522__176 (.L_HI(net176));
 sg13g2_tiehi _7991__177 (.L_HI(net177));
 sg13g2_tiehi _7989__178 (.L_HI(net178));
 sg13g2_tiehi _8521__179 (.L_HI(net179));
 sg13g2_tiehi _7988__180 (.L_HI(net180));
 sg13g2_tiehi _7979__181 (.L_HI(net181));
 sg13g2_tiehi _8520__182 (.L_HI(net182));
 sg13g2_tiehi _7968__183 (.L_HI(net183));
 sg13g2_tiehi _7966__184 (.L_HI(net184));
 sg13g2_tiehi _8519__185 (.L_HI(net185));
 sg13g2_tiehi _7952__186 (.L_HI(net186));
 sg13g2_tiehi _8518__187 (.L_HI(net187));
 sg13g2_tiehi _7950__188 (.L_HI(net188));
 sg13g2_tiehi _8517__189 (.L_HI(net189));
 sg13g2_tiehi _7948__190 (.L_HI(net190));
 sg13g2_tiehi _7946__191 (.L_HI(net191));
 sg13g2_tiehi _7942__192 (.L_HI(net192));
 sg13g2_tiehi _8516__193 (.L_HI(net193));
 sg13g2_tiehi _7939__194 (.L_HI(net194));
 sg13g2_tiehi _7938__195 (.L_HI(net195));
 sg13g2_tiehi _7937__196 (.L_HI(net196));
 sg13g2_tiehi _7936__197 (.L_HI(net197));
 sg13g2_tiehi _7935__198 (.L_HI(net198));
 sg13g2_tiehi _7934__199 (.L_HI(net199));
 sg13g2_tiehi _7933__200 (.L_HI(net200));
 sg13g2_tiehi _7932__201 (.L_HI(net201));
 sg13g2_tiehi _7931__202 (.L_HI(net202));
 sg13g2_tiehi _7929__203 (.L_HI(net203));
 sg13g2_tiehi _7928__204 (.L_HI(net204));
 sg13g2_tiehi _8515__205 (.L_HI(net205));
 sg13g2_tiehi _7927__206 (.L_HI(net206));
 sg13g2_tiehi _7902__207 (.L_HI(net207));
 sg13g2_tiehi _7901__208 (.L_HI(net208));
 sg13g2_tiehi _7900__209 (.L_HI(net209));
 sg13g2_tiehi _7899__210 (.L_HI(net210));
 sg13g2_tiehi _8100__211 (.L_HI(net211));
 sg13g2_tiehi _7898__212 (.L_HI(net212));
 sg13g2_tiehi _7897__213 (.L_HI(net213));
 sg13g2_tiehi _8219__214 (.L_HI(net214));
 sg13g2_tiehi _7896__215 (.L_HI(net215));
 sg13g2_tiehi _7895__216 (.L_HI(net216));
 sg13g2_tiehi _7894__217 (.L_HI(net217));
 sg13g2_tiehi _7893__218 (.L_HI(net218));
 sg13g2_tiehi _7892__219 (.L_HI(net219));
 sg13g2_tiehi _7891__220 (.L_HI(net220));
 sg13g2_tiehi _7890__221 (.L_HI(net221));
 sg13g2_tiehi _7889__222 (.L_HI(net222));
 sg13g2_tiehi _8514__223 (.L_HI(net223));
 sg13g2_tiehi _8248__224 (.L_HI(net224));
 sg13g2_tiehi _8513__225 (.L_HI(net225));
 sg13g2_tiehi _8512__226 (.L_HI(net226));
 sg13g2_tiehi _8511__227 (.L_HI(net227));
 sg13g2_tiehi _8510__228 (.L_HI(net228));
 sg13g2_tiehi _8509__229 (.L_HI(net229));
 sg13g2_tiehi _8508__230 (.L_HI(net230));
 sg13g2_tiehi _8507__231 (.L_HI(net231));
 sg13g2_tiehi _8506__232 (.L_HI(net232));
 sg13g2_tiehi _8505__233 (.L_HI(net233));
 sg13g2_tiehi _8504__234 (.L_HI(net234));
 sg13g2_tiehi _8503__235 (.L_HI(net235));
 sg13g2_tiehi _8502__236 (.L_HI(net236));
 sg13g2_tiehi _8501__237 (.L_HI(net237));
 sg13g2_tiehi _8500__238 (.L_HI(net238));
 sg13g2_tiehi _8499__239 (.L_HI(net239));
 sg13g2_tiehi _8498__240 (.L_HI(net240));
 sg13g2_tiehi _8497__241 (.L_HI(net241));
 sg13g2_tiehi _8496__242 (.L_HI(net242));
 sg13g2_tiehi _8495__243 (.L_HI(net243));
 sg13g2_tiehi _8494__244 (.L_HI(net244));
 sg13g2_tiehi _8493__245 (.L_HI(net245));
 sg13g2_tiehi _8492__246 (.L_HI(net246));
 sg13g2_tiehi _8491__247 (.L_HI(net247));
 sg13g2_tiehi _8490__248 (.L_HI(net248));
 sg13g2_tiehi _8489__249 (.L_HI(net249));
 sg13g2_tiehi _8488__250 (.L_HI(net250));
 sg13g2_tiehi _8487__251 (.L_HI(net251));
 sg13g2_tiehi _8486__252 (.L_HI(net252));
 sg13g2_tiehi _8485__253 (.L_HI(net253));
 sg13g2_tiehi _8484__254 (.L_HI(net254));
 sg13g2_tiehi _8483__255 (.L_HI(net255));
 sg13g2_tiehi _8482__256 (.L_HI(net256));
 sg13g2_tiehi _8481__257 (.L_HI(net257));
 sg13g2_tiehi _8480__258 (.L_HI(net258));
 sg13g2_tiehi _8479__259 (.L_HI(net259));
 sg13g2_tiehi _8478__260 (.L_HI(net260));
 sg13g2_tiehi _8477__261 (.L_HI(net261));
 sg13g2_tiehi _8476__262 (.L_HI(net262));
 sg13g2_tiehi _8475__263 (.L_HI(net263));
 sg13g2_tiehi _8474__264 (.L_HI(net264));
 sg13g2_tiehi _8473__265 (.L_HI(net265));
 sg13g2_tiehi _8472__266 (.L_HI(net266));
 sg13g2_tiehi _8471__267 (.L_HI(net267));
 sg13g2_tiehi _8470__268 (.L_HI(net268));
 sg13g2_tiehi _8469__269 (.L_HI(net269));
 sg13g2_tiehi _8468__270 (.L_HI(net270));
 sg13g2_tiehi _8467__271 (.L_HI(net271));
 sg13g2_tiehi _8466__272 (.L_HI(net272));
 sg13g2_tiehi _8465__273 (.L_HI(net273));
 sg13g2_tiehi _8464__274 (.L_HI(net274));
 sg13g2_tiehi _8463__275 (.L_HI(net275));
 sg13g2_tiehi _8462__276 (.L_HI(net276));
 sg13g2_tiehi _8461__277 (.L_HI(net277));
 sg13g2_tiehi _8448__278 (.L_HI(net278));
 sg13g2_tiehi _8447__279 (.L_HI(net279));
 sg13g2_tiehi _8446__280 (.L_HI(net280));
 sg13g2_tiehi _8445__281 (.L_HI(net281));
 sg13g2_tiehi _8444__282 (.L_HI(net282));
 sg13g2_tiehi _8443__283 (.L_HI(net283));
 sg13g2_tiehi _8442__284 (.L_HI(net284));
 sg13g2_tiehi _8441__285 (.L_HI(net285));
 sg13g2_tiehi _8636__286 (.L_HI(net286));
 sg13g2_tiehi _8432__287 (.L_HI(net287));
 sg13g2_tiehi _8431__288 (.L_HI(net288));
 sg13g2_tiehi _8430__289 (.L_HI(net289));
 sg13g2_tiehi _8429__290 (.L_HI(net290));
 sg13g2_tiehi _8428__291 (.L_HI(net291));
 sg13g2_tiehi _8427__292 (.L_HI(net292));
 sg13g2_tiehi _8426__293 (.L_HI(net293));
 sg13g2_tiehi _8425__294 (.L_HI(net294));
 sg13g2_tiehi _8424__295 (.L_HI(net295));
 sg13g2_tiehi _8423__296 (.L_HI(net296));
 sg13g2_tiehi _8422__297 (.L_HI(net297));
 sg13g2_tiehi _8421__298 (.L_HI(net298));
 sg13g2_tiehi _8420__299 (.L_HI(net299));
 sg13g2_tiehi _8419__300 (.L_HI(net300));
 sg13g2_tiehi _8418__301 (.L_HI(net301));
 sg13g2_tiehi _8417__302 (.L_HI(net302));
 sg13g2_tiehi _8406__303 (.L_HI(net303));
 sg13g2_tiehi _8635__304 (.L_HI(net304));
 sg13g2_tiehi _8400__305 (.L_HI(net305));
 sg13g2_tiehi _8399__306 (.L_HI(net306));
 sg13g2_tiehi _8398__307 (.L_HI(net307));
 sg13g2_tiehi _8397__308 (.L_HI(net308));
 sg13g2_tiehi _8396__309 (.L_HI(net309));
 sg13g2_tiehi _8395__310 (.L_HI(net310));
 sg13g2_tiehi _8394__311 (.L_HI(net311));
 sg13g2_tiehi _8386__312 (.L_HI(net312));
 sg13g2_tiehi _8385__313 (.L_HI(net313));
 sg13g2_tiehi _8382__314 (.L_HI(net314));
 sg13g2_tiehi _8381__315 (.L_HI(net315));
 sg13g2_tiehi _8380__316 (.L_HI(net316));
 sg13g2_tiehi _8379__317 (.L_HI(net317));
 sg13g2_tiehi _8378__318 (.L_HI(net318));
 sg13g2_tiehi _8377__319 (.L_HI(net319));
 sg13g2_tiehi _8376__320 (.L_HI(net320));
 sg13g2_tiehi _8375__321 (.L_HI(net321));
 sg13g2_tiehi _8374__322 (.L_HI(net322));
 sg13g2_tiehi _8373__323 (.L_HI(net323));
 sg13g2_tiehi _8372__324 (.L_HI(net324));
 sg13g2_tiehi _8371__325 (.L_HI(net325));
 sg13g2_tiehi _8339__326 (.L_HI(net326));
 sg13g2_tiehi _8370__327 (.L_HI(net327));
 sg13g2_tiehi _8369__328 (.L_HI(net328));
 sg13g2_tiehi _8368__329 (.L_HI(net329));
 sg13g2_tiehi _8367__330 (.L_HI(net330));
 sg13g2_tiehi _8366__331 (.L_HI(net331));
 sg13g2_tiehi _8365__332 (.L_HI(net332));
 sg13g2_tiehi _8364__333 (.L_HI(net333));
 sg13g2_tiehi _8363__334 (.L_HI(net334));
 sg13g2_tiehi _8362__335 (.L_HI(net335));
 sg13g2_tiehi _8361__336 (.L_HI(net336));
 sg13g2_tiehi _8360__337 (.L_HI(net337));
 sg13g2_tiehi _8359__338 (.L_HI(net338));
 sg13g2_tiehi _8358__339 (.L_HI(net339));
 sg13g2_tiehi _8401__340 (.L_HI(net340));
 sg13g2_tiehi _8357__341 (.L_HI(net341));
 sg13g2_tiehi _8356__342 (.L_HI(net342));
 sg13g2_tiehi _8404__343 (.L_HI(net343));
 sg13g2_tiehi _8407__344 (.L_HI(net344));
 sg13g2_tiehi _8355__345 (.L_HI(net345));
 sg13g2_tiehi _8354__346 (.L_HI(net346));
 sg13g2_tiehi _8353__347 (.L_HI(net347));
 sg13g2_tiehi _8352__348 (.L_HI(net348));
 sg13g2_tiehi _8351__349 (.L_HI(net349));
 sg13g2_tiehi _8350__350 (.L_HI(net350));
 sg13g2_tiehi _8349__351 (.L_HI(net351));
 sg13g2_tiehi _8348__352 (.L_HI(net352));
 sg13g2_tiehi _8347__353 (.L_HI(net353));
 sg13g2_tiehi _8346__354 (.L_HI(net354));
 sg13g2_tiehi _8345__355 (.L_HI(net355));
 sg13g2_tiehi _8344__356 (.L_HI(net356));
 sg13g2_tiehi _8343__357 (.L_HI(net357));
 sg13g2_tiehi _8342__358 (.L_HI(net358));
 sg13g2_tiehi _8341__359 (.L_HI(net359));
 sg13g2_tiehi _8338__360 (.L_HI(net360));
 sg13g2_tiehi _8337__361 (.L_HI(net361));
 sg13g2_tiehi _8336__362 (.L_HI(net362));
 sg13g2_tiehi _8335__363 (.L_HI(net363));
 sg13g2_tiehi _8334__364 (.L_HI(net364));
 sg13g2_tiehi _8333__365 (.L_HI(net365));
 sg13g2_tiehi _8332__366 (.L_HI(net366));
 sg13g2_tiehi _8331__367 (.L_HI(net367));
 sg13g2_tiehi _8330__368 (.L_HI(net368));
 sg13g2_tiehi _8329__369 (.L_HI(net369));
 sg13g2_tiehi _8328__370 (.L_HI(net370));
 sg13g2_tiehi _8327__371 (.L_HI(net371));
 sg13g2_tiehi _8326__372 (.L_HI(net372));
 sg13g2_tiehi _8325__373 (.L_HI(net373));
 sg13g2_tiehi _8324__374 (.L_HI(net374));
 sg13g2_tiehi _8323__375 (.L_HI(net375));
 sg13g2_tiehi _8322__376 (.L_HI(net376));
 sg13g2_tiehi _8415__377 (.L_HI(net377));
 sg13g2_tiehi _8449__378 (.L_HI(net378));
 sg13g2_tiehi _8321__379 (.L_HI(net379));
 sg13g2_tiehi _8320__380 (.L_HI(net380));
 sg13g2_tiehi _8319__381 (.L_HI(net381));
 sg13g2_tiehi _8318__382 (.L_HI(net382));
 sg13g2_tiehi _8317__383 (.L_HI(net383));
 sg13g2_tiehi _8316__384 (.L_HI(net384));
 sg13g2_tiehi _8315__385 (.L_HI(net385));
 sg13g2_tiehi _8314__386 (.L_HI(net386));
 sg13g2_tiehi _8313__387 (.L_HI(net387));
 sg13g2_tiehi _8312__388 (.L_HI(net388));
 sg13g2_tiehi _8311__389 (.L_HI(net389));
 sg13g2_tiehi _8310__390 (.L_HI(net390));
 sg13g2_tiehi _8309__391 (.L_HI(net391));
 sg13g2_tiehi _8308__392 (.L_HI(net392));
 sg13g2_tiehi _8307__393 (.L_HI(net393));
 sg13g2_tiehi _8306__394 (.L_HI(net394));
 sg13g2_tiehi _8305__395 (.L_HI(net395));
 sg13g2_tiehi _8304__396 (.L_HI(net396));
 sg13g2_tiehi _8303__397 (.L_HI(net397));
 sg13g2_tiehi _8302__398 (.L_HI(net398));
 sg13g2_tiehi _8301__399 (.L_HI(net399));
 sg13g2_tiehi _8300__400 (.L_HI(net400));
 sg13g2_tiehi _8299__401 (.L_HI(net401));
 sg13g2_tiehi _8298__402 (.L_HI(net402));
 sg13g2_tiehi _8297__403 (.L_HI(net403));
 sg13g2_tiehi _8296__404 (.L_HI(net404));
 sg13g2_tiehi _8295__405 (.L_HI(net405));
 sg13g2_tiehi _8294__406 (.L_HI(net406));
 sg13g2_tiehi _8293__407 (.L_HI(net407));
 sg13g2_tiehi _8292__408 (.L_HI(net408));
 sg13g2_tiehi _8291__409 (.L_HI(net409));
 sg13g2_tiehi _8290__410 (.L_HI(net410));
 sg13g2_tiehi _8289__411 (.L_HI(net411));
 sg13g2_tiehi _8288__412 (.L_HI(net412));
 sg13g2_tiehi _8287__413 (.L_HI(net413));
 sg13g2_tiehi _8286__414 (.L_HI(net414));
 sg13g2_tiehi _8285__415 (.L_HI(net415));
 sg13g2_tiehi _8284__416 (.L_HI(net416));
 sg13g2_tiehi _8283__417 (.L_HI(net417));
 sg13g2_tiehi _8282__418 (.L_HI(net418));
 sg13g2_tiehi _8281__419 (.L_HI(net419));
 sg13g2_tiehi _8280__420 (.L_HI(net420));
 sg13g2_tiehi _8279__421 (.L_HI(net421));
 sg13g2_tiehi _8278__422 (.L_HI(net422));
 sg13g2_tiehi _8277__423 (.L_HI(net423));
 sg13g2_tiehi _8276__424 (.L_HI(net424));
 sg13g2_tiehi _8275__425 (.L_HI(net425));
 sg13g2_tiehi _8274__426 (.L_HI(net426));
 sg13g2_tiehi _8273__427 (.L_HI(net427));
 sg13g2_tiehi _8272__428 (.L_HI(net428));
 sg13g2_tiehi _8271__429 (.L_HI(net429));
 sg13g2_tiehi _8270__430 (.L_HI(net430));
 sg13g2_tiehi _8269__431 (.L_HI(net431));
 sg13g2_tiehi _8268__432 (.L_HI(net432));
 sg13g2_tiehi _8267__433 (.L_HI(net433));
 sg13g2_tiehi _8266__434 (.L_HI(net434));
 sg13g2_tiehi _8265__435 (.L_HI(net435));
 sg13g2_tiehi _8264__436 (.L_HI(net436));
 sg13g2_tiehi _8263__437 (.L_HI(net437));
 sg13g2_tiehi _8262__438 (.L_HI(net438));
 sg13g2_tiehi _8261__439 (.L_HI(net439));
 sg13g2_tiehi _8260__440 (.L_HI(net440));
 sg13g2_tiehi _8259__441 (.L_HI(net441));
 sg13g2_tiehi _8258__442 (.L_HI(net442));
 sg13g2_tiehi _8257__443 (.L_HI(net443));
 sg13g2_tiehi _8256__444 (.L_HI(net444));
 sg13g2_tiehi _8524__445 (.L_HI(net445));
 sg13g2_tiehi _8525__446 (.L_HI(net446));
 sg13g2_tiehi _8526__447 (.L_HI(net447));
 sg13g2_tiehi _8527__448 (.L_HI(net448));
 sg13g2_tiehi _8528__449 (.L_HI(net449));
 sg13g2_tiehi _8529__450 (.L_HI(net450));
 sg13g2_tiehi _8530__451 (.L_HI(net451));
 sg13g2_tiehi _8531__452 (.L_HI(net452));
 sg13g2_tiehi _8532__453 (.L_HI(net453));
 sg13g2_tiehi _8533__454 (.L_HI(net454));
 sg13g2_tiehi _8534__455 (.L_HI(net455));
 sg13g2_tiehi _8535__456 (.L_HI(net456));
 sg13g2_tiehi _8536__457 (.L_HI(net457));
 sg13g2_tiehi _8537__458 (.L_HI(net458));
 sg13g2_tiehi _8538__459 (.L_HI(net459));
 sg13g2_tiehi _8539__460 (.L_HI(net460));
 sg13g2_tiehi _8540__461 (.L_HI(net461));
 sg13g2_tiehi _8541__462 (.L_HI(net462));
 sg13g2_tiehi _8542__463 (.L_HI(net463));
 sg13g2_tiehi _8543__464 (.L_HI(net464));
 sg13g2_tiehi _8544__465 (.L_HI(net465));
 sg13g2_tiehi _8545__466 (.L_HI(net466));
 sg13g2_tiehi _8553__467 (.L_HI(net467));
 sg13g2_tiehi _8554__468 (.L_HI(net468));
 sg13g2_tiehi _8555__469 (.L_HI(net469));
 sg13g2_tiehi _8556__470 (.L_HI(net470));
 sg13g2_tiehi _8557__471 (.L_HI(net471));
 sg13g2_tiehi _8558__472 (.L_HI(net472));
 sg13g2_tiehi _8559__473 (.L_HI(net473));
 sg13g2_tiehi _8560__474 (.L_HI(net474));
 sg13g2_tiehi _8255__475 (.L_HI(net475));
 sg13g2_tiehi _8583__476 (.L_HI(net476));
 sg13g2_tiehi _8584__477 (.L_HI(net477));
 sg13g2_tiehi _8585__478 (.L_HI(net478));
 sg13g2_tiehi _8586__479 (.L_HI(net479));
 sg13g2_tiehi _8587__480 (.L_HI(net480));
 sg13g2_tiehi _8588__481 (.L_HI(net481));
 sg13g2_tiehi _8589__482 (.L_HI(net482));
 sg13g2_tiehi _8590__483 (.L_HI(net483));
 sg13g2_tiehi _8591__484 (.L_HI(net484));
 sg13g2_tiehi _8592__485 (.L_HI(net485));
 sg13g2_tiehi _8593__486 (.L_HI(net486));
 sg13g2_tiehi _8594__487 (.L_HI(net487));
 sg13g2_tiehi _8595__488 (.L_HI(net488));
 sg13g2_tiehi _8596__489 (.L_HI(net489));
 sg13g2_tiehi _8597__490 (.L_HI(net490));
 sg13g2_tiehi _8598__491 (.L_HI(net491));
 sg13g2_tiehi _8599__492 (.L_HI(net492));
 sg13g2_tiehi _8600__493 (.L_HI(net493));
 sg13g2_tiehi _8601__494 (.L_HI(net494));
 sg13g2_tiehi _8602__495 (.L_HI(net495));
 sg13g2_tiehi _8603__496 (.L_HI(net496));
 sg13g2_tiehi _8604__497 (.L_HI(net497));
 sg13g2_tiehi _8605__498 (.L_HI(net498));
 sg13g2_tiehi _8606__499 (.L_HI(net499));
 sg13g2_tiehi _8607__500 (.L_HI(net500));
 sg13g2_tiehi _8608__501 (.L_HI(net501));
 sg13g2_tiehi _8609__502 (.L_HI(net502));
 sg13g2_tiehi _8610__503 (.L_HI(net503));
 sg13g2_tiehi _8611__504 (.L_HI(net504));
 sg13g2_tiehi _8612__505 (.L_HI(net505));
 sg13g2_tiehi _8613__506 (.L_HI(net506));
 sg13g2_tiehi _8614__507 (.L_HI(net507));
 sg13g2_tiehi _8615__508 (.L_HI(net508));
 sg13g2_tiehi _8616__509 (.L_HI(net509));
 sg13g2_tiehi _8617__510 (.L_HI(net510));
 sg13g2_tiehi _8618__511 (.L_HI(net511));
 sg13g2_tiehi _8619__512 (.L_HI(net512));
 sg13g2_tiehi _8620__513 (.L_HI(net513));
 sg13g2_tiehi _8621__514 (.L_HI(net514));
 sg13g2_tiehi _8622__515 (.L_HI(net515));
 sg13g2_tiehi _8623__516 (.L_HI(net516));
 sg13g2_tiehi _8624__517 (.L_HI(net517));
 sg13g2_tiehi _8625__518 (.L_HI(net518));
 sg13g2_tiehi _8626__519 (.L_HI(net519));
 sg13g2_tiehi _8627__520 (.L_HI(net520));
 sg13g2_tiehi _8628__521 (.L_HI(net521));
 sg13g2_tiehi _8254__522 (.L_HI(net522));
 sg13g2_tiehi _8253__523 (.L_HI(net523));
 sg13g2_tiehi _8252__524 (.L_HI(net524));
 sg13g2_tiehi _8247__525 (.L_HI(net525));
 sg13g2_tiehi _8634__526 (.L_HI(net526));
 sg13g2_tiehi _8629__527 (.L_HI(net527));
 sg13g2_inv_1 _4530__1 (.Y(net528),
    .A(clknet_1_1__leaf_clk));
 sg13g2_buf_2 _9161_ (.A(\usbfunction0.scl_usbgpiophy0.n6496_o ),
    .X(uio_oe[6]));
 sg13g2_buf_2 _9162_ (.A(\usbfunction0.scl_usbgpiophy0.n6496_o ),
    .X(uio_oe[7]));
 sg13g2_buf_1 _9163_ (.A(n106_o),
    .X(uio_out[0]));
 sg13g2_buf_1 _9164_ (.A(n118_o),
    .X(uio_out[2]));
 sg13g2_buf_1 _9165_ (.A(n124_o),
    .X(uio_out[3]));
 sg13g2_buf_1 _9166_ (.A(n130_o),
    .X(uio_out[4]));
 sg13g2_buf_1 _9167_ (.A(n136_o),
    .X(uio_out[5]));
 sg13g2_buf_2 _9168_ (.A(\usbfunction0.scl_usbgpiophy0.n6500_o ),
    .X(uio_out[6]));
 sg13g2_buf_2 _9169_ (.A(\usbfunction0.scl_usbgpiophy0.n6503_o ),
    .X(uio_out[7]));
 sg13g2_buf_1 _9170_ (.A(s_m_io10_out),
    .X(uo_out[2]));
 sg13g2_buf_1 _9171_ (.A(s_m_io11_out),
    .X(uo_out[3]));
 sg13g2_buf_1 _9172_ (.A(s_m_io12_out),
    .X(uo_out[4]));
 sg13g2_buf_1 _9173_ (.A(s_m_io13_out),
    .X(uo_out[5]));
 sg13g2_buf_1 _9174_ (.A(s_m_io14_out),
    .X(uo_out[6]));
 sg13g2_buf_1 _9175_ (.A(s_m_io15_out),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout1173 (.A(net1174),
    .X(net1173));
 sg13g2_buf_1 fanout1174 (.A(net1175),
    .X(net1174));
 sg13g2_buf_2 fanout1175 (.A(\scl_fifo0.n2697_o[3] ),
    .X(net1175));
 sg13g2_buf_2 fanout1176 (.A(net1178),
    .X(net1176));
 sg13g2_buf_2 fanout1177 (.A(net1178),
    .X(net1177));
 sg13g2_buf_2 fanout1178 (.A(net1179),
    .X(net1178));
 sg13g2_buf_4 fanout1179 (.X(net1179),
    .A(_1652_));
 sg13g2_buf_4 fanout1180 (.X(net1180),
    .A(net1182));
 sg13g2_buf_2 fanout1181 (.A(net1182),
    .X(net1181));
 sg13g2_buf_2 fanout1182 (.A(\scl_fifo0.n2697_o[2] ),
    .X(net1182));
 sg13g2_buf_2 fanout1183 (.A(_3068_),
    .X(net1183));
 sg13g2_buf_2 fanout1184 (.A(_3068_),
    .X(net1184));
 sg13g2_buf_2 fanout1185 (.A(_3002_),
    .X(net1185));
 sg13g2_buf_2 fanout1186 (.A(_3002_),
    .X(net1186));
 sg13g2_buf_2 fanout1187 (.A(_2724_),
    .X(net1187));
 sg13g2_buf_2 fanout1188 (.A(_2724_),
    .X(net1188));
 sg13g2_buf_2 fanout1189 (.A(net1190),
    .X(net1189));
 sg13g2_buf_4 fanout1190 (.X(net1190),
    .A(_1347_));
 sg13g2_buf_2 fanout1191 (.A(net1195),
    .X(net1191));
 sg13g2_buf_2 fanout1192 (.A(net1195),
    .X(net1192));
 sg13g2_buf_2 fanout1193 (.A(net1194),
    .X(net1193));
 sg13g2_buf_2 fanout1194 (.A(net1195),
    .X(net1194));
 sg13g2_buf_2 fanout1195 (.A(\scl_fifo0.n2697_o[1] ),
    .X(net1195));
 sg13g2_buf_2 fanout1196 (.A(_3092_),
    .X(net1196));
 sg13g2_buf_2 fanout1197 (.A(_3092_),
    .X(net1197));
 sg13g2_buf_2 fanout1198 (.A(_3084_),
    .X(net1198));
 sg13g2_buf_2 fanout1199 (.A(_3084_),
    .X(net1199));
 sg13g2_buf_2 fanout1200 (.A(_3076_),
    .X(net1200));
 sg13g2_buf_2 fanout1201 (.A(_3076_),
    .X(net1201));
 sg13g2_buf_2 fanout1202 (.A(_3060_),
    .X(net1202));
 sg13g2_buf_2 fanout1203 (.A(_3060_),
    .X(net1203));
 sg13g2_buf_2 fanout1204 (.A(_3052_),
    .X(net1204));
 sg13g2_buf_2 fanout1205 (.A(_3052_),
    .X(net1205));
 sg13g2_buf_2 fanout1206 (.A(net1207),
    .X(net1206));
 sg13g2_buf_2 fanout1207 (.A(_3044_),
    .X(net1207));
 sg13g2_buf_2 fanout1208 (.A(_3035_),
    .X(net1208));
 sg13g2_buf_2 fanout1209 (.A(_3035_),
    .X(net1209));
 sg13g2_buf_2 fanout1210 (.A(_3027_),
    .X(net1210));
 sg13g2_buf_2 fanout1211 (.A(_3027_),
    .X(net1211));
 sg13g2_buf_2 fanout1212 (.A(net1214),
    .X(net1212));
 sg13g2_buf_1 fanout1213 (.A(net1214),
    .X(net1213));
 sg13g2_buf_2 fanout1214 (.A(_3019_),
    .X(net1214));
 sg13g2_buf_2 fanout1215 (.A(net1216),
    .X(net1215));
 sg13g2_buf_4 fanout1216 (.X(net1216),
    .A(_3011_));
 sg13g2_buf_2 fanout1217 (.A(net1218),
    .X(net1217));
 sg13g2_buf_2 fanout1218 (.A(_2994_),
    .X(net1218));
 sg13g2_buf_2 fanout1219 (.A(_2985_),
    .X(net1219));
 sg13g2_buf_2 fanout1220 (.A(_2985_),
    .X(net1220));
 sg13g2_buf_2 fanout1221 (.A(_2767_),
    .X(net1221));
 sg13g2_buf_2 fanout1222 (.A(_2767_),
    .X(net1222));
 sg13g2_buf_2 fanout1223 (.A(_1995_),
    .X(net1223));
 sg13g2_buf_4 fanout1224 (.X(net1224),
    .A(_1995_));
 sg13g2_buf_4 fanout1225 (.X(net1225),
    .A(net1226));
 sg13g2_buf_4 fanout1226 (.X(net1226),
    .A(net1229));
 sg13g2_buf_4 fanout1227 (.X(net1227),
    .A(net1228));
 sg13g2_buf_4 fanout1228 (.X(net1228),
    .A(net1229));
 sg13g2_buf_2 fanout1229 (.A(net1234),
    .X(net1229));
 sg13g2_buf_4 fanout1230 (.X(net1230),
    .A(net1232));
 sg13g2_buf_4 fanout1231 (.X(net1231),
    .A(net1232));
 sg13g2_buf_4 fanout1232 (.X(net1232),
    .A(net1234));
 sg13g2_buf_4 fanout1233 (.X(net1233),
    .A(net1234));
 sg13g2_buf_2 fanout1234 (.A(_1342_),
    .X(net1234));
 sg13g2_buf_2 fanout1235 (.A(net1236),
    .X(net1235));
 sg13g2_buf_1 fanout1236 (.A(net1237),
    .X(net1236));
 sg13g2_buf_4 fanout1237 (.X(net1237),
    .A(_1341_));
 sg13g2_buf_2 fanout1238 (.A(net1240),
    .X(net1238));
 sg13g2_buf_1 fanout1239 (.A(net1240),
    .X(net1239));
 sg13g2_buf_2 fanout1240 (.A(_1341_),
    .X(net1240));
 sg13g2_buf_4 fanout1241 (.X(net1241),
    .A(_0919_));
 sg13g2_buf_4 fanout1242 (.X(net1242),
    .A(net1243));
 sg13g2_buf_2 fanout1243 (.A(_2772_),
    .X(net1243));
 sg13g2_buf_2 fanout1244 (.A(_2761_),
    .X(net1244));
 sg13g2_buf_2 fanout1245 (.A(_2761_),
    .X(net1245));
 sg13g2_buf_4 fanout1246 (.X(net1246),
    .A(net1248));
 sg13g2_buf_2 fanout1247 (.A(net1248),
    .X(net1247));
 sg13g2_buf_2 fanout1248 (.A(_2755_),
    .X(net1248));
 sg13g2_buf_4 fanout1249 (.X(net1249),
    .A(_2749_));
 sg13g2_buf_4 fanout1250 (.X(net1250),
    .A(_2749_));
 sg13g2_buf_4 fanout1251 (.X(net1251),
    .A(_2743_));
 sg13g2_buf_4 fanout1252 (.X(net1252),
    .A(_2743_));
 sg13g2_buf_4 fanout1253 (.X(net1253),
    .A(_2735_));
 sg13g2_buf_2 fanout1254 (.A(_2735_),
    .X(net1254));
 sg13g2_buf_4 fanout1255 (.X(net1255),
    .A(net1256));
 sg13g2_buf_4 fanout1256 (.X(net1256),
    .A(_2729_));
 sg13g2_buf_2 fanout1257 (.A(_1989_),
    .X(net1257));
 sg13g2_buf_2 fanout1258 (.A(_1989_),
    .X(net1258));
 sg13g2_buf_2 fanout1259 (.A(net1260),
    .X(net1259));
 sg13g2_buf_2 fanout1260 (.A(_0920_),
    .X(net1260));
 sg13g2_buf_4 fanout1261 (.X(net1261),
    .A(_1317_));
 sg13g2_buf_2 fanout1262 (.A(_1317_),
    .X(net1262));
 sg13g2_buf_2 fanout1263 (.A(net1264),
    .X(net1263));
 sg13g2_buf_2 fanout1264 (.A(_1718_),
    .X(net1264));
 sg13g2_buf_2 fanout1265 (.A(_1215_),
    .X(net1265));
 sg13g2_buf_4 fanout1266 (.X(net1266),
    .A(\scl_fifo1.n6238_o[3] ));
 sg13g2_buf_2 fanout1267 (.A(_1711_),
    .X(net1267));
 sg13g2_buf_4 fanout1268 (.X(net1268),
    .A(_1702_));
 sg13g2_buf_2 fanout1269 (.A(_1214_),
    .X(net1269));
 sg13g2_buf_2 fanout1270 (.A(net1271),
    .X(net1270));
 sg13g2_buf_2 fanout1271 (.A(_1213_),
    .X(net1271));
 sg13g2_buf_2 fanout1272 (.A(net1273),
    .X(net1272));
 sg13g2_buf_4 fanout1273 (.X(net1273),
    .A(\scl_fifo1.n6238_o[2] ));
 sg13g2_buf_2 fanout1274 (.A(_1055_),
    .X(net1274));
 sg13g2_buf_2 fanout1275 (.A(net1276),
    .X(net1275));
 sg13g2_buf_2 fanout1276 (.A(net1277),
    .X(net1276));
 sg13g2_buf_2 fanout1277 (.A(_1695_),
    .X(net1277));
 sg13g2_buf_2 fanout1278 (.A(net1279),
    .X(net1278));
 sg13g2_buf_2 fanout1279 (.A(_1694_),
    .X(net1279));
 sg13g2_buf_2 fanout1280 (.A(_1064_),
    .X(net1280));
 sg13g2_buf_2 fanout1281 (.A(_1064_),
    .X(net1281));
 sg13g2_buf_2 fanout1282 (.A(net1283),
    .X(net1282));
 sg13g2_buf_4 fanout1283 (.X(net1283),
    .A(net1287));
 sg13g2_buf_2 fanout1284 (.A(net1286),
    .X(net1284));
 sg13g2_buf_1 fanout1285 (.A(net1286),
    .X(net1285));
 sg13g2_buf_2 fanout1286 (.A(net1287),
    .X(net1286));
 sg13g2_buf_2 fanout1287 (.A(net1293),
    .X(net1287));
 sg13g2_buf_4 fanout1288 (.X(net1288),
    .A(net1293));
 sg13g2_buf_1 fanout1289 (.A(net1293),
    .X(net1289));
 sg13g2_buf_2 fanout1290 (.A(net1292),
    .X(net1290));
 sg13g2_buf_2 fanout1291 (.A(net1292),
    .X(net1291));
 sg13g2_buf_2 fanout1292 (.A(net1293),
    .X(net1292));
 sg13g2_buf_2 fanout1293 (.A(\scl_fifo1.n6238_o[0] ),
    .X(net1293));
 sg13g2_buf_2 fanout1294 (.A(net1295),
    .X(net1294));
 sg13g2_buf_2 fanout1295 (.A(\scl_fifo1.n6238_o[1] ),
    .X(net1295));
 sg13g2_buf_2 fanout1296 (.A(net1299),
    .X(net1296));
 sg13g2_buf_1 fanout1297 (.A(net1299),
    .X(net1297));
 sg13g2_buf_2 fanout1298 (.A(net1299),
    .X(net1298));
 sg13g2_buf_2 fanout1299 (.A(\scl_fifo1.n6238_o[1] ),
    .X(net1299));
 sg13g2_buf_2 fanout1300 (.A(net1304),
    .X(net1300));
 sg13g2_buf_2 fanout1301 (.A(net1304),
    .X(net1301));
 sg13g2_buf_2 fanout1302 (.A(net1304),
    .X(net1302));
 sg13g2_buf_2 fanout1303 (.A(net1304),
    .X(net1303));
 sg13g2_buf_2 fanout1304 (.A(\scl_fifo1.n6238_o[1] ),
    .X(net1304));
 sg13g2_buf_4 fanout1305 (.X(net1305),
    .A(net1307));
 sg13g2_buf_1 fanout1306 (.A(net1307),
    .X(net1306));
 sg13g2_buf_1 fanout1307 (.A(_1686_),
    .X(net1307));
 sg13g2_buf_4 fanout1308 (.X(net1308),
    .A(net1310));
 sg13g2_buf_1 fanout1309 (.A(net1310),
    .X(net1309));
 sg13g2_buf_2 fanout1310 (.A(_1685_),
    .X(net1310));
 sg13g2_buf_2 fanout1311 (.A(net1312),
    .X(net1311));
 sg13g2_buf_4 fanout1312 (.X(net1312),
    .A(net1313));
 sg13g2_buf_2 fanout1313 (.A(_1678_),
    .X(net1313));
 sg13g2_buf_2 fanout1314 (.A(_1677_),
    .X(net1314));
 sg13g2_buf_2 fanout1315 (.A(_1677_),
    .X(net1315));
 sg13g2_buf_4 fanout1316 (.X(net1316),
    .A(_1666_));
 sg13g2_buf_2 fanout1317 (.A(net1320),
    .X(net1317));
 sg13g2_buf_2 fanout1318 (.A(net1320),
    .X(net1318));
 sg13g2_buf_2 fanout1319 (.A(net1320),
    .X(net1319));
 sg13g2_buf_2 fanout1320 (.A(net1325),
    .X(net1320));
 sg13g2_buf_2 fanout1321 (.A(net1325),
    .X(net1321));
 sg13g2_buf_2 fanout1322 (.A(net1324),
    .X(net1322));
 sg13g2_buf_2 fanout1323 (.A(net1324),
    .X(net1323));
 sg13g2_buf_2 fanout1324 (.A(net1325),
    .X(net1324));
 sg13g2_buf_2 fanout1325 (.A(_1059_),
    .X(net1325));
 sg13g2_buf_4 fanout1326 (.X(net1326),
    .A(_2920_));
 sg13g2_buf_4 fanout1327 (.X(net1327),
    .A(_2916_));
 sg13g2_buf_4 fanout1328 (.X(net1328),
    .A(_2886_));
 sg13g2_buf_4 fanout1329 (.X(net1329),
    .A(_1654_));
 sg13g2_buf_2 fanout1330 (.A(_1654_),
    .X(net1330));
 sg13g2_buf_2 fanout1331 (.A(net1332),
    .X(net1331));
 sg13g2_buf_2 fanout1332 (.A(net1333),
    .X(net1332));
 sg13g2_buf_2 fanout1333 (.A(_3183_),
    .X(net1333));
 sg13g2_buf_4 fanout1334 (.X(net1334),
    .A(net1335));
 sg13g2_buf_2 fanout1335 (.A(_3100_),
    .X(net1335));
 sg13g2_buf_2 fanout1336 (.A(_2972_),
    .X(net1336));
 sg13g2_buf_4 fanout1337 (.X(net1337),
    .A(_2912_));
 sg13g2_buf_2 fanout1338 (.A(net1339),
    .X(net1338));
 sg13g2_buf_2 fanout1339 (.A(_2908_),
    .X(net1339));
 sg13g2_buf_4 fanout1340 (.X(net1340),
    .A(net1341));
 sg13g2_buf_2 fanout1341 (.A(_2904_),
    .X(net1341));
 sg13g2_buf_4 fanout1342 (.X(net1342),
    .A(_2900_));
 sg13g2_buf_4 fanout1343 (.X(net1343),
    .A(_2895_));
 sg13g2_buf_4 fanout1344 (.X(net1344),
    .A(net1345));
 sg13g2_buf_2 fanout1345 (.A(_2890_),
    .X(net1345));
 sg13g2_buf_4 fanout1346 (.X(net1346),
    .A(_2881_));
 sg13g2_buf_4 fanout1347 (.X(net1347),
    .A(_2876_));
 sg13g2_buf_4 fanout1348 (.X(net1348),
    .A(_1873_));
 sg13g2_buf_2 fanout1349 (.A(_1873_),
    .X(net1349));
 sg13g2_buf_4 fanout1350 (.X(net1350),
    .A(_1545_));
 sg13g2_buf_2 fanout1351 (.A(net1354),
    .X(net1351));
 sg13g2_buf_2 fanout1352 (.A(net1354),
    .X(net1352));
 sg13g2_buf_1 fanout1353 (.A(net1354),
    .X(net1353));
 sg13g2_buf_2 fanout1354 (.A(_2957_),
    .X(net1354));
 sg13g2_buf_4 fanout1355 (.X(net1355),
    .A(_2871_));
 sg13g2_buf_4 fanout1356 (.X(net1356),
    .A(_2866_));
 sg13g2_buf_4 fanout1357 (.X(net1357),
    .A(_2861_));
 sg13g2_buf_1 fanout1358 (.A(_2861_),
    .X(net1358));
 sg13g2_buf_2 fanout1359 (.A(_2597_),
    .X(net1359));
 sg13g2_buf_1 fanout1360 (.A(_2597_),
    .X(net1360));
 sg13g2_buf_2 fanout1361 (.A(_1856_),
    .X(net1361));
 sg13g2_buf_2 fanout1362 (.A(_1846_),
    .X(net1362));
 sg13g2_buf_4 fanout1363 (.X(net1363),
    .A(_1987_));
 sg13g2_buf_2 fanout1364 (.A(_1848_),
    .X(net1364));
 sg13g2_buf_2 fanout1365 (.A(net1367),
    .X(net1365));
 sg13g2_buf_1 fanout1366 (.A(net1367),
    .X(net1366));
 sg13g2_buf_2 fanout1367 (.A(_1019_),
    .X(net1367));
 sg13g2_buf_4 fanout1368 (.X(net1368),
    .A(_1516_));
 sg13g2_buf_2 fanout1369 (.A(net1370),
    .X(net1369));
 sg13g2_buf_2 fanout1370 (.A(net1371),
    .X(net1370));
 sg13g2_buf_2 fanout1371 (.A(_1165_),
    .X(net1371));
 sg13g2_buf_2 fanout1372 (.A(_3182_),
    .X(net1372));
 sg13g2_buf_2 fanout1373 (.A(_2655_),
    .X(net1373));
 sg13g2_buf_2 fanout1374 (.A(_2596_),
    .X(net1374));
 sg13g2_buf_2 fanout1375 (.A(net1376),
    .X(net1375));
 sg13g2_buf_2 fanout1376 (.A(net1377),
    .X(net1376));
 sg13g2_buf_2 fanout1377 (.A(_1399_),
    .X(net1377));
 sg13g2_buf_4 fanout1378 (.X(net1378),
    .A(net1379));
 sg13g2_buf_1 fanout1379 (.A(net1380),
    .X(net1379));
 sg13g2_buf_2 fanout1380 (.A(_1390_),
    .X(net1380));
 sg13g2_buf_2 fanout1381 (.A(\s_m_pushdata_endpoint[1] ),
    .X(net1381));
 sg13g2_buf_2 fanout1382 (.A(net1383),
    .X(net1382));
 sg13g2_buf_2 fanout1383 (.A(net1384),
    .X(net1383));
 sg13g2_buf_2 fanout1384 (.A(net1385),
    .X(net1384));
 sg13g2_buf_4 fanout1385 (.X(net1385),
    .A(_1002_));
 sg13g2_buf_2 fanout1386 (.A(_0787_),
    .X(net1386));
 sg13g2_buf_2 fanout1387 (.A(net1388),
    .X(net1387));
 sg13g2_buf_2 fanout1388 (.A(_1770_),
    .X(net1388));
 sg13g2_buf_4 fanout1389 (.X(net1389),
    .A(net1391));
 sg13g2_buf_2 fanout1390 (.A(net1391),
    .X(net1390));
 sg13g2_buf_4 fanout1391 (.X(net1391),
    .A(_1406_));
 sg13g2_buf_4 fanout1392 (.X(net1392),
    .A(_1039_));
 sg13g2_buf_2 fanout1393 (.A(_1038_),
    .X(net1393));
 sg13g2_buf_2 fanout1394 (.A(_1028_),
    .X(net1394));
 sg13g2_buf_2 fanout1395 (.A(_1028_),
    .X(net1395));
 sg13g2_buf_4 fanout1396 (.X(net1396),
    .A(net1397));
 sg13g2_buf_2 fanout1397 (.A(_0993_),
    .X(net1397));
 sg13g2_buf_2 fanout1398 (.A(_0784_),
    .X(net1398));
 sg13g2_buf_4 fanout1399 (.X(net1399),
    .A(_2809_));
 sg13g2_buf_2 fanout1400 (.A(_2774_),
    .X(net1400));
 sg13g2_buf_2 fanout1401 (.A(_2774_),
    .X(net1401));
 sg13g2_buf_2 fanout1402 (.A(net1403),
    .X(net1402));
 sg13g2_buf_4 fanout1403 (.X(net1403),
    .A(net1404));
 sg13g2_buf_2 fanout1404 (.A(_1724_),
    .X(net1404));
 sg13g2_buf_2 fanout1405 (.A(net1406),
    .X(net1405));
 sg13g2_buf_2 fanout1406 (.A(_1094_),
    .X(net1406));
 sg13g2_buf_2 fanout1407 (.A(_3181_),
    .X(net1407));
 sg13g2_buf_4 fanout1408 (.X(net1408),
    .A(net1409));
 sg13g2_buf_1 fanout1409 (.A(_3177_),
    .X(net1409));
 sg13g2_buf_4 fanout1410 (.X(net1410),
    .A(_2838_));
 sg13g2_buf_2 fanout1411 (.A(net1412),
    .X(net1411));
 sg13g2_buf_2 fanout1412 (.A(_2593_),
    .X(net1412));
 sg13g2_buf_2 fanout1413 (.A(_2591_),
    .X(net1413));
 sg13g2_buf_2 fanout1414 (.A(_1206_),
    .X(net1414));
 sg13g2_buf_4 fanout1415 (.X(net1415),
    .A(_1371_));
 sg13g2_buf_2 fanout1416 (.A(net1417),
    .X(net1416));
 sg13g2_buf_1 fanout1417 (.A(_1069_),
    .X(net1417));
 sg13g2_buf_2 fanout1418 (.A(net1420),
    .X(net1418));
 sg13g2_buf_2 fanout1419 (.A(net1420),
    .X(net1419));
 sg13g2_buf_2 fanout1420 (.A(_0943_),
    .X(net1420));
 sg13g2_buf_2 fanout1421 (.A(net1422),
    .X(net1421));
 sg13g2_buf_4 fanout1422 (.X(net1422),
    .A(_0942_));
 sg13g2_buf_4 fanout1423 (.X(net1423),
    .A(net1425));
 sg13g2_buf_2 fanout1424 (.A(net1425),
    .X(net1424));
 sg13g2_buf_4 fanout1425 (.X(net1425),
    .A(_0942_));
 sg13g2_buf_4 fanout1426 (.X(net1426),
    .A(_0941_));
 sg13g2_buf_2 fanout1427 (.A(_0940_),
    .X(net1427));
 sg13g2_buf_2 fanout1428 (.A(_0938_),
    .X(net1428));
 sg13g2_buf_4 fanout1429 (.X(net1429),
    .A(net1433));
 sg13g2_buf_4 fanout1430 (.X(net1430),
    .A(net1431));
 sg13g2_buf_2 fanout1431 (.A(net1432),
    .X(net1431));
 sg13g2_buf_2 fanout1432 (.A(net1433),
    .X(net1432));
 sg13g2_buf_2 fanout1433 (.A(_0811_),
    .X(net1433));
 sg13g2_buf_4 fanout1434 (.X(net1434),
    .A(_0804_));
 sg13g2_buf_2 fanout1435 (.A(_0803_),
    .X(net1435));
 sg13g2_buf_2 fanout1436 (.A(net1437),
    .X(net1436));
 sg13g2_buf_2 fanout1437 (.A(\usbfunction0.scl_usbgpiophy0.scl_recoverdatadifferential0.scl_recoverdatadifferential_equalsampling_sky1300.n7861_o ),
    .X(net1437));
 sg13g2_buf_4 fanout1438 (.X(net1438),
    .A(_3218_));
 sg13g2_buf_2 fanout1439 (.A(_3218_),
    .X(net1439));
 sg13g2_buf_4 fanout1440 (.X(net1440),
    .A(net1441));
 sg13g2_buf_2 fanout1441 (.A(net1442),
    .X(net1441));
 sg13g2_buf_2 fanout1442 (.A(net1443),
    .X(net1442));
 sg13g2_buf_4 fanout1443 (.X(net1443),
    .A(_3218_));
 sg13g2_buf_2 fanout1444 (.A(net1449),
    .X(net1444));
 sg13g2_buf_2 fanout1445 (.A(net1449),
    .X(net1445));
 sg13g2_buf_4 fanout1446 (.X(net1446),
    .A(net1447));
 sg13g2_buf_2 fanout1447 (.A(net1448),
    .X(net1447));
 sg13g2_buf_4 fanout1448 (.X(net1448),
    .A(net1449));
 sg13g2_buf_4 fanout1449 (.X(net1449),
    .A(_3217_));
 sg13g2_buf_2 fanout1450 (.A(_3217_),
    .X(net1450));
 sg13g2_buf_4 fanout1451 (.X(net1451),
    .A(_0731_));
 sg13g2_buf_4 fanout1452 (.X(net1452),
    .A(net1454));
 sg13g2_buf_2 fanout1453 (.A(net1454),
    .X(net1453));
 sg13g2_buf_4 fanout1454 (.X(net1454),
    .A(_0688_));
 sg13g2_buf_4 fanout1455 (.X(net1455),
    .A(net1456));
 sg13g2_buf_2 fanout1456 (.A(net1457),
    .X(net1456));
 sg13g2_buf_4 fanout1457 (.X(net1457),
    .A(_0687_));
 sg13g2_buf_4 fanout1458 (.X(net1458),
    .A(net1459));
 sg13g2_buf_4 fanout1459 (.X(net1459),
    .A(net1460));
 sg13g2_buf_4 fanout1460 (.X(net1460),
    .A(_0685_));
 sg13g2_buf_2 fanout1461 (.A(\scl_uartrx0.s_m_value[1] ),
    .X(net1461));
 sg13g2_buf_4 fanout1462 (.X(net1462),
    .A(net1464));
 sg13g2_buf_2 fanout1463 (.A(net1464),
    .X(net1463));
 sg13g2_buf_4 fanout1464 (.X(net1464),
    .A(net1631));
 sg13g2_buf_2 fanout1465 (.A(net1466),
    .X(net1465));
 sg13g2_buf_4 fanout1466 (.X(net1466),
    .A(net1467));
 sg13g2_buf_2 fanout1467 (.A(net1681),
    .X(net1467));
 sg13g2_buf_2 fanout1468 (.A(net1470),
    .X(net1468));
 sg13g2_buf_1 fanout1469 (.A(net1470),
    .X(net1469));
 sg13g2_buf_4 fanout1470 (.X(net1470),
    .A(net1715));
 sg13g2_buf_4 fanout1471 (.X(net1471),
    .A(net1473));
 sg13g2_buf_2 fanout1472 (.A(net1473),
    .X(net1472));
 sg13g2_buf_4 fanout1473 (.X(net1473),
    .A(net1712));
 sg13g2_buf_2 fanout1474 (.A(net1476),
    .X(net1474));
 sg13g2_buf_2 fanout1475 (.A(net1476),
    .X(net1475));
 sg13g2_buf_4 fanout1476 (.X(net1476),
    .A(net1864));
 sg13g2_buf_2 fanout1477 (.A(net1594),
    .X(net1477));
 sg13g2_buf_2 fanout1478 (.A(net1645),
    .X(net1478));
 sg13g2_buf_2 fanout1479 (.A(net1645),
    .X(net1479));
 sg13g2_buf_2 fanout1480 (.A(net1664),
    .X(net1480));
 sg13g2_buf_1 fanout1481 (.A(\usbfunction0.n1360_o[1] ),
    .X(net1481));
 sg13g2_buf_4 fanout1482 (.X(net1482),
    .A(net1052));
 sg13g2_buf_4 fanout1483 (.X(net1483),
    .A(net790));
 sg13g2_buf_4 fanout1484 (.X(net1484),
    .A(net966));
 sg13g2_buf_2 fanout1485 (.A(net974),
    .X(net1485));
 sg13g2_buf_2 fanout1486 (.A(net1172),
    .X(net1486));
 sg13g2_buf_4 fanout1487 (.X(net1487),
    .A(net767));
 sg13g2_buf_2 fanout1488 (.A(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.s_m_value[1] ),
    .X(net1488));
 sg13g2_buf_4 fanout1489 (.X(net1489),
    .A(net1491));
 sg13g2_buf_2 fanout1490 (.A(net1491),
    .X(net1490));
 sg13g2_buf_2 fanout1491 (.A(\usbfunction0.functionreset0.n6708_q ),
    .X(net1491));
 sg13g2_buf_4 fanout1492 (.X(net1492),
    .A(\scl_bitbangengine0.n3179_o ));
 sg13g2_buf_4 fanout1493 (.X(net1493),
    .A(net1494));
 sg13g2_buf_2 fanout1494 (.A(\scl_bitbangengine0.n3257_o ),
    .X(net1494));
 sg13g2_buf_2 fanout1495 (.A(net1496),
    .X(net1495));
 sg13g2_buf_2 fanout1496 (.A(net1497),
    .X(net1496));
 sg13g2_buf_4 fanout1497 (.X(net1497),
    .A(\scl_bitbangengine0.n3740_o ));
 sg13g2_buf_4 fanout1498 (.X(net1498),
    .A(\scl_bitbangengine0.n3737_o ));
 sg13g2_buf_2 fanout1499 (.A(net1500),
    .X(net1499));
 sg13g2_buf_2 fanout1500 (.A(net1501),
    .X(net1500));
 sg13g2_buf_2 fanout1501 (.A(\scl_bitbangengine0.n3198_o ),
    .X(net1501));
 sg13g2_buf_4 fanout1502 (.X(net1502),
    .A(\scl_bitbangengine0.n3230_o ));
 sg13g2_buf_2 fanout1503 (.A(net1892),
    .X(net1503));
 sg13g2_buf_4 fanout1504 (.X(net1504),
    .A(net11));
 sg13g2_buf_4 fanout1505 (.X(net1505),
    .A(net1510));
 sg13g2_buf_4 fanout1506 (.X(net1506),
    .A(net1510));
 sg13g2_buf_4 fanout1507 (.X(net1507),
    .A(net1508));
 sg13g2_buf_4 fanout1508 (.X(net1508),
    .A(net1509));
 sg13g2_buf_4 fanout1509 (.X(net1509),
    .A(net1510));
 sg13g2_buf_4 fanout1510 (.X(net1510),
    .A(net1535));
 sg13g2_buf_4 fanout1511 (.X(net1511),
    .A(net1512));
 sg13g2_buf_2 fanout1512 (.A(net1523),
    .X(net1512));
 sg13g2_buf_4 fanout1513 (.X(net1513),
    .A(net1514));
 sg13g2_buf_2 fanout1514 (.A(net1523),
    .X(net1514));
 sg13g2_buf_4 fanout1515 (.X(net1515),
    .A(net1519));
 sg13g2_buf_4 fanout1516 (.X(net1516),
    .A(net1518));
 sg13g2_buf_4 fanout1517 (.X(net1517),
    .A(net1518));
 sg13g2_buf_4 fanout1518 (.X(net1518),
    .A(net1519));
 sg13g2_buf_2 fanout1519 (.A(net1523),
    .X(net1519));
 sg13g2_buf_4 fanout1520 (.X(net1520),
    .A(net1522));
 sg13g2_buf_4 fanout1521 (.X(net1521),
    .A(net1522));
 sg13g2_buf_4 fanout1522 (.X(net1522),
    .A(net1523));
 sg13g2_buf_2 fanout1523 (.A(net1535),
    .X(net1523));
 sg13g2_buf_4 fanout1524 (.X(net1524),
    .A(net1526));
 sg13g2_buf_2 fanout1525 (.A(net1526),
    .X(net1525));
 sg13g2_buf_4 fanout1526 (.X(net1526),
    .A(net1529));
 sg13g2_buf_4 fanout1527 (.X(net1527),
    .A(net1528));
 sg13g2_buf_4 fanout1528 (.X(net1528),
    .A(net1529));
 sg13g2_buf_2 fanout1529 (.A(net1535),
    .X(net1529));
 sg13g2_buf_4 fanout1530 (.X(net1530),
    .A(net1534));
 sg13g2_buf_4 fanout1531 (.X(net1531),
    .A(net1534));
 sg13g2_buf_4 fanout1532 (.X(net1532),
    .A(net1533));
 sg13g2_buf_4 fanout1533 (.X(net1533),
    .A(net1534));
 sg13g2_buf_2 fanout1534 (.A(net1535),
    .X(net1534));
 sg13g2_buf_4 fanout1535 (.X(net1535),
    .A(rst_n));
 sg13g2_buf_4 fanout1536 (.X(net1536),
    .A(net1549));
 sg13g2_buf_4 fanout1537 (.X(net1537),
    .A(net1549));
 sg13g2_buf_4 fanout1538 (.X(net1538),
    .A(net1539));
 sg13g2_buf_2 fanout1539 (.A(net1540),
    .X(net1539));
 sg13g2_buf_2 fanout1540 (.A(net1549),
    .X(net1540));
 sg13g2_buf_4 fanout1541 (.X(net1541),
    .A(net1542));
 sg13g2_buf_4 fanout1542 (.X(net1542),
    .A(net1548));
 sg13g2_buf_4 fanout1543 (.X(net1543),
    .A(net1547));
 sg13g2_buf_2 fanout1544 (.A(net1547),
    .X(net1544));
 sg13g2_buf_4 fanout1545 (.X(net1545),
    .A(net1546));
 sg13g2_buf_4 fanout1546 (.X(net1546),
    .A(net1547));
 sg13g2_buf_2 fanout1547 (.A(net1548),
    .X(net1547));
 sg13g2_buf_4 fanout1548 (.X(net1548),
    .A(net1549));
 sg13g2_buf_2 fanout1549 (.A(rst_n),
    .X(net1549));
 sg13g2_buf_4 fanout1550 (.X(net1550),
    .A(net1552));
 sg13g2_buf_4 fanout1551 (.X(net1551),
    .A(net1552));
 sg13g2_buf_2 fanout1552 (.A(net1554),
    .X(net1552));
 sg13g2_buf_4 fanout1553 (.X(net1553),
    .A(net1554));
 sg13g2_buf_2 fanout1554 (.A(net1559),
    .X(net1554));
 sg13g2_buf_4 fanout1555 (.X(net1555),
    .A(net1559));
 sg13g2_buf_4 fanout1556 (.X(net1556),
    .A(net1559));
 sg13g2_buf_4 fanout1557 (.X(net1557),
    .A(net1558));
 sg13g2_buf_4 fanout1558 (.X(net1558),
    .A(net1559));
 sg13g2_buf_2 fanout1559 (.A(rst_n),
    .X(net1559));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_4 input11 (.X(net11),
    .A(uio_in[2]));
 sg13g2_buf_2 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_2 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[7]),
    .X(net16));
 sg13g2_tiehi _8234__17 (.L_HI(net17));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(delaynet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_buf_2 clkbuf_leaf_0_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_0_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_1_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_1_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_2_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_2_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_3_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_3_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_4_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_4_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_5_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_5_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_6_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_6_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_7_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_7_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_8_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_8_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_9_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_9_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_10_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_10_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_11_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_11_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_12_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_12_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_13_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_13_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_14_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_14_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_15_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_15_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_16_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_16_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_17_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_17_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_18_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_18_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_19_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_19_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_20_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_20_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_21_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_21_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_22_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_22_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_23_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_23_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_24_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_24_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_25_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_25_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_26_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_26_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_27_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_27_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_28_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_28_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_29_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_29_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_30_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_30_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_31_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_31_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_32_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_32_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_33_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_33_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_34_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_34_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_35_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_35_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_36_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_36_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_37_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_37_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_38_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_38_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_39_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_39_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_40_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_40_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_41_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_41_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_42_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_42_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_43_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_43_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_44_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_44_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_45_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_45_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_46_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_46_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_47_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_47_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_48_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_48_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_49_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_49_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_50_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_50_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_51_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_51_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_52_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_52_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_53_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_53_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_54_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_54_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_55_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_55_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_56_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_56_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_57_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_57_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_58_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_58_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_59_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_59_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_60_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_60_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_61_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_61_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_62_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_62_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_63_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_63_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_64_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_64_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_65_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_65_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_66_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_66_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_67_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_67_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_68_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_68_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_69_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_69_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_70_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_70_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_71_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_71_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_72_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_72_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_73_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_73_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_74_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_74_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_75_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_75_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_76_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_76_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_77_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_77_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_78_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_78_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_79_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_79_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_80_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_80_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_81_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_81_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_82_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_82_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_83_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_83_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_84_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_84_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_85_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_85_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_86_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_86_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_87_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_87_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_88_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_88_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_89_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_89_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_90_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_90_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_91_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_91_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_92_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_92_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_93_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_93_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_94_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_94_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_95_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_95_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_96_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_96_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_97_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_97_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_98_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_98_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_99_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_99_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_100_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_100_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_101_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_101_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_102_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_102_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_103_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_103_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_104_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_104_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_105_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_105_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_106_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_106_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_107_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_107_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_108_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_108_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_109_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_109_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_110_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_110_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_111_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_111_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_112_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_112_clk_regs));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_buf_2 clkbuf_5_0__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_1__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_2__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_2__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_3__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_4__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_4__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_5__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_6__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_6__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_7__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_8__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_8__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_9__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_10__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_10__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_11__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_12__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_12__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_13__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_14__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_14__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_15__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_15__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_16__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_16__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_17__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_18__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_18__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_19__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_20__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_20__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_21__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_22__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_22__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_23__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_23__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_24__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_24__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_25__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_26__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_26__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_27__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_28__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_28__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_29__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_29__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_30__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_30__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_31__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_31__leaf_clk_regs));
 sg13g2_buf_2 clkload0 (.A(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_2 clkload1 (.A(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_2 clkload2 (.A(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_2 clkload3 (.A(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_2 clkload4 (.A(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_2 clkload5 (.A(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_2 clkload6 (.A(clknet_5_15__leaf_clk_regs));
 sg13g2_buf_2 clkload7 (.A(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_2 clkload8 (.A(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_2 clkload9 (.A(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_2 clkload10 (.A(clknet_5_23__leaf_clk_regs));
 sg13g2_buf_2 clkload11 (.A(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_2 clkload12 (.A(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_2 clkload13 (.A(clknet_5_29__leaf_clk_regs));
 sg13g2_buf_2 clkload14 (.A(clknet_5_31__leaf_clk_regs));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_112_clk_regs));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_111_clk_regs));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_8_clk_regs));
 sg13g2_inv_4 clkload18 (.A(clknet_leaf_9_clk_regs));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_106_clk_regs));
 sg13g2_inv_1 clkload20 (.A(clknet_leaf_108_clk_regs));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_107_clk_regs));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_15_clk_regs));
 sg13g2_inv_2 clkload23 (.A(clknet_leaf_24_clk_regs));
 sg13g2_inv_1 clkload24 (.A(clknet_leaf_25_clk_regs));
 sg13g2_inv_4 clkload25 (.A(clknet_leaf_26_clk_regs));
 sg13g2_inv_2 clkload26 (.A(clknet_leaf_33_clk_regs));
 sg13g2_inv_4 clkload27 (.A(clknet_leaf_34_clk_regs));
 sg13g2_inv_4 clkload28 (.A(clknet_leaf_43_clk_regs));
 sg13g2_inv_2 clkload29 (.A(clknet_leaf_42_clk_regs));
 sg13g2_inv_4 clkload30 (.A(clknet_leaf_35_clk_regs));
 sg13g2_inv_2 clkload31 (.A(clknet_leaf_38_clk_regs));
 sg13g2_inv_1 clkload32 (.A(clknet_leaf_95_clk_regs));
 sg13g2_inv_4 clkload33 (.A(clknet_leaf_91_clk_regs));
 sg13g2_inv_1 clkload34 (.A(clknet_leaf_96_clk_regs));
 sg13g2_inv_4 clkload35 (.A(clknet_leaf_97_clk_regs));
 sg13g2_inv_2 clkload36 (.A(clknet_leaf_98_clk_regs));
 sg13g2_inv_4 clkload37 (.A(clknet_leaf_78_clk_regs));
 sg13g2_inv_4 clkload38 (.A(clknet_leaf_87_clk_regs));
 sg13g2_inv_2 clkload39 (.A(clknet_leaf_70_clk_regs));
 sg13g2_inv_1 clkload40 (.A(clknet_leaf_81_clk_regs));
 sg13g2_inv_4 clkload41 (.A(clknet_leaf_45_clk_regs));
 sg13g2_inv_1 clkload42 (.A(clknet_leaf_47_clk_regs));
 sg13g2_inv_8 clkload43 (.A(clknet_leaf_74_clk_regs));
 sg13g2_inv_4 clkload44 (.A(clknet_leaf_53_clk_regs));
 sg13g2_inv_1 clkload45 (.A(clknet_leaf_50_clk_regs));
 sg13g2_inv_1 clkload46 (.A(clknet_leaf_71_clk_regs));
 sg13g2_inv_2 clkload47 (.A(clknet_leaf_67_clk_regs));
 sg13g2_inv_1 clkload48 (.A(clknet_leaf_68_clk_regs));
 sg13g2_inv_8 clkload49 (.A(clknet_leaf_58_clk_regs));
 sg13g2_inv_1 clkload50 (.A(clknet_leaf_59_clk_regs));
 sg13g2_buf_2 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(delaynet_1_clk));
 sg13g2_buf_2 delaybuf_1_clk (.A(delaynet_1_clk),
    .X(clknet_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\usbfunction0.s_m_rx_sop ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold2 (.A(\usbfunction0.s_m_rx_data[5] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold3 (.A(\usbfunction0.s_m_rx_data[2] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold4 (.A(\usbfunction0.s_m_rx_data[4] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold5 (.A(\usbfunction0.s_m_rx_data[3] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold6 (.A(\usbfunction0.s_m_rx_data[6] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold7 (.A(\usbfunction0.s_m_rx_data[0] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold8 (.A(\usbfunction0.scl_usbgpiophy0.scl_extendwidth0.scl_counter0.n7984_q[0] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold9 (.A(_1518_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold10 (.A(\usbfunction0.scl_usbgpiophy0.n6533_o ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold11 (.A(\usbfunction0.s_m_rx_data[1] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0152_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold13 (.A(\s_m_status_linestate[1] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0158_),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold15 (.A(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.scl_counter0.n8088_o[0] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold16 (.A(\s_m_status_linestate[0] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold17 (.A(\usbfunction0.scl_usbgpiophy0.scl_pulseextender1.scl_counter0.n8282_q[0] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold18 (.A(\usbfunction0.scl_usbgpiophy0.scl_pulseextender1.scl_counter0.n8260_o[0] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0041_),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold20 (.A(\usbfunction0.rxstream0.n6755_o ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold21 (.A(\usbfunction0.n2334_o[0] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0675_),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold23 (.A(\scl_uartrx0.n6053_o ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0183_),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0045_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold26 (.A(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.scl_counter0.n8088_o[2] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0150_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0177_),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold29 (.A(\usbfunction0.scl_usbgpiophy0.scl_pulseextender1.scl_counter0.n8282_q[1] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold30 (.A(\usbfunction0.scl_usbgpiophy0.n6405_o ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0184_),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0149_),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold33 (.A(\usbfunction0.scl_usbgpiophy0.scl_pulseextender0.scl_counter0.n8243_q[0] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold34 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[5][3] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold35 (.A(\scl_streamarbiter_2.n6192_q ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold36 (.A(\scl_streamarbiter_2.n6171_o ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold37 (.A(\scl_bitbangengine0.s_m_value[1] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold38 (.A(_2694_),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0215_),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold40 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[5][0] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold41 (.A(\usbfunction0.scl_usbgpiophy0.n6651_q ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold42 (.A(_2572_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold43 (.A(\usbfunction0.scl_usbgpiophy0.n6553_o ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold44 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[1][0] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold45 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[9][0] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold46 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[9][1] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold47 (.A(\scl_bitbangengine0.n3865_o ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0255_),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold49 (.A(\scl_fifo0.n2711_o[3] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold50 (.A(_2850_),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0288_),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0154_),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold53 (.A(\scl_fifo1.n6233_o[3] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold54 (.A(\usbfunction0.functionreset0.n6707_q[0] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold55 (.A(\usbfunction0.functionreset0.n6674_o[0] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold56 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[13][0] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold57 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[13][1] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold58 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[13][3] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold59 (.A(\usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8209_q[2] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold60 (.A(_2543_),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold61 (.A(\usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8195_o[2] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold62 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[9][3] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold63 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[5][1] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold64 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[1][3] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold65 (.A(s_m_io14_out),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold66 (.A(s_m_io15_out),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0231_),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold68 (.A(s_m_io13_out),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold69 (.A(\scl_uartrx0.n6119_q ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold70 (.A(\usbfunction0.scl_usbgpiophy0.n6653_q ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0420_),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold72 (.A(\usbfunction0.scl_usbgpiophy0.scl_decodenrzi0.scl_counter0.n7944_q[2] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold73 (.A(_3115_),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold74 (.A(\usbfunction0.functionreset0.n6707_q[9] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold75 (.A(\usbfunction0.functionreset0.n6674_o[9] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold76 (.A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[0] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0571_),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold78 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[8][1] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold79 (.A(\usbfunction0.scl_usbgpiophy0.scl_extendwidth0.scl_counter0.n7984_q[2] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold80 (.A(\usbfunction0.scl_usbgpiophy0.scl_extendwidth0.scl_counter0.n7961_o[2] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold81 (.A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[15] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold82 (.A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[0] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold83 (.A(\scl_uarttx0.scl_baudrategenerator0.n6878_o[0] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold84 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[1][1] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0398_),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold86 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[14][1] ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0302_),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold88 (.A(\usbfunction0.scl_usbgpiophy0.s_out_2[6] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0565_),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold90 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[12][3] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold91 (.A(\usbfunction0.scl_usbgpiophy0.s_out_2[1] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0560_),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold93 (.A(\usbfunction0.n2639_q ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0191_),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold95 (.A(\usbfunction0.n2644_q[15] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold96 (.A(\usbfunction0.n2433_o[15] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold97 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[4][3] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold98 (.A(\usbfunction0.scl_usbgpiophy0.scl_pulseextender1.n7775_q ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0156_),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold100 (.A(_3108_),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold101 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[8][1] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold102 (.A(\usbfunction0.n2644_q[9] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold103 (.A(\usbfunction0.n2433_o[9] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold104 (.A(\usbfunction0.scl_usbgpiophy0.s_out_2[2] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0561_),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold106 (.A(s_m_io10_out),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold107 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[10][1] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold108 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[11][1] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold109 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[0][1] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0342_),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0174_),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0587_),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold113 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[15][1] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0197_),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold115 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[11][4] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold116 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[8][0] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold117 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[11][3] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold118 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[7][3] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold119 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[10][0] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0333_),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold121 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[8][3] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0153_),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold123 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[14][3] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0304_),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold125 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[0][0] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold126 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[0][0] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold127 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[0][3] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold128 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[7][4] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold129 (.A(\scl_fifo0.n2711_o[2] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold130 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[2][0] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold131 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[3][6] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0111_),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold133 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[4][0] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold134 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[6][1] ),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold135 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[7][2] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold136 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[3][1] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0390_),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold138 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[3][4] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0173_),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0567_),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold141 (.A(\scl_fifo0.n2711_o[0] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0285_),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold143 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[14][0] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0301_),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold145 (.A(\s_out_3[0] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold146 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[15][7] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0203_),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold148 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[11][7] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0107_),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold150 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[2][3] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold151 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[3][7] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0396_),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold153 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[8][3] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold154 (.A(\scl_bitbangengine0.n3241_o ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0253_),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold156 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[8][5] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold157 (.A(\s_out_3[7] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold158 (.A(\scl_fifo0.n2711_o[1] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0286_),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold160 (.A(\s_out_3[1] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0300_),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold162 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[6][3] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold163 (.A(\usbfunction0.n2644_q[13] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold164 (.A(\usbfunction0.n2433_o[13] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold165 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[11][0] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold166 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[3][5] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0394_),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold168 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[15][4] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0200_),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold170 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[3][0] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0105_),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold172 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[12][0] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold173 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[15][5] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0201_),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold175 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[7][0] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0116_),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold177 (.A(s_m_io9_out),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold178 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[10][3] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold179 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[11][1] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold180 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[3][2] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold181 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[4][7] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold182 (.A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[14] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold183 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[2][1] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0406_),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0109_),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold186 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[7][7] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold187 (.A(\s_out_3[4] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold188 (.A(_2835_),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0262_),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold190 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[6][0] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold191 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[7][1] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold192 (.A(\scl_bitbangengine0.scl_counter0.n6975_q[0] ),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold193 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[4][1] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold194 (.A(\usbfunction0.scl_usbgpiophy0.s_out_2[0] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0559_),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold196 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[11][5] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold197 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[12][1] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0108_),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold199 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[3][3] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold200 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[11][6] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold201 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[15][4] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold202 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[8][0] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold203 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[7][6] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold204 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[12][2] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold205 (.A(\scl_bitbangengine0.n5920_q[18] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0602_),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold207 (.A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[13] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold208 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[15][2] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold209 (.A(s_m_io2_en),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold210 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[7][3] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold211 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[5][3] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold212 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[7][5] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold213 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[12][1] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold214 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[0][2] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold215 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[8][7] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold216 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[15][0] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0196_),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold218 (.A(\scl_bitbangengine0.n5902_q ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold219 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[9][6] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold220 (.A(s_m_match_delayed1),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0421_),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0110_),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold223 (.A(\scl_bitbangengine0.s_m_value[0] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0214_),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold225 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[14][6] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold226 (.A(n347_q),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold227 (.A(_2857_),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold228 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[8][6] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold229 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[3][3] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold230 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[6][5] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold231 (.A(s_m_io1_en),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold232 (.A(\usbfunction0.n2644_q[7] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold233 (.A(\usbfunction0.n2433_o[7] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold234 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[14][0] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold235 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[3][4] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold236 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[14][6] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold237 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[3][1] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold238 (.A(\s_m_packetdata_2_rewired[8] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0606_),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold240 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[8][4] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold241 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[11][7] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold242 (.A(\usbfunction0.n2644_q[10] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold243 (.A(\usbfunction0.n2433_o[10] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold244 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[11][2] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold245 (.A(\usbfunction0.n2644_q[8] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold246 (.A(\usbfunction0.n2433_o[8] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold247 (.A(\usbfunction0.n2644_q[6] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold248 (.A(\usbfunction0.n2433_o[6] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold249 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[2][0] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold250 (.A(\usbfunction0.scl_usbgpiophy0.scl_decodenrzi0.n7166_q ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold251 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[13][4] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold252 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[4][4] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold253 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[1][6] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold254 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[14][7] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold255 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[12][3] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0157_),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold257 (.A(_2519_),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold258 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[2][5] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold259 (.A(\s_out_3[2] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0218_),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold261 (.A(\usbfunction0.n2481_o[26] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0640_),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold263 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[10][5] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold264 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[7][5] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold265 (.A(\usbfunction0.functionreset0.n6707_q[3] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold266 (.A(_2158_),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold267 (.A(\usbfunction0.functionreset0.n6674_o[3] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold268 (.A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[7] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0577_),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold270 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[7][6] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold271 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[15][7] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold272 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[12][5] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold273 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[1][1] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold274 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[15][3] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold275 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[9][4] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold276 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[0][4] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold277 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[13][1] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold278 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[5][5] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold279 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[2][1] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold280 (.A(\usbfunction0.functionreset0.in_unnamed_2[1] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold281 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[15][3] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0199_),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold283 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[3][2] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold284 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[15][1] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold285 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[11][5] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold286 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[4][3] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold287 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[13][0] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold288 (.A(\usbfunction0.n2644_q[14] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold289 (.A(\usbfunction0.n2433_o[14] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold290 (.A(\scl_bitbangengine0.n5921_q[6] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold291 (.A(s_m_io2_out),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0114_),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold293 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[12][4] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold294 (.A(\scl_bitbangengine0.n3663_o[2] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold295 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[10][2] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold296 (.A(s_m_io4_en),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold297 (.A(_0252_),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0112_),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold299 (.A(_0164_),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold300 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[5][6] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold301 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[14][3] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold302 (.A(\scl_bitbangengine0.n5921_q[2] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold303 (.A(\usbfunction0.scl_usbgpiophy0.s_out_2[7] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0566_),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold305 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[13][3] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold306 (.A(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.in_in_valid ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold307 (.A(_2528_),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold308 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[0][3] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold309 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[6][0] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold310 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[10][0] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0104_),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0103_),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold313 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[7][1] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0102_),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold315 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[9][1] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold316 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[0][5] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold317 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[1][0] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold318 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[12][7] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold319 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[15][5] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold320 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[15][0] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold321 (.A(s_m_io0_en),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold322 (.A(_2842_),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0275_),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold324 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[6][1] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold325 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[8][2] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold326 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[11][0] ),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold327 (.A(\scl_bitbangengine0.n3663_o[6] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold328 (.A(_0271_),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold329 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[10][7] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold330 (.A(\scl_bitbangengine0.n5923_q ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold331 (.A(_0230_),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold332 (.A(s_m_io1_opendrain),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold333 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[4][1] ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold334 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[9][2] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold335 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[2][2] ),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold336 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[14][1] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0113_),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold338 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[9][0] ),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold339 (.A(\s_out_3[5] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0219_),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold341 (.A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[12] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold342 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[1][3] ),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold343 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[7][4] ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold344 (.A(\usbfunction0.n2481_o[55] ),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0661_),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold346 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[7][7] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold347 (.A(\n353_q[0] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold348 (.A(\n352_o[0] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold349 (.A(\scl_uartrx0.n6074_o ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold350 (.A(_0106_),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold351 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[15][2] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold352 (.A(\scl_bitbangengine0.n5920_q[14] ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold353 (.A(_0598_),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold354 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[10][4] ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold355 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[4][2] ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold356 (.A(s_m_io0_out),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0256_),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold358 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[1][5] ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold359 (.A(s_m_io0_opendrain),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold360 (.A(_2818_),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold361 (.A(_0250_),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold362 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[9][7] ),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold363 (.A(\scl_fifo1.n6323_q[2] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold364 (.A(\scl_fifo1.n6239_o[2] ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold365 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[0][6] ),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold366 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[1][2] ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold367 (.A(\usbfunction0.scl_usbgpiophy0.scl_addeopdeferred0.scl_eraselastbeat0.n8041_q ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold368 (.A(\usbfunction0.n2644_q[1] ),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold369 (.A(\usbfunction0.n2433_o[1] ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold370 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[13][5] ),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold371 (.A(\usbfunction0.n2644_q[5] ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold372 (.A(\usbfunction0.n2433_o[5] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold373 (.A(\usbfunction0.scl_usbgpiophy0.s_out_2[4] ),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold374 (.A(_0563_),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold375 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[5][0] ),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold376 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[12][6] ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold377 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[6][3] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold378 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[13][7] ),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold379 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[2][3] ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold380 (.A(\usbfunction0.n2644_q[11] ),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold381 (.A(\usbfunction0.n2433_o[11] ),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0115_),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold383 (.A(\usbfunction0.n2637_q ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold384 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[3][7] ),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold385 (.A(\scl_bitbangengine0.n5904_q ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold386 (.A(_0241_),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold387 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[14][4] ),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold388 (.A(_0147_),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold389 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[11][6] ),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold390 (.A(\usbfunction0.n2651_q[7] ),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold391 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[4][0] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold392 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[5][7] ),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold393 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[7][2] ),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold394 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[14][2] ),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold395 (.A(\scl_bitbangengine0.s_m_value[2] ),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold396 (.A(_0216_),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold397 (.A(\usbfunction0.n2644_q[4] ),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold398 (.A(\usbfunction0.n2433_o[4] ),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold399 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[0][7] ),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold400 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[6][7] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold401 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[5][1] ),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold402 (.A(_0134_),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold403 (.A(\scl_bitbangengine0.n5462_o[0] ),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold404 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[2][7] ),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold405 (.A(\usbfunction0.functionreset0.in_unnamed_2[3] ),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold406 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[1][5] ),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold407 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[9][2] ),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold408 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[6][2] ),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold409 (.A(\scl_uartrx0.n6090_o ),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold410 (.A(\usbfunction0.n2644_q[12] ),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold411 (.A(\usbfunction0.n2433_o[12] ),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold412 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[1][4] ),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold413 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[1][7] ),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold414 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[13][6] ),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold415 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[15][6] ),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold416 (.A(n153_o),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold417 (.A(_0244_),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold418 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[9][7] ),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold419 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[3][6] ),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold420 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[10][1] ),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold421 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[5][2] ),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold422 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[9][3] ),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold423 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[11][4] ),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold424 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[11][3] ),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold425 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[13][4] ),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold426 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[12][0] ),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold427 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[0][1] ),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold428 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[11][2] ),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold429 (.A(\usbfunction0.functionreset0.in_unnamed_2[2] ),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold430 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[13][5] ),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold431 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[14][5] ),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold432 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[6][4] ),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold433 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[4][6] ),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold434 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[9][5] ),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold435 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[13][2] ),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold436 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[6][6] ),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold437 (.A(\usbfunction0.n2481_o[25] ),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold438 (.A(_0631_),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold439 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[13][2] ),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold440 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[2][6] ),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold441 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[5][6] ),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold442 (.A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[5] ),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold443 (.A(_0575_),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold444 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[5][4] ),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold445 (.A(\usbfunction0.n2481_o[24] ),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold446 (.A(_0630_),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold447 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[9][4] ),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold448 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[2][4] ),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold449 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[5][2] ),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold450 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[1][2] ),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold451 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[10][6] ),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold452 (.A(s_m_io5_en),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold453 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[9][5] ),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold454 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[13][7] ),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold455 (.A(\usbfunction0.scl_usbgpiophy0.scl_addeopdeferred0.n7349_q ),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold456 (.A(_0080_),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold457 (.A(_1930_),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold458 (.A(\scl_bitbangengine0.n5917_q ),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold459 (.A(_0257_),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold460 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[4][5] ),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold461 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[13][6] ),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold462 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[7][0] ),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold463 (.A(\scl_uarttx0.n2884_o ),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold464 (.A(\scl_uarttx0.scl_counter0.n6919_o[3] ),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold465 (.A(s_m_io5_opendrain),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold466 (.A(_0245_),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold467 (.A(\usbfunction0.n2645_q[2] ),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold468 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[3][0] ),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold469 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[5][5] ),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold470 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[1][4] ),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold471 (.A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[9] ),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold472 (.A(_0579_),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold473 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[5][7] ),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold474 (.A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[3] ),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold475 (.A(_0573_),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold476 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[1][7] ),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold477 (.A(\usbfunction0.scl_usbgpiophy0.scl_pulseextender0.n7750_q ),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold478 (.A(\usbfunction0.scl_usbgpiophy0.scl_pulseextender0.n7741_o ),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold479 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[3][5] ),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold480 (.A(\usbfunction0.scl_usbgpiophy0.s_out_2[3] ),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold481 (.A(_0562_),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold482 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[15][6] ),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold483 (.A(_0202_),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold484 (.A(s_m_io12_out),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold485 (.A(\scl_bitbangengine0.n5903_q ),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold486 (.A(\usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8209_q[0] ),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold487 (.A(s_m_io11_out),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold488 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[10][3] ),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold489 (.A(\usbfunction0.n2481_o[51] ),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold490 (.A(_0657_),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold491 (.A(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7657_q ),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold492 (.A(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7634_o ),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold493 (.A(\scl_bitbangengine0.n5909_q ),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold494 (.A(\usbfunction0.scl_usbgpiophy0.n6411_o ),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold495 (.A(_0155_),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold496 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[1][6] ),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold497 (.A(_0129_),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold498 (.A(\scl_fifo0.n2697_o[4] ),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold499 (.A(\usbfunction0.n2644_q[2] ),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold500 (.A(\usbfunction0.n2433_o[2] ),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold501 (.A(\usbfunction0.scl_usbgpiophy0.scl_decodenrzi0.scl_counter0.n7944_q[1] ),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold502 (.A(s_m_io2_opendrain),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold503 (.A(_0261_),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold504 (.A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[4] ),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold505 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[5][4] ),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold506 (.A(\usbfunction0.scl_usbgpiophy0.scl_pulseextender0.scl_counter0.n8243_q[1] ),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold507 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[10][6] ),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold508 (.A(\scl_bitbangengine0.n5920_q[6] ),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold509 (.A(_0207_),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold510 (.A(_0076_),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold511 (.A(_1923_),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold512 (.A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[11] ),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold513 (.A(\usbfunction0.n2642_q[1] ),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold514 (.A(\s_m_pushdata_endpoint[1] ),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold515 (.A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[6] ),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold516 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[6][2] ),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold517 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[4][4] ),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold518 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[10][7] ),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold519 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[6][6] ),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold520 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[9][6] ),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold521 (.A(\usbfunction0.n2481_o[52] ),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold522 (.A(_0658_),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold523 (.A(\usbfunction0.n2481_o[27] ),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold524 (.A(_0633_),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold525 (.A(\scl_bitbangengine0.n5920_q[19] ),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold526 (.A(_0603_),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold527 (.A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[2] ),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold528 (.A(_0572_),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold529 (.A(\scl_fifo0.n2700_o ),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold530 (.A(_0289_),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold531 (.A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[10] ),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold532 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[14][7] ),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold533 (.A(_0308_),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold534 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[10][2] ),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold535 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[12][7] ),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold536 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[10][4] ),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold537 (.A(\scl_bitbangengine0.n5907_q ),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold538 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[8][2] ),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold539 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[2][6] ),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold540 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[10][5] ),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold541 (.A(\n353_q[1] ),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold542 (.A(\n352_o[1] ),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold543 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[12][4] ),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold544 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[6][7] ),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold545 (.A(\n353_q[15] ),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold546 (.A(_0820_),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold547 (.A(\usbfunction0.scl_usbgpiophy0.s_out_2[5] ),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold548 (.A(_0564_),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold549 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[4][6] ),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold550 (.A(_0066_),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold551 (.A(_1904_),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold552 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[8][4] ),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold553 (.A(\n353_q[5] ),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold554 (.A(\n352_o[5] ),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold555 (.A(\usbfunction0.n2481_o[36] ),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold556 (.A(_0650_),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold557 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[0][5] ),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold558 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[6][4] ),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold559 (.A(\scl_bitbangengine0.n5918_q ),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold560 (.A(_0248_),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold561 (.A(\usbfunction0.scl_usbgpiophy0.s_linein ),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold562 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[0][6] ),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold563 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[8][6] ),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold564 (.A(\usbfunction0.n2481_o[29] ),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold565 (.A(_0643_),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold566 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[12][5] ),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold567 (.A(\usbfunction0.scl_usbgpiophy0.n6649_q ),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold568 (.A(\usbfunction0.s_m_rx_eop ),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold569 (.A(\s_out_3[3] ),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold570 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[0][2] ),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold571 (.A(\n353_q[3] ),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold572 (.A(\n352_o[3] ),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold573 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[2][4] ),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold574 (.A(\scl_bitbangengine0.n5920_q[10] ),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold575 (.A(_0570_),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold576 (.A(\scl_fifo1.n6323_q[4] ),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold577 (.A(\scl_fifo1.n6239_o[4] ),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold578 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[12][2] ),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold579 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[4][5] ),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold580 (.A(\usbfunction0.n2481_o[39] ),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold581 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[4][2] ),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold582 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[8][7] ),
    .X(net1111));
 sg13g2_dlygate4sd3_1 hold583 (.A(\n353_q[6] ),
    .X(net1112));
 sg13g2_dlygate4sd3_1 hold584 (.A(\n352_o[6] ),
    .X(net1113));
 sg13g2_dlygate4sd3_1 hold585 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[2][2] ),
    .X(net1114));
 sg13g2_dlygate4sd3_1 hold586 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[6][5] ),
    .X(net1115));
 sg13g2_dlygate4sd3_1 hold587 (.A(\scl_bitbangengine0.s_m_value_2[1] ),
    .X(net1116));
 sg13g2_dlygate4sd3_1 hold588 (.A(_0194_),
    .X(net1117));
 sg13g2_dlygate4sd3_1 hold589 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[4][7] ),
    .X(net1118));
 sg13g2_dlygate4sd3_1 hold590 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[12][6] ),
    .X(net1119));
 sg13g2_dlygate4sd3_1 hold591 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[14][2] ),
    .X(net1120));
 sg13g2_dlygate4sd3_1 hold592 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[8][5] ),
    .X(net1121));
 sg13g2_dlygate4sd3_1 hold593 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[14][5] ),
    .X(net1122));
 sg13g2_dlygate4sd3_1 hold594 (.A(_0306_),
    .X(net1123));
 sg13g2_dlygate4sd3_1 hold595 (.A(\s_m_pushdata_data[3] ),
    .X(net1124));
 sg13g2_dlygate4sd3_1 hold596 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[14][4] ),
    .X(net1125));
 sg13g2_dlygate4sd3_1 hold597 (.A(_0305_),
    .X(net1126));
 sg13g2_dlygate4sd3_1 hold598 (.A(\usbfunction0.n2644_q[3] ),
    .X(net1127));
 sg13g2_dlygate4sd3_1 hold599 (.A(\usbfunction0.n2433_o[3] ),
    .X(net1128));
 sg13g2_dlygate4sd3_1 hold600 (.A(s_m_io5_out),
    .X(net1129));
 sg13g2_dlygate4sd3_1 hold601 (.A(_2817_),
    .X(net1130));
 sg13g2_dlygate4sd3_1 hold602 (.A(_0249_),
    .X(net1131));
 sg13g2_dlygate4sd3_1 hold603 (.A(\usbfunction0.scl_usbgpiophy0.scl_reducewidth0.s_m_value[2] ),
    .X(net1132));
 sg13g2_dlygate4sd3_1 hold604 (.A(_2853_),
    .X(net1133));
 sg13g2_dlygate4sd3_1 hold605 (.A(_0291_),
    .X(net1134));
 sg13g2_dlygate4sd3_1 hold606 (.A(_0139_),
    .X(net1135));
 sg13g2_dlygate4sd3_1 hold607 (.A(\scl_bitbangengine0.n5462_o[5] ),
    .X(net1136));
 sg13g2_dlygate4sd3_1 hold608 (.A(\n353_q[9] ),
    .X(net1137));
 sg13g2_dlygate4sd3_1 hold609 (.A(_0828_),
    .X(net1138));
 sg13g2_dlygate4sd3_1 hold610 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[2][5] ),
    .X(net1139));
 sg13g2_dlygate4sd3_1 hold611 (.A(_0410_),
    .X(net1140));
 sg13g2_dlygate4sd3_1 hold612 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[0][7] ),
    .X(net1141));
 sg13g2_dlygate4sd3_1 hold613 (.A(\usbfunction0.scl_usbgpiophy0.scl_extendwidth0.scl_counter0.n7984_q[1] ),
    .X(net1142));
 sg13g2_dlygate4sd3_1 hold614 (.A(\usbfunction0.scl_usbgpiophy0.scl_extendwidth0.scl_counter0.n7961_o[1] ),
    .X(net1143));
 sg13g2_dlygate4sd3_1 hold615 (.A(\scl_fifo1.n6323_q[1] ),
    .X(net1144));
 sg13g2_dlygate4sd3_1 hold616 (.A(_0280_),
    .X(net1145));
 sg13g2_dlygate4sd3_1 hold617 (.A(_0135_),
    .X(net1146));
 sg13g2_dlygate4sd3_1 hold618 (.A(\scl_bitbangengine0.n5462_o[1] ),
    .X(net1147));
 sg13g2_dlygate4sd3_1 hold619 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[2][7] ),
    .X(net1148));
 sg13g2_dlygate4sd3_1 hold620 (.A(\n353_q[4] ),
    .X(net1149));
 sg13g2_dlygate4sd3_1 hold621 (.A(\n352_o[4] ),
    .X(net1150));
 sg13g2_dlygate4sd3_1 hold622 (.A(\scl_bitbangengine0.n5920_q[11] ),
    .X(net1151));
 sg13g2_dlygate4sd3_1 hold623 (.A(_0595_),
    .X(net1152));
 sg13g2_dlygate4sd3_1 hold624 (.A(_0146_),
    .X(net1153));
 sg13g2_dlygate4sd3_1 hold625 (.A(\usbfunction0.n2098_o ),
    .X(net1154));
 sg13g2_dlygate4sd3_1 hold626 (.A(\usbfunction0.n2481_o[28] ),
    .X(net1155));
 sg13g2_dlygate4sd3_1 hold627 (.A(_0634_),
    .X(net1156));
 sg13g2_dlygate4sd3_1 hold628 (.A(_0082_),
    .X(net1157));
 sg13g2_dlygate4sd3_1 hold629 (.A(_0680_),
    .X(net1158));
 sg13g2_dlygate4sd3_1 hold630 (.A(\usbfunction0.n2481_o[54] ),
    .X(net1159));
 sg13g2_dlygate4sd3_1 hold631 (.A(_0660_),
    .X(net1160));
 sg13g2_dlygate4sd3_1 hold632 (.A(\s_m_packetdata_2_rewired[14] ),
    .X(net1161));
 sg13g2_dlygate4sd3_1 hold633 (.A(_0612_),
    .X(net1162));
 sg13g2_dlygate4sd3_1 hold634 (.A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.n7250_q[8] ),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold635 (.A(\scl_fifo1.n6321_q[4] ),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold636 (.A(_1045_),
    .X(net1165));
 sg13g2_dlygate4sd3_1 hold637 (.A(\scl_bitbangengine0.n5910_q ),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold638 (.A(_2803_),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold639 (.A(_0128_),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold640 (.A(\scl_fifo0.n2746_o ),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold641 (.A(\usbfunction0.scl_usbgpiophy0.n6449_o ),
    .X(net1170));
 sg13g2_dlygate4sd3_1 hold642 (.A(_0027_),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold643 (.A(\s_m_packetdata_2_rewired[9] ),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold644 (.A(_0607_),
    .X(net1560));
 sg13g2_dlygate4sd3_1 hold645 (.A(_0161_),
    .X(net1561));
 sg13g2_dlygate4sd3_1 hold646 (.A(_0190_),
    .X(net1562));
 sg13g2_dlygate4sd3_1 hold647 (.A(_0136_),
    .X(net1563));
 sg13g2_dlygate4sd3_1 hold648 (.A(\scl_bitbangengine0.n5462_o[2] ),
    .X(net1564));
 sg13g2_dlygate4sd3_1 hold649 (.A(\s_m_packetdata_2_rewired[23] ),
    .X(net1565));
 sg13g2_dlygate4sd3_1 hold650 (.A(_0621_),
    .X(net1566));
 sg13g2_dlygate4sd3_1 hold651 (.A(\scl_uartrx0.s_m_value[2] ),
    .X(net1567));
 sg13g2_dlygate4sd3_1 hold652 (.A(_0681_),
    .X(net1568));
 sg13g2_dlygate4sd3_1 hold653 (.A(\scl_fifo0.scl_memory0.physical_memory0.memory[0][4] ),
    .X(net1569));
 sg13g2_dlygate4sd3_1 hold654 (.A(\usbfunction0.n2631_q ),
    .X(net1570));
 sg13g2_dlygate4sd3_1 hold655 (.A(\scl_bitbangengine0.n5920_q[15] ),
    .X(net1571));
 sg13g2_dlygate4sd3_1 hold656 (.A(_0599_),
    .X(net1572));
 sg13g2_dlygate4sd3_1 hold657 (.A(\n353_q[2] ),
    .X(net1573));
 sg13g2_dlygate4sd3_1 hold658 (.A(\n352_o[2] ),
    .X(net1574));
 sg13g2_dlygate4sd3_1 hold659 (.A(\usbfunction0.functionreset0.in_unnamed_2[0] ),
    .X(net1575));
 sg13g2_dlygate4sd3_1 hold660 (.A(_1660_),
    .X(net1576));
 sg13g2_dlygate4sd3_1 hold661 (.A(\scl_bitbangengine0.n5920_q[16] ),
    .X(net1577));
 sg13g2_dlygate4sd3_1 hold662 (.A(\s_m_packetdata_2_rewired[2] ),
    .X(net1578));
 sg13g2_dlygate4sd3_1 hold663 (.A(_0608_),
    .X(net1579));
 sg13g2_dlygate4sd3_1 hold664 (.A(\scl_bitbangengine0.n5921_q[3] ),
    .X(net1580));
 sg13g2_dlygate4sd3_1 hold665 (.A(_0160_),
    .X(net1581));
 sg13g2_dlygate4sd3_1 hold666 (.A(_2533_),
    .X(net1582));
 sg13g2_dlygate4sd3_1 hold667 (.A(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.scl_counter0.n8128_o[1] ),
    .X(net1583));
 sg13g2_dlygate4sd3_1 hold668 (.A(\scl_bitbangengine0.n5920_q[13] ),
    .X(net1584));
 sg13g2_dlygate4sd3_1 hold669 (.A(_0074_),
    .X(net1585));
 sg13g2_dlygate4sd3_1 hold670 (.A(_1918_),
    .X(net1586));
 sg13g2_dlygate4sd3_1 hold671 (.A(\scl_bitbangengine0.n5921_q[5] ),
    .X(net1587));
 sg13g2_dlygate4sd3_1 hold672 (.A(_0037_),
    .X(net1588));
 sg13g2_dlygate4sd3_1 hold673 (.A(_1961_),
    .X(net1589));
 sg13g2_dlygate4sd3_1 hold674 (.A(_0138_),
    .X(net1590));
 sg13g2_dlygate4sd3_1 hold675 (.A(\scl_bitbangengine0.n5462_o[4] ),
    .X(net1591));
 sg13g2_dlygate4sd3_1 hold676 (.A(\usbfunction0.n2481_o[53] ),
    .X(net1592));
 sg13g2_dlygate4sd3_1 hold677 (.A(_0659_),
    .X(net1593));
 sg13g2_dlygate4sd3_1 hold678 (.A(\usbfunction0.n1360_o[3] ),
    .X(net1594));
 sg13g2_dlygate4sd3_1 hold679 (.A(\s_m_packetdata_2_rewired[21] ),
    .X(net1595));
 sg13g2_dlygate4sd3_1 hold680 (.A(\usbfunction0.n1083_o[5] ),
    .X(net1596));
 sg13g2_dlygate4sd3_1 hold681 (.A(\usbfunction0.n2481_o[22] ),
    .X(net1597));
 sg13g2_dlygate4sd3_1 hold682 (.A(_0636_),
    .X(net1598));
 sg13g2_dlygate4sd3_1 hold683 (.A(\usbfunction0.n2481_o[23] ),
    .X(net1599));
 sg13g2_dlygate4sd3_1 hold684 (.A(_0064_),
    .X(net1600));
 sg13g2_dlygate4sd3_1 hold685 (.A(_1900_),
    .X(net1601));
 sg13g2_dlygate4sd3_1 hold686 (.A(\usbfunction0.n2644_q[0] ),
    .X(net1602));
 sg13g2_dlygate4sd3_1 hold687 (.A(\scl_fifo1.n6323_q[3] ),
    .X(net1603));
 sg13g2_dlygate4sd3_1 hold688 (.A(\scl_fifo1.n6239_o[3] ),
    .X(net1604));
 sg13g2_dlygate4sd3_1 hold689 (.A(\scl_bitbangengine0.n5920_q[2] ),
    .X(net1605));
 sg13g2_dlygate4sd3_1 hold690 (.A(_0417_),
    .X(net1606));
 sg13g2_dlygate4sd3_1 hold691 (.A(_0077_),
    .X(net1607));
 sg13g2_dlygate4sd3_1 hold692 (.A(_1926_),
    .X(net1608));
 sg13g2_dlygate4sd3_1 hold693 (.A(\scl_bitbangengine0.scl_counter0.n6954_o[14] ),
    .X(net1609));
 sg13g2_dlygate4sd3_1 hold694 (.A(\n353_q[16] ),
    .X(net1610));
 sg13g2_dlygate4sd3_1 hold695 (.A(\scl_fifo1.n6323_q[0] ),
    .X(net1611));
 sg13g2_dlygate4sd3_1 hold696 (.A(\scl_fifo1.n6239_o[0] ),
    .X(net1612));
 sg13g2_dlygate4sd3_1 hold697 (.A(\usbfunction0.n2640_q[2] ),
    .X(net1613));
 sg13g2_dlygate4sd3_1 hold698 (.A(_0189_),
    .X(net1614));
 sg13g2_dlygate4sd3_1 hold699 (.A(\usbfunction0.n2481_o[32] ),
    .X(net1615));
 sg13g2_dlygate4sd3_1 hold700 (.A(_0646_),
    .X(net1616));
 sg13g2_dlygate4sd3_1 hold701 (.A(\s_m_packetdata_2_rewired[22] ),
    .X(net1617));
 sg13g2_dlygate4sd3_1 hold702 (.A(\scl_fifo1.n6321_q[0] ),
    .X(net1618));
 sg13g2_dlygate4sd3_1 hold703 (.A(_0042_),
    .X(net1619));
 sg13g2_dlygate4sd3_1 hold704 (.A(_0784_),
    .X(net1620));
 sg13g2_dlygate4sd3_1 hold705 (.A(_0140_),
    .X(net1621));
 sg13g2_dlygate4sd3_1 hold706 (.A(\scl_bitbangengine0.n5462_o[6] ),
    .X(net1622));
 sg13g2_dlygate4sd3_1 hold707 (.A(\usbfunction0.n2481_o[30] ),
    .X(net1623));
 sg13g2_dlygate4sd3_1 hold708 (.A(_0644_),
    .X(net1624));
 sg13g2_dlygate4sd3_1 hold709 (.A(\usbfunction0.n1360_o[0] ),
    .X(net1625));
 sg13g2_dlygate4sd3_1 hold710 (.A(_1745_),
    .X(net1626));
 sg13g2_dlygate4sd3_1 hold711 (.A(\s_m_packetdata_2_rewired[7] ),
    .X(net1627));
 sg13g2_dlygate4sd3_1 hold712 (.A(_0613_),
    .X(net1628));
 sg13g2_dlygate4sd3_1 hold713 (.A(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7656_q ),
    .X(net1629));
 sg13g2_dlygate4sd3_1 hold714 (.A(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7508_o ),
    .X(net1630));
 sg13g2_dlygate4sd3_1 hold715 (.A(\s_m_pushdata_data[7] ),
    .X(net1631));
 sg13g2_dlygate4sd3_1 hold716 (.A(\s_m_packetdata_2_rewired[4] ),
    .X(net1632));
 sg13g2_dlygate4sd3_1 hold717 (.A(_0610_),
    .X(net1633));
 sg13g2_dlygate4sd3_1 hold718 (.A(_0148_),
    .X(net1634));
 sg13g2_dlygate4sd3_1 hold719 (.A(\usbfunction0.n2481_o[37] ),
    .X(net1635));
 sg13g2_dlygate4sd3_1 hold720 (.A(_0651_),
    .X(net1636));
 sg13g2_dlygate4sd3_1 hold721 (.A(\usbfunction0.scl_usbgpiophy0.bitstuff0.scl_counter0.n8209_q[1] ),
    .X(net1637));
 sg13g2_dlygate4sd3_1 hold722 (.A(\s_out_3[6] ),
    .X(net1638));
 sg13g2_dlygate4sd3_1 hold723 (.A(_0260_),
    .X(net1639));
 sg13g2_dlygate4sd3_1 hold724 (.A(\usbfunction0.scl_usbgpiophy0.n6437_o ),
    .X(net1640));
 sg13g2_dlygate4sd3_1 hold725 (.A(_0130_),
    .X(net1641));
 sg13g2_dlygate4sd3_1 hold726 (.A(\scl_uarttx0.n2856_o[2] ),
    .X(net1642));
 sg13g2_dlygate4sd3_1 hold727 (.A(_0176_),
    .X(net1643));
 sg13g2_dlygate4sd3_1 hold728 (.A(\usbfunction0.n2481_o[21] ),
    .X(net1644));
 sg13g2_dlygate4sd3_1 hold729 (.A(\usbfunction0.n1360_o[2] ),
    .X(net1645));
 sg13g2_dlygate4sd3_1 hold730 (.A(\scl_bitbangengine0.n5920_q[17] ),
    .X(net1646));
 sg13g2_dlygate4sd3_1 hold731 (.A(\usbfunction0.functionreset0.n6707_q[4] ),
    .X(net1647));
 sg13g2_dlygate4sd3_1 hold732 (.A(_2161_),
    .X(net1648));
 sg13g2_dlygate4sd3_1 hold733 (.A(\usbfunction0.n1360_o[0] ),
    .X(net1649));
 sg13g2_dlygate4sd3_1 hold734 (.A(\usbfunction0.n2481_o[33] ),
    .X(net1650));
 sg13g2_dlygate4sd3_1 hold735 (.A(\scl_bitbangengine0.n5924_q[7] ),
    .X(net1651));
 sg13g2_dlygate4sd3_1 hold736 (.A(\scl_bitbangengine0.n5462_o[7] ),
    .X(net1652));
 sg13g2_dlygate4sd3_1 hold737 (.A(\scl_bitbangengine0.n5921_q[7] ),
    .X(net1653));
 sg13g2_dlygate4sd3_1 hold738 (.A(\usbfunction0.n2640_q[1] ),
    .X(net1654));
 sg13g2_dlygate4sd3_1 hold739 (.A(_0188_),
    .X(net1655));
 sg13g2_dlygate4sd3_1 hold740 (.A(\usbfunction0.n1583_o[2] ),
    .X(net1656));
 sg13g2_dlygate4sd3_1 hold741 (.A(_0062_),
    .X(net1657));
 sg13g2_dlygate4sd3_1 hold742 (.A(_1898_),
    .X(net1658));
 sg13g2_dlygate4sd3_1 hold743 (.A(\scl_bitbangengine0.scl_counter0.n6954_o[2] ),
    .X(net1659));
 sg13g2_dlygate4sd3_1 hold744 (.A(\n353_q[14] ),
    .X(net1660));
 sg13g2_dlygate4sd3_1 hold745 (.A(_0071_),
    .X(net1661));
 sg13g2_dlygate4sd3_1 hold746 (.A(_1913_),
    .X(net1662));
 sg13g2_dlygate4sd3_1 hold747 (.A(_0137_),
    .X(net1663));
 sg13g2_dlygate4sd3_1 hold748 (.A(\usbfunction0.n1360_o[1] ),
    .X(net1664));
 sg13g2_dlygate4sd3_1 hold749 (.A(s_m_io4_opendrain),
    .X(net1665));
 sg13g2_dlygate4sd3_1 hold750 (.A(_0251_),
    .X(net1666));
 sg13g2_dlygate4sd3_1 hold751 (.A(\usbfunction0.n1583_o[1] ),
    .X(net1667));
 sg13g2_dlygate4sd3_1 hold752 (.A(\scl_bitbangengine0.n3663_o[5] ),
    .X(net1668));
 sg13g2_dlygate4sd3_1 hold753 (.A(s_m_io3_en),
    .X(net1669));
 sg13g2_dlygate4sd3_1 hold754 (.A(\usbfunction0.scl_usbgpiophy0.s_m_last ),
    .X(net1670));
 sg13g2_dlygate4sd3_1 hold755 (.A(\usbfunction0.functionreset0.n6707_q[8] ),
    .X(net1671));
 sg13g2_dlygate4sd3_1 hold756 (.A(_2169_),
    .X(net1672));
 sg13g2_dlygate4sd3_1 hold757 (.A(\scl_bitbangengine0.s_m_value_2[0] ),
    .X(net1673));
 sg13g2_dlygate4sd3_1 hold758 (.A(_2582_),
    .X(net1674));
 sg13g2_dlygate4sd3_1 hold759 (.A(\s_m_packetdata_2_rewired[3] ),
    .X(net1675));
 sg13g2_dlygate4sd3_1 hold760 (.A(_0609_),
    .X(net1676));
 sg13g2_dlygate4sd3_1 hold761 (.A(\usbfunction0.functionreset0.n6707_q[1] ),
    .X(net1677));
 sg13g2_dlygate4sd3_1 hold762 (.A(\usbfunction0.functionreset0.n6674_o[1] ),
    .X(net1678));
 sg13g2_dlygate4sd3_1 hold763 (.A(\usbfunction0.functionreset0.n6707_q[5] ),
    .X(net1679));
 sg13g2_dlygate4sd3_1 hold764 (.A(_2163_),
    .X(net1680));
 sg13g2_dlygate4sd3_1 hold765 (.A(\s_m_pushdata_data[6] ),
    .X(net1681));
 sg13g2_dlygate4sd3_1 hold766 (.A(_0159_),
    .X(net1682));
 sg13g2_dlygate4sd3_1 hold767 (.A(\usbfunction0.functionreset0.n6707_q[6] ),
    .X(net1683));
 sg13g2_dlygate4sd3_1 hold768 (.A(_2165_),
    .X(net1684));
 sg13g2_dlygate4sd3_1 hold769 (.A(\usbfunction0.n2481_o[38] ),
    .X(net1685));
 sg13g2_dlygate4sd3_1 hold770 (.A(_0652_),
    .X(net1686));
 sg13g2_dlygate4sd3_1 hold771 (.A(\usbfunction0.functionreset0.in_unnamed_3[6] ),
    .X(net1687));
 sg13g2_dlygate4sd3_1 hold772 (.A(\usbfunction0.n2481_o[17] ),
    .X(net1688));
 sg13g2_dlygate4sd3_1 hold773 (.A(_0623_),
    .X(net1689));
 sg13g2_dlygate4sd3_1 hold774 (.A(s_m_io3_opendrain),
    .X(net1690));
 sg13g2_dlygate4sd3_1 hold775 (.A(\usbfunction0.n2481_o[35] ),
    .X(net1691));
 sg13g2_dlygate4sd3_1 hold776 (.A(\scl_bitbangengine0.n3336_o ),
    .X(net1692));
 sg13g2_dlygate4sd3_1 hold777 (.A(\scl_bitbangengine0.n3663_o[8] ),
    .X(net1693));
 sg13g2_dlygate4sd3_1 hold778 (.A(\usbfunction0.n2640_q[0] ),
    .X(net1694));
 sg13g2_dlygate4sd3_1 hold779 (.A(_0187_),
    .X(net1695));
 sg13g2_dlygate4sd3_1 hold780 (.A(\s_m_packetdata_2_rewired[13] ),
    .X(net1696));
 sg13g2_dlygate4sd3_1 hold781 (.A(\usbfunction0.n1581_o[0] ),
    .X(net1697));
 sg13g2_dlygate4sd3_1 hold782 (.A(_3237_),
    .X(net1698));
 sg13g2_dlygate4sd3_1 hold783 (.A(_0671_),
    .X(net1699));
 sg13g2_dlygate4sd3_1 hold784 (.A(\usbfunction0.functionreset0.n6707_q[7] ),
    .X(net1700));
 sg13g2_dlygate4sd3_1 hold785 (.A(_2167_),
    .X(net1701));
 sg13g2_dlygate4sd3_1 hold786 (.A(\s_m_packetdata_2_rewired[5] ),
    .X(net1702));
 sg13g2_dlygate4sd3_1 hold787 (.A(\usbfunction0.n1359_o[0] ),
    .X(net1703));
 sg13g2_dlygate4sd3_1 hold788 (.A(_0673_),
    .X(net1704));
 sg13g2_dlygate4sd3_1 hold789 (.A(_0065_),
    .X(net1705));
 sg13g2_dlygate4sd3_1 hold790 (.A(_1902_),
    .X(net1706));
 sg13g2_dlygate4sd3_1 hold791 (.A(\scl_bitbangengine0.scl_counter0.n6954_o[4] ),
    .X(net1707));
 sg13g2_dlygate4sd3_1 hold792 (.A(\scl_bitbangengine0.n3663_o[3] ),
    .X(net1708));
 sg13g2_dlygate4sd3_1 hold793 (.A(\usbfunction0.n2651_q[0] ),
    .X(net1709));
 sg13g2_dlygate4sd3_1 hold794 (.A(\usbfunction0.n1583_o[3] ),
    .X(net1710));
 sg13g2_dlygate4sd3_1 hold795 (.A(\scl_bitbangengine0.n5921_q[1] ),
    .X(net1711));
 sg13g2_dlygate4sd3_1 hold796 (.A(\s_m_pushdata_data[4] ),
    .X(net1712));
 sg13g2_dlygate4sd3_1 hold797 (.A(\usbfunction0.scl_usbgpiophy0.scl_addeopdeferred0.scl_eraselastbeat0.n8042_q ),
    .X(net1713));
 sg13g2_dlygate4sd3_1 hold798 (.A(\usbfunction0.scl_usbgpiophy0.scl_addeopdeferred0.scl_eraselastbeat0.n8008_o ),
    .X(net1714));
 sg13g2_dlygate4sd3_1 hold799 (.A(\s_m_pushdata_data[5] ),
    .X(net1715));
 sg13g2_dlygate4sd3_1 hold800 (.A(\scl_bitbangengine0.n5920_q[5] ),
    .X(net1716));
 sg13g2_dlygate4sd3_1 hold801 (.A(\scl_uartrx0.s_m_value[0] ),
    .X(net1717));
 sg13g2_dlygate4sd3_1 hold802 (.A(_0679_),
    .X(net1718));
 sg13g2_dlygate4sd3_1 hold803 (.A(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.s_m_value[3] ),
    .X(net1719));
 sg13g2_dlygate4sd3_1 hold804 (.A(_2538_),
    .X(net1720));
 sg13g2_dlygate4sd3_1 hold805 (.A(\usbfunction0.n2481_o[34] ),
    .X(net1721));
 sg13g2_dlygate4sd3_1 hold806 (.A(\scl_bitbangengine0.n5920_q[1] ),
    .X(net1722));
 sg13g2_dlygate4sd3_1 hold807 (.A(_0416_),
    .X(net1723));
 sg13g2_dlygate4sd3_1 hold808 (.A(\usbfunction0.n2635_q[1] ),
    .X(net1724));
 sg13g2_dlygate4sd3_1 hold809 (.A(_0419_),
    .X(net1725));
 sg13g2_dlygate4sd3_1 hold810 (.A(\scl_bitbangengine0.n5920_q[9] ),
    .X(net1726));
 sg13g2_dlygate4sd3_1 hold811 (.A(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.s_m_value[2] ),
    .X(net1727));
 sg13g2_dlygate4sd3_1 hold812 (.A(_0067_),
    .X(net1728));
 sg13g2_dlygate4sd3_1 hold813 (.A(_1907_),
    .X(net1729));
 sg13g2_dlygate4sd3_1 hold814 (.A(\scl_bitbangengine0.scl_counter0.n6954_o[6] ),
    .X(net1730));
 sg13g2_dlygate4sd3_1 hold815 (.A(\usbfunction0.n1359_o[1] ),
    .X(net1731));
 sg13g2_dlygate4sd3_1 hold816 (.A(_3240_),
    .X(net1732));
 sg13g2_dlygate4sd3_1 hold817 (.A(\usbfunction0.n2313_o[2] ),
    .X(net1733));
 sg13g2_dlygate4sd3_1 hold818 (.A(_0677_),
    .X(net1734));
 sg13g2_dlygate4sd3_1 hold819 (.A(\usbfunction0.scl_usbgpiophy0.combinedbitcrc0.in_unnamed ),
    .X(net1735));
 sg13g2_dlygate4sd3_1 hold820 (.A(_0422_),
    .X(net1736));
 sg13g2_dlygate4sd3_1 hold821 (.A(\scl_uarttx0.n2856_o[0] ),
    .X(net1737));
 sg13g2_dlygate4sd3_1 hold822 (.A(\scl_uarttx0.scl_counter0.n6919_o[0] ),
    .X(net1738));
 sg13g2_dlygate4sd3_1 hold823 (.A(\s_m_packetdata_2_rewired[12] ),
    .X(net1739));
 sg13g2_dlygate4sd3_1 hold824 (.A(_0618_),
    .X(net1740));
 sg13g2_dlygate4sd3_1 hold825 (.A(\usbfunction0.n2635_q[0] ),
    .X(net1741));
 sg13g2_dlygate4sd3_1 hold826 (.A(_3236_),
    .X(net1742));
 sg13g2_dlygate4sd3_1 hold827 (.A(_0670_),
    .X(net1743));
 sg13g2_dlygate4sd3_1 hold828 (.A(\usbfunction0.scl_usbgpiophy0.scl_recoverdatadifferential0.scl_recoverdatadifferential_equalsampling_sky1300.detectsingleended0.n9022_q ),
    .X(net1744));
 sg13g2_dlygate4sd3_1 hold829 (.A(\scl_bitbangengine0.n3663_o[7] ),
    .X(net1745));
 sg13g2_dlygate4sd3_1 hold830 (.A(_0072_),
    .X(net1746));
 sg13g2_dlygate4sd3_1 hold831 (.A(_1916_),
    .X(net1747));
 sg13g2_dlygate4sd3_1 hold832 (.A(\scl_bitbangengine0.scl_counter0.n6954_o[10] ),
    .X(net1748));
 sg13g2_dlygate4sd3_1 hold833 (.A(_0069_),
    .X(net1749));
 sg13g2_dlygate4sd3_1 hold834 (.A(_1909_),
    .X(net1750));
 sg13g2_dlygate4sd3_1 hold835 (.A(\scl_bitbangengine0.n5898_q[2] ),
    .X(net1751));
 sg13g2_dlygate4sd3_1 hold836 (.A(\usbfunction0.n2636_q ),
    .X(net1752));
 sg13g2_dlygate4sd3_1 hold837 (.A(\usbfunction0.n1583_o[5] ),
    .X(net1753));
 sg13g2_dlygate4sd3_1 hold838 (.A(\usbfunction0.functionreset0.n6707_q[2] ),
    .X(net1754));
 sg13g2_dlygate4sd3_1 hold839 (.A(_2157_),
    .X(net1755));
 sg13g2_dlygate4sd3_1 hold840 (.A(\usbfunction0.n2481_o[18] ),
    .X(net1756));
 sg13g2_dlygate4sd3_1 hold841 (.A(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.s_m_value[1] ),
    .X(net1757));
 sg13g2_dlygate4sd3_1 hold842 (.A(_2547_),
    .X(net1758));
 sg13g2_dlygate4sd3_1 hold843 (.A(\s_m_packetdata_2_rewired[20] ),
    .X(net1759));
 sg13g2_dlygate4sd3_1 hold844 (.A(\usbfunction0.n1083_o[4] ),
    .X(net1760));
 sg13g2_dlygate4sd3_1 hold845 (.A(\scl_bitbangengine0.n5921_q[4] ),
    .X(net1761));
 sg13g2_dlygate4sd3_1 hold846 (.A(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7654_q[0] ),
    .X(net1762));
 sg13g2_dlygate4sd3_1 hold847 (.A(_0604_),
    .X(net1763));
 sg13g2_dlygate4sd3_1 hold848 (.A(\usbfunction0.scl_usbgpiophy0.n6646_q ),
    .X(net1764));
 sg13g2_dlygate4sd3_1 hold849 (.A(\usbfunction0.n2642_q[2] ),
    .X(net1765));
 sg13g2_dlygate4sd3_1 hold850 (.A(\scl_bitbangengine0.n5920_q[12] ),
    .X(net1766));
 sg13g2_dlygate4sd3_1 hold851 (.A(\s_m_packetdata_2_rewired[18] ),
    .X(net1767));
 sg13g2_dlygate4sd3_1 hold852 (.A(\usbfunction0.n1583_o[4] ),
    .X(net1768));
 sg13g2_dlygate4sd3_1 hold853 (.A(\scl_fifo1.n6267_o ),
    .X(net1769));
 sg13g2_dlygate4sd3_1 hold854 (.A(\scl_fifo1.n6287_o ),
    .X(net1770));
 sg13g2_dlygate4sd3_1 hold855 (.A(\usbfunction0.n2652_q[3] ),
    .X(net1771));
 sg13g2_dlygate4sd3_1 hold856 (.A(\usbfunction0.n2481_o[20] ),
    .X(net1772));
 sg13g2_dlygate4sd3_1 hold857 (.A(\scl_bitbangengine0.n3663_o[1] ),
    .X(net1773));
 sg13g2_dlygate4sd3_1 hold858 (.A(\scl_bitbangengine0.n5920_q[4] ),
    .X(net1774));
 sg13g2_dlygate4sd3_1 hold859 (.A(\n353_q[17] ),
    .X(net1775));
 sg13g2_dlygate4sd3_1 hold860 (.A(\usbfunction0.n1583_o[6] ),
    .X(net1776));
 sg13g2_dlygate4sd3_1 hold861 (.A(_0094_),
    .X(net1777));
 sg13g2_dlygate4sd3_1 hold862 (.A(\scl_bitbangengine0.n5920_q[3] ),
    .X(net1778));
 sg13g2_dlygate4sd3_1 hold863 (.A(\scl_bitbangengine0.n3663_o[4] ),
    .X(net1779));
 sg13g2_dlygate4sd3_1 hold864 (.A(_0269_),
    .X(net1780));
 sg13g2_dlygate4sd3_1 hold865 (.A(_0079_),
    .X(net1781));
 sg13g2_dlygate4sd3_1 hold866 (.A(_1928_),
    .X(net1782));
 sg13g2_dlygate4sd3_1 hold867 (.A(\usbfunction0.n2481_o[19] ),
    .X(net1783));
 sg13g2_dlygate4sd3_1 hold868 (.A(_0625_),
    .X(net1784));
 sg13g2_dlygate4sd3_1 hold869 (.A(\scl_bitbangengine0.s_m_value_2[2] ),
    .X(net1785));
 sg13g2_dlygate4sd3_1 hold870 (.A(\scl_bitbangengine0.n5920_q[7] ),
    .X(net1786));
 sg13g2_dlygate4sd3_1 hold871 (.A(_0208_),
    .X(net1787));
 sg13g2_dlygate4sd3_1 hold872 (.A(\usbfunction0.functionreset0.in_unnamed_3[2] ),
    .X(net1788));
 sg13g2_dlygate4sd3_1 hold873 (.A(\usbfunction0.functionreset0.in_unnamed_3[1] ),
    .X(net1789));
 sg13g2_dlygate4sd3_1 hold874 (.A(_0962_),
    .X(net1790));
 sg13g2_dlygate4sd3_1 hold875 (.A(\usbfunction0.n1083_o[1] ),
    .X(net1791));
 sg13g2_dlygate4sd3_1 hold876 (.A(\n353_q[8] ),
    .X(net1792));
 sg13g2_dlygate4sd3_1 hold877 (.A(\n353_q[19] ),
    .X(net1793));
 sg13g2_dlygate4sd3_1 hold878 (.A(\s_m_packetdata_2_rewired[10] ),
    .X(net1794));
 sg13g2_dlygate4sd3_1 hold879 (.A(\usbfunction0.n2642_q[3] ),
    .X(net1795));
 sg13g2_dlygate4sd3_1 hold880 (.A(_0075_),
    .X(net1796));
 sg13g2_dlygate4sd3_1 hold881 (.A(_1921_),
    .X(net1797));
 sg13g2_dlygate4sd3_1 hold882 (.A(\usbfunction0.n1583_o[0] ),
    .X(net1798));
 sg13g2_dlygate4sd3_1 hold883 (.A(_0092_),
    .X(net1799));
 sg13g2_dlygate4sd3_1 hold884 (.A(\scl_bitbangengine0.n5898_q[3] ),
    .X(net1800));
 sg13g2_dlygate4sd3_1 hold885 (.A(\scl_bitbangengine0.n5911_q ),
    .X(net1801));
 sg13g2_dlygate4sd3_1 hold886 (.A(_0259_),
    .X(net1802));
 sg13g2_dlygate4sd3_1 hold887 (.A(s_m_packetdata_2_bit_16),
    .X(net1803));
 sg13g2_dlygate4sd3_1 hold888 (.A(\n353_q[18] ),
    .X(net1804));
 sg13g2_dlygate4sd3_1 hold889 (.A(\n352_o[18] ),
    .X(net1805));
 sg13g2_dlygate4sd3_1 hold890 (.A(\usbfunction0.n1581_o[1] ),
    .X(net1806));
 sg13g2_dlygate4sd3_1 hold891 (.A(_3238_),
    .X(net1807));
 sg13g2_dlygate4sd3_1 hold892 (.A(_0672_),
    .X(net1808));
 sg13g2_dlygate4sd3_1 hold893 (.A(\usbfunction0.functionreset0.in_unnamed_3[0] ),
    .X(net1809));
 sg13g2_dlygate4sd3_1 hold894 (.A(\n353_q[7] ),
    .X(net1810));
 sg13g2_dlygate4sd3_1 hold895 (.A(n349_q),
    .X(net1811));
 sg13g2_dlygate4sd3_1 hold896 (.A(_0087_),
    .X(net1812));
 sg13g2_dlygate4sd3_1 hold897 (.A(_0070_),
    .X(net1813));
 sg13g2_dlygate4sd3_1 hold898 (.A(_1911_),
    .X(net1814));
 sg13g2_dlygate4sd3_1 hold899 (.A(\scl_bitbangengine0.scl_counter0.n6954_o[8] ),
    .X(net1815));
 sg13g2_dlygate4sd3_1 hold900 (.A(\n353_q[13] ),
    .X(net1816));
 sg13g2_dlygate4sd3_1 hold901 (.A(\usbfunction0.n2313_o[1] ),
    .X(net1817));
 sg13g2_dlygate4sd3_1 hold902 (.A(_3250_),
    .X(net1818));
 sg13g2_dlygate4sd3_1 hold903 (.A(_0676_),
    .X(net1819));
 sg13g2_dlygate4sd3_1 hold904 (.A(\usbfunction0.scl_usbgpiophy0.generatetxcrcappend0.n7654_q[1] ),
    .X(net1820));
 sg13g2_dlygate4sd3_1 hold905 (.A(_3215_),
    .X(net1821));
 sg13g2_dlygate4sd3_1 hold906 (.A(_0091_),
    .X(net1822));
 sg13g2_dlygate4sd3_1 hold907 (.A(_1603_),
    .X(net1823));
 sg13g2_dlygate4sd3_1 hold908 (.A(\usbfunction0.functionreset0.in_unnamed[6] ),
    .X(net1824));
 sg13g2_dlygate4sd3_1 hold909 (.A(\usbfunction0.n665_o[6] ),
    .X(net1825));
 sg13g2_dlygate4sd3_1 hold910 (.A(\usbfunction0.n2481_o[16] ),
    .X(net1826));
 sg13g2_dlygate4sd3_1 hold911 (.A(\usbfunction0.functionreset0.in_unnamed[1] ),
    .X(net1827));
 sg13g2_dlygate4sd3_1 hold912 (.A(\usbfunction0.n665_o[1] ),
    .X(net1828));
 sg13g2_dlygate4sd3_1 hold913 (.A(\n353_q[20] ),
    .X(net1829));
 sg13g2_dlygate4sd3_1 hold914 (.A(\s_m_packetdata_2_rewired[11] ),
    .X(net1830));
 sg13g2_dlygate4sd3_1 hold915 (.A(_0617_),
    .X(net1831));
 sg13g2_dlygate4sd3_1 hold916 (.A(s_m_io4_out),
    .X(net1832));
 sg13g2_dlygate4sd3_1 hold917 (.A(_0254_),
    .X(net1833));
 sg13g2_dlygate4sd3_1 hold918 (.A(n351_q),
    .X(net1834));
 sg13g2_dlygate4sd3_1 hold919 (.A(\n353_q[10] ),
    .X(net1835));
 sg13g2_dlygate4sd3_1 hold920 (.A(_0123_),
    .X(net1836));
 sg13g2_dlygate4sd3_1 hold921 (.A(_0175_),
    .X(net1837));
 sg13g2_dlygate4sd3_1 hold922 (.A(_0089_),
    .X(net1838));
 sg13g2_dlygate4sd3_1 hold923 (.A(\usbfunction0.n2648_q[0] ),
    .X(net1839));
 sg13g2_dlygate4sd3_1 hold924 (.A(_0090_),
    .X(net1840));
 sg13g2_dlygate4sd3_1 hold925 (.A(\usbfunction0.n2653_q[0] ),
    .X(net1841));
 sg13g2_dlygate4sd3_1 hold926 (.A(\scl_uartrx0.n5991_o ),
    .X(net1842));
 sg13g2_dlygate4sd3_1 hold927 (.A(\usbfunction0.functionreset0.in_unnamed_3[3] ),
    .X(net1843));
 sg13g2_dlygate4sd3_1 hold928 (.A(\usbfunction0.n1083_o[3] ),
    .X(net1844));
 sg13g2_dlygate4sd3_1 hold929 (.A(\usbfunction0.functionreset0.in_unnamed_3[4] ),
    .X(net1845));
 sg13g2_dlygate4sd3_1 hold930 (.A(_0981_),
    .X(net1846));
 sg13g2_dlygate4sd3_1 hold931 (.A(\usbfunction0.n665_o[4] ),
    .X(net1847));
 sg13g2_dlygate4sd3_1 hold932 (.A(\scl_uarttx0.n2856_o[1] ),
    .X(net1848));
 sg13g2_dlygate4sd3_1 hold933 (.A(\scl_uarttx0.scl_counter0.n6919_o[1] ),
    .X(net1849));
 sg13g2_dlygate4sd3_1 hold934 (.A(_0101_),
    .X(net1850));
 sg13g2_dlygate4sd3_1 hold935 (.A(\scl_bitbangengine0.n3663_o[0] ),
    .X(net1851));
 sg13g2_dlygate4sd3_1 hold936 (.A(\n353_q[12] ),
    .X(net1852));
 sg13g2_dlygate4sd3_1 hold937 (.A(_0061_),
    .X(net1853));
 sg13g2_dlygate4sd3_1 hold938 (.A(\usbfunction0.n2313_o[3] ),
    .X(net1854));
 sg13g2_dlygate4sd3_1 hold939 (.A(_3253_),
    .X(net1855));
 sg13g2_dlygate4sd3_1 hold940 (.A(_0678_),
    .X(net1856));
 sg13g2_dlygate4sd3_1 hold941 (.A(\n353_q[23] ),
    .X(net1857));
 sg13g2_dlygate4sd3_1 hold942 (.A(_0125_),
    .X(net1858));
 sg13g2_dlygate4sd3_1 hold943 (.A(\n353_q[11] ),
    .X(net1859));
 sg13g2_dlygate4sd3_1 hold944 (.A(\n352_o[11] ),
    .X(net1860));
 sg13g2_dlygate4sd3_1 hold945 (.A(\scl_bitbangengine0.n3258_o ),
    .X(net1861));
 sg13g2_dlygate4sd3_1 hold946 (.A(_2700_),
    .X(net1862));
 sg13g2_dlygate4sd3_1 hold947 (.A(_0095_),
    .X(net1863));
 sg13g2_dlygate4sd3_1 hold948 (.A(\s_m_pushdata_data[2] ),
    .X(net1864));
 sg13g2_dlygate4sd3_1 hold949 (.A(_0088_),
    .X(net1865));
 sg13g2_dlygate4sd3_1 hold950 (.A(\scl_bitbangengine0.n3817_o ),
    .X(net1866));
 sg13g2_dlygate4sd3_1 hold951 (.A(\scl_bitbangengine0.n5920_q[8] ),
    .X(net1867));
 sg13g2_dlygate4sd3_1 hold952 (.A(\scl_bitbangengine0.scl_counter0.n6975_q[1] ),
    .X(net1868));
 sg13g2_dlygate4sd3_1 hold953 (.A(\n353_q[22] ),
    .X(net1869));
 sg13g2_dlygate4sd3_1 hold954 (.A(\usbfunction0.n2634_q[3] ),
    .X(net1870));
 sg13g2_dlygate4sd3_1 hold955 (.A(\n353_q[21] ),
    .X(net1871));
 sg13g2_dlygate4sd3_1 hold956 (.A(\s_m_pushdata_data[1] ),
    .X(net1872));
 sg13g2_dlygate4sd3_1 hold957 (.A(\usbfunction0.n2651_q[6] ),
    .X(net1873));
 sg13g2_dlygate4sd3_1 hold958 (.A(\usbfunction0.n2642_q[0] ),
    .X(net1874));
 sg13g2_dlygate4sd3_1 hold959 (.A(\s_m_pushdata_data[0] ),
    .X(net1875));
 sg13g2_dlygate4sd3_1 hold960 (.A(\usbfunction0.functionreset0.in_unnamed[2] ),
    .X(net1876));
 sg13g2_dlygate4sd3_1 hold961 (.A(s_m_io3_out),
    .X(net1877));
 sg13g2_dlygate4sd3_1 hold962 (.A(\usbfunction0.scl_usbgpiophy0.scl_insertbeat0.n7369_o ),
    .X(net1878));
 sg13g2_dlygate4sd3_1 hold963 (.A(\usbfunction0.scl_usbgpiophy0.scl_addeopdeferred0.n7339_o ),
    .X(net1879));
 sg13g2_dlygate4sd3_1 hold964 (.A(s_m_packetdata_2_bit_17),
    .X(net1880));
 sg13g2_dlygate4sd3_1 hold965 (.A(\usbfunction0.n2652_q[7] ),
    .X(net1881));
 sg13g2_dlygate4sd3_1 hold966 (.A(_0096_),
    .X(net1882));
 sg13g2_dlygate4sd3_1 hold967 (.A(\usbfunction0.functionreset0.in_unnamed[3] ),
    .X(net1883));
 sg13g2_dlygate4sd3_1 hold968 (.A(\usbfunction0.n665_o[3] ),
    .X(net1884));
 sg13g2_dlygate4sd3_1 hold969 (.A(\usbfunction0.functionreset0.in_unnamed[0] ),
    .X(net1885));
 sg13g2_dlygate4sd3_1 hold970 (.A(\usbfunction0.functionreset0.in_unnamed[5] ),
    .X(net1886));
 sg13g2_dlygate4sd3_1 hold971 (.A(\usbfunction0.n665_o[5] ),
    .X(net1887));
 sg13g2_dlygate4sd3_1 hold972 (.A(\usbfunction0.n2634_q[1] ),
    .X(net1888));
 sg13g2_dlygate4sd3_1 hold973 (.A(\scl_bitbangengine0.n5920_q[0] ),
    .X(net1889));
 sg13g2_dlygate4sd3_1 hold974 (.A(s_m_io1_out),
    .X(net1890));
 sg13g2_dlygate4sd3_1 hold975 (.A(_2801_),
    .X(net1891));
 sg13g2_dlygate4sd3_1 hold976 (.A(\scl_bitbangengine0.n5898_q[0] ),
    .X(net1892));
 sg13g2_dlygate4sd3_1 hold977 (.A(_0210_),
    .X(net1893));
 sg13g2_dlygate4sd3_1 hold978 (.A(\usbfunction0.n2651_q[5] ),
    .X(net1894));
 sg13g2_dlygate4sd3_1 hold979 (.A(\scl_fifo1.scl_memory0.physical_memory0.memory[12][1] ),
    .X(net1895));
 sg13g2_dlygate4sd3_1 hold980 (.A(_0101_),
    .X(net1896));
 sg13g2_dlygate4sd3_1 hold981 (.A(\usbfunction0.n2650_q[0] ),
    .X(net1897));
 sg13g2_dlygate4sd3_1 hold982 (.A(\scl_bitbangengine0.n5898_q[1] ),
    .X(net1898));
 sg13g2_dlygate4sd3_1 hold983 (.A(\usbfunction0.n2651_q[4] ),
    .X(net1899));
 sg13g2_dlygate4sd3_1 hold984 (.A(_0098_),
    .X(net1900));
 sg13g2_dlygate4sd3_1 hold985 (.A(\scl_uarttx0.scl_baudrategenerator0.n6874_o[3] ),
    .X(net1901));
 sg13g2_dlygate4sd3_1 hold986 (.A(\usbfunction0.n1359_o[0] ),
    .X(net1902));
 sg13g2_dlygate4sd3_1 hold987 (.A(\scl_bitbangengine0.n3817_o ),
    .X(net1903));
 sg13g2_dlygate4sd3_1 hold988 (.A(s_m_packetdata_2_bit_16),
    .X(net1904));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_4 FILLER_2_350 ();
 sg13g2_fill_1 FILLER_2_354 ();
 sg13g2_fill_1 FILLER_2_359 ();
 sg13g2_fill_2 FILLER_2_364 ();
 sg13g2_fill_1 FILLER_2_370 ();
 sg13g2_decap_8 FILLER_2_397 ();
 sg13g2_decap_8 FILLER_2_404 ();
 sg13g2_decap_8 FILLER_2_411 ();
 sg13g2_decap_8 FILLER_2_418 ();
 sg13g2_decap_8 FILLER_2_425 ();
 sg13g2_decap_8 FILLER_2_432 ();
 sg13g2_decap_8 FILLER_2_439 ();
 sg13g2_decap_8 FILLER_2_446 ();
 sg13g2_decap_8 FILLER_2_453 ();
 sg13g2_decap_4 FILLER_2_460 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_fill_1 FILLER_2_497 ();
 sg13g2_fill_2 FILLER_2_502 ();
 sg13g2_fill_1 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_531 ();
 sg13g2_decap_8 FILLER_2_538 ();
 sg13g2_decap_8 FILLER_2_545 ();
 sg13g2_decap_8 FILLER_2_552 ();
 sg13g2_decap_8 FILLER_2_559 ();
 sg13g2_decap_8 FILLER_2_566 ();
 sg13g2_decap_8 FILLER_2_573 ();
 sg13g2_decap_8 FILLER_2_580 ();
 sg13g2_decap_8 FILLER_2_587 ();
 sg13g2_decap_8 FILLER_2_594 ();
 sg13g2_decap_8 FILLER_2_601 ();
 sg13g2_decap_8 FILLER_2_608 ();
 sg13g2_decap_8 FILLER_2_615 ();
 sg13g2_decap_8 FILLER_2_622 ();
 sg13g2_decap_8 FILLER_2_629 ();
 sg13g2_decap_8 FILLER_2_636 ();
 sg13g2_decap_8 FILLER_2_643 ();
 sg13g2_decap_8 FILLER_2_650 ();
 sg13g2_decap_8 FILLER_2_657 ();
 sg13g2_decap_8 FILLER_2_664 ();
 sg13g2_decap_8 FILLER_2_671 ();
 sg13g2_decap_8 FILLER_2_678 ();
 sg13g2_decap_8 FILLER_2_685 ();
 sg13g2_decap_8 FILLER_2_692 ();
 sg13g2_decap_8 FILLER_2_699 ();
 sg13g2_decap_8 FILLER_2_706 ();
 sg13g2_decap_8 FILLER_2_713 ();
 sg13g2_decap_8 FILLER_2_720 ();
 sg13g2_decap_8 FILLER_2_727 ();
 sg13g2_decap_8 FILLER_2_734 ();
 sg13g2_decap_8 FILLER_2_741 ();
 sg13g2_decap_8 FILLER_2_748 ();
 sg13g2_decap_8 FILLER_2_755 ();
 sg13g2_decap_8 FILLER_2_762 ();
 sg13g2_decap_8 FILLER_2_769 ();
 sg13g2_decap_8 FILLER_2_776 ();
 sg13g2_decap_8 FILLER_2_783 ();
 sg13g2_decap_8 FILLER_2_790 ();
 sg13g2_decap_8 FILLER_2_797 ();
 sg13g2_decap_8 FILLER_2_804 ();
 sg13g2_decap_8 FILLER_2_811 ();
 sg13g2_decap_8 FILLER_2_818 ();
 sg13g2_decap_8 FILLER_2_825 ();
 sg13g2_decap_8 FILLER_2_832 ();
 sg13g2_decap_8 FILLER_2_839 ();
 sg13g2_decap_8 FILLER_2_846 ();
 sg13g2_decap_8 FILLER_2_853 ();
 sg13g2_fill_2 FILLER_2_860 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_4 FILLER_3_315 ();
 sg13g2_decap_4 FILLER_3_384 ();
 sg13g2_fill_2 FILLER_3_414 ();
 sg13g2_decap_4 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_424 ();
 sg13g2_decap_8 FILLER_3_452 ();
 sg13g2_fill_1 FILLER_3_459 ();
 sg13g2_fill_2 FILLER_3_490 ();
 sg13g2_fill_1 FILLER_3_492 ();
 sg13g2_decap_8 FILLER_3_527 ();
 sg13g2_decap_8 FILLER_3_534 ();
 sg13g2_decap_8 FILLER_3_541 ();
 sg13g2_fill_1 FILLER_3_548 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_327 ();
 sg13g2_decap_4 FILLER_4_338 ();
 sg13g2_fill_1 FILLER_4_352 ();
 sg13g2_fill_2 FILLER_4_362 ();
 sg13g2_fill_1 FILLER_4_372 ();
 sg13g2_fill_2 FILLER_4_403 ();
 sg13g2_fill_2 FILLER_4_479 ();
 sg13g2_fill_1 FILLER_4_481 ();
 sg13g2_fill_2 FILLER_4_500 ();
 sg13g2_fill_2 FILLER_4_521 ();
 sg13g2_decap_4 FILLER_4_532 ();
 sg13g2_fill_2 FILLER_4_536 ();
 sg13g2_decap_8 FILLER_4_573 ();
 sg13g2_decap_8 FILLER_4_580 ();
 sg13g2_decap_8 FILLER_4_587 ();
 sg13g2_decap_8 FILLER_4_594 ();
 sg13g2_decap_8 FILLER_4_601 ();
 sg13g2_decap_8 FILLER_4_608 ();
 sg13g2_decap_8 FILLER_4_615 ();
 sg13g2_decap_8 FILLER_4_622 ();
 sg13g2_decap_8 FILLER_4_629 ();
 sg13g2_decap_8 FILLER_4_636 ();
 sg13g2_decap_8 FILLER_4_643 ();
 sg13g2_decap_8 FILLER_4_650 ();
 sg13g2_decap_8 FILLER_4_657 ();
 sg13g2_decap_8 FILLER_4_664 ();
 sg13g2_decap_8 FILLER_4_671 ();
 sg13g2_decap_8 FILLER_4_678 ();
 sg13g2_decap_8 FILLER_4_685 ();
 sg13g2_decap_8 FILLER_4_692 ();
 sg13g2_decap_8 FILLER_4_699 ();
 sg13g2_decap_8 FILLER_4_706 ();
 sg13g2_decap_8 FILLER_4_713 ();
 sg13g2_decap_8 FILLER_4_720 ();
 sg13g2_decap_8 FILLER_4_727 ();
 sg13g2_decap_8 FILLER_4_734 ();
 sg13g2_decap_8 FILLER_4_741 ();
 sg13g2_decap_8 FILLER_4_748 ();
 sg13g2_decap_8 FILLER_4_755 ();
 sg13g2_decap_8 FILLER_4_762 ();
 sg13g2_decap_8 FILLER_4_769 ();
 sg13g2_decap_8 FILLER_4_776 ();
 sg13g2_decap_8 FILLER_4_783 ();
 sg13g2_decap_8 FILLER_4_790 ();
 sg13g2_decap_8 FILLER_4_797 ();
 sg13g2_decap_8 FILLER_4_804 ();
 sg13g2_decap_8 FILLER_4_811 ();
 sg13g2_decap_8 FILLER_4_818 ();
 sg13g2_decap_8 FILLER_4_825 ();
 sg13g2_decap_8 FILLER_4_832 ();
 sg13g2_decap_8 FILLER_4_839 ();
 sg13g2_decap_8 FILLER_4_846 ();
 sg13g2_decap_8 FILLER_4_853 ();
 sg13g2_fill_2 FILLER_4_860 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_fill_1 FILLER_5_359 ();
 sg13g2_fill_1 FILLER_5_380 ();
 sg13g2_fill_2 FILLER_5_394 ();
 sg13g2_decap_4 FILLER_5_413 ();
 sg13g2_fill_2 FILLER_5_460 ();
 sg13g2_fill_1 FILLER_5_462 ();
 sg13g2_fill_2 FILLER_5_469 ();
 sg13g2_fill_1 FILLER_5_471 ();
 sg13g2_fill_2 FILLER_5_541 ();
 sg13g2_fill_1 FILLER_5_543 ();
 sg13g2_decap_8 FILLER_5_583 ();
 sg13g2_decap_8 FILLER_5_590 ();
 sg13g2_decap_8 FILLER_5_597 ();
 sg13g2_decap_8 FILLER_5_604 ();
 sg13g2_decap_8 FILLER_5_611 ();
 sg13g2_decap_8 FILLER_5_618 ();
 sg13g2_decap_8 FILLER_5_625 ();
 sg13g2_decap_8 FILLER_5_632 ();
 sg13g2_decap_8 FILLER_5_639 ();
 sg13g2_decap_8 FILLER_5_646 ();
 sg13g2_decap_8 FILLER_5_653 ();
 sg13g2_decap_8 FILLER_5_660 ();
 sg13g2_decap_8 FILLER_5_667 ();
 sg13g2_decap_8 FILLER_5_674 ();
 sg13g2_decap_8 FILLER_5_681 ();
 sg13g2_decap_8 FILLER_5_688 ();
 sg13g2_decap_8 FILLER_5_695 ();
 sg13g2_decap_8 FILLER_5_702 ();
 sg13g2_decap_8 FILLER_5_709 ();
 sg13g2_decap_8 FILLER_5_716 ();
 sg13g2_decap_8 FILLER_5_723 ();
 sg13g2_decap_8 FILLER_5_730 ();
 sg13g2_decap_8 FILLER_5_737 ();
 sg13g2_decap_8 FILLER_5_744 ();
 sg13g2_decap_8 FILLER_5_751 ();
 sg13g2_decap_8 FILLER_5_758 ();
 sg13g2_decap_8 FILLER_5_765 ();
 sg13g2_decap_8 FILLER_5_772 ();
 sg13g2_decap_8 FILLER_5_779 ();
 sg13g2_decap_8 FILLER_5_786 ();
 sg13g2_decap_8 FILLER_5_793 ();
 sg13g2_decap_8 FILLER_5_800 ();
 sg13g2_decap_8 FILLER_5_807 ();
 sg13g2_decap_8 FILLER_5_814 ();
 sg13g2_decap_8 FILLER_5_821 ();
 sg13g2_decap_8 FILLER_5_828 ();
 sg13g2_decap_8 FILLER_5_835 ();
 sg13g2_decap_8 FILLER_5_842 ();
 sg13g2_decap_8 FILLER_5_849 ();
 sg13g2_decap_4 FILLER_5_856 ();
 sg13g2_fill_2 FILLER_5_860 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_fill_2 FILLER_6_301 ();
 sg13g2_fill_1 FILLER_6_303 ();
 sg13g2_fill_2 FILLER_6_313 ();
 sg13g2_decap_8 FILLER_6_330 ();
 sg13g2_decap_8 FILLER_6_337 ();
 sg13g2_fill_1 FILLER_6_344 ();
 sg13g2_fill_2 FILLER_6_361 ();
 sg13g2_fill_2 FILLER_6_398 ();
 sg13g2_fill_2 FILLER_6_414 ();
 sg13g2_fill_1 FILLER_6_416 ();
 sg13g2_decap_4 FILLER_6_431 ();
 sg13g2_fill_2 FILLER_6_435 ();
 sg13g2_fill_2 FILLER_6_460 ();
 sg13g2_fill_1 FILLER_6_462 ();
 sg13g2_decap_4 FILLER_6_467 ();
 sg13g2_fill_1 FILLER_6_471 ();
 sg13g2_decap_4 FILLER_6_476 ();
 sg13g2_decap_4 FILLER_6_484 ();
 sg13g2_fill_2 FILLER_6_488 ();
 sg13g2_decap_4 FILLER_6_495 ();
 sg13g2_fill_2 FILLER_6_499 ();
 sg13g2_fill_1 FILLER_6_508 ();
 sg13g2_decap_4 FILLER_6_522 ();
 sg13g2_decap_4 FILLER_6_530 ();
 sg13g2_fill_2 FILLER_6_564 ();
 sg13g2_fill_1 FILLER_6_566 ();
 sg13g2_decap_8 FILLER_6_593 ();
 sg13g2_decap_8 FILLER_6_600 ();
 sg13g2_decap_8 FILLER_6_607 ();
 sg13g2_decap_8 FILLER_6_614 ();
 sg13g2_decap_8 FILLER_6_621 ();
 sg13g2_decap_8 FILLER_6_628 ();
 sg13g2_decap_8 FILLER_6_635 ();
 sg13g2_decap_8 FILLER_6_642 ();
 sg13g2_decap_8 FILLER_6_649 ();
 sg13g2_decap_8 FILLER_6_656 ();
 sg13g2_decap_8 FILLER_6_663 ();
 sg13g2_decap_8 FILLER_6_670 ();
 sg13g2_decap_8 FILLER_6_677 ();
 sg13g2_decap_8 FILLER_6_684 ();
 sg13g2_decap_8 FILLER_6_691 ();
 sg13g2_decap_8 FILLER_6_698 ();
 sg13g2_decap_8 FILLER_6_705 ();
 sg13g2_decap_8 FILLER_6_712 ();
 sg13g2_decap_8 FILLER_6_719 ();
 sg13g2_decap_8 FILLER_6_726 ();
 sg13g2_decap_8 FILLER_6_733 ();
 sg13g2_decap_8 FILLER_6_740 ();
 sg13g2_decap_8 FILLER_6_747 ();
 sg13g2_decap_8 FILLER_6_754 ();
 sg13g2_decap_8 FILLER_6_761 ();
 sg13g2_decap_8 FILLER_6_768 ();
 sg13g2_decap_8 FILLER_6_775 ();
 sg13g2_decap_8 FILLER_6_782 ();
 sg13g2_decap_8 FILLER_6_789 ();
 sg13g2_decap_8 FILLER_6_796 ();
 sg13g2_decap_8 FILLER_6_803 ();
 sg13g2_decap_8 FILLER_6_810 ();
 sg13g2_decap_8 FILLER_6_817 ();
 sg13g2_decap_8 FILLER_6_824 ();
 sg13g2_decap_8 FILLER_6_831 ();
 sg13g2_decap_8 FILLER_6_838 ();
 sg13g2_decap_8 FILLER_6_845 ();
 sg13g2_decap_8 FILLER_6_852 ();
 sg13g2_fill_2 FILLER_6_859 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_fill_1 FILLER_7_334 ();
 sg13g2_fill_2 FILLER_7_361 ();
 sg13g2_decap_8 FILLER_7_409 ();
 sg13g2_decap_4 FILLER_7_416 ();
 sg13g2_fill_1 FILLER_7_420 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_fill_2 FILLER_7_435 ();
 sg13g2_fill_2 FILLER_7_471 ();
 sg13g2_fill_2 FILLER_7_495 ();
 sg13g2_fill_1 FILLER_7_505 ();
 sg13g2_fill_2 FILLER_7_540 ();
 sg13g2_fill_1 FILLER_7_542 ();
 sg13g2_fill_1 FILLER_7_556 ();
 sg13g2_decap_8 FILLER_7_601 ();
 sg13g2_decap_8 FILLER_7_608 ();
 sg13g2_decap_8 FILLER_7_615 ();
 sg13g2_decap_4 FILLER_7_622 ();
 sg13g2_fill_2 FILLER_7_626 ();
 sg13g2_decap_8 FILLER_7_632 ();
 sg13g2_decap_8 FILLER_7_639 ();
 sg13g2_decap_8 FILLER_7_646 ();
 sg13g2_decap_8 FILLER_7_653 ();
 sg13g2_decap_8 FILLER_7_660 ();
 sg13g2_decap_8 FILLER_7_667 ();
 sg13g2_decap_8 FILLER_7_674 ();
 sg13g2_decap_8 FILLER_7_681 ();
 sg13g2_decap_8 FILLER_7_688 ();
 sg13g2_decap_8 FILLER_7_695 ();
 sg13g2_decap_8 FILLER_7_702 ();
 sg13g2_decap_8 FILLER_7_709 ();
 sg13g2_decap_8 FILLER_7_716 ();
 sg13g2_decap_8 FILLER_7_723 ();
 sg13g2_decap_8 FILLER_7_730 ();
 sg13g2_decap_8 FILLER_7_737 ();
 sg13g2_decap_8 FILLER_7_744 ();
 sg13g2_decap_8 FILLER_7_751 ();
 sg13g2_decap_8 FILLER_7_758 ();
 sg13g2_decap_8 FILLER_7_765 ();
 sg13g2_decap_8 FILLER_7_772 ();
 sg13g2_decap_8 FILLER_7_779 ();
 sg13g2_decap_8 FILLER_7_786 ();
 sg13g2_decap_8 FILLER_7_793 ();
 sg13g2_decap_8 FILLER_7_800 ();
 sg13g2_decap_8 FILLER_7_807 ();
 sg13g2_decap_8 FILLER_7_814 ();
 sg13g2_decap_8 FILLER_7_821 ();
 sg13g2_decap_8 FILLER_7_828 ();
 sg13g2_decap_8 FILLER_7_835 ();
 sg13g2_decap_8 FILLER_7_842 ();
 sg13g2_decap_8 FILLER_7_849 ();
 sg13g2_decap_4 FILLER_7_856 ();
 sg13g2_fill_2 FILLER_7_860 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_4 FILLER_8_112 ();
 sg13g2_fill_2 FILLER_8_116 ();
 sg13g2_decap_8 FILLER_8_127 ();
 sg13g2_decap_8 FILLER_8_134 ();
 sg13g2_decap_8 FILLER_8_141 ();
 sg13g2_decap_8 FILLER_8_148 ();
 sg13g2_decap_8 FILLER_8_155 ();
 sg13g2_decap_8 FILLER_8_162 ();
 sg13g2_decap_8 FILLER_8_169 ();
 sg13g2_decap_8 FILLER_8_176 ();
 sg13g2_decap_8 FILLER_8_183 ();
 sg13g2_decap_8 FILLER_8_190 ();
 sg13g2_decap_8 FILLER_8_197 ();
 sg13g2_decap_8 FILLER_8_204 ();
 sg13g2_decap_8 FILLER_8_211 ();
 sg13g2_decap_8 FILLER_8_218 ();
 sg13g2_decap_8 FILLER_8_225 ();
 sg13g2_decap_8 FILLER_8_232 ();
 sg13g2_decap_8 FILLER_8_239 ();
 sg13g2_decap_8 FILLER_8_246 ();
 sg13g2_decap_8 FILLER_8_253 ();
 sg13g2_decap_8 FILLER_8_260 ();
 sg13g2_decap_8 FILLER_8_267 ();
 sg13g2_decap_8 FILLER_8_274 ();
 sg13g2_fill_1 FILLER_8_281 ();
 sg13g2_fill_2 FILLER_8_308 ();
 sg13g2_fill_1 FILLER_8_331 ();
 sg13g2_fill_1 FILLER_8_444 ();
 sg13g2_fill_2 FILLER_8_454 ();
 sg13g2_fill_1 FILLER_8_456 ();
 sg13g2_fill_2 FILLER_8_474 ();
 sg13g2_fill_1 FILLER_8_476 ();
 sg13g2_fill_1 FILLER_8_493 ();
 sg13g2_fill_1 FILLER_8_498 ();
 sg13g2_fill_2 FILLER_8_511 ();
 sg13g2_fill_1 FILLER_8_513 ();
 sg13g2_fill_1 FILLER_8_535 ();
 sg13g2_fill_2 FILLER_8_551 ();
 sg13g2_decap_8 FILLER_8_612 ();
 sg13g2_fill_2 FILLER_8_646 ();
 sg13g2_fill_2 FILLER_8_662 ();
 sg13g2_decap_8 FILLER_8_681 ();
 sg13g2_decap_8 FILLER_8_688 ();
 sg13g2_decap_4 FILLER_8_695 ();
 sg13g2_fill_1 FILLER_8_699 ();
 sg13g2_decap_8 FILLER_8_704 ();
 sg13g2_decap_8 FILLER_8_711 ();
 sg13g2_decap_8 FILLER_8_718 ();
 sg13g2_decap_8 FILLER_8_725 ();
 sg13g2_decap_8 FILLER_8_732 ();
 sg13g2_decap_8 FILLER_8_739 ();
 sg13g2_decap_8 FILLER_8_746 ();
 sg13g2_decap_8 FILLER_8_753 ();
 sg13g2_decap_8 FILLER_8_760 ();
 sg13g2_decap_8 FILLER_8_767 ();
 sg13g2_decap_8 FILLER_8_774 ();
 sg13g2_decap_8 FILLER_8_781 ();
 sg13g2_decap_8 FILLER_8_788 ();
 sg13g2_decap_8 FILLER_8_795 ();
 sg13g2_decap_8 FILLER_8_802 ();
 sg13g2_decap_8 FILLER_8_809 ();
 sg13g2_decap_8 FILLER_8_816 ();
 sg13g2_decap_8 FILLER_8_823 ();
 sg13g2_decap_8 FILLER_8_830 ();
 sg13g2_decap_8 FILLER_8_837 ();
 sg13g2_decap_8 FILLER_8_844 ();
 sg13g2_decap_8 FILLER_8_851 ();
 sg13g2_decap_4 FILLER_8_858 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_fill_2 FILLER_9_56 ();
 sg13g2_fill_1 FILLER_9_58 ();
 sg13g2_decap_8 FILLER_9_64 ();
 sg13g2_fill_1 FILLER_9_71 ();
 sg13g2_decap_8 FILLER_9_81 ();
 sg13g2_decap_8 FILLER_9_88 ();
 sg13g2_decap_8 FILLER_9_95 ();
 sg13g2_decap_4 FILLER_9_102 ();
 sg13g2_fill_2 FILLER_9_132 ();
 sg13g2_decap_4 FILLER_9_143 ();
 sg13g2_decap_8 FILLER_9_151 ();
 sg13g2_decap_4 FILLER_9_158 ();
 sg13g2_fill_1 FILLER_9_162 ();
 sg13g2_fill_1 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_263 ();
 sg13g2_decap_8 FILLER_9_270 ();
 sg13g2_decap_8 FILLER_9_277 ();
 sg13g2_decap_8 FILLER_9_284 ();
 sg13g2_decap_8 FILLER_9_291 ();
 sg13g2_fill_1 FILLER_9_298 ();
 sg13g2_fill_2 FILLER_9_308 ();
 sg13g2_fill_1 FILLER_9_310 ();
 sg13g2_fill_1 FILLER_9_331 ();
 sg13g2_fill_2 FILLER_9_414 ();
 sg13g2_fill_1 FILLER_9_416 ();
 sg13g2_fill_1 FILLER_9_450 ();
 sg13g2_fill_1 FILLER_9_469 ();
 sg13g2_decap_4 FILLER_9_474 ();
 sg13g2_fill_2 FILLER_9_478 ();
 sg13g2_fill_2 FILLER_9_495 ();
 sg13g2_fill_2 FILLER_9_504 ();
 sg13g2_fill_1 FILLER_9_506 ();
 sg13g2_fill_1 FILLER_9_512 ();
 sg13g2_fill_2 FILLER_9_539 ();
 sg13g2_fill_2 FILLER_9_561 ();
 sg13g2_fill_1 FILLER_9_563 ();
 sg13g2_fill_1 FILLER_9_590 ();
 sg13g2_fill_2 FILLER_9_601 ();
 sg13g2_fill_1 FILLER_9_616 ();
 sg13g2_fill_1 FILLER_9_653 ();
 sg13g2_fill_1 FILLER_9_680 ();
 sg13g2_fill_2 FILLER_9_695 ();
 sg13g2_fill_1 FILLER_9_697 ();
 sg13g2_decap_8 FILLER_9_724 ();
 sg13g2_decap_8 FILLER_9_731 ();
 sg13g2_decap_8 FILLER_9_738 ();
 sg13g2_decap_8 FILLER_9_745 ();
 sg13g2_decap_8 FILLER_9_752 ();
 sg13g2_decap_8 FILLER_9_759 ();
 sg13g2_decap_8 FILLER_9_766 ();
 sg13g2_decap_8 FILLER_9_773 ();
 sg13g2_decap_8 FILLER_9_780 ();
 sg13g2_decap_8 FILLER_9_787 ();
 sg13g2_decap_8 FILLER_9_794 ();
 sg13g2_decap_8 FILLER_9_801 ();
 sg13g2_decap_8 FILLER_9_808 ();
 sg13g2_decap_8 FILLER_9_815 ();
 sg13g2_decap_8 FILLER_9_822 ();
 sg13g2_decap_8 FILLER_9_829 ();
 sg13g2_decap_8 FILLER_9_836 ();
 sg13g2_decap_8 FILLER_9_843 ();
 sg13g2_decap_8 FILLER_9_850 ();
 sg13g2_decap_4 FILLER_9_857 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_4 FILLER_10_42 ();
 sg13g2_fill_2 FILLER_10_46 ();
 sg13g2_fill_1 FILLER_10_88 ();
 sg13g2_fill_2 FILLER_10_99 ();
 sg13g2_fill_1 FILLER_10_111 ();
 sg13g2_decap_8 FILLER_10_162 ();
 sg13g2_fill_1 FILLER_10_169 ();
 sg13g2_decap_4 FILLER_10_206 ();
 sg13g2_decap_8 FILLER_10_236 ();
 sg13g2_decap_4 FILLER_10_243 ();
 sg13g2_fill_1 FILLER_10_247 ();
 sg13g2_decap_8 FILLER_10_283 ();
 sg13g2_fill_1 FILLER_10_290 ();
 sg13g2_fill_2 FILLER_10_377 ();
 sg13g2_fill_1 FILLER_10_400 ();
 sg13g2_decap_4 FILLER_10_410 ();
 sg13g2_fill_1 FILLER_10_414 ();
 sg13g2_fill_2 FILLER_10_499 ();
 sg13g2_fill_1 FILLER_10_501 ();
 sg13g2_fill_2 FILLER_10_532 ();
 sg13g2_fill_1 FILLER_10_534 ();
 sg13g2_fill_2 FILLER_10_554 ();
 sg13g2_fill_2 FILLER_10_590 ();
 sg13g2_fill_1 FILLER_10_592 ();
 sg13g2_decap_8 FILLER_10_734 ();
 sg13g2_decap_8 FILLER_10_741 ();
 sg13g2_decap_8 FILLER_10_748 ();
 sg13g2_decap_8 FILLER_10_755 ();
 sg13g2_decap_8 FILLER_10_762 ();
 sg13g2_decap_8 FILLER_10_769 ();
 sg13g2_decap_8 FILLER_10_776 ();
 sg13g2_decap_8 FILLER_10_783 ();
 sg13g2_decap_8 FILLER_10_790 ();
 sg13g2_decap_8 FILLER_10_797 ();
 sg13g2_decap_8 FILLER_10_804 ();
 sg13g2_decap_8 FILLER_10_811 ();
 sg13g2_decap_8 FILLER_10_818 ();
 sg13g2_decap_8 FILLER_10_825 ();
 sg13g2_decap_8 FILLER_10_832 ();
 sg13g2_decap_8 FILLER_10_839 ();
 sg13g2_decap_8 FILLER_10_846 ();
 sg13g2_decap_8 FILLER_10_853 ();
 sg13g2_fill_2 FILLER_10_860 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_4 FILLER_11_7 ();
 sg13g2_fill_1 FILLER_11_11 ();
 sg13g2_fill_1 FILLER_11_88 ();
 sg13g2_fill_1 FILLER_11_115 ();
 sg13g2_decap_4 FILLER_11_142 ();
 sg13g2_fill_2 FILLER_11_146 ();
 sg13g2_fill_2 FILLER_11_156 ();
 sg13g2_fill_1 FILLER_11_168 ();
 sg13g2_decap_4 FILLER_11_182 ();
 sg13g2_fill_2 FILLER_11_229 ();
 sg13g2_fill_1 FILLER_11_231 ();
 sg13g2_fill_2 FILLER_11_251 ();
 sg13g2_fill_1 FILLER_11_253 ();
 sg13g2_fill_1 FILLER_11_315 ();
 sg13g2_fill_2 FILLER_11_325 ();
 sg13g2_fill_2 FILLER_11_346 ();
 sg13g2_fill_1 FILLER_11_348 ();
 sg13g2_fill_1 FILLER_11_353 ();
 sg13g2_fill_2 FILLER_11_373 ();
 sg13g2_fill_1 FILLER_11_379 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_440 ();
 sg13g2_decap_8 FILLER_11_447 ();
 sg13g2_decap_8 FILLER_11_454 ();
 sg13g2_fill_2 FILLER_11_461 ();
 sg13g2_fill_1 FILLER_11_463 ();
 sg13g2_fill_2 FILLER_11_480 ();
 sg13g2_fill_1 FILLER_11_482 ();
 sg13g2_decap_4 FILLER_11_491 ();
 sg13g2_fill_1 FILLER_11_500 ();
 sg13g2_fill_1 FILLER_11_505 ();
 sg13g2_fill_2 FILLER_11_533 ();
 sg13g2_decap_4 FILLER_11_543 ();
 sg13g2_decap_8 FILLER_11_565 ();
 sg13g2_fill_1 FILLER_11_572 ();
 sg13g2_fill_2 FILLER_11_589 ();
 sg13g2_fill_1 FILLER_11_591 ();
 sg13g2_fill_2 FILLER_11_642 ();
 sg13g2_fill_1 FILLER_11_680 ();
 sg13g2_fill_1 FILLER_11_708 ();
 sg13g2_decap_8 FILLER_11_745 ();
 sg13g2_decap_8 FILLER_11_752 ();
 sg13g2_decap_8 FILLER_11_759 ();
 sg13g2_decap_8 FILLER_11_766 ();
 sg13g2_decap_8 FILLER_11_773 ();
 sg13g2_decap_8 FILLER_11_780 ();
 sg13g2_decap_8 FILLER_11_787 ();
 sg13g2_decap_8 FILLER_11_794 ();
 sg13g2_decap_8 FILLER_11_801 ();
 sg13g2_decap_8 FILLER_11_808 ();
 sg13g2_decap_8 FILLER_11_815 ();
 sg13g2_decap_8 FILLER_11_822 ();
 sg13g2_decap_8 FILLER_11_829 ();
 sg13g2_decap_8 FILLER_11_836 ();
 sg13g2_decap_8 FILLER_11_843 ();
 sg13g2_decap_8 FILLER_11_850 ();
 sg13g2_decap_4 FILLER_11_857 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_4 FILLER_12_7 ();
 sg13g2_fill_1 FILLER_12_11 ();
 sg13g2_fill_2 FILLER_12_45 ();
 sg13g2_fill_2 FILLER_12_57 ();
 sg13g2_fill_2 FILLER_12_141 ();
 sg13g2_fill_1 FILLER_12_143 ();
 sg13g2_fill_1 FILLER_12_148 ();
 sg13g2_fill_1 FILLER_12_270 ();
 sg13g2_fill_2 FILLER_12_289 ();
 sg13g2_fill_1 FILLER_12_291 ();
 sg13g2_fill_1 FILLER_12_305 ();
 sg13g2_fill_1 FILLER_12_330 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_407 ();
 sg13g2_fill_2 FILLER_12_440 ();
 sg13g2_fill_1 FILLER_12_442 ();
 sg13g2_fill_2 FILLER_12_487 ();
 sg13g2_fill_1 FILLER_12_489 ();
 sg13g2_fill_2 FILLER_12_550 ();
 sg13g2_fill_1 FILLER_12_552 ();
 sg13g2_decap_4 FILLER_12_562 ();
 sg13g2_fill_1 FILLER_12_566 ();
 sg13g2_fill_2 FILLER_12_598 ();
 sg13g2_fill_1 FILLER_12_600 ();
 sg13g2_fill_1 FILLER_12_640 ();
 sg13g2_fill_1 FILLER_12_660 ();
 sg13g2_fill_1 FILLER_12_671 ();
 sg13g2_decap_8 FILLER_12_755 ();
 sg13g2_decap_8 FILLER_12_762 ();
 sg13g2_decap_8 FILLER_12_769 ();
 sg13g2_decap_8 FILLER_12_776 ();
 sg13g2_decap_8 FILLER_12_783 ();
 sg13g2_decap_8 FILLER_12_790 ();
 sg13g2_decap_8 FILLER_12_797 ();
 sg13g2_decap_8 FILLER_12_804 ();
 sg13g2_decap_8 FILLER_12_811 ();
 sg13g2_decap_8 FILLER_12_818 ();
 sg13g2_decap_8 FILLER_12_825 ();
 sg13g2_decap_8 FILLER_12_832 ();
 sg13g2_decap_8 FILLER_12_839 ();
 sg13g2_decap_8 FILLER_12_846 ();
 sg13g2_decap_8 FILLER_12_853 ();
 sg13g2_fill_2 FILLER_12_860 ();
 sg13g2_decap_4 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_4 ();
 sg13g2_fill_1 FILLER_13_32 ();
 sg13g2_fill_2 FILLER_13_43 ();
 sg13g2_fill_1 FILLER_13_59 ();
 sg13g2_fill_1 FILLER_13_86 ();
 sg13g2_fill_1 FILLER_13_110 ();
 sg13g2_decap_8 FILLER_13_173 ();
 sg13g2_fill_1 FILLER_13_193 ();
 sg13g2_fill_1 FILLER_13_198 ();
 sg13g2_fill_2 FILLER_13_212 ();
 sg13g2_fill_1 FILLER_13_214 ();
 sg13g2_decap_4 FILLER_13_219 ();
 sg13g2_fill_1 FILLER_13_292 ();
 sg13g2_fill_1 FILLER_13_333 ();
 sg13g2_decap_4 FILLER_13_346 ();
 sg13g2_fill_2 FILLER_13_350 ();
 sg13g2_fill_1 FILLER_13_359 ();
 sg13g2_fill_1 FILLER_13_365 ();
 sg13g2_fill_2 FILLER_13_382 ();
 sg13g2_fill_1 FILLER_13_388 ();
 sg13g2_fill_1 FILLER_13_436 ();
 sg13g2_fill_1 FILLER_13_474 ();
 sg13g2_fill_1 FILLER_13_493 ();
 sg13g2_fill_1 FILLER_13_507 ();
 sg13g2_fill_1 FILLER_13_512 ();
 sg13g2_fill_1 FILLER_13_526 ();
 sg13g2_fill_1 FILLER_13_540 ();
 sg13g2_decap_4 FILLER_13_549 ();
 sg13g2_fill_1 FILLER_13_579 ();
 sg13g2_fill_2 FILLER_13_599 ();
 sg13g2_fill_1 FILLER_13_601 ();
 sg13g2_fill_1 FILLER_13_611 ();
 sg13g2_fill_2 FILLER_13_621 ();
 sg13g2_fill_1 FILLER_13_623 ();
 sg13g2_fill_2 FILLER_13_671 ();
 sg13g2_fill_2 FILLER_13_711 ();
 sg13g2_fill_1 FILLER_13_713 ();
 sg13g2_decap_8 FILLER_13_750 ();
 sg13g2_decap_8 FILLER_13_757 ();
 sg13g2_decap_8 FILLER_13_764 ();
 sg13g2_decap_8 FILLER_13_771 ();
 sg13g2_decap_8 FILLER_13_778 ();
 sg13g2_decap_8 FILLER_13_785 ();
 sg13g2_decap_8 FILLER_13_792 ();
 sg13g2_decap_8 FILLER_13_799 ();
 sg13g2_decap_8 FILLER_13_806 ();
 sg13g2_decap_8 FILLER_13_813 ();
 sg13g2_decap_8 FILLER_13_820 ();
 sg13g2_decap_8 FILLER_13_827 ();
 sg13g2_decap_8 FILLER_13_834 ();
 sg13g2_decap_8 FILLER_13_841 ();
 sg13g2_decap_8 FILLER_13_848 ();
 sg13g2_decap_8 FILLER_13_855 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_28 ();
 sg13g2_fill_1 FILLER_14_30 ();
 sg13g2_fill_2 FILLER_14_40 ();
 sg13g2_fill_2 FILLER_14_123 ();
 sg13g2_fill_2 FILLER_14_158 ();
 sg13g2_fill_1 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_213 ();
 sg13g2_fill_2 FILLER_14_228 ();
 sg13g2_fill_2 FILLER_14_254 ();
 sg13g2_fill_2 FILLER_14_306 ();
 sg13g2_fill_1 FILLER_14_308 ();
 sg13g2_fill_2 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_4 FILLER_14_357 ();
 sg13g2_fill_1 FILLER_14_361 ();
 sg13g2_fill_2 FILLER_14_367 ();
 sg13g2_fill_2 FILLER_14_382 ();
 sg13g2_decap_4 FILLER_14_411 ();
 sg13g2_fill_1 FILLER_14_431 ();
 sg13g2_fill_2 FILLER_14_437 ();
 sg13g2_fill_1 FILLER_14_468 ();
 sg13g2_fill_1 FILLER_14_483 ();
 sg13g2_fill_1 FILLER_14_512 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_fill_2 FILLER_14_588 ();
 sg13g2_fill_1 FILLER_14_590 ();
 sg13g2_fill_1 FILLER_14_627 ();
 sg13g2_fill_2 FILLER_14_663 ();
 sg13g2_fill_2 FILLER_14_675 ();
 sg13g2_fill_1 FILLER_14_677 ();
 sg13g2_fill_2 FILLER_14_713 ();
 sg13g2_fill_1 FILLER_14_715 ();
 sg13g2_fill_2 FILLER_14_726 ();
 sg13g2_decap_8 FILLER_14_758 ();
 sg13g2_decap_8 FILLER_14_765 ();
 sg13g2_decap_8 FILLER_14_772 ();
 sg13g2_decap_8 FILLER_14_779 ();
 sg13g2_decap_8 FILLER_14_786 ();
 sg13g2_decap_8 FILLER_14_793 ();
 sg13g2_decap_8 FILLER_14_800 ();
 sg13g2_decap_8 FILLER_14_807 ();
 sg13g2_decap_8 FILLER_14_814 ();
 sg13g2_decap_8 FILLER_14_821 ();
 sg13g2_decap_8 FILLER_14_828 ();
 sg13g2_decap_8 FILLER_14_835 ();
 sg13g2_decap_8 FILLER_14_842 ();
 sg13g2_decap_8 FILLER_14_849 ();
 sg13g2_decap_4 FILLER_14_856 ();
 sg13g2_fill_2 FILLER_14_860 ();
 sg13g2_fill_2 FILLER_15_26 ();
 sg13g2_fill_1 FILLER_15_28 ();
 sg13g2_fill_2 FILLER_15_39 ();
 sg13g2_fill_2 FILLER_15_50 ();
 sg13g2_fill_1 FILLER_15_75 ();
 sg13g2_fill_2 FILLER_15_109 ();
 sg13g2_fill_1 FILLER_15_111 ();
 sg13g2_fill_2 FILLER_15_126 ();
 sg13g2_fill_1 FILLER_15_128 ();
 sg13g2_fill_2 FILLER_15_155 ();
 sg13g2_fill_1 FILLER_15_157 ();
 sg13g2_fill_2 FILLER_15_184 ();
 sg13g2_fill_1 FILLER_15_206 ();
 sg13g2_fill_1 FILLER_15_233 ();
 sg13g2_fill_2 FILLER_15_275 ();
 sg13g2_fill_1 FILLER_15_277 ();
 sg13g2_fill_1 FILLER_15_306 ();
 sg13g2_fill_2 FILLER_15_370 ();
 sg13g2_fill_2 FILLER_15_398 ();
 sg13g2_fill_2 FILLER_15_490 ();
 sg13g2_fill_1 FILLER_15_492 ();
 sg13g2_fill_2 FILLER_15_519 ();
 sg13g2_fill_1 FILLER_15_521 ();
 sg13g2_decap_8 FILLER_15_526 ();
 sg13g2_fill_2 FILLER_15_533 ();
 sg13g2_fill_2 FILLER_15_608 ();
 sg13g2_fill_1 FILLER_15_651 ();
 sg13g2_fill_1 FILLER_15_661 ();
 sg13g2_fill_1 FILLER_15_695 ();
 sg13g2_decap_8 FILLER_15_765 ();
 sg13g2_decap_8 FILLER_15_772 ();
 sg13g2_decap_8 FILLER_15_779 ();
 sg13g2_decap_8 FILLER_15_786 ();
 sg13g2_decap_8 FILLER_15_793 ();
 sg13g2_decap_8 FILLER_15_800 ();
 sg13g2_decap_8 FILLER_15_807 ();
 sg13g2_decap_8 FILLER_15_814 ();
 sg13g2_decap_8 FILLER_15_821 ();
 sg13g2_decap_8 FILLER_15_828 ();
 sg13g2_decap_8 FILLER_15_835 ();
 sg13g2_decap_8 FILLER_15_842 ();
 sg13g2_decap_8 FILLER_15_849 ();
 sg13g2_decap_4 FILLER_15_856 ();
 sg13g2_fill_2 FILLER_15_860 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_86 ();
 sg13g2_fill_2 FILLER_16_130 ();
 sg13g2_fill_1 FILLER_16_132 ();
 sg13g2_fill_2 FILLER_16_138 ();
 sg13g2_fill_1 FILLER_16_144 ();
 sg13g2_fill_2 FILLER_16_160 ();
 sg13g2_fill_1 FILLER_16_162 ();
 sg13g2_fill_2 FILLER_16_207 ();
 sg13g2_fill_1 FILLER_16_209 ();
 sg13g2_fill_1 FILLER_16_233 ();
 sg13g2_fill_2 FILLER_16_278 ();
 sg13g2_fill_1 FILLER_16_280 ();
 sg13g2_fill_2 FILLER_16_316 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_4 FILLER_16_347 ();
 sg13g2_fill_2 FILLER_16_351 ();
 sg13g2_fill_1 FILLER_16_370 ();
 sg13g2_fill_2 FILLER_16_375 ();
 sg13g2_fill_1 FILLER_16_427 ();
 sg13g2_fill_1 FILLER_16_432 ();
 sg13g2_fill_1 FILLER_16_462 ();
 sg13g2_decap_4 FILLER_16_494 ();
 sg13g2_fill_1 FILLER_16_498 ();
 sg13g2_decap_4 FILLER_16_503 ();
 sg13g2_fill_2 FILLER_16_516 ();
 sg13g2_fill_1 FILLER_16_527 ();
 sg13g2_fill_2 FILLER_16_544 ();
 sg13g2_fill_1 FILLER_16_546 ();
 sg13g2_fill_1 FILLER_16_560 ();
 sg13g2_fill_1 FILLER_16_597 ();
 sg13g2_fill_2 FILLER_16_629 ();
 sg13g2_fill_1 FILLER_16_631 ();
 sg13g2_fill_1 FILLER_16_668 ();
 sg13g2_fill_2 FILLER_16_678 ();
 sg13g2_fill_1 FILLER_16_680 ();
 sg13g2_fill_2 FILLER_16_708 ();
 sg13g2_decap_8 FILLER_16_773 ();
 sg13g2_decap_8 FILLER_16_780 ();
 sg13g2_decap_8 FILLER_16_787 ();
 sg13g2_decap_8 FILLER_16_794 ();
 sg13g2_decap_8 FILLER_16_801 ();
 sg13g2_decap_8 FILLER_16_808 ();
 sg13g2_decap_8 FILLER_16_815 ();
 sg13g2_decap_8 FILLER_16_822 ();
 sg13g2_decap_8 FILLER_16_829 ();
 sg13g2_decap_8 FILLER_16_836 ();
 sg13g2_decap_8 FILLER_16_843 ();
 sg13g2_decap_8 FILLER_16_850 ();
 sg13g2_decap_4 FILLER_16_857 ();
 sg13g2_fill_1 FILLER_16_861 ();
 sg13g2_fill_2 FILLER_17_43 ();
 sg13g2_fill_1 FILLER_17_45 ();
 sg13g2_fill_2 FILLER_17_81 ();
 sg13g2_fill_2 FILLER_17_107 ();
 sg13g2_fill_1 FILLER_17_109 ();
 sg13g2_fill_1 FILLER_17_119 ();
 sg13g2_fill_1 FILLER_17_133 ();
 sg13g2_decap_4 FILLER_17_147 ();
 sg13g2_fill_2 FILLER_17_168 ();
 sg13g2_fill_1 FILLER_17_170 ();
 sg13g2_fill_2 FILLER_17_202 ();
 sg13g2_fill_2 FILLER_17_235 ();
 sg13g2_fill_2 FILLER_17_259 ();
 sg13g2_fill_2 FILLER_17_271 ();
 sg13g2_fill_2 FILLER_17_282 ();
 sg13g2_fill_2 FILLER_17_293 ();
 sg13g2_fill_2 FILLER_17_305 ();
 sg13g2_fill_1 FILLER_17_312 ();
 sg13g2_decap_4 FILLER_17_335 ();
 sg13g2_fill_1 FILLER_17_339 ();
 sg13g2_fill_2 FILLER_17_350 ();
 sg13g2_fill_2 FILLER_17_383 ();
 sg13g2_fill_2 FILLER_17_389 ();
 sg13g2_fill_1 FILLER_17_391 ();
 sg13g2_fill_1 FILLER_17_396 ();
 sg13g2_fill_2 FILLER_17_405 ();
 sg13g2_fill_1 FILLER_17_416 ();
 sg13g2_fill_2 FILLER_17_452 ();
 sg13g2_fill_1 FILLER_17_454 ();
 sg13g2_fill_2 FILLER_17_499 ();
 sg13g2_fill_2 FILLER_17_536 ();
 sg13g2_fill_1 FILLER_17_538 ();
 sg13g2_fill_1 FILLER_17_548 ();
 sg13g2_fill_2 FILLER_17_595 ();
 sg13g2_fill_2 FILLER_17_613 ();
 sg13g2_fill_1 FILLER_17_615 ();
 sg13g2_fill_1 FILLER_17_697 ();
 sg13g2_decap_8 FILLER_17_778 ();
 sg13g2_decap_8 FILLER_17_785 ();
 sg13g2_decap_8 FILLER_17_792 ();
 sg13g2_decap_8 FILLER_17_799 ();
 sg13g2_decap_8 FILLER_17_806 ();
 sg13g2_decap_8 FILLER_17_813 ();
 sg13g2_decap_8 FILLER_17_820 ();
 sg13g2_decap_8 FILLER_17_827 ();
 sg13g2_decap_8 FILLER_17_834 ();
 sg13g2_decap_8 FILLER_17_841 ();
 sg13g2_decap_8 FILLER_17_848 ();
 sg13g2_decap_8 FILLER_17_855 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_37 ();
 sg13g2_fill_2 FILLER_18_64 ();
 sg13g2_decap_4 FILLER_18_151 ();
 sg13g2_decap_8 FILLER_18_178 ();
 sg13g2_fill_1 FILLER_18_185 ();
 sg13g2_fill_2 FILLER_18_190 ();
 sg13g2_decap_8 FILLER_18_214 ();
 sg13g2_decap_4 FILLER_18_221 ();
 sg13g2_fill_2 FILLER_18_364 ();
 sg13g2_fill_2 FILLER_18_370 ();
 sg13g2_fill_1 FILLER_18_372 ();
 sg13g2_decap_8 FILLER_18_377 ();
 sg13g2_fill_1 FILLER_18_384 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_fill_2 FILLER_18_449 ();
 sg13g2_fill_1 FILLER_18_475 ();
 sg13g2_fill_2 FILLER_18_507 ();
 sg13g2_fill_2 FILLER_18_558 ();
 sg13g2_fill_1 FILLER_18_576 ();
 sg13g2_fill_2 FILLER_18_582 ();
 sg13g2_fill_2 FILLER_18_650 ();
 sg13g2_fill_2 FILLER_18_714 ();
 sg13g2_fill_1 FILLER_18_716 ();
 sg13g2_fill_1 FILLER_18_727 ();
 sg13g2_fill_1 FILLER_18_737 ();
 sg13g2_decap_8 FILLER_18_778 ();
 sg13g2_decap_8 FILLER_18_785 ();
 sg13g2_decap_8 FILLER_18_792 ();
 sg13g2_decap_8 FILLER_18_799 ();
 sg13g2_decap_8 FILLER_18_806 ();
 sg13g2_decap_8 FILLER_18_813 ();
 sg13g2_decap_8 FILLER_18_820 ();
 sg13g2_decap_8 FILLER_18_827 ();
 sg13g2_decap_8 FILLER_18_834 ();
 sg13g2_decap_8 FILLER_18_841 ();
 sg13g2_decap_8 FILLER_18_848 ();
 sg13g2_decap_8 FILLER_18_855 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_7 ();
 sg13g2_fill_1 FILLER_19_9 ();
 sg13g2_fill_2 FILLER_19_23 ();
 sg13g2_fill_1 FILLER_19_43 ();
 sg13g2_fill_2 FILLER_19_72 ();
 sg13g2_fill_2 FILLER_19_83 ();
 sg13g2_fill_1 FILLER_19_85 ();
 sg13g2_fill_2 FILLER_19_95 ();
 sg13g2_fill_2 FILLER_19_110 ();
 sg13g2_fill_2 FILLER_19_117 ();
 sg13g2_fill_1 FILLER_19_119 ();
 sg13g2_fill_2 FILLER_19_130 ();
 sg13g2_decap_4 FILLER_19_168 ();
 sg13g2_fill_1 FILLER_19_207 ();
 sg13g2_fill_2 FILLER_19_244 ();
 sg13g2_fill_1 FILLER_19_285 ();
 sg13g2_fill_2 FILLER_19_320 ();
 sg13g2_fill_2 FILLER_19_336 ();
 sg13g2_fill_1 FILLER_19_338 ();
 sg13g2_fill_2 FILLER_19_402 ();
 sg13g2_fill_1 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_418 ();
 sg13g2_fill_2 FILLER_19_441 ();
 sg13g2_fill_2 FILLER_19_452 ();
 sg13g2_fill_2 FILLER_19_531 ();
 sg13g2_fill_1 FILLER_19_533 ();
 sg13g2_fill_2 FILLER_19_546 ();
 sg13g2_fill_1 FILLER_19_548 ();
 sg13g2_decap_4 FILLER_19_552 ();
 sg13g2_fill_1 FILLER_19_556 ();
 sg13g2_fill_1 FILLER_19_568 ();
 sg13g2_fill_1 FILLER_19_586 ();
 sg13g2_fill_1 FILLER_19_591 ();
 sg13g2_fill_1 FILLER_19_598 ();
 sg13g2_fill_2 FILLER_19_611 ();
 sg13g2_fill_2 FILLER_19_654 ();
 sg13g2_fill_1 FILLER_19_739 ();
 sg13g2_fill_1 FILLER_19_755 ();
 sg13g2_decap_8 FILLER_19_782 ();
 sg13g2_decap_8 FILLER_19_789 ();
 sg13g2_decap_8 FILLER_19_796 ();
 sg13g2_decap_8 FILLER_19_803 ();
 sg13g2_decap_8 FILLER_19_810 ();
 sg13g2_decap_8 FILLER_19_817 ();
 sg13g2_decap_8 FILLER_19_824 ();
 sg13g2_decap_8 FILLER_19_831 ();
 sg13g2_decap_8 FILLER_19_838 ();
 sg13g2_decap_8 FILLER_19_845 ();
 sg13g2_decap_8 FILLER_19_852 ();
 sg13g2_fill_2 FILLER_19_859 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_fill_1 FILLER_20_26 ();
 sg13g2_fill_1 FILLER_20_37 ();
 sg13g2_fill_2 FILLER_20_107 ();
 sg13g2_fill_2 FILLER_20_128 ();
 sg13g2_decap_4 FILLER_20_161 ();
 sg13g2_fill_1 FILLER_20_165 ();
 sg13g2_fill_2 FILLER_20_225 ();
 sg13g2_fill_1 FILLER_20_227 ();
 sg13g2_fill_2 FILLER_20_237 ();
 sg13g2_fill_1 FILLER_20_273 ();
 sg13g2_decap_4 FILLER_20_304 ();
 sg13g2_decap_8 FILLER_20_368 ();
 sg13g2_fill_1 FILLER_20_375 ();
 sg13g2_fill_2 FILLER_20_412 ();
 sg13g2_fill_1 FILLER_20_463 ();
 sg13g2_fill_1 FILLER_20_481 ();
 sg13g2_fill_2 FILLER_20_516 ();
 sg13g2_decap_8 FILLER_20_555 ();
 sg13g2_fill_1 FILLER_20_573 ();
 sg13g2_fill_2 FILLER_20_586 ();
 sg13g2_fill_1 FILLER_20_588 ();
 sg13g2_fill_2 FILLER_20_601 ();
 sg13g2_fill_1 FILLER_20_603 ();
 sg13g2_fill_2 FILLER_20_657 ();
 sg13g2_fill_1 FILLER_20_702 ();
 sg13g2_fill_2 FILLER_20_712 ();
 sg13g2_fill_1 FILLER_20_714 ();
 sg13g2_decap_8 FILLER_20_786 ();
 sg13g2_decap_8 FILLER_20_793 ();
 sg13g2_decap_8 FILLER_20_800 ();
 sg13g2_decap_8 FILLER_20_807 ();
 sg13g2_decap_8 FILLER_20_814 ();
 sg13g2_fill_2 FILLER_20_821 ();
 sg13g2_fill_1 FILLER_20_823 ();
 sg13g2_decap_8 FILLER_20_828 ();
 sg13g2_decap_8 FILLER_20_835 ();
 sg13g2_decap_8 FILLER_20_842 ();
 sg13g2_decap_8 FILLER_20_849 ();
 sg13g2_decap_4 FILLER_20_856 ();
 sg13g2_fill_2 FILLER_20_860 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_4 ();
 sg13g2_fill_2 FILLER_21_73 ();
 sg13g2_fill_1 FILLER_21_75 ();
 sg13g2_fill_1 FILLER_21_80 ();
 sg13g2_fill_2 FILLER_21_104 ();
 sg13g2_fill_1 FILLER_21_106 ();
 sg13g2_fill_2 FILLER_21_116 ();
 sg13g2_fill_1 FILLER_21_124 ();
 sg13g2_fill_2 FILLER_21_130 ();
 sg13g2_decap_8 FILLER_21_214 ();
 sg13g2_decap_4 FILLER_21_221 ();
 sg13g2_fill_2 FILLER_21_225 ();
 sg13g2_fill_2 FILLER_21_264 ();
 sg13g2_fill_2 FILLER_21_305 ();
 sg13g2_decap_4 FILLER_21_311 ();
 sg13g2_fill_2 FILLER_21_350 ();
 sg13g2_fill_2 FILLER_21_392 ();
 sg13g2_fill_2 FILLER_21_420 ();
 sg13g2_fill_1 FILLER_21_422 ();
 sg13g2_fill_2 FILLER_21_437 ();
 sg13g2_fill_1 FILLER_21_439 ();
 sg13g2_fill_1 FILLER_21_472 ();
 sg13g2_fill_2 FILLER_21_513 ();
 sg13g2_fill_1 FILLER_21_555 ();
 sg13g2_decap_4 FILLER_21_576 ();
 sg13g2_fill_2 FILLER_21_605 ();
 sg13g2_fill_2 FILLER_21_611 ();
 sg13g2_fill_2 FILLER_21_623 ();
 sg13g2_fill_1 FILLER_21_625 ();
 sg13g2_fill_2 FILLER_21_720 ();
 sg13g2_fill_2 FILLER_21_767 ();
 sg13g2_fill_1 FILLER_21_769 ();
 sg13g2_decap_8 FILLER_21_800 ();
 sg13g2_decap_4 FILLER_21_807 ();
 sg13g2_fill_1 FILLER_21_811 ();
 sg13g2_decap_8 FILLER_21_839 ();
 sg13g2_decap_8 FILLER_21_846 ();
 sg13g2_decap_8 FILLER_21_853 ();
 sg13g2_fill_2 FILLER_21_860 ();
 sg13g2_decap_4 FILLER_22_40 ();
 sg13g2_fill_1 FILLER_22_44 ();
 sg13g2_fill_2 FILLER_22_59 ();
 sg13g2_fill_1 FILLER_22_61 ();
 sg13g2_fill_2 FILLER_22_70 ();
 sg13g2_fill_2 FILLER_22_107 ();
 sg13g2_fill_1 FILLER_22_109 ();
 sg13g2_fill_2 FILLER_22_120 ();
 sg13g2_fill_1 FILLER_22_122 ();
 sg13g2_fill_2 FILLER_22_149 ();
 sg13g2_fill_2 FILLER_22_183 ();
 sg13g2_fill_1 FILLER_22_185 ();
 sg13g2_decap_4 FILLER_22_199 ();
 sg13g2_fill_1 FILLER_22_203 ();
 sg13g2_fill_1 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_248 ();
 sg13g2_fill_1 FILLER_22_255 ();
 sg13g2_fill_2 FILLER_22_290 ();
 sg13g2_fill_2 FILLER_22_326 ();
 sg13g2_fill_2 FILLER_22_368 ();
 sg13g2_fill_1 FILLER_22_370 ();
 sg13g2_fill_2 FILLER_22_423 ();
 sg13g2_fill_2 FILLER_22_434 ();
 sg13g2_decap_8 FILLER_22_481 ();
 sg13g2_fill_2 FILLER_22_488 ();
 sg13g2_decap_8 FILLER_22_509 ();
 sg13g2_fill_2 FILLER_22_526 ();
 sg13g2_fill_1 FILLER_22_564 ();
 sg13g2_fill_1 FILLER_22_579 ();
 sg13g2_fill_2 FILLER_22_607 ();
 sg13g2_fill_1 FILLER_22_651 ();
 sg13g2_decap_4 FILLER_22_666 ();
 sg13g2_decap_4 FILLER_22_679 ();
 sg13g2_fill_2 FILLER_22_693 ();
 sg13g2_fill_2 FILLER_22_744 ();
 sg13g2_fill_1 FILLER_22_755 ();
 sg13g2_fill_1 FILLER_22_792 ();
 sg13g2_fill_2 FILLER_22_807 ();
 sg13g2_decap_4 FILLER_22_857 ();
 sg13g2_fill_1 FILLER_22_861 ();
 sg13g2_fill_2 FILLER_23_80 ();
 sg13g2_fill_2 FILLER_23_91 ();
 sg13g2_decap_4 FILLER_23_203 ();
 sg13g2_fill_1 FILLER_23_225 ();
 sg13g2_fill_2 FILLER_23_252 ();
 sg13g2_fill_1 FILLER_23_289 ();
 sg13g2_fill_1 FILLER_23_299 ();
 sg13g2_fill_2 FILLER_23_308 ();
 sg13g2_fill_2 FILLER_23_384 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_415 ();
 sg13g2_fill_1 FILLER_23_422 ();
 sg13g2_decap_4 FILLER_23_438 ();
 sg13g2_decap_8 FILLER_23_456 ();
 sg13g2_fill_2 FILLER_23_463 ();
 sg13g2_decap_8 FILLER_23_474 ();
 sg13g2_fill_1 FILLER_23_481 ();
 sg13g2_fill_2 FILLER_23_485 ();
 sg13g2_fill_2 FILLER_23_526 ();
 sg13g2_fill_1 FILLER_23_528 ();
 sg13g2_decap_4 FILLER_23_534 ();
 sg13g2_fill_1 FILLER_23_538 ();
 sg13g2_decap_8 FILLER_23_544 ();
 sg13g2_fill_2 FILLER_23_556 ();
 sg13g2_decap_8 FILLER_23_603 ();
 sg13g2_fill_1 FILLER_23_610 ();
 sg13g2_fill_1 FILLER_23_621 ();
 sg13g2_decap_8 FILLER_23_626 ();
 sg13g2_fill_2 FILLER_23_633 ();
 sg13g2_decap_8 FILLER_23_640 ();
 sg13g2_fill_1 FILLER_23_647 ();
 sg13g2_decap_4 FILLER_23_684 ();
 sg13g2_fill_2 FILLER_23_714 ();
 sg13g2_fill_1 FILLER_23_716 ();
 sg13g2_fill_1 FILLER_23_772 ();
 sg13g2_fill_2 FILLER_23_832 ();
 sg13g2_fill_1 FILLER_23_834 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_4 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_18 ();
 sg13g2_fill_1 FILLER_24_56 ();
 sg13g2_fill_2 FILLER_24_62 ();
 sg13g2_fill_2 FILLER_24_73 ();
 sg13g2_fill_1 FILLER_24_75 ();
 sg13g2_fill_1 FILLER_24_90 ();
 sg13g2_fill_2 FILLER_24_100 ();
 sg13g2_fill_2 FILLER_24_110 ();
 sg13g2_fill_2 FILLER_24_135 ();
 sg13g2_fill_2 FILLER_24_145 ();
 sg13g2_fill_1 FILLER_24_162 ();
 sg13g2_fill_1 FILLER_24_195 ();
 sg13g2_decap_8 FILLER_24_232 ();
 sg13g2_decap_4 FILLER_24_245 ();
 sg13g2_fill_2 FILLER_24_309 ();
 sg13g2_fill_1 FILLER_24_345 ();
 sg13g2_fill_2 FILLER_24_351 ();
 sg13g2_fill_2 FILLER_24_357 ();
 sg13g2_fill_2 FILLER_24_423 ();
 sg13g2_fill_1 FILLER_24_490 ();
 sg13g2_fill_2 FILLER_24_504 ();
 sg13g2_fill_2 FILLER_24_510 ();
 sg13g2_fill_1 FILLER_24_512 ();
 sg13g2_fill_1 FILLER_24_534 ();
 sg13g2_fill_1 FILLER_24_561 ();
 sg13g2_fill_2 FILLER_24_576 ();
 sg13g2_fill_2 FILLER_24_583 ();
 sg13g2_fill_2 FILLER_24_599 ();
 sg13g2_fill_1 FILLER_24_653 ();
 sg13g2_fill_1 FILLER_24_690 ();
 sg13g2_fill_2 FILLER_24_696 ();
 sg13g2_fill_1 FILLER_24_698 ();
 sg13g2_fill_2 FILLER_24_737 ();
 sg13g2_fill_2 FILLER_24_748 ();
 sg13g2_fill_1 FILLER_24_750 ();
 sg13g2_fill_1 FILLER_24_777 ();
 sg13g2_fill_2 FILLER_24_837 ();
 sg13g2_fill_1 FILLER_24_839 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_91 ();
 sg13g2_fill_2 FILLER_25_102 ();
 sg13g2_fill_1 FILLER_25_130 ();
 sg13g2_decap_4 FILLER_25_166 ();
 sg13g2_decap_4 FILLER_25_176 ();
 sg13g2_decap_4 FILLER_25_197 ();
 sg13g2_fill_2 FILLER_25_207 ();
 sg13g2_fill_1 FILLER_25_209 ();
 sg13g2_fill_1 FILLER_25_221 ();
 sg13g2_decap_8 FILLER_25_225 ();
 sg13g2_fill_2 FILLER_25_232 ();
 sg13g2_fill_1 FILLER_25_234 ();
 sg13g2_fill_2 FILLER_25_266 ();
 sg13g2_fill_1 FILLER_25_292 ();
 sg13g2_fill_2 FILLER_25_334 ();
 sg13g2_fill_1 FILLER_25_336 ();
 sg13g2_fill_1 FILLER_25_342 ();
 sg13g2_fill_2 FILLER_25_409 ();
 sg13g2_fill_1 FILLER_25_424 ();
 sg13g2_fill_1 FILLER_25_443 ();
 sg13g2_decap_8 FILLER_25_464 ();
 sg13g2_decap_8 FILLER_25_471 ();
 sg13g2_decap_4 FILLER_25_478 ();
 sg13g2_fill_1 FILLER_25_494 ();
 sg13g2_fill_1 FILLER_25_521 ();
 sg13g2_decap_8 FILLER_25_531 ();
 sg13g2_fill_1 FILLER_25_538 ();
 sg13g2_fill_2 FILLER_25_568 ();
 sg13g2_fill_2 FILLER_25_605 ();
 sg13g2_fill_1 FILLER_25_607 ();
 sg13g2_decap_8 FILLER_25_624 ();
 sg13g2_decap_4 FILLER_25_631 ();
 sg13g2_fill_1 FILLER_25_635 ();
 sg13g2_decap_8 FILLER_25_644 ();
 sg13g2_fill_2 FILLER_25_664 ();
 sg13g2_fill_2 FILLER_25_699 ();
 sg13g2_fill_1 FILLER_25_749 ();
 sg13g2_fill_2 FILLER_25_776 ();
 sg13g2_fill_1 FILLER_25_809 ();
 sg13g2_fill_1 FILLER_25_824 ();
 sg13g2_fill_1 FILLER_25_861 ();
 sg13g2_fill_2 FILLER_26_36 ();
 sg13g2_fill_1 FILLER_26_57 ();
 sg13g2_decap_4 FILLER_26_87 ();
 sg13g2_fill_1 FILLER_26_136 ();
 sg13g2_fill_2 FILLER_26_145 ();
 sg13g2_decap_4 FILLER_26_166 ();
 sg13g2_fill_1 FILLER_26_176 ();
 sg13g2_fill_2 FILLER_26_195 ();
 sg13g2_fill_1 FILLER_26_217 ();
 sg13g2_fill_2 FILLER_26_244 ();
 sg13g2_fill_2 FILLER_26_273 ();
 sg13g2_fill_2 FILLER_26_288 ();
 sg13g2_fill_1 FILLER_26_336 ();
 sg13g2_fill_1 FILLER_26_347 ();
 sg13g2_fill_1 FILLER_26_407 ();
 sg13g2_fill_1 FILLER_26_428 ();
 sg13g2_fill_2 FILLER_26_442 ();
 sg13g2_fill_1 FILLER_26_534 ();
 sg13g2_fill_1 FILLER_26_594 ();
 sg13g2_fill_2 FILLER_26_605 ();
 sg13g2_fill_1 FILLER_26_607 ();
 sg13g2_decap_8 FILLER_26_631 ();
 sg13g2_decap_4 FILLER_26_648 ();
 sg13g2_fill_1 FILLER_26_652 ();
 sg13g2_decap_4 FILLER_26_658 ();
 sg13g2_fill_1 FILLER_26_662 ();
 sg13g2_fill_2 FILLER_26_721 ();
 sg13g2_fill_2 FILLER_26_729 ();
 sg13g2_fill_1 FILLER_26_731 ();
 sg13g2_fill_1 FILLER_26_739 ();
 sg13g2_fill_1 FILLER_26_846 ();
 sg13g2_fill_1 FILLER_26_861 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_7 ();
 sg13g2_fill_1 FILLER_27_9 ();
 sg13g2_decap_4 FILLER_27_44 ();
 sg13g2_decap_4 FILLER_27_74 ();
 sg13g2_decap_4 FILLER_27_166 ();
 sg13g2_fill_1 FILLER_27_170 ();
 sg13g2_fill_1 FILLER_27_185 ();
 sg13g2_fill_2 FILLER_27_200 ();
 sg13g2_fill_2 FILLER_27_296 ();
 sg13g2_fill_1 FILLER_27_298 ();
 sg13g2_fill_2 FILLER_27_321 ();
 sg13g2_fill_1 FILLER_27_341 ();
 sg13g2_fill_2 FILLER_27_364 ();
 sg13g2_fill_1 FILLER_27_366 ();
 sg13g2_fill_2 FILLER_27_436 ();
 sg13g2_decap_4 FILLER_27_443 ();
 sg13g2_fill_1 FILLER_27_447 ();
 sg13g2_fill_1 FILLER_27_455 ();
 sg13g2_fill_1 FILLER_27_468 ();
 sg13g2_fill_2 FILLER_27_493 ();
 sg13g2_decap_4 FILLER_27_562 ();
 sg13g2_fill_1 FILLER_27_570 ();
 sg13g2_fill_2 FILLER_27_588 ();
 sg13g2_fill_2 FILLER_27_612 ();
 sg13g2_fill_1 FILLER_27_614 ();
 sg13g2_fill_2 FILLER_27_693 ();
 sg13g2_fill_1 FILLER_27_695 ();
 sg13g2_fill_2 FILLER_27_708 ();
 sg13g2_fill_1 FILLER_27_710 ();
 sg13g2_fill_1 FILLER_27_753 ();
 sg13g2_fill_2 FILLER_27_780 ();
 sg13g2_fill_1 FILLER_27_782 ();
 sg13g2_fill_1 FILLER_27_805 ();
 sg13g2_fill_1 FILLER_28_26 ();
 sg13g2_fill_1 FILLER_28_32 ();
 sg13g2_fill_2 FILLER_28_52 ();
 sg13g2_fill_1 FILLER_28_58 ();
 sg13g2_decap_4 FILLER_28_63 ();
 sg13g2_fill_2 FILLER_28_67 ();
 sg13g2_decap_4 FILLER_28_78 ();
 sg13g2_fill_1 FILLER_28_82 ();
 sg13g2_decap_8 FILLER_28_114 ();
 sg13g2_decap_8 FILLER_28_134 ();
 sg13g2_decap_8 FILLER_28_149 ();
 sg13g2_fill_2 FILLER_28_156 ();
 sg13g2_fill_1 FILLER_28_158 ();
 sg13g2_fill_1 FILLER_28_168 ();
 sg13g2_fill_1 FILLER_28_187 ();
 sg13g2_fill_1 FILLER_28_223 ();
 sg13g2_fill_2 FILLER_28_250 ();
 sg13g2_fill_1 FILLER_28_252 ();
 sg13g2_fill_2 FILLER_28_261 ();
 sg13g2_fill_2 FILLER_28_276 ();
 sg13g2_fill_2 FILLER_28_342 ();
 sg13g2_fill_1 FILLER_28_430 ();
 sg13g2_fill_2 FILLER_28_485 ();
 sg13g2_fill_2 FILLER_28_492 ();
 sg13g2_decap_8 FILLER_28_512 ();
 sg13g2_fill_2 FILLER_28_519 ();
 sg13g2_decap_4 FILLER_28_538 ();
 sg13g2_fill_1 FILLER_28_590 ();
 sg13g2_decap_4 FILLER_28_596 ();
 sg13g2_fill_2 FILLER_28_608 ();
 sg13g2_fill_2 FILLER_28_623 ();
 sg13g2_fill_1 FILLER_28_625 ();
 sg13g2_fill_2 FILLER_28_644 ();
 sg13g2_fill_1 FILLER_28_646 ();
 sg13g2_decap_8 FILLER_28_651 ();
 sg13g2_fill_2 FILLER_28_658 ();
 sg13g2_fill_1 FILLER_28_660 ();
 sg13g2_fill_1 FILLER_28_669 ();
 sg13g2_decap_4 FILLER_28_697 ();
 sg13g2_fill_2 FILLER_28_701 ();
 sg13g2_fill_2 FILLER_28_708 ();
 sg13g2_fill_1 FILLER_28_732 ();
 sg13g2_fill_2 FILLER_28_749 ();
 sg13g2_fill_1 FILLER_28_751 ();
 sg13g2_fill_1 FILLER_28_757 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_61 ();
 sg13g2_fill_2 FILLER_29_67 ();
 sg13g2_fill_1 FILLER_29_69 ();
 sg13g2_fill_1 FILLER_29_79 ();
 sg13g2_fill_2 FILLER_29_85 ();
 sg13g2_fill_2 FILLER_29_137 ();
 sg13g2_decap_4 FILLER_29_180 ();
 sg13g2_decap_4 FILLER_29_189 ();
 sg13g2_fill_1 FILLER_29_193 ();
 sg13g2_decap_4 FILLER_29_259 ();
 sg13g2_fill_1 FILLER_29_263 ();
 sg13g2_fill_2 FILLER_29_272 ();
 sg13g2_fill_1 FILLER_29_300 ();
 sg13g2_fill_1 FILLER_29_314 ();
 sg13g2_fill_2 FILLER_29_341 ();
 sg13g2_fill_1 FILLER_29_343 ();
 sg13g2_fill_2 FILLER_29_352 ();
 sg13g2_fill_1 FILLER_29_354 ();
 sg13g2_fill_2 FILLER_29_364 ();
 sg13g2_fill_2 FILLER_29_389 ();
 sg13g2_fill_2 FILLER_29_422 ();
 sg13g2_decap_4 FILLER_29_457 ();
 sg13g2_fill_2 FILLER_29_461 ();
 sg13g2_fill_2 FILLER_29_487 ();
 sg13g2_fill_1 FILLER_29_489 ();
 sg13g2_decap_4 FILLER_29_525 ();
 sg13g2_fill_1 FILLER_29_529 ();
 sg13g2_decap_8 FILLER_29_562 ();
 sg13g2_decap_8 FILLER_29_569 ();
 sg13g2_decap_4 FILLER_29_576 ();
 sg13g2_fill_2 FILLER_29_580 ();
 sg13g2_fill_1 FILLER_29_596 ();
 sg13g2_decap_4 FILLER_29_638 ();
 sg13g2_fill_1 FILLER_29_642 ();
 sg13g2_fill_2 FILLER_29_647 ();
 sg13g2_fill_2 FILLER_29_668 ();
 sg13g2_fill_1 FILLER_29_675 ();
 sg13g2_fill_1 FILLER_29_714 ();
 sg13g2_fill_2 FILLER_29_729 ();
 sg13g2_decap_4 FILLER_29_817 ();
 sg13g2_fill_1 FILLER_29_831 ();
 sg13g2_decap_4 FILLER_29_858 ();
 sg13g2_fill_1 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_187 ();
 sg13g2_decap_8 FILLER_30_202 ();
 sg13g2_fill_1 FILLER_30_209 ();
 sg13g2_fill_2 FILLER_30_231 ();
 sg13g2_fill_1 FILLER_30_233 ();
 sg13g2_fill_2 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_260 ();
 sg13g2_fill_1 FILLER_30_329 ();
 sg13g2_fill_2 FILLER_30_350 ();
 sg13g2_fill_1 FILLER_30_352 ();
 sg13g2_fill_1 FILLER_30_379 ();
 sg13g2_fill_1 FILLER_30_393 ();
 sg13g2_fill_2 FILLER_30_416 ();
 sg13g2_fill_2 FILLER_30_427 ();
 sg13g2_fill_2 FILLER_30_440 ();
 sg13g2_fill_1 FILLER_30_442 ();
 sg13g2_decap_4 FILLER_30_455 ();
 sg13g2_fill_2 FILLER_30_468 ();
 sg13g2_fill_1 FILLER_30_470 ();
 sg13g2_fill_1 FILLER_30_509 ();
 sg13g2_decap_8 FILLER_30_514 ();
 sg13g2_fill_1 FILLER_30_521 ();
 sg13g2_decap_8 FILLER_30_532 ();
 sg13g2_fill_1 FILLER_30_539 ();
 sg13g2_fill_2 FILLER_30_553 ();
 sg13g2_fill_1 FILLER_30_591 ();
 sg13g2_fill_1 FILLER_30_601 ();
 sg13g2_fill_2 FILLER_30_605 ();
 sg13g2_fill_1 FILLER_30_622 ();
 sg13g2_decap_4 FILLER_30_628 ();
 sg13g2_fill_2 FILLER_30_658 ();
 sg13g2_fill_1 FILLER_30_674 ();
 sg13g2_decap_8 FILLER_30_700 ();
 sg13g2_fill_2 FILLER_30_707 ();
 sg13g2_fill_2 FILLER_30_775 ();
 sg13g2_fill_1 FILLER_30_813 ();
 sg13g2_fill_1 FILLER_30_846 ();
 sg13g2_decap_4 FILLER_30_857 ();
 sg13g2_fill_1 FILLER_30_861 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_4 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_15 ();
 sg13g2_fill_1 FILLER_31_57 ();
 sg13g2_fill_1 FILLER_31_81 ();
 sg13g2_fill_2 FILLER_31_114 ();
 sg13g2_fill_1 FILLER_31_116 ();
 sg13g2_fill_2 FILLER_31_141 ();
 sg13g2_fill_1 FILLER_31_143 ();
 sg13g2_fill_1 FILLER_31_186 ();
 sg13g2_fill_1 FILLER_31_195 ();
 sg13g2_decap_4 FILLER_31_213 ();
 sg13g2_fill_2 FILLER_31_248 ();
 sg13g2_fill_1 FILLER_31_284 ();
 sg13g2_fill_2 FILLER_31_317 ();
 sg13g2_fill_2 FILLER_31_373 ();
 sg13g2_fill_1 FILLER_31_467 ();
 sg13g2_fill_2 FILLER_31_494 ();
 sg13g2_decap_4 FILLER_31_509 ();
 sg13g2_fill_1 FILLER_31_539 ();
 sg13g2_fill_2 FILLER_31_559 ();
 sg13g2_fill_1 FILLER_31_561 ();
 sg13g2_fill_1 FILLER_31_571 ();
 sg13g2_fill_2 FILLER_31_603 ();
 sg13g2_fill_2 FILLER_31_626 ();
 sg13g2_fill_1 FILLER_31_628 ();
 sg13g2_fill_2 FILLER_31_634 ();
 sg13g2_fill_1 FILLER_31_636 ();
 sg13g2_fill_2 FILLER_31_641 ();
 sg13g2_fill_1 FILLER_31_643 ();
 sg13g2_fill_1 FILLER_31_652 ();
 sg13g2_fill_1 FILLER_31_677 ();
 sg13g2_fill_2 FILLER_31_744 ();
 sg13g2_fill_1 FILLER_31_746 ();
 sg13g2_fill_2 FILLER_31_783 ();
 sg13g2_fill_1 FILLER_31_794 ();
 sg13g2_fill_1 FILLER_31_838 ();
 sg13g2_decap_4 FILLER_31_857 ();
 sg13g2_fill_1 FILLER_31_861 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_38 ();
 sg13g2_fill_1 FILLER_32_54 ();
 sg13g2_fill_2 FILLER_32_114 ();
 sg13g2_fill_2 FILLER_32_152 ();
 sg13g2_fill_2 FILLER_32_190 ();
 sg13g2_fill_1 FILLER_32_192 ();
 sg13g2_fill_2 FILLER_32_201 ();
 sg13g2_fill_1 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_228 ();
 sg13g2_fill_1 FILLER_32_235 ();
 sg13g2_decap_8 FILLER_32_241 ();
 sg13g2_decap_4 FILLER_32_248 ();
 sg13g2_fill_2 FILLER_32_252 ();
 sg13g2_fill_2 FILLER_32_330 ();
 sg13g2_fill_2 FILLER_32_353 ();
 sg13g2_fill_1 FILLER_32_355 ();
 sg13g2_fill_1 FILLER_32_377 ();
 sg13g2_fill_1 FILLER_32_404 ();
 sg13g2_decap_4 FILLER_32_530 ();
 sg13g2_decap_4 FILLER_32_619 ();
 sg13g2_fill_1 FILLER_32_623 ();
 sg13g2_fill_1 FILLER_32_632 ();
 sg13g2_decap_4 FILLER_32_659 ();
 sg13g2_decap_8 FILLER_32_689 ();
 sg13g2_fill_1 FILLER_32_696 ();
 sg13g2_fill_1 FILLER_32_759 ();
 sg13g2_fill_2 FILLER_32_818 ();
 sg13g2_fill_1 FILLER_32_820 ();
 sg13g2_decap_4 FILLER_32_858 ();
 sg13g2_fill_1 FILLER_33_26 ();
 sg13g2_fill_2 FILLER_33_37 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_4 FILLER_33_56 ();
 sg13g2_fill_2 FILLER_33_60 ();
 sg13g2_fill_2 FILLER_33_84 ();
 sg13g2_fill_2 FILLER_33_106 ();
 sg13g2_fill_1 FILLER_33_108 ();
 sg13g2_fill_1 FILLER_33_151 ();
 sg13g2_fill_2 FILLER_33_165 ();
 sg13g2_decap_4 FILLER_33_208 ();
 sg13g2_fill_2 FILLER_33_236 ();
 sg13g2_decap_4 FILLER_33_264 ();
 sg13g2_fill_1 FILLER_33_268 ();
 sg13g2_fill_2 FILLER_33_331 ();
 sg13g2_fill_2 FILLER_33_355 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_decap_4 FILLER_33_389 ();
 sg13g2_fill_2 FILLER_33_422 ();
 sg13g2_fill_1 FILLER_33_424 ();
 sg13g2_decap_8 FILLER_33_504 ();
 sg13g2_fill_1 FILLER_33_511 ();
 sg13g2_fill_1 FILLER_33_588 ();
 sg13g2_fill_2 FILLER_33_594 ();
 sg13g2_fill_2 FILLER_33_614 ();
 sg13g2_decap_4 FILLER_33_639 ();
 sg13g2_decap_4 FILLER_33_669 ();
 sg13g2_fill_2 FILLER_33_677 ();
 sg13g2_fill_1 FILLER_33_684 ();
 sg13g2_fill_1 FILLER_33_727 ();
 sg13g2_fill_2 FILLER_33_742 ();
 sg13g2_fill_1 FILLER_33_744 ();
 sg13g2_fill_1 FILLER_33_765 ();
 sg13g2_fill_2 FILLER_33_860 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_46 ();
 sg13g2_fill_1 FILLER_34_50 ();
 sg13g2_fill_1 FILLER_34_105 ();
 sg13g2_fill_2 FILLER_34_111 ();
 sg13g2_fill_1 FILLER_34_168 ();
 sg13g2_fill_2 FILLER_34_174 ();
 sg13g2_fill_1 FILLER_34_176 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_4 FILLER_34_203 ();
 sg13g2_fill_1 FILLER_34_207 ();
 sg13g2_decap_4 FILLER_34_263 ();
 sg13g2_fill_2 FILLER_34_398 ();
 sg13g2_decap_4 FILLER_34_406 ();
 sg13g2_fill_2 FILLER_34_410 ();
 sg13g2_fill_2 FILLER_34_452 ();
 sg13g2_decap_4 FILLER_34_504 ();
 sg13g2_fill_1 FILLER_34_508 ();
 sg13g2_decap_8 FILLER_34_517 ();
 sg13g2_fill_2 FILLER_34_524 ();
 sg13g2_fill_2 FILLER_34_549 ();
 sg13g2_fill_1 FILLER_34_551 ();
 sg13g2_fill_2 FILLER_34_578 ();
 sg13g2_fill_1 FILLER_34_606 ();
 sg13g2_fill_2 FILLER_34_616 ();
 sg13g2_decap_4 FILLER_34_635 ();
 sg13g2_fill_2 FILLER_34_648 ();
 sg13g2_fill_1 FILLER_34_650 ();
 sg13g2_decap_4 FILLER_34_668 ();
 sg13g2_fill_1 FILLER_34_672 ();
 sg13g2_fill_1 FILLER_34_730 ();
 sg13g2_fill_2 FILLER_34_783 ();
 sg13g2_fill_1 FILLER_34_785 ();
 sg13g2_decap_4 FILLER_34_843 ();
 sg13g2_decap_4 FILLER_34_858 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_18 ();
 sg13g2_fill_1 FILLER_35_33 ();
 sg13g2_fill_1 FILLER_35_53 ();
 sg13g2_fill_2 FILLER_35_71 ();
 sg13g2_fill_1 FILLER_35_85 ();
 sg13g2_fill_1 FILLER_35_100 ();
 sg13g2_fill_2 FILLER_35_113 ();
 sg13g2_fill_1 FILLER_35_115 ();
 sg13g2_fill_2 FILLER_35_124 ();
 sg13g2_fill_1 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_134 ();
 sg13g2_fill_1 FILLER_35_141 ();
 sg13g2_decap_4 FILLER_35_146 ();
 sg13g2_decap_4 FILLER_35_214 ();
 sg13g2_fill_1 FILLER_35_252 ();
 sg13g2_fill_1 FILLER_35_279 ();
 sg13g2_fill_1 FILLER_35_330 ();
 sg13g2_fill_2 FILLER_35_345 ();
 sg13g2_fill_1 FILLER_35_347 ();
 sg13g2_fill_2 FILLER_35_377 ();
 sg13g2_fill_1 FILLER_35_379 ();
 sg13g2_fill_1 FILLER_35_388 ();
 sg13g2_fill_2 FILLER_35_394 ();
 sg13g2_fill_1 FILLER_35_396 ();
 sg13g2_fill_2 FILLER_35_557 ();
 sg13g2_fill_1 FILLER_35_559 ();
 sg13g2_decap_8 FILLER_35_566 ();
 sg13g2_fill_1 FILLER_35_573 ();
 sg13g2_fill_1 FILLER_35_583 ();
 sg13g2_fill_2 FILLER_35_588 ();
 sg13g2_fill_1 FILLER_35_590 ();
 sg13g2_fill_1 FILLER_35_595 ();
 sg13g2_decap_8 FILLER_35_600 ();
 sg13g2_decap_8 FILLER_35_607 ();
 sg13g2_decap_8 FILLER_35_614 ();
 sg13g2_fill_2 FILLER_35_621 ();
 sg13g2_fill_1 FILLER_35_623 ();
 sg13g2_decap_4 FILLER_35_634 ();
 sg13g2_fill_2 FILLER_35_638 ();
 sg13g2_fill_2 FILLER_35_644 ();
 sg13g2_fill_1 FILLER_35_660 ();
 sg13g2_fill_1 FILLER_35_709 ();
 sg13g2_fill_2 FILLER_35_772 ();
 sg13g2_fill_1 FILLER_35_774 ();
 sg13g2_fill_1 FILLER_35_832 ();
 sg13g2_fill_1 FILLER_36_109 ();
 sg13g2_fill_1 FILLER_36_132 ();
 sg13g2_fill_1 FILLER_36_137 ();
 sg13g2_decap_4 FILLER_36_152 ();
 sg13g2_decap_4 FILLER_36_161 ();
 sg13g2_fill_2 FILLER_36_165 ();
 sg13g2_fill_2 FILLER_36_181 ();
 sg13g2_fill_1 FILLER_36_192 ();
 sg13g2_decap_4 FILLER_36_254 ();
 sg13g2_fill_2 FILLER_36_291 ();
 sg13g2_fill_1 FILLER_36_293 ();
 sg13g2_fill_1 FILLER_36_311 ();
 sg13g2_fill_2 FILLER_36_399 ();
 sg13g2_fill_1 FILLER_36_401 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_432 ();
 sg13g2_decap_8 FILLER_36_518 ();
 sg13g2_fill_2 FILLER_36_525 ();
 sg13g2_fill_1 FILLER_36_544 ();
 sg13g2_fill_2 FILLER_36_558 ();
 sg13g2_decap_4 FILLER_36_569 ();
 sg13g2_fill_1 FILLER_36_599 ();
 sg13g2_fill_1 FILLER_36_608 ();
 sg13g2_fill_2 FILLER_36_626 ();
 sg13g2_fill_1 FILLER_36_628 ();
 sg13g2_fill_1 FILLER_36_655 ();
 sg13g2_decap_4 FILLER_36_661 ();
 sg13g2_decap_8 FILLER_36_673 ();
 sg13g2_fill_2 FILLER_36_689 ();
 sg13g2_fill_2 FILLER_36_766 ();
 sg13g2_fill_1 FILLER_36_768 ();
 sg13g2_fill_2 FILLER_36_785 ();
 sg13g2_fill_2 FILLER_36_850 ();
 sg13g2_fill_1 FILLER_36_852 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_2 ();
 sg13g2_decap_8 FILLER_37_38 ();
 sg13g2_fill_1 FILLER_37_45 ();
 sg13g2_fill_2 FILLER_37_85 ();
 sg13g2_fill_1 FILLER_37_87 ();
 sg13g2_decap_8 FILLER_37_97 ();
 sg13g2_fill_1 FILLER_37_104 ();
 sg13g2_fill_2 FILLER_37_109 ();
 sg13g2_fill_2 FILLER_37_126 ();
 sg13g2_fill_2 FILLER_37_133 ();
 sg13g2_fill_1 FILLER_37_145 ();
 sg13g2_decap_4 FILLER_37_202 ();
 sg13g2_decap_4 FILLER_37_245 ();
 sg13g2_fill_2 FILLER_37_249 ();
 sg13g2_fill_2 FILLER_37_295 ();
 sg13g2_fill_1 FILLER_37_297 ();
 sg13g2_fill_1 FILLER_37_364 ();
 sg13g2_fill_2 FILLER_37_400 ();
 sg13g2_fill_1 FILLER_37_444 ();
 sg13g2_fill_1 FILLER_37_462 ();
 sg13g2_fill_2 FILLER_37_508 ();
 sg13g2_fill_1 FILLER_37_591 ();
 sg13g2_decap_4 FILLER_37_618 ();
 sg13g2_decap_4 FILLER_37_648 ();
 sg13g2_fill_1 FILLER_37_652 ();
 sg13g2_fill_2 FILLER_37_662 ();
 sg13g2_fill_1 FILLER_37_664 ();
 sg13g2_decap_4 FILLER_37_691 ();
 sg13g2_fill_1 FILLER_37_695 ();
 sg13g2_fill_2 FILLER_37_811 ();
 sg13g2_fill_2 FILLER_37_859 ();
 sg13g2_fill_1 FILLER_37_861 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_4 FILLER_38_7 ();
 sg13g2_decap_4 FILLER_38_29 ();
 sg13g2_fill_2 FILLER_38_38 ();
 sg13g2_fill_1 FILLER_38_44 ();
 sg13g2_fill_2 FILLER_38_49 ();
 sg13g2_fill_1 FILLER_38_60 ();
 sg13g2_fill_2 FILLER_38_65 ();
 sg13g2_fill_2 FILLER_38_76 ();
 sg13g2_fill_2 FILLER_38_83 ();
 sg13g2_fill_1 FILLER_38_85 ();
 sg13g2_decap_8 FILLER_38_96 ();
 sg13g2_fill_1 FILLER_38_103 ();
 sg13g2_fill_2 FILLER_38_112 ();
 sg13g2_fill_1 FILLER_38_114 ();
 sg13g2_fill_2 FILLER_38_146 ();
 sg13g2_fill_1 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_168 ();
 sg13g2_fill_2 FILLER_38_185 ();
 sg13g2_decap_8 FILLER_38_195 ();
 sg13g2_fill_2 FILLER_38_202 ();
 sg13g2_fill_1 FILLER_38_204 ();
 sg13g2_fill_1 FILLER_38_215 ();
 sg13g2_fill_2 FILLER_38_294 ();
 sg13g2_fill_2 FILLER_38_306 ();
 sg13g2_fill_2 FILLER_38_466 ();
 sg13g2_fill_2 FILLER_38_477 ();
 sg13g2_fill_1 FILLER_38_479 ();
 sg13g2_fill_1 FILLER_38_489 ();
 sg13g2_fill_2 FILLER_38_499 ();
 sg13g2_fill_1 FILLER_38_501 ();
 sg13g2_decap_8 FILLER_38_510 ();
 sg13g2_decap_4 FILLER_38_517 ();
 sg13g2_decap_4 FILLER_38_525 ();
 sg13g2_fill_1 FILLER_38_529 ();
 sg13g2_decap_8 FILLER_38_554 ();
 sg13g2_fill_1 FILLER_38_561 ();
 sg13g2_decap_8 FILLER_38_575 ();
 sg13g2_decap_8 FILLER_38_582 ();
 sg13g2_fill_2 FILLER_38_589 ();
 sg13g2_fill_2 FILLER_38_596 ();
 sg13g2_decap_4 FILLER_38_616 ();
 sg13g2_fill_2 FILLER_38_620 ();
 sg13g2_fill_1 FILLER_38_627 ();
 sg13g2_fill_2 FILLER_38_642 ();
 sg13g2_fill_2 FILLER_38_660 ();
 sg13g2_fill_1 FILLER_38_662 ();
 sg13g2_decap_4 FILLER_38_684 ();
 sg13g2_fill_1 FILLER_38_735 ();
 sg13g2_decap_8 FILLER_38_793 ();
 sg13g2_decap_8 FILLER_38_800 ();
 sg13g2_fill_1 FILLER_38_807 ();
 sg13g2_fill_2 FILLER_38_834 ();
 sg13g2_fill_2 FILLER_39_66 ();
 sg13g2_fill_1 FILLER_39_68 ();
 sg13g2_fill_2 FILLER_39_109 ();
 sg13g2_decap_8 FILLER_39_121 ();
 sg13g2_fill_2 FILLER_39_158 ();
 sg13g2_fill_1 FILLER_39_196 ();
 sg13g2_fill_1 FILLER_39_214 ();
 sg13g2_decap_8 FILLER_39_225 ();
 sg13g2_fill_1 FILLER_39_232 ();
 sg13g2_fill_2 FILLER_39_246 ();
 sg13g2_fill_1 FILLER_39_248 ();
 sg13g2_fill_2 FILLER_39_266 ();
 sg13g2_fill_1 FILLER_39_344 ();
 sg13g2_fill_2 FILLER_39_374 ();
 sg13g2_fill_2 FILLER_39_406 ();
 sg13g2_fill_1 FILLER_39_422 ();
 sg13g2_fill_2 FILLER_39_453 ();
 sg13g2_fill_1 FILLER_39_469 ();
 sg13g2_decap_8 FILLER_39_519 ();
 sg13g2_decap_8 FILLER_39_526 ();
 sg13g2_fill_2 FILLER_39_533 ();
 sg13g2_fill_1 FILLER_39_562 ();
 sg13g2_decap_4 FILLER_39_569 ();
 sg13g2_fill_2 FILLER_39_587 ();
 sg13g2_fill_2 FILLER_39_644 ();
 sg13g2_fill_1 FILLER_39_646 ();
 sg13g2_decap_4 FILLER_39_663 ();
 sg13g2_fill_1 FILLER_39_741 ();
 sg13g2_fill_2 FILLER_39_753 ();
 sg13g2_decap_4 FILLER_39_767 ();
 sg13g2_decap_4 FILLER_39_797 ();
 sg13g2_decap_4 FILLER_39_814 ();
 sg13g2_fill_2 FILLER_39_818 ();
 sg13g2_decap_4 FILLER_40_0 ();
 sg13g2_decap_4 FILLER_40_42 ();
 sg13g2_fill_2 FILLER_40_46 ();
 sg13g2_fill_2 FILLER_40_57 ();
 sg13g2_fill_2 FILLER_40_97 ();
 sg13g2_fill_1 FILLER_40_99 ();
 sg13g2_fill_1 FILLER_40_122 ();
 sg13g2_fill_1 FILLER_40_131 ();
 sg13g2_fill_1 FILLER_40_154 ();
 sg13g2_fill_1 FILLER_40_196 ();
 sg13g2_fill_2 FILLER_40_236 ();
 sg13g2_fill_1 FILLER_40_238 ();
 sg13g2_fill_2 FILLER_40_303 ();
 sg13g2_fill_2 FILLER_40_313 ();
 sg13g2_fill_1 FILLER_40_385 ();
 sg13g2_fill_1 FILLER_40_468 ();
 sg13g2_fill_2 FILLER_40_492 ();
 sg13g2_fill_1 FILLER_40_510 ();
 sg13g2_decap_4 FILLER_40_537 ();
 sg13g2_fill_1 FILLER_40_541 ();
 sg13g2_decap_8 FILLER_40_550 ();
 sg13g2_fill_2 FILLER_40_557 ();
 sg13g2_fill_2 FILLER_40_567 ();
 sg13g2_fill_1 FILLER_40_569 ();
 sg13g2_decap_8 FILLER_40_574 ();
 sg13g2_decap_8 FILLER_40_581 ();
 sg13g2_fill_2 FILLER_40_605 ();
 sg13g2_decap_4 FILLER_40_613 ();
 sg13g2_fill_1 FILLER_40_617 ();
 sg13g2_fill_1 FILLER_40_638 ();
 sg13g2_decap_4 FILLER_40_653 ();
 sg13g2_decap_8 FILLER_40_670 ();
 sg13g2_fill_2 FILLER_40_677 ();
 sg13g2_decap_8 FILLER_40_711 ();
 sg13g2_decap_4 FILLER_40_718 ();
 sg13g2_fill_1 FILLER_40_739 ();
 sg13g2_fill_2 FILLER_40_749 ();
 sg13g2_fill_2 FILLER_40_764 ();
 sg13g2_fill_1 FILLER_40_766 ();
 sg13g2_fill_2 FILLER_40_790 ();
 sg13g2_fill_1 FILLER_40_792 ();
 sg13g2_fill_2 FILLER_40_824 ();
 sg13g2_fill_2 FILLER_40_830 ();
 sg13g2_decap_8 FILLER_41_26 ();
 sg13g2_fill_1 FILLER_41_33 ();
 sg13g2_decap_4 FILLER_41_74 ();
 sg13g2_fill_2 FILLER_41_78 ();
 sg13g2_fill_2 FILLER_41_98 ();
 sg13g2_fill_1 FILLER_41_100 ();
 sg13g2_fill_1 FILLER_41_144 ();
 sg13g2_fill_1 FILLER_41_158 ();
 sg13g2_fill_1 FILLER_41_194 ();
 sg13g2_fill_2 FILLER_41_205 ();
 sg13g2_fill_1 FILLER_41_246 ();
 sg13g2_fill_1 FILLER_41_252 ();
 sg13g2_fill_1 FILLER_41_312 ();
 sg13g2_fill_2 FILLER_41_327 ();
 sg13g2_fill_1 FILLER_41_341 ();
 sg13g2_fill_2 FILLER_41_379 ();
 sg13g2_fill_2 FILLER_41_407 ();
 sg13g2_fill_1 FILLER_41_409 ();
 sg13g2_fill_2 FILLER_41_424 ();
 sg13g2_fill_1 FILLER_41_426 ();
 sg13g2_fill_2 FILLER_41_441 ();
 sg13g2_fill_2 FILLER_41_461 ();
 sg13g2_fill_1 FILLER_41_495 ();
 sg13g2_decap_4 FILLER_41_512 ();
 sg13g2_fill_1 FILLER_41_516 ();
 sg13g2_decap_8 FILLER_41_526 ();
 sg13g2_decap_8 FILLER_41_533 ();
 sg13g2_fill_2 FILLER_41_540 ();
 sg13g2_fill_1 FILLER_41_570 ();
 sg13g2_fill_1 FILLER_41_587 ();
 sg13g2_fill_1 FILLER_41_596 ();
 sg13g2_decap_4 FILLER_41_626 ();
 sg13g2_fill_1 FILLER_41_630 ();
 sg13g2_fill_1 FILLER_41_640 ();
 sg13g2_decap_4 FILLER_41_661 ();
 sg13g2_fill_1 FILLER_41_665 ();
 sg13g2_fill_2 FILLER_41_692 ();
 sg13g2_fill_1 FILLER_41_731 ();
 sg13g2_fill_1 FILLER_41_801 ();
 sg13g2_decap_8 FILLER_41_818 ();
 sg13g2_fill_2 FILLER_41_825 ();
 sg13g2_fill_1 FILLER_41_827 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_7 ();
 sg13g2_fill_1 FILLER_42_9 ();
 sg13g2_fill_2 FILLER_42_33 ();
 sg13g2_fill_1 FILLER_42_35 ();
 sg13g2_decap_4 FILLER_42_50 ();
 sg13g2_fill_1 FILLER_42_54 ();
 sg13g2_fill_2 FILLER_42_100 ();
 sg13g2_fill_1 FILLER_42_102 ();
 sg13g2_decap_8 FILLER_42_122 ();
 sg13g2_fill_2 FILLER_42_223 ();
 sg13g2_fill_1 FILLER_42_251 ();
 sg13g2_fill_1 FILLER_42_296 ();
 sg13g2_fill_1 FILLER_42_304 ();
 sg13g2_fill_2 FILLER_42_352 ();
 sg13g2_fill_1 FILLER_42_378 ();
 sg13g2_fill_2 FILLER_42_388 ();
 sg13g2_fill_1 FILLER_42_390 ();
 sg13g2_fill_1 FILLER_42_433 ();
 sg13g2_fill_1 FILLER_42_472 ();
 sg13g2_fill_1 FILLER_42_507 ();
 sg13g2_fill_2 FILLER_42_534 ();
 sg13g2_fill_2 FILLER_42_556 ();
 sg13g2_fill_1 FILLER_42_558 ();
 sg13g2_fill_2 FILLER_42_573 ();
 sg13g2_fill_2 FILLER_42_588 ();
 sg13g2_fill_2 FILLER_42_602 ();
 sg13g2_fill_1 FILLER_42_625 ();
 sg13g2_decap_8 FILLER_42_642 ();
 sg13g2_fill_2 FILLER_42_649 ();
 sg13g2_decap_8 FILLER_42_668 ();
 sg13g2_fill_2 FILLER_42_675 ();
 sg13g2_decap_4 FILLER_42_703 ();
 sg13g2_fill_1 FILLER_42_707 ();
 sg13g2_fill_2 FILLER_42_716 ();
 sg13g2_decap_8 FILLER_42_743 ();
 sg13g2_decap_4 FILLER_42_750 ();
 sg13g2_fill_1 FILLER_42_754 ();
 sg13g2_fill_2 FILLER_42_767 ();
 sg13g2_decap_4 FILLER_42_773 ();
 sg13g2_fill_2 FILLER_42_777 ();
 sg13g2_fill_2 FILLER_42_804 ();
 sg13g2_fill_1 FILLER_42_810 ();
 sg13g2_decap_8 FILLER_42_828 ();
 sg13g2_decap_8 FILLER_42_835 ();
 sg13g2_decap_4 FILLER_42_842 ();
 sg13g2_fill_2 FILLER_42_846 ();
 sg13g2_fill_1 FILLER_42_861 ();
 sg13g2_decap_8 FILLER_43_26 ();
 sg13g2_fill_2 FILLER_43_72 ();
 sg13g2_decap_4 FILLER_43_84 ();
 sg13g2_fill_2 FILLER_43_88 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_4 FILLER_43_133 ();
 sg13g2_fill_2 FILLER_43_167 ();
 sg13g2_fill_2 FILLER_43_250 ();
 sg13g2_fill_1 FILLER_43_252 ();
 sg13g2_fill_2 FILLER_43_262 ();
 sg13g2_fill_1 FILLER_43_264 ();
 sg13g2_fill_2 FILLER_43_273 ();
 sg13g2_fill_1 FILLER_43_275 ();
 sg13g2_fill_1 FILLER_43_312 ();
 sg13g2_fill_2 FILLER_43_334 ();
 sg13g2_fill_2 FILLER_43_420 ();
 sg13g2_fill_1 FILLER_43_443 ();
 sg13g2_fill_2 FILLER_43_484 ();
 sg13g2_decap_8 FILLER_43_512 ();
 sg13g2_fill_1 FILLER_43_519 ();
 sg13g2_decap_8 FILLER_43_529 ();
 sg13g2_decap_8 FILLER_43_536 ();
 sg13g2_fill_2 FILLER_43_573 ();
 sg13g2_fill_1 FILLER_43_575 ();
 sg13g2_decap_4 FILLER_43_614 ();
 sg13g2_fill_1 FILLER_43_627 ();
 sg13g2_fill_1 FILLER_43_650 ();
 sg13g2_decap_8 FILLER_43_672 ();
 sg13g2_decap_8 FILLER_43_679 ();
 sg13g2_decap_8 FILLER_43_686 ();
 sg13g2_decap_4 FILLER_43_693 ();
 sg13g2_fill_2 FILLER_43_720 ();
 sg13g2_fill_1 FILLER_43_722 ();
 sg13g2_fill_2 FILLER_43_799 ();
 sg13g2_fill_2 FILLER_43_827 ();
 sg13g2_fill_1 FILLER_43_829 ();
 sg13g2_fill_1 FILLER_43_856 ();
 sg13g2_fill_1 FILLER_43_861 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_4 FILLER_44_7 ();
 sg13g2_decap_4 FILLER_44_15 ();
 sg13g2_fill_1 FILLER_44_19 ();
 sg13g2_fill_2 FILLER_44_30 ();
 sg13g2_decap_4 FILLER_44_57 ();
 sg13g2_fill_1 FILLER_44_61 ();
 sg13g2_decap_8 FILLER_44_97 ();
 sg13g2_decap_8 FILLER_44_104 ();
 sg13g2_fill_1 FILLER_44_165 ();
 sg13g2_fill_1 FILLER_44_255 ();
 sg13g2_fill_2 FILLER_44_271 ();
 sg13g2_fill_1 FILLER_44_273 ();
 sg13g2_fill_1 FILLER_44_309 ();
 sg13g2_fill_1 FILLER_44_333 ();
 sg13g2_fill_2 FILLER_44_380 ();
 sg13g2_fill_2 FILLER_44_396 ();
 sg13g2_fill_1 FILLER_44_473 ();
 sg13g2_fill_1 FILLER_44_500 ();
 sg13g2_fill_2 FILLER_44_518 ();
 sg13g2_fill_1 FILLER_44_520 ();
 sg13g2_decap_8 FILLER_44_525 ();
 sg13g2_decap_8 FILLER_44_532 ();
 sg13g2_fill_2 FILLER_44_539 ();
 sg13g2_fill_2 FILLER_44_550 ();
 sg13g2_decap_8 FILLER_44_583 ();
 sg13g2_fill_1 FILLER_44_609 ();
 sg13g2_decap_4 FILLER_44_615 ();
 sg13g2_fill_1 FILLER_44_619 ();
 sg13g2_fill_1 FILLER_44_625 ();
 sg13g2_fill_2 FILLER_44_645 ();
 sg13g2_fill_1 FILLER_44_647 ();
 sg13g2_decap_8 FILLER_44_664 ();
 sg13g2_decap_8 FILLER_44_671 ();
 sg13g2_decap_8 FILLER_44_678 ();
 sg13g2_decap_8 FILLER_44_689 ();
 sg13g2_fill_2 FILLER_44_696 ();
 sg13g2_fill_1 FILLER_44_698 ();
 sg13g2_fill_1 FILLER_44_709 ();
 sg13g2_decap_8 FILLER_44_727 ();
 sg13g2_decap_4 FILLER_44_734 ();
 sg13g2_fill_2 FILLER_44_738 ();
 sg13g2_decap_4 FILLER_44_752 ();
 sg13g2_fill_2 FILLER_44_766 ();
 sg13g2_fill_1 FILLER_44_794 ();
 sg13g2_fill_1 FILLER_44_816 ();
 sg13g2_decap_8 FILLER_44_830 ();
 sg13g2_decap_4 FILLER_44_837 ();
 sg13g2_fill_1 FILLER_44_861 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_58 ();
 sg13g2_decap_4 FILLER_45_65 ();
 sg13g2_fill_2 FILLER_45_69 ();
 sg13g2_decap_4 FILLER_45_116 ();
 sg13g2_fill_2 FILLER_45_120 ();
 sg13g2_fill_2 FILLER_45_126 ();
 sg13g2_fill_1 FILLER_45_128 ();
 sg13g2_fill_1 FILLER_45_173 ();
 sg13g2_fill_1 FILLER_45_183 ();
 sg13g2_fill_1 FILLER_45_214 ();
 sg13g2_fill_2 FILLER_45_255 ();
 sg13g2_fill_2 FILLER_45_266 ();
 sg13g2_fill_1 FILLER_45_268 ();
 sg13g2_fill_2 FILLER_45_295 ();
 sg13g2_fill_1 FILLER_45_297 ();
 sg13g2_fill_1 FILLER_45_331 ();
 sg13g2_fill_1 FILLER_45_403 ();
 sg13g2_fill_1 FILLER_45_445 ();
 sg13g2_fill_2 FILLER_45_468 ();
 sg13g2_fill_1 FILLER_45_475 ();
 sg13g2_fill_2 FILLER_45_508 ();
 sg13g2_fill_2 FILLER_45_536 ();
 sg13g2_fill_1 FILLER_45_538 ();
 sg13g2_fill_1 FILLER_45_549 ();
 sg13g2_decap_8 FILLER_45_559 ();
 sg13g2_fill_2 FILLER_45_566 ();
 sg13g2_fill_2 FILLER_45_591 ();
 sg13g2_fill_2 FILLER_45_597 ();
 sg13g2_fill_1 FILLER_45_603 ();
 sg13g2_fill_1 FILLER_45_619 ();
 sg13g2_fill_2 FILLER_45_638 ();
 sg13g2_fill_1 FILLER_45_640 ();
 sg13g2_decap_4 FILLER_45_669 ();
 sg13g2_fill_2 FILLER_45_673 ();
 sg13g2_decap_8 FILLER_45_723 ();
 sg13g2_fill_2 FILLER_45_730 ();
 sg13g2_fill_1 FILLER_45_732 ();
 sg13g2_fill_2 FILLER_45_741 ();
 sg13g2_fill_2 FILLER_45_751 ();
 sg13g2_fill_1 FILLER_45_753 ();
 sg13g2_decap_4 FILLER_45_780 ();
 sg13g2_fill_2 FILLER_45_784 ();
 sg13g2_fill_1 FILLER_45_861 ();
 sg13g2_fill_1 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_19 ();
 sg13g2_fill_1 FILLER_46_21 ();
 sg13g2_fill_1 FILLER_46_27 ();
 sg13g2_fill_1 FILLER_46_56 ();
 sg13g2_fill_2 FILLER_46_109 ();
 sg13g2_fill_1 FILLER_46_140 ();
 sg13g2_fill_1 FILLER_46_177 ();
 sg13g2_fill_2 FILLER_46_348 ();
 sg13g2_fill_2 FILLER_46_395 ();
 sg13g2_fill_1 FILLER_46_397 ();
 sg13g2_fill_1 FILLER_46_433 ();
 sg13g2_fill_2 FILLER_46_465 ();
 sg13g2_fill_1 FILLER_46_493 ();
 sg13g2_decap_8 FILLER_46_527 ();
 sg13g2_fill_2 FILLER_46_534 ();
 sg13g2_fill_1 FILLER_46_536 ();
 sg13g2_fill_1 FILLER_46_566 ();
 sg13g2_fill_2 FILLER_46_586 ();
 sg13g2_fill_2 FILLER_46_597 ();
 sg13g2_fill_1 FILLER_46_599 ();
 sg13g2_fill_1 FILLER_46_625 ();
 sg13g2_fill_1 FILLER_46_644 ();
 sg13g2_fill_2 FILLER_46_663 ();
 sg13g2_decap_8 FILLER_46_669 ();
 sg13g2_fill_2 FILLER_46_761 ();
 sg13g2_fill_2 FILLER_46_768 ();
 sg13g2_decap_8 FILLER_46_775 ();
 sg13g2_fill_2 FILLER_46_782 ();
 sg13g2_fill_1 FILLER_46_784 ();
 sg13g2_decap_8 FILLER_46_792 ();
 sg13g2_decap_4 FILLER_46_799 ();
 sg13g2_decap_4 FILLER_46_808 ();
 sg13g2_fill_2 FILLER_46_812 ();
 sg13g2_fill_2 FILLER_46_838 ();
 sg13g2_fill_2 FILLER_46_845 ();
 sg13g2_decap_8 FILLER_46_855 ();
 sg13g2_fill_2 FILLER_47_34 ();
 sg13g2_fill_2 FILLER_47_53 ();
 sg13g2_fill_1 FILLER_47_55 ();
 sg13g2_fill_2 FILLER_47_65 ();
 sg13g2_fill_1 FILLER_47_89 ();
 sg13g2_fill_1 FILLER_47_95 ();
 sg13g2_fill_1 FILLER_47_130 ();
 sg13g2_fill_2 FILLER_47_157 ();
 sg13g2_fill_1 FILLER_47_185 ();
 sg13g2_fill_1 FILLER_47_212 ();
 sg13g2_fill_2 FILLER_47_262 ();
 sg13g2_fill_1 FILLER_47_273 ();
 sg13g2_fill_2 FILLER_47_288 ();
 sg13g2_fill_2 FILLER_47_306 ();
 sg13g2_fill_2 FILLER_47_341 ();
 sg13g2_fill_1 FILLER_47_369 ();
 sg13g2_fill_2 FILLER_47_421 ();
 sg13g2_fill_2 FILLER_47_462 ();
 sg13g2_fill_2 FILLER_47_493 ();
 sg13g2_fill_2 FILLER_47_511 ();
 sg13g2_fill_1 FILLER_47_531 ();
 sg13g2_decap_8 FILLER_47_536 ();
 sg13g2_fill_2 FILLER_47_543 ();
 sg13g2_decap_8 FILLER_47_565 ();
 sg13g2_decap_4 FILLER_47_572 ();
 sg13g2_fill_2 FILLER_47_576 ();
 sg13g2_decap_4 FILLER_47_603 ();
 sg13g2_decap_4 FILLER_47_611 ();
 sg13g2_fill_1 FILLER_47_615 ();
 sg13g2_decap_8 FILLER_47_637 ();
 sg13g2_fill_2 FILLER_47_644 ();
 sg13g2_fill_2 FILLER_47_651 ();
 sg13g2_fill_2 FILLER_47_658 ();
 sg13g2_fill_1 FILLER_47_664 ();
 sg13g2_decap_4 FILLER_47_691 ();
 sg13g2_fill_1 FILLER_47_695 ();
 sg13g2_decap_8 FILLER_47_709 ();
 sg13g2_decap_8 FILLER_47_716 ();
 sg13g2_decap_8 FILLER_47_723 ();
 sg13g2_decap_8 FILLER_47_730 ();
 sg13g2_fill_2 FILLER_47_776 ();
 sg13g2_fill_1 FILLER_47_778 ();
 sg13g2_decap_8 FILLER_47_802 ();
 sg13g2_fill_2 FILLER_47_809 ();
 sg13g2_fill_2 FILLER_47_837 ();
 sg13g2_fill_2 FILLER_47_860 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_4 FILLER_48_30 ();
 sg13g2_fill_2 FILLER_48_50 ();
 sg13g2_fill_1 FILLER_48_52 ();
 sg13g2_fill_2 FILLER_48_58 ();
 sg13g2_fill_1 FILLER_48_153 ();
 sg13g2_fill_1 FILLER_48_167 ();
 sg13g2_fill_2 FILLER_48_315 ();
 sg13g2_fill_2 FILLER_48_333 ();
 sg13g2_fill_2 FILLER_48_367 ();
 sg13g2_fill_2 FILLER_48_443 ();
 sg13g2_fill_2 FILLER_48_460 ();
 sg13g2_fill_1 FILLER_48_467 ();
 sg13g2_fill_1 FILLER_48_496 ();
 sg13g2_fill_2 FILLER_48_509 ();
 sg13g2_fill_1 FILLER_48_511 ();
 sg13g2_fill_2 FILLER_48_577 ();
 sg13g2_fill_1 FILLER_48_583 ();
 sg13g2_fill_2 FILLER_48_615 ();
 sg13g2_decap_8 FILLER_48_635 ();
 sg13g2_fill_1 FILLER_48_642 ();
 sg13g2_decap_4 FILLER_48_651 ();
 sg13g2_fill_1 FILLER_48_655 ();
 sg13g2_fill_2 FILLER_48_690 ();
 sg13g2_fill_1 FILLER_48_692 ();
 sg13g2_fill_2 FILLER_48_706 ();
 sg13g2_decap_4 FILLER_48_763 ();
 sg13g2_fill_2 FILLER_48_767 ();
 sg13g2_decap_8 FILLER_48_773 ();
 sg13g2_fill_2 FILLER_48_780 ();
 sg13g2_fill_2 FILLER_48_787 ();
 sg13g2_fill_2 FILLER_48_805 ();
 sg13g2_fill_1 FILLER_48_828 ();
 sg13g2_decap_8 FILLER_48_855 ();
 sg13g2_fill_2 FILLER_49_45 ();
 sg13g2_decap_8 FILLER_49_51 ();
 sg13g2_fill_1 FILLER_49_77 ();
 sg13g2_fill_1 FILLER_49_91 ();
 sg13g2_fill_2 FILLER_49_127 ();
 sg13g2_fill_1 FILLER_49_164 ();
 sg13g2_fill_1 FILLER_49_196 ();
 sg13g2_fill_2 FILLER_49_206 ();
 sg13g2_fill_1 FILLER_49_315 ();
 sg13g2_fill_2 FILLER_49_338 ();
 sg13g2_fill_1 FILLER_49_340 ();
 sg13g2_fill_1 FILLER_49_355 ();
 sg13g2_fill_1 FILLER_49_383 ();
 sg13g2_fill_2 FILLER_49_406 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_fill_2 FILLER_49_488 ();
 sg13g2_fill_1 FILLER_49_490 ();
 sg13g2_fill_1 FILLER_49_501 ();
 sg13g2_fill_1 FILLER_49_531 ();
 sg13g2_decap_8 FILLER_49_567 ();
 sg13g2_fill_1 FILLER_49_574 ();
 sg13g2_decap_4 FILLER_49_611 ();
 sg13g2_fill_1 FILLER_49_623 ();
 sg13g2_decap_4 FILLER_49_658 ();
 sg13g2_decap_8 FILLER_49_678 ();
 sg13g2_fill_1 FILLER_49_685 ();
 sg13g2_decap_8 FILLER_49_715 ();
 sg13g2_decap_8 FILLER_49_722 ();
 sg13g2_decap_4 FILLER_49_760 ();
 sg13g2_decap_8 FILLER_49_773 ();
 sg13g2_decap_8 FILLER_49_780 ();
 sg13g2_fill_2 FILLER_49_805 ();
 sg13g2_fill_1 FILLER_49_807 ();
 sg13g2_fill_2 FILLER_49_822 ();
 sg13g2_fill_1 FILLER_49_824 ();
 sg13g2_decap_8 FILLER_49_851 ();
 sg13g2_decap_4 FILLER_49_858 ();
 sg13g2_decap_4 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_4 ();
 sg13g2_fill_2 FILLER_50_71 ();
 sg13g2_fill_2 FILLER_50_104 ();
 sg13g2_fill_1 FILLER_50_144 ();
 sg13g2_fill_2 FILLER_50_154 ();
 sg13g2_fill_1 FILLER_50_229 ();
 sg13g2_decap_8 FILLER_50_233 ();
 sg13g2_fill_2 FILLER_50_240 ();
 sg13g2_fill_1 FILLER_50_314 ();
 sg13g2_fill_1 FILLER_50_338 ();
 sg13g2_fill_2 FILLER_50_347 ();
 sg13g2_fill_1 FILLER_50_375 ();
 sg13g2_fill_1 FILLER_50_491 ();
 sg13g2_fill_1 FILLER_50_499 ();
 sg13g2_fill_1 FILLER_50_577 ();
 sg13g2_decap_8 FILLER_50_613 ();
 sg13g2_fill_1 FILLER_50_620 ();
 sg13g2_fill_1 FILLER_50_626 ();
 sg13g2_decap_8 FILLER_50_634 ();
 sg13g2_decap_8 FILLER_50_641 ();
 sg13g2_decap_8 FILLER_50_648 ();
 sg13g2_decap_8 FILLER_50_655 ();
 sg13g2_fill_2 FILLER_50_662 ();
 sg13g2_fill_1 FILLER_50_664 ();
 sg13g2_decap_8 FILLER_50_683 ();
 sg13g2_decap_4 FILLER_50_690 ();
 sg13g2_fill_2 FILLER_50_694 ();
 sg13g2_decap_8 FILLER_50_711 ();
 sg13g2_decap_8 FILLER_50_718 ();
 sg13g2_decap_8 FILLER_50_835 ();
 sg13g2_decap_8 FILLER_50_842 ();
 sg13g2_decap_8 FILLER_50_849 ();
 sg13g2_decap_4 FILLER_50_856 ();
 sg13g2_fill_2 FILLER_50_860 ();
 sg13g2_fill_1 FILLER_51_38 ();
 sg13g2_fill_1 FILLER_51_53 ();
 sg13g2_fill_1 FILLER_51_91 ();
 sg13g2_fill_2 FILLER_51_116 ();
 sg13g2_fill_2 FILLER_51_175 ();
 sg13g2_fill_2 FILLER_51_211 ();
 sg13g2_decap_8 FILLER_51_239 ();
 sg13g2_fill_1 FILLER_51_246 ();
 sg13g2_fill_1 FILLER_51_265 ();
 sg13g2_fill_2 FILLER_51_289 ();
 sg13g2_fill_2 FILLER_51_340 ();
 sg13g2_fill_2 FILLER_51_355 ();
 sg13g2_fill_1 FILLER_51_357 ();
 sg13g2_fill_2 FILLER_51_364 ();
 sg13g2_fill_1 FILLER_51_366 ();
 sg13g2_fill_1 FILLER_51_410 ();
 sg13g2_decap_8 FILLER_51_599 ();
 sg13g2_decap_8 FILLER_51_606 ();
 sg13g2_decap_4 FILLER_51_613 ();
 sg13g2_decap_4 FILLER_51_656 ();
 sg13g2_fill_1 FILLER_51_729 ();
 sg13g2_fill_2 FILLER_51_754 ();
 sg13g2_fill_1 FILLER_51_756 ();
 sg13g2_decap_8 FILLER_51_776 ();
 sg13g2_decap_8 FILLER_51_783 ();
 sg13g2_decap_8 FILLER_51_803 ();
 sg13g2_decap_8 FILLER_51_810 ();
 sg13g2_decap_8 FILLER_51_817 ();
 sg13g2_decap_8 FILLER_51_824 ();
 sg13g2_decap_8 FILLER_51_831 ();
 sg13g2_decap_8 FILLER_51_838 ();
 sg13g2_decap_8 FILLER_51_845 ();
 sg13g2_decap_8 FILLER_51_852 ();
 sg13g2_fill_2 FILLER_51_859 ();
 sg13g2_fill_1 FILLER_51_861 ();
 sg13g2_fill_1 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_32 ();
 sg13g2_fill_1 FILLER_52_40 ();
 sg13g2_fill_2 FILLER_52_48 ();
 sg13g2_fill_1 FILLER_52_56 ();
 sg13g2_fill_2 FILLER_52_71 ();
 sg13g2_fill_2 FILLER_52_103 ();
 sg13g2_fill_2 FILLER_52_197 ();
 sg13g2_fill_1 FILLER_52_199 ();
 sg13g2_decap_8 FILLER_52_238 ();
 sg13g2_fill_2 FILLER_52_245 ();
 sg13g2_fill_1 FILLER_52_273 ();
 sg13g2_fill_2 FILLER_52_283 ();
 sg13g2_fill_1 FILLER_52_312 ();
 sg13g2_fill_1 FILLER_52_358 ();
 sg13g2_fill_2 FILLER_52_389 ();
 sg13g2_fill_1 FILLER_52_391 ();
 sg13g2_fill_2 FILLER_52_411 ();
 sg13g2_fill_1 FILLER_52_413 ();
 sg13g2_fill_2 FILLER_52_488 ();
 sg13g2_fill_2 FILLER_52_505 ();
 sg13g2_fill_1 FILLER_52_507 ();
 sg13g2_fill_2 FILLER_52_534 ();
 sg13g2_fill_1 FILLER_52_536 ();
 sg13g2_decap_4 FILLER_52_580 ();
 sg13g2_decap_4 FILLER_52_588 ();
 sg13g2_fill_1 FILLER_52_592 ();
 sg13g2_decap_8 FILLER_52_597 ();
 sg13g2_fill_2 FILLER_52_604 ();
 sg13g2_fill_1 FILLER_52_606 ();
 sg13g2_fill_2 FILLER_52_629 ();
 sg13g2_fill_1 FILLER_52_657 ();
 sg13g2_decap_4 FILLER_52_662 ();
 sg13g2_fill_1 FILLER_52_666 ();
 sg13g2_decap_8 FILLER_52_683 ();
 sg13g2_decap_8 FILLER_52_690 ();
 sg13g2_decap_8 FILLER_52_697 ();
 sg13g2_decap_8 FILLER_52_704 ();
 sg13g2_decap_8 FILLER_52_711 ();
 sg13g2_fill_2 FILLER_52_743 ();
 sg13g2_fill_1 FILLER_52_751 ();
 sg13g2_decap_8 FILLER_52_756 ();
 sg13g2_fill_2 FILLER_52_763 ();
 sg13g2_decap_8 FILLER_52_777 ();
 sg13g2_fill_2 FILLER_52_784 ();
 sg13g2_fill_1 FILLER_52_786 ();
 sg13g2_decap_8 FILLER_52_813 ();
 sg13g2_decap_8 FILLER_52_820 ();
 sg13g2_decap_8 FILLER_52_827 ();
 sg13g2_decap_8 FILLER_52_834 ();
 sg13g2_decap_8 FILLER_52_841 ();
 sg13g2_decap_8 FILLER_52_848 ();
 sg13g2_decap_8 FILLER_52_855 ();
 sg13g2_fill_1 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_32 ();
 sg13g2_fill_1 FILLER_53_62 ();
 sg13g2_fill_2 FILLER_53_68 ();
 sg13g2_fill_1 FILLER_53_111 ();
 sg13g2_fill_2 FILLER_53_168 ();
 sg13g2_fill_1 FILLER_53_170 ();
 sg13g2_fill_2 FILLER_53_193 ();
 sg13g2_fill_1 FILLER_53_195 ();
 sg13g2_fill_1 FILLER_53_218 ();
 sg13g2_fill_1 FILLER_53_254 ();
 sg13g2_fill_2 FILLER_53_374 ();
 sg13g2_fill_1 FILLER_53_376 ();
 sg13g2_fill_2 FILLER_53_444 ();
 sg13g2_fill_1 FILLER_53_446 ();
 sg13g2_fill_2 FILLER_53_465 ();
 sg13g2_fill_2 FILLER_53_471 ();
 sg13g2_fill_2 FILLER_53_534 ();
 sg13g2_fill_1 FILLER_53_536 ();
 sg13g2_fill_2 FILLER_53_555 ();
 sg13g2_decap_4 FILLER_53_576 ();
 sg13g2_fill_2 FILLER_53_580 ();
 sg13g2_decap_8 FILLER_53_592 ();
 sg13g2_decap_8 FILLER_53_599 ();
 sg13g2_fill_1 FILLER_53_606 ();
 sg13g2_fill_1 FILLER_53_624 ();
 sg13g2_fill_1 FILLER_53_661 ();
 sg13g2_fill_1 FILLER_53_717 ();
 sg13g2_decap_8 FILLER_53_726 ();
 sg13g2_decap_8 FILLER_53_733 ();
 sg13g2_fill_2 FILLER_53_740 ();
 sg13g2_decap_8 FILLER_53_757 ();
 sg13g2_fill_2 FILLER_53_764 ();
 sg13g2_fill_1 FILLER_53_792 ();
 sg13g2_decap_8 FILLER_53_811 ();
 sg13g2_decap_8 FILLER_53_818 ();
 sg13g2_decap_8 FILLER_53_825 ();
 sg13g2_decap_8 FILLER_53_832 ();
 sg13g2_decap_8 FILLER_53_839 ();
 sg13g2_decap_8 FILLER_53_846 ();
 sg13g2_decap_8 FILLER_53_853 ();
 sg13g2_fill_2 FILLER_53_860 ();
 sg13g2_fill_2 FILLER_54_57 ();
 sg13g2_fill_1 FILLER_54_82 ();
 sg13g2_fill_2 FILLER_54_100 ();
 sg13g2_fill_1 FILLER_54_102 ();
 sg13g2_fill_1 FILLER_54_117 ();
 sg13g2_fill_1 FILLER_54_167 ();
 sg13g2_fill_2 FILLER_54_194 ();
 sg13g2_fill_1 FILLER_54_203 ();
 sg13g2_decap_4 FILLER_54_254 ();
 sg13g2_fill_1 FILLER_54_299 ();
 sg13g2_fill_2 FILLER_54_343 ();
 sg13g2_fill_1 FILLER_54_359 ();
 sg13g2_fill_2 FILLER_54_370 ();
 sg13g2_decap_8 FILLER_54_393 ();
 sg13g2_decap_4 FILLER_54_400 ();
 sg13g2_fill_2 FILLER_54_425 ();
 sg13g2_fill_1 FILLER_54_427 ();
 sg13g2_fill_2 FILLER_54_482 ();
 sg13g2_fill_2 FILLER_54_488 ();
 sg13g2_fill_2 FILLER_54_503 ();
 sg13g2_fill_2 FILLER_54_509 ();
 sg13g2_fill_1 FILLER_54_511 ();
 sg13g2_fill_2 FILLER_54_564 ();
 sg13g2_fill_1 FILLER_54_566 ();
 sg13g2_fill_2 FILLER_54_640 ();
 sg13g2_fill_2 FILLER_54_667 ();
 sg13g2_decap_4 FILLER_54_743 ();
 sg13g2_decap_8 FILLER_54_761 ();
 sg13g2_decap_4 FILLER_54_787 ();
 sg13g2_fill_1 FILLER_54_791 ();
 sg13g2_decap_8 FILLER_54_804 ();
 sg13g2_decap_8 FILLER_54_811 ();
 sg13g2_decap_8 FILLER_54_818 ();
 sg13g2_decap_8 FILLER_54_825 ();
 sg13g2_decap_8 FILLER_54_832 ();
 sg13g2_decap_8 FILLER_54_839 ();
 sg13g2_decap_8 FILLER_54_846 ();
 sg13g2_decap_8 FILLER_54_853 ();
 sg13g2_fill_2 FILLER_54_860 ();
 sg13g2_fill_2 FILLER_55_26 ();
 sg13g2_fill_2 FILLER_55_48 ();
 sg13g2_fill_1 FILLER_55_50 ();
 sg13g2_fill_2 FILLER_55_61 ();
 sg13g2_fill_2 FILLER_55_68 ();
 sg13g2_fill_1 FILLER_55_108 ();
 sg13g2_fill_1 FILLER_55_141 ();
 sg13g2_fill_1 FILLER_55_174 ();
 sg13g2_fill_2 FILLER_55_201 ();
 sg13g2_fill_1 FILLER_55_208 ();
 sg13g2_fill_1 FILLER_55_240 ();
 sg13g2_fill_2 FILLER_55_246 ();
 sg13g2_fill_2 FILLER_55_256 ();
 sg13g2_decap_4 FILLER_55_263 ();
 sg13g2_fill_2 FILLER_55_271 ();
 sg13g2_decap_4 FILLER_55_278 ();
 sg13g2_fill_1 FILLER_55_282 ();
 sg13g2_fill_2 FILLER_55_286 ();
 sg13g2_fill_1 FILLER_55_288 ();
 sg13g2_fill_1 FILLER_55_308 ();
 sg13g2_fill_2 FILLER_55_377 ();
 sg13g2_fill_1 FILLER_55_413 ();
 sg13g2_decap_8 FILLER_55_449 ();
 sg13g2_decap_8 FILLER_55_456 ();
 sg13g2_fill_2 FILLER_55_463 ();
 sg13g2_fill_1 FILLER_55_465 ();
 sg13g2_fill_2 FILLER_55_528 ();
 sg13g2_fill_1 FILLER_55_530 ();
 sg13g2_fill_2 FILLER_55_571 ();
 sg13g2_fill_2 FILLER_55_597 ();
 sg13g2_fill_1 FILLER_55_625 ();
 sg13g2_decap_4 FILLER_55_663 ();
 sg13g2_fill_2 FILLER_55_667 ();
 sg13g2_fill_1 FILLER_55_731 ();
 sg13g2_fill_2 FILLER_55_744 ();
 sg13g2_fill_1 FILLER_55_762 ();
 sg13g2_fill_2 FILLER_55_782 ();
 sg13g2_fill_1 FILLER_55_784 ();
 sg13g2_decap_8 FILLER_55_811 ();
 sg13g2_decap_8 FILLER_55_818 ();
 sg13g2_decap_8 FILLER_55_825 ();
 sg13g2_decap_8 FILLER_55_832 ();
 sg13g2_decap_8 FILLER_55_839 ();
 sg13g2_decap_8 FILLER_55_846 ();
 sg13g2_decap_8 FILLER_55_853 ();
 sg13g2_fill_2 FILLER_55_860 ();
 sg13g2_fill_2 FILLER_56_52 ();
 sg13g2_fill_1 FILLER_56_54 ();
 sg13g2_fill_2 FILLER_56_72 ();
 sg13g2_fill_1 FILLER_56_74 ();
 sg13g2_fill_2 FILLER_56_80 ();
 sg13g2_fill_1 FILLER_56_92 ();
 sg13g2_fill_2 FILLER_56_124 ();
 sg13g2_fill_1 FILLER_56_126 ();
 sg13g2_fill_1 FILLER_56_165 ();
 sg13g2_fill_2 FILLER_56_186 ();
 sg13g2_fill_1 FILLER_56_188 ();
 sg13g2_fill_2 FILLER_56_194 ();
 sg13g2_fill_1 FILLER_56_196 ();
 sg13g2_fill_2 FILLER_56_206 ();
 sg13g2_fill_1 FILLER_56_208 ();
 sg13g2_fill_1 FILLER_56_248 ();
 sg13g2_fill_2 FILLER_56_254 ();
 sg13g2_fill_1 FILLER_56_256 ();
 sg13g2_fill_2 FILLER_56_315 ();
 sg13g2_fill_1 FILLER_56_317 ();
 sg13g2_fill_1 FILLER_56_347 ();
 sg13g2_fill_2 FILLER_56_366 ();
 sg13g2_fill_2 FILLER_56_449 ();
 sg13g2_decap_8 FILLER_56_457 ();
 sg13g2_decap_8 FILLER_56_470 ();
 sg13g2_decap_8 FILLER_56_481 ();
 sg13g2_decap_8 FILLER_56_488 ();
 sg13g2_decap_8 FILLER_56_495 ();
 sg13g2_fill_1 FILLER_56_502 ();
 sg13g2_fill_2 FILLER_56_519 ();
 sg13g2_fill_1 FILLER_56_531 ();
 sg13g2_fill_1 FILLER_56_541 ();
 sg13g2_fill_2 FILLER_56_564 ();
 sg13g2_fill_1 FILLER_56_566 ();
 sg13g2_decap_8 FILLER_56_621 ();
 sg13g2_decap_8 FILLER_56_628 ();
 sg13g2_fill_2 FILLER_56_635 ();
 sg13g2_fill_1 FILLER_56_637 ();
 sg13g2_decap_4 FILLER_56_646 ();
 sg13g2_fill_2 FILLER_56_650 ();
 sg13g2_fill_2 FILLER_56_695 ();
 sg13g2_fill_1 FILLER_56_789 ();
 sg13g2_decap_8 FILLER_56_803 ();
 sg13g2_decap_8 FILLER_56_810 ();
 sg13g2_decap_8 FILLER_56_817 ();
 sg13g2_decap_8 FILLER_56_824 ();
 sg13g2_decap_8 FILLER_56_831 ();
 sg13g2_decap_8 FILLER_56_838 ();
 sg13g2_decap_8 FILLER_56_845 ();
 sg13g2_decap_8 FILLER_56_852 ();
 sg13g2_fill_2 FILLER_56_859 ();
 sg13g2_fill_1 FILLER_56_861 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_2 ();
 sg13g2_fill_1 FILLER_57_87 ();
 sg13g2_fill_2 FILLER_57_108 ();
 sg13g2_fill_1 FILLER_57_124 ();
 sg13g2_fill_2 FILLER_57_133 ();
 sg13g2_fill_2 FILLER_57_141 ();
 sg13g2_fill_2 FILLER_57_169 ();
 sg13g2_fill_1 FILLER_57_171 ();
 sg13g2_fill_2 FILLER_57_207 ();
 sg13g2_fill_1 FILLER_57_209 ();
 sg13g2_fill_1 FILLER_57_214 ();
 sg13g2_fill_1 FILLER_57_229 ();
 sg13g2_fill_2 FILLER_57_252 ();
 sg13g2_fill_2 FILLER_57_281 ();
 sg13g2_fill_1 FILLER_57_320 ();
 sg13g2_fill_2 FILLER_57_347 ();
 sg13g2_fill_1 FILLER_57_381 ();
 sg13g2_fill_2 FILLER_57_391 ();
 sg13g2_decap_4 FILLER_57_433 ();
 sg13g2_decap_4 FILLER_57_463 ();
 sg13g2_decap_4 FILLER_57_528 ();
 sg13g2_fill_1 FILLER_57_589 ();
 sg13g2_fill_2 FILLER_57_613 ();
 sg13g2_decap_8 FILLER_57_628 ();
 sg13g2_fill_1 FILLER_57_635 ();
 sg13g2_decap_8 FILLER_57_644 ();
 sg13g2_decap_8 FILLER_57_651 ();
 sg13g2_decap_8 FILLER_57_658 ();
 sg13g2_decap_4 FILLER_57_665 ();
 sg13g2_decap_4 FILLER_57_685 ();
 sg13g2_fill_2 FILLER_57_689 ();
 sg13g2_decap_4 FILLER_57_726 ();
 sg13g2_fill_1 FILLER_57_764 ();
 sg13g2_decap_8 FILLER_57_783 ();
 sg13g2_decap_8 FILLER_57_790 ();
 sg13g2_decap_8 FILLER_57_797 ();
 sg13g2_decap_8 FILLER_57_804 ();
 sg13g2_decap_8 FILLER_57_811 ();
 sg13g2_decap_8 FILLER_57_818 ();
 sg13g2_decap_8 FILLER_57_825 ();
 sg13g2_decap_8 FILLER_57_832 ();
 sg13g2_decap_8 FILLER_57_839 ();
 sg13g2_decap_8 FILLER_57_846 ();
 sg13g2_decap_8 FILLER_57_853 ();
 sg13g2_fill_2 FILLER_57_860 ();
 sg13g2_fill_2 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_37 ();
 sg13g2_fill_2 FILLER_58_57 ();
 sg13g2_fill_1 FILLER_58_91 ();
 sg13g2_fill_2 FILLER_58_115 ();
 sg13g2_fill_1 FILLER_58_117 ();
 sg13g2_fill_1 FILLER_58_141 ();
 sg13g2_fill_1 FILLER_58_191 ();
 sg13g2_fill_1 FILLER_58_224 ();
 sg13g2_fill_1 FILLER_58_349 ();
 sg13g2_fill_2 FILLER_58_360 ();
 sg13g2_fill_2 FILLER_58_385 ();
 sg13g2_fill_2 FILLER_58_415 ();
 sg13g2_decap_4 FILLER_58_443 ();
 sg13g2_fill_1 FILLER_58_447 ();
 sg13g2_decap_4 FILLER_58_458 ();
 sg13g2_fill_1 FILLER_58_462 ();
 sg13g2_fill_1 FILLER_58_477 ();
 sg13g2_fill_1 FILLER_58_482 ();
 sg13g2_fill_2 FILLER_58_516 ();
 sg13g2_fill_1 FILLER_58_547 ();
 sg13g2_fill_2 FILLER_58_564 ();
 sg13g2_fill_1 FILLER_58_566 ();
 sg13g2_fill_2 FILLER_58_605 ();
 sg13g2_decap_8 FILLER_58_695 ();
 sg13g2_fill_2 FILLER_58_702 ();
 sg13g2_fill_1 FILLER_58_704 ();
 sg13g2_fill_2 FILLER_58_756 ();
 sg13g2_decap_8 FILLER_58_763 ();
 sg13g2_decap_8 FILLER_58_775 ();
 sg13g2_decap_8 FILLER_58_782 ();
 sg13g2_decap_8 FILLER_58_789 ();
 sg13g2_decap_8 FILLER_58_796 ();
 sg13g2_decap_8 FILLER_58_803 ();
 sg13g2_decap_8 FILLER_58_810 ();
 sg13g2_decap_8 FILLER_58_817 ();
 sg13g2_decap_8 FILLER_58_824 ();
 sg13g2_decap_8 FILLER_58_831 ();
 sg13g2_decap_8 FILLER_58_838 ();
 sg13g2_decap_8 FILLER_58_845 ();
 sg13g2_decap_8 FILLER_58_852 ();
 sg13g2_fill_2 FILLER_58_859 ();
 sg13g2_fill_1 FILLER_58_861 ();
 sg13g2_fill_2 FILLER_59_26 ();
 sg13g2_fill_1 FILLER_59_28 ();
 sg13g2_fill_1 FILLER_59_60 ();
 sg13g2_fill_2 FILLER_59_78 ();
 sg13g2_fill_1 FILLER_59_80 ();
 sg13g2_fill_2 FILLER_59_127 ();
 sg13g2_fill_1 FILLER_59_189 ();
 sg13g2_fill_1 FILLER_59_218 ();
 sg13g2_fill_1 FILLER_59_225 ();
 sg13g2_fill_2 FILLER_59_239 ();
 sg13g2_fill_1 FILLER_59_257 ();
 sg13g2_fill_2 FILLER_59_299 ();
 sg13g2_fill_1 FILLER_59_341 ();
 sg13g2_fill_2 FILLER_59_366 ();
 sg13g2_fill_1 FILLER_59_373 ();
 sg13g2_fill_1 FILLER_59_410 ();
 sg13g2_fill_2 FILLER_59_425 ();
 sg13g2_fill_1 FILLER_59_427 ();
 sg13g2_fill_1 FILLER_59_498 ();
 sg13g2_fill_2 FILLER_59_539 ();
 sg13g2_fill_1 FILLER_59_576 ();
 sg13g2_decap_4 FILLER_59_627 ();
 sg13g2_fill_2 FILLER_59_644 ();
 sg13g2_fill_1 FILLER_59_646 ();
 sg13g2_decap_4 FILLER_59_726 ();
 sg13g2_fill_1 FILLER_59_730 ();
 sg13g2_fill_2 FILLER_59_783 ();
 sg13g2_fill_2 FILLER_59_794 ();
 sg13g2_fill_2 FILLER_59_810 ();
 sg13g2_fill_1 FILLER_59_812 ();
 sg13g2_decap_8 FILLER_59_821 ();
 sg13g2_decap_8 FILLER_59_828 ();
 sg13g2_decap_8 FILLER_59_835 ();
 sg13g2_decap_8 FILLER_59_842 ();
 sg13g2_decap_8 FILLER_59_849 ();
 sg13g2_decap_4 FILLER_59_856 ();
 sg13g2_fill_2 FILLER_59_860 ();
 sg13g2_fill_2 FILLER_60_22 ();
 sg13g2_fill_1 FILLER_60_81 ();
 sg13g2_fill_2 FILLER_60_95 ();
 sg13g2_fill_2 FILLER_60_120 ();
 sg13g2_fill_2 FILLER_60_149 ();
 sg13g2_fill_1 FILLER_60_151 ();
 sg13g2_fill_1 FILLER_60_162 ();
 sg13g2_fill_1 FILLER_60_181 ();
 sg13g2_fill_1 FILLER_60_193 ();
 sg13g2_fill_1 FILLER_60_204 ();
 sg13g2_fill_1 FILLER_60_249 ();
 sg13g2_fill_1 FILLER_60_267 ();
 sg13g2_fill_1 FILLER_60_334 ();
 sg13g2_fill_2 FILLER_60_361 ();
 sg13g2_fill_1 FILLER_60_363 ();
 sg13g2_fill_2 FILLER_60_437 ();
 sg13g2_fill_1 FILLER_60_439 ();
 sg13g2_fill_1 FILLER_60_449 ();
 sg13g2_fill_2 FILLER_60_469 ();
 sg13g2_decap_8 FILLER_60_475 ();
 sg13g2_fill_1 FILLER_60_482 ();
 sg13g2_decap_4 FILLER_60_542 ();
 sg13g2_fill_2 FILLER_60_546 ();
 sg13g2_fill_1 FILLER_60_592 ();
 sg13g2_fill_2 FILLER_60_653 ();
 sg13g2_fill_1 FILLER_60_655 ();
 sg13g2_decap_4 FILLER_60_666 ();
 sg13g2_fill_1 FILLER_60_670 ();
 sg13g2_fill_2 FILLER_60_706 ();
 sg13g2_fill_2 FILLER_60_753 ();
 sg13g2_fill_2 FILLER_60_773 ();
 sg13g2_fill_1 FILLER_60_801 ();
 sg13g2_decap_8 FILLER_60_828 ();
 sg13g2_decap_8 FILLER_60_835 ();
 sg13g2_decap_8 FILLER_60_842 ();
 sg13g2_decap_8 FILLER_60_849 ();
 sg13g2_decap_4 FILLER_60_856 ();
 sg13g2_fill_2 FILLER_60_860 ();
 sg13g2_fill_2 FILLER_61_31 ();
 sg13g2_fill_1 FILLER_61_33 ();
 sg13g2_fill_2 FILLER_61_96 ();
 sg13g2_fill_1 FILLER_61_98 ();
 sg13g2_fill_2 FILLER_61_122 ();
 sg13g2_fill_1 FILLER_61_124 ();
 sg13g2_fill_2 FILLER_61_131 ();
 sg13g2_fill_1 FILLER_61_133 ();
 sg13g2_fill_1 FILLER_61_161 ();
 sg13g2_fill_2 FILLER_61_171 ();
 sg13g2_fill_1 FILLER_61_234 ();
 sg13g2_fill_2 FILLER_61_269 ();
 sg13g2_fill_1 FILLER_61_281 ();
 sg13g2_fill_2 FILLER_61_313 ();
 sg13g2_fill_1 FILLER_61_315 ();
 sg13g2_fill_1 FILLER_61_352 ();
 sg13g2_fill_1 FILLER_61_377 ();
 sg13g2_fill_1 FILLER_61_413 ();
 sg13g2_fill_1 FILLER_61_428 ();
 sg13g2_fill_1 FILLER_61_438 ();
 sg13g2_decap_4 FILLER_61_444 ();
 sg13g2_fill_1 FILLER_61_448 ();
 sg13g2_decap_4 FILLER_61_457 ();
 sg13g2_fill_2 FILLER_61_461 ();
 sg13g2_fill_1 FILLER_61_489 ();
 sg13g2_fill_2 FILLER_61_495 ();
 sg13g2_fill_1 FILLER_61_497 ();
 sg13g2_fill_1 FILLER_61_508 ();
 sg13g2_fill_1 FILLER_61_556 ();
 sg13g2_fill_2 FILLER_61_565 ();
 sg13g2_fill_1 FILLER_61_567 ();
 sg13g2_fill_2 FILLER_61_586 ();
 sg13g2_fill_1 FILLER_61_588 ();
 sg13g2_decap_8 FILLER_61_658 ();
 sg13g2_decap_4 FILLER_61_665 ();
 sg13g2_fill_1 FILLER_61_674 ();
 sg13g2_decap_8 FILLER_61_720 ();
 sg13g2_fill_2 FILLER_61_727 ();
 sg13g2_decap_4 FILLER_61_781 ();
 sg13g2_fill_1 FILLER_61_785 ();
 sg13g2_fill_1 FILLER_61_790 ();
 sg13g2_fill_2 FILLER_61_805 ();
 sg13g2_fill_1 FILLER_61_807 ();
 sg13g2_decap_8 FILLER_61_848 ();
 sg13g2_decap_8 FILLER_61_855 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_25 ();
 sg13g2_fill_2 FILLER_62_42 ();
 sg13g2_fill_1 FILLER_62_44 ();
 sg13g2_fill_2 FILLER_62_78 ();
 sg13g2_fill_1 FILLER_62_80 ();
 sg13g2_fill_1 FILLER_62_107 ();
 sg13g2_fill_2 FILLER_62_115 ();
 sg13g2_fill_1 FILLER_62_117 ();
 sg13g2_fill_1 FILLER_62_140 ();
 sg13g2_fill_2 FILLER_62_150 ();
 sg13g2_fill_2 FILLER_62_165 ();
 sg13g2_fill_1 FILLER_62_167 ();
 sg13g2_fill_2 FILLER_62_211 ();
 sg13g2_fill_2 FILLER_62_239 ();
 sg13g2_fill_1 FILLER_62_241 ();
 sg13g2_fill_2 FILLER_62_260 ();
 sg13g2_fill_1 FILLER_62_262 ();
 sg13g2_fill_2 FILLER_62_272 ();
 sg13g2_fill_2 FILLER_62_355 ();
 sg13g2_fill_1 FILLER_62_357 ();
 sg13g2_fill_1 FILLER_62_397 ();
 sg13g2_fill_2 FILLER_62_412 ();
 sg13g2_fill_2 FILLER_62_466 ();
 sg13g2_fill_1 FILLER_62_492 ();
 sg13g2_fill_2 FILLER_62_498 ();
 sg13g2_fill_1 FILLER_62_543 ();
 sg13g2_fill_1 FILLER_62_552 ();
 sg13g2_fill_2 FILLER_62_580 ();
 sg13g2_decap_8 FILLER_62_617 ();
 sg13g2_decap_4 FILLER_62_624 ();
 sg13g2_fill_2 FILLER_62_628 ();
 sg13g2_fill_2 FILLER_62_725 ();
 sg13g2_fill_1 FILLER_62_727 ();
 sg13g2_decap_4 FILLER_62_739 ();
 sg13g2_fill_2 FILLER_62_760 ();
 sg13g2_fill_2 FILLER_62_788 ();
 sg13g2_fill_1 FILLER_62_800 ();
 sg13g2_decap_8 FILLER_62_845 ();
 sg13g2_decap_8 FILLER_62_852 ();
 sg13g2_fill_2 FILLER_62_859 ();
 sg13g2_fill_1 FILLER_62_861 ();
 sg13g2_fill_1 FILLER_63_44 ();
 sg13g2_fill_2 FILLER_63_94 ();
 sg13g2_fill_1 FILLER_63_96 ();
 sg13g2_fill_2 FILLER_63_112 ();
 sg13g2_fill_1 FILLER_63_114 ();
 sg13g2_fill_1 FILLER_63_136 ();
 sg13g2_fill_1 FILLER_63_158 ();
 sg13g2_fill_1 FILLER_63_164 ();
 sg13g2_fill_1 FILLER_63_169 ();
 sg13g2_fill_2 FILLER_63_189 ();
 sg13g2_fill_1 FILLER_63_195 ();
 sg13g2_fill_1 FILLER_63_213 ();
 sg13g2_fill_2 FILLER_63_245 ();
 sg13g2_fill_2 FILLER_63_257 ();
 sg13g2_fill_1 FILLER_63_259 ();
 sg13g2_fill_2 FILLER_63_278 ();
 sg13g2_fill_1 FILLER_63_280 ();
 sg13g2_fill_2 FILLER_63_311 ();
 sg13g2_fill_1 FILLER_63_313 ();
 sg13g2_fill_2 FILLER_63_319 ();
 sg13g2_fill_1 FILLER_63_321 ();
 sg13g2_fill_2 FILLER_63_341 ();
 sg13g2_fill_2 FILLER_63_430 ();
 sg13g2_fill_2 FILLER_63_441 ();
 sg13g2_fill_2 FILLER_63_452 ();
 sg13g2_fill_1 FILLER_63_497 ();
 sg13g2_fill_2 FILLER_63_522 ();
 sg13g2_fill_1 FILLER_63_524 ();
 sg13g2_fill_1 FILLER_63_534 ();
 sg13g2_fill_2 FILLER_63_561 ();
 sg13g2_fill_1 FILLER_63_563 ();
 sg13g2_fill_1 FILLER_63_595 ();
 sg13g2_fill_2 FILLER_63_644 ();
 sg13g2_fill_1 FILLER_63_646 ();
 sg13g2_fill_2 FILLER_63_652 ();
 sg13g2_fill_1 FILLER_63_654 ();
 sg13g2_decap_4 FILLER_63_668 ();
 sg13g2_fill_1 FILLER_63_672 ();
 sg13g2_fill_2 FILLER_63_678 ();
 sg13g2_fill_2 FILLER_63_703 ();
 sg13g2_decap_8 FILLER_63_740 ();
 sg13g2_fill_1 FILLER_63_747 ();
 sg13g2_fill_1 FILLER_63_753 ();
 sg13g2_fill_1 FILLER_63_763 ();
 sg13g2_fill_2 FILLER_63_773 ();
 sg13g2_fill_1 FILLER_63_789 ();
 sg13g2_decap_8 FILLER_63_795 ();
 sg13g2_fill_2 FILLER_63_802 ();
 sg13g2_fill_2 FILLER_63_808 ();
 sg13g2_fill_2 FILLER_63_833 ();
 sg13g2_fill_1 FILLER_63_861 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_89 ();
 sg13g2_fill_1 FILLER_64_91 ();
 sg13g2_fill_2 FILLER_64_127 ();
 sg13g2_fill_1 FILLER_64_129 ();
 sg13g2_fill_1 FILLER_64_153 ();
 sg13g2_fill_1 FILLER_64_160 ();
 sg13g2_fill_2 FILLER_64_203 ();
 sg13g2_fill_1 FILLER_64_205 ();
 sg13g2_fill_2 FILLER_64_230 ();
 sg13g2_fill_2 FILLER_64_259 ();
 sg13g2_fill_1 FILLER_64_261 ();
 sg13g2_fill_2 FILLER_64_271 ();
 sg13g2_fill_2 FILLER_64_278 ();
 sg13g2_fill_2 FILLER_64_310 ();
 sg13g2_fill_1 FILLER_64_312 ();
 sg13g2_fill_2 FILLER_64_343 ();
 sg13g2_fill_2 FILLER_64_368 ();
 sg13g2_fill_1 FILLER_64_370 ();
 sg13g2_fill_2 FILLER_64_408 ();
 sg13g2_fill_1 FILLER_64_410 ();
 sg13g2_fill_1 FILLER_64_419 ();
 sg13g2_fill_2 FILLER_64_450 ();
 sg13g2_fill_1 FILLER_64_478 ();
 sg13g2_fill_2 FILLER_64_489 ();
 sg13g2_fill_1 FILLER_64_491 ();
 sg13g2_decap_4 FILLER_64_542 ();
 sg13g2_fill_1 FILLER_64_546 ();
 sg13g2_fill_1 FILLER_64_556 ();
 sg13g2_decap_4 FILLER_64_562 ();
 sg13g2_fill_2 FILLER_64_583 ();
 sg13g2_fill_1 FILLER_64_585 ();
 sg13g2_fill_2 FILLER_64_591 ();
 sg13g2_fill_1 FILLER_64_593 ();
 sg13g2_decap_8 FILLER_64_602 ();
 sg13g2_fill_1 FILLER_64_609 ();
 sg13g2_fill_2 FILLER_64_715 ();
 sg13g2_fill_1 FILLER_64_717 ();
 sg13g2_fill_1 FILLER_64_753 ();
 sg13g2_fill_1 FILLER_64_810 ();
 sg13g2_fill_1 FILLER_64_842 ();
 sg13g2_decap_8 FILLER_64_852 ();
 sg13g2_fill_2 FILLER_64_859 ();
 sg13g2_fill_1 FILLER_64_861 ();
 sg13g2_fill_2 FILLER_65_26 ();
 sg13g2_fill_1 FILLER_65_129 ();
 sg13g2_fill_2 FILLER_65_152 ();
 sg13g2_fill_1 FILLER_65_164 ();
 sg13g2_fill_2 FILLER_65_211 ();
 sg13g2_fill_1 FILLER_65_213 ();
 sg13g2_fill_1 FILLER_65_227 ();
 sg13g2_fill_1 FILLER_65_262 ();
 sg13g2_fill_2 FILLER_65_285 ();
 sg13g2_fill_1 FILLER_65_344 ();
 sg13g2_fill_1 FILLER_65_397 ();
 sg13g2_fill_2 FILLER_65_429 ();
 sg13g2_decap_4 FILLER_65_452 ();
 sg13g2_fill_2 FILLER_65_456 ();
 sg13g2_fill_2 FILLER_65_463 ();
 sg13g2_fill_1 FILLER_65_465 ();
 sg13g2_fill_2 FILLER_65_516 ();
 sg13g2_decap_8 FILLER_65_574 ();
 sg13g2_decap_8 FILLER_65_602 ();
 sg13g2_fill_2 FILLER_65_609 ();
 sg13g2_fill_2 FILLER_65_616 ();
 sg13g2_fill_1 FILLER_65_638 ();
 sg13g2_fill_2 FILLER_65_661 ();
 sg13g2_fill_1 FILLER_65_676 ();
 sg13g2_fill_2 FILLER_65_687 ();
 sg13g2_fill_2 FILLER_65_723 ();
 sg13g2_fill_2 FILLER_65_735 ();
 sg13g2_fill_2 FILLER_65_742 ();
 sg13g2_decap_8 FILLER_65_806 ();
 sg13g2_fill_1 FILLER_65_813 ();
 sg13g2_fill_2 FILLER_65_832 ();
 sg13g2_fill_2 FILLER_65_843 ();
 sg13g2_fill_2 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_24 ();
 sg13g2_fill_1 FILLER_66_80 ();
 sg13g2_fill_2 FILLER_66_109 ();
 sg13g2_fill_1 FILLER_66_111 ();
 sg13g2_fill_1 FILLER_66_138 ();
 sg13g2_fill_2 FILLER_66_148 ();
 sg13g2_fill_1 FILLER_66_172 ();
 sg13g2_fill_1 FILLER_66_207 ();
 sg13g2_fill_1 FILLER_66_241 ();
 sg13g2_fill_1 FILLER_66_257 ();
 sg13g2_fill_1 FILLER_66_267 ();
 sg13g2_fill_2 FILLER_66_314 ();
 sg13g2_fill_1 FILLER_66_402 ();
 sg13g2_fill_2 FILLER_66_411 ();
 sg13g2_fill_1 FILLER_66_413 ();
 sg13g2_fill_2 FILLER_66_472 ();
 sg13g2_fill_2 FILLER_66_484 ();
 sg13g2_fill_2 FILLER_66_499 ();
 sg13g2_fill_1 FILLER_66_501 ();
 sg13g2_fill_1 FILLER_66_517 ();
 sg13g2_fill_1 FILLER_66_541 ();
 sg13g2_fill_2 FILLER_66_551 ();
 sg13g2_fill_1 FILLER_66_553 ();
 sg13g2_fill_2 FILLER_66_568 ();
 sg13g2_fill_2 FILLER_66_590 ();
 sg13g2_fill_1 FILLER_66_592 ();
 sg13g2_decap_8 FILLER_66_607 ();
 sg13g2_fill_2 FILLER_66_614 ();
 sg13g2_fill_1 FILLER_66_616 ();
 sg13g2_fill_2 FILLER_66_629 ();
 sg13g2_fill_1 FILLER_66_631 ();
 sg13g2_decap_4 FILLER_66_637 ();
 sg13g2_fill_2 FILLER_66_641 ();
 sg13g2_fill_1 FILLER_66_674 ();
 sg13g2_decap_4 FILLER_66_734 ();
 sg13g2_fill_2 FILLER_66_756 ();
 sg13g2_fill_1 FILLER_66_762 ();
 sg13g2_decap_8 FILLER_66_768 ();
 sg13g2_fill_2 FILLER_66_775 ();
 sg13g2_fill_1 FILLER_66_797 ();
 sg13g2_fill_1 FILLER_66_803 ();
 sg13g2_fill_2 FILLER_66_832 ();
 sg13g2_fill_1 FILLER_66_834 ();
 sg13g2_fill_1 FILLER_66_861 ();
 sg13g2_fill_1 FILLER_67_53 ();
 sg13g2_fill_2 FILLER_67_67 ();
 sg13g2_fill_1 FILLER_67_69 ();
 sg13g2_fill_2 FILLER_67_75 ();
 sg13g2_fill_2 FILLER_67_122 ();
 sg13g2_fill_1 FILLER_67_124 ();
 sg13g2_fill_2 FILLER_67_183 ();
 sg13g2_fill_1 FILLER_67_185 ();
 sg13g2_fill_2 FILLER_67_214 ();
 sg13g2_fill_2 FILLER_67_228 ();
 sg13g2_fill_2 FILLER_67_238 ();
 sg13g2_fill_1 FILLER_67_319 ();
 sg13g2_fill_1 FILLER_67_394 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_fill_1 FILLER_67_423 ();
 sg13g2_fill_2 FILLER_67_452 ();
 sg13g2_fill_2 FILLER_67_511 ();
 sg13g2_fill_2 FILLER_67_518 ();
 sg13g2_fill_2 FILLER_67_539 ();
 sg13g2_fill_1 FILLER_67_546 ();
 sg13g2_fill_2 FILLER_67_562 ();
 sg13g2_fill_1 FILLER_67_564 ();
 sg13g2_fill_2 FILLER_67_571 ();
 sg13g2_fill_2 FILLER_67_591 ();
 sg13g2_fill_1 FILLER_67_593 ();
 sg13g2_decap_4 FILLER_67_610 ();
 sg13g2_decap_4 FILLER_67_634 ();
 sg13g2_fill_1 FILLER_67_638 ();
 sg13g2_decap_8 FILLER_67_643 ();
 sg13g2_fill_2 FILLER_67_650 ();
 sg13g2_fill_1 FILLER_67_652 ();
 sg13g2_fill_1 FILLER_67_661 ();
 sg13g2_fill_1 FILLER_67_684 ();
 sg13g2_fill_2 FILLER_67_746 ();
 sg13g2_fill_1 FILLER_67_748 ();
 sg13g2_fill_1 FILLER_67_754 ();
 sg13g2_decap_4 FILLER_67_826 ();
 sg13g2_fill_1 FILLER_67_830 ();
 sg13g2_decap_4 FILLER_67_857 ();
 sg13g2_fill_1 FILLER_67_861 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_2 ();
 sg13g2_fill_1 FILLER_68_21 ();
 sg13g2_fill_2 FILLER_68_102 ();
 sg13g2_fill_1 FILLER_68_113 ();
 sg13g2_fill_1 FILLER_68_214 ();
 sg13g2_fill_2 FILLER_68_265 ();
 sg13g2_fill_2 FILLER_68_284 ();
 sg13g2_fill_2 FILLER_68_292 ();
 sg13g2_fill_1 FILLER_68_294 ();
 sg13g2_fill_2 FILLER_68_300 ();
 sg13g2_fill_1 FILLER_68_302 ();
 sg13g2_fill_1 FILLER_68_338 ();
 sg13g2_fill_2 FILLER_68_435 ();
 sg13g2_fill_1 FILLER_68_437 ();
 sg13g2_fill_1 FILLER_68_447 ();
 sg13g2_fill_2 FILLER_68_458 ();
 sg13g2_fill_2 FILLER_68_473 ();
 sg13g2_fill_2 FILLER_68_484 ();
 sg13g2_fill_2 FILLER_68_517 ();
 sg13g2_fill_2 FILLER_68_565 ();
 sg13g2_fill_1 FILLER_68_567 ();
 sg13g2_fill_2 FILLER_68_585 ();
 sg13g2_fill_1 FILLER_68_587 ();
 sg13g2_fill_1 FILLER_68_602 ();
 sg13g2_fill_2 FILLER_68_615 ();
 sg13g2_fill_1 FILLER_68_617 ();
 sg13g2_fill_2 FILLER_68_627 ();
 sg13g2_decap_4 FILLER_68_664 ();
 sg13g2_fill_1 FILLER_68_668 ();
 sg13g2_decap_4 FILLER_68_674 ();
 sg13g2_fill_2 FILLER_68_701 ();
 sg13g2_fill_2 FILLER_68_720 ();
 sg13g2_fill_2 FILLER_68_731 ();
 sg13g2_fill_2 FILLER_68_737 ();
 sg13g2_fill_1 FILLER_68_739 ();
 sg13g2_decap_8 FILLER_68_758 ();
 sg13g2_fill_2 FILLER_68_778 ();
 sg13g2_fill_1 FILLER_68_793 ();
 sg13g2_decap_4 FILLER_68_799 ();
 sg13g2_decap_4 FILLER_68_811 ();
 sg13g2_fill_1 FILLER_68_815 ();
 sg13g2_fill_2 FILLER_68_831 ();
 sg13g2_fill_1 FILLER_68_833 ();
 sg13g2_fill_2 FILLER_68_838 ();
 sg13g2_fill_1 FILLER_68_840 ();
 sg13g2_decap_4 FILLER_68_858 ();
 sg13g2_fill_2 FILLER_69_26 ();
 sg13g2_fill_1 FILLER_69_46 ();
 sg13g2_fill_1 FILLER_69_117 ();
 sg13g2_fill_1 FILLER_69_132 ();
 sg13g2_fill_2 FILLER_69_165 ();
 sg13g2_fill_1 FILLER_69_167 ();
 sg13g2_fill_2 FILLER_69_173 ();
 sg13g2_fill_2 FILLER_69_188 ();
 sg13g2_fill_1 FILLER_69_190 ();
 sg13g2_fill_1 FILLER_69_247 ();
 sg13g2_fill_2 FILLER_69_303 ();
 sg13g2_fill_1 FILLER_69_322 ();
 sg13g2_fill_2 FILLER_69_357 ();
 sg13g2_fill_2 FILLER_69_396 ();
 sg13g2_fill_1 FILLER_69_398 ();
 sg13g2_fill_2 FILLER_69_415 ();
 sg13g2_fill_1 FILLER_69_417 ();
 sg13g2_fill_2 FILLER_69_471 ();
 sg13g2_fill_1 FILLER_69_481 ();
 sg13g2_fill_2 FILLER_69_495 ();
 sg13g2_fill_1 FILLER_69_497 ();
 sg13g2_fill_1 FILLER_69_520 ();
 sg13g2_fill_1 FILLER_69_534 ();
 sg13g2_fill_1 FILLER_69_558 ();
 sg13g2_fill_2 FILLER_69_568 ();
 sg13g2_fill_1 FILLER_69_570 ();
 sg13g2_fill_2 FILLER_69_585 ();
 sg13g2_fill_1 FILLER_69_587 ();
 sg13g2_fill_2 FILLER_69_613 ();
 sg13g2_fill_1 FILLER_69_628 ();
 sg13g2_decap_4 FILLER_69_643 ();
 sg13g2_fill_1 FILLER_69_647 ();
 sg13g2_decap_4 FILLER_69_658 ();
 sg13g2_fill_2 FILLER_69_662 ();
 sg13g2_fill_2 FILLER_69_716 ();
 sg13g2_fill_2 FILLER_69_732 ();
 sg13g2_fill_1 FILLER_69_734 ();
 sg13g2_fill_1 FILLER_69_749 ();
 sg13g2_fill_1 FILLER_69_754 ();
 sg13g2_decap_8 FILLER_69_759 ();
 sg13g2_decap_4 FILLER_69_766 ();
 sg13g2_decap_8 FILLER_69_849 ();
 sg13g2_decap_4 FILLER_69_856 ();
 sg13g2_fill_2 FILLER_69_860 ();
 sg13g2_fill_2 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_2 ();
 sg13g2_fill_1 FILLER_70_25 ();
 sg13g2_fill_2 FILLER_70_54 ();
 sg13g2_fill_1 FILLER_70_82 ();
 sg13g2_fill_2 FILLER_70_109 ();
 sg13g2_fill_1 FILLER_70_207 ();
 sg13g2_fill_1 FILLER_70_226 ();
 sg13g2_fill_2 FILLER_70_296 ();
 sg13g2_fill_1 FILLER_70_360 ();
 sg13g2_fill_2 FILLER_70_396 ();
 sg13g2_fill_1 FILLER_70_424 ();
 sg13g2_fill_1 FILLER_70_439 ();
 sg13g2_fill_2 FILLER_70_452 ();
 sg13g2_fill_1 FILLER_70_454 ();
 sg13g2_fill_2 FILLER_70_460 ();
 sg13g2_fill_2 FILLER_70_506 ();
 sg13g2_fill_1 FILLER_70_508 ();
 sg13g2_decap_4 FILLER_70_579 ();
 sg13g2_fill_1 FILLER_70_583 ();
 sg13g2_fill_1 FILLER_70_588 ();
 sg13g2_fill_1 FILLER_70_593 ();
 sg13g2_decap_8 FILLER_70_609 ();
 sg13g2_fill_1 FILLER_70_616 ();
 sg13g2_fill_2 FILLER_70_639 ();
 sg13g2_fill_2 FILLER_70_676 ();
 sg13g2_fill_1 FILLER_70_686 ();
 sg13g2_fill_1 FILLER_70_718 ();
 sg13g2_fill_1 FILLER_70_732 ();
 sg13g2_fill_2 FILLER_70_737 ();
 sg13g2_fill_2 FILLER_70_792 ();
 sg13g2_fill_2 FILLER_70_807 ();
 sg13g2_fill_2 FILLER_70_818 ();
 sg13g2_fill_1 FILLER_70_820 ();
 sg13g2_fill_1 FILLER_70_861 ();
 sg13g2_fill_1 FILLER_71_61 ();
 sg13g2_fill_2 FILLER_71_80 ();
 sg13g2_fill_1 FILLER_71_109 ();
 sg13g2_fill_1 FILLER_71_218 ();
 sg13g2_fill_1 FILLER_71_243 ();
 sg13g2_fill_1 FILLER_71_261 ();
 sg13g2_fill_2 FILLER_71_290 ();
 sg13g2_fill_1 FILLER_71_305 ();
 sg13g2_fill_1 FILLER_71_341 ();
 sg13g2_fill_2 FILLER_71_387 ();
 sg13g2_fill_2 FILLER_71_424 ();
 sg13g2_fill_2 FILLER_71_489 ();
 sg13g2_fill_1 FILLER_71_491 ();
 sg13g2_fill_1 FILLER_71_524 ();
 sg13g2_fill_1 FILLER_71_538 ();
 sg13g2_fill_2 FILLER_71_558 ();
 sg13g2_fill_2 FILLER_71_564 ();
 sg13g2_decap_8 FILLER_71_640 ();
 sg13g2_fill_2 FILLER_71_660 ();
 sg13g2_fill_1 FILLER_71_662 ();
 sg13g2_fill_1 FILLER_71_672 ();
 sg13g2_decap_4 FILLER_71_678 ();
 sg13g2_fill_1 FILLER_71_723 ();
 sg13g2_fill_2 FILLER_71_778 ();
 sg13g2_fill_2 FILLER_71_794 ();
 sg13g2_fill_2 FILLER_71_801 ();
 sg13g2_fill_1 FILLER_71_847 ();
 sg13g2_decap_4 FILLER_71_857 ();
 sg13g2_fill_1 FILLER_71_861 ();
 sg13g2_fill_2 FILLER_72_0 ();
 sg13g2_fill_1 FILLER_72_2 ();
 sg13g2_fill_1 FILLER_72_74 ();
 sg13g2_fill_2 FILLER_72_89 ();
 sg13g2_fill_1 FILLER_72_91 ();
 sg13g2_fill_1 FILLER_72_148 ();
 sg13g2_fill_1 FILLER_72_163 ();
 sg13g2_fill_2 FILLER_72_242 ();
 sg13g2_fill_1 FILLER_72_244 ();
 sg13g2_fill_2 FILLER_72_255 ();
 sg13g2_fill_1 FILLER_72_288 ();
 sg13g2_fill_2 FILLER_72_370 ();
 sg13g2_fill_1 FILLER_72_388 ();
 sg13g2_fill_2 FILLER_72_397 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_fill_1 FILLER_72_413 ();
 sg13g2_fill_1 FILLER_72_440 ();
 sg13g2_fill_1 FILLER_72_454 ();
 sg13g2_fill_1 FILLER_72_489 ();
 sg13g2_fill_2 FILLER_72_495 ();
 sg13g2_fill_1 FILLER_72_497 ();
 sg13g2_fill_2 FILLER_72_538 ();
 sg13g2_fill_1 FILLER_72_540 ();
 sg13g2_fill_1 FILLER_72_581 ();
 sg13g2_decap_4 FILLER_72_600 ();
 sg13g2_decap_4 FILLER_72_608 ();
 sg13g2_fill_2 FILLER_72_612 ();
 sg13g2_fill_2 FILLER_72_618 ();
 sg13g2_fill_1 FILLER_72_620 ();
 sg13g2_fill_1 FILLER_72_625 ();
 sg13g2_fill_2 FILLER_72_636 ();
 sg13g2_fill_1 FILLER_72_638 ();
 sg13g2_fill_1 FILLER_72_713 ();
 sg13g2_fill_2 FILLER_72_724 ();
 sg13g2_fill_1 FILLER_72_744 ();
 sg13g2_fill_2 FILLER_72_780 ();
 sg13g2_fill_1 FILLER_72_782 ();
 sg13g2_fill_1 FILLER_72_813 ();
 sg13g2_decap_8 FILLER_72_828 ();
 sg13g2_decap_8 FILLER_72_852 ();
 sg13g2_fill_2 FILLER_72_859 ();
 sg13g2_fill_1 FILLER_72_861 ();
 sg13g2_fill_2 FILLER_73_40 ();
 sg13g2_fill_1 FILLER_73_42 ();
 sg13g2_fill_2 FILLER_73_65 ();
 sg13g2_fill_1 FILLER_73_183 ();
 sg13g2_fill_1 FILLER_73_215 ();
 sg13g2_fill_2 FILLER_73_230 ();
 sg13g2_fill_1 FILLER_73_316 ();
 sg13g2_fill_2 FILLER_73_330 ();
 sg13g2_fill_2 FILLER_73_435 ();
 sg13g2_fill_1 FILLER_73_437 ();
 sg13g2_fill_2 FILLER_73_443 ();
 sg13g2_fill_1 FILLER_73_445 ();
 sg13g2_fill_2 FILLER_73_476 ();
 sg13g2_fill_2 FILLER_73_483 ();
 sg13g2_decap_8 FILLER_73_499 ();
 sg13g2_fill_2 FILLER_73_506 ();
 sg13g2_fill_1 FILLER_73_508 ();
 sg13g2_decap_8 FILLER_73_513 ();
 sg13g2_decap_4 FILLER_73_520 ();
 sg13g2_fill_2 FILLER_73_524 ();
 sg13g2_fill_1 FILLER_73_530 ();
 sg13g2_fill_1 FILLER_73_535 ();
 sg13g2_fill_1 FILLER_73_550 ();
 sg13g2_decap_8 FILLER_73_555 ();
 sg13g2_decap_4 FILLER_73_562 ();
 sg13g2_fill_1 FILLER_73_575 ();
 sg13g2_fill_2 FILLER_73_700 ();
 sg13g2_fill_1 FILLER_73_702 ();
 sg13g2_fill_2 FILLER_73_738 ();
 sg13g2_fill_1 FILLER_73_740 ();
 sg13g2_fill_2 FILLER_73_746 ();
 sg13g2_fill_1 FILLER_73_748 ();
 sg13g2_fill_2 FILLER_73_776 ();
 sg13g2_fill_1 FILLER_73_778 ();
 sg13g2_fill_2 FILLER_73_798 ();
 sg13g2_fill_1 FILLER_73_800 ();
 sg13g2_decap_8 FILLER_73_853 ();
 sg13g2_fill_2 FILLER_73_860 ();
 sg13g2_fill_2 FILLER_74_43 ();
 sg13g2_fill_2 FILLER_74_65 ();
 sg13g2_fill_2 FILLER_74_157 ();
 sg13g2_fill_1 FILLER_74_159 ();
 sg13g2_fill_1 FILLER_74_177 ();
 sg13g2_fill_2 FILLER_74_193 ();
 sg13g2_fill_2 FILLER_74_298 ();
 sg13g2_fill_2 FILLER_74_314 ();
 sg13g2_fill_1 FILLER_74_351 ();
 sg13g2_fill_1 FILLER_74_368 ();
 sg13g2_fill_2 FILLER_74_392 ();
 sg13g2_fill_1 FILLER_74_407 ();
 sg13g2_fill_1 FILLER_74_413 ();
 sg13g2_fill_2 FILLER_74_419 ();
 sg13g2_fill_2 FILLER_74_465 ();
 sg13g2_fill_1 FILLER_74_493 ();
 sg13g2_fill_1 FILLER_74_499 ();
 sg13g2_fill_1 FILLER_74_504 ();
 sg13g2_fill_2 FILLER_74_509 ();
 sg13g2_fill_1 FILLER_74_511 ();
 sg13g2_fill_1 FILLER_74_565 ();
 sg13g2_fill_2 FILLER_74_592 ();
 sg13g2_fill_1 FILLER_74_594 ();
 sg13g2_fill_2 FILLER_74_609 ();
 sg13g2_fill_1 FILLER_74_639 ();
 sg13g2_fill_2 FILLER_74_730 ();
 sg13g2_fill_1 FILLER_74_736 ();
 sg13g2_fill_2 FILLER_74_745 ();
 sg13g2_fill_2 FILLER_74_819 ();
 sg13g2_decap_4 FILLER_74_857 ();
 sg13g2_fill_1 FILLER_74_861 ();
 sg13g2_fill_1 FILLER_75_18 ();
 sg13g2_fill_2 FILLER_75_64 ();
 sg13g2_fill_2 FILLER_75_122 ();
 sg13g2_fill_1 FILLER_75_124 ();
 sg13g2_fill_2 FILLER_75_191 ();
 sg13g2_fill_1 FILLER_75_193 ();
 sg13g2_fill_1 FILLER_75_225 ();
 sg13g2_fill_1 FILLER_75_278 ();
 sg13g2_fill_1 FILLER_75_305 ();
 sg13g2_fill_2 FILLER_75_319 ();
 sg13g2_fill_1 FILLER_75_321 ();
 sg13g2_fill_2 FILLER_75_414 ();
 sg13g2_fill_2 FILLER_75_482 ();
 sg13g2_fill_1 FILLER_75_484 ();
 sg13g2_fill_2 FILLER_75_533 ();
 sg13g2_fill_1 FILLER_75_548 ();
 sg13g2_fill_2 FILLER_75_564 ();
 sg13g2_fill_1 FILLER_75_566 ();
 sg13g2_fill_1 FILLER_75_575 ();
 sg13g2_fill_2 FILLER_75_589 ();
 sg13g2_fill_2 FILLER_75_609 ();
 sg13g2_fill_1 FILLER_75_611 ();
 sg13g2_fill_2 FILLER_75_651 ();
 sg13g2_fill_2 FILLER_75_661 ();
 sg13g2_fill_1 FILLER_75_672 ();
 sg13g2_fill_1 FILLER_75_691 ();
 sg13g2_decap_8 FILLER_75_705 ();
 sg13g2_fill_1 FILLER_75_712 ();
 sg13g2_fill_2 FILLER_75_761 ();
 sg13g2_fill_1 FILLER_75_772 ();
 sg13g2_decap_8 FILLER_75_824 ();
 sg13g2_decap_8 FILLER_75_831 ();
 sg13g2_fill_2 FILLER_75_838 ();
 sg13g2_fill_1 FILLER_75_840 ();
 sg13g2_decap_8 FILLER_75_854 ();
 sg13g2_fill_1 FILLER_75_861 ();
 sg13g2_fill_1 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_36 ();
 sg13g2_fill_1 FILLER_76_110 ();
 sg13g2_fill_2 FILLER_76_119 ();
 sg13g2_fill_1 FILLER_76_121 ();
 sg13g2_fill_1 FILLER_76_157 ();
 sg13g2_fill_1 FILLER_76_337 ();
 sg13g2_fill_2 FILLER_76_356 ();
 sg13g2_fill_1 FILLER_76_389 ();
 sg13g2_fill_1 FILLER_76_416 ();
 sg13g2_fill_1 FILLER_76_426 ();
 sg13g2_fill_2 FILLER_76_431 ();
 sg13g2_fill_2 FILLER_76_512 ();
 sg13g2_fill_2 FILLER_76_527 ();
 sg13g2_fill_1 FILLER_76_529 ();
 sg13g2_fill_2 FILLER_76_535 ();
 sg13g2_fill_1 FILLER_76_537 ();
 sg13g2_fill_1 FILLER_76_543 ();
 sg13g2_decap_4 FILLER_76_549 ();
 sg13g2_fill_1 FILLER_76_553 ();
 sg13g2_fill_2 FILLER_76_604 ();
 sg13g2_decap_4 FILLER_76_645 ();
 sg13g2_fill_2 FILLER_76_649 ();
 sg13g2_fill_1 FILLER_76_656 ();
 sg13g2_fill_1 FILLER_76_722 ();
 sg13g2_fill_1 FILLER_76_736 ();
 sg13g2_fill_2 FILLER_76_752 ();
 sg13g2_fill_1 FILLER_76_754 ();
 sg13g2_fill_2 FILLER_76_768 ();
 sg13g2_fill_1 FILLER_76_794 ();
 sg13g2_decap_8 FILLER_76_816 ();
 sg13g2_decap_8 FILLER_76_823 ();
 sg13g2_decap_8 FILLER_76_830 ();
 sg13g2_decap_8 FILLER_76_837 ();
 sg13g2_decap_8 FILLER_76_844 ();
 sg13g2_decap_8 FILLER_76_851 ();
 sg13g2_decap_4 FILLER_76_858 ();
 sg13g2_fill_1 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_19 ();
 sg13g2_fill_2 FILLER_77_46 ();
 sg13g2_fill_1 FILLER_77_48 ();
 sg13g2_fill_2 FILLER_77_113 ();
 sg13g2_fill_2 FILLER_77_150 ();
 sg13g2_fill_1 FILLER_77_152 ();
 sg13g2_fill_2 FILLER_77_197 ();
 sg13g2_fill_2 FILLER_77_255 ();
 sg13g2_fill_2 FILLER_77_302 ();
 sg13g2_fill_1 FILLER_77_304 ();
 sg13g2_fill_2 FILLER_77_336 ();
 sg13g2_fill_1 FILLER_77_338 ();
 sg13g2_fill_1 FILLER_77_348 ();
 sg13g2_fill_2 FILLER_77_393 ();
 sg13g2_fill_2 FILLER_77_443 ();
 sg13g2_fill_2 FILLER_77_454 ();
 sg13g2_fill_2 FILLER_77_495 ();
 sg13g2_fill_1 FILLER_77_497 ();
 sg13g2_decap_4 FILLER_77_549 ();
 sg13g2_fill_2 FILLER_77_553 ();
 sg13g2_fill_1 FILLER_77_560 ();
 sg13g2_fill_1 FILLER_77_586 ();
 sg13g2_fill_2 FILLER_77_646 ();
 sg13g2_fill_1 FILLER_77_648 ();
 sg13g2_fill_2 FILLER_77_684 ();
 sg13g2_fill_1 FILLER_77_686 ();
 sg13g2_fill_2 FILLER_77_708 ();
 sg13g2_fill_2 FILLER_77_745 ();
 sg13g2_decap_8 FILLER_77_825 ();
 sg13g2_decap_8 FILLER_77_832 ();
 sg13g2_decap_8 FILLER_77_839 ();
 sg13g2_decap_8 FILLER_77_846 ();
 sg13g2_decap_8 FILLER_77_853 ();
 sg13g2_fill_2 FILLER_77_860 ();
 sg13g2_fill_1 FILLER_78_60 ();
 sg13g2_fill_1 FILLER_78_70 ();
 sg13g2_fill_2 FILLER_78_100 ();
 sg13g2_fill_1 FILLER_78_102 ();
 sg13g2_fill_1 FILLER_78_168 ();
 sg13g2_fill_2 FILLER_78_191 ();
 sg13g2_fill_1 FILLER_78_267 ();
 sg13g2_fill_2 FILLER_78_299 ();
 sg13g2_fill_2 FILLER_78_307 ();
 sg13g2_fill_1 FILLER_78_309 ();
 sg13g2_fill_2 FILLER_78_336 ();
 sg13g2_fill_1 FILLER_78_338 ();
 sg13g2_fill_1 FILLER_78_348 ();
 sg13g2_fill_2 FILLER_78_406 ();
 sg13g2_fill_1 FILLER_78_413 ();
 sg13g2_fill_2 FILLER_78_429 ();
 sg13g2_fill_2 FILLER_78_448 ();
 sg13g2_fill_1 FILLER_78_467 ();
 sg13g2_fill_1 FILLER_78_498 ();
 sg13g2_fill_1 FILLER_78_525 ();
 sg13g2_fill_2 FILLER_78_534 ();
 sg13g2_decap_4 FILLER_78_545 ();
 sg13g2_fill_2 FILLER_78_549 ();
 sg13g2_fill_1 FILLER_78_577 ();
 sg13g2_fill_2 FILLER_78_587 ();
 sg13g2_fill_1 FILLER_78_589 ();
 sg13g2_decap_4 FILLER_78_625 ();
 sg13g2_decap_4 FILLER_78_655 ();
 sg13g2_fill_1 FILLER_78_659 ();
 sg13g2_fill_2 FILLER_78_664 ();
 sg13g2_decap_8 FILLER_78_670 ();
 sg13g2_fill_2 FILLER_78_677 ();
 sg13g2_fill_1 FILLER_78_679 ();
 sg13g2_decap_4 FILLER_78_720 ();
 sg13g2_fill_1 FILLER_78_729 ();
 sg13g2_decap_4 FILLER_78_734 ();
 sg13g2_fill_1 FILLER_78_738 ();
 sg13g2_decap_8 FILLER_78_748 ();
 sg13g2_fill_2 FILLER_78_755 ();
 sg13g2_fill_1 FILLER_78_757 ();
 sg13g2_decap_8 FILLER_78_762 ();
 sg13g2_decap_8 FILLER_78_769 ();
 sg13g2_fill_2 FILLER_78_776 ();
 sg13g2_fill_1 FILLER_78_778 ();
 sg13g2_decap_4 FILLER_78_783 ();
 sg13g2_fill_1 FILLER_78_787 ();
 sg13g2_decap_8 FILLER_78_797 ();
 sg13g2_fill_2 FILLER_78_804 ();
 sg13g2_decap_8 FILLER_78_815 ();
 sg13g2_decap_8 FILLER_78_822 ();
 sg13g2_decap_8 FILLER_78_829 ();
 sg13g2_decap_8 FILLER_78_836 ();
 sg13g2_decap_8 FILLER_78_843 ();
 sg13g2_decap_8 FILLER_78_850 ();
 sg13g2_decap_4 FILLER_78_857 ();
 sg13g2_fill_1 FILLER_78_861 ();
 sg13g2_fill_1 FILLER_79_166 ();
 sg13g2_fill_1 FILLER_79_207 ();
 sg13g2_fill_1 FILLER_79_303 ();
 sg13g2_fill_2 FILLER_79_349 ();
 sg13g2_fill_1 FILLER_79_410 ();
 sg13g2_fill_2 FILLER_79_441 ();
 sg13g2_fill_2 FILLER_79_492 ();
 sg13g2_fill_2 FILLER_79_503 ();
 sg13g2_fill_1 FILLER_79_505 ();
 sg13g2_fill_1 FILLER_79_541 ();
 sg13g2_fill_2 FILLER_79_564 ();
 sg13g2_fill_1 FILLER_79_566 ();
 sg13g2_fill_2 FILLER_79_581 ();
 sg13g2_fill_1 FILLER_79_583 ();
 sg13g2_decap_8 FILLER_79_657 ();
 sg13g2_decap_8 FILLER_79_664 ();
 sg13g2_decap_8 FILLER_79_671 ();
 sg13g2_decap_8 FILLER_79_678 ();
 sg13g2_decap_8 FILLER_79_685 ();
 sg13g2_decap_4 FILLER_79_692 ();
 sg13g2_decap_8 FILLER_79_700 ();
 sg13g2_decap_8 FILLER_79_707 ();
 sg13g2_decap_8 FILLER_79_714 ();
 sg13g2_decap_8 FILLER_79_721 ();
 sg13g2_decap_8 FILLER_79_728 ();
 sg13g2_decap_8 FILLER_79_735 ();
 sg13g2_decap_8 FILLER_79_742 ();
 sg13g2_decap_8 FILLER_79_749 ();
 sg13g2_decap_8 FILLER_79_756 ();
 sg13g2_decap_8 FILLER_79_763 ();
 sg13g2_decap_8 FILLER_79_770 ();
 sg13g2_decap_8 FILLER_79_777 ();
 sg13g2_decap_8 FILLER_79_784 ();
 sg13g2_decap_8 FILLER_79_791 ();
 sg13g2_decap_8 FILLER_79_798 ();
 sg13g2_decap_8 FILLER_79_805 ();
 sg13g2_decap_8 FILLER_79_812 ();
 sg13g2_decap_8 FILLER_79_819 ();
 sg13g2_decap_8 FILLER_79_826 ();
 sg13g2_decap_8 FILLER_79_833 ();
 sg13g2_decap_8 FILLER_79_840 ();
 sg13g2_decap_8 FILLER_79_847 ();
 sg13g2_decap_8 FILLER_79_854 ();
 sg13g2_fill_1 FILLER_79_861 ();
 sg13g2_fill_2 FILLER_80_0 ();
 sg13g2_fill_1 FILLER_80_2 ();
 sg13g2_fill_1 FILLER_80_43 ();
 sg13g2_fill_2 FILLER_80_70 ();
 sg13g2_fill_2 FILLER_80_90 ();
 sg13g2_fill_2 FILLER_80_133 ();
 sg13g2_fill_1 FILLER_80_175 ();
 sg13g2_fill_2 FILLER_80_185 ();
 sg13g2_fill_1 FILLER_80_296 ();
 sg13g2_fill_2 FILLER_80_311 ();
 sg13g2_fill_2 FILLER_80_471 ();
 sg13g2_fill_2 FILLER_80_499 ();
 sg13g2_fill_1 FILLER_80_535 ();
 sg13g2_fill_1 FILLER_80_606 ();
 sg13g2_decap_8 FILLER_80_646 ();
 sg13g2_decap_8 FILLER_80_653 ();
 sg13g2_decap_8 FILLER_80_660 ();
 sg13g2_decap_8 FILLER_80_667 ();
 sg13g2_decap_8 FILLER_80_674 ();
 sg13g2_decap_8 FILLER_80_681 ();
 sg13g2_decap_8 FILLER_80_688 ();
 sg13g2_decap_8 FILLER_80_695 ();
 sg13g2_decap_8 FILLER_80_702 ();
 sg13g2_decap_8 FILLER_80_709 ();
 sg13g2_decap_8 FILLER_80_716 ();
 sg13g2_decap_8 FILLER_80_723 ();
 sg13g2_decap_8 FILLER_80_730 ();
 sg13g2_decap_8 FILLER_80_737 ();
 sg13g2_decap_8 FILLER_80_744 ();
 sg13g2_decap_8 FILLER_80_751 ();
 sg13g2_decap_8 FILLER_80_758 ();
 sg13g2_decap_8 FILLER_80_765 ();
 sg13g2_decap_8 FILLER_80_772 ();
 sg13g2_decap_8 FILLER_80_779 ();
 sg13g2_decap_8 FILLER_80_786 ();
 sg13g2_decap_8 FILLER_80_793 ();
 sg13g2_decap_8 FILLER_80_800 ();
 sg13g2_decap_8 FILLER_80_807 ();
 sg13g2_decap_8 FILLER_80_814 ();
 sg13g2_decap_8 FILLER_80_821 ();
 sg13g2_decap_8 FILLER_80_828 ();
 sg13g2_decap_8 FILLER_80_835 ();
 sg13g2_decap_8 FILLER_80_842 ();
 sg13g2_decap_8 FILLER_80_849 ();
 sg13g2_decap_4 FILLER_80_856 ();
 sg13g2_fill_2 FILLER_80_860 ();
endmodule

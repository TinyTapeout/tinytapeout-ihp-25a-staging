module tt_um_Esteban_Oman_Mendoza_maze_2024_top (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire Hertz_4;
 wire Hertz_60;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire _463_;
 wire _464_;
 wire _465_;
 wire _466_;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire \counter[0] ;
 wire \counter[10] ;
 wire \counter[11] ;
 wire \counter[12] ;
 wire \counter[13] ;
 wire \counter[14] ;
 wire \counter[15] ;
 wire \counter[16] ;
 wire \counter[17] ;
 wire \counter[18] ;
 wire \counter[19] ;
 wire \counter[1] ;
 wire \counter[20] ;
 wire \counter[21] ;
 wire \counter[22] ;
 wire \counter[23] ;
 wire \counter[24] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire \display_sel[0] ;
 wire \display_sel[1] ;
 wire \display_sel[2] ;
 wire \next_state[0] ;
 wire \next_state[1] ;
 wire \next_state[2] ;
 wire \next_state[3] ;
 wire \next_state[4] ;
 wire \next_state[5] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire \state[4] ;
 wire \state[5] ;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire clknet_0_clk;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net1;
 wire net2;
 wire net3;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;

 sg13g2_inv_1 _473_ (.Y(_427_),
    .A(\state[4] ));
 sg13g2_inv_1 _474_ (.Y(_428_),
    .A(net135));
 sg13g2_inv_2 _475_ (.Y(_429_),
    .A(net133));
 sg13g2_inv_1 _476_ (.Y(_430_),
    .A(_002_));
 sg13g2_inv_1 _477_ (.Y(_431_),
    .A(_003_));
 sg13g2_inv_1 _478_ (.Y(_432_),
    .A(_005_));
 sg13g2_inv_2 _479_ (.Y(_433_),
    .A(net141));
 sg13g2_inv_1 _480_ (.Y(_034_),
    .A(net142));
 sg13g2_inv_1 _481_ (.Y(_035_),
    .A(net45));
 sg13g2_inv_1 _482_ (.Y(_036_),
    .A(net61));
 sg13g2_nor2_1 _483_ (.A(\display_sel[0] ),
    .B(\display_sel[1] ),
    .Y(_037_));
 sg13g2_and2_2 _484_ (.A(_001_),
    .B(_037_),
    .X(_038_));
 sg13g2_nand2b_1 _485_ (.Y(uio_out[0]),
    .B(_038_),
    .A_N(\display_sel[2] ));
 sg13g2_nand2b_1 _486_ (.Y(_039_),
    .B(\display_sel[1] ),
    .A_N(\display_sel[0] ));
 sg13g2_or2_1 _487_ (.X(uio_out[2]),
    .B(_039_),
    .A(\display_sel[2] ));
 sg13g2_nand2b_1 _488_ (.Y(_040_),
    .B(\display_sel[0] ),
    .A_N(\display_sel[1] ));
 sg13g2_a21oi_1 _489_ (.A1(_039_),
    .A2(_040_),
    .Y(_041_),
    .B1(\display_sel[2] ));
 sg13g2_nand2_1 _490_ (.Y(_042_),
    .A(\display_sel[0] ),
    .B(\display_sel[1] ));
 sg13g2_or2_2 _491_ (.X(uio_out[3]),
    .B(_042_),
    .A(\display_sel[2] ));
 sg13g2_nand2_1 _492_ (.Y(_043_),
    .A(\display_sel[2] ),
    .B(_037_));
 sg13g2_nand2_1 _493_ (.Y(_044_),
    .A(uio_out[3]),
    .B(_043_));
 sg13g2_nor3_1 _494_ (.A(_038_),
    .B(_041_),
    .C(_044_),
    .Y(_045_));
 sg13g2_nor2b_1 _495_ (.A(\display_sel[1] ),
    .B_N(_033_),
    .Y(_046_));
 sg13g2_a21oi_1 _496_ (.A1(\display_sel[1] ),
    .A2(_001_),
    .Y(_047_),
    .B1(_046_));
 sg13g2_nand2b_1 _497_ (.Y(uio_out[1]),
    .B(_047_),
    .A_N(_045_));
 sg13g2_nand2b_1 _498_ (.Y(uio_out[4]),
    .B(_037_),
    .A_N(_001_));
 sg13g2_nor2b_2 _499_ (.A(net126),
    .B_N(net124),
    .Y(_048_));
 sg13g2_nand2_1 _500_ (.Y(_049_),
    .A(net125),
    .B(_427_));
 sg13g2_nor2b_2 _501_ (.A(net129),
    .B_N(net131),
    .Y(_050_));
 sg13g2_nand2b_2 _502_ (.Y(_051_),
    .B(net130),
    .A_N(net128));
 sg13g2_nor2_1 _503_ (.A(net136),
    .B(net134),
    .Y(_052_));
 sg13g2_or2_2 _504_ (.X(_053_),
    .B(\state[1] ),
    .A(net135));
 sg13g2_nor2_2 _505_ (.A(net123),
    .B(_053_),
    .Y(_054_));
 sg13g2_and2_2 _506_ (.A(_048_),
    .B(_054_),
    .X(_055_));
 sg13g2_nand2_2 _507_ (.Y(_056_),
    .A(_048_),
    .B(_054_));
 sg13g2_nand2b_2 _508_ (.Y(_057_),
    .B(_056_),
    .A_N(_043_));
 sg13g2_o21ai_1 _509_ (.B1(net124),
    .Y(_058_),
    .A1(net126),
    .A2(net127));
 sg13g2_nand2_1 _510_ (.Y(_059_),
    .A(net124),
    .B(net127));
 sg13g2_and3_1 _511_ (.X(_060_),
    .A(net124),
    .B(net126),
    .C(net127));
 sg13g2_a21oi_2 _512_ (.B1(_060_),
    .Y(_061_),
    .A2(net121),
    .A1(_430_));
 sg13g2_a21o_1 _513_ (.A2(net121),
    .A1(_430_),
    .B1(_060_),
    .X(_062_));
 sg13g2_a21o_1 _514_ (.A2(net126),
    .A1(net124),
    .B1(net127),
    .X(_063_));
 sg13g2_nand2_1 _515_ (.Y(_064_),
    .A(_059_),
    .B(_063_));
 sg13g2_a21oi_1 _516_ (.A1(_059_),
    .A2(_063_),
    .Y(_065_),
    .B1(net132));
 sg13g2_a21o_1 _517_ (.A2(_063_),
    .A1(_059_),
    .B1(net132),
    .X(_066_));
 sg13g2_nor2_1 _518_ (.A(_061_),
    .B(_065_),
    .Y(_067_));
 sg13g2_nand2_1 _519_ (.Y(_068_),
    .A(_062_),
    .B(_066_));
 sg13g2_nor2_2 _520_ (.A(net127),
    .B(net132),
    .Y(_069_));
 sg13g2_or2_2 _521_ (.X(_070_),
    .B(net130),
    .A(net128));
 sg13g2_nand2_1 _522_ (.Y(_071_),
    .A(_431_),
    .B(net121));
 sg13g2_a22oi_1 _523_ (.Y(_072_),
    .B1(_062_),
    .B2(_066_),
    .A2(net121),
    .A1(_431_));
 sg13g2_o21ai_1 _524_ (.B1(_071_),
    .Y(_073_),
    .A1(_061_),
    .A2(_065_));
 sg13g2_o21ai_1 _525_ (.B1(_061_),
    .Y(_074_),
    .A1(_069_),
    .A2(_071_));
 sg13g2_nor3_1 _526_ (.A(_061_),
    .B(_065_),
    .C(_071_),
    .Y(_075_));
 sg13g2_a21o_2 _527_ (.A2(_074_),
    .A1(_068_),
    .B1(_075_),
    .X(_076_));
 sg13g2_a21o_1 _528_ (.A2(_073_),
    .A1(_004_),
    .B1(_064_),
    .X(_077_));
 sg13g2_nand3_1 _529_ (.B(_064_),
    .C(_073_),
    .A(_004_),
    .Y(_078_));
 sg13g2_and2_1 _530_ (.A(_077_),
    .B(_078_),
    .X(_079_));
 sg13g2_xnor2_1 _531_ (.Y(_080_),
    .A(net132),
    .B(_073_));
 sg13g2_xnor2_1 _532_ (.Y(_081_),
    .A(net132),
    .B(_072_));
 sg13g2_a22oi_1 _533_ (.Y(_082_),
    .B1(_080_),
    .B2(_429_),
    .A2(_078_),
    .A1(_077_));
 sg13g2_nor2_1 _534_ (.A(_076_),
    .B(_082_),
    .Y(_083_));
 sg13g2_or2_2 _535_ (.X(_084_),
    .B(_082_),
    .A(_076_));
 sg13g2_a22oi_1 _536_ (.Y(_085_),
    .B1(_080_),
    .B2(_005_),
    .A2(_078_),
    .A1(_077_));
 sg13g2_a21o_1 _537_ (.A2(_074_),
    .A1(_068_),
    .B1(_085_),
    .X(_086_));
 sg13g2_o21ai_1 _538_ (.B1(_076_),
    .Y(_087_),
    .A1(_075_),
    .A2(_085_));
 sg13g2_o21ai_1 _539_ (.B1(_087_),
    .Y(_088_),
    .A1(_083_),
    .A2(_086_));
 sg13g2_o21ai_1 _540_ (.B1(_076_),
    .Y(_089_),
    .A1(net133),
    .A2(_081_));
 sg13g2_a21oi_2 _541_ (.B1(_082_),
    .Y(_090_),
    .A2(_089_),
    .A1(_079_));
 sg13g2_inv_1 _542_ (.Y(_091_),
    .A(_090_));
 sg13g2_o21ai_1 _543_ (.B1(net133),
    .Y(_092_),
    .A1(_076_),
    .A2(_082_));
 sg13g2_or3_1 _544_ (.A(net133),
    .B(_076_),
    .C(_082_),
    .X(_093_));
 sg13g2_nand2_1 _545_ (.Y(_094_),
    .A(_092_),
    .B(_093_));
 sg13g2_and2_1 _546_ (.A(_092_),
    .B(_093_),
    .X(_095_));
 sg13g2_nand3_1 _547_ (.B(_092_),
    .C(_093_),
    .A(net136),
    .Y(_096_));
 sg13g2_o21ai_1 _548_ (.B1(_005_),
    .Y(_097_),
    .A1(_076_),
    .A2(_082_));
 sg13g2_xnor2_1 _549_ (.Y(_098_),
    .A(_080_),
    .B(_097_));
 sg13g2_xnor2_1 _550_ (.Y(_099_),
    .A(_081_),
    .B(_097_));
 sg13g2_nand2_1 _551_ (.Y(_100_),
    .A(_096_),
    .B(_098_));
 sg13g2_a21oi_1 _552_ (.A1(_096_),
    .A2(_098_),
    .Y(_101_),
    .B1(_091_));
 sg13g2_nor4_1 _553_ (.A(_006_),
    .B(_090_),
    .C(_095_),
    .D(_099_),
    .Y(_102_));
 sg13g2_a21o_1 _554_ (.A2(_093_),
    .A1(_092_),
    .B1(net136),
    .X(_103_));
 sg13g2_nor2_1 _555_ (.A(_098_),
    .B(_103_),
    .Y(_104_));
 sg13g2_nor4_1 _556_ (.A(_088_),
    .B(_101_),
    .C(_102_),
    .D(_104_),
    .Y(_105_));
 sg13g2_nor2_1 _557_ (.A(\counter[24] ),
    .B(_056_),
    .Y(_106_));
 sg13g2_nor2b_2 _558_ (.A(_106_),
    .B_N(net146),
    .Y(_107_));
 sg13g2_o21ai_1 _559_ (.B1(net146),
    .Y(_108_),
    .A1(\counter[24] ),
    .A2(_056_));
 sg13g2_a21oi_1 _560_ (.A1(net140),
    .A2(_056_),
    .Y(_109_),
    .B1(_108_));
 sg13g2_nor3_1 _561_ (.A(\display_sel[2] ),
    .B(_040_),
    .C(_109_),
    .Y(_110_));
 sg13g2_a21o_1 _562_ (.A2(_108_),
    .A1(_044_),
    .B1(_045_),
    .X(_111_));
 sg13g2_a21oi_1 _563_ (.A1(net141),
    .A2(_056_),
    .Y(_112_),
    .B1(_108_));
 sg13g2_nor2_1 _564_ (.A(uio_out[2]),
    .B(_112_),
    .Y(_113_));
 sg13g2_nor3_2 _565_ (.A(_110_),
    .B(_111_),
    .C(_113_),
    .Y(_114_));
 sg13g2_a21oi_1 _566_ (.A1(_058_),
    .A2(_072_),
    .Y(_115_),
    .B1(_083_));
 sg13g2_nor2_2 _567_ (.A(uio_out[3]),
    .B(_055_),
    .Y(_116_));
 sg13g2_nor2_1 _568_ (.A(_058_),
    .B(_067_),
    .Y(_117_));
 sg13g2_o21ai_1 _569_ (.B1(_116_),
    .Y(_118_),
    .A1(_084_),
    .A2(_117_));
 sg13g2_o21ai_1 _570_ (.B1(_114_),
    .Y(_119_),
    .A1(_115_),
    .A2(_118_));
 sg13g2_and2_2 _571_ (.A(net135),
    .B(net134),
    .X(_120_));
 sg13g2_nand2_2 _572_ (.Y(_121_),
    .A(\state[0] ),
    .B(\state[1] ));
 sg13g2_xor2_1 _573_ (.B(net133),
    .A(net136),
    .X(_122_));
 sg13g2_mux2_1 _574_ (.A0(net135),
    .A1(_122_),
    .S(net123),
    .X(_123_));
 sg13g2_nor2b_1 _575_ (.A(net130),
    .B_N(net128),
    .Y(_124_));
 sg13g2_nand2b_2 _576_ (.Y(_125_),
    .B(net129),
    .A_N(net130));
 sg13g2_nand3b_1 _577_ (.B(net128),
    .C(net135),
    .Y(_126_),
    .A_N(net130));
 sg13g2_nor2_2 _578_ (.A(net125),
    .B(net126),
    .Y(_127_));
 sg13g2_or2_1 _579_ (.X(_128_),
    .B(net126),
    .A(net125));
 sg13g2_and2_1 _580_ (.A(_126_),
    .B(_127_),
    .X(_129_));
 sg13g2_nor2_2 _581_ (.A(net125),
    .B(_427_),
    .Y(_130_));
 sg13g2_nand2b_1 _582_ (.Y(_131_),
    .B(net126),
    .A_N(net124));
 sg13g2_and2_1 _583_ (.A(net128),
    .B(net130),
    .X(_132_));
 sg13g2_nand2_2 _584_ (.Y(_133_),
    .A(net128),
    .B(net130));
 sg13g2_and2_1 _585_ (.A(_006_),
    .B(_132_),
    .X(_134_));
 sg13g2_a21oi_1 _586_ (.A1(net136),
    .A2(net133),
    .Y(_135_),
    .B1(net127));
 sg13g2_nor2_2 _587_ (.A(_428_),
    .B(net134),
    .Y(_136_));
 sg13g2_nand2b_2 _588_ (.Y(_137_),
    .B(net135),
    .A_N(\state[1] ));
 sg13g2_nor2_1 _589_ (.A(_125_),
    .B(net118),
    .Y(_138_));
 sg13g2_nand2_1 _590_ (.Y(_139_),
    .A(_124_),
    .B(_130_));
 sg13g2_nor3_2 _591_ (.A(_125_),
    .B(net117),
    .C(_137_),
    .Y(_140_));
 sg13g2_nand3_1 _592_ (.B(_002_),
    .C(_004_),
    .A(net124),
    .Y(_141_));
 sg13g2_o21ai_1 _593_ (.B1(_141_),
    .Y(_142_),
    .A1(net122),
    .A2(net118));
 sg13g2_nand2_2 _594_ (.Y(_143_),
    .A(_135_),
    .B(_142_));
 sg13g2_a221oi_1 _595_ (.B2(_134_),
    .C1(_140_),
    .B1(_130_),
    .A1(_123_),
    .Y(_144_),
    .A2(_129_));
 sg13g2_nand2_2 _596_ (.Y(_145_),
    .A(net140),
    .B(net143));
 sg13g2_nand2_1 _597_ (.Y(_146_),
    .A(net141),
    .B(net143));
 sg13g2_o21ai_1 _598_ (.B1(net143),
    .Y(_147_),
    .A1(net141),
    .A2(net140));
 sg13g2_nand2_2 _599_ (.Y(_148_),
    .A(_145_),
    .B(_146_));
 sg13g2_a21o_1 _600_ (.A2(_144_),
    .A1(_143_),
    .B1(_148_),
    .X(_149_));
 sg13g2_nand2_1 _601_ (.Y(_150_),
    .A(net133),
    .B(net131));
 sg13g2_a21o_1 _602_ (.A2(net132),
    .A1(net133),
    .B1(net136),
    .X(_151_));
 sg13g2_o21ai_1 _603_ (.B1(_151_),
    .Y(_152_),
    .A1(_069_),
    .A2(_135_));
 sg13g2_a22oi_1 _604_ (.Y(_153_),
    .B1(_132_),
    .B2(_006_),
    .A2(_124_),
    .A1(_120_));
 sg13g2_a21oi_2 _605_ (.B1(_427_),
    .Y(_154_),
    .A2(_153_),
    .A1(_152_));
 sg13g2_and2_1 _606_ (.A(net127),
    .B(_005_),
    .X(_155_));
 sg13g2_a221oi_1 _607_ (.B2(_050_),
    .C1(_155_),
    .B1(_120_),
    .A1(net122),
    .Y(_156_),
    .A2(_069_));
 sg13g2_o21ai_1 _608_ (.B1(_003_),
    .Y(_157_),
    .A1(net126),
    .A2(_156_));
 sg13g2_nor2_1 _609_ (.A(_154_),
    .B(_157_),
    .Y(_158_));
 sg13g2_or3_1 _610_ (.A(_146_),
    .B(_154_),
    .C(_157_),
    .X(_159_));
 sg13g2_nor2_2 _611_ (.A(_433_),
    .B(_145_),
    .Y(_160_));
 sg13g2_inv_1 _612_ (.Y(_161_),
    .A(_160_));
 sg13g2_xor2_1 _613_ (.B(net130),
    .A(net128),
    .X(_162_));
 sg13g2_o21ai_1 _614_ (.B1(_126_),
    .Y(_163_),
    .A1(_432_),
    .A2(_162_));
 sg13g2_a22oi_1 _615_ (.Y(_164_),
    .B1(net123),
    .B2(_122_),
    .A2(net131),
    .A1(_429_));
 sg13g2_nand2_2 _616_ (.Y(_165_),
    .A(_054_),
    .B(_127_));
 sg13g2_and4_1 _617_ (.A(net124),
    .B(_002_),
    .C(_053_),
    .D(_069_),
    .X(_166_));
 sg13g2_inv_1 _618_ (.Y(_167_),
    .A(_166_));
 sg13g2_a221oi_1 _619_ (.B2(_130_),
    .C1(_166_),
    .B1(_164_),
    .A1(_127_),
    .Y(_168_),
    .A2(_163_));
 sg13g2_nand2_1 _620_ (.Y(_169_),
    .A(_165_),
    .B(_168_));
 sg13g2_a21o_1 _621_ (.A2(_168_),
    .A1(_165_),
    .B1(_145_),
    .X(_170_));
 sg13g2_o21ai_1 _622_ (.B1(net127),
    .Y(_171_),
    .A1(net131),
    .A2(_122_));
 sg13g2_and2_1 _623_ (.A(net131),
    .B(_122_),
    .X(_172_));
 sg13g2_a221oi_1 _624_ (.B2(_428_),
    .C1(net118),
    .B1(_069_),
    .A1(_432_),
    .Y(_173_),
    .A2(_050_));
 sg13g2_o21ai_1 _625_ (.B1(_173_),
    .Y(_174_),
    .A1(_171_),
    .A2(_172_));
 sg13g2_nor2_2 _626_ (.A(net135),
    .B(_429_),
    .Y(_175_));
 sg13g2_nand2b_2 _627_ (.Y(_176_),
    .B(net134),
    .A_N(net135));
 sg13g2_o21ai_1 _628_ (.B1(_127_),
    .Y(_177_),
    .A1(net116),
    .A2(_176_));
 sg13g2_a21o_1 _629_ (.A2(_171_),
    .A1(_150_),
    .B1(_177_),
    .X(_178_));
 sg13g2_and3_1 _630_ (.X(_179_),
    .A(_167_),
    .B(_174_),
    .C(_178_));
 sg13g2_a21oi_2 _631_ (.B1(_160_),
    .Y(_180_),
    .A2(_170_),
    .A1(_159_));
 sg13g2_o21ai_1 _632_ (.B1(_149_),
    .Y(_181_),
    .A1(_161_),
    .A2(_179_));
 sg13g2_nor2_1 _633_ (.A(_180_),
    .B(_181_),
    .Y(_182_));
 sg13g2_or2_1 _634_ (.X(_183_),
    .B(_181_),
    .A(_180_));
 sg13g2_nor2_1 _635_ (.A(net140),
    .B(_146_),
    .Y(_184_));
 sg13g2_nand4_1 _636_ (.B(_174_),
    .C(_178_),
    .A(_167_),
    .Y(_185_),
    .D(_184_));
 sg13g2_o21ai_1 _637_ (.B1(_160_),
    .Y(_186_),
    .A1(_154_),
    .A2(_157_));
 sg13g2_nand3_1 _638_ (.B(_143_),
    .C(_144_),
    .A(_433_),
    .Y(_187_));
 sg13g2_and4_1 _639_ (.A(_148_),
    .B(_185_),
    .C(_186_),
    .D(_187_),
    .X(_188_));
 sg13g2_a21oi_1 _640_ (.A1(_165_),
    .A2(_168_),
    .Y(_189_),
    .B1(_148_));
 sg13g2_nor2_1 _641_ (.A(_188_),
    .B(_189_),
    .Y(_190_));
 sg13g2_nor4_1 _642_ (.A(_180_),
    .B(_181_),
    .C(_188_),
    .D(_189_),
    .Y(_191_));
 sg13g2_o21ai_1 _643_ (.B1(_433_),
    .Y(_192_),
    .A1(_154_),
    .A2(_157_));
 sg13g2_nand3_1 _644_ (.B(_144_),
    .C(_145_),
    .A(_143_),
    .Y(_193_));
 sg13g2_nand3_1 _645_ (.B(_165_),
    .C(_168_),
    .A(_160_),
    .Y(_194_));
 sg13g2_and3_1 _646_ (.X(_195_),
    .A(_148_),
    .B(_193_),
    .C(_194_));
 sg13g2_and4_1 _647_ (.A(_148_),
    .B(_192_),
    .C(_193_),
    .D(_194_),
    .X(_196_));
 sg13g2_nor2_1 _648_ (.A(_148_),
    .B(_179_),
    .Y(_197_));
 sg13g2_nor2_1 _649_ (.A(_196_),
    .B(_197_),
    .Y(_198_));
 sg13g2_nor3_1 _650_ (.A(_148_),
    .B(_154_),
    .C(_157_),
    .Y(_199_));
 sg13g2_nor2_1 _651_ (.A(net141),
    .B(_145_),
    .Y(_200_));
 sg13g2_nand4_1 _652_ (.B(_174_),
    .C(_178_),
    .A(_167_),
    .Y(_201_),
    .D(_200_));
 sg13g2_nand3_1 _653_ (.B(_144_),
    .C(_160_),
    .A(_143_),
    .Y(_202_));
 sg13g2_nand3_1 _654_ (.B(_168_),
    .C(_184_),
    .A(_165_),
    .Y(_203_));
 sg13g2_and4_1 _655_ (.A(_148_),
    .B(_201_),
    .C(_202_),
    .D(_203_),
    .X(_204_));
 sg13g2_nor2_1 _656_ (.A(_199_),
    .B(_204_),
    .Y(_205_));
 sg13g2_a221oi_1 _657_ (.B2(_198_),
    .C1(_204_),
    .B1(_191_),
    .A1(_147_),
    .Y(_206_),
    .A2(_158_));
 sg13g2_o21ai_1 _658_ (.B1(_107_),
    .Y(_207_),
    .A1(_055_),
    .A2(_206_));
 sg13g2_a21oi_1 _659_ (.A1(_038_),
    .A2(_207_),
    .Y(_208_),
    .B1(_119_));
 sg13g2_o21ai_1 _660_ (.B1(_208_),
    .Y(uo_out[0]),
    .A1(_057_),
    .A2(_105_));
 sg13g2_and2_1 _661_ (.A(_096_),
    .B(_099_),
    .X(_209_));
 sg13g2_nand2_1 _662_ (.Y(_210_),
    .A(_096_),
    .B(_099_));
 sg13g2_a21oi_1 _663_ (.A1(_006_),
    .A2(_094_),
    .Y(_211_),
    .B1(_090_));
 sg13g2_a221oi_1 _664_ (.B2(_211_),
    .C1(_088_),
    .B1(_209_),
    .A1(_090_),
    .Y(_212_),
    .A2(_100_));
 sg13g2_a21oi_1 _665_ (.A1(_041_),
    .A2(_108_),
    .Y(_213_),
    .B1(_111_));
 sg13g2_o21ai_1 _666_ (.B1(_116_),
    .Y(_214_),
    .A1(_073_),
    .A2(_084_));
 sg13g2_a21o_1 _667_ (.A2(_084_),
    .A1(_067_),
    .B1(_058_),
    .X(_215_));
 sg13g2_a21oi_1 _668_ (.A1(_067_),
    .A2(_084_),
    .Y(_216_),
    .B1(net121));
 sg13g2_o21ai_1 _669_ (.B1(_213_),
    .Y(_217_),
    .A1(_214_),
    .A2(_215_));
 sg13g2_nor4_1 _670_ (.A(_196_),
    .B(_197_),
    .C(_199_),
    .D(_204_),
    .Y(_218_));
 sg13g2_a221oi_1 _671_ (.B2(_218_),
    .C1(_188_),
    .B1(_182_),
    .A1(_147_),
    .Y(_219_),
    .A2(_169_));
 sg13g2_o21ai_1 _672_ (.B1(_107_),
    .Y(_220_),
    .A1(_055_),
    .A2(_219_));
 sg13g2_a21oi_1 _673_ (.A1(_038_),
    .A2(_220_),
    .Y(_221_),
    .B1(_217_));
 sg13g2_o21ai_1 _674_ (.B1(_221_),
    .Y(uo_out[1]),
    .A1(_057_),
    .A2(_212_));
 sg13g2_nor4_1 _675_ (.A(net136),
    .B(_090_),
    .C(_094_),
    .D(_099_),
    .Y(_222_));
 sg13g2_nor3_1 _676_ (.A(_088_),
    .B(_101_),
    .C(_222_),
    .Y(_223_));
 sg13g2_nand2_1 _677_ (.Y(_224_),
    .A(net121),
    .B(_073_));
 sg13g2_nand4_1 _678_ (.B(_073_),
    .C(_083_),
    .A(net121),
    .Y(_225_),
    .D(_116_));
 sg13g2_nand3_1 _679_ (.B(net146),
    .C(_055_),
    .A(\counter[24] ),
    .Y(_226_));
 sg13g2_nand2_1 _680_ (.Y(_227_),
    .A(_038_),
    .B(_226_));
 sg13g2_and3_1 _681_ (.X(_228_),
    .A(_213_),
    .B(_225_),
    .C(_227_));
 sg13g2_o21ai_1 _682_ (.B1(_228_),
    .Y(uo_out[2]),
    .A1(_057_),
    .A2(_223_));
 sg13g2_a21oi_1 _683_ (.A1(_096_),
    .A2(_103_),
    .Y(_229_),
    .B1(_098_));
 sg13g2_nor4_1 _684_ (.A(_088_),
    .B(_101_),
    .C(_102_),
    .D(_229_),
    .Y(_230_));
 sg13g2_a22oi_1 _685_ (.Y(_231_),
    .B1(_084_),
    .B2(_117_),
    .A2(_073_),
    .A1(net121));
 sg13g2_nand2_1 _686_ (.Y(_232_),
    .A(_116_),
    .B(_224_));
 sg13g2_nand2b_1 _687_ (.Y(_233_),
    .B(_231_),
    .A_N(_118_));
 sg13g2_and3_1 _688_ (.X(_234_),
    .A(_114_),
    .B(_227_),
    .C(_233_));
 sg13g2_o21ai_1 _689_ (.B1(_234_),
    .Y(uo_out[3]),
    .A1(_057_),
    .A2(_230_));
 sg13g2_a21o_1 _690_ (.A2(_098_),
    .A1(_006_),
    .B1(_091_),
    .X(_235_));
 sg13g2_a221oi_1 _691_ (.B2(_099_),
    .C1(_088_),
    .B1(_094_),
    .A1(net136),
    .Y(_236_),
    .A2(_091_));
 sg13g2_a21o_1 _692_ (.A2(_236_),
    .A1(_235_),
    .B1(_057_),
    .X(_237_));
 sg13g2_nand4_1 _693_ (.B(_118_),
    .C(_227_),
    .A(_114_),
    .Y(uo_out[4]),
    .D(_237_));
 sg13g2_a221oi_1 _694_ (.B2(_211_),
    .C1(_088_),
    .B1(_210_),
    .A1(_090_),
    .Y(_238_),
    .A2(_100_));
 sg13g2_o21ai_1 _695_ (.B1(_114_),
    .Y(_239_),
    .A1(_214_),
    .A2(_216_));
 sg13g2_a21oi_1 _696_ (.A1(_190_),
    .A2(_218_),
    .Y(_240_),
    .B1(_183_));
 sg13g2_o21ai_1 _697_ (.B1(_107_),
    .Y(_241_),
    .A1(_055_),
    .A2(_240_));
 sg13g2_a21oi_1 _698_ (.A1(_038_),
    .A2(_241_),
    .Y(_242_),
    .B1(_239_));
 sg13g2_o21ai_1 _699_ (.B1(_242_),
    .Y(uo_out[5]),
    .A1(_057_),
    .A2(_238_));
 sg13g2_a21oi_1 _700_ (.A1(_095_),
    .A2(_098_),
    .Y(_243_),
    .B1(_090_));
 sg13g2_a221oi_1 _701_ (.B2(_243_),
    .C1(_088_),
    .B1(_210_),
    .A1(_090_),
    .Y(_244_),
    .A2(_100_));
 sg13g2_a21oi_1 _702_ (.A1(_041_),
    .A2(_226_),
    .Y(_245_),
    .B1(_111_));
 sg13g2_o21ai_1 _703_ (.B1(_245_),
    .Y(_246_),
    .A1(_216_),
    .A2(_232_));
 sg13g2_a221oi_1 _704_ (.B2(_191_),
    .C1(_197_),
    .B1(_205_),
    .A1(_192_),
    .Y(_247_),
    .A2(_195_));
 sg13g2_o21ai_1 _705_ (.B1(_107_),
    .Y(_248_),
    .A1(_055_),
    .A2(_247_));
 sg13g2_a21oi_1 _706_ (.A1(_038_),
    .A2(_248_),
    .Y(_249_),
    .B1(_246_));
 sg13g2_o21ai_1 _707_ (.B1(_249_),
    .Y(uo_out[6]),
    .A1(_057_),
    .A2(_244_));
 sg13g2_nor2_2 _708_ (.A(net2),
    .B(net142),
    .Y(_250_));
 sg13g2_or2_2 _709_ (.X(_251_),
    .B(net142),
    .A(net140));
 sg13g2_nand2_1 _710_ (.Y(_252_),
    .A(net1),
    .B(_034_));
 sg13g2_nand2_2 _711_ (.Y(_253_),
    .A(net1),
    .B(_250_));
 sg13g2_nor2b_2 _712_ (.A(net142),
    .B_N(net140),
    .Y(_254_));
 sg13g2_inv_1 _713_ (.Y(_255_),
    .A(_254_));
 sg13g2_nor2_2 _714_ (.A(net1),
    .B(net142),
    .Y(_256_));
 sg13g2_nand2_2 _715_ (.Y(_257_),
    .A(_433_),
    .B(_034_));
 sg13g2_nand2_1 _716_ (.Y(_258_),
    .A(net140),
    .B(_256_));
 sg13g2_nand2_2 _717_ (.Y(_259_),
    .A(_253_),
    .B(net139));
 sg13g2_nor2_1 _718_ (.A(_125_),
    .B(net120),
    .Y(_260_));
 sg13g2_nor2_2 _719_ (.A(_049_),
    .B(_070_),
    .Y(_261_));
 sg13g2_nand2_2 _720_ (.Y(_262_),
    .A(_048_),
    .B(_069_));
 sg13g2_nand2_2 _721_ (.Y(_263_),
    .A(_069_),
    .B(_130_));
 sg13g2_a21oi_1 _722_ (.A1(_262_),
    .A2(_263_),
    .Y(_264_),
    .B1(_121_));
 sg13g2_a21oi_1 _723_ (.A1(_136_),
    .A2(net115),
    .Y(_265_),
    .B1(_264_));
 sg13g2_nand3_1 _724_ (.B(_127_),
    .C(_136_),
    .A(_050_),
    .Y(_266_));
 sg13g2_nor2_2 _725_ (.A(_433_),
    .B(_255_),
    .Y(_267_));
 sg13g2_nand2_1 _726_ (.Y(_268_),
    .A(net141),
    .B(_254_));
 sg13g2_nor2_2 _727_ (.A(net141),
    .B(_251_),
    .Y(_269_));
 sg13g2_nand2_2 _728_ (.Y(_270_),
    .A(_433_),
    .B(_250_));
 sg13g2_nor2_1 _729_ (.A(_267_),
    .B(_269_),
    .Y(_271_));
 sg13g2_nor3_1 _730_ (.A(_140_),
    .B(_267_),
    .C(net137),
    .Y(_272_));
 sg13g2_nand2_2 _731_ (.Y(_273_),
    .A(_127_),
    .B(_175_));
 sg13g2_nor2_1 _732_ (.A(_162_),
    .B(_273_),
    .Y(_274_));
 sg13g2_nor2_2 _733_ (.A(_176_),
    .B(_263_),
    .Y(_275_));
 sg13g2_nor3_1 _734_ (.A(_271_),
    .B(_274_),
    .C(_275_),
    .Y(_276_));
 sg13g2_a21oi_1 _735_ (.A1(_266_),
    .A2(_272_),
    .Y(_277_),
    .B1(_276_));
 sg13g2_nand3_1 _736_ (.B(_175_),
    .C(net137),
    .A(_138_),
    .Y(_278_));
 sg13g2_nor3_2 _737_ (.A(_053_),
    .B(_125_),
    .C(net119),
    .Y(_279_));
 sg13g2_nand2_1 _738_ (.Y(_280_),
    .A(net122),
    .B(net115));
 sg13g2_o21ai_1 _739_ (.B1(_278_),
    .Y(_281_),
    .A1(net142),
    .A2(_280_));
 sg13g2_nor2_1 _740_ (.A(_053_),
    .B(_139_),
    .Y(_282_));
 sg13g2_nand2_1 _741_ (.Y(_283_),
    .A(net122),
    .B(_138_));
 sg13g2_a21oi_1 _742_ (.A1(_251_),
    .A2(_257_),
    .Y(_284_),
    .B1(_283_));
 sg13g2_nor2_1 _743_ (.A(_070_),
    .B(net120),
    .Y(_285_));
 sg13g2_nor4_2 _744_ (.A(_070_),
    .B(_121_),
    .C(net119),
    .Y(_286_),
    .D(net137));
 sg13g2_nor4_1 _745_ (.A(_277_),
    .B(_281_),
    .C(_284_),
    .D(_286_),
    .Y(_287_));
 sg13g2_o21ai_1 _746_ (.B1(_287_),
    .Y(_288_),
    .A1(_259_),
    .A2(_265_));
 sg13g2_nor3_1 _747_ (.A(_121_),
    .B(net119),
    .C(_133_),
    .Y(_289_));
 sg13g2_nand2_1 _748_ (.Y(_290_),
    .A(_257_),
    .B(_289_));
 sg13g2_nor3_2 _749_ (.A(_053_),
    .B(net118),
    .C(_133_),
    .Y(_291_));
 sg13g2_nor3_2 _750_ (.A(_121_),
    .B(net117),
    .C(net116),
    .Y(_292_));
 sg13g2_a22oi_1 _751_ (.Y(_293_),
    .B1(_292_),
    .B2(net142),
    .A2(_291_),
    .A1(_267_));
 sg13g2_nor3_2 _752_ (.A(_429_),
    .B(_126_),
    .C(net118),
    .Y(_294_));
 sg13g2_nand3_1 _753_ (.B(net138),
    .C(_294_),
    .A(_253_),
    .Y(_295_));
 sg13g2_nor3_2 _754_ (.A(_051_),
    .B(_121_),
    .C(net119),
    .Y(_296_));
 sg13g2_nand3_1 _755_ (.B(_120_),
    .C(_127_),
    .A(_050_),
    .Y(_297_));
 sg13g2_nand2_1 _756_ (.Y(_298_),
    .A(_255_),
    .B(_296_));
 sg13g2_nand4_1 _757_ (.B(_293_),
    .C(_295_),
    .A(_290_),
    .Y(_299_),
    .D(_298_));
 sg13g2_nor3_1 _758_ (.A(_053_),
    .B(net119),
    .C(net116),
    .Y(_300_));
 sg13g2_nand2_1 _759_ (.Y(_301_),
    .A(_259_),
    .B(_300_));
 sg13g2_nor3_2 _760_ (.A(_051_),
    .B(_053_),
    .C(net118),
    .Y(_302_));
 sg13g2_nand2_1 _761_ (.Y(_303_),
    .A(_256_),
    .B(_302_));
 sg13g2_nand3_1 _762_ (.B(_261_),
    .C(_267_),
    .A(net122),
    .Y(_304_));
 sg13g2_nand3_1 _763_ (.B(_132_),
    .C(_136_),
    .A(_130_),
    .Y(_305_));
 sg13g2_nand2b_1 _764_ (.Y(_306_),
    .B(_257_),
    .A_N(_305_));
 sg13g2_nand4_1 _765_ (.B(_303_),
    .C(_304_),
    .A(_301_),
    .Y(_307_),
    .D(_306_));
 sg13g2_nor3_2 _766_ (.A(_051_),
    .B(net117),
    .C(_176_),
    .Y(_308_));
 sg13g2_a21oi_1 _767_ (.A1(_175_),
    .A2(_261_),
    .Y(_309_),
    .B1(_308_));
 sg13g2_nor2_1 _768_ (.A(_053_),
    .B(_263_),
    .Y(_310_));
 sg13g2_nor2b_1 _769_ (.A(_273_),
    .B_N(_162_),
    .Y(_311_));
 sg13g2_nor2_1 _770_ (.A(net123),
    .B(_273_),
    .Y(_312_));
 sg13g2_o21ai_1 _771_ (.B1(_256_),
    .Y(_313_),
    .A1(_310_),
    .A2(_311_));
 sg13g2_o21ai_1 _772_ (.B1(_313_),
    .Y(_314_),
    .A1(_252_),
    .A2(_309_));
 sg13g2_nor4_1 _773_ (.A(_288_),
    .B(_299_),
    .C(_307_),
    .D(_314_),
    .Y(_315_));
 sg13g2_nor3_2 _774_ (.A(net123),
    .B(_121_),
    .C(net117),
    .Y(_316_));
 sg13g2_nor3_2 _775_ (.A(_070_),
    .B(net119),
    .C(_137_),
    .Y(_317_));
 sg13g2_a22oi_1 _776_ (.Y(_318_),
    .B1(_317_),
    .B2(_252_),
    .A2(net115),
    .A1(_120_));
 sg13g2_nand2b_1 _777_ (.Y(_319_),
    .B(_318_),
    .A_N(_316_));
 sg13g2_nor3_2 _778_ (.A(net117),
    .B(net116),
    .C(_176_),
    .Y(_320_));
 sg13g2_a21oi_1 _779_ (.A1(_175_),
    .A2(net115),
    .Y(_321_),
    .B1(_320_));
 sg13g2_o21ai_1 _780_ (.B1(_321_),
    .Y(_322_),
    .A1(_176_),
    .A2(_262_));
 sg13g2_a22oi_1 _781_ (.Y(_323_),
    .B1(_322_),
    .B2(_254_),
    .A2(_319_),
    .A1(_251_));
 sg13g2_nor3_2 _782_ (.A(_429_),
    .B(net120),
    .C(net116),
    .Y(_324_));
 sg13g2_a21oi_2 _783_ (.B1(_300_),
    .Y(_325_),
    .A2(_260_),
    .A1(_136_));
 sg13g2_nor2b_1 _784_ (.A(_324_),
    .B_N(_325_),
    .Y(_326_));
 sg13g2_a21oi_1 _785_ (.A1(_052_),
    .A2(_261_),
    .Y(_327_),
    .B1(_055_));
 sg13g2_nor3_2 _786_ (.A(net134),
    .B(net123),
    .C(net120),
    .Y(_328_));
 sg13g2_nor2_1 _787_ (.A(net122),
    .B(_262_),
    .Y(_329_));
 sg13g2_nand2_1 _788_ (.Y(_330_),
    .A(net134),
    .B(net115));
 sg13g2_o21ai_1 _789_ (.B1(_330_),
    .Y(_331_),
    .A1(net123),
    .A2(_273_));
 sg13g2_nor4_1 _790_ (.A(_130_),
    .B(_328_),
    .C(_329_),
    .D(_331_),
    .Y(_332_));
 sg13g2_nand4_1 _791_ (.B(_326_),
    .C(_327_),
    .A(_297_),
    .Y(_333_),
    .D(_332_));
 sg13g2_nor3_2 _792_ (.A(net120),
    .B(net116),
    .C(_137_),
    .Y(_334_));
 sg13g2_nor3_1 _793_ (.A(net122),
    .B(_070_),
    .C(net119),
    .Y(_335_));
 sg13g2_nor4_1 _794_ (.A(_253_),
    .B(_279_),
    .C(_334_),
    .D(_335_),
    .Y(_336_));
 sg13g2_nand2b_1 _795_ (.Y(_337_),
    .B(_336_),
    .A_N(_333_));
 sg13g2_nor3_1 _796_ (.A(net123),
    .B(net117),
    .C(_137_),
    .Y(_338_));
 sg13g2_nand3_1 _797_ (.B(_130_),
    .C(_136_),
    .A(_050_),
    .Y(_339_));
 sg13g2_nor3_1 _798_ (.A(net128),
    .B(net117),
    .C(_137_),
    .Y(_340_));
 sg13g2_nor2_1 _799_ (.A(_137_),
    .B(_262_),
    .Y(_341_));
 sg13g2_o21ai_1 _800_ (.B1(_253_),
    .Y(_342_),
    .A1(_334_),
    .A2(_341_));
 sg13g2_o21ai_1 _801_ (.B1(_342_),
    .Y(_343_),
    .A1(net143),
    .A2(_165_));
 sg13g2_o21ai_1 _802_ (.B1(_255_),
    .Y(_344_),
    .A1(_340_),
    .A2(_343_));
 sg13g2_nand4_1 _803_ (.B(_323_),
    .C(_337_),
    .A(_315_),
    .Y(_434_),
    .D(_344_));
 sg13g2_nor3_1 _804_ (.A(_137_),
    .B(net139),
    .C(_263_),
    .Y(_345_));
 sg13g2_o21ai_1 _805_ (.B1(_259_),
    .Y(_346_),
    .A1(_334_),
    .A2(_345_));
 sg13g2_o21ai_1 _806_ (.B1(net139),
    .Y(_347_),
    .A1(_264_),
    .A2(_320_));
 sg13g2_o21ai_1 _807_ (.B1(_279_),
    .Y(_348_),
    .A1(_250_),
    .A2(_256_));
 sg13g2_o21ai_1 _808_ (.B1(_348_),
    .Y(_349_),
    .A1(_257_),
    .A2(_305_));
 sg13g2_a221oi_1 _809_ (.B2(_257_),
    .C1(_349_),
    .B1(_311_),
    .A1(_270_),
    .Y(_350_),
    .A2(_275_));
 sg13g2_nor3_1 _810_ (.A(_176_),
    .B(_259_),
    .C(_262_),
    .Y(_351_));
 sg13g2_a21o_1 _811_ (.A2(_317_),
    .A1(_250_),
    .B1(_351_),
    .X(_352_));
 sg13g2_a221oi_1 _812_ (.B2(_253_),
    .C1(_352_),
    .B1(_308_),
    .A1(_271_),
    .Y(_353_),
    .A2(_274_));
 sg13g2_and4_1 _813_ (.A(_346_),
    .B(_347_),
    .C(_350_),
    .D(_353_),
    .X(_354_));
 sg13g2_nand2_1 _814_ (.Y(_355_),
    .A(_270_),
    .B(_316_));
 sg13g2_nand3b_1 _815_ (.B(_303_),
    .C(_355_),
    .Y(_356_),
    .A_N(_286_));
 sg13g2_a22oi_1 _816_ (.Y(_357_),
    .B1(_282_),
    .B2(_256_),
    .A2(net137),
    .A1(_140_));
 sg13g2_a22oi_1 _817_ (.Y(_358_),
    .B1(net115),
    .B2(_120_),
    .A2(_175_),
    .A1(_138_));
 sg13g2_o21ai_1 _818_ (.B1(_357_),
    .Y(_359_),
    .A1(_269_),
    .A2(_358_));
 sg13g2_nor3_1 _819_ (.A(_299_),
    .B(_356_),
    .C(_359_),
    .Y(_360_));
 sg13g2_o21ai_1 _820_ (.B1(_339_),
    .Y(_361_),
    .A1(net141),
    .A2(_325_));
 sg13g2_o21ai_1 _821_ (.B1(_254_),
    .Y(_362_),
    .A1(_341_),
    .A2(_361_));
 sg13g2_o21ai_1 _822_ (.B1(_269_),
    .Y(_363_),
    .A1(_310_),
    .A2(_328_));
 sg13g2_nand4_1 _823_ (.B(_360_),
    .C(_362_),
    .A(_354_),
    .Y(_435_),
    .D(_363_));
 sg13g2_o21ai_1 _824_ (.B1(_268_),
    .Y(_364_),
    .A1(_291_),
    .A2(_296_));
 sg13g2_nor3_1 _825_ (.A(net134),
    .B(net119),
    .C(net116),
    .Y(_365_));
 sg13g2_o21ai_1 _826_ (.B1(net138),
    .Y(_366_),
    .A1(_289_),
    .A2(_365_));
 sg13g2_nor2_1 _827_ (.A(net139),
    .B(_283_),
    .Y(_367_));
 sg13g2_nor2_1 _828_ (.A(_251_),
    .B(_280_),
    .Y(_368_));
 sg13g2_nor4_1 _829_ (.A(_338_),
    .B(_345_),
    .C(_367_),
    .D(_368_),
    .Y(_369_));
 sg13g2_nor2b_1 _830_ (.A(_305_),
    .B_N(net138),
    .Y(_370_));
 sg13g2_nor2_1 _831_ (.A(_320_),
    .B(_370_),
    .Y(_371_));
 sg13g2_o21ai_1 _832_ (.B1(_270_),
    .Y(_372_),
    .A1(_302_),
    .A2(_312_));
 sg13g2_nor2b_1 _833_ (.A(_275_),
    .B_N(_330_),
    .Y(_373_));
 sg13g2_o21ai_1 _834_ (.B1(_372_),
    .Y(_374_),
    .A1(_270_),
    .A2(_373_));
 sg13g2_o21ai_1 _835_ (.B1(_056_),
    .Y(_375_),
    .A1(net116),
    .A2(_273_));
 sg13g2_nor4_1 _836_ (.A(_292_),
    .B(_308_),
    .C(_328_),
    .D(_375_),
    .Y(_376_));
 sg13g2_nand2_1 _837_ (.Y(_377_),
    .A(_259_),
    .B(_294_));
 sg13g2_nand3_1 _838_ (.B(_376_),
    .C(_377_),
    .A(_355_),
    .Y(_378_));
 sg13g2_nor4_1 _839_ (.A(_320_),
    .B(_370_),
    .C(_374_),
    .D(_378_),
    .Y(_379_));
 sg13g2_nand4_1 _840_ (.B(_366_),
    .C(_369_),
    .A(_364_),
    .Y(_436_),
    .D(_379_));
 sg13g2_nor3_1 _841_ (.A(net122),
    .B(net138),
    .C(_262_),
    .Y(_380_));
 sg13g2_a21o_1 _842_ (.A2(_292_),
    .A1(net142),
    .B1(_380_),
    .X(_381_));
 sg13g2_nor2_1 _843_ (.A(net138),
    .B(_339_),
    .Y(_382_));
 sg13g2_nor2_1 _844_ (.A(_139_),
    .B(net137),
    .Y(_383_));
 sg13g2_a21o_1 _845_ (.A2(net115),
    .A1(_122_),
    .B1(_294_),
    .X(_384_));
 sg13g2_a22oi_1 _846_ (.Y(_385_),
    .B1(_383_),
    .B2(_122_),
    .A2(_282_),
    .A1(_257_));
 sg13g2_o21ai_1 _847_ (.B1(_385_),
    .Y(_386_),
    .A1(_259_),
    .A2(_280_));
 sg13g2_a21oi_1 _848_ (.A1(_267_),
    .A2(_296_),
    .Y(_387_),
    .B1(_386_));
 sg13g2_or3_1 _849_ (.A(_270_),
    .B(_316_),
    .C(_335_),
    .X(_388_));
 sg13g2_o21ai_1 _850_ (.B1(_388_),
    .Y(_389_),
    .A1(net137),
    .A2(_324_));
 sg13g2_a21oi_1 _851_ (.A1(net138),
    .A2(_384_),
    .Y(_390_),
    .B1(_381_));
 sg13g2_nor2_1 _852_ (.A(_365_),
    .B(_382_),
    .Y(_391_));
 sg13g2_a221oi_1 _853_ (.B2(_275_),
    .C1(_291_),
    .B1(net137),
    .A1(_120_),
    .Y(_392_),
    .A2(net115));
 sg13g2_and4_1 _854_ (.A(_387_),
    .B(_389_),
    .C(_391_),
    .D(_392_),
    .X(_393_));
 sg13g2_nand4_1 _855_ (.B(_371_),
    .C(_390_),
    .A(_303_),
    .Y(_437_),
    .D(_393_));
 sg13g2_o21ai_1 _856_ (.B1(net138),
    .Y(_394_),
    .A1(_302_),
    .A2(_340_));
 sg13g2_o21ai_1 _857_ (.B1(net137),
    .Y(_395_),
    .A1(_312_),
    .A2(_324_));
 sg13g2_a22oi_1 _858_ (.Y(_396_),
    .B1(_137_),
    .B2(_069_),
    .A2(_132_),
    .A1(_121_));
 sg13g2_nor4_1 _859_ (.A(_294_),
    .B(_308_),
    .C(_316_),
    .D(_383_),
    .Y(_397_));
 sg13g2_o21ai_1 _860_ (.B1(_397_),
    .Y(_398_),
    .A1(net117),
    .A2(_396_));
 sg13g2_nor2_1 _861_ (.A(_381_),
    .B(_398_),
    .Y(_399_));
 sg13g2_nand3_1 _862_ (.B(_395_),
    .C(_399_),
    .A(_394_),
    .Y(_438_));
 sg13g2_nand2_1 _863_ (.Y(_400_),
    .A(_278_),
    .B(_327_));
 sg13g2_a221oi_1 _864_ (.B2(net138),
    .C1(_400_),
    .B1(_329_),
    .A1(_034_),
    .Y(_401_),
    .A2(_292_));
 sg13g2_o21ai_1 _865_ (.B1(_401_),
    .Y(_439_),
    .A1(net140),
    .A2(_357_));
 sg13g2_and2_1 _866_ (.A(net144),
    .B(\counter[15] ),
    .X(Hertz_60));
 sg13g2_and2_2 _867_ (.A(net146),
    .B(\counter[23] ),
    .X(Hertz_4));
 sg13g2_nor4_2 _868_ (.A(_279_),
    .B(_285_),
    .C(_333_),
    .Y(_000_),
    .D(_334_));
 sg13g2_xor2_1 _869_ (.B(net50),
    .A(\counter[1] ),
    .X(_017_));
 sg13g2_nand3_1 _870_ (.B(net50),
    .C(net63),
    .A(\counter[1] ),
    .Y(_402_));
 sg13g2_a21o_1 _871_ (.A2(net50),
    .A1(\counter[1] ),
    .B1(net63),
    .X(_403_));
 sg13g2_and2_1 _872_ (.A(_402_),
    .B(net64),
    .X(_023_));
 sg13g2_and4_1 _873_ (.A(\counter[1] ),
    .B(\counter[0] ),
    .C(\counter[2] ),
    .D(net32),
    .X(_404_));
 sg13g2_xnor2_1 _874_ (.Y(_024_),
    .A(net32),
    .B(_402_));
 sg13g2_and2_1 _875_ (.A(\counter[4] ),
    .B(_404_),
    .X(_405_));
 sg13g2_xor2_1 _876_ (.B(_404_),
    .A(net41),
    .X(_025_));
 sg13g2_xor2_1 _877_ (.B(_405_),
    .A(net37),
    .X(_026_));
 sg13g2_nand4_1 _878_ (.B(net37),
    .C(net59),
    .A(net41),
    .Y(_406_),
    .D(_404_));
 sg13g2_a21o_1 _879_ (.A2(_405_),
    .A1(net37),
    .B1(net59),
    .X(_407_));
 sg13g2_and2_1 _880_ (.A(_406_),
    .B(net60),
    .X(_027_));
 sg13g2_xnor2_1 _881_ (.Y(_028_),
    .A(net45),
    .B(_406_));
 sg13g2_nor3_2 _882_ (.A(_035_),
    .B(_036_),
    .C(_406_),
    .Y(_408_));
 sg13g2_o21ai_1 _883_ (.B1(_036_),
    .Y(_409_),
    .A1(_035_),
    .A2(_406_));
 sg13g2_nor2b_1 _884_ (.A(_408_),
    .B_N(_409_),
    .Y(_029_));
 sg13g2_xor2_1 _885_ (.B(_408_),
    .A(net47),
    .X(_030_));
 sg13g2_and3_2 _886_ (.X(_410_),
    .A(net47),
    .B(net29),
    .C(_408_));
 sg13g2_a21oi_1 _887_ (.A1(\counter[9] ),
    .A2(_408_),
    .Y(_411_),
    .B1(net29));
 sg13g2_nor2_1 _888_ (.A(_410_),
    .B(net30),
    .Y(_007_));
 sg13g2_xor2_1 _889_ (.B(_410_),
    .A(net53),
    .X(_008_));
 sg13g2_nand3_1 _890_ (.B(net66),
    .C(_410_),
    .A(net53),
    .Y(_412_));
 sg13g2_a21o_1 _891_ (.A2(_410_),
    .A1(net53),
    .B1(net66),
    .X(_413_));
 sg13g2_and2_1 _892_ (.A(_412_),
    .B(_413_),
    .X(_009_));
 sg13g2_and4_1 _893_ (.A(net67),
    .B(\counter[12] ),
    .C(net27),
    .D(_410_),
    .X(_414_));
 sg13g2_xnor2_1 _894_ (.Y(_010_),
    .A(net27),
    .B(_412_));
 sg13g2_xor2_1 _895_ (.B(_414_),
    .A(net39),
    .X(_011_));
 sg13g2_nand3_1 _896_ (.B(net39),
    .C(net68),
    .A(net34),
    .Y(_415_));
 sg13g2_inv_1 _897_ (.Y(_416_),
    .A(_415_));
 sg13g2_a21oi_1 _898_ (.A1(\counter[14] ),
    .A2(_414_),
    .Y(_417_),
    .B1(net34));
 sg13g2_nor2_1 _899_ (.A(_416_),
    .B(net35),
    .Y(_012_));
 sg13g2_xnor2_1 _900_ (.Y(_013_),
    .A(net49),
    .B(_415_));
 sg13g2_nand2_1 _901_ (.Y(_418_),
    .A(net49),
    .B(net22));
 sg13g2_nor2_2 _902_ (.A(_415_),
    .B(_418_),
    .Y(_419_));
 sg13g2_a21oi_1 _903_ (.A1(\counter[16] ),
    .A2(_416_),
    .Y(_420_),
    .B1(net22));
 sg13g2_nor2_1 _904_ (.A(_419_),
    .B(net23),
    .Y(_014_));
 sg13g2_xor2_1 _905_ (.B(_419_),
    .A(net52),
    .X(_015_));
 sg13g2_nand3_1 _906_ (.B(net62),
    .C(_419_),
    .A(net52),
    .Y(_421_));
 sg13g2_a21o_1 _907_ (.A2(_419_),
    .A1(net52),
    .B1(net62),
    .X(_422_));
 sg13g2_and2_1 _908_ (.A(_421_),
    .B(_422_),
    .X(_016_));
 sg13g2_and4_2 _909_ (.A(net52),
    .B(\counter[19] ),
    .C(net25),
    .D(_419_),
    .X(_423_));
 sg13g2_xnor2_1 _910_ (.Y(_018_),
    .A(net25),
    .B(_421_));
 sg13g2_xor2_1 _911_ (.B(_423_),
    .A(net54),
    .X(_019_));
 sg13g2_nand3_1 _912_ (.B(net56),
    .C(_423_),
    .A(net54),
    .Y(_424_));
 sg13g2_a21o_1 _913_ (.A2(_423_),
    .A1(net54),
    .B1(net56),
    .X(_425_));
 sg13g2_and2_1 _914_ (.A(_424_),
    .B(_425_),
    .X(_020_));
 sg13g2_nand4_1 _915_ (.B(net54),
    .C(net56),
    .A(net43),
    .Y(_426_),
    .D(_423_));
 sg13g2_xnor2_1 _916_ (.Y(_021_),
    .A(net43),
    .B(_424_));
 sg13g2_xnor2_1 _917_ (.Y(_022_),
    .A(\counter[24] ),
    .B(net57));
 sg13g2_nand2_1 _918_ (.Y(_031_),
    .A(_039_),
    .B(_040_));
 sg13g2_xnor2_1 _919_ (.Y(_032_),
    .A(\display_sel[2] ),
    .B(_042_));
 sg13g2_dllrq_1 _920_ (.D(_434_),
    .GATE_N(_000_),
    .RESET_B(net3),
    .Q(\next_state[0] ));
 sg13g2_dllrq_1 _921_ (.D(_435_),
    .GATE_N(_000_),
    .RESET_B(net4),
    .Q(\next_state[1] ));
 sg13g2_dllrq_1 _922_ (.D(_436_),
    .GATE_N(_000_),
    .RESET_B(net5),
    .Q(\next_state[2] ));
 sg13g2_dllrq_1 _923_ (.D(_437_),
    .GATE_N(_000_),
    .RESET_B(net6),
    .Q(\next_state[3] ));
 sg13g2_dllrq_1 _924_ (.D(_438_),
    .GATE_N(_000_),
    .RESET_B(net7),
    .Q(\next_state[4] ));
 sg13g2_dllrq_1 _925_ (.D(_439_),
    .GATE_N(_000_),
    .RESET_B(net8),
    .Q(\next_state[5] ));
 sg13g2_dfrbp_1 _926_ (.CLK(Hertz_60),
    .RESET_B(net144),
    .D(_033_),
    .Q_N(_033_),
    .Q(\display_sel[0] ));
 sg13g2_dfrbp_1 _927_ (.CLK(Hertz_60),
    .RESET_B(net144),
    .D(_031_),
    .Q_N(_441_),
    .Q(\display_sel[1] ));
 sg13g2_dfrbp_1 _928_ (.CLK(Hertz_60),
    .RESET_B(net144),
    .D(_032_),
    .Q_N(_001_),
    .Q(\display_sel[2] ));
 sg13g2_dfrbp_1 _929_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net149),
    .D(net21),
    .Q_N(_440_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 _930_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net149),
    .D(net51),
    .Q_N(_442_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 _931_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net149),
    .D(net65),
    .Q_N(_443_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 _932_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net149),
    .D(net33),
    .Q_N(_444_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 _933_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net149),
    .D(net42),
    .Q_N(_445_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 _934_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net148),
    .D(net38),
    .Q_N(_446_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 _935_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net148),
    .D(_027_),
    .Q_N(_447_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 _936_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net148),
    .D(net46),
    .Q_N(_448_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 _937_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net147),
    .D(_029_),
    .Q_N(_449_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 _938_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net147),
    .D(net48),
    .Q_N(_450_),
    .Q(\counter[9] ));
 sg13g2_dfrbp_1 _939_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net147),
    .D(net31),
    .Q_N(_451_),
    .Q(\counter[10] ));
 sg13g2_dfrbp_1 _940_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net145),
    .D(_008_),
    .Q_N(_452_),
    .Q(\counter[11] ));
 sg13g2_dfrbp_1 _941_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net145),
    .D(_009_),
    .Q_N(_453_),
    .Q(\counter[12] ));
 sg13g2_dfrbp_1 _942_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net145),
    .D(net28),
    .Q_N(_454_),
    .Q(\counter[13] ));
 sg13g2_dfrbp_1 _943_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net144),
    .D(net40),
    .Q_N(_455_),
    .Q(\counter[14] ));
 sg13g2_dfrbp_1 _944_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net144),
    .D(net36),
    .Q_N(_456_),
    .Q(\counter[15] ));
 sg13g2_dfrbp_1 _945_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net144),
    .D(_013_),
    .Q_N(_457_),
    .Q(\counter[16] ));
 sg13g2_dfrbp_1 _946_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net144),
    .D(net24),
    .Q_N(_458_),
    .Q(\counter[17] ));
 sg13g2_dfrbp_1 _947_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net145),
    .D(_015_),
    .Q_N(_459_),
    .Q(\counter[18] ));
 sg13g2_dfrbp_1 _948_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net145),
    .D(_016_),
    .Q_N(_460_),
    .Q(\counter[19] ));
 sg13g2_dfrbp_1 _949_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net145),
    .D(net26),
    .Q_N(_461_),
    .Q(\counter[20] ));
 sg13g2_dfrbp_1 _950_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net145),
    .D(net55),
    .Q_N(_462_),
    .Q(\counter[21] ));
 sg13g2_dfrbp_1 _951_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net145),
    .D(_020_),
    .Q_N(_463_),
    .Q(\counter[22] ));
 sg13g2_dfrbp_1 _952_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net147),
    .D(net44),
    .Q_N(_464_),
    .Q(\counter[23] ));
 sg13g2_dfrbp_1 _953_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net146),
    .D(net58),
    .Q_N(_465_),
    .Q(\counter[24] ));
 sg13g2_dfrbp_1 _954_ (.CLK(Hertz_4),
    .RESET_B(net148),
    .D(\next_state[0] ),
    .Q_N(_006_),
    .Q(\state[0] ));
 sg13g2_dfrbp_1 _955_ (.CLK(Hertz_4),
    .RESET_B(net148),
    .D(\next_state[1] ),
    .Q_N(_005_),
    .Q(\state[1] ));
 sg13g2_dfrbp_1 _956_ (.CLK(Hertz_4),
    .RESET_B(net146),
    .D(\next_state[2] ),
    .Q_N(_004_),
    .Q(\state[2] ));
 sg13g2_dfrbp_1 _957_ (.CLK(Hertz_4),
    .RESET_B(net148),
    .D(\next_state[3] ),
    .Q_N(_466_),
    .Q(\state[3] ));
 sg13g2_dfrbp_1 _958_ (.CLK(Hertz_4),
    .RESET_B(net148),
    .D(\next_state[4] ),
    .Q_N(_002_),
    .Q(\state[4] ));
 sg13g2_dfrbp_1 _959_ (.CLK(Hertz_4),
    .RESET_B(net148),
    .D(\next_state[5] ),
    .Q_N(_003_),
    .Q(\state[5] ));
 sg13g2_tiehi _921__4 (.L_HI(net4));
 sg13g2_tiehi _922__5 (.L_HI(net5));
 sg13g2_tiehi _923__6 (.L_HI(net6));
 sg13g2_tiehi _924__7 (.L_HI(net7));
 sg13g2_tiehi _925__8 (.L_HI(net8));
 sg13g2_tiehi tt_um_Esteban_Oman_Mendoza_maze_2024_top_9 (.L_HI(net9));
 sg13g2_tiehi tt_um_Esteban_Oman_Mendoza_maze_2024_top_10 (.L_HI(net10));
 sg13g2_tiehi tt_um_Esteban_Oman_Mendoza_maze_2024_top_11 (.L_HI(net11));
 sg13g2_tiehi tt_um_Esteban_Oman_Mendoza_maze_2024_top_12 (.L_HI(net12));
 sg13g2_tiehi tt_um_Esteban_Oman_Mendoza_maze_2024_top_13 (.L_HI(net13));
 sg13g2_tiehi tt_um_Esteban_Oman_Mendoza_maze_2024_top_14 (.L_HI(net14));
 sg13g2_tiehi tt_um_Esteban_Oman_Mendoza_maze_2024_top_15 (.L_HI(net15));
 sg13g2_tiehi tt_um_Esteban_Oman_Mendoza_maze_2024_top_16 (.L_HI(net16));
 sg13g2_tiehi tt_um_Esteban_Oman_Mendoza_maze_2024_top_17 (.L_HI(net17));
 sg13g2_tiehi tt_um_Esteban_Oman_Mendoza_maze_2024_top_18 (.L_HI(net18));
 sg13g2_tiehi tt_um_Esteban_Oman_Mendoza_maze_2024_top_19 (.L_HI(net19));
 sg13g2_tiehi tt_um_Esteban_Oman_Mendoza_maze_2024_top_20 (.L_HI(net20));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 fanout115 (.A(_260_),
    .X(net115));
 sg13g2_buf_4 fanout116 (.X(net116),
    .A(_133_));
 sg13g2_buf_4 fanout117 (.X(net117),
    .A(net118));
 sg13g2_buf_4 fanout118 (.X(net118),
    .A(_131_));
 sg13g2_buf_2 fanout119 (.A(net120),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_128_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_058_),
    .X(net121));
 sg13g2_buf_4 fanout122 (.X(net122),
    .A(_052_));
 sg13g2_buf_4 fanout123 (.X(net123),
    .A(_051_));
 sg13g2_buf_2 fanout124 (.A(\state[5] ),
    .X(net124));
 sg13g2_buf_1 fanout125 (.A(\state[5] ),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(\state[4] ),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(net129),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(net129),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(\state[3] ),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(net131),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(net132),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(\state[2] ),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(net134),
    .X(net133));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(\state[1] ));
 sg13g2_buf_2 fanout135 (.A(\state[0] ),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(\state[0] ),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_269_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_258_),
    .X(net138));
 sg13g2_buf_1 fanout139 (.A(_258_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(net2),
    .X(net140));
 sg13g2_buf_4 fanout141 (.X(net141),
    .A(net1));
 sg13g2_buf_4 fanout142 (.X(net142),
    .A(net143));
 sg13g2_buf_2 fanout143 (.A(ui_in[0]),
    .X(net143));
 sg13g2_buf_4 fanout144 (.X(net144),
    .A(net146));
 sg13g2_buf_4 fanout145 (.X(net145),
    .A(net146));
 sg13g2_buf_4 fanout146 (.X(net146),
    .A(net150));
 sg13g2_buf_2 fanout147 (.A(net150),
    .X(net147));
 sg13g2_buf_4 fanout148 (.X(net148),
    .A(net150));
 sg13g2_buf_4 fanout149 (.X(net149),
    .A(net150));
 sg13g2_buf_2 fanout150 (.A(rst_n),
    .X(net150));
 sg13g2_buf_1 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_tiehi _920__3 (.L_HI(net3));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_2_2__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_440_),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold2 (.A(\counter[17] ),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold3 (.A(_420_),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold4 (.A(_014_),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold5 (.A(\counter[20] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold6 (.A(_018_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold7 (.A(\counter[13] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold8 (.A(_010_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold9 (.A(\counter[10] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold10 (.A(_411_),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold11 (.A(_007_),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold12 (.A(\counter[3] ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold13 (.A(_024_),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold14 (.A(\counter[15] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold15 (.A(_417_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold16 (.A(_012_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold17 (.A(\counter[5] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold18 (.A(_026_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold19 (.A(\counter[14] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold20 (.A(_011_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold21 (.A(\counter[4] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold22 (.A(_025_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold23 (.A(\counter[23] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold24 (.A(_021_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold25 (.A(\counter[7] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold26 (.A(_028_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold27 (.A(\counter[9] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold28 (.A(_030_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold29 (.A(\counter[16] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold30 (.A(\counter[0] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold31 (.A(_017_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold32 (.A(\counter[18] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold33 (.A(\counter[11] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold34 (.A(\counter[21] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold35 (.A(_019_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold36 (.A(\counter[22] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold37 (.A(_426_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold38 (.A(_022_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold39 (.A(\counter[6] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold40 (.A(_407_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold41 (.A(\counter[8] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold42 (.A(\counter[19] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold43 (.A(\counter[2] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold44 (.A(_403_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold45 (.A(_023_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold46 (.A(\counter[12] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold47 (.A(\counter[11] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold48 (.A(_414_),
    .X(net68));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_4 FILLER_18_210 ();
 sg13g2_fill_2 FILLER_18_214 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_4 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_257 ();
 sg13g2_decap_8 FILLER_18_264 ();
 sg13g2_decap_8 FILLER_18_271 ();
 sg13g2_decap_8 FILLER_18_278 ();
 sg13g2_decap_8 FILLER_18_285 ();
 sg13g2_decap_8 FILLER_18_292 ();
 sg13g2_decap_8 FILLER_18_299 ();
 sg13g2_decap_8 FILLER_18_306 ();
 sg13g2_decap_8 FILLER_18_313 ();
 sg13g2_decap_8 FILLER_18_320 ();
 sg13g2_decap_8 FILLER_18_327 ();
 sg13g2_decap_8 FILLER_18_334 ();
 sg13g2_decap_8 FILLER_18_341 ();
 sg13g2_decap_8 FILLER_18_348 ();
 sg13g2_decap_8 FILLER_18_355 ();
 sg13g2_decap_8 FILLER_18_362 ();
 sg13g2_decap_8 FILLER_18_369 ();
 sg13g2_decap_8 FILLER_18_376 ();
 sg13g2_decap_8 FILLER_18_383 ();
 sg13g2_decap_8 FILLER_18_390 ();
 sg13g2_decap_8 FILLER_18_397 ();
 sg13g2_decap_4 FILLER_18_404 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_fill_1 FILLER_19_182 ();
 sg13g2_fill_1 FILLER_19_240 ();
 sg13g2_decap_8 FILLER_19_267 ();
 sg13g2_decap_8 FILLER_19_274 ();
 sg13g2_decap_8 FILLER_19_281 ();
 sg13g2_decap_8 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_295 ();
 sg13g2_decap_8 FILLER_19_302 ();
 sg13g2_decap_8 FILLER_19_309 ();
 sg13g2_decap_8 FILLER_19_316 ();
 sg13g2_decap_8 FILLER_19_323 ();
 sg13g2_decap_8 FILLER_19_330 ();
 sg13g2_decap_8 FILLER_19_337 ();
 sg13g2_decap_8 FILLER_19_344 ();
 sg13g2_decap_8 FILLER_19_351 ();
 sg13g2_decap_8 FILLER_19_358 ();
 sg13g2_decap_8 FILLER_19_365 ();
 sg13g2_decap_8 FILLER_19_372 ();
 sg13g2_decap_8 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_4 FILLER_20_91 ();
 sg13g2_fill_1 FILLER_20_95 ();
 sg13g2_decap_8 FILLER_20_104 ();
 sg13g2_decap_8 FILLER_20_111 ();
 sg13g2_decap_8 FILLER_20_118 ();
 sg13g2_decap_8 FILLER_20_125 ();
 sg13g2_decap_8 FILLER_20_132 ();
 sg13g2_decap_8 FILLER_20_139 ();
 sg13g2_decap_8 FILLER_20_146 ();
 sg13g2_decap_4 FILLER_20_153 ();
 sg13g2_fill_2 FILLER_20_157 ();
 sg13g2_decap_8 FILLER_20_167 ();
 sg13g2_decap_8 FILLER_20_174 ();
 sg13g2_fill_2 FILLER_20_181 ();
 sg13g2_decap_8 FILLER_20_191 ();
 sg13g2_fill_1 FILLER_20_198 ();
 sg13g2_fill_2 FILLER_20_251 ();
 sg13g2_decap_8 FILLER_20_279 ();
 sg13g2_decap_8 FILLER_20_286 ();
 sg13g2_decap_8 FILLER_20_293 ();
 sg13g2_decap_8 FILLER_20_300 ();
 sg13g2_decap_8 FILLER_20_307 ();
 sg13g2_decap_8 FILLER_20_314 ();
 sg13g2_decap_8 FILLER_20_321 ();
 sg13g2_decap_8 FILLER_20_328 ();
 sg13g2_decap_8 FILLER_20_335 ();
 sg13g2_decap_8 FILLER_20_342 ();
 sg13g2_decap_8 FILLER_20_349 ();
 sg13g2_decap_8 FILLER_20_356 ();
 sg13g2_decap_8 FILLER_20_363 ();
 sg13g2_decap_8 FILLER_20_370 ();
 sg13g2_decap_8 FILLER_20_377 ();
 sg13g2_decap_8 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_fill_2 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_117 ();
 sg13g2_decap_8 FILLER_21_124 ();
 sg13g2_decap_4 FILLER_21_131 ();
 sg13g2_fill_2 FILLER_21_135 ();
 sg13g2_decap_4 FILLER_21_150 ();
 sg13g2_fill_1 FILLER_21_154 ();
 sg13g2_decap_4 FILLER_21_181 ();
 sg13g2_fill_1 FILLER_21_185 ();
 sg13g2_fill_1 FILLER_21_198 ();
 sg13g2_decap_4 FILLER_21_215 ();
 sg13g2_decap_8 FILLER_21_281 ();
 sg13g2_decap_8 FILLER_21_288 ();
 sg13g2_decap_8 FILLER_21_295 ();
 sg13g2_decap_8 FILLER_21_302 ();
 sg13g2_decap_8 FILLER_21_309 ();
 sg13g2_decap_8 FILLER_21_316 ();
 sg13g2_decap_8 FILLER_21_323 ();
 sg13g2_decap_8 FILLER_21_330 ();
 sg13g2_decap_8 FILLER_21_337 ();
 sg13g2_decap_8 FILLER_21_344 ();
 sg13g2_decap_8 FILLER_21_351 ();
 sg13g2_decap_8 FILLER_21_358 ();
 sg13g2_decap_8 FILLER_21_365 ();
 sg13g2_decap_8 FILLER_21_372 ();
 sg13g2_decap_8 FILLER_21_379 ();
 sg13g2_decap_8 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_393 ();
 sg13g2_decap_8 FILLER_21_400 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_fill_2 FILLER_22_105 ();
 sg13g2_decap_4 FILLER_22_182 ();
 sg13g2_decap_4 FILLER_22_248 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_fill_2 FILLER_23_70 ();
 sg13g2_fill_1 FILLER_23_72 ();
 sg13g2_fill_1 FILLER_23_104 ();
 sg13g2_decap_4 FILLER_23_131 ();
 sg13g2_fill_1 FILLER_23_135 ();
 sg13g2_fill_1 FILLER_23_195 ();
 sg13g2_decap_8 FILLER_23_284 ();
 sg13g2_decap_8 FILLER_23_291 ();
 sg13g2_decap_8 FILLER_23_298 ();
 sg13g2_decap_8 FILLER_23_305 ();
 sg13g2_decap_8 FILLER_23_312 ();
 sg13g2_decap_8 FILLER_23_319 ();
 sg13g2_decap_8 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_333 ();
 sg13g2_decap_8 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_347 ();
 sg13g2_decap_8 FILLER_23_354 ();
 sg13g2_decap_8 FILLER_23_361 ();
 sg13g2_decap_8 FILLER_23_368 ();
 sg13g2_decap_8 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_fill_2 FILLER_24_63 ();
 sg13g2_fill_1 FILLER_24_65 ();
 sg13g2_fill_2 FILLER_24_82 ();
 sg13g2_fill_1 FILLER_24_84 ();
 sg13g2_fill_2 FILLER_24_94 ();
 sg13g2_fill_1 FILLER_24_96 ();
 sg13g2_decap_4 FILLER_24_114 ();
 sg13g2_fill_2 FILLER_24_144 ();
 sg13g2_fill_2 FILLER_24_189 ();
 sg13g2_fill_1 FILLER_24_191 ();
 sg13g2_fill_1 FILLER_24_201 ();
 sg13g2_fill_1 FILLER_24_223 ();
 sg13g2_decap_4 FILLER_24_250 ();
 sg13g2_decap_8 FILLER_24_285 ();
 sg13g2_decap_8 FILLER_24_292 ();
 sg13g2_fill_1 FILLER_24_299 ();
 sg13g2_decap_4 FILLER_24_305 ();
 sg13g2_fill_2 FILLER_24_309 ();
 sg13g2_decap_8 FILLER_24_327 ();
 sg13g2_decap_8 FILLER_24_334 ();
 sg13g2_decap_8 FILLER_24_341 ();
 sg13g2_decap_8 FILLER_24_348 ();
 sg13g2_decap_8 FILLER_24_355 ();
 sg13g2_decap_8 FILLER_24_362 ();
 sg13g2_decap_8 FILLER_24_369 ();
 sg13g2_decap_8 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_24_383 ();
 sg13g2_decap_8 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_fill_2 FILLER_25_63 ();
 sg13g2_fill_1 FILLER_25_99 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_fill_2 FILLER_25_245 ();
 sg13g2_fill_1 FILLER_25_247 ();
 sg13g2_decap_4 FILLER_25_274 ();
 sg13g2_fill_2 FILLER_25_278 ();
 sg13g2_decap_4 FILLER_25_358 ();
 sg13g2_fill_1 FILLER_25_362 ();
 sg13g2_decap_8 FILLER_25_379 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_4 FILLER_26_63 ();
 sg13g2_fill_1 FILLER_26_67 ();
 sg13g2_fill_2 FILLER_26_173 ();
 sg13g2_fill_1 FILLER_26_180 ();
 sg13g2_fill_1 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_198 ();
 sg13g2_fill_2 FILLER_26_205 ();
 sg13g2_decap_8 FILLER_26_212 ();
 sg13g2_decap_8 FILLER_26_219 ();
 sg13g2_decap_8 FILLER_26_226 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_254 ();
 sg13g2_decap_4 FILLER_26_261 ();
 sg13g2_fill_2 FILLER_26_265 ();
 sg13g2_decap_8 FILLER_26_272 ();
 sg13g2_fill_1 FILLER_26_279 ();
 sg13g2_decap_8 FILLER_26_286 ();
 sg13g2_decap_4 FILLER_26_293 ();
 sg13g2_fill_1 FILLER_26_297 ();
 sg13g2_fill_2 FILLER_26_303 ();
 sg13g2_fill_1 FILLER_26_305 ();
 sg13g2_decap_8 FILLER_26_312 ();
 sg13g2_decap_4 FILLER_26_319 ();
 sg13g2_fill_1 FILLER_26_323 ();
 sg13g2_decap_8 FILLER_26_328 ();
 sg13g2_decap_4 FILLER_26_335 ();
 sg13g2_decap_4 FILLER_26_343 ();
 sg13g2_fill_2 FILLER_26_347 ();
 sg13g2_fill_2 FILLER_26_362 ();
 sg13g2_decap_8 FILLER_26_388 ();
 sg13g2_decap_8 FILLER_26_395 ();
 sg13g2_decap_8 FILLER_26_402 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_fill_2 FILLER_27_70 ();
 sg13g2_fill_1 FILLER_27_127 ();
 sg13g2_fill_2 FILLER_27_186 ();
 sg13g2_decap_8 FILLER_27_202 ();
 sg13g2_decap_4 FILLER_27_209 ();
 sg13g2_fill_2 FILLER_27_213 ();
 sg13g2_fill_1 FILLER_27_223 ();
 sg13g2_decap_4 FILLER_27_250 ();
 sg13g2_fill_2 FILLER_27_254 ();
 sg13g2_fill_1 FILLER_27_271 ();
 sg13g2_fill_2 FILLER_27_294 ();
 sg13g2_decap_4 FILLER_27_318 ();
 sg13g2_fill_1 FILLER_27_347 ();
 sg13g2_fill_2 FILLER_27_357 ();
 sg13g2_fill_1 FILLER_27_359 ();
 sg13g2_fill_2 FILLER_27_372 ();
 sg13g2_decap_8 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_27_396 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_4 FILLER_28_63 ();
 sg13g2_fill_2 FILLER_28_120 ();
 sg13g2_decap_8 FILLER_28_172 ();
 sg13g2_decap_8 FILLER_28_179 ();
 sg13g2_fill_2 FILLER_28_186 ();
 sg13g2_fill_1 FILLER_28_188 ();
 sg13g2_decap_4 FILLER_28_194 ();
 sg13g2_fill_2 FILLER_28_198 ();
 sg13g2_decap_4 FILLER_28_212 ();
 sg13g2_fill_1 FILLER_28_216 ();
 sg13g2_decap_4 FILLER_28_223 ();
 sg13g2_fill_2 FILLER_28_247 ();
 sg13g2_fill_1 FILLER_28_249 ();
 sg13g2_decap_4 FILLER_28_263 ();
 sg13g2_decap_4 FILLER_28_278 ();
 sg13g2_fill_1 FILLER_28_282 ();
 sg13g2_decap_8 FILLER_28_291 ();
 sg13g2_decap_8 FILLER_28_298 ();
 sg13g2_fill_2 FILLER_28_305 ();
 sg13g2_decap_8 FILLER_28_312 ();
 sg13g2_decap_4 FILLER_28_319 ();
 sg13g2_fill_2 FILLER_28_323 ();
 sg13g2_decap_4 FILLER_28_343 ();
 sg13g2_decap_4 FILLER_28_356 ();
 sg13g2_fill_1 FILLER_28_360 ();
 sg13g2_decap_4 FILLER_28_365 ();
 sg13g2_fill_1 FILLER_28_369 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_4 FILLER_29_63 ();
 sg13g2_fill_2 FILLER_29_136 ();
 sg13g2_fill_2 FILLER_29_183 ();
 sg13g2_fill_2 FILLER_29_193 ();
 sg13g2_decap_8 FILLER_29_215 ();
 sg13g2_decap_4 FILLER_29_222 ();
 sg13g2_fill_1 FILLER_29_226 ();
 sg13g2_fill_2 FILLER_29_232 ();
 sg13g2_fill_1 FILLER_29_239 ();
 sg13g2_decap_4 FILLER_29_248 ();
 sg13g2_fill_2 FILLER_29_252 ();
 sg13g2_fill_2 FILLER_29_258 ();
 sg13g2_fill_2 FILLER_29_272 ();
 sg13g2_fill_1 FILLER_29_274 ();
 sg13g2_decap_4 FILLER_29_301 ();
 sg13g2_fill_1 FILLER_29_305 ();
 sg13g2_fill_1 FILLER_29_310 ();
 sg13g2_decap_8 FILLER_29_321 ();
 sg13g2_fill_1 FILLER_29_328 ();
 sg13g2_decap_8 FILLER_29_333 ();
 sg13g2_fill_2 FILLER_29_340 ();
 sg13g2_decap_4 FILLER_29_351 ();
 sg13g2_decap_4 FILLER_29_369 ();
 sg13g2_fill_1 FILLER_29_373 ();
 sg13g2_decap_8 FILLER_29_380 ();
 sg13g2_decap_8 FILLER_29_387 ();
 sg13g2_decap_8 FILLER_29_394 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_4 FILLER_30_63 ();
 sg13g2_fill_1 FILLER_30_137 ();
 sg13g2_decap_8 FILLER_30_144 ();
 sg13g2_fill_2 FILLER_30_151 ();
 sg13g2_fill_1 FILLER_30_153 ();
 sg13g2_decap_8 FILLER_30_173 ();
 sg13g2_fill_2 FILLER_30_180 ();
 sg13g2_fill_1 FILLER_30_203 ();
 sg13g2_fill_1 FILLER_30_226 ();
 sg13g2_fill_2 FILLER_30_240 ();
 sg13g2_fill_1 FILLER_30_242 ();
 sg13g2_fill_1 FILLER_30_251 ();
 sg13g2_fill_2 FILLER_30_258 ();
 sg13g2_decap_8 FILLER_30_277 ();
 sg13g2_decap_4 FILLER_30_290 ();
 sg13g2_decap_8 FILLER_30_298 ();
 sg13g2_fill_1 FILLER_30_359 ();
 sg13g2_fill_2 FILLER_30_365 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_4 FILLER_31_77 ();
 sg13g2_fill_2 FILLER_31_81 ();
 sg13g2_fill_1 FILLER_31_92 ();
 sg13g2_fill_2 FILLER_31_124 ();
 sg13g2_fill_1 FILLER_31_126 ();
 sg13g2_fill_2 FILLER_31_152 ();
 sg13g2_fill_2 FILLER_31_159 ();
 sg13g2_fill_1 FILLER_31_161 ();
 sg13g2_decap_4 FILLER_31_167 ();
 sg13g2_fill_2 FILLER_31_178 ();
 sg13g2_fill_2 FILLER_31_187 ();
 sg13g2_fill_2 FILLER_31_206 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_4 FILLER_31_246 ();
 sg13g2_fill_1 FILLER_31_250 ();
 sg13g2_fill_2 FILLER_31_258 ();
 sg13g2_fill_1 FILLER_31_260 ();
 sg13g2_fill_2 FILLER_31_305 ();
 sg13g2_fill_1 FILLER_31_307 ();
 sg13g2_fill_2 FILLER_31_320 ();
 sg13g2_fill_1 FILLER_31_322 ();
 sg13g2_decap_4 FILLER_31_333 ();
 sg13g2_fill_1 FILLER_31_337 ();
 sg13g2_decap_4 FILLER_31_343 ();
 sg13g2_fill_1 FILLER_31_347 ();
 sg13g2_decap_4 FILLER_31_352 ();
 sg13g2_fill_2 FILLER_31_356 ();
 sg13g2_decap_4 FILLER_31_368 ();
 sg13g2_fill_1 FILLER_31_372 ();
 sg13g2_decap_8 FILLER_31_386 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_fill_2 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_fill_1 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_128 ();
 sg13g2_fill_2 FILLER_32_159 ();
 sg13g2_fill_2 FILLER_32_193 ();
 sg13g2_fill_1 FILLER_32_195 ();
 sg13g2_fill_1 FILLER_32_202 ();
 sg13g2_fill_2 FILLER_32_208 ();
 sg13g2_fill_1 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_216 ();
 sg13g2_fill_2 FILLER_32_223 ();
 sg13g2_fill_2 FILLER_32_250 ();
 sg13g2_fill_1 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_272 ();
 sg13g2_fill_2 FILLER_32_279 ();
 sg13g2_fill_1 FILLER_32_291 ();
 sg13g2_decap_8 FILLER_32_304 ();
 sg13g2_decap_4 FILLER_32_330 ();
 sg13g2_fill_1 FILLER_32_334 ();
 sg13g2_fill_1 FILLER_32_340 ();
 sg13g2_fill_2 FILLER_32_362 ();
 sg13g2_fill_1 FILLER_32_390 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_fill_2 FILLER_33_91 ();
 sg13g2_fill_1 FILLER_33_93 ();
 sg13g2_decap_8 FILLER_33_120 ();
 sg13g2_decap_4 FILLER_33_127 ();
 sg13g2_fill_1 FILLER_33_131 ();
 sg13g2_fill_2 FILLER_33_138 ();
 sg13g2_decap_4 FILLER_33_154 ();
 sg13g2_decap_4 FILLER_33_162 ();
 sg13g2_fill_2 FILLER_33_171 ();
 sg13g2_fill_1 FILLER_33_178 ();
 sg13g2_decap_8 FILLER_33_183 ();
 sg13g2_decap_8 FILLER_33_220 ();
 sg13g2_fill_1 FILLER_33_227 ();
 sg13g2_decap_8 FILLER_33_242 ();
 sg13g2_decap_4 FILLER_33_257 ();
 sg13g2_fill_2 FILLER_33_279 ();
 sg13g2_fill_1 FILLER_33_281 ();
 sg13g2_decap_8 FILLER_33_288 ();
 sg13g2_fill_2 FILLER_33_295 ();
 sg13g2_fill_1 FILLER_33_297 ();
 sg13g2_fill_1 FILLER_33_302 ();
 sg13g2_decap_4 FILLER_33_312 ();
 sg13g2_fill_1 FILLER_33_316 ();
 sg13g2_fill_2 FILLER_33_338 ();
 sg13g2_fill_2 FILLER_33_371 ();
 sg13g2_fill_1 FILLER_33_373 ();
 sg13g2_fill_1 FILLER_33_384 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_4 FILLER_34_70 ();
 sg13g2_fill_2 FILLER_34_105 ();
 sg13g2_fill_1 FILLER_34_107 ();
 sg13g2_fill_2 FILLER_34_126 ();
 sg13g2_fill_1 FILLER_34_128 ();
 sg13g2_decap_4 FILLER_34_149 ();
 sg13g2_fill_1 FILLER_34_153 ();
 sg13g2_fill_2 FILLER_34_159 ();
 sg13g2_fill_2 FILLER_34_168 ();
 sg13g2_decap_4 FILLER_34_195 ();
 sg13g2_fill_1 FILLER_34_199 ();
 sg13g2_decap_8 FILLER_34_212 ();
 sg13g2_decap_8 FILLER_34_219 ();
 sg13g2_decap_4 FILLER_34_226 ();
 sg13g2_fill_1 FILLER_34_230 ();
 sg13g2_fill_2 FILLER_34_248 ();
 sg13g2_fill_1 FILLER_34_250 ();
 sg13g2_fill_2 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_272 ();
 sg13g2_fill_2 FILLER_34_279 ();
 sg13g2_decap_4 FILLER_34_317 ();
 sg13g2_fill_1 FILLER_34_321 ();
 sg13g2_decap_4 FILLER_34_349 ();
 sg13g2_fill_1 FILLER_34_353 ();
 sg13g2_decap_4 FILLER_34_359 ();
 sg13g2_decap_8 FILLER_34_368 ();
 sg13g2_fill_2 FILLER_34_375 ();
 sg13g2_fill_1 FILLER_34_377 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_4 FILLER_35_70 ();
 sg13g2_fill_1 FILLER_35_74 ();
 sg13g2_fill_2 FILLER_35_117 ();
 sg13g2_fill_1 FILLER_35_140 ();
 sg13g2_fill_2 FILLER_35_150 ();
 sg13g2_fill_2 FILLER_35_165 ();
 sg13g2_fill_2 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_194 ();
 sg13g2_fill_1 FILLER_35_211 ();
 sg13g2_decap_4 FILLER_35_220 ();
 sg13g2_fill_1 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_246 ();
 sg13g2_fill_2 FILLER_35_271 ();
 sg13g2_fill_1 FILLER_35_273 ();
 sg13g2_fill_1 FILLER_35_280 ();
 sg13g2_decap_4 FILLER_35_293 ();
 sg13g2_fill_2 FILLER_35_309 ();
 sg13g2_decap_4 FILLER_35_317 ();
 sg13g2_fill_1 FILLER_35_321 ();
 sg13g2_decap_8 FILLER_35_341 ();
 sg13g2_decap_4 FILLER_35_348 ();
 sg13g2_fill_1 FILLER_35_368 ();
 sg13g2_decap_8 FILLER_35_394 ();
 sg13g2_decap_8 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_fill_2 FILLER_36_99 ();
 sg13g2_fill_1 FILLER_36_101 ();
 sg13g2_decap_4 FILLER_36_106 ();
 sg13g2_fill_2 FILLER_36_110 ();
 sg13g2_decap_4 FILLER_36_132 ();
 sg13g2_decap_4 FILLER_36_150 ();
 sg13g2_fill_1 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_160 ();
 sg13g2_decap_8 FILLER_36_167 ();
 sg13g2_decap_4 FILLER_36_174 ();
 sg13g2_fill_2 FILLER_36_178 ();
 sg13g2_decap_4 FILLER_36_189 ();
 sg13g2_fill_2 FILLER_36_193 ();
 sg13g2_fill_2 FILLER_36_248 ();
 sg13g2_fill_2 FILLER_36_256 ();
 sg13g2_fill_1 FILLER_36_258 ();
 sg13g2_decap_8 FILLER_36_268 ();
 sg13g2_fill_2 FILLER_36_275 ();
 sg13g2_fill_1 FILLER_36_277 ();
 sg13g2_fill_2 FILLER_36_283 ();
 sg13g2_fill_1 FILLER_36_285 ();
 sg13g2_decap_4 FILLER_36_295 ();
 sg13g2_fill_2 FILLER_36_299 ();
 sg13g2_decap_8 FILLER_36_306 ();
 sg13g2_decap_4 FILLER_36_313 ();
 sg13g2_fill_2 FILLER_36_317 ();
 sg13g2_fill_1 FILLER_36_324 ();
 sg13g2_decap_4 FILLER_36_333 ();
 sg13g2_fill_1 FILLER_36_337 ();
 sg13g2_decap_4 FILLER_36_351 ();
 sg13g2_fill_2 FILLER_36_355 ();
 sg13g2_fill_1 FILLER_36_361 ();
 sg13g2_fill_2 FILLER_36_371 ();
 sg13g2_fill_1 FILLER_36_373 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_4 FILLER_37_175 ();
 sg13g2_fill_1 FILLER_37_179 ();
 sg13g2_fill_1 FILLER_37_224 ();
 sg13g2_fill_2 FILLER_37_240 ();
 sg13g2_fill_1 FILLER_37_242 ();
 sg13g2_decap_8 FILLER_37_271 ();
 sg13g2_decap_4 FILLER_37_278 ();
 sg13g2_decap_8 FILLER_37_286 ();
 sg13g2_decap_4 FILLER_37_293 ();
 sg13g2_fill_1 FILLER_37_297 ();
 sg13g2_fill_2 FILLER_37_358 ();
 sg13g2_fill_1 FILLER_37_367 ();
 sg13g2_decap_8 FILLER_37_383 ();
 sg13g2_decap_8 FILLER_37_390 ();
 sg13g2_decap_8 FILLER_37_397 ();
 sg13g2_decap_4 FILLER_37_404 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_fill_2 FILLER_38_182 ();
 sg13g2_fill_1 FILLER_38_184 ();
 sg13g2_decap_4 FILLER_38_193 ();
 sg13g2_fill_1 FILLER_38_197 ();
 sg13g2_decap_8 FILLER_38_202 ();
 sg13g2_decap_8 FILLER_38_209 ();
 sg13g2_fill_2 FILLER_38_216 ();
 sg13g2_fill_1 FILLER_38_218 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_decap_4 FILLER_38_229 ();
 sg13g2_decap_8 FILLER_38_253 ();
 sg13g2_decap_8 FILLER_38_260 ();
 sg13g2_decap_8 FILLER_38_267 ();
 sg13g2_decap_8 FILLER_38_274 ();
 sg13g2_decap_8 FILLER_38_281 ();
 sg13g2_decap_8 FILLER_38_288 ();
 sg13g2_decap_8 FILLER_38_295 ();
 sg13g2_decap_4 FILLER_38_302 ();
 sg13g2_decap_4 FILLER_38_317 ();
 sg13g2_decap_8 FILLER_38_341 ();
 sg13g2_fill_1 FILLER_38_348 ();
 sg13g2_decap_8 FILLER_38_370 ();
 sg13g2_decap_8 FILLER_38_377 ();
 sg13g2_decap_8 FILLER_38_384 ();
 sg13g2_decap_8 FILLER_38_391 ();
 sg13g2_decap_8 FILLER_38_398 ();
 sg13g2_decap_4 FILLER_38_405 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[5] = net17;
 assign uio_out[6] = net18;
 assign uio_out[7] = net19;
 assign uo_out[7] = net20;
endmodule

module tt_um_gamepad_pmod_demo (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire clknet_0_clk;
 wire \driver.decoder.data_reg[0] ;
 wire \driver.decoder.data_reg[10] ;
 wire \driver.decoder.data_reg[11] ;
 wire \driver.decoder.data_reg[1] ;
 wire \driver.decoder.data_reg[2] ;
 wire \driver.decoder.data_reg[3] ;
 wire \driver.decoder.data_reg[4] ;
 wire \driver.decoder.data_reg[5] ;
 wire \driver.decoder.data_reg[6] ;
 wire \driver.decoder.data_reg[7] ;
 wire \driver.decoder.data_reg[8] ;
 wire \driver.decoder.data_reg[9] ;
 wire \driver.driver.pmod_clk_prev ;
 wire \driver.driver.pmod_clk_sync[0] ;
 wire \driver.driver.pmod_clk_sync[1] ;
 wire \driver.driver.pmod_data_sync[0] ;
 wire \driver.driver.pmod_data_sync[1] ;
 wire \driver.driver.pmod_latch_prev ;
 wire \driver.driver.pmod_latch_sync[0] ;
 wire \driver.driver.pmod_latch_sync[1] ;
 wire \driver.driver.shift_reg[0] ;
 wire \driver.driver.shift_reg[10] ;
 wire \driver.driver.shift_reg[11] ;
 wire \driver.driver.shift_reg[1] ;
 wire \driver.driver.shift_reg[2] ;
 wire \driver.driver.shift_reg[3] ;
 wire \driver.driver.shift_reg[4] ;
 wire \driver.driver.shift_reg[5] ;
 wire \driver.driver.shift_reg[6] ;
 wire \driver.driver.shift_reg[7] ;
 wire \driver.driver.shift_reg[8] ;
 wire \driver.driver.shift_reg[9] ;
 wire hsync;
 wire \pix_x[0] ;
 wire \pix_x[1] ;
 wire \pix_x[2] ;
 wire \pix_x[3] ;
 wire \pix_x[4] ;
 wire \pix_x[5] ;
 wire \pix_x[6] ;
 wire \pix_x[7] ;
 wire \pix_x[8] ;
 wire \pix_x[9] ;
 wire \pix_y[0] ;
 wire \pix_y[1] ;
 wire \pix_y[2] ;
 wire \pix_y[3] ;
 wire \pix_y[4] ;
 wire \pix_y[5] ;
 wire \pix_y[6] ;
 wire \pix_y[7] ;
 wire \pix_y[8] ;
 wire \pix_y[9] ;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire \vga_sync_gen.vsync ;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;

 sg13g2_inv_1 _0579_ (.Y(_0070_),
    .A(net122));
 sg13g2_inv_1 _0580_ (.Y(_0071_),
    .A(net94));
 sg13g2_inv_1 _0581_ (.Y(_0072_),
    .A(net120));
 sg13g2_inv_1 _0582_ (.Y(_0073_),
    .A(net104));
 sg13g2_inv_1 _0583_ (.Y(_0074_),
    .A(net134));
 sg13g2_inv_1 _0584_ (.Y(_0075_),
    .A(net110));
 sg13g2_inv_1 _0585_ (.Y(_0076_),
    .A(net132));
 sg13g2_inv_1 _0586_ (.Y(_0077_),
    .A(net124));
 sg13g2_inv_1 _0587_ (.Y(_0078_),
    .A(net128));
 sg13g2_inv_1 _0588_ (.Y(_0079_),
    .A(net108));
 sg13g2_inv_1 _0589_ (.Y(_0080_),
    .A(\driver.driver.shift_reg[0] ));
 sg13g2_inv_1 _0590_ (.Y(_0081_),
    .A(net85));
 sg13g2_inv_1 _0591_ (.Y(_0082_),
    .A(net80));
 sg13g2_inv_1 _0592_ (.Y(_0083_),
    .A(net92));
 sg13g2_inv_1 _0593_ (.Y(_0084_),
    .A(net181));
 sg13g2_inv_1 _0594_ (.Y(_0085_),
    .A(\pix_y[6] ));
 sg13g2_inv_1 _0595_ (.Y(_0086_),
    .A(\pix_y[2] ));
 sg13g2_inv_1 _0596_ (.Y(_0087_),
    .A(net193));
 sg13g2_inv_1 _0597_ (.Y(_0088_),
    .A(\pix_x[4] ));
 sg13g2_inv_1 _0598_ (.Y(_0089_),
    .A(net197));
 sg13g2_inv_1 _0599_ (.Y(_0090_),
    .A(net198));
 sg13g2_inv_1 _0600_ (.Y(_0091_),
    .A(_0006_));
 sg13g2_inv_1 _0601_ (.Y(_0092_),
    .A(net211));
 sg13g2_inv_1 _0602_ (.Y(_0093_),
    .A(net98));
 sg13g2_inv_1 _0603_ (.Y(_0094_),
    .A(net114));
 sg13g2_inv_1 _0604_ (.Y(_0095_),
    .A(net118));
 sg13g2_inv_1 _0605_ (.Y(_0096_),
    .A(net116));
 sg13g2_inv_1 _0606_ (.Y(_0097_),
    .A(net90));
 sg13g2_inv_1 _0607_ (.Y(_0098_),
    .A(net100));
 sg13g2_inv_1 _0608_ (.Y(_0099_),
    .A(net102));
 sg13g2_inv_1 _0609_ (.Y(_0100_),
    .A(net96));
 sg13g2_inv_1 _0610_ (.Y(_0101_),
    .A(net106));
 sg13g2_inv_1 _0611_ (.Y(_0102_),
    .A(net130));
 sg13g2_inv_1 _0612_ (.Y(_0103_),
    .A(net126));
 sg13g2_inv_1 _0613_ (.Y(_0104_),
    .A(net112));
 sg13g2_and2_1 _0614_ (.A(\pix_y[7] ),
    .B(\pix_y[6] ),
    .X(_0105_));
 sg13g2_nand2_2 _0615_ (.Y(_0106_),
    .A(net182),
    .B(\pix_y[6] ));
 sg13g2_nand2b_1 _0616_ (.Y(_0107_),
    .B(net188),
    .A_N(net189));
 sg13g2_nand3b_1 _0617_ (.B(net193),
    .C(net184),
    .Y(_0108_),
    .A_N(net186));
 sg13g2_nand2b_1 _0618_ (.Y(_0109_),
    .B(net181),
    .A_N(\pix_y[9] ));
 sg13g2_nor4_2 _0619_ (.A(_0106_),
    .B(_0107_),
    .C(net208),
    .Y(_0001_),
    .D(_0109_));
 sg13g2_nor2_1 _0620_ (.A(net196),
    .B(\pix_x[5] ),
    .Y(_0110_));
 sg13g2_nor3_2 _0621_ (.A(\pix_x[6] ),
    .B(net196),
    .C(\pix_x[5] ),
    .Y(_0111_));
 sg13g2_nor2b_1 _0622_ (.A(\pix_x[8] ),
    .B_N(net151),
    .Y(_0112_));
 sg13g2_nand2b_1 _0623_ (.Y(_0113_),
    .B(net194),
    .A_N(\pix_x[8] ));
 sg13g2_nand2_1 _0624_ (.Y(_0114_),
    .A(net195),
    .B(net201));
 sg13g2_nand2_2 _0625_ (.Y(_0115_),
    .A(net196),
    .B(\pix_x[5] ));
 sg13g2_nand2_2 _0626_ (.Y(_0116_),
    .A(net195),
    .B(\pix_x[6] ));
 sg13g2_nor2_1 _0627_ (.A(_0115_),
    .B(_0116_),
    .Y(_0117_));
 sg13g2_nor3_1 _0628_ (.A(_0111_),
    .B(net202),
    .C(_0117_),
    .Y(_0000_));
 sg13g2_nor2_2 _0629_ (.A(\pix_x[7] ),
    .B(\pix_x[6] ),
    .Y(_0118_));
 sg13g2_nand2_1 _0630_ (.Y(_0119_),
    .A(_0110_),
    .B(_0118_));
 sg13g2_nor2b_1 _0631_ (.A(\pix_x[5] ),
    .B_N(net196),
    .Y(_0120_));
 sg13g2_and2_1 _0632_ (.A(_0118_),
    .B(_0120_),
    .X(_0121_));
 sg13g2_nand2_1 _0633_ (.Y(_0122_),
    .A(_0118_),
    .B(_0120_));
 sg13g2_nor2_1 _0634_ (.A(net136),
    .B(\pix_x[1] ),
    .Y(_0123_));
 sg13g2_nor3_1 _0635_ (.A(\pix_x[0] ),
    .B(\pix_x[2] ),
    .C(\pix_x[1] ),
    .Y(_0124_));
 sg13g2_and2_1 _0636_ (.A(\pix_x[3] ),
    .B(_0124_),
    .X(_0125_));
 sg13g2_nand2_1 _0637_ (.Y(_0126_),
    .A(\pix_x[3] ),
    .B(_0124_));
 sg13g2_a21oi_1 _0638_ (.A1(\pix_x[3] ),
    .A2(_0124_),
    .Y(_0127_),
    .B1(_0003_));
 sg13g2_o21ai_1 _0639_ (.B1(_0119_),
    .Y(_0128_),
    .A1(_0122_),
    .A2(_0127_));
 sg13g2_and2_2 _0640_ (.A(net184),
    .B(net185),
    .X(_0129_));
 sg13g2_nand2_2 _0641_ (.Y(_0130_),
    .A(net183),
    .B(net186));
 sg13g2_nor2_1 _0642_ (.A(net181),
    .B(\pix_y[9] ),
    .Y(_0131_));
 sg13g2_or2_1 _0643_ (.X(_0132_),
    .B(\pix_y[9] ),
    .A(net181));
 sg13g2_nand3_1 _0644_ (.B(_0129_),
    .C(_0131_),
    .A(_0105_),
    .Y(_0133_));
 sg13g2_nand2b_1 _0645_ (.Y(_0134_),
    .B(\pix_x[8] ),
    .A_N(net194));
 sg13g2_nor4_2 _0646_ (.A(_0106_),
    .B(_0130_),
    .C(_0132_),
    .Y(_0135_),
    .D(_0134_));
 sg13g2_nand2_1 _0647_ (.Y(_0136_),
    .A(_0121_),
    .B(_0125_));
 sg13g2_nor2_2 _0648_ (.A(\pix_x[8] ),
    .B(net194),
    .Y(_0137_));
 sg13g2_and3_1 _0649_ (.X(_0138_),
    .A(_0003_),
    .B(_0110_),
    .C(_0118_));
 sg13g2_o21ai_1 _0650_ (.B1(_0126_),
    .Y(_0139_),
    .A1(_0137_),
    .A2(_0138_));
 sg13g2_and4_2 _0651_ (.A(_0128_),
    .B(_0135_),
    .C(_0136_),
    .D(_0139_),
    .X(_0140_));
 sg13g2_or2_2 _0652_ (.X(_0141_),
    .B(net216),
    .A(net193));
 sg13g2_a21oi_1 _0653_ (.A1(net189),
    .A2(_0141_),
    .Y(_0142_),
    .B1(net188));
 sg13g2_nand3b_1 _0654_ (.B(\pix_y[6] ),
    .C(net184),
    .Y(_0143_),
    .A_N(\pix_y[7] ));
 sg13g2_nor2_1 _0655_ (.A(net185),
    .B(_0143_),
    .Y(_0144_));
 sg13g2_a21oi_1 _0656_ (.A1(\pix_y[6] ),
    .A2(_0091_),
    .Y(_0145_),
    .B1(\pix_y[7] ));
 sg13g2_a21o_1 _0657_ (.A2(_0144_),
    .A1(_0142_),
    .B1(_0145_),
    .X(_0146_));
 sg13g2_nor3_1 _0658_ (.A(_0086_),
    .B(net188),
    .C(_0141_),
    .Y(_0147_));
 sg13g2_nand2_1 _0659_ (.Y(_0148_),
    .A(_0144_),
    .B(_0147_));
 sg13g2_nand2_1 _0660_ (.Y(_0149_),
    .A(\pix_y[6] ),
    .B(_0129_));
 sg13g2_nor2_1 _0661_ (.A(net182),
    .B(_0132_),
    .Y(_0150_));
 sg13g2_o21ai_1 _0662_ (.B1(_0150_),
    .Y(_0151_),
    .A1(_0142_),
    .A2(_0149_));
 sg13g2_nor3_1 _0663_ (.A(net182),
    .B(_0085_),
    .C(_0130_),
    .Y(_0152_));
 sg13g2_a221oi_1 _0664_ (.B2(_0147_),
    .C1(_0151_),
    .B1(_0152_),
    .A1(_0146_),
    .Y(_0153_),
    .A2(_0148_));
 sg13g2_nor2b_2 _0665_ (.A(net196),
    .B_N(\pix_x[5] ),
    .Y(_0154_));
 sg13g2_nand2b_1 _0666_ (.Y(_0155_),
    .B(\pix_x[5] ),
    .A_N(net196));
 sg13g2_or4_1 _0667_ (.A(\pix_x[0] ),
    .B(net197),
    .C(\pix_x[2] ),
    .D(\pix_x[1] ),
    .X(_0156_));
 sg13g2_o21ai_1 _0668_ (.B1(_0007_),
    .Y(_0157_),
    .A1(_0155_),
    .A2(_0156_));
 sg13g2_and4_1 _0669_ (.A(_0115_),
    .B(_0118_),
    .C(_0137_),
    .D(_0157_),
    .X(_0158_));
 sg13g2_and2_2 _0670_ (.A(_0153_),
    .B(_0158_),
    .X(_0159_));
 sg13g2_nand2_2 _0671_ (.Y(_0160_),
    .A(_0153_),
    .B(_0158_));
 sg13g2_nor2b_1 _0672_ (.A(\pix_x[7] ),
    .B_N(\pix_x[6] ),
    .Y(_0161_));
 sg13g2_nand2_1 _0673_ (.Y(_0162_),
    .A(_0120_),
    .B(_0161_));
 sg13g2_nor2_1 _0674_ (.A(_0113_),
    .B(_0162_),
    .Y(_0163_));
 sg13g2_nand2_1 _0675_ (.Y(_0164_),
    .A(_0153_),
    .B(_0163_));
 sg13g2_o21ai_1 _0676_ (.B1(_0153_),
    .Y(_0165_),
    .A1(_0158_),
    .A2(_0163_));
 sg13g2_nand2_1 _0677_ (.Y(_0166_),
    .A(_0160_),
    .B(net164));
 sg13g2_xor2_1 _0678_ (.B(net187),
    .A(net185),
    .X(_0167_));
 sg13g2_nand2_1 _0679_ (.Y(_0168_),
    .A(net185),
    .B(net189));
 sg13g2_o21ai_1 _0680_ (.B1(_0168_),
    .Y(_0169_),
    .A1(net189),
    .A2(_0167_));
 sg13g2_nor2_1 _0681_ (.A(_0143_),
    .B(_0169_),
    .Y(_0170_));
 sg13g2_nand3b_1 _0682_ (.B(_0170_),
    .C(_0011_),
    .Y(_0171_),
    .A_N(net162));
 sg13g2_nor4_2 _0683_ (.A(net182),
    .B(\pix_y[6] ),
    .C(_0109_),
    .Y(_0172_),
    .D(_0129_));
 sg13g2_o21ai_1 _0684_ (.B1(_0008_),
    .Y(_0173_),
    .A1(_0107_),
    .A2(_0141_));
 sg13g2_mux2_1 _0685_ (.A0(net184),
    .A1(net185),
    .S(_0173_),
    .X(_0174_));
 sg13g2_and4_1 _0686_ (.A(_0115_),
    .B(_0137_),
    .C(_0157_),
    .D(_0161_),
    .X(_0175_));
 sg13g2_nand3_1 _0687_ (.B(_0174_),
    .C(_0175_),
    .A(_0172_),
    .Y(_0176_));
 sg13g2_nand2_1 _0688_ (.Y(_0177_),
    .A(_0112_),
    .B(_0118_));
 sg13g2_nor2_1 _0689_ (.A(_0113_),
    .B(_0119_),
    .Y(_0178_));
 sg13g2_and3_1 _0690_ (.X(_0179_),
    .A(_0172_),
    .B(_0174_),
    .C(_0178_));
 sg13g2_nand3_1 _0691_ (.B(_0174_),
    .C(_0178_),
    .A(_0172_),
    .Y(_0180_));
 sg13g2_a21oi_1 _0692_ (.A1(net168),
    .A2(_0180_),
    .Y(_0181_),
    .B1(_0167_));
 sg13g2_a21oi_1 _0693_ (.A1(net183),
    .A2(_0006_),
    .Y(_0182_),
    .B1(_0009_));
 sg13g2_a21o_1 _0694_ (.A2(_0129_),
    .A1(net188),
    .B1(_0182_),
    .X(_0183_));
 sg13g2_nand2_1 _0695_ (.Y(_0184_),
    .A(_0006_),
    .B(_0009_));
 sg13g2_a22oi_1 _0696_ (.Y(_0185_),
    .B1(_0184_),
    .B2(net183),
    .A2(net188),
    .A1(net186));
 sg13g2_nand2_1 _0697_ (.Y(_0186_),
    .A(_0011_),
    .B(_0012_));
 sg13g2_nor4_1 _0698_ (.A(_0084_),
    .B(_0183_),
    .C(_0185_),
    .D(_0186_),
    .Y(_0187_));
 sg13g2_nor3_2 _0699_ (.A(net183),
    .B(_0106_),
    .C(_0132_),
    .Y(_0188_));
 sg13g2_xor2_1 _0700_ (.B(_0173_),
    .A(net185),
    .X(_0189_));
 sg13g2_nand3_1 _0701_ (.B(_0188_),
    .C(_0189_),
    .A(_0175_),
    .Y(_0190_));
 sg13g2_and3_2 _0702_ (.X(_0191_),
    .A(_0178_),
    .B(_0188_),
    .C(_0189_));
 sg13g2_nand3_1 _0703_ (.B(_0188_),
    .C(_0189_),
    .A(_0178_),
    .Y(_0192_));
 sg13g2_nand2_1 _0704_ (.Y(_0193_),
    .A(net167),
    .B(net166));
 sg13g2_nand2_1 _0705_ (.Y(_0194_),
    .A(net181),
    .B(_0010_));
 sg13g2_xnor2_1 _0706_ (.Y(_0195_),
    .A(_0011_),
    .B(_0194_));
 sg13g2_nand4_1 _0707_ (.B(_0105_),
    .C(_0167_),
    .A(_0006_),
    .Y(_0196_),
    .D(_0195_));
 sg13g2_nor3_1 _0708_ (.A(net184),
    .B(net185),
    .C(net187),
    .Y(_0197_));
 sg13g2_xor2_1 _0709_ (.B(_0197_),
    .A(\pix_y[8] ),
    .X(_0198_));
 sg13g2_nor2_1 _0710_ (.A(_0196_),
    .B(_0198_),
    .Y(_0199_));
 sg13g2_nor2_1 _0711_ (.A(net181),
    .B(net182),
    .Y(_0200_));
 sg13g2_xnor2_1 _0712_ (.Y(_0201_),
    .A(net182),
    .B(net148));
 sg13g2_xnor2_1 _0713_ (.Y(_0202_),
    .A(\pix_y[9] ),
    .B(_0194_));
 sg13g2_or4_1 _0714_ (.A(_0149_),
    .B(_0200_),
    .C(_0201_),
    .D(_0202_),
    .X(_0203_));
 sg13g2_a21oi_1 _0715_ (.A1(\pix_y[8] ),
    .A2(_0105_),
    .Y(_0204_),
    .B1(_0203_));
 sg13g2_a221oi_1 _0716_ (.B2(_0199_),
    .C1(_0204_),
    .B1(_0193_),
    .A1(_0181_),
    .Y(_0205_),
    .A2(_0187_));
 sg13g2_nand2_1 _0717_ (.Y(_0206_),
    .A(_0171_),
    .B(net160));
 sg13g2_nand2_2 _0718_ (.Y(_0207_),
    .A(net169),
    .B(net167));
 sg13g2_and4_2 _0719_ (.A(_0105_),
    .B(_0129_),
    .C(_0131_),
    .D(_0137_),
    .X(_0208_));
 sg13g2_and3_1 _0720_ (.X(_0209_),
    .A(net195),
    .B(_0111_),
    .C(_0208_));
 sg13g2_nand3_1 _0721_ (.B(_0111_),
    .C(_0208_),
    .A(net195),
    .Y(_0210_));
 sg13g2_and2_1 _0722_ (.A(_0110_),
    .B(_0161_),
    .X(_0211_));
 sg13g2_and2_2 _0723_ (.A(_0208_),
    .B(_0211_),
    .X(_0212_));
 sg13g2_nand2_2 _0724_ (.Y(_0213_),
    .A(_0208_),
    .B(_0211_));
 sg13g2_nor2_1 _0725_ (.A(_0140_),
    .B(_0212_),
    .Y(_0214_));
 sg13g2_nor3_2 _0726_ (.A(_0133_),
    .B(_0155_),
    .C(_0177_),
    .Y(_0215_));
 sg13g2_nor2_2 _0727_ (.A(_0179_),
    .B(_0215_),
    .Y(_0216_));
 sg13g2_or2_1 _0728_ (.X(_0217_),
    .B(_0215_),
    .A(_0179_));
 sg13g2_nor2b_2 _0729_ (.A(_0116_),
    .B_N(_0135_),
    .Y(_0218_));
 sg13g2_and2_2 _0730_ (.A(_0154_),
    .B(_0218_),
    .X(_0219_));
 sg13g2_nand2_1 _0731_ (.Y(_0220_),
    .A(_0154_),
    .B(_0218_));
 sg13g2_nor2_2 _0732_ (.A(_0191_),
    .B(_0219_),
    .Y(_0221_));
 sg13g2_nand3_1 _0733_ (.B(_0216_),
    .C(_0221_),
    .A(_0164_),
    .Y(_0222_));
 sg13g2_nand3_1 _0734_ (.B(_0111_),
    .C(_0208_),
    .A(net195),
    .Y(_0223_));
 sg13g2_and2_1 _0735_ (.A(net167),
    .B(_0223_),
    .X(_0224_));
 sg13g2_nand3_1 _0736_ (.B(net167),
    .C(_0223_),
    .A(net168),
    .Y(_0225_));
 sg13g2_and4_1 _0737_ (.A(_0128_),
    .B(_0135_),
    .C(_0136_),
    .D(_0139_),
    .X(_0226_));
 sg13g2_or3_2 _0738_ (.A(_0212_),
    .B(_0225_),
    .C(_0226_),
    .X(_0227_));
 sg13g2_nor2_1 _0739_ (.A(_0159_),
    .B(_0227_),
    .Y(_0228_));
 sg13g2_or3_1 _0740_ (.A(_0133_),
    .B(_0155_),
    .C(_0177_),
    .X(_0229_));
 sg13g2_nand4_1 _0741_ (.B(\pix_x[6] ),
    .C(_0135_),
    .A(net195),
    .Y(_0230_),
    .D(_0154_));
 sg13g2_nand4_1 _0742_ (.B(net166),
    .C(_0220_),
    .A(_0180_),
    .Y(_0231_),
    .D(_0229_));
 sg13g2_or2_1 _0743_ (.X(_0232_),
    .B(_0231_),
    .A(_0225_));
 sg13g2_nand4_1 _0744_ (.B(_0135_),
    .C(_0136_),
    .A(_0128_),
    .Y(_0233_),
    .D(_0139_));
 sg13g2_nand2_1 _0745_ (.Y(_0234_),
    .A(_0213_),
    .B(_0233_));
 sg13g2_nor3_2 _0746_ (.A(_0225_),
    .B(_0231_),
    .C(_0234_),
    .Y(_0235_));
 sg13g2_nor4_1 _0747_ (.A(_0166_),
    .B(net160),
    .C(_0232_),
    .D(_0234_),
    .Y(_0236_));
 sg13g2_nand3b_1 _0748_ (.B(_0235_),
    .C(net163),
    .Y(_0237_),
    .A_N(net160));
 sg13g2_xor2_1 _0749_ (.B(net162),
    .A(_0013_),
    .X(_0238_));
 sg13g2_o21ai_1 _0750_ (.B1(_0086_),
    .Y(_0239_),
    .A1(_0225_),
    .A2(_0231_));
 sg13g2_mux2_1 _0751_ (.A0(_0238_),
    .A1(\pix_y[2] ),
    .S(_0232_),
    .X(_0240_));
 sg13g2_o21ai_1 _0752_ (.B1(_0239_),
    .Y(_0241_),
    .A1(_0232_),
    .A2(_0238_));
 sg13g2_a21oi_1 _0753_ (.A1(net190),
    .A2(_0237_),
    .Y(_0242_),
    .B1(net155));
 sg13g2_nand2_1 _0754_ (.Y(_0243_),
    .A(_0213_),
    .B(_0229_));
 sg13g2_nand4_1 _0755_ (.B(_0180_),
    .C(net167),
    .A(net168),
    .Y(_0244_),
    .D(net166));
 sg13g2_nand2_1 _0756_ (.Y(_0245_),
    .A(_0008_),
    .B(_0244_));
 sg13g2_o21ai_1 _0757_ (.B1(net187),
    .Y(_0246_),
    .A1(net189),
    .A2(net162));
 sg13g2_or3_1 _0758_ (.A(net189),
    .B(net187),
    .C(net162),
    .X(_0247_));
 sg13g2_a21o_1 _0759_ (.A2(_0247_),
    .A1(_0246_),
    .B1(_0244_),
    .X(_0248_));
 sg13g2_and2_1 _0760_ (.A(_0245_),
    .B(_0248_),
    .X(_0249_));
 sg13g2_nand2_1 _0761_ (.Y(_0250_),
    .A(_0245_),
    .B(_0248_));
 sg13g2_nor2_1 _0762_ (.A(_0140_),
    .B(_0159_),
    .Y(_0251_));
 sg13g2_nand2_1 _0763_ (.Y(_0252_),
    .A(_0216_),
    .B(_0251_));
 sg13g2_nand3_1 _0764_ (.B(_0216_),
    .C(_0251_),
    .A(net164),
    .Y(_0253_));
 sg13g2_nor2_1 _0765_ (.A(_0159_),
    .B(_0226_),
    .Y(_0254_));
 sg13g2_and3_1 _0766_ (.X(_0255_),
    .A(_0160_),
    .B(net161),
    .C(_0233_));
 sg13g2_and4_1 _0767_ (.A(_0160_),
    .B(net164),
    .C(net161),
    .D(_0233_),
    .X(_0256_));
 sg13g2_a22oi_1 _0768_ (.Y(_0257_),
    .B1(_0256_),
    .B2(net166),
    .A2(net160),
    .A1(_0171_));
 sg13g2_or2_1 _0769_ (.X(_0258_),
    .B(_0257_),
    .A(net190));
 sg13g2_a21oi_1 _0770_ (.A1(_0242_),
    .A2(_0258_),
    .Y(_0259_),
    .B1(net154));
 sg13g2_a21oi_2 _0771_ (.B1(net178),
    .Y(_0260_),
    .A2(net160),
    .A1(_0171_));
 sg13g2_a21oi_1 _0772_ (.A1(_0171_),
    .A2(net160),
    .Y(_0261_),
    .B1(net168));
 sg13g2_nor2_1 _0773_ (.A(_0179_),
    .B(_0243_),
    .Y(_0262_));
 sg13g2_nand2b_2 _0774_ (.Y(_0263_),
    .B(_0180_),
    .A_N(_0243_));
 sg13g2_and4_1 _0775_ (.A(net162),
    .B(net168),
    .C(_0213_),
    .D(net161),
    .X(_0264_));
 sg13g2_a21oi_1 _0776_ (.A1(_0171_),
    .A2(_0205_),
    .Y(_0265_),
    .B1(_0264_));
 sg13g2_a21o_1 _0777_ (.A2(_0260_),
    .A1(_0191_),
    .B1(_0265_),
    .X(_0266_));
 sg13g2_a22oi_1 _0778_ (.Y(_0267_),
    .B1(_0266_),
    .B2(net155),
    .A2(_0261_),
    .A1(_0242_));
 sg13g2_nand2b_1 _0779_ (.Y(_0268_),
    .B(_0169_),
    .A_N(net162));
 sg13g2_a21oi_1 _0780_ (.A1(_0014_),
    .A2(net162),
    .Y(_0269_),
    .B1(_0244_));
 sg13g2_a221oi_1 _0781_ (.B2(_0269_),
    .C1(_0181_),
    .B1(_0268_),
    .A1(_0167_),
    .Y(_0270_),
    .A2(_0193_));
 sg13g2_nor2_2 _0782_ (.A(\pix_x[1] ),
    .B(_0270_),
    .Y(_0271_));
 sg13g2_inv_1 _0783_ (.Y(_0272_),
    .A(_0271_));
 sg13g2_nand3_1 _0784_ (.B(net164),
    .C(_0262_),
    .A(net191),
    .Y(_0273_));
 sg13g2_and4_1 _0785_ (.A(net192),
    .B(_0160_),
    .C(net164),
    .D(_0262_),
    .X(_0274_));
 sg13g2_a21oi_1 _0786_ (.A1(_0224_),
    .A2(_0274_),
    .Y(_0275_),
    .B1(net156));
 sg13g2_nand2_1 _0787_ (.Y(_0276_),
    .A(net178),
    .B(net167));
 sg13g2_nor2_1 _0788_ (.A(_0263_),
    .B(_0276_),
    .Y(_0277_));
 sg13g2_nand2_2 _0789_ (.Y(_0278_),
    .A(net163),
    .B(_0221_));
 sg13g2_inv_1 _0790_ (.Y(_0279_),
    .A(_0278_));
 sg13g2_a221oi_1 _0791_ (.B2(_0279_),
    .C1(net156),
    .B1(_0277_),
    .A1(_0224_),
    .Y(_0280_),
    .A2(_0274_));
 sg13g2_nand2_1 _0792_ (.Y(_0281_),
    .A(net191),
    .B(_0190_));
 sg13g2_nor2_1 _0793_ (.A(_0231_),
    .B(_0281_),
    .Y(_0282_));
 sg13g2_and2_1 _0794_ (.A(net163),
    .B(_0214_),
    .X(_0283_));
 sg13g2_and3_1 _0795_ (.X(_0284_),
    .A(net179),
    .B(net164),
    .C(net161));
 sg13g2_a221oi_1 _0796_ (.B2(_0160_),
    .C1(net158),
    .B1(_0284_),
    .A1(_0282_),
    .Y(_0285_),
    .A2(_0283_));
 sg13g2_o21ai_1 _0797_ (.B1(_0206_),
    .Y(_0286_),
    .A1(_0280_),
    .A2(_0285_));
 sg13g2_nand2_1 _0798_ (.Y(_0287_),
    .A(net159),
    .B(_0271_));
 sg13g2_a221oi_1 _0799_ (.B2(net154),
    .C1(_0272_),
    .B1(_0286_),
    .A1(_0259_),
    .Y(_0288_),
    .A2(_0267_));
 sg13g2_nand2_1 _0800_ (.Y(_0289_),
    .A(_0192_),
    .B(_0210_));
 sg13g2_nand3_1 _0801_ (.B(_0223_),
    .C(_0274_),
    .A(net166),
    .Y(_0290_));
 sg13g2_nor4_1 _0802_ (.A(_0159_),
    .B(_0207_),
    .C(_0212_),
    .D(_0219_),
    .Y(_0291_));
 sg13g2_a21o_1 _0803_ (.A2(_0291_),
    .A1(_0180_),
    .B1(net192),
    .X(_0292_));
 sg13g2_a21o_1 _0804_ (.A2(_0292_),
    .A1(_0290_),
    .B1(net153),
    .X(_0293_));
 sg13g2_a21oi_1 _0805_ (.A1(_0223_),
    .A2(_0256_),
    .Y(_0294_),
    .B1(net190));
 sg13g2_nor2b_1 _0806_ (.A(_0294_),
    .B_N(_0254_),
    .Y(_0295_));
 sg13g2_a21oi_1 _0807_ (.A1(net153),
    .A2(_0295_),
    .Y(_0296_),
    .B1(net156));
 sg13g2_nor4_1 _0808_ (.A(net179),
    .B(_0207_),
    .C(_0212_),
    .D(_0278_),
    .Y(_0297_));
 sg13g2_a21oi_1 _0809_ (.A1(_0223_),
    .A2(_0255_),
    .Y(_0298_),
    .B1(net192));
 sg13g2_or3_1 _0810_ (.A(net153),
    .B(_0297_),
    .C(_0298_),
    .X(_0299_));
 sg13g2_nand3_1 _0811_ (.B(_0210_),
    .C(_0221_),
    .A(_0160_),
    .Y(_0300_));
 sg13g2_a21oi_1 _0812_ (.A1(net191),
    .A2(_0253_),
    .Y(_0301_),
    .B1(_0300_));
 sg13g2_a21oi_1 _0813_ (.A1(net152),
    .A2(_0301_),
    .Y(_0302_),
    .B1(net158));
 sg13g2_nor2b_2 _0814_ (.A(_0270_),
    .B_N(\pix_x[1] ),
    .Y(_0303_));
 sg13g2_nand2_1 _0815_ (.Y(_0304_),
    .A(net159),
    .B(_0303_));
 sg13g2_a221oi_1 _0816_ (.B2(_0302_),
    .C1(_0304_),
    .B1(_0299_),
    .A1(_0293_),
    .Y(_0305_),
    .A2(_0296_));
 sg13g2_or3_1 _0817_ (.A(_0090_),
    .B(_0288_),
    .C(_0305_),
    .X(_0306_));
 sg13g2_nand2_1 _0818_ (.Y(_0307_),
    .A(net178),
    .B(_0264_));
 sg13g2_nand2_1 _0819_ (.Y(_0308_),
    .A(net169),
    .B(_0251_));
 sg13g2_nand4_1 _0820_ (.B(net164),
    .C(net169),
    .A(net191),
    .Y(_0309_),
    .D(_0255_));
 sg13g2_nand3_1 _0821_ (.B(_0307_),
    .C(_0309_),
    .A(net156),
    .Y(_0310_));
 sg13g2_nor2_1 _0822_ (.A(net180),
    .B(_0191_),
    .Y(_0311_));
 sg13g2_nor3_1 _0823_ (.A(_0219_),
    .B(_0227_),
    .C(_0311_),
    .Y(_0312_));
 sg13g2_a21oi_1 _0824_ (.A1(net157),
    .A2(_0312_),
    .Y(_0313_),
    .B1(net153));
 sg13g2_nand2_1 _0825_ (.Y(_0314_),
    .A(net161),
    .B(_0283_));
 sg13g2_o21ai_1 _0826_ (.B1(_0275_),
    .Y(_0315_),
    .A1(_0276_),
    .A2(_0314_));
 sg13g2_nand2_1 _0827_ (.Y(_0316_),
    .A(net179),
    .B(_0180_));
 sg13g2_nor2_1 _0828_ (.A(_0278_),
    .B(_0316_),
    .Y(_0317_));
 sg13g2_nor3_1 _0829_ (.A(_0227_),
    .B(net157),
    .C(_0317_),
    .Y(_0318_));
 sg13g2_nor2_1 _0830_ (.A(_0250_),
    .B(_0318_),
    .Y(_0319_));
 sg13g2_a221oi_1 _0831_ (.B2(_0319_),
    .C1(_0304_),
    .B1(_0315_),
    .A1(_0310_),
    .Y(_0320_),
    .A2(_0313_));
 sg13g2_nor3_1 _0832_ (.A(_0191_),
    .B(_0219_),
    .C(_0316_),
    .Y(_0321_));
 sg13g2_and4_1 _0833_ (.A(net167),
    .B(_0210_),
    .C(_0213_),
    .D(_0229_),
    .X(_0322_));
 sg13g2_a22oi_1 _0834_ (.Y(_0323_),
    .B1(_0321_),
    .B2(_0322_),
    .A2(_0235_),
    .A1(net192));
 sg13g2_or2_1 _0835_ (.X(_0324_),
    .B(_0323_),
    .A(net154));
 sg13g2_nor2_1 _0836_ (.A(net190),
    .B(_0278_),
    .Y(_0325_));
 sg13g2_a21oi_1 _0837_ (.A1(net190),
    .A2(_0151_),
    .Y(_0326_),
    .B1(_0325_));
 sg13g2_a21oi_1 _0838_ (.A1(net154),
    .A2(_0326_),
    .Y(_0327_),
    .B1(net157));
 sg13g2_a21o_1 _0839_ (.A2(_0151_),
    .A1(net180),
    .B1(_0311_),
    .X(_0328_));
 sg13g2_nor2b_1 _0840_ (.A(_0231_),
    .B_N(net168),
    .Y(_0329_));
 sg13g2_a21oi_1 _0841_ (.A1(net190),
    .A2(_0329_),
    .Y(_0330_),
    .B1(_0235_));
 sg13g2_mux2_1 _0842_ (.A0(_0328_),
    .A1(_0330_),
    .S(net154),
    .X(_0331_));
 sg13g2_a221oi_1 _0843_ (.B2(net157),
    .C1(_0287_),
    .B1(_0331_),
    .A1(_0324_),
    .Y(_0332_),
    .A2(_0327_));
 sg13g2_or3_1 _0844_ (.A(net198),
    .B(_0320_),
    .C(_0332_),
    .X(_0333_));
 sg13g2_nand4_1 _0845_ (.B(net197),
    .C(_0306_),
    .A(_0088_),
    .Y(_0334_),
    .D(_0333_));
 sg13g2_nand2_1 _0846_ (.Y(_0335_),
    .A(net196),
    .B(_0089_));
 sg13g2_nor3_1 _0847_ (.A(_0225_),
    .B(_0263_),
    .C(_0278_),
    .Y(_0336_));
 sg13g2_a21o_1 _0848_ (.A2(_0336_),
    .A1(net159),
    .B1(net190),
    .X(_0337_));
 sg13g2_a21oi_1 _0849_ (.A1(net190),
    .A2(_0237_),
    .Y(_0338_),
    .B1(net157));
 sg13g2_nor3_1 _0850_ (.A(_0005_),
    .B(net166),
    .C(net155),
    .Y(_0339_));
 sg13g2_a221oi_1 _0851_ (.B2(net159),
    .C1(net154),
    .B1(_0339_),
    .A1(_0337_),
    .Y(_0340_),
    .A2(_0338_));
 sg13g2_nor2_1 _0852_ (.A(net191),
    .B(_0221_),
    .Y(_0341_));
 sg13g2_a21oi_1 _0853_ (.A1(net159),
    .A2(_0341_),
    .Y(_0342_),
    .B1(net157));
 sg13g2_nor3_1 _0854_ (.A(_0207_),
    .B(_0217_),
    .C(_0278_),
    .Y(_0343_));
 sg13g2_a221oi_1 _0855_ (.B2(_0343_),
    .C1(net155),
    .B1(_0260_),
    .A1(net178),
    .Y(_0344_),
    .A2(_0236_));
 sg13g2_o21ai_1 _0856_ (.B1(net152),
    .Y(_0345_),
    .A1(_0342_),
    .A2(_0344_));
 sg13g2_nand3b_1 _0857_ (.B(_0345_),
    .C(_0303_),
    .Y(_0346_),
    .A_N(_0340_));
 sg13g2_and3_1 _0858_ (.X(_0347_),
    .A(net168),
    .B(net161),
    .C(_0223_));
 sg13g2_a21oi_1 _0859_ (.A1(_0171_),
    .A2(net160),
    .Y(_0348_),
    .B1(_0347_));
 sg13g2_a221oi_1 _0860_ (.B2(net178),
    .C1(net157),
    .B1(_0348_),
    .A1(_0252_),
    .Y(_0349_),
    .A2(_0260_));
 sg13g2_nor3_1 _0861_ (.A(_0219_),
    .B(_0227_),
    .C(_0316_),
    .Y(_0350_));
 sg13g2_a221oi_1 _0862_ (.B2(net159),
    .C1(net155),
    .B1(_0350_),
    .A1(_0191_),
    .Y(_0351_),
    .A2(_0260_));
 sg13g2_o21ai_1 _0863_ (.B1(_0250_),
    .Y(_0352_),
    .A1(_0349_),
    .A2(_0351_));
 sg13g2_a221oi_1 _0864_ (.B2(_0206_),
    .C1(net157),
    .B1(_0341_),
    .A1(_0228_),
    .Y(_0353_),
    .A2(_0260_));
 sg13g2_nor2_1 _0865_ (.A(_0140_),
    .B(_0209_),
    .Y(_0354_));
 sg13g2_a22oi_1 _0866_ (.Y(_0355_),
    .B1(_0354_),
    .B2(_0284_),
    .A2(_0322_),
    .A1(net191));
 sg13g2_a21oi_1 _0867_ (.A1(net159),
    .A2(_0355_),
    .Y(_0356_),
    .B1(net155));
 sg13g2_o21ai_1 _0868_ (.B1(net152),
    .Y(_0357_),
    .A1(_0353_),
    .A2(_0356_));
 sg13g2_nand3_1 _0869_ (.B(_0352_),
    .C(_0357_),
    .A(_0271_),
    .Y(_0358_));
 sg13g2_nand3_1 _0870_ (.B(_0346_),
    .C(_0358_),
    .A(net198),
    .Y(_0359_));
 sg13g2_a22oi_1 _0871_ (.Y(_0360_),
    .B1(_0347_),
    .B2(net180),
    .A2(net160),
    .A1(_0171_));
 sg13g2_nand3_1 _0872_ (.B(net166),
    .C(_0347_),
    .A(net162),
    .Y(_0361_));
 sg13g2_and3_1 _0873_ (.X(_0362_),
    .A(net155),
    .B(_0360_),
    .C(_0361_));
 sg13g2_a221oi_1 _0874_ (.B2(_0242_),
    .C1(_0362_),
    .B1(_0258_),
    .A1(_0245_),
    .Y(_0363_),
    .A2(_0248_));
 sg13g2_o21ai_1 _0875_ (.B1(_0273_),
    .Y(_0364_),
    .A1(net191),
    .A2(_0222_));
 sg13g2_and3_1 _0876_ (.X(_0365_),
    .A(_0224_),
    .B(net158),
    .C(_0364_));
 sg13g2_nand4_1 _0877_ (.B(net161),
    .C(_0221_),
    .A(net164),
    .Y(_0366_),
    .D(_0354_));
 sg13g2_nor2b_1 _0878_ (.A(_0284_),
    .B_N(_0366_),
    .Y(_0367_));
 sg13g2_o21ai_1 _0879_ (.B1(net159),
    .Y(_0368_),
    .A1(net158),
    .A2(_0367_));
 sg13g2_o21ai_1 _0880_ (.B1(net152),
    .Y(_0369_),
    .A1(_0365_),
    .A2(_0368_));
 sg13g2_nand3b_1 _0881_ (.B(_0369_),
    .C(_0303_),
    .Y(_0370_),
    .A_N(_0363_));
 sg13g2_or2_1 _0882_ (.X(_0371_),
    .B(_0290_),
    .A(_0207_));
 sg13g2_nand4_1 _0883_ (.B(_0180_),
    .C(_0223_),
    .A(net168),
    .Y(_0372_),
    .D(_0230_));
 sg13g2_o21ai_1 _0884_ (.B1(net178),
    .Y(_0373_),
    .A1(_0166_),
    .A2(_0372_));
 sg13g2_a21o_1 _0885_ (.A2(_0373_),
    .A1(_0371_),
    .B1(net152),
    .X(_0374_));
 sg13g2_a21oi_1 _0886_ (.A1(net179),
    .A2(_0314_),
    .Y(_0375_),
    .B1(_0308_));
 sg13g2_a21oi_1 _0887_ (.A1(net152),
    .A2(_0375_),
    .Y(_0376_),
    .B1(net156));
 sg13g2_nand2_1 _0888_ (.Y(_0377_),
    .A(net166),
    .B(_0291_));
 sg13g2_nor2_1 _0889_ (.A(net178),
    .B(_0209_),
    .Y(_0378_));
 sg13g2_nand4_1 _0890_ (.B(net161),
    .C(_0221_),
    .A(net169),
    .Y(_0379_),
    .D(_0283_));
 sg13g2_a22oi_1 _0891_ (.Y(_0380_),
    .B1(_0378_),
    .B2(_0379_),
    .A2(_0377_),
    .A1(net178));
 sg13g2_and2_1 _0892_ (.A(_0254_),
    .B(_0277_),
    .X(_0381_));
 sg13g2_nand4_1 _0893_ (.B(net169),
    .C(_0210_),
    .A(net163),
    .Y(_0382_),
    .D(_0221_));
 sg13g2_a21oi_1 _0894_ (.A1(net191),
    .A2(_0382_),
    .Y(_0383_),
    .B1(_0381_));
 sg13g2_o21ai_1 _0895_ (.B1(net155),
    .Y(_0384_),
    .A1(net152),
    .A2(_0383_));
 sg13g2_a21oi_1 _0896_ (.A1(net152),
    .A2(_0380_),
    .Y(_0385_),
    .B1(_0384_));
 sg13g2_a21o_1 _0897_ (.A2(_0376_),
    .A1(_0374_),
    .B1(_0287_),
    .X(_0386_));
 sg13g2_o21ai_1 _0898_ (.B1(_0370_),
    .Y(_0387_),
    .A1(_0385_),
    .A2(_0386_));
 sg13g2_o21ai_1 _0899_ (.B1(_0359_),
    .Y(_0388_),
    .A1(net198),
    .A2(_0387_));
 sg13g2_a221oi_1 _0900_ (.B2(_0089_),
    .C1(_0092_),
    .B1(_0388_),
    .A1(_0334_),
    .Y(_0389_),
    .A2(_0335_));
 sg13g2_nand2_1 _0901_ (.Y(_0390_),
    .A(_0140_),
    .B(_0389_));
 sg13g2_nand3_1 _0902_ (.B(_0140_),
    .C(_0389_),
    .A(net106),
    .Y(_0391_));
 sg13g2_a21oi_1 _0903_ (.A1(_0306_),
    .A2(_0333_),
    .Y(_0392_),
    .B1(net197));
 sg13g2_a21oi_1 _0904_ (.A1(net197),
    .A2(_0388_),
    .Y(_0393_),
    .B1(_0392_));
 sg13g2_nor2_1 _0905_ (.A(_0100_),
    .B(net169),
    .Y(_0394_));
 sg13g2_a21oi_1 _0906_ (.A1(\driver.decoder.data_reg[10] ),
    .A2(_0218_),
    .Y(_0395_),
    .B1(_0394_));
 sg13g2_o21ai_1 _0907_ (.B1(_0395_),
    .Y(_0396_),
    .A1(_0099_),
    .A2(net167));
 sg13g2_a21o_1 _0908_ (.A2(_0159_),
    .A1(\driver.decoder.data_reg[1] ),
    .B1(_0396_),
    .X(_0397_));
 sg13g2_nor3_1 _0909_ (.A(\pix_x[5] ),
    .B(_0002_),
    .C(_0164_),
    .Y(_0398_));
 sg13g2_a22oi_1 _0910_ (.Y(_0399_),
    .B1(_0215_),
    .B2(\driver.decoder.data_reg[3] ),
    .A2(_0209_),
    .A1(\driver.decoder.data_reg[4] ));
 sg13g2_inv_1 _0911_ (.Y(_0400_),
    .A(_0399_));
 sg13g2_a221oi_1 _0912_ (.B2(\driver.decoder.data_reg[5] ),
    .C1(_0400_),
    .B1(_0212_),
    .A1(\driver.decoder.data_reg[2] ),
    .Y(_0401_),
    .A2(_0191_));
 sg13g2_o21ai_1 _0913_ (.B1(_0401_),
    .Y(_0402_),
    .A1(_0103_),
    .A2(_0180_));
 sg13g2_a221oi_1 _0914_ (.B2(net205),
    .C1(_0402_),
    .B1(_0398_),
    .A1(_0154_),
    .Y(_0403_),
    .A2(_0397_));
 sg13g2_nand2b_1 _0915_ (.Y(_0404_),
    .B(_0393_),
    .A_N(_0403_));
 sg13g2_nor2_1 _0916_ (.A(_0127_),
    .B(_0162_),
    .Y(_0405_));
 sg13g2_nor2_1 _0917_ (.A(_0211_),
    .B(_0405_),
    .Y(_0406_));
 sg13g2_o21ai_1 _0918_ (.B1(_0135_),
    .Y(_0407_),
    .A1(_0126_),
    .A2(_0162_));
 sg13g2_a21oi_1 _0919_ (.A1(_0003_),
    .A2(_0211_),
    .Y(_0408_),
    .B1(_0118_));
 sg13g2_nor2_1 _0920_ (.A(_0125_),
    .B(_0408_),
    .Y(_0409_));
 sg13g2_nor3_1 _0921_ (.A(_0406_),
    .B(_0407_),
    .C(_0409_),
    .Y(_0410_));
 sg13g2_nand3_1 _0922_ (.B(_0389_),
    .C(_0410_),
    .A(net130),
    .Y(_0411_));
 sg13g2_nand3_1 _0923_ (.B(_0404_),
    .C(_0411_),
    .A(_0391_),
    .Y(_0412_));
 sg13g2_nor4_2 _0924_ (.A(_0101_),
    .B(_0102_),
    .C(_0103_),
    .Y(_0413_),
    .D(_0104_));
 sg13g2_nand4_1 _0925_ (.B(net100),
    .C(net102),
    .A(net90),
    .Y(_0414_),
    .D(net96));
 sg13g2_nand3_1 _0926_ (.B(net114),
    .C(net118),
    .A(net98),
    .Y(_0415_));
 sg13g2_nor3_2 _0927_ (.A(_0096_),
    .B(_0414_),
    .C(_0415_),
    .Y(_0416_));
 sg13g2_nand2_1 _0928_ (.Y(_0417_),
    .A(_0413_),
    .B(_0416_));
 sg13g2_o21ai_1 _0929_ (.B1(_0154_),
    .Y(_0418_),
    .A1(_0159_),
    .A2(_0207_));
 sg13g2_nor4_1 _0930_ (.A(_0219_),
    .B(_0263_),
    .C(_0289_),
    .D(_0398_),
    .Y(_0419_));
 sg13g2_nand2_1 _0931_ (.Y(_0420_),
    .A(_0418_),
    .B(_0419_));
 sg13g2_a22oi_1 _0932_ (.Y(_0421_),
    .B1(_0420_),
    .B2(_0393_),
    .A2(_0410_),
    .A1(_0389_));
 sg13g2_nand3_1 _0933_ (.B(net183),
    .C(_0105_),
    .A(net181),
    .Y(_0422_));
 sg13g2_nand2_1 _0934_ (.Y(_0423_),
    .A(net206),
    .B(net194));
 sg13g2_nand2b_1 _0935_ (.Y(_0424_),
    .B(net199),
    .A_N(\pix_y[9] ));
 sg13g2_a21oi_1 _0936_ (.A1(net195),
    .A2(net194),
    .Y(_0425_),
    .B1(_0424_));
 sg13g2_nand3_1 _0937_ (.B(_0423_),
    .C(_0425_),
    .A(_0422_),
    .Y(_0426_));
 sg13g2_a221oi_1 _0938_ (.B2(_0390_),
    .C1(_0426_),
    .B1(_0421_),
    .A1(_0412_),
    .Y(_0017_),
    .A2(_0417_));
 sg13g2_nor2b_1 _0939_ (.A(\driver.driver.pmod_latch_prev ),
    .B_N(\driver.driver.pmod_latch_sync[1] ),
    .Y(_0427_));
 sg13g2_nor2b_1 _0940_ (.A(net176),
    .B_N(net200),
    .Y(_0428_));
 sg13g2_a22oi_1 _0941_ (.Y(_0018_),
    .B1(net173),
    .B2(_0094_),
    .A2(net177),
    .A1(_0080_));
 sg13g2_a22oi_1 _0942_ (.Y(_0019_),
    .B1(net172),
    .B2(_0093_),
    .A2(net177),
    .A1(_0079_));
 sg13g2_a22oi_1 _0943_ (.Y(_0020_),
    .B1(net172),
    .B2(_0096_),
    .A2(net176),
    .A1(_0078_));
 sg13g2_a22oi_1 _0944_ (.Y(_0021_),
    .B1(net173),
    .B2(_0095_),
    .A2(net177),
    .A1(_0077_));
 sg13g2_a22oi_1 _0945_ (.Y(_0022_),
    .B1(net173),
    .B2(_0098_),
    .A2(net177),
    .A1(_0076_));
 sg13g2_a22oi_1 _0946_ (.Y(_0023_),
    .B1(net173),
    .B2(_0097_),
    .A2(net177),
    .A1(_0075_));
 sg13g2_a22oi_1 _0947_ (.Y(_0024_),
    .B1(net172),
    .B2(_0100_),
    .A2(net176),
    .A1(_0074_));
 sg13g2_a22oi_1 _0948_ (.Y(_0025_),
    .B1(net172),
    .B2(_0099_),
    .A2(net176),
    .A1(_0073_));
 sg13g2_a22oi_1 _0949_ (.Y(_0026_),
    .B1(net172),
    .B2(_0102_),
    .A2(net176),
    .A1(_0072_));
 sg13g2_a22oi_1 _0950_ (.Y(_0027_),
    .B1(net172),
    .B2(_0101_),
    .A2(net176),
    .A1(_0071_));
 sg13g2_a22oi_1 _0951_ (.Y(_0028_),
    .B1(net172),
    .B2(_0104_),
    .A2(net176),
    .A1(_0070_));
 sg13g2_a22oi_1 _0952_ (.Y(_0029_),
    .B1(net172),
    .B2(_0103_),
    .A2(net176),
    .A1(_0083_));
 sg13g2_and2_2 _0953_ (.A(net136),
    .B(\pix_x[1] ),
    .X(_0429_));
 sg13g2_and3_1 _0954_ (.X(_0430_),
    .A(net197),
    .B(net198),
    .C(_0429_));
 sg13g2_nand3_1 _0955_ (.B(net198),
    .C(_0429_),
    .A(net197),
    .Y(_0431_));
 sg13g2_nand4_1 _0956_ (.B(net194),
    .C(_0121_),
    .A(\pix_x[8] ),
    .Y(_0432_),
    .D(_0430_));
 sg13g2_and2_2 _0957_ (.A(net199),
    .B(_0432_),
    .X(_0433_));
 sg13g2_nand2_1 _0958_ (.Y(_0434_),
    .A(net199),
    .B(_0432_));
 sg13g2_and2_1 _0959_ (.A(net79),
    .B(_0433_),
    .X(_0030_));
 sg13g2_nor3_1 _0960_ (.A(net137),
    .B(_0429_),
    .C(_0434_),
    .Y(_0031_));
 sg13g2_o21ai_1 _0961_ (.B1(net199),
    .Y(_0435_),
    .A1(net198),
    .A2(_0429_));
 sg13g2_a21oi_1 _0962_ (.A1(net198),
    .A2(_0429_),
    .Y(_0032_),
    .B1(_0435_));
 sg13g2_nor2b_1 _0963_ (.A(net87),
    .B_N(_0429_),
    .Y(_0436_));
 sg13g2_xnor2_1 _0964_ (.Y(_0437_),
    .A(net197),
    .B(_0436_));
 sg13g2_nor2_1 _0965_ (.A(_0434_),
    .B(net88),
    .Y(_0033_));
 sg13g2_xnor2_1 _0966_ (.Y(_0438_),
    .A(net89),
    .B(_0431_));
 sg13g2_nor2_1 _0967_ (.A(net165),
    .B(_0438_),
    .Y(_0034_));
 sg13g2_nor2_2 _0968_ (.A(_0115_),
    .B(_0431_),
    .Y(_0439_));
 sg13g2_a21oi_1 _0969_ (.A1(net196),
    .A2(_0430_),
    .Y(_0440_),
    .B1(net203));
 sg13g2_nor3_1 _0970_ (.A(net165),
    .B(_0439_),
    .C(net204),
    .Y(_0035_));
 sg13g2_o21ai_1 _0971_ (.B1(_0433_),
    .Y(_0441_),
    .A1(net210),
    .A2(_0439_));
 sg13g2_a21oi_1 _0972_ (.A1(net210),
    .A2(_0439_),
    .Y(_0036_),
    .B1(_0441_));
 sg13g2_a21oi_1 _0973_ (.A1(net210),
    .A2(_0439_),
    .Y(_0442_),
    .B1(net195));
 sg13g2_nor3_2 _0974_ (.A(_0115_),
    .B(_0116_),
    .C(_0431_),
    .Y(_0443_));
 sg13g2_nor3_1 _0975_ (.A(net165),
    .B(_0442_),
    .C(_0443_),
    .Y(_0037_));
 sg13g2_nor2_1 _0976_ (.A(net206),
    .B(_0443_),
    .Y(_0444_));
 sg13g2_and2_1 _0977_ (.A(net206),
    .B(_0443_),
    .X(_0445_));
 sg13g2_nor3_1 _0978_ (.A(net165),
    .B(_0444_),
    .C(_0445_),
    .Y(_0038_));
 sg13g2_a21oi_1 _0979_ (.A1(net194),
    .A2(_0445_),
    .Y(_0446_),
    .B1(net165));
 sg13g2_o21ai_1 _0980_ (.B1(_0446_),
    .Y(_0447_),
    .A1(net194),
    .A2(_0445_));
 sg13g2_inv_1 _0981_ (.Y(_0039_),
    .A(_0447_));
 sg13g2_a221oi_1 _0982_ (.B2(_0390_),
    .C1(_0426_),
    .B1(_0421_),
    .A1(_0413_),
    .Y(_0041_),
    .A2(_0416_));
 sg13g2_nor2b_1 _0983_ (.A(_0412_),
    .B_N(_0041_),
    .Y(_0040_));
 sg13g2_and2_1 _0984_ (.A(net200),
    .B(net1),
    .X(_0042_));
 sg13g2_and2_1 _0985_ (.A(net200),
    .B(net83),
    .X(_0043_));
 sg13g2_nand2_1 _0986_ (.Y(_0448_),
    .A(\pix_y[0] ),
    .B(_0433_));
 sg13g2_nor3_1 _0987_ (.A(\pix_y[8] ),
    .B(net183),
    .C(net185),
    .Y(_0449_));
 sg13g2_nor4_1 _0988_ (.A(net182),
    .B(\pix_y[6] ),
    .C(_0086_),
    .D(_0141_),
    .Y(_0450_));
 sg13g2_nand4_1 _0989_ (.B(net187),
    .C(_0449_),
    .A(\pix_y[9] ),
    .Y(_0451_),
    .D(_0450_));
 sg13g2_nand2_1 _0990_ (.Y(_0452_),
    .A(net199),
    .B(_0451_));
 sg13g2_or2_2 _0991_ (.X(_0453_),
    .B(_0452_),
    .A(_0432_));
 sg13g2_o21ai_1 _0992_ (.B1(_0448_),
    .Y(_0044_),
    .A1(_0082_),
    .A2(_0453_));
 sg13g2_nand2_1 _0993_ (.Y(_0454_),
    .A(net193),
    .B(net216));
 sg13g2_nand3b_1 _0994_ (.B(_0454_),
    .C(_0141_),
    .Y(_0455_),
    .A_N(_0453_));
 sg13g2_o21ai_1 _0995_ (.B1(_0455_),
    .Y(_0045_),
    .A1(net180),
    .A2(net165));
 sg13g2_nor2_1 _0996_ (.A(_0433_),
    .B(_0454_),
    .Y(_0456_));
 sg13g2_and2_2 _0997_ (.A(net165),
    .B(_0452_),
    .X(_0457_));
 sg13g2_xnor2_1 _0998_ (.Y(_0458_),
    .A(net189),
    .B(_0456_));
 sg13g2_nor2_1 _0999_ (.A(_0457_),
    .B(net217),
    .Y(_0046_));
 sg13g2_nand2_1 _1000_ (.Y(_0459_),
    .A(net187),
    .B(_0433_));
 sg13g2_nor2_1 _1001_ (.A(net144),
    .B(_0454_),
    .Y(_0460_));
 sg13g2_xnor2_1 _1002_ (.Y(_0461_),
    .A(net187),
    .B(net145));
 sg13g2_o21ai_1 _1003_ (.B1(_0459_),
    .Y(_0047_),
    .A1(_0453_),
    .A2(net146));
 sg13g2_nand4_1 _1004_ (.B(net187),
    .C(net193),
    .A(net189),
    .Y(_0462_),
    .D(\pix_y[0] ));
 sg13g2_nor2_1 _1005_ (.A(_0433_),
    .B(_0462_),
    .Y(_0463_));
 sg13g2_xnor2_1 _1006_ (.Y(_0464_),
    .A(net186),
    .B(_0463_));
 sg13g2_nor2_1 _1007_ (.A(_0457_),
    .B(net213),
    .Y(_0048_));
 sg13g2_nand2_1 _1008_ (.Y(_0465_),
    .A(net183),
    .B(_0433_));
 sg13g2_nor2_1 _1009_ (.A(net141),
    .B(_0462_),
    .Y(_0466_));
 sg13g2_xnor2_1 _1010_ (.Y(_0467_),
    .A(net183),
    .B(_0466_));
 sg13g2_o21ai_1 _1011_ (.B1(_0465_),
    .Y(_0049_),
    .A1(_0453_),
    .A2(net142));
 sg13g2_nor2_1 _1012_ (.A(_0130_),
    .B(_0462_),
    .Y(_0468_));
 sg13g2_nand2_1 _1013_ (.Y(_0469_),
    .A(net165),
    .B(_0468_));
 sg13g2_xnor2_1 _1014_ (.Y(_0470_),
    .A(_0085_),
    .B(_0469_));
 sg13g2_nor2_1 _1015_ (.A(_0457_),
    .B(_0470_),
    .Y(_0050_));
 sg13g2_nand3b_1 _1016_ (.B(_0469_),
    .C(net182),
    .Y(_0471_),
    .A_N(_0457_));
 sg13g2_nand2_1 _1017_ (.Y(_0472_),
    .A(_0201_),
    .B(_0468_));
 sg13g2_o21ai_1 _1018_ (.B1(_0471_),
    .Y(_0051_),
    .A1(_0453_),
    .A2(net149));
 sg13g2_nor2_1 _1019_ (.A(_0106_),
    .B(_0469_),
    .Y(_0473_));
 sg13g2_xnor2_1 _1020_ (.Y(_0474_),
    .A(net181),
    .B(_0473_));
 sg13g2_nor2_1 _1021_ (.A(_0457_),
    .B(_0474_),
    .Y(_0052_));
 sg13g2_nand2_1 _1022_ (.Y(_0475_),
    .A(\pix_y[9] ),
    .B(_0433_));
 sg13g2_nor4_1 _1023_ (.A(net138),
    .B(_0106_),
    .C(_0130_),
    .D(_0462_),
    .Y(_0476_));
 sg13g2_xnor2_1 _1024_ (.Y(_0477_),
    .A(\pix_y[9] ),
    .B(_0476_));
 sg13g2_o21ai_1 _1025_ (.B1(_0475_),
    .Y(_0053_),
    .A1(_0453_),
    .A2(net139));
 sg13g2_nor2b_1 _1026_ (.A(\driver.driver.pmod_clk_prev ),
    .B_N(\driver.driver.pmod_clk_sync[1] ),
    .Y(_0478_));
 sg13g2_nor2b_1 _1027_ (.A(net174),
    .B_N(net200),
    .Y(_0479_));
 sg13g2_a22oi_1 _1028_ (.Y(_0054_),
    .B1(net170),
    .B2(_0080_),
    .A2(net174),
    .A1(_0081_));
 sg13g2_a22oi_1 _1029_ (.Y(_0055_),
    .B1(net170),
    .B2(_0079_),
    .A2(net174),
    .A1(_0080_));
 sg13g2_a22oi_1 _1030_ (.Y(_0056_),
    .B1(net170),
    .B2(_0078_),
    .A2(net175),
    .A1(_0079_));
 sg13g2_a22oi_1 _1031_ (.Y(_0057_),
    .B1(net171),
    .B2(_0077_),
    .A2(net175),
    .A1(_0078_));
 sg13g2_a22oi_1 _1032_ (.Y(_0058_),
    .B1(net171),
    .B2(_0076_),
    .A2(net175),
    .A1(_0077_));
 sg13g2_a22oi_1 _1033_ (.Y(_0059_),
    .B1(net171),
    .B2(_0075_),
    .A2(net175),
    .A1(_0076_));
 sg13g2_a22oi_1 _1034_ (.Y(_0060_),
    .B1(net171),
    .B2(_0074_),
    .A2(net175),
    .A1(_0075_));
 sg13g2_a22oi_1 _1035_ (.Y(_0061_),
    .B1(net170),
    .B2(_0073_),
    .A2(net174),
    .A1(_0074_));
 sg13g2_a22oi_1 _1036_ (.Y(_0062_),
    .B1(net170),
    .B2(_0072_),
    .A2(net174),
    .A1(_0073_));
 sg13g2_a22oi_1 _1037_ (.Y(_0063_),
    .B1(net170),
    .B2(_0071_),
    .A2(net174),
    .A1(_0072_));
 sg13g2_a22oi_1 _1038_ (.Y(_0064_),
    .B1(net170),
    .B2(_0070_),
    .A2(net174),
    .A1(_0071_));
 sg13g2_a22oi_1 _1039_ (.Y(_0065_),
    .B1(net170),
    .B2(_0083_),
    .A2(net174),
    .A1(_0070_));
 sg13g2_and2_1 _1040_ (.A(net200),
    .B(net3),
    .X(_0066_));
 sg13g2_and2_1 _1041_ (.A(net199),
    .B(net84),
    .X(_0067_));
 sg13g2_and2_1 _1042_ (.A(net199),
    .B(net2),
    .X(_0068_));
 sg13g2_and2_1 _1043_ (.A(net199),
    .B(net82),
    .X(_0069_));
 sg13g2_dfrbp_1 _1044_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net47),
    .D(_0017_),
    .Q_N(_0518_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _1045_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net64),
    .D(net115),
    .Q_N(_0517_),
    .Q(\driver.decoder.data_reg[0] ));
 sg13g2_dfrbp_1 _1046_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net62),
    .D(net99),
    .Q_N(_0516_),
    .Q(\driver.decoder.data_reg[1] ));
 sg13g2_dfrbp_1 _1047_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net57),
    .D(net117),
    .Q_N(_0515_),
    .Q(\driver.decoder.data_reg[2] ));
 sg13g2_dfrbp_1 _1048_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net55),
    .D(net119),
    .Q_N(_0514_),
    .Q(\driver.decoder.data_reg[3] ));
 sg13g2_dfrbp_1 _1049_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net53),
    .D(net101),
    .Q_N(_0513_),
    .Q(\driver.decoder.data_reg[4] ));
 sg13g2_dfrbp_1 _1050_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net51),
    .D(net91),
    .Q_N(_0512_),
    .Q(\driver.decoder.data_reg[5] ));
 sg13g2_dfrbp_1 _1051_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net49),
    .D(net97),
    .Q_N(_0511_),
    .Q(\driver.decoder.data_reg[6] ));
 sg13g2_dfrbp_1 _1052_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net46),
    .D(net103),
    .Q_N(_0510_),
    .Q(\driver.decoder.data_reg[7] ));
 sg13g2_dfrbp_1 _1053_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net44),
    .D(net131),
    .Q_N(_0509_),
    .Q(\driver.decoder.data_reg[8] ));
 sg13g2_dfrbp_1 _1054_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net42),
    .D(net107),
    .Q_N(_0508_),
    .Q(\driver.decoder.data_reg[9] ));
 sg13g2_dfrbp_1 _1055_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net40),
    .D(net113),
    .Q_N(_0507_),
    .Q(\driver.decoder.data_reg[10] ));
 sg13g2_dfrbp_1 _1056_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net38),
    .D(net127),
    .Q_N(_0506_),
    .Q(\driver.decoder.data_reg[11] ));
 sg13g2_dfrbp_1 _1057_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net36),
    .D(_0030_),
    .Q_N(_0016_),
    .Q(\pix_x[0] ));
 sg13g2_dfrbp_1 _1058_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net35),
    .D(_0031_),
    .Q_N(_0505_),
    .Q(\pix_x[1] ));
 sg13g2_dfrbp_1 _1059_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net34),
    .D(_0032_),
    .Q_N(_0004_),
    .Q(\pix_x[2] ));
 sg13g2_dfrbp_1 _1060_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net33),
    .D(_0033_),
    .Q_N(_0003_),
    .Q(\pix_x[3] ));
 sg13g2_dfrbp_1 _1061_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net32),
    .D(_0034_),
    .Q_N(_0002_),
    .Q(\pix_x[4] ));
 sg13g2_dfrbp_1 _1062_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net31),
    .D(_0035_),
    .Q_N(_0007_),
    .Q(\pix_x[5] ));
 sg13g2_dfrbp_1 _1063_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net30),
    .D(_0036_),
    .Q_N(_0504_),
    .Q(\pix_x[6] ));
 sg13g2_dfrbp_1 _1064_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net29),
    .D(_0037_),
    .Q_N(_0503_),
    .Q(\pix_x[7] ));
 sg13g2_dfrbp_1 _1065_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net28),
    .D(_0038_),
    .Q_N(_0502_),
    .Q(\pix_x[8] ));
 sg13g2_dfrbp_1 _1066_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net27),
    .D(_0039_),
    .Q_N(_0501_),
    .Q(\pix_x[9] ));
 sg13g2_dfrbp_1 _1067_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net26),
    .D(_0040_),
    .Q_N(_0500_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _1068_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net25),
    .D(_0041_),
    .Q_N(_0499_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _1069_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net24),
    .D(_0042_),
    .Q_N(_0498_),
    .Q(\driver.driver.pmod_latch_sync[0] ));
 sg13g2_dfrbp_1 _1070_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net58),
    .D(_0043_),
    .Q_N(_0519_),
    .Q(\driver.driver.pmod_latch_sync[1] ));
 sg13g2_dfrbp_1 _1071_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net23),
    .D(_0000_),
    .Q_N(_0497_),
    .Q(hsync));
 sg13g2_dfrbp_1 _1072_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net22),
    .D(net81),
    .Q_N(_0015_),
    .Q(\pix_y[0] ));
 sg13g2_dfrbp_1 _1073_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net20),
    .D(_0045_),
    .Q_N(_0005_),
    .Q(\pix_y[1] ));
 sg13g2_dfrbp_1 _1074_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net75),
    .D(_0046_),
    .Q_N(_0013_),
    .Q(\pix_y[2] ));
 sg13g2_dfrbp_1 _1075_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net73),
    .D(net147),
    .Q_N(_0008_),
    .Q(\pix_y[3] ));
 sg13g2_dfrbp_1 _1076_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net71),
    .D(_0048_),
    .Q_N(_0014_),
    .Q(\pix_y[4] ));
 sg13g2_dfrbp_1 _1077_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net69),
    .D(net143),
    .Q_N(_0006_),
    .Q(\pix_y[5] ));
 sg13g2_dfrbp_1 _1078_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net67),
    .D(_0050_),
    .Q_N(_0009_),
    .Q(\pix_y[6] ));
 sg13g2_dfrbp_1 _1079_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net65),
    .D(net150),
    .Q_N(_0012_),
    .Q(\pix_y[7] ));
 sg13g2_dfrbp_1 _1080_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net61),
    .D(_0052_),
    .Q_N(_0010_),
    .Q(\pix_y[8] ));
 sg13g2_dfrbp_1 _1081_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net59),
    .D(net140),
    .Q_N(_0011_),
    .Q(\pix_y[9] ));
 sg13g2_dfrbp_1 _1082_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net60),
    .D(net209),
    .Q_N(_0520_),
    .Q(\vga_sync_gen.vsync ));
 sg13g2_dfrbp_1 _1083_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net66),
    .D(net77),
    .Q_N(_0521_),
    .Q(\driver.driver.pmod_clk_prev ));
 sg13g2_dfrbp_1 _1084_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net54),
    .D(net78),
    .Q_N(_0496_),
    .Q(\driver.driver.pmod_latch_prev ));
 sg13g2_dfrbp_1 _1085_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net50),
    .D(net86),
    .Q_N(_0495_),
    .Q(\driver.driver.shift_reg[0] ));
 sg13g2_dfrbp_1 _1086_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net45),
    .D(net109),
    .Q_N(_0494_),
    .Q(\driver.driver.shift_reg[1] ));
 sg13g2_dfrbp_1 _1087_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net41),
    .D(net129),
    .Q_N(_0493_),
    .Q(\driver.driver.shift_reg[2] ));
 sg13g2_dfrbp_1 _1088_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net37),
    .D(net125),
    .Q_N(_0492_),
    .Q(\driver.driver.shift_reg[3] ));
 sg13g2_dfrbp_1 _1089_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net76),
    .D(net133),
    .Q_N(_0491_),
    .Q(\driver.driver.shift_reg[4] ));
 sg13g2_dfrbp_1 _1090_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net72),
    .D(net111),
    .Q_N(_0490_),
    .Q(\driver.driver.shift_reg[5] ));
 sg13g2_dfrbp_1 _1091_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net68),
    .D(net135),
    .Q_N(_0489_),
    .Q(\driver.driver.shift_reg[6] ));
 sg13g2_dfrbp_1 _1092_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net63),
    .D(net105),
    .Q_N(_0488_),
    .Q(\driver.driver.shift_reg[7] ));
 sg13g2_dfrbp_1 _1093_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net52),
    .D(net121),
    .Q_N(_0487_),
    .Q(\driver.driver.shift_reg[8] ));
 sg13g2_dfrbp_1 _1094_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net43),
    .D(net95),
    .Q_N(_0486_),
    .Q(\driver.driver.shift_reg[9] ));
 sg13g2_dfrbp_1 _1095_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net21),
    .D(net123),
    .Q_N(_0485_),
    .Q(\driver.driver.shift_reg[10] ));
 sg13g2_dfrbp_1 _1096_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net70),
    .D(net93),
    .Q_N(_0484_),
    .Q(\driver.driver.shift_reg[11] ));
 sg13g2_dfrbp_1 _1097_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net56),
    .D(_0066_),
    .Q_N(_0483_),
    .Q(\driver.driver.pmod_data_sync[0] ));
 sg13g2_dfrbp_1 _1098_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net48),
    .D(_0067_),
    .Q_N(_0482_),
    .Q(\driver.driver.pmod_data_sync[1] ));
 sg13g2_dfrbp_1 _1099_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net39),
    .D(_0068_),
    .Q_N(_0481_),
    .Q(\driver.driver.pmod_clk_sync[0] ));
 sg13g2_dfrbp_1 _1100_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net74),
    .D(_0069_),
    .Q_N(_0480_),
    .Q(\driver.driver.pmod_clk_sync[1] ));
 sg13g2_tiehi _1095__21 (.L_HI(net21));
 sg13g2_tiehi _1072__22 (.L_HI(net22));
 sg13g2_tiehi _1071__23 (.L_HI(net23));
 sg13g2_tiehi _1069__24 (.L_HI(net24));
 sg13g2_tiehi _1068__25 (.L_HI(net25));
 sg13g2_tiehi _1067__26 (.L_HI(net26));
 sg13g2_tiehi _1066__27 (.L_HI(net27));
 sg13g2_tiehi _1065__28 (.L_HI(net28));
 sg13g2_tiehi _1064__29 (.L_HI(net29));
 sg13g2_tiehi _1063__30 (.L_HI(net30));
 sg13g2_tiehi _1062__31 (.L_HI(net31));
 sg13g2_tiehi _1061__32 (.L_HI(net32));
 sg13g2_tiehi _1060__33 (.L_HI(net33));
 sg13g2_tiehi _1059__34 (.L_HI(net34));
 sg13g2_tiehi _1058__35 (.L_HI(net35));
 sg13g2_tiehi _1057__36 (.L_HI(net36));
 sg13g2_tiehi _1088__37 (.L_HI(net37));
 sg13g2_tiehi _1056__38 (.L_HI(net38));
 sg13g2_tiehi _1099__39 (.L_HI(net39));
 sg13g2_tiehi _1055__40 (.L_HI(net40));
 sg13g2_tiehi _1087__41 (.L_HI(net41));
 sg13g2_tiehi _1054__42 (.L_HI(net42));
 sg13g2_tiehi _1094__43 (.L_HI(net43));
 sg13g2_tiehi _1053__44 (.L_HI(net44));
 sg13g2_tiehi _1086__45 (.L_HI(net45));
 sg13g2_tiehi _1052__46 (.L_HI(net46));
 sg13g2_tiehi _1044__47 (.L_HI(net47));
 sg13g2_tiehi _1098__48 (.L_HI(net48));
 sg13g2_tiehi _1051__49 (.L_HI(net49));
 sg13g2_tiehi _1085__50 (.L_HI(net50));
 sg13g2_tiehi _1050__51 (.L_HI(net51));
 sg13g2_tiehi _1093__52 (.L_HI(net52));
 sg13g2_tiehi _1049__53 (.L_HI(net53));
 sg13g2_tiehi _1084__54 (.L_HI(net54));
 sg13g2_tiehi _1048__55 (.L_HI(net55));
 sg13g2_tiehi _1097__56 (.L_HI(net56));
 sg13g2_tiehi _1047__57 (.L_HI(net57));
 sg13g2_tiehi _1070__58 (.L_HI(net58));
 sg13g2_tiehi _1081__59 (.L_HI(net59));
 sg13g2_tiehi _1082__60 (.L_HI(net60));
 sg13g2_tiehi _1080__61 (.L_HI(net61));
 sg13g2_tiehi _1046__62 (.L_HI(net62));
 sg13g2_tiehi _1092__63 (.L_HI(net63));
 sg13g2_tiehi _1045__64 (.L_HI(net64));
 sg13g2_tiehi _1079__65 (.L_HI(net65));
 sg13g2_tiehi _1083__66 (.L_HI(net66));
 sg13g2_tiehi _1078__67 (.L_HI(net67));
 sg13g2_tiehi _1091__68 (.L_HI(net68));
 sg13g2_tiehi _1077__69 (.L_HI(net69));
 sg13g2_tiehi _1096__70 (.L_HI(net70));
 sg13g2_tiehi _1076__71 (.L_HI(net71));
 sg13g2_tiehi _1090__72 (.L_HI(net72));
 sg13g2_tiehi _1075__73 (.L_HI(net73));
 sg13g2_tiehi _1100__74 (.L_HI(net74));
 sg13g2_tiehi _1074__75 (.L_HI(net75));
 sg13g2_tiehi _1089__76 (.L_HI(net76));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_gamepad_pmod_demo_5 (.L_LO(net5));
 sg13g2_tielo tt_um_gamepad_pmod_demo_6 (.L_LO(net6));
 sg13g2_tielo tt_um_gamepad_pmod_demo_7 (.L_LO(net7));
 sg13g2_tielo tt_um_gamepad_pmod_demo_8 (.L_LO(net8));
 sg13g2_tielo tt_um_gamepad_pmod_demo_9 (.L_LO(net9));
 sg13g2_tielo tt_um_gamepad_pmod_demo_10 (.L_LO(net10));
 sg13g2_tielo tt_um_gamepad_pmod_demo_11 (.L_LO(net11));
 sg13g2_tielo tt_um_gamepad_pmod_demo_12 (.L_LO(net12));
 sg13g2_tielo tt_um_gamepad_pmod_demo_13 (.L_LO(net13));
 sg13g2_tielo tt_um_gamepad_pmod_demo_14 (.L_LO(net14));
 sg13g2_tielo tt_um_gamepad_pmod_demo_15 (.L_LO(net15));
 sg13g2_tielo tt_um_gamepad_pmod_demo_16 (.L_LO(net16));
 sg13g2_tielo tt_um_gamepad_pmod_demo_17 (.L_LO(net17));
 sg13g2_tielo tt_um_gamepad_pmod_demo_18 (.L_LO(net18));
 sg13g2_tielo tt_um_gamepad_pmod_demo_19 (.L_LO(net19));
 sg13g2_tiehi _1073__20 (.L_HI(net20));
 sg13g2_buf_1 _1174_ (.A(uo_out[6]),
    .X(uo_out[0]));
 sg13g2_buf_1 _1175_ (.A(uo_out[5]),
    .X(uo_out[1]));
 sg13g2_buf_1 _1176_ (.A(uo_out[6]),
    .X(uo_out[2]));
 sg13g2_buf_1 _1177_ (.A(\vga_sync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _1178_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout152 (.A(net154),
    .X(net152));
 sg13g2_buf_1 fanout153 (.A(net154),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_0249_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_0241_),
    .X(net155));
 sg13g2_buf_1 fanout156 (.A(_0241_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_0240_),
    .X(net157));
 sg13g2_buf_1 fanout158 (.A(_0240_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_0206_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_0205_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_0216_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_0165_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_0165_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_0164_),
    .X(net164));
 sg13g2_buf_4 fanout165 (.X(net165),
    .A(_0434_));
 sg13g2_buf_2 fanout166 (.A(_0192_),
    .X(net166));
 sg13g2_buf_4 fanout167 (.X(net167),
    .A(_0190_));
 sg13g2_buf_2 fanout168 (.A(_0176_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_0176_),
    .X(net169));
 sg13g2_buf_4 fanout170 (.X(net170),
    .A(_0479_));
 sg13g2_buf_1 fanout171 (.A(_0479_),
    .X(net171));
 sg13g2_buf_4 fanout172 (.X(net172),
    .A(_0428_));
 sg13g2_buf_2 fanout173 (.A(_0428_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_0478_),
    .X(net174));
 sg13g2_buf_1 fanout175 (.A(_0478_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_0427_),
    .X(net176));
 sg13g2_buf_1 fanout177 (.A(_0427_),
    .X(net177));
 sg13g2_buf_4 fanout178 (.X(net178),
    .A(net180));
 sg13g2_buf_1 fanout179 (.A(net180),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_0087_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(net218),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(\pix_y[7] ),
    .X(net182));
 sg13g2_buf_4 fanout183 (.X(net183),
    .A(\pix_y[5] ));
 sg13g2_buf_1 fanout184 (.A(\pix_y[5] ),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(net186),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(net212),
    .X(net186));
 sg13g2_buf_4 fanout187 (.X(net187),
    .A(\pix_y[3] ));
 sg13g2_buf_1 fanout188 (.A(\pix_y[3] ),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(\pix_y[2] ),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(net192),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(net192),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(net193),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(net207),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(net151),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(net215),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(\pix_x[4] ),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(\pix_x[3] ),
    .X(net197));
 sg13g2_buf_4 fanout198 (.X(net198),
    .A(net214));
 sg13g2_buf_4 fanout199 (.X(net199),
    .A(rst_n));
 sg13g2_buf_1 fanout200 (.A(rst_n),
    .X(net200));
 sg13g2_buf_1 input1 (.A(ui_in[4]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[5]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[6]),
    .X(net3));
 sg13g2_tielo tt_um_gamepad_pmod_demo_4 (.L_LO(net4));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\driver.driver.pmod_clk_sync[1] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold2 (.A(\driver.driver.pmod_latch_sync[1] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0016_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0015_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0044_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold6 (.A(\driver.driver.pmod_clk_sync[0] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold7 (.A(\driver.driver.pmod_latch_sync[0] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold8 (.A(\driver.driver.pmod_data_sync[0] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold9 (.A(\driver.driver.pmod_data_sync[1] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0054_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0004_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0437_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0002_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold14 (.A(\driver.decoder.data_reg[5] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0023_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold16 (.A(\driver.driver.shift_reg[11] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0065_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold18 (.A(\driver.driver.shift_reg[9] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0063_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold20 (.A(\driver.decoder.data_reg[6] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0024_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold22 (.A(\driver.decoder.data_reg[1] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0019_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold24 (.A(\driver.decoder.data_reg[4] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0022_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold26 (.A(\driver.decoder.data_reg[7] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0025_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold28 (.A(\driver.driver.shift_reg[7] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0061_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold30 (.A(\driver.decoder.data_reg[9] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0027_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold32 (.A(\driver.driver.shift_reg[1] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0055_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold34 (.A(\driver.driver.shift_reg[5] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0059_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold36 (.A(\driver.decoder.data_reg[10] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0028_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold38 (.A(\driver.decoder.data_reg[0] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0018_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold40 (.A(\driver.decoder.data_reg[2] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0020_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold42 (.A(\driver.decoder.data_reg[3] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0021_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold44 (.A(\driver.driver.shift_reg[8] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0062_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold46 (.A(\driver.driver.shift_reg[10] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0064_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold48 (.A(\driver.driver.shift_reg[3] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0057_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold50 (.A(\driver.decoder.data_reg[11] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0029_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold52 (.A(\driver.driver.shift_reg[2] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0056_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold54 (.A(\driver.decoder.data_reg[8] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0026_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold56 (.A(\driver.driver.shift_reg[4] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0058_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold58 (.A(\driver.driver.shift_reg[6] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0060_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold60 (.A(\pix_x[0] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0123_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0010_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0477_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0053_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0014_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0467_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0049_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0013_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0460_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0461_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0047_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0009_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0472_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0051_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold75 (.A(\pix_x[9] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0112_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0114_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold78 (.A(\pix_x[5] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0440_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold80 (.A(\driver.decoder.data_reg[0] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold81 (.A(\pix_x[8] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold82 (.A(\pix_y[1] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0108_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0001_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold85 (.A(\pix_x[6] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0007_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold87 (.A(\pix_y[4] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0464_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold89 (.A(\pix_x[2] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold90 (.A(\pix_x[7] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold91 (.A(\pix_y[0] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0458_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold93 (.A(\pix_y[8] ),
    .X(net218));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_fill_1 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_97 ();
 sg13g2_decap_8 FILLER_17_104 ();
 sg13g2_decap_8 FILLER_17_111 ();
 sg13g2_decap_8 FILLER_17_118 ();
 sg13g2_decap_8 FILLER_17_125 ();
 sg13g2_decap_8 FILLER_17_132 ();
 sg13g2_decap_8 FILLER_17_139 ();
 sg13g2_decap_8 FILLER_17_146 ();
 sg13g2_decap_8 FILLER_17_153 ();
 sg13g2_decap_8 FILLER_17_160 ();
 sg13g2_decap_8 FILLER_17_167 ();
 sg13g2_decap_8 FILLER_17_174 ();
 sg13g2_decap_8 FILLER_17_181 ();
 sg13g2_decap_8 FILLER_17_188 ();
 sg13g2_decap_8 FILLER_17_195 ();
 sg13g2_decap_8 FILLER_17_202 ();
 sg13g2_decap_8 FILLER_17_209 ();
 sg13g2_decap_8 FILLER_17_216 ();
 sg13g2_decap_8 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_230 ();
 sg13g2_decap_8 FILLER_17_237 ();
 sg13g2_decap_8 FILLER_17_244 ();
 sg13g2_decap_8 FILLER_17_251 ();
 sg13g2_decap_8 FILLER_17_258 ();
 sg13g2_decap_8 FILLER_17_265 ();
 sg13g2_decap_8 FILLER_17_272 ();
 sg13g2_decap_8 FILLER_17_279 ();
 sg13g2_decap_8 FILLER_17_286 ();
 sg13g2_decap_8 FILLER_17_293 ();
 sg13g2_decap_8 FILLER_17_300 ();
 sg13g2_decap_8 FILLER_17_307 ();
 sg13g2_decap_8 FILLER_17_314 ();
 sg13g2_decap_8 FILLER_17_321 ();
 sg13g2_decap_8 FILLER_17_328 ();
 sg13g2_decap_8 FILLER_17_335 ();
 sg13g2_decap_8 FILLER_17_342 ();
 sg13g2_decap_8 FILLER_17_349 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_decap_8 FILLER_17_363 ();
 sg13g2_decap_8 FILLER_17_370 ();
 sg13g2_decap_8 FILLER_17_377 ();
 sg13g2_decap_8 FILLER_17_384 ();
 sg13g2_decap_8 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_17_398 ();
 sg13g2_decap_4 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_fill_1 FILLER_18_57 ();
 sg13g2_fill_2 FILLER_18_74 ();
 sg13g2_fill_1 FILLER_18_76 ();
 sg13g2_fill_2 FILLER_18_92 ();
 sg13g2_decap_4 FILLER_18_107 ();
 sg13g2_decap_8 FILLER_18_115 ();
 sg13g2_decap_8 FILLER_18_122 ();
 sg13g2_fill_1 FILLER_18_129 ();
 sg13g2_decap_8 FILLER_18_135 ();
 sg13g2_decap_4 FILLER_18_142 ();
 sg13g2_decap_4 FILLER_18_150 ();
 sg13g2_fill_2 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_166 ();
 sg13g2_decap_8 FILLER_18_173 ();
 sg13g2_decap_8 FILLER_18_180 ();
 sg13g2_decap_8 FILLER_18_187 ();
 sg13g2_decap_8 FILLER_18_199 ();
 sg13g2_decap_8 FILLER_18_206 ();
 sg13g2_fill_2 FILLER_18_213 ();
 sg13g2_fill_1 FILLER_18_219 ();
 sg13g2_fill_1 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_235 ();
 sg13g2_decap_8 FILLER_18_242 ();
 sg13g2_decap_8 FILLER_18_249 ();
 sg13g2_decap_8 FILLER_18_256 ();
 sg13g2_decap_8 FILLER_18_263 ();
 sg13g2_decap_8 FILLER_18_270 ();
 sg13g2_decap_8 FILLER_18_277 ();
 sg13g2_decap_8 FILLER_18_284 ();
 sg13g2_decap_8 FILLER_18_291 ();
 sg13g2_decap_8 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_305 ();
 sg13g2_decap_8 FILLER_18_312 ();
 sg13g2_decap_8 FILLER_18_319 ();
 sg13g2_decap_8 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_333 ();
 sg13g2_decap_8 FILLER_18_340 ();
 sg13g2_decap_8 FILLER_18_347 ();
 sg13g2_decap_8 FILLER_18_354 ();
 sg13g2_decap_8 FILLER_18_361 ();
 sg13g2_decap_8 FILLER_18_368 ();
 sg13g2_decap_8 FILLER_18_375 ();
 sg13g2_decap_8 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_18_389 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_4 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_fill_1 FILLER_19_68 ();
 sg13g2_fill_1 FILLER_19_126 ();
 sg13g2_fill_1 FILLER_19_170 ();
 sg13g2_fill_2 FILLER_19_176 ();
 sg13g2_fill_1 FILLER_19_178 ();
 sg13g2_fill_2 FILLER_19_187 ();
 sg13g2_fill_2 FILLER_19_240 ();
 sg13g2_decap_8 FILLER_19_251 ();
 sg13g2_decap_4 FILLER_19_258 ();
 sg13g2_fill_1 FILLER_19_262 ();
 sg13g2_decap_8 FILLER_19_268 ();
 sg13g2_decap_8 FILLER_19_275 ();
 sg13g2_decap_8 FILLER_19_282 ();
 sg13g2_decap_8 FILLER_19_289 ();
 sg13g2_decap_8 FILLER_19_296 ();
 sg13g2_decap_8 FILLER_19_303 ();
 sg13g2_decap_8 FILLER_19_310 ();
 sg13g2_decap_8 FILLER_19_317 ();
 sg13g2_decap_8 FILLER_19_324 ();
 sg13g2_decap_8 FILLER_19_331 ();
 sg13g2_decap_8 FILLER_19_338 ();
 sg13g2_decap_8 FILLER_19_345 ();
 sg13g2_decap_8 FILLER_19_352 ();
 sg13g2_decap_8 FILLER_19_359 ();
 sg13g2_decap_8 FILLER_19_366 ();
 sg13g2_decap_8 FILLER_19_373 ();
 sg13g2_decap_8 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_4 FILLER_20_32 ();
 sg13g2_fill_1 FILLER_20_36 ();
 sg13g2_fill_2 FILLER_20_125 ();
 sg13g2_decap_8 FILLER_20_150 ();
 sg13g2_fill_2 FILLER_20_157 ();
 sg13g2_fill_2 FILLER_20_164 ();
 sg13g2_fill_1 FILLER_20_179 ();
 sg13g2_decap_8 FILLER_20_200 ();
 sg13g2_decap_8 FILLER_20_207 ();
 sg13g2_decap_4 FILLER_20_214 ();
 sg13g2_fill_2 FILLER_20_218 ();
 sg13g2_decap_4 FILLER_20_234 ();
 sg13g2_fill_2 FILLER_20_247 ();
 sg13g2_fill_1 FILLER_20_258 ();
 sg13g2_decap_8 FILLER_20_275 ();
 sg13g2_decap_8 FILLER_20_282 ();
 sg13g2_decap_8 FILLER_20_289 ();
 sg13g2_decap_8 FILLER_20_296 ();
 sg13g2_decap_8 FILLER_20_303 ();
 sg13g2_decap_8 FILLER_20_310 ();
 sg13g2_decap_8 FILLER_20_317 ();
 sg13g2_decap_8 FILLER_20_324 ();
 sg13g2_decap_8 FILLER_20_331 ();
 sg13g2_decap_8 FILLER_20_338 ();
 sg13g2_decap_8 FILLER_20_345 ();
 sg13g2_decap_8 FILLER_20_352 ();
 sg13g2_decap_8 FILLER_20_359 ();
 sg13g2_decap_8 FILLER_20_366 ();
 sg13g2_decap_8 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_fill_2 FILLER_21_21 ();
 sg13g2_fill_1 FILLER_21_58 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_fill_1 FILLER_21_105 ();
 sg13g2_decap_4 FILLER_21_119 ();
 sg13g2_fill_1 FILLER_21_123 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_157 ();
 sg13g2_decap_4 FILLER_21_164 ();
 sg13g2_fill_2 FILLER_21_168 ();
 sg13g2_fill_2 FILLER_21_189 ();
 sg13g2_fill_1 FILLER_21_191 ();
 sg13g2_decap_8 FILLER_21_209 ();
 sg13g2_fill_1 FILLER_21_216 ();
 sg13g2_fill_2 FILLER_21_237 ();
 sg13g2_fill_1 FILLER_21_239 ();
 sg13g2_fill_2 FILLER_21_249 ();
 sg13g2_fill_1 FILLER_21_251 ();
 sg13g2_decap_4 FILLER_21_257 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_4 FILLER_22_21 ();
 sg13g2_fill_2 FILLER_22_25 ();
 sg13g2_fill_1 FILLER_22_44 ();
 sg13g2_fill_2 FILLER_22_68 ();
 sg13g2_decap_4 FILLER_22_74 ();
 sg13g2_fill_1 FILLER_22_90 ();
 sg13g2_fill_2 FILLER_22_108 ();
 sg13g2_decap_4 FILLER_22_123 ();
 sg13g2_fill_2 FILLER_22_127 ();
 sg13g2_decap_4 FILLER_22_134 ();
 sg13g2_fill_2 FILLER_22_169 ();
 sg13g2_fill_1 FILLER_22_189 ();
 sg13g2_fill_2 FILLER_22_207 ();
 sg13g2_fill_2 FILLER_22_216 ();
 sg13g2_decap_4 FILLER_22_228 ();
 sg13g2_fill_1 FILLER_22_232 ();
 sg13g2_fill_2 FILLER_22_241 ();
 sg13g2_decap_4 FILLER_22_248 ();
 sg13g2_fill_1 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_4 FILLER_23_21 ();
 sg13g2_fill_2 FILLER_23_25 ();
 sg13g2_fill_2 FILLER_23_35 ();
 sg13g2_fill_1 FILLER_23_45 ();
 sg13g2_decap_4 FILLER_23_76 ();
 sg13g2_fill_2 FILLER_23_85 ();
 sg13g2_fill_1 FILLER_23_93 ();
 sg13g2_fill_1 FILLER_23_121 ();
 sg13g2_decap_8 FILLER_23_146 ();
 sg13g2_fill_2 FILLER_23_153 ();
 sg13g2_fill_2 FILLER_23_189 ();
 sg13g2_fill_1 FILLER_23_191 ();
 sg13g2_decap_4 FILLER_23_207 ();
 sg13g2_fill_2 FILLER_23_235 ();
 sg13g2_decap_8 FILLER_23_257 ();
 sg13g2_decap_4 FILLER_23_269 ();
 sg13g2_decap_8 FILLER_23_290 ();
 sg13g2_decap_8 FILLER_23_297 ();
 sg13g2_decap_8 FILLER_23_304 ();
 sg13g2_decap_8 FILLER_23_311 ();
 sg13g2_decap_8 FILLER_23_318 ();
 sg13g2_decap_8 FILLER_23_325 ();
 sg13g2_decap_8 FILLER_23_332 ();
 sg13g2_decap_8 FILLER_23_339 ();
 sg13g2_decap_8 FILLER_23_346 ();
 sg13g2_decap_8 FILLER_23_353 ();
 sg13g2_decap_8 FILLER_23_360 ();
 sg13g2_decap_8 FILLER_23_367 ();
 sg13g2_decap_8 FILLER_23_374 ();
 sg13g2_decap_8 FILLER_23_381 ();
 sg13g2_decap_8 FILLER_23_388 ();
 sg13g2_decap_8 FILLER_23_395 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_4 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_18 ();
 sg13g2_fill_1 FILLER_24_80 ();
 sg13g2_fill_2 FILLER_24_94 ();
 sg13g2_decap_4 FILLER_24_123 ();
 sg13g2_fill_2 FILLER_24_127 ();
 sg13g2_fill_2 FILLER_24_158 ();
 sg13g2_fill_1 FILLER_24_160 ();
 sg13g2_fill_1 FILLER_24_165 ();
 sg13g2_fill_2 FILLER_24_181 ();
 sg13g2_decap_4 FILLER_24_187 ();
 sg13g2_fill_1 FILLER_24_191 ();
 sg13g2_fill_1 FILLER_24_197 ();
 sg13g2_decap_8 FILLER_24_216 ();
 sg13g2_fill_1 FILLER_24_223 ();
 sg13g2_decap_4 FILLER_24_229 ();
 sg13g2_decap_4 FILLER_24_254 ();
 sg13g2_fill_2 FILLER_24_258 ();
 sg13g2_fill_2 FILLER_24_265 ();
 sg13g2_decap_8 FILLER_24_289 ();
 sg13g2_decap_8 FILLER_24_296 ();
 sg13g2_decap_8 FILLER_24_303 ();
 sg13g2_decap_8 FILLER_24_310 ();
 sg13g2_decap_8 FILLER_24_317 ();
 sg13g2_decap_8 FILLER_24_324 ();
 sg13g2_decap_8 FILLER_24_331 ();
 sg13g2_decap_8 FILLER_24_338 ();
 sg13g2_decap_8 FILLER_24_345 ();
 sg13g2_decap_8 FILLER_24_352 ();
 sg13g2_decap_8 FILLER_24_359 ();
 sg13g2_decap_8 FILLER_24_366 ();
 sg13g2_decap_8 FILLER_24_373 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_fill_2 FILLER_25_28 ();
 sg13g2_fill_2 FILLER_25_38 ();
 sg13g2_fill_1 FILLER_25_94 ();
 sg13g2_fill_2 FILLER_25_105 ();
 sg13g2_fill_1 FILLER_25_107 ();
 sg13g2_decap_4 FILLER_25_118 ();
 sg13g2_decap_8 FILLER_25_137 ();
 sg13g2_decap_8 FILLER_25_144 ();
 sg13g2_decap_8 FILLER_25_151 ();
 sg13g2_fill_2 FILLER_25_158 ();
 sg13g2_decap_4 FILLER_25_165 ();
 sg13g2_fill_2 FILLER_25_169 ();
 sg13g2_fill_2 FILLER_25_177 ();
 sg13g2_fill_1 FILLER_25_184 ();
 sg13g2_fill_2 FILLER_25_197 ();
 sg13g2_fill_1 FILLER_25_199 ();
 sg13g2_decap_4 FILLER_25_215 ();
 sg13g2_fill_2 FILLER_25_219 ();
 sg13g2_decap_4 FILLER_25_239 ();
 sg13g2_decap_8 FILLER_25_289 ();
 sg13g2_decap_8 FILLER_25_296 ();
 sg13g2_decap_8 FILLER_25_303 ();
 sg13g2_decap_8 FILLER_25_310 ();
 sg13g2_decap_8 FILLER_25_317 ();
 sg13g2_decap_8 FILLER_25_324 ();
 sg13g2_decap_8 FILLER_25_331 ();
 sg13g2_decap_8 FILLER_25_338 ();
 sg13g2_decap_8 FILLER_25_345 ();
 sg13g2_decap_8 FILLER_25_352 ();
 sg13g2_decap_8 FILLER_25_359 ();
 sg13g2_decap_8 FILLER_25_366 ();
 sg13g2_fill_2 FILLER_25_373 ();
 sg13g2_fill_1 FILLER_25_375 ();
 sg13g2_decap_4 FILLER_25_380 ();
 sg13g2_fill_1 FILLER_25_384 ();
 sg13g2_decap_4 FILLER_25_389 ();
 sg13g2_fill_2 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_fill_1 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_4 FILLER_26_14 ();
 sg13g2_fill_1 FILLER_26_51 ();
 sg13g2_decap_8 FILLER_26_137 ();
 sg13g2_decap_8 FILLER_26_144 ();
 sg13g2_fill_1 FILLER_26_173 ();
 sg13g2_fill_2 FILLER_26_179 ();
 sg13g2_fill_1 FILLER_26_181 ();
 sg13g2_fill_1 FILLER_26_204 ();
 sg13g2_fill_1 FILLER_26_212 ();
 sg13g2_decap_4 FILLER_26_220 ();
 sg13g2_fill_1 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_234 ();
 sg13g2_decap_8 FILLER_26_241 ();
 sg13g2_fill_1 FILLER_26_253 ();
 sg13g2_fill_2 FILLER_26_259 ();
 sg13g2_fill_1 FILLER_26_269 ();
 sg13g2_decap_8 FILLER_26_282 ();
 sg13g2_decap_8 FILLER_26_289 ();
 sg13g2_decap_8 FILLER_26_296 ();
 sg13g2_decap_8 FILLER_26_303 ();
 sg13g2_decap_8 FILLER_26_310 ();
 sg13g2_fill_1 FILLER_26_317 ();
 sg13g2_decap_4 FILLER_26_321 ();
 sg13g2_fill_2 FILLER_26_328 ();
 sg13g2_fill_2 FILLER_26_336 ();
 sg13g2_fill_1 FILLER_26_352 ();
 sg13g2_fill_1 FILLER_26_357 ();
 sg13g2_fill_2 FILLER_26_365 ();
 sg13g2_fill_1 FILLER_26_370 ();
 sg13g2_fill_2 FILLER_26_381 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_83 ();
 sg13g2_decap_8 FILLER_27_90 ();
 sg13g2_fill_2 FILLER_27_97 ();
 sg13g2_decap_4 FILLER_27_108 ();
 sg13g2_fill_1 FILLER_27_112 ();
 sg13g2_fill_1 FILLER_27_117 ();
 sg13g2_decap_4 FILLER_27_123 ();
 sg13g2_fill_2 FILLER_27_127 ();
 sg13g2_decap_4 FILLER_27_137 ();
 sg13g2_decap_8 FILLER_27_167 ();
 sg13g2_decap_8 FILLER_27_190 ();
 sg13g2_decap_8 FILLER_27_197 ();
 sg13g2_fill_1 FILLER_27_204 ();
 sg13g2_decap_4 FILLER_27_208 ();
 sg13g2_fill_2 FILLER_27_212 ();
 sg13g2_fill_1 FILLER_27_240 ();
 sg13g2_fill_2 FILLER_27_246 ();
 sg13g2_fill_2 FILLER_27_269 ();
 sg13g2_decap_8 FILLER_27_286 ();
 sg13g2_fill_1 FILLER_27_293 ();
 sg13g2_fill_1 FILLER_27_301 ();
 sg13g2_fill_1 FILLER_27_345 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_4 FILLER_28_28 ();
 sg13g2_fill_2 FILLER_28_77 ();
 sg13g2_fill_2 FILLER_28_91 ();
 sg13g2_fill_1 FILLER_28_93 ();
 sg13g2_fill_1 FILLER_28_120 ();
 sg13g2_fill_2 FILLER_28_135 ();
 sg13g2_decap_4 FILLER_28_141 ();
 sg13g2_fill_2 FILLER_28_162 ();
 sg13g2_fill_1 FILLER_28_164 ();
 sg13g2_fill_2 FILLER_28_171 ();
 sg13g2_fill_1 FILLER_28_173 ();
 sg13g2_fill_2 FILLER_28_179 ();
 sg13g2_decap_4 FILLER_28_198 ();
 sg13g2_fill_1 FILLER_28_202 ();
 sg13g2_fill_2 FILLER_28_215 ();
 sg13g2_fill_1 FILLER_28_217 ();
 sg13g2_fill_2 FILLER_28_226 ();
 sg13g2_fill_2 FILLER_28_233 ();
 sg13g2_decap_4 FILLER_28_241 ();
 sg13g2_decap_4 FILLER_28_251 ();
 sg13g2_fill_1 FILLER_28_255 ();
 sg13g2_fill_2 FILLER_28_268 ();
 sg13g2_fill_1 FILLER_28_285 ();
 sg13g2_fill_1 FILLER_28_366 ();
 sg13g2_fill_1 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_fill_2 FILLER_29_42 ();
 sg13g2_fill_1 FILLER_29_44 ();
 sg13g2_fill_1 FILLER_29_80 ();
 sg13g2_fill_1 FILLER_29_87 ();
 sg13g2_decap_4 FILLER_29_92 ();
 sg13g2_fill_1 FILLER_29_96 ();
 sg13g2_fill_1 FILLER_29_107 ();
 sg13g2_fill_2 FILLER_29_113 ();
 sg13g2_fill_1 FILLER_29_126 ();
 sg13g2_decap_4 FILLER_29_148 ();
 sg13g2_fill_1 FILLER_29_152 ();
 sg13g2_fill_2 FILLER_29_160 ();
 sg13g2_fill_2 FILLER_29_176 ();
 sg13g2_fill_1 FILLER_29_178 ();
 sg13g2_decap_8 FILLER_29_183 ();
 sg13g2_fill_1 FILLER_29_190 ();
 sg13g2_fill_2 FILLER_29_204 ();
 sg13g2_decap_8 FILLER_29_246 ();
 sg13g2_decap_8 FILLER_29_253 ();
 sg13g2_fill_1 FILLER_29_279 ();
 sg13g2_fill_2 FILLER_29_301 ();
 sg13g2_fill_2 FILLER_29_398 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_fill_2 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_74 ();
 sg13g2_fill_2 FILLER_30_81 ();
 sg13g2_fill_1 FILLER_30_88 ();
 sg13g2_fill_1 FILLER_30_103 ();
 sg13g2_fill_2 FILLER_30_140 ();
 sg13g2_fill_1 FILLER_30_154 ();
 sg13g2_fill_2 FILLER_30_168 ();
 sg13g2_fill_1 FILLER_30_170 ();
 sg13g2_decap_4 FILLER_30_180 ();
 sg13g2_fill_2 FILLER_30_184 ();
 sg13g2_decap_4 FILLER_30_221 ();
 sg13g2_decap_4 FILLER_30_243 ();
 sg13g2_fill_1 FILLER_30_280 ();
 sg13g2_fill_1 FILLER_30_371 ();
 sg13g2_fill_2 FILLER_30_378 ();
 sg13g2_fill_2 FILLER_30_398 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_fill_2 FILLER_31_103 ();
 sg13g2_fill_1 FILLER_31_105 ();
 sg13g2_fill_2 FILLER_31_115 ();
 sg13g2_fill_1 FILLER_31_117 ();
 sg13g2_fill_1 FILLER_31_143 ();
 sg13g2_fill_1 FILLER_31_152 ();
 sg13g2_fill_1 FILLER_31_158 ();
 sg13g2_fill_2 FILLER_31_168 ();
 sg13g2_fill_1 FILLER_31_170 ();
 sg13g2_decap_8 FILLER_31_192 ();
 sg13g2_decap_8 FILLER_31_199 ();
 sg13g2_decap_8 FILLER_31_206 ();
 sg13g2_fill_2 FILLER_31_213 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_fill_2 FILLER_31_245 ();
 sg13g2_fill_1 FILLER_31_247 ();
 sg13g2_fill_1 FILLER_31_274 ();
 sg13g2_fill_1 FILLER_31_308 ();
 sg13g2_fill_2 FILLER_31_337 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_4 FILLER_32_28 ();
 sg13g2_fill_2 FILLER_32_32 ();
 sg13g2_fill_2 FILLER_32_79 ();
 sg13g2_fill_1 FILLER_32_95 ();
 sg13g2_fill_2 FILLER_32_152 ();
 sg13g2_fill_1 FILLER_32_154 ();
 sg13g2_fill_2 FILLER_32_187 ();
 sg13g2_fill_2 FILLER_32_230 ();
 sg13g2_fill_1 FILLER_32_232 ();
 sg13g2_fill_2 FILLER_32_238 ();
 sg13g2_fill_1 FILLER_32_316 ();
 sg13g2_fill_2 FILLER_32_326 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_4 FILLER_33_49 ();
 sg13g2_fill_2 FILLER_33_53 ();
 sg13g2_fill_1 FILLER_33_81 ();
 sg13g2_fill_1 FILLER_33_105 ();
 sg13g2_fill_2 FILLER_33_111 ();
 sg13g2_fill_1 FILLER_33_113 ();
 sg13g2_fill_1 FILLER_33_157 ();
 sg13g2_fill_2 FILLER_33_176 ();
 sg13g2_fill_2 FILLER_33_200 ();
 sg13g2_fill_1 FILLER_33_202 ();
 sg13g2_fill_2 FILLER_33_229 ();
 sg13g2_fill_1 FILLER_33_335 ();
 sg13g2_fill_2 FILLER_33_359 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_4 FILLER_34_67 ();
 sg13g2_fill_1 FILLER_34_71 ();
 sg13g2_fill_1 FILLER_34_115 ();
 sg13g2_fill_2 FILLER_34_140 ();
 sg13g2_decap_4 FILLER_34_184 ();
 sg13g2_fill_1 FILLER_34_196 ();
 sg13g2_fill_2 FILLER_34_210 ();
 sg13g2_fill_1 FILLER_34_298 ();
 sg13g2_fill_1 FILLER_34_325 ();
 sg13g2_fill_1 FILLER_34_340 ();
 sg13g2_fill_2 FILLER_34_367 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_fill_2 FILLER_35_84 ();
 sg13g2_fill_1 FILLER_35_86 ();
 sg13g2_fill_2 FILLER_35_117 ();
 sg13g2_fill_1 FILLER_35_119 ();
 sg13g2_fill_2 FILLER_35_146 ();
 sg13g2_fill_1 FILLER_35_148 ();
 sg13g2_decap_4 FILLER_35_184 ();
 sg13g2_fill_1 FILLER_35_188 ();
 sg13g2_decap_4 FILLER_35_218 ();
 sg13g2_decap_4 FILLER_35_226 ();
 sg13g2_fill_1 FILLER_35_230 ();
 sg13g2_decap_8 FILLER_35_235 ();
 sg13g2_fill_1 FILLER_35_312 ();
 sg13g2_fill_1 FILLER_35_322 ();
 sg13g2_fill_1 FILLER_35_328 ();
 sg13g2_fill_1 FILLER_35_337 ();
 sg13g2_fill_2 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_4 FILLER_36_98 ();
 sg13g2_fill_2 FILLER_36_106 ();
 sg13g2_fill_2 FILLER_36_116 ();
 sg13g2_fill_1 FILLER_36_118 ();
 sg13g2_fill_1 FILLER_36_137 ();
 sg13g2_decap_8 FILLER_36_197 ();
 sg13g2_decap_4 FILLER_36_204 ();
 sg13g2_fill_1 FILLER_36_208 ();
 sg13g2_fill_2 FILLER_36_244 ();
 sg13g2_fill_1 FILLER_36_246 ();
 sg13g2_fill_2 FILLER_36_284 ();
 sg13g2_fill_1 FILLER_36_341 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_4 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_162 ();
 sg13g2_decap_8 FILLER_37_169 ();
 sg13g2_fill_1 FILLER_37_176 ();
 sg13g2_decap_8 FILLER_37_181 ();
 sg13g2_decap_8 FILLER_37_188 ();
 sg13g2_decap_8 FILLER_37_195 ();
 sg13g2_decap_8 FILLER_37_202 ();
 sg13g2_decap_8 FILLER_37_209 ();
 sg13g2_decap_4 FILLER_37_216 ();
 sg13g2_fill_1 FILLER_37_220 ();
 sg13g2_fill_1 FILLER_37_247 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_fill_2 FILLER_38_222 ();
 sg13g2_fill_1 FILLER_38_224 ();
 sg13g2_fill_2 FILLER_38_229 ();
 sg13g2_fill_1 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_fill_1 FILLER_38_243 ();
 sg13g2_fill_1 FILLER_38_346 ();
 sg13g2_fill_1 FILLER_38_373 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net4;
 assign uio_oe[1] = net5;
 assign uio_oe[2] = net6;
 assign uio_oe[3] = net7;
 assign uio_oe[4] = net8;
 assign uio_oe[5] = net9;
 assign uio_oe[6] = net10;
 assign uio_oe[7] = net11;
 assign uio_out[0] = net12;
 assign uio_out[1] = net13;
 assign uio_out[2] = net14;
 assign uio_out[3] = net15;
 assign uio_out[4] = net16;
 assign uio_out[5] = net17;
 assign uio_out[6] = net18;
 assign uio_out[7] = net19;
endmodule

module tt_um_pyamnihc_dummy_counter (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire count_en_db_r;
 wire \count_en_p[0] ;
 wire \count_en_p[1] ;
 wire \count_en_p[2] ;
 wire \count_en_p[3] ;
 wire count_en_r;
 wire \counter_db_r[0] ;
 wire \counter_db_r[1] ;
 wire \counter_db_r[2] ;
 wire \counter_db_r[3] ;
 wire \counter_r[0] ;
 wire \counter_r[10] ;
 wire \counter_r[11] ;
 wire \counter_r[12] ;
 wire \counter_r[13] ;
 wire \counter_r[14] ;
 wire \counter_r[15] ;
 wire \counter_r[1] ;
 wire \counter_r[2] ;
 wire \counter_r[3] ;
 wire \counter_r[4] ;
 wire \counter_r[5] ;
 wire \counter_r[6] ;
 wire \counter_r[7] ;
 wire \counter_r[8] ;
 wire \counter_r[9] ;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire clknet_0_clk;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;

 sg13g2_inv_1 _0490_ (.Y(_0439_),
    .A(net114));
 sg13g2_inv_1 _0491_ (.Y(_0440_),
    .A(\counter_r[2] ));
 sg13g2_inv_1 _0492_ (.Y(_0441_),
    .A(net36));
 sg13g2_and2_2 _0493_ (.A(net5),
    .B(net2),
    .X(_0442_));
 sg13g2_nand2_1 _0494_ (.Y(_0443_),
    .A(net5),
    .B(net2));
 sg13g2_nand3_1 _0495_ (.B(net120),
    .C(_0442_),
    .A(_0006_),
    .Y(_0444_));
 sg13g2_o21ai_1 _0496_ (.B1(_0444_),
    .Y(uo_out[0]),
    .A1(_0439_),
    .A2(net120));
 sg13g2_nor2_1 _0497_ (.A(net120),
    .B(net113),
    .Y(_0445_));
 sg13g2_and3_1 _0498_ (.X(_0446_),
    .A(net3),
    .B(net6),
    .C(_0442_));
 sg13g2_a22oi_1 _0499_ (.Y(_0447_),
    .B1(net6),
    .B2(net2),
    .A2(net3),
    .A1(net5));
 sg13g2_nor2_1 _0500_ (.A(_0446_),
    .B(_0447_),
    .Y(_0448_));
 sg13g2_or2_2 _0501_ (.X(_0449_),
    .B(_0447_),
    .A(_0446_));
 sg13g2_nand2_1 _0502_ (.Y(_0450_),
    .A(_0006_),
    .B(net108));
 sg13g2_nand2_1 _0503_ (.Y(_0451_),
    .A(net115),
    .B(net51));
 sg13g2_xor2_1 _0504_ (.B(net113),
    .A(net114),
    .X(_0452_));
 sg13g2_xnor2_1 _0505_ (.Y(_0453_),
    .A(net114),
    .B(net113));
 sg13g2_nor2_2 _0506_ (.A(_0443_),
    .B(_0453_),
    .Y(_0454_));
 sg13g2_nand3_1 _0507_ (.B(net108),
    .C(_0454_),
    .A(_0006_),
    .Y(_0455_));
 sg13g2_xor2_1 _0508_ (.B(_0454_),
    .A(_0450_),
    .X(_0456_));
 sg13g2_a21oi_2 _0509_ (.B1(_0445_),
    .Y(uo_out[1]),
    .A2(_0456_),
    .A1(net120));
 sg13g2_nand2_1 _0510_ (.Y(_0457_),
    .A(net2),
    .B(net7));
 sg13g2_and4_1 _0511_ (.A(net5),
    .B(net3),
    .C(net6),
    .D(net4),
    .X(_0458_));
 sg13g2_nand4_1 _0512_ (.B(net3),
    .C(net6),
    .A(net5),
    .Y(_0459_),
    .D(net4));
 sg13g2_a22oi_1 _0513_ (.Y(_0460_),
    .B1(net4),
    .B2(net5),
    .A2(net6),
    .A1(net3));
 sg13g2_o21ai_1 _0514_ (.B1(_0457_),
    .Y(_0461_),
    .A1(_0458_),
    .A2(_0460_));
 sg13g2_or3_1 _0515_ (.A(_0457_),
    .B(_0458_),
    .C(_0460_),
    .X(_0462_));
 sg13g2_nand3_1 _0516_ (.B(_0461_),
    .C(_0462_),
    .A(_0446_),
    .Y(_0463_));
 sg13g2_a21o_2 _0517_ (.A2(_0462_),
    .A1(_0461_),
    .B1(_0446_),
    .X(_0464_));
 sg13g2_and2_1 _0518_ (.A(net107),
    .B(_0464_),
    .X(_0465_));
 sg13g2_nand2_2 _0519_ (.Y(_0466_),
    .A(net107),
    .B(_0464_));
 sg13g2_nand3_1 _0520_ (.B(net107),
    .C(_0464_),
    .A(_0452_),
    .Y(_0024_));
 sg13g2_nor2_1 _0521_ (.A(_0450_),
    .B(_0024_),
    .Y(_0025_));
 sg13g2_a22oi_1 _0522_ (.Y(_0026_),
    .B1(_0465_),
    .B2(_0006_),
    .A2(_0452_),
    .A1(net109));
 sg13g2_or2_1 _0523_ (.X(_0027_),
    .B(_0026_),
    .A(_0025_));
 sg13g2_nand3_1 _0524_ (.B(net113),
    .C(\counter_r[2] ),
    .A(net115),
    .Y(_0028_));
 sg13g2_xnor2_1 _0525_ (.Y(_0029_),
    .A(\counter_r[2] ),
    .B(_0451_));
 sg13g2_xnor2_1 _0526_ (.Y(_0030_),
    .A(_0440_),
    .B(_0451_));
 sg13g2_nor2_1 _0527_ (.A(_0443_),
    .B(_0030_),
    .Y(_0031_));
 sg13g2_inv_1 _0528_ (.Y(_0032_),
    .A(_0031_));
 sg13g2_xnor2_1 _0529_ (.Y(_0033_),
    .A(_0027_),
    .B(_0031_));
 sg13g2_nand2b_1 _0530_ (.Y(_0034_),
    .B(_0033_),
    .A_N(_0455_));
 sg13g2_xnor2_1 _0531_ (.Y(_0035_),
    .A(_0455_),
    .B(_0033_));
 sg13g2_nand2_1 _0532_ (.Y(_0036_),
    .A(net120),
    .B(_0035_));
 sg13g2_o21ai_1 _0533_ (.B1(_0036_),
    .Y(uo_out[2]),
    .A1(net119),
    .A2(_0440_));
 sg13g2_nor2_1 _0534_ (.A(net119),
    .B(\counter_r[3] ),
    .Y(_0037_));
 sg13g2_and4_1 _0535_ (.A(net114),
    .B(net113),
    .C(\counter_r[2] ),
    .D(\counter_r[3] ),
    .X(_0038_));
 sg13g2_nand4_1 _0536_ (.B(net113),
    .C(\counter_r[2] ),
    .A(net114),
    .Y(_0039_),
    .D(\counter_r[3] ));
 sg13g2_xnor2_1 _0537_ (.Y(_0040_),
    .A(\counter_r[3] ),
    .B(_0028_));
 sg13g2_xor2_1 _0538_ (.B(_0028_),
    .A(\counter_r[3] ),
    .X(_0041_));
 sg13g2_nor2_1 _0539_ (.A(_0449_),
    .B(_0030_),
    .Y(_0042_));
 sg13g2_o21ai_1 _0540_ (.B1(_0459_),
    .Y(_0043_),
    .A1(_0457_),
    .A2(_0460_));
 sg13g2_nand2_1 _0541_ (.Y(_0044_),
    .A(net4),
    .B(net7));
 sg13g2_and4_1 _0542_ (.A(net3),
    .B(net6),
    .C(net4),
    .D(net7),
    .X(_0045_));
 sg13g2_a22oi_1 _0543_ (.Y(_0046_),
    .B1(net7),
    .B2(net3),
    .A2(net4),
    .A1(net6));
 sg13g2_nor2_1 _0544_ (.A(_0045_),
    .B(_0046_),
    .Y(_0047_));
 sg13g2_nand2_1 _0545_ (.Y(_0048_),
    .A(_0043_),
    .B(_0047_));
 sg13g2_xnor2_1 _0546_ (.Y(_0049_),
    .A(_0043_),
    .B(_0047_));
 sg13g2_xor2_1 _0547_ (.B(_0049_),
    .A(_0463_),
    .X(_0050_));
 sg13g2_xnor2_1 _0548_ (.Y(_0051_),
    .A(_0463_),
    .B(_0049_));
 sg13g2_nor3_1 _0549_ (.A(net115),
    .B(_0024_),
    .C(net101),
    .Y(_0052_));
 sg13g2_o21ai_1 _0550_ (.B1(_0024_),
    .Y(_0053_),
    .A1(net114),
    .A2(net102));
 sg13g2_nor2b_1 _0551_ (.A(_0052_),
    .B_N(_0053_),
    .Y(_0054_));
 sg13g2_xnor2_1 _0552_ (.Y(_0055_),
    .A(_0042_),
    .B(_0054_));
 sg13g2_or3_1 _0553_ (.A(_0450_),
    .B(_0024_),
    .C(_0055_),
    .X(_0056_));
 sg13g2_xor2_1 _0554_ (.B(_0055_),
    .A(_0025_),
    .X(_0057_));
 sg13g2_o21ai_1 _0555_ (.B1(_0057_),
    .Y(_0058_),
    .A1(net116),
    .A2(_0041_));
 sg13g2_or3_1 _0556_ (.A(net116),
    .B(_0041_),
    .C(_0057_),
    .X(_0059_));
 sg13g2_and2_1 _0557_ (.A(_0058_),
    .B(_0059_),
    .X(_0060_));
 sg13g2_o21ai_1 _0558_ (.B1(_0034_),
    .Y(_0061_),
    .A1(_0027_),
    .A2(_0032_));
 sg13g2_xnor2_1 _0559_ (.Y(_0062_),
    .A(_0060_),
    .B(_0061_));
 sg13g2_a21oi_2 _0560_ (.B1(_0037_),
    .Y(uo_out[3]),
    .A2(_0062_),
    .A1(net119));
 sg13g2_nor2_1 _0561_ (.A(_0004_),
    .B(_0039_),
    .Y(_0063_));
 sg13g2_xnor2_1 _0562_ (.Y(_0064_),
    .A(_0004_),
    .B(_0038_));
 sg13g2_xnor2_1 _0563_ (.Y(_0065_),
    .A(_0004_),
    .B(_0039_));
 sg13g2_a21oi_2 _0564_ (.B1(_0044_),
    .Y(_0066_),
    .A2(net6),
    .A1(net3));
 sg13g2_o21ai_1 _0565_ (.B1(_0048_),
    .Y(_0067_),
    .A1(_0463_),
    .A2(_0049_));
 sg13g2_xor2_1 _0566_ (.B(_0067_),
    .A(_0066_),
    .X(_0068_));
 sg13g2_xnor2_1 _0567_ (.Y(_0069_),
    .A(_0066_),
    .B(_0067_));
 sg13g2_nor4_2 _0568_ (.A(net114),
    .B(net116),
    .C(_0065_),
    .Y(_0070_),
    .D(_0069_));
 sg13g2_a22oi_1 _0569_ (.Y(_0071_),
    .B1(net97),
    .B2(_0439_),
    .A2(net106),
    .A1(_0442_));
 sg13g2_nor2_1 _0570_ (.A(_0070_),
    .B(_0071_),
    .Y(_0072_));
 sg13g2_a21oi_1 _0571_ (.A1(_0042_),
    .A2(_0053_),
    .Y(_0073_),
    .B1(_0052_));
 sg13g2_nor2_1 _0572_ (.A(_0449_),
    .B(_0041_),
    .Y(_0074_));
 sg13g2_nand3_1 _0573_ (.B(_0464_),
    .C(_0029_),
    .A(net107),
    .Y(_0075_));
 sg13g2_nor3_1 _0574_ (.A(_0453_),
    .B(net101),
    .C(_0075_),
    .Y(_0076_));
 sg13g2_nand4_1 _0575_ (.B(net104),
    .C(_0029_),
    .A(_0452_),
    .Y(_0077_),
    .D(_0050_));
 sg13g2_o21ai_1 _0576_ (.B1(_0075_),
    .Y(_0078_),
    .A1(_0453_),
    .A2(net101));
 sg13g2_and3_1 _0577_ (.X(_0079_),
    .A(_0074_),
    .B(_0077_),
    .C(_0078_));
 sg13g2_a21oi_1 _0578_ (.A1(_0077_),
    .A2(_0078_),
    .Y(_0080_),
    .B1(_0074_));
 sg13g2_nor3_1 _0579_ (.A(_0073_),
    .B(_0079_),
    .C(_0080_),
    .Y(_0081_));
 sg13g2_o21ai_1 _0580_ (.B1(_0073_),
    .Y(_0082_),
    .A1(_0079_),
    .A2(_0080_));
 sg13g2_nor2b_1 _0581_ (.A(_0081_),
    .B_N(_0082_),
    .Y(_0083_));
 sg13g2_xnor2_1 _0582_ (.Y(_0084_),
    .A(_0072_),
    .B(_0083_));
 sg13g2_a21o_1 _0583_ (.A2(_0059_),
    .A1(_0056_),
    .B1(_0084_),
    .X(_0085_));
 sg13g2_nand3_1 _0584_ (.B(_0059_),
    .C(_0084_),
    .A(_0056_),
    .Y(_0086_));
 sg13g2_and4_1 _0585_ (.A(_0060_),
    .B(_0061_),
    .C(_0085_),
    .D(_0086_),
    .X(_0087_));
 sg13g2_a22oi_1 _0586_ (.Y(_0088_),
    .B1(_0085_),
    .B2(_0086_),
    .A2(_0061_),
    .A1(_0060_));
 sg13g2_nor2_1 _0587_ (.A(_0087_),
    .B(_0088_),
    .Y(_0089_));
 sg13g2_mux2_1 _0588_ (.A0(\counter_r[4] ),
    .A1(_0089_),
    .S(net119),
    .X(uo_out[4]));
 sg13g2_a21oi_1 _0589_ (.A1(_0072_),
    .A2(_0082_),
    .Y(_0090_),
    .B1(_0081_));
 sg13g2_a21oi_2 _0590_ (.B1(_0045_),
    .Y(_0091_),
    .A2(_0067_),
    .A1(_0066_));
 sg13g2_nor2_1 _0591_ (.A(net114),
    .B(net96),
    .Y(_0092_));
 sg13g2_xor2_1 _0592_ (.B(_0063_),
    .A(\counter_r[5] ),
    .X(_0093_));
 sg13g2_xnor2_1 _0593_ (.Y(_0094_),
    .A(net54),
    .B(_0063_));
 sg13g2_nand2_1 _0594_ (.Y(_0095_),
    .A(_0442_),
    .B(net99));
 sg13g2_nand3_1 _0595_ (.B(net97),
    .C(net100),
    .A(_0454_),
    .Y(_0096_));
 sg13g2_o21ai_1 _0596_ (.B1(_0095_),
    .Y(_0097_),
    .A1(_0453_),
    .A2(_0069_));
 sg13g2_nand3_1 _0597_ (.B(_0096_),
    .C(_0097_),
    .A(_0092_),
    .Y(_0098_));
 sg13g2_a21o_1 _0598_ (.A2(_0097_),
    .A1(_0096_),
    .B1(_0092_),
    .X(_0099_));
 sg13g2_a21oi_1 _0599_ (.A1(_0074_),
    .A2(_0078_),
    .Y(_0100_),
    .B1(_0076_));
 sg13g2_nand2_1 _0600_ (.Y(_0101_),
    .A(net108),
    .B(net105));
 sg13g2_nand3_1 _0601_ (.B(_0464_),
    .C(_0040_),
    .A(net107),
    .Y(_0102_));
 sg13g2_nand4_1 _0602_ (.B(_0029_),
    .C(_0040_),
    .A(net104),
    .Y(_0103_),
    .D(_0050_));
 sg13g2_a22oi_1 _0603_ (.Y(_0104_),
    .B1(_0050_),
    .B2(_0029_),
    .A2(_0040_),
    .A1(net104));
 sg13g2_o21ai_1 _0604_ (.B1(_0102_),
    .Y(_0105_),
    .A1(_0030_),
    .A2(net101));
 sg13g2_and4_1 _0605_ (.A(net108),
    .B(net105),
    .C(_0103_),
    .D(_0105_),
    .X(_0106_));
 sg13g2_a22oi_1 _0606_ (.Y(_0107_),
    .B1(_0103_),
    .B2(_0105_),
    .A2(net105),
    .A1(net108));
 sg13g2_nor3_1 _0607_ (.A(_0100_),
    .B(_0106_),
    .C(_0107_),
    .Y(_0108_));
 sg13g2_or3_1 _0608_ (.A(_0100_),
    .B(_0106_),
    .C(_0107_),
    .X(_0109_));
 sg13g2_o21ai_1 _0609_ (.B1(_0100_),
    .Y(_0110_),
    .A1(_0106_),
    .A2(_0107_));
 sg13g2_and4_1 _0610_ (.A(_0098_),
    .B(_0099_),
    .C(_0109_),
    .D(_0110_),
    .X(_0111_));
 sg13g2_a22oi_1 _0611_ (.Y(_0112_),
    .B1(_0109_),
    .B2(_0110_),
    .A2(_0099_),
    .A1(_0098_));
 sg13g2_nor3_1 _0612_ (.A(_0090_),
    .B(_0111_),
    .C(_0112_),
    .Y(_0113_));
 sg13g2_or3_1 _0613_ (.A(_0090_),
    .B(_0111_),
    .C(_0112_),
    .X(_0114_));
 sg13g2_o21ai_1 _0614_ (.B1(_0090_),
    .Y(_0115_),
    .A1(_0111_),
    .A2(_0112_));
 sg13g2_and3_1 _0615_ (.X(_0116_),
    .A(_0070_),
    .B(_0114_),
    .C(_0115_));
 sg13g2_a21oi_1 _0616_ (.A1(_0114_),
    .A2(_0115_),
    .Y(_0117_),
    .B1(_0070_));
 sg13g2_nor3_1 _0617_ (.A(_0085_),
    .B(_0116_),
    .C(_0117_),
    .Y(_0118_));
 sg13g2_o21ai_1 _0618_ (.B1(_0085_),
    .Y(_0119_),
    .A1(_0116_),
    .A2(_0117_));
 sg13g2_nor2b_1 _0619_ (.A(_0118_),
    .B_N(_0119_),
    .Y(_0120_));
 sg13g2_xnor2_1 _0620_ (.Y(_0121_),
    .A(_0087_),
    .B(_0120_));
 sg13g2_nor2_1 _0621_ (.A(net119),
    .B(\counter_r[5] ),
    .Y(_0122_));
 sg13g2_a21oi_2 _0622_ (.B1(_0122_),
    .Y(uo_out[5]),
    .A2(_0121_),
    .A1(net119));
 sg13g2_nor2_1 _0623_ (.A(_0113_),
    .B(_0116_),
    .Y(_0123_));
 sg13g2_and2_1 _0624_ (.A(_0096_),
    .B(_0098_),
    .X(_0124_));
 sg13g2_nor2_1 _0625_ (.A(_0108_),
    .B(_0111_),
    .Y(_0125_));
 sg13g2_nor2_1 _0626_ (.A(_0453_),
    .B(net96),
    .Y(_0126_));
 sg13g2_nand2b_1 _0627_ (.Y(_0127_),
    .B(_0452_),
    .A_N(net96));
 sg13g2_and2_1 _0628_ (.A(\counter_r[4] ),
    .B(\counter_r[5] ),
    .X(_0128_));
 sg13g2_and2_2 _0629_ (.A(_0038_),
    .B(_0128_),
    .X(_0129_));
 sg13g2_and2_2 _0630_ (.A(\counter_r[6] ),
    .B(_0129_),
    .X(_0130_));
 sg13g2_xor2_1 _0631_ (.B(_0129_),
    .A(\counter_r[6] ),
    .X(_0131_));
 sg13g2_xnor2_1 _0632_ (.Y(_0132_),
    .A(\counter_r[6] ),
    .B(_0129_));
 sg13g2_nand2_1 _0633_ (.Y(_0133_),
    .A(net97),
    .B(_0131_));
 sg13g2_nor2_1 _0634_ (.A(net116),
    .B(_0132_),
    .Y(_0134_));
 sg13g2_nand3_1 _0635_ (.B(net98),
    .C(_0134_),
    .A(_0029_),
    .Y(_0135_));
 sg13g2_a21o_1 _0636_ (.A2(net98),
    .A1(_0029_),
    .B1(_0134_),
    .X(_0136_));
 sg13g2_nand3_1 _0637_ (.B(_0135_),
    .C(_0136_),
    .A(_0126_),
    .Y(_0137_));
 sg13g2_a21o_1 _0638_ (.A2(_0136_),
    .A1(_0135_),
    .B1(_0126_),
    .X(_0138_));
 sg13g2_a21o_1 _0639_ (.A2(_0136_),
    .A1(_0135_),
    .B1(_0127_),
    .X(_0139_));
 sg13g2_nand3_1 _0640_ (.B(_0135_),
    .C(_0136_),
    .A(_0127_),
    .Y(_0140_));
 sg13g2_o21ai_1 _0641_ (.B1(_0103_),
    .Y(_0141_),
    .A1(_0101_),
    .A2(_0104_));
 sg13g2_nor2_1 _0642_ (.A(_0449_),
    .B(_0094_),
    .Y(_0142_));
 sg13g2_nand2_1 _0643_ (.Y(_0143_),
    .A(net108),
    .B(net99));
 sg13g2_nand3_1 _0644_ (.B(_0464_),
    .C(net105),
    .A(net107),
    .Y(_0144_));
 sg13g2_nor3_1 _0645_ (.A(net101),
    .B(_0065_),
    .C(_0102_),
    .Y(_0145_));
 sg13g2_nand4_1 _0646_ (.B(_0040_),
    .C(net103),
    .A(net104),
    .Y(_0146_),
    .D(net105));
 sg13g2_a22oi_1 _0647_ (.Y(_0147_),
    .B1(net105),
    .B2(net104),
    .A2(net103),
    .A1(_0040_));
 sg13g2_o21ai_1 _0648_ (.B1(_0144_),
    .Y(_0148_),
    .A1(_0041_),
    .A2(net101));
 sg13g2_nand3_1 _0649_ (.B(_0146_),
    .C(_0148_),
    .A(_0142_),
    .Y(_0149_));
 sg13g2_o21ai_1 _0650_ (.B1(_0143_),
    .Y(_0150_),
    .A1(_0145_),
    .A2(_0147_));
 sg13g2_nand3_1 _0651_ (.B(_0149_),
    .C(_0150_),
    .A(_0141_),
    .Y(_0151_));
 sg13g2_a21o_1 _0652_ (.A2(_0150_),
    .A1(_0149_),
    .B1(_0141_),
    .X(_0152_));
 sg13g2_nand4_1 _0653_ (.B(_0138_),
    .C(_0151_),
    .A(_0137_),
    .Y(_0153_),
    .D(_0152_));
 sg13g2_a22oi_1 _0654_ (.Y(_0154_),
    .B1(_0151_),
    .B2(_0152_),
    .A2(_0140_),
    .A1(_0139_));
 sg13g2_nand4_1 _0655_ (.B(_0140_),
    .C(_0151_),
    .A(_0139_),
    .Y(_0155_),
    .D(_0152_));
 sg13g2_nand2b_2 _0656_ (.Y(_0156_),
    .B(_0155_),
    .A_N(_0154_));
 sg13g2_nand2b_1 _0657_ (.Y(_0157_),
    .B(_0156_),
    .A_N(_0125_));
 sg13g2_xnor2_1 _0658_ (.Y(_0158_),
    .A(_0125_),
    .B(_0156_));
 sg13g2_nand2b_1 _0659_ (.Y(_0159_),
    .B(_0158_),
    .A_N(_0124_));
 sg13g2_xnor2_1 _0660_ (.Y(_0160_),
    .A(_0124_),
    .B(_0158_));
 sg13g2_nor2b_1 _0661_ (.A(_0123_),
    .B_N(_0160_),
    .Y(_0161_));
 sg13g2_xnor2_1 _0662_ (.Y(_0162_),
    .A(_0123_),
    .B(_0160_));
 sg13g2_a21o_1 _0663_ (.A2(_0119_),
    .A1(_0087_),
    .B1(_0118_),
    .X(_0163_));
 sg13g2_xor2_1 _0664_ (.B(_0163_),
    .A(_0162_),
    .X(_0164_));
 sg13g2_mux2_1 _0665_ (.A0(\counter_r[6] ),
    .A1(_0164_),
    .S(net119),
    .X(uo_out[6]));
 sg13g2_a21oi_1 _0666_ (.A1(_0162_),
    .A2(_0163_),
    .Y(_0165_),
    .B1(_0161_));
 sg13g2_nand2_1 _0667_ (.Y(_0166_),
    .A(_0157_),
    .B(_0159_));
 sg13g2_nand2_1 _0668_ (.Y(_0167_),
    .A(_0135_),
    .B(_0137_));
 sg13g2_nor2_1 _0669_ (.A(_0030_),
    .B(net96),
    .Y(_0168_));
 sg13g2_nand2b_1 _0670_ (.Y(_0169_),
    .B(_0029_),
    .A_N(net96));
 sg13g2_and2_1 _0671_ (.A(\counter_r[7] ),
    .B(_0130_),
    .X(_0170_));
 sg13g2_nand4_1 _0672_ (.B(\counter_r[7] ),
    .C(_0038_),
    .A(\counter_r[6] ),
    .Y(_0171_),
    .D(_0128_));
 sg13g2_xor2_1 _0673_ (.B(_0130_),
    .A(\counter_r[7] ),
    .X(_0172_));
 sg13g2_xnor2_1 _0674_ (.Y(_0173_),
    .A(\counter_r[7] ),
    .B(_0130_));
 sg13g2_nor2_2 _0675_ (.A(_0069_),
    .B(_0173_),
    .Y(_0174_));
 sg13g2_nor2_1 _0676_ (.A(net116),
    .B(_0173_),
    .Y(_0175_));
 sg13g2_nand3_1 _0677_ (.B(net98),
    .C(_0175_),
    .A(_0040_),
    .Y(_0176_));
 sg13g2_a21o_1 _0678_ (.A2(net98),
    .A1(_0040_),
    .B1(_0175_),
    .X(_0177_));
 sg13g2_nand3_1 _0679_ (.B(_0176_),
    .C(_0177_),
    .A(_0168_),
    .Y(_0178_));
 sg13g2_a21o_1 _0680_ (.A2(_0177_),
    .A1(_0176_),
    .B1(_0168_),
    .X(_0179_));
 sg13g2_a21o_1 _0681_ (.A2(_0177_),
    .A1(_0176_),
    .B1(_0169_),
    .X(_0180_));
 sg13g2_nand3_1 _0682_ (.B(_0176_),
    .C(_0177_),
    .A(_0169_),
    .Y(_0181_));
 sg13g2_a21oi_1 _0683_ (.A1(_0142_),
    .A2(_0148_),
    .Y(_0182_),
    .B1(_0145_));
 sg13g2_o21ai_1 _0684_ (.B1(_0146_),
    .Y(_0183_),
    .A1(_0143_),
    .A2(_0147_));
 sg13g2_nor2_1 _0685_ (.A(_0449_),
    .B(_0132_),
    .Y(_0184_));
 sg13g2_nand2_1 _0686_ (.Y(_0185_),
    .A(net108),
    .B(_0131_));
 sg13g2_nand3_1 _0687_ (.B(_0464_),
    .C(net99),
    .A(net107),
    .Y(_0186_));
 sg13g2_nor3_2 _0688_ (.A(net101),
    .B(_0065_),
    .C(_0186_),
    .Y(_0187_));
 sg13g2_nand4_1 _0689_ (.B(net103),
    .C(net105),
    .A(net104),
    .Y(_0188_),
    .D(net99));
 sg13g2_a22oi_1 _0690_ (.Y(_0189_),
    .B1(net99),
    .B2(net104),
    .A2(net105),
    .A1(net103));
 sg13g2_o21ai_1 _0691_ (.B1(_0186_),
    .Y(_0190_),
    .A1(net101),
    .A2(_0065_));
 sg13g2_nor3_1 _0692_ (.A(_0185_),
    .B(_0187_),
    .C(_0189_),
    .Y(_0191_));
 sg13g2_nand3_1 _0693_ (.B(_0188_),
    .C(_0190_),
    .A(_0184_),
    .Y(_0192_));
 sg13g2_a21oi_1 _0694_ (.A1(_0188_),
    .A2(_0190_),
    .Y(_0193_),
    .B1(_0184_));
 sg13g2_o21ai_1 _0695_ (.B1(_0185_),
    .Y(_0194_),
    .A1(_0187_),
    .A2(_0189_));
 sg13g2_nand3_1 _0696_ (.B(_0192_),
    .C(_0194_),
    .A(_0183_),
    .Y(_0195_));
 sg13g2_o21ai_1 _0697_ (.B1(_0182_),
    .Y(_0196_),
    .A1(_0191_),
    .A2(_0193_));
 sg13g2_nand3_1 _0698_ (.B(_0192_),
    .C(_0194_),
    .A(_0182_),
    .Y(_0197_));
 sg13g2_o21ai_1 _0699_ (.B1(_0183_),
    .Y(_0198_),
    .A1(_0191_),
    .A2(_0193_));
 sg13g2_nand4_1 _0700_ (.B(_0179_),
    .C(_0195_),
    .A(_0178_),
    .Y(_0199_),
    .D(_0196_));
 sg13g2_nand4_1 _0701_ (.B(_0179_),
    .C(_0197_),
    .A(_0178_),
    .Y(_0200_),
    .D(_0198_));
 sg13g2_nand4_1 _0702_ (.B(_0181_),
    .C(_0195_),
    .A(_0180_),
    .Y(_0201_),
    .D(_0196_));
 sg13g2_a22oi_1 _0703_ (.Y(_0202_),
    .B1(_0200_),
    .B2(_0201_),
    .A2(_0153_),
    .A1(_0151_));
 sg13g2_nand4_1 _0704_ (.B(_0153_),
    .C(_0200_),
    .A(_0151_),
    .Y(_0203_),
    .D(_0201_));
 sg13g2_nand2b_1 _0705_ (.Y(_0204_),
    .B(_0203_),
    .A_N(_0202_));
 sg13g2_xnor2_1 _0706_ (.Y(_0205_),
    .A(_0167_),
    .B(_0204_));
 sg13g2_nor2_1 _0707_ (.A(_0166_),
    .B(_0205_),
    .Y(_0206_));
 sg13g2_xnor2_1 _0708_ (.Y(_0207_),
    .A(_0166_),
    .B(_0205_));
 sg13g2_nor2_1 _0709_ (.A(net118),
    .B(\counter_r[7] ),
    .Y(_0208_));
 sg13g2_xnor2_1 _0710_ (.Y(_0209_),
    .A(_0165_),
    .B(_0207_));
 sg13g2_a21oi_1 _0711_ (.A1(net119),
    .A2(_0209_),
    .Y(uo_out[7]),
    .B1(_0208_));
 sg13g2_nor2_1 _0712_ (.A(net118),
    .B(\counter_r[8] ),
    .Y(_0210_));
 sg13g2_and2_1 _0713_ (.A(_0176_),
    .B(_0178_),
    .X(_0211_));
 sg13g2_nor2_1 _0714_ (.A(_0041_),
    .B(net96),
    .Y(_0212_));
 sg13g2_nand2b_1 _0715_ (.Y(_0213_),
    .B(_0040_),
    .A_N(net96));
 sg13g2_nor2_1 _0716_ (.A(_0005_),
    .B(_0171_),
    .Y(_0214_));
 sg13g2_xor2_1 _0717_ (.B(_0171_),
    .A(_0005_),
    .X(_0215_));
 sg13g2_xnor2_1 _0718_ (.Y(_0216_),
    .A(_0005_),
    .B(_0171_));
 sg13g2_nand2_1 _0719_ (.Y(_0217_),
    .A(net97),
    .B(_0215_));
 sg13g2_nor2_1 _0720_ (.A(net116),
    .B(_0216_),
    .Y(_0218_));
 sg13g2_nand2_1 _0721_ (.Y(_0219_),
    .A(_0442_),
    .B(_0215_));
 sg13g2_nor3_2 _0722_ (.A(_0065_),
    .B(_0069_),
    .C(_0219_),
    .Y(_0220_));
 sg13g2_nand3_1 _0723_ (.B(net97),
    .C(_0218_),
    .A(net106),
    .Y(_0221_));
 sg13g2_a21oi_1 _0724_ (.A1(net106),
    .A2(net97),
    .Y(_0222_),
    .B1(_0218_));
 sg13g2_o21ai_1 _0725_ (.B1(_0219_),
    .Y(_0223_),
    .A1(_0065_),
    .A2(_0069_));
 sg13g2_nand3_1 _0726_ (.B(_0221_),
    .C(_0223_),
    .A(_0212_),
    .Y(_0224_));
 sg13g2_o21ai_1 _0727_ (.B1(_0213_),
    .Y(_0225_),
    .A1(_0220_),
    .A2(_0222_));
 sg13g2_o21ai_1 _0728_ (.B1(_0212_),
    .Y(_0226_),
    .A1(_0220_),
    .A2(_0222_));
 sg13g2_nand3_1 _0729_ (.B(_0221_),
    .C(_0223_),
    .A(_0213_),
    .Y(_0227_));
 sg13g2_a21oi_1 _0730_ (.A1(_0184_),
    .A2(_0190_),
    .Y(_0228_),
    .B1(_0187_));
 sg13g2_o21ai_1 _0731_ (.B1(_0188_),
    .Y(_0229_),
    .A1(_0185_),
    .A2(_0189_));
 sg13g2_nor2_1 _0732_ (.A(_0449_),
    .B(_0173_),
    .Y(_0230_));
 sg13g2_nand2_1 _0733_ (.Y(_0231_),
    .A(net108),
    .B(_0172_));
 sg13g2_and3_1 _0734_ (.X(_0232_),
    .A(net107),
    .B(_0464_),
    .C(_0131_));
 sg13g2_nor3_2 _0735_ (.A(_0051_),
    .B(_0132_),
    .C(_0186_),
    .Y(_0233_));
 sg13g2_nand3_1 _0736_ (.B(net99),
    .C(_0232_),
    .A(net103),
    .Y(_0234_));
 sg13g2_a21oi_1 _0737_ (.A1(net103),
    .A2(net99),
    .Y(_0235_),
    .B1(_0232_));
 sg13g2_a21o_1 _0738_ (.A2(net99),
    .A1(net103),
    .B1(_0232_),
    .X(_0236_));
 sg13g2_nor3_1 _0739_ (.A(_0231_),
    .B(_0233_),
    .C(_0235_),
    .Y(_0237_));
 sg13g2_nand3_1 _0740_ (.B(_0234_),
    .C(_0236_),
    .A(_0230_),
    .Y(_0238_));
 sg13g2_a21oi_1 _0741_ (.A1(_0234_),
    .A2(_0236_),
    .Y(_0239_),
    .B1(_0230_));
 sg13g2_o21ai_1 _0742_ (.B1(_0231_),
    .Y(_0240_),
    .A1(_0233_),
    .A2(_0235_));
 sg13g2_nand3_1 _0743_ (.B(_0238_),
    .C(_0240_),
    .A(_0229_),
    .Y(_0241_));
 sg13g2_o21ai_1 _0744_ (.B1(_0228_),
    .Y(_0242_),
    .A1(_0237_),
    .A2(_0239_));
 sg13g2_nand3_1 _0745_ (.B(_0238_),
    .C(_0240_),
    .A(_0228_),
    .Y(_0243_));
 sg13g2_o21ai_1 _0746_ (.B1(_0229_),
    .Y(_0244_),
    .A1(_0237_),
    .A2(_0239_));
 sg13g2_nand4_1 _0747_ (.B(_0225_),
    .C(_0241_),
    .A(_0224_),
    .Y(_0245_),
    .D(_0242_));
 sg13g2_nand4_1 _0748_ (.B(_0225_),
    .C(_0243_),
    .A(_0224_),
    .Y(_0246_),
    .D(_0244_));
 sg13g2_nand4_1 _0749_ (.B(_0227_),
    .C(_0241_),
    .A(_0226_),
    .Y(_0247_),
    .D(_0242_));
 sg13g2_a22oi_1 _0750_ (.Y(_0248_),
    .B1(_0246_),
    .B2(_0247_),
    .A2(_0199_),
    .A1(_0195_));
 sg13g2_and4_1 _0751_ (.A(_0195_),
    .B(_0199_),
    .C(_0246_),
    .D(_0247_),
    .X(_0249_));
 sg13g2_o21ai_1 _0752_ (.B1(_0211_),
    .Y(_0250_),
    .A1(_0248_),
    .A2(_0249_));
 sg13g2_or3_1 _0753_ (.A(_0211_),
    .B(_0248_),
    .C(_0249_),
    .X(_0251_));
 sg13g2_nand2_1 _0754_ (.Y(_0252_),
    .A(_0250_),
    .B(_0251_));
 sg13g2_a21o_1 _0755_ (.A2(_0203_),
    .A1(_0167_),
    .B1(_0202_),
    .X(_0253_));
 sg13g2_nand3_1 _0756_ (.B(_0251_),
    .C(_0253_),
    .A(_0250_),
    .Y(_0254_));
 sg13g2_xnor2_1 _0757_ (.Y(_0255_),
    .A(_0252_),
    .B(_0253_));
 sg13g2_a221oi_1 _0758_ (.B2(_0205_),
    .C1(_0161_),
    .B1(_0166_),
    .A1(_0162_),
    .Y(_0256_),
    .A2(_0163_));
 sg13g2_or2_1 _0759_ (.X(_0257_),
    .B(_0256_),
    .A(_0206_));
 sg13g2_nor2_2 _0760_ (.A(_0206_),
    .B(_0256_),
    .Y(_0258_));
 sg13g2_nand2_1 _0761_ (.Y(_0259_),
    .A(_0255_),
    .B(_0258_));
 sg13g2_xnor2_1 _0762_ (.Y(_0260_),
    .A(_0255_),
    .B(_0258_));
 sg13g2_a21oi_2 _0763_ (.B1(_0210_),
    .Y(uio_out[0]),
    .A2(_0260_),
    .A1(net118));
 sg13g2_nor2b_2 _0764_ (.A(_0248_),
    .B_N(_0251_),
    .Y(_0261_));
 sg13g2_a21oi_1 _0765_ (.A1(_0212_),
    .A2(_0223_),
    .Y(_0262_),
    .B1(_0220_));
 sg13g2_nor2_1 _0766_ (.A(_0065_),
    .B(net95),
    .Y(_0263_));
 sg13g2_nand2b_1 _0767_ (.Y(_0264_),
    .B(net106),
    .A_N(net95));
 sg13g2_xnor2_1 _0768_ (.Y(_0265_),
    .A(\counter_r[9] ),
    .B(_0214_));
 sg13g2_nor2_1 _0769_ (.A(_0069_),
    .B(_0265_),
    .Y(_0266_));
 sg13g2_nor2_1 _0770_ (.A(net116),
    .B(_0265_),
    .Y(_0267_));
 sg13g2_nor3_2 _0771_ (.A(_0069_),
    .B(_0095_),
    .C(_0265_),
    .Y(_0268_));
 sg13g2_a21oi_2 _0772_ (.B1(_0267_),
    .Y(_0269_),
    .A2(net100),
    .A1(net97));
 sg13g2_or3_1 _0773_ (.A(_0264_),
    .B(_0268_),
    .C(_0269_),
    .X(_0270_));
 sg13g2_o21ai_1 _0774_ (.B1(_0264_),
    .Y(_0271_),
    .A1(_0268_),
    .A2(_0269_));
 sg13g2_o21ai_1 _0775_ (.B1(_0263_),
    .Y(_0272_),
    .A1(_0268_),
    .A2(_0269_));
 sg13g2_or3_1 _0776_ (.A(_0263_),
    .B(_0268_),
    .C(_0269_),
    .X(_0273_));
 sg13g2_a21oi_1 _0777_ (.A1(_0230_),
    .A2(_0236_),
    .Y(_0274_),
    .B1(_0233_));
 sg13g2_o21ai_1 _0778_ (.B1(_0234_),
    .Y(_0275_),
    .A1(_0231_),
    .A2(_0235_));
 sg13g2_nand2_1 _0779_ (.Y(_0276_),
    .A(net109),
    .B(_0215_));
 sg13g2_nor2_1 _0780_ (.A(net102),
    .B(_0173_),
    .Y(_0277_));
 sg13g2_nor4_2 _0781_ (.A(_0466_),
    .B(net102),
    .C(_0132_),
    .Y(_0278_),
    .D(_0173_));
 sg13g2_a22oi_1 _0782_ (.Y(_0279_),
    .B1(_0172_),
    .B2(net104),
    .A2(_0131_),
    .A1(net103));
 sg13g2_or3_2 _0783_ (.A(_0276_),
    .B(_0278_),
    .C(_0279_),
    .X(_0280_));
 sg13g2_o21ai_1 _0784_ (.B1(_0276_),
    .Y(_0281_),
    .A1(_0278_),
    .A2(_0279_));
 sg13g2_nand3_1 _0785_ (.B(_0280_),
    .C(_0281_),
    .A(_0275_),
    .Y(_0282_));
 sg13g2_a21o_1 _0786_ (.A2(_0281_),
    .A1(_0280_),
    .B1(_0275_),
    .X(_0283_));
 sg13g2_nand3_1 _0787_ (.B(_0280_),
    .C(_0281_),
    .A(_0274_),
    .Y(_0284_));
 sg13g2_a21o_1 _0788_ (.A2(_0281_),
    .A1(_0280_),
    .B1(_0274_),
    .X(_0285_));
 sg13g2_nand4_1 _0789_ (.B(_0271_),
    .C(_0282_),
    .A(_0270_),
    .Y(_0286_),
    .D(_0283_));
 sg13g2_nand4_1 _0790_ (.B(_0271_),
    .C(_0284_),
    .A(_0270_),
    .Y(_0287_),
    .D(_0285_));
 sg13g2_nand4_1 _0791_ (.B(_0273_),
    .C(_0282_),
    .A(_0272_),
    .Y(_0288_),
    .D(_0283_));
 sg13g2_a22oi_1 _0792_ (.Y(_0289_),
    .B1(_0287_),
    .B2(_0288_),
    .A2(_0245_),
    .A1(_0241_));
 sg13g2_and4_1 _0793_ (.A(_0241_),
    .B(_0245_),
    .C(_0287_),
    .D(_0288_),
    .X(_0290_));
 sg13g2_or3_1 _0794_ (.A(_0262_),
    .B(_0289_),
    .C(_0290_),
    .X(_0291_));
 sg13g2_o21ai_1 _0795_ (.B1(_0262_),
    .Y(_0292_),
    .A1(_0289_),
    .A2(_0290_));
 sg13g2_nand2_1 _0796_ (.Y(_0293_),
    .A(_0291_),
    .B(_0292_));
 sg13g2_nand2_1 _0797_ (.Y(_0294_),
    .A(_0261_),
    .B(_0293_));
 sg13g2_xor2_1 _0798_ (.B(_0293_),
    .A(_0261_),
    .X(_0295_));
 sg13g2_and2_1 _0799_ (.A(_0254_),
    .B(_0259_),
    .X(_0296_));
 sg13g2_xnor2_1 _0800_ (.Y(_0297_),
    .A(_0295_),
    .B(_0296_));
 sg13g2_mux2_1 _0801_ (.A0(\counter_r[9] ),
    .A1(_0297_),
    .S(net117),
    .X(uio_out[1]));
 sg13g2_o21ai_1 _0802_ (.B1(_0254_),
    .Y(_0298_),
    .A1(_0261_),
    .A2(_0293_));
 sg13g2_and3_1 _0803_ (.X(_0299_),
    .A(_0255_),
    .B(_0258_),
    .C(_0295_));
 sg13g2_a21o_1 _0804_ (.A2(_0298_),
    .A1(_0294_),
    .B1(_0299_),
    .X(_0300_));
 sg13g2_nor2b_1 _0805_ (.A(_0289_),
    .B_N(_0291_),
    .Y(_0301_));
 sg13g2_nand2b_1 _0806_ (.Y(_0302_),
    .B(_0270_),
    .A_N(_0268_));
 sg13g2_nand2_1 _0807_ (.Y(_0303_),
    .A(_0282_),
    .B(_0286_));
 sg13g2_and3_1 _0808_ (.X(_0304_),
    .A(\counter_r[8] ),
    .B(\counter_r[9] ),
    .C(_0170_));
 sg13g2_nand3_1 _0809_ (.B(\counter_r[9] ),
    .C(_0170_),
    .A(\counter_r[8] ),
    .Y(_0305_));
 sg13g2_o21ai_1 _0810_ (.B1(_0133_),
    .Y(_0306_),
    .A1(net116),
    .A2(_0305_));
 sg13g2_nand2b_1 _0811_ (.Y(_0307_),
    .B(net100),
    .A_N(net95));
 sg13g2_nor2b_1 _0812_ (.A(_0307_),
    .B_N(_0306_),
    .Y(_0308_));
 sg13g2_xor2_1 _0813_ (.B(_0307_),
    .A(_0306_),
    .X(_0309_));
 sg13g2_nand2b_1 _0814_ (.Y(_0310_),
    .B(_0280_),
    .A_N(_0278_));
 sg13g2_nor2_1 _0815_ (.A(_0449_),
    .B(_0265_),
    .Y(_0311_));
 sg13g2_nor2_1 _0816_ (.A(net102),
    .B(_0216_),
    .Y(_0312_));
 sg13g2_nor2_2 _0817_ (.A(_0466_),
    .B(_0216_),
    .Y(_0313_));
 sg13g2_and2_1 _0818_ (.A(_0277_),
    .B(_0313_),
    .X(_0314_));
 sg13g2_or2_1 _0819_ (.X(_0315_),
    .B(_0313_),
    .A(_0277_));
 sg13g2_xnor2_1 _0820_ (.Y(_0316_),
    .A(_0277_),
    .B(_0313_));
 sg13g2_xnor2_1 _0821_ (.Y(_0317_),
    .A(_0311_),
    .B(_0316_));
 sg13g2_nand2_1 _0822_ (.Y(_0318_),
    .A(_0310_),
    .B(_0317_));
 sg13g2_xnor2_1 _0823_ (.Y(_0319_),
    .A(_0310_),
    .B(_0317_));
 sg13g2_xor2_1 _0824_ (.B(_0319_),
    .A(_0309_),
    .X(_0320_));
 sg13g2_and2_1 _0825_ (.A(_0303_),
    .B(_0320_),
    .X(_0321_));
 sg13g2_or2_1 _0826_ (.X(_0322_),
    .B(_0320_),
    .A(_0303_));
 sg13g2_xnor2_1 _0827_ (.Y(_0323_),
    .A(_0303_),
    .B(_0320_));
 sg13g2_xnor2_1 _0828_ (.Y(_0324_),
    .A(_0302_),
    .B(_0323_));
 sg13g2_nor2b_1 _0829_ (.A(_0301_),
    .B_N(_0324_),
    .Y(_0325_));
 sg13g2_xnor2_1 _0830_ (.Y(_0326_),
    .A(_0301_),
    .B(_0324_));
 sg13g2_xnor2_1 _0831_ (.Y(_0327_),
    .A(_0300_),
    .B(_0326_));
 sg13g2_nor2_1 _0832_ (.A(net118),
    .B(\counter_r[10] ),
    .Y(_0328_));
 sg13g2_a21oi_2 _0833_ (.B1(_0328_),
    .Y(uio_out[2]),
    .A2(_0327_),
    .A1(net118));
 sg13g2_nor2_1 _0834_ (.A(net117),
    .B(\counter_r[11] ),
    .Y(_0329_));
 sg13g2_a21oi_1 _0835_ (.A1(_0300_),
    .A2(_0326_),
    .Y(_0330_),
    .B1(_0325_));
 sg13g2_a21oi_2 _0836_ (.B1(_0321_),
    .Y(_0331_),
    .A2(_0322_),
    .A1(_0302_));
 sg13g2_o21ai_1 _0837_ (.B1(_0318_),
    .Y(_0332_),
    .A1(_0309_),
    .A2(_0319_));
 sg13g2_nor2_1 _0838_ (.A(net95),
    .B(_0132_),
    .Y(_0333_));
 sg13g2_and2_1 _0839_ (.A(_0174_),
    .B(_0333_),
    .X(_0334_));
 sg13g2_xor2_1 _0840_ (.B(_0333_),
    .A(_0174_),
    .X(_0335_));
 sg13g2_a21oi_1 _0841_ (.A1(_0311_),
    .A2(_0315_),
    .Y(_0336_),
    .B1(_0314_));
 sg13g2_nand2_1 _0842_ (.Y(_0337_),
    .A(net109),
    .B(_0304_));
 sg13g2_or2_1 _0843_ (.X(_0338_),
    .B(_0265_),
    .A(net102));
 sg13g2_nor2_1 _0844_ (.A(_0466_),
    .B(_0265_),
    .Y(_0339_));
 sg13g2_nand2_1 _0845_ (.Y(_0340_),
    .A(_0312_),
    .B(_0339_));
 sg13g2_xnor2_1 _0846_ (.Y(_0341_),
    .A(_0312_),
    .B(_0339_));
 sg13g2_or2_1 _0847_ (.X(_0342_),
    .B(_0341_),
    .A(_0337_));
 sg13g2_xnor2_1 _0848_ (.Y(_0343_),
    .A(_0337_),
    .B(_0341_));
 sg13g2_nor2_1 _0849_ (.A(_0336_),
    .B(_0343_),
    .Y(_0344_));
 sg13g2_xor2_1 _0850_ (.B(_0343_),
    .A(_0336_),
    .X(_0345_));
 sg13g2_xor2_1 _0851_ (.B(_0345_),
    .A(_0335_),
    .X(_0346_));
 sg13g2_and2_1 _0852_ (.A(_0332_),
    .B(_0346_),
    .X(_0347_));
 sg13g2_xor2_1 _0853_ (.B(_0346_),
    .A(_0332_),
    .X(_0348_));
 sg13g2_xnor2_1 _0854_ (.Y(_0349_),
    .A(_0308_),
    .B(_0348_));
 sg13g2_nand2_1 _0855_ (.Y(_0350_),
    .A(_0331_),
    .B(_0349_));
 sg13g2_or2_1 _0856_ (.X(_0351_),
    .B(_0349_),
    .A(_0331_));
 sg13g2_xor2_1 _0857_ (.B(_0349_),
    .A(_0331_),
    .X(_0352_));
 sg13g2_xor2_1 _0858_ (.B(_0352_),
    .A(_0330_),
    .X(_0353_));
 sg13g2_a21oi_2 _0859_ (.B1(_0329_),
    .Y(uio_out[3]),
    .A2(_0353_),
    .A1(net118));
 sg13g2_nor2_1 _0860_ (.A(net117),
    .B(\counter_r[12] ),
    .Y(_0354_));
 sg13g2_a21o_1 _0861_ (.A2(_0348_),
    .A1(_0308_),
    .B1(_0347_),
    .X(_0355_));
 sg13g2_a21oi_1 _0862_ (.A1(_0335_),
    .A2(_0345_),
    .Y(_0356_),
    .B1(_0344_));
 sg13g2_o21ai_1 _0863_ (.B1(_0338_),
    .Y(_0357_),
    .A1(_0466_),
    .A2(_0305_));
 sg13g2_nor3_1 _0864_ (.A(_0466_),
    .B(_0305_),
    .C(_0338_),
    .Y(_0358_));
 sg13g2_a21oi_1 _0865_ (.A1(_0340_),
    .A2(_0342_),
    .Y(_0359_),
    .B1(_0358_));
 sg13g2_a21o_1 _0866_ (.A2(_0342_),
    .A1(_0340_),
    .B1(_0358_),
    .X(_0360_));
 sg13g2_nand2_1 _0867_ (.Y(_0361_),
    .A(_0357_),
    .B(_0360_));
 sg13g2_o21ai_1 _0868_ (.B1(_0217_),
    .Y(_0362_),
    .A1(net95),
    .A2(_0173_));
 sg13g2_nor2_1 _0869_ (.A(net95),
    .B(_0216_),
    .Y(_0363_));
 sg13g2_nand2_1 _0870_ (.Y(_0364_),
    .A(_0174_),
    .B(_0363_));
 sg13g2_and2_1 _0871_ (.A(_0362_),
    .B(_0364_),
    .X(_0365_));
 sg13g2_xnor2_1 _0872_ (.Y(_0366_),
    .A(_0361_),
    .B(_0365_));
 sg13g2_nand2b_1 _0873_ (.Y(_0367_),
    .B(_0366_),
    .A_N(_0356_));
 sg13g2_xnor2_1 _0874_ (.Y(_0368_),
    .A(_0356_),
    .B(_0366_));
 sg13g2_nand2_1 _0875_ (.Y(_0369_),
    .A(_0334_),
    .B(_0368_));
 sg13g2_xnor2_1 _0876_ (.Y(_0370_),
    .A(_0334_),
    .B(_0368_));
 sg13g2_nor2b_1 _0877_ (.A(_0370_),
    .B_N(_0355_),
    .Y(_0371_));
 sg13g2_xnor2_1 _0878_ (.Y(_0372_),
    .A(_0355_),
    .B(_0370_));
 sg13g2_nand4_1 _0879_ (.B(_0295_),
    .C(_0326_),
    .A(_0255_),
    .Y(_0373_),
    .D(_0352_));
 sg13g2_nand4_1 _0880_ (.B(_0298_),
    .C(_0326_),
    .A(_0294_),
    .Y(_0374_),
    .D(_0352_));
 sg13g2_nand2_1 _0881_ (.Y(_0375_),
    .A(_0325_),
    .B(_0350_));
 sg13g2_and3_1 _0882_ (.X(_0376_),
    .A(_0351_),
    .B(_0374_),
    .C(_0375_));
 sg13g2_o21ai_1 _0883_ (.B1(_0376_),
    .Y(_0377_),
    .A1(_0257_),
    .A2(_0373_));
 sg13g2_xnor2_1 _0884_ (.Y(_0378_),
    .A(_0372_),
    .B(_0377_));
 sg13g2_a21oi_2 _0885_ (.B1(_0354_),
    .Y(uio_out[4]),
    .A2(_0378_),
    .A1(net117));
 sg13g2_nand2_1 _0886_ (.Y(_0379_),
    .A(_0367_),
    .B(_0369_));
 sg13g2_nor3_1 _0887_ (.A(net102),
    .B(_0305_),
    .C(_0313_),
    .Y(_0380_));
 sg13g2_nor2_1 _0888_ (.A(net95),
    .B(_0265_),
    .Y(_0381_));
 sg13g2_nand2_1 _0889_ (.Y(_0382_),
    .A(_0266_),
    .B(_0363_));
 sg13g2_xnor2_1 _0890_ (.Y(_0383_),
    .A(_0266_),
    .B(_0363_));
 sg13g2_nor4_1 _0891_ (.A(net102),
    .B(_0305_),
    .C(_0313_),
    .D(_0383_),
    .Y(_0384_));
 sg13g2_xnor2_1 _0892_ (.Y(_0385_),
    .A(_0380_),
    .B(_0383_));
 sg13g2_a21oi_1 _0893_ (.A1(_0357_),
    .A2(_0365_),
    .Y(_0386_),
    .B1(_0359_));
 sg13g2_inv_1 _0894_ (.Y(_0387_),
    .A(_0386_));
 sg13g2_nand2_1 _0895_ (.Y(_0388_),
    .A(_0385_),
    .B(_0387_));
 sg13g2_xor2_1 _0896_ (.B(_0386_),
    .A(_0385_),
    .X(_0389_));
 sg13g2_xnor2_1 _0897_ (.Y(_0390_),
    .A(_0364_),
    .B(_0389_));
 sg13g2_nand3_1 _0898_ (.B(_0369_),
    .C(_0390_),
    .A(_0367_),
    .Y(_0391_));
 sg13g2_a21oi_1 _0899_ (.A1(_0367_),
    .A2(_0369_),
    .Y(_0392_),
    .B1(_0390_));
 sg13g2_xnor2_1 _0900_ (.Y(_0393_),
    .A(_0379_),
    .B(_0390_));
 sg13g2_a21oi_1 _0901_ (.A1(_0372_),
    .A2(_0377_),
    .Y(_0394_),
    .B1(_0371_));
 sg13g2_xnor2_1 _0902_ (.Y(_0395_),
    .A(_0393_),
    .B(_0394_));
 sg13g2_mux2_1 _0903_ (.A0(\counter_r[13] ),
    .A1(_0395_),
    .S(net117),
    .X(uio_out[5]));
 sg13g2_and2_1 _0904_ (.A(_0372_),
    .B(_0393_),
    .X(_0396_));
 sg13g2_a221oi_1 _0905_ (.B2(_0377_),
    .C1(_0392_),
    .B1(_0396_),
    .A1(_0371_),
    .Y(_0397_),
    .A2(_0391_));
 sg13g2_nor2_1 _0906_ (.A(_0358_),
    .B(_0384_),
    .Y(_0398_));
 sg13g2_nand2_1 _0907_ (.Y(_0399_),
    .A(net97),
    .B(_0304_));
 sg13g2_xnor2_1 _0908_ (.Y(_0400_),
    .A(_0381_),
    .B(_0399_));
 sg13g2_inv_1 _0909_ (.Y(_0401_),
    .A(_0400_));
 sg13g2_xnor2_1 _0910_ (.Y(_0402_),
    .A(_0398_),
    .B(_0400_));
 sg13g2_nand2b_1 _0911_ (.Y(_0403_),
    .B(_0402_),
    .A_N(_0382_));
 sg13g2_xnor2_1 _0912_ (.Y(_0404_),
    .A(_0382_),
    .B(_0402_));
 sg13g2_o21ai_1 _0913_ (.B1(_0388_),
    .Y(_0405_),
    .A1(_0364_),
    .A2(_0389_));
 sg13g2_nand2_1 _0914_ (.Y(_0406_),
    .A(_0404_),
    .B(_0405_));
 sg13g2_nor2_1 _0915_ (.A(_0404_),
    .B(_0405_),
    .Y(_0407_));
 sg13g2_xor2_1 _0916_ (.B(_0405_),
    .A(_0404_),
    .X(_0408_));
 sg13g2_xnor2_1 _0917_ (.Y(_0409_),
    .A(_0397_),
    .B(_0408_));
 sg13g2_mux2_1 _0918_ (.A0(\counter_r[14] ),
    .A1(_0409_),
    .S(net117),
    .X(uio_out[6]));
 sg13g2_o21ai_1 _0919_ (.B1(_0406_),
    .Y(_0410_),
    .A1(_0397_),
    .A2(_0407_));
 sg13g2_o21ai_1 _0920_ (.B1(_0403_),
    .Y(_0411_),
    .A1(_0398_),
    .A2(_0401_));
 sg13g2_nand3b_1 _0921_ (.B(_0217_),
    .C(_0304_),
    .Y(_0412_),
    .A_N(net95));
 sg13g2_xnor2_1 _0922_ (.Y(_0413_),
    .A(_0411_),
    .B(_0412_));
 sg13g2_xnor2_1 _0923_ (.Y(_0414_),
    .A(_0410_),
    .B(_0413_));
 sg13g2_nor2_1 _0924_ (.A(net117),
    .B(\counter_r[15] ),
    .Y(_0415_));
 sg13g2_a21oi_1 _0925_ (.A1(net117),
    .A2(_0414_),
    .Y(uio_out[7]),
    .B1(_0415_));
 sg13g2_xnor2_1 _0926_ (.Y(_0416_),
    .A(net34),
    .B(net112));
 sg13g2_inv_1 _0927_ (.Y(_0417_),
    .A(_0416_));
 sg13g2_nor2_1 _0928_ (.A(net20),
    .B(_0416_),
    .Y(_0000_));
 sg13g2_xnor2_1 _0929_ (.Y(_0418_),
    .A(net43),
    .B(net20));
 sg13g2_nor2_1 _0930_ (.A(_0416_),
    .B(_0418_),
    .Y(_0001_));
 sg13g2_a21oi_1 _0931_ (.A1(\counter_db_r[1] ),
    .A2(net20),
    .Y(_0419_),
    .B1(net22));
 sg13g2_and3_1 _0932_ (.X(_0420_),
    .A(\counter_db_r[1] ),
    .B(net20),
    .C(net22));
 sg13g2_nor3_1 _0933_ (.A(_0416_),
    .B(net23),
    .C(_0420_),
    .Y(_0002_));
 sg13g2_nand2_1 _0934_ (.Y(_0421_),
    .A(net41),
    .B(_0420_));
 sg13g2_o21ai_1 _0935_ (.B1(_0417_),
    .Y(_0422_),
    .A1(net41),
    .A2(_0420_));
 sg13g2_nor2b_1 _0936_ (.A(net42),
    .B_N(_0421_),
    .Y(_0003_));
 sg13g2_nand2_1 _0937_ (.Y(_0423_),
    .A(net45),
    .B(net111));
 sg13g2_o21ai_1 _0938_ (.B1(_0423_),
    .Y(_0007_),
    .A1(_0439_),
    .A2(net111));
 sg13g2_nor2_1 _0939_ (.A(net113),
    .B(net112),
    .Y(_0424_));
 sg13g2_a21oi_1 _0940_ (.A1(net112),
    .A2(_0453_),
    .Y(_0008_),
    .B1(_0424_));
 sg13g2_nand4_1 _0941_ (.B(net113),
    .C(\counter_r[2] ),
    .A(net115),
    .Y(_0425_),
    .D(net112));
 sg13g2_o21ai_1 _0942_ (.B1(_0425_),
    .Y(_0426_),
    .A1(\counter_r[2] ),
    .A2(net112));
 sg13g2_a21oi_1 _0943_ (.A1(_0440_),
    .A2(net52),
    .Y(_0009_),
    .B1(_0426_));
 sg13g2_xnor2_1 _0944_ (.Y(_0010_),
    .A(net57),
    .B(_0425_));
 sg13g2_nor2_1 _0945_ (.A(net33),
    .B(net111),
    .Y(_0427_));
 sg13g2_a21oi_1 _0946_ (.A1(net110),
    .A2(_0065_),
    .Y(_0011_),
    .B1(_0427_));
 sg13g2_nor2_1 _0947_ (.A(net54),
    .B(net111),
    .Y(_0428_));
 sg13g2_a21oi_1 _0948_ (.A1(net111),
    .A2(_0094_),
    .Y(_0012_),
    .B1(_0428_));
 sg13g2_nand2_1 _0949_ (.Y(_0429_),
    .A(net111),
    .B(_0130_));
 sg13g2_a21oi_1 _0950_ (.A1(net110),
    .A2(_0129_),
    .Y(_0430_),
    .B1(net50));
 sg13g2_a21oi_1 _0951_ (.A1(net110),
    .A2(_0130_),
    .Y(_0013_),
    .B1(_0430_));
 sg13g2_xnor2_1 _0952_ (.Y(_0014_),
    .A(net55),
    .B(_0429_));
 sg13g2_nor2_1 _0953_ (.A(net47),
    .B(net110),
    .Y(_0431_));
 sg13g2_a21oi_1 _0954_ (.A1(net110),
    .A2(_0216_),
    .Y(_0015_),
    .B1(_0431_));
 sg13g2_nor2_1 _0955_ (.A(net49),
    .B(net110),
    .Y(_0432_));
 sg13g2_a21oi_1 _0956_ (.A1(net110),
    .A2(_0265_),
    .Y(_0016_),
    .B1(_0432_));
 sg13g2_nand4_1 _0957_ (.B(\counter_r[9] ),
    .C(net110),
    .A(\counter_r[8] ),
    .Y(_0433_),
    .D(_0170_));
 sg13g2_nor2_1 _0958_ (.A(_0441_),
    .B(_0433_),
    .Y(_0434_));
 sg13g2_xnor2_1 _0959_ (.Y(_0017_),
    .A(net36),
    .B(_0433_));
 sg13g2_xor2_1 _0960_ (.B(_0434_),
    .A(net38),
    .X(_0018_));
 sg13g2_a21oi_1 _0961_ (.A1(\counter_r[11] ),
    .A2(_0434_),
    .Y(_0435_),
    .B1(net30));
 sg13g2_and3_1 _0962_ (.X(_0436_),
    .A(net38),
    .B(net30),
    .C(_0434_));
 sg13g2_nor2_1 _0963_ (.A(net31),
    .B(_0436_),
    .Y(_0019_));
 sg13g2_xor2_1 _0964_ (.B(_0436_),
    .A(net40),
    .X(_0020_));
 sg13g2_a21oi_1 _0965_ (.A1(\counter_r[13] ),
    .A2(_0436_),
    .Y(_0437_),
    .B1(net27));
 sg13g2_nand3_1 _0966_ (.B(net27),
    .C(_0436_),
    .A(\counter_r[13] ),
    .Y(_0438_));
 sg13g2_nor2b_1 _0967_ (.A(net28),
    .B_N(_0438_),
    .Y(_0021_));
 sg13g2_xnor2_1 _0968_ (.Y(_0022_),
    .A(net25),
    .B(_0438_));
 sg13g2_mux2_1 _0969_ (.A0(net34),
    .A1(net112),
    .S(_0421_),
    .X(_0023_));
 sg13g2_dfrbp_1 _0970_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net126),
    .D(net46),
    .Q_N(_0006_),
    .Q(\counter_r[0] ));
 sg13g2_dfrbp_1 _0971_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net125),
    .D(_0008_),
    .Q_N(_0480_),
    .Q(\counter_r[1] ));
 sg13g2_dfrbp_1 _0972_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net126),
    .D(net53),
    .Q_N(_0479_),
    .Q(\counter_r[2] ));
 sg13g2_dfrbp_1 _0973_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net126),
    .D(net58),
    .Q_N(_0478_),
    .Q(\counter_r[3] ));
 sg13g2_dfrbp_1 _0974_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net123),
    .D(_0011_),
    .Q_N(_0004_),
    .Q(\counter_r[4] ));
 sg13g2_dfrbp_1 _0975_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net123),
    .D(_0012_),
    .Q_N(_0477_),
    .Q(\counter_r[5] ));
 sg13g2_dfrbp_1 _0976_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net123),
    .D(_0013_),
    .Q_N(_0476_),
    .Q(\counter_r[6] ));
 sg13g2_dfrbp_1 _0977_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net123),
    .D(_0014_),
    .Q_N(_0475_),
    .Q(\counter_r[7] ));
 sg13g2_dfrbp_1 _0978_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net122),
    .D(net48),
    .Q_N(_0005_),
    .Q(\counter_r[8] ));
 sg13g2_dfrbp_1 _0979_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net122),
    .D(_0016_),
    .Q_N(_0474_),
    .Q(\counter_r[9] ));
 sg13g2_dfrbp_1 _0980_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net122),
    .D(net37),
    .Q_N(_0473_),
    .Q(\counter_r[10] ));
 sg13g2_dfrbp_1 _0981_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net122),
    .D(net39),
    .Q_N(_0472_),
    .Q(\counter_r[11] ));
 sg13g2_dfrbp_1 _0982_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net122),
    .D(net32),
    .Q_N(_0471_),
    .Q(\counter_r[12] ));
 sg13g2_dfrbp_1 _0983_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net122),
    .D(_0020_),
    .Q_N(_0470_),
    .Q(\counter_r[13] ));
 sg13g2_dfrbp_1 _0984_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net122),
    .D(net29),
    .Q_N(_0469_),
    .Q(\counter_r[14] ));
 sg13g2_dfrbp_1 _0985_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net122),
    .D(net26),
    .Q_N(_0481_),
    .Q(\counter_r[15] ));
 sg13g2_dfrbp_1 _0986_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net124),
    .D(net21),
    .Q_N(_0482_),
    .Q(\counter_db_r[0] ));
 sg13g2_dfrbp_1 _0987_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net124),
    .D(net44),
    .Q_N(_0483_),
    .Q(\counter_db_r[1] ));
 sg13g2_dfrbp_1 _0988_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net124),
    .D(net24),
    .Q_N(_0484_),
    .Q(\counter_db_r[2] ));
 sg13g2_dfrbp_1 _0989_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net124),
    .D(_0003_),
    .Q_N(_0485_),
    .Q(\counter_db_r[3] ));
 sg13g2_dfrbp_1 _0990_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net125),
    .D(net1),
    .Q_N(_0486_),
    .Q(\count_en_p[0] ));
 sg13g2_dfrbp_1 _0991_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net124),
    .D(net16),
    .Q_N(_0487_),
    .Q(\count_en_p[1] ));
 sg13g2_dfrbp_1 _0992_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net124),
    .D(net17),
    .Q_N(_0488_),
    .Q(\count_en_p[2] ));
 sg13g2_dfrbp_1 _0993_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net124),
    .D(net18),
    .Q_N(_0468_),
    .Q(\count_en_p[3] ));
 sg13g2_dfrbp_1 _0994_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net124),
    .D(net35),
    .Q_N(_0489_),
    .Q(count_en_db_r));
 sg13g2_dfrbp_1 _0995_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net125),
    .D(net19),
    .Q_N(_0467_),
    .Q(count_en_r));
 sg13g2_tiehi tt_um_pyamnihc_dummy_counter_9 (.L_HI(net9));
 sg13g2_tiehi tt_um_pyamnihc_dummy_counter_10 (.L_HI(net10));
 sg13g2_tiehi tt_um_pyamnihc_dummy_counter_11 (.L_HI(net11));
 sg13g2_tiehi tt_um_pyamnihc_dummy_counter_12 (.L_HI(net12));
 sg13g2_tiehi tt_um_pyamnihc_dummy_counter_13 (.L_HI(net13));
 sg13g2_tiehi tt_um_pyamnihc_dummy_counter_14 (.L_HI(net14));
 sg13g2_tiehi tt_um_pyamnihc_dummy_counter_15 (.L_HI(net15));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 fanout95 (.A(_0091_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_0091_),
    .X(net96));
 sg13g2_buf_4 fanout97 (.X(net97),
    .A(_0068_));
 sg13g2_buf_1 fanout98 (.A(_0068_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(net100),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_0093_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(net102),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_0051_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_0050_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_0465_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(net106),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_0064_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_0463_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(net109),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_0448_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(net111),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(net112),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(net56),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(net51),
    .X(net113));
 sg13g2_buf_4 fanout114 (.X(net114),
    .A(\counter_r[0] ));
 sg13g2_buf_1 fanout115 (.A(\counter_r[0] ),
    .X(net115));
 sg13g2_buf_4 fanout116 (.X(net116),
    .A(_0443_));
 sg13g2_buf_2 fanout117 (.A(net121),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(net121),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(net121),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(net121),
    .X(net120));
 sg13g2_buf_1 fanout121 (.A(ui_in[1]),
    .X(net121));
 sg13g2_buf_4 fanout122 (.X(net122),
    .A(rst_n));
 sg13g2_buf_2 fanout123 (.A(rst_n),
    .X(net123));
 sg13g2_buf_4 fanout124 (.X(net124),
    .A(net125));
 sg13g2_buf_2 fanout125 (.A(net126),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(rst_n),
    .X(net126));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[4]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[5]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[6]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[7]),
    .X(net7));
 sg13g2_tiehi tt_um_pyamnihc_dummy_counter_8 (.L_HI(net8));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\count_en_p[0] ),
    .X(net16));
 sg13g2_dlygate4sd3_1 hold2 (.A(\count_en_p[1] ),
    .X(net17));
 sg13g2_dlygate4sd3_1 hold3 (.A(\count_en_p[2] ),
    .X(net18));
 sg13g2_dlygate4sd3_1 hold4 (.A(\count_en_p[3] ),
    .X(net19));
 sg13g2_dlygate4sd3_1 hold5 (.A(\counter_db_r[0] ),
    .X(net20));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0000_),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold7 (.A(\counter_db_r[2] ),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0419_),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0002_),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold10 (.A(\counter_r[15] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0022_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold12 (.A(\counter_r[14] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0437_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0021_),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold15 (.A(\counter_r[12] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0435_),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0019_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold18 (.A(\counter_r[4] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold19 (.A(count_en_r),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0023_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold21 (.A(\counter_r[10] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0017_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold23 (.A(\counter_r[11] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0018_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold25 (.A(\counter_r[13] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold26 (.A(\counter_db_r[3] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0422_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold28 (.A(\counter_db_r[1] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0001_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0006_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0007_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold32 (.A(\counter_r[8] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0015_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold34 (.A(\counter_r[9] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold35 (.A(\counter_r[6] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold36 (.A(\counter_r[1] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0451_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0009_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold39 (.A(\counter_r[5] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold40 (.A(\counter_r[7] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold41 (.A(count_en_db_r),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold42 (.A(\counter_r[3] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0010_),
    .X(net58));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_fill_2 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_160 ();
 sg13g2_decap_8 FILLER_19_167 ();
 sg13g2_decap_4 FILLER_19_174 ();
 sg13g2_fill_1 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_202 ();
 sg13g2_decap_8 FILLER_19_209 ();
 sg13g2_fill_2 FILLER_19_216 ();
 sg13g2_fill_1 FILLER_19_218 ();
 sg13g2_decap_4 FILLER_19_229 ();
 sg13g2_decap_8 FILLER_19_244 ();
 sg13g2_decap_8 FILLER_19_251 ();
 sg13g2_fill_2 FILLER_19_258 ();
 sg13g2_fill_1 FILLER_19_260 ();
 sg13g2_decap_8 FILLER_19_267 ();
 sg13g2_decap_8 FILLER_19_274 ();
 sg13g2_decap_8 FILLER_19_281 ();
 sg13g2_decap_8 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_295 ();
 sg13g2_decap_8 FILLER_19_302 ();
 sg13g2_decap_8 FILLER_19_309 ();
 sg13g2_decap_8 FILLER_19_316 ();
 sg13g2_decap_8 FILLER_19_323 ();
 sg13g2_decap_8 FILLER_19_330 ();
 sg13g2_decap_8 FILLER_19_337 ();
 sg13g2_decap_8 FILLER_19_344 ();
 sg13g2_decap_8 FILLER_19_351 ();
 sg13g2_decap_8 FILLER_19_358 ();
 sg13g2_decap_8 FILLER_19_365 ();
 sg13g2_decap_8 FILLER_19_372 ();
 sg13g2_decap_8 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_fill_2 FILLER_20_133 ();
 sg13g2_fill_2 FILLER_20_152 ();
 sg13g2_fill_2 FILLER_20_167 ();
 sg13g2_fill_1 FILLER_20_169 ();
 sg13g2_decap_8 FILLER_20_183 ();
 sg13g2_fill_1 FILLER_20_190 ();
 sg13g2_decap_8 FILLER_20_205 ();
 sg13g2_fill_1 FILLER_20_212 ();
 sg13g2_decap_8 FILLER_20_283 ();
 sg13g2_decap_8 FILLER_20_290 ();
 sg13g2_decap_8 FILLER_20_297 ();
 sg13g2_decap_8 FILLER_20_304 ();
 sg13g2_decap_8 FILLER_20_311 ();
 sg13g2_decap_8 FILLER_20_318 ();
 sg13g2_decap_8 FILLER_20_325 ();
 sg13g2_decap_8 FILLER_20_332 ();
 sg13g2_decap_8 FILLER_20_339 ();
 sg13g2_decap_8 FILLER_20_346 ();
 sg13g2_decap_8 FILLER_20_353 ();
 sg13g2_decap_8 FILLER_20_360 ();
 sg13g2_decap_8 FILLER_20_367 ();
 sg13g2_decap_8 FILLER_20_374 ();
 sg13g2_decap_8 FILLER_20_381 ();
 sg13g2_decap_8 FILLER_20_388 ();
 sg13g2_decap_8 FILLER_20_395 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_4 FILLER_21_131 ();
 sg13g2_fill_1 FILLER_21_135 ();
 sg13g2_decap_4 FILLER_21_144 ();
 sg13g2_fill_1 FILLER_21_148 ();
 sg13g2_decap_8 FILLER_21_158 ();
 sg13g2_decap_8 FILLER_21_165 ();
 sg13g2_fill_1 FILLER_21_172 ();
 sg13g2_fill_1 FILLER_21_178 ();
 sg13g2_decap_4 FILLER_21_185 ();
 sg13g2_fill_1 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_4 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_4 FILLER_21_231 ();
 sg13g2_fill_2 FILLER_21_235 ();
 sg13g2_fill_2 FILLER_21_246 ();
 sg13g2_decap_8 FILLER_21_253 ();
 sg13g2_fill_2 FILLER_21_260 ();
 sg13g2_fill_1 FILLER_21_262 ();
 sg13g2_fill_2 FILLER_21_274 ();
 sg13g2_decap_8 FILLER_21_288 ();
 sg13g2_decap_8 FILLER_21_295 ();
 sg13g2_decap_8 FILLER_21_302 ();
 sg13g2_decap_8 FILLER_21_309 ();
 sg13g2_decap_8 FILLER_21_316 ();
 sg13g2_decap_8 FILLER_21_323 ();
 sg13g2_decap_8 FILLER_21_330 ();
 sg13g2_decap_8 FILLER_21_337 ();
 sg13g2_decap_8 FILLER_21_344 ();
 sg13g2_decap_8 FILLER_21_351 ();
 sg13g2_decap_8 FILLER_21_358 ();
 sg13g2_decap_8 FILLER_21_365 ();
 sg13g2_decap_8 FILLER_21_372 ();
 sg13g2_decap_8 FILLER_21_379 ();
 sg13g2_decap_8 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_393 ();
 sg13g2_decap_8 FILLER_21_400 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_4 FILLER_22_91 ();
 sg13g2_fill_2 FILLER_22_95 ();
 sg13g2_fill_2 FILLER_22_105 ();
 sg13g2_fill_1 FILLER_22_120 ();
 sg13g2_fill_2 FILLER_22_134 ();
 sg13g2_fill_1 FILLER_22_136 ();
 sg13g2_decap_4 FILLER_22_163 ();
 sg13g2_fill_2 FILLER_22_188 ();
 sg13g2_decap_4 FILLER_22_205 ();
 sg13g2_decap_4 FILLER_22_229 ();
 sg13g2_decap_4 FILLER_22_254 ();
 sg13g2_fill_2 FILLER_22_258 ();
 sg13g2_decap_4 FILLER_22_272 ();
 sg13g2_fill_2 FILLER_22_283 ();
 sg13g2_fill_1 FILLER_22_285 ();
 sg13g2_decap_8 FILLER_22_298 ();
 sg13g2_decap_8 FILLER_22_305 ();
 sg13g2_decap_8 FILLER_22_312 ();
 sg13g2_decap_8 FILLER_22_319 ();
 sg13g2_decap_8 FILLER_22_326 ();
 sg13g2_decap_8 FILLER_22_333 ();
 sg13g2_decap_8 FILLER_22_340 ();
 sg13g2_decap_8 FILLER_22_347 ();
 sg13g2_decap_8 FILLER_22_354 ();
 sg13g2_decap_8 FILLER_22_361 ();
 sg13g2_decap_8 FILLER_22_368 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_129 ();
 sg13g2_decap_4 FILLER_23_136 ();
 sg13g2_decap_4 FILLER_23_160 ();
 sg13g2_fill_1 FILLER_23_164 ();
 sg13g2_decap_8 FILLER_23_170 ();
 sg13g2_fill_1 FILLER_23_177 ();
 sg13g2_fill_2 FILLER_23_183 ();
 sg13g2_fill_1 FILLER_23_185 ();
 sg13g2_decap_8 FILLER_23_205 ();
 sg13g2_fill_1 FILLER_23_212 ();
 sg13g2_decap_4 FILLER_23_229 ();
 sg13g2_fill_2 FILLER_23_233 ();
 sg13g2_fill_1 FILLER_23_257 ();
 sg13g2_fill_1 FILLER_23_265 ();
 sg13g2_fill_2 FILLER_23_274 ();
 sg13g2_fill_1 FILLER_23_276 ();
 sg13g2_fill_2 FILLER_23_287 ();
 sg13g2_fill_1 FILLER_23_289 ();
 sg13g2_decap_8 FILLER_23_302 ();
 sg13g2_decap_8 FILLER_23_309 ();
 sg13g2_decap_8 FILLER_23_316 ();
 sg13g2_decap_8 FILLER_23_323 ();
 sg13g2_decap_8 FILLER_23_330 ();
 sg13g2_decap_8 FILLER_23_337 ();
 sg13g2_decap_8 FILLER_23_344 ();
 sg13g2_decap_8 FILLER_23_351 ();
 sg13g2_decap_8 FILLER_23_358 ();
 sg13g2_decap_8 FILLER_23_365 ();
 sg13g2_decap_8 FILLER_23_372 ();
 sg13g2_decap_8 FILLER_23_379 ();
 sg13g2_decap_8 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_fill_2 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_86 ();
 sg13g2_fill_2 FILLER_24_93 ();
 sg13g2_fill_1 FILLER_24_95 ();
 sg13g2_fill_2 FILLER_24_101 ();
 sg13g2_fill_1 FILLER_24_103 ();
 sg13g2_fill_2 FILLER_24_108 ();
 sg13g2_fill_1 FILLER_24_110 ();
 sg13g2_fill_2 FILLER_24_116 ();
 sg13g2_decap_8 FILLER_24_125 ();
 sg13g2_decap_4 FILLER_24_132 ();
 sg13g2_fill_2 FILLER_24_136 ();
 sg13g2_decap_4 FILLER_24_158 ();
 sg13g2_fill_2 FILLER_24_181 ();
 sg13g2_fill_1 FILLER_24_183 ();
 sg13g2_decap_8 FILLER_24_211 ();
 sg13g2_decap_8 FILLER_24_218 ();
 sg13g2_fill_2 FILLER_24_225 ();
 sg13g2_fill_1 FILLER_24_227 ();
 sg13g2_decap_4 FILLER_24_232 ();
 sg13g2_fill_2 FILLER_24_250 ();
 sg13g2_fill_1 FILLER_24_252 ();
 sg13g2_fill_1 FILLER_24_258 ();
 sg13g2_decap_8 FILLER_24_264 ();
 sg13g2_fill_2 FILLER_24_271 ();
 sg13g2_fill_1 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_fill_2 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_333 ();
 sg13g2_decap_8 FILLER_24_340 ();
 sg13g2_decap_8 FILLER_24_347 ();
 sg13g2_decap_8 FILLER_24_354 ();
 sg13g2_decap_8 FILLER_24_361 ();
 sg13g2_decap_8 FILLER_24_368 ();
 sg13g2_decap_8 FILLER_24_375 ();
 sg13g2_decap_8 FILLER_24_382 ();
 sg13g2_decap_8 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_4 FILLER_24_403 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_4 FILLER_25_70 ();
 sg13g2_fill_2 FILLER_25_74 ();
 sg13g2_fill_1 FILLER_25_92 ();
 sg13g2_decap_8 FILLER_25_114 ();
 sg13g2_fill_1 FILLER_25_121 ();
 sg13g2_decap_4 FILLER_25_142 ();
 sg13g2_fill_1 FILLER_25_146 ();
 sg13g2_decap_8 FILLER_25_158 ();
 sg13g2_fill_1 FILLER_25_189 ();
 sg13g2_fill_1 FILLER_25_194 ();
 sg13g2_decap_8 FILLER_25_205 ();
 sg13g2_fill_2 FILLER_25_212 ();
 sg13g2_fill_1 FILLER_25_214 ();
 sg13g2_fill_1 FILLER_25_234 ();
 sg13g2_decap_4 FILLER_25_240 ();
 sg13g2_decap_4 FILLER_25_270 ();
 sg13g2_fill_1 FILLER_25_274 ();
 sg13g2_fill_2 FILLER_25_285 ();
 sg13g2_fill_1 FILLER_25_287 ();
 sg13g2_fill_2 FILLER_25_312 ();
 sg13g2_fill_1 FILLER_25_314 ();
 sg13g2_decap_8 FILLER_25_341 ();
 sg13g2_decap_8 FILLER_25_348 ();
 sg13g2_decap_8 FILLER_25_355 ();
 sg13g2_decap_8 FILLER_25_362 ();
 sg13g2_decap_8 FILLER_25_369 ();
 sg13g2_decap_8 FILLER_25_376 ();
 sg13g2_decap_8 FILLER_25_383 ();
 sg13g2_decap_8 FILLER_25_390 ();
 sg13g2_decap_8 FILLER_25_397 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_fill_2 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_88 ();
 sg13g2_fill_2 FILLER_26_95 ();
 sg13g2_fill_1 FILLER_26_97 ();
 sg13g2_decap_8 FILLER_26_111 ();
 sg13g2_fill_2 FILLER_26_118 ();
 sg13g2_fill_1 FILLER_26_120 ();
 sg13g2_fill_2 FILLER_26_140 ();
 sg13g2_fill_1 FILLER_26_142 ();
 sg13g2_fill_2 FILLER_26_160 ();
 sg13g2_fill_1 FILLER_26_162 ();
 sg13g2_fill_2 FILLER_26_176 ();
 sg13g2_fill_1 FILLER_26_178 ();
 sg13g2_fill_2 FILLER_26_193 ();
 sg13g2_decap_8 FILLER_26_216 ();
 sg13g2_fill_2 FILLER_26_223 ();
 sg13g2_decap_4 FILLER_26_246 ();
 sg13g2_fill_2 FILLER_26_250 ();
 sg13g2_fill_1 FILLER_26_257 ();
 sg13g2_decap_8 FILLER_26_263 ();
 sg13g2_fill_1 FILLER_26_270 ();
 sg13g2_decap_4 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_296 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_fill_2 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_338 ();
 sg13g2_decap_8 FILLER_26_345 ();
 sg13g2_decap_8 FILLER_26_352 ();
 sg13g2_decap_8 FILLER_26_359 ();
 sg13g2_decap_8 FILLER_26_366 ();
 sg13g2_decap_8 FILLER_26_373 ();
 sg13g2_decap_8 FILLER_26_380 ();
 sg13g2_decap_8 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_fill_1 FILLER_27_70 ();
 sg13g2_decap_4 FILLER_27_92 ();
 sg13g2_decap_4 FILLER_27_121 ();
 sg13g2_fill_1 FILLER_27_125 ();
 sg13g2_decap_4 FILLER_27_140 ();
 sg13g2_fill_2 FILLER_27_144 ();
 sg13g2_fill_2 FILLER_27_160 ();
 sg13g2_fill_1 FILLER_27_162 ();
 sg13g2_fill_2 FILLER_27_168 ();
 sg13g2_fill_2 FILLER_27_182 ();
 sg13g2_fill_1 FILLER_27_184 ();
 sg13g2_decap_4 FILLER_27_189 ();
 sg13g2_fill_1 FILLER_27_193 ();
 sg13g2_decap_4 FILLER_27_214 ();
 sg13g2_decap_4 FILLER_27_236 ();
 sg13g2_fill_2 FILLER_27_240 ();
 sg13g2_decap_4 FILLER_27_268 ();
 sg13g2_fill_2 FILLER_27_272 ();
 sg13g2_decap_8 FILLER_27_288 ();
 sg13g2_fill_2 FILLER_27_295 ();
 sg13g2_fill_2 FILLER_27_322 ();
 sg13g2_decap_8 FILLER_27_340 ();
 sg13g2_decap_8 FILLER_27_347 ();
 sg13g2_decap_8 FILLER_27_354 ();
 sg13g2_decap_8 FILLER_27_361 ();
 sg13g2_decap_8 FILLER_27_368 ();
 sg13g2_decap_8 FILLER_27_375 ();
 sg13g2_decap_8 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_27_396 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_4 FILLER_28_70 ();
 sg13g2_fill_2 FILLER_28_74 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_fill_1 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_115 ();
 sg13g2_fill_2 FILLER_28_122 ();
 sg13g2_fill_1 FILLER_28_124 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_fill_2 FILLER_28_147 ();
 sg13g2_fill_1 FILLER_28_149 ();
 sg13g2_fill_1 FILLER_28_156 ();
 sg13g2_fill_2 FILLER_28_165 ();
 sg13g2_fill_1 FILLER_28_171 ();
 sg13g2_fill_2 FILLER_28_180 ();
 sg13g2_decap_4 FILLER_28_190 ();
 sg13g2_decap_4 FILLER_28_199 ();
 sg13g2_fill_2 FILLER_28_215 ();
 sg13g2_fill_1 FILLER_28_217 ();
 sg13g2_decap_4 FILLER_28_233 ();
 sg13g2_decap_8 FILLER_28_241 ();
 sg13g2_decap_8 FILLER_28_263 ();
 sg13g2_fill_1 FILLER_28_270 ();
 sg13g2_decap_8 FILLER_28_294 ();
 sg13g2_decap_4 FILLER_28_311 ();
 sg13g2_decap_8 FILLER_28_335 ();
 sg13g2_decap_8 FILLER_28_342 ();
 sg13g2_decap_8 FILLER_28_349 ();
 sg13g2_decap_8 FILLER_28_356 ();
 sg13g2_decap_8 FILLER_28_363 ();
 sg13g2_decap_8 FILLER_28_370 ();
 sg13g2_decap_8 FILLER_28_377 ();
 sg13g2_decap_8 FILLER_28_384 ();
 sg13g2_decap_8 FILLER_28_391 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_fill_2 FILLER_29_95 ();
 sg13g2_fill_1 FILLER_29_97 ();
 sg13g2_decap_8 FILLER_29_111 ();
 sg13g2_fill_2 FILLER_29_118 ();
 sg13g2_fill_1 FILLER_29_120 ();
 sg13g2_fill_2 FILLER_29_139 ();
 sg13g2_fill_1 FILLER_29_141 ();
 sg13g2_fill_1 FILLER_29_158 ();
 sg13g2_decap_8 FILLER_29_163 ();
 sg13g2_decap_8 FILLER_29_170 ();
 sg13g2_decap_4 FILLER_29_177 ();
 sg13g2_fill_2 FILLER_29_189 ();
 sg13g2_fill_1 FILLER_29_191 ();
 sg13g2_fill_2 FILLER_29_205 ();
 sg13g2_fill_1 FILLER_29_207 ();
 sg13g2_decap_8 FILLER_29_228 ();
 sg13g2_fill_2 FILLER_29_235 ();
 sg13g2_fill_1 FILLER_29_237 ();
 sg13g2_decap_8 FILLER_29_260 ();
 sg13g2_decap_8 FILLER_29_267 ();
 sg13g2_fill_1 FILLER_29_274 ();
 sg13g2_decap_8 FILLER_29_286 ();
 sg13g2_fill_1 FILLER_29_293 ();
 sg13g2_decap_4 FILLER_29_298 ();
 sg13g2_decap_8 FILLER_29_320 ();
 sg13g2_decap_8 FILLER_29_327 ();
 sg13g2_decap_8 FILLER_29_334 ();
 sg13g2_decap_8 FILLER_29_341 ();
 sg13g2_decap_8 FILLER_29_348 ();
 sg13g2_decap_8 FILLER_29_355 ();
 sg13g2_decap_8 FILLER_29_362 ();
 sg13g2_decap_8 FILLER_29_369 ();
 sg13g2_decap_8 FILLER_29_376 ();
 sg13g2_decap_8 FILLER_29_383 ();
 sg13g2_decap_8 FILLER_29_390 ();
 sg13g2_decap_8 FILLER_29_397 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_4 FILLER_30_63 ();
 sg13g2_fill_2 FILLER_30_67 ();
 sg13g2_fill_1 FILLER_30_96 ();
 sg13g2_fill_2 FILLER_30_125 ();
 sg13g2_fill_1 FILLER_30_127 ();
 sg13g2_decap_4 FILLER_30_137 ();
 sg13g2_fill_1 FILLER_30_150 ();
 sg13g2_fill_2 FILLER_30_175 ();
 sg13g2_fill_1 FILLER_30_177 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_fill_2 FILLER_30_189 ();
 sg13g2_fill_1 FILLER_30_191 ();
 sg13g2_decap_8 FILLER_30_204 ();
 sg13g2_decap_4 FILLER_30_211 ();
 sg13g2_fill_1 FILLER_30_215 ();
 sg13g2_decap_4 FILLER_30_258 ();
 sg13g2_fill_2 FILLER_30_274 ();
 sg13g2_fill_1 FILLER_30_276 ();
 sg13g2_decap_4 FILLER_30_304 ();
 sg13g2_decap_8 FILLER_30_319 ();
 sg13g2_decap_8 FILLER_30_326 ();
 sg13g2_decap_8 FILLER_30_333 ();
 sg13g2_decap_8 FILLER_30_340 ();
 sg13g2_decap_8 FILLER_30_347 ();
 sg13g2_decap_8 FILLER_30_354 ();
 sg13g2_decap_8 FILLER_30_361 ();
 sg13g2_decap_8 FILLER_30_368 ();
 sg13g2_decap_8 FILLER_30_375 ();
 sg13g2_decap_8 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_30_389 ();
 sg13g2_decap_8 FILLER_30_396 ();
 sg13g2_decap_4 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_fill_1 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_92 ();
 sg13g2_decap_8 FILLER_31_99 ();
 sg13g2_fill_2 FILLER_31_106 ();
 sg13g2_decap_4 FILLER_31_117 ();
 sg13g2_fill_1 FILLER_31_121 ();
 sg13g2_fill_1 FILLER_31_143 ();
 sg13g2_decap_4 FILLER_31_152 ();
 sg13g2_fill_2 FILLER_31_156 ();
 sg13g2_decap_4 FILLER_31_162 ();
 sg13g2_fill_1 FILLER_31_166 ();
 sg13g2_fill_2 FILLER_31_186 ();
 sg13g2_decap_4 FILLER_31_209 ();
 sg13g2_fill_1 FILLER_31_213 ();
 sg13g2_decap_8 FILLER_31_233 ();
 sg13g2_decap_8 FILLER_31_240 ();
 sg13g2_fill_1 FILLER_31_247 ();
 sg13g2_decap_8 FILLER_31_275 ();
 sg13g2_fill_2 FILLER_31_282 ();
 sg13g2_fill_1 FILLER_31_284 ();
 sg13g2_decap_8 FILLER_31_290 ();
 sg13g2_fill_2 FILLER_31_297 ();
 sg13g2_fill_1 FILLER_31_304 ();
 sg13g2_decap_8 FILLER_31_323 ();
 sg13g2_decap_8 FILLER_31_330 ();
 sg13g2_fill_1 FILLER_31_337 ();
 sg13g2_decap_8 FILLER_31_342 ();
 sg13g2_decap_8 FILLER_31_349 ();
 sg13g2_decap_8 FILLER_31_356 ();
 sg13g2_decap_8 FILLER_31_363 ();
 sg13g2_decap_8 FILLER_31_370 ();
 sg13g2_decap_8 FILLER_31_377 ();
 sg13g2_decap_8 FILLER_31_384 ();
 sg13g2_decap_8 FILLER_31_391 ();
 sg13g2_decap_8 FILLER_31_398 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_fill_2 FILLER_32_56 ();
 sg13g2_fill_1 FILLER_32_58 ();
 sg13g2_decap_4 FILLER_32_68 ();
 sg13g2_decap_4 FILLER_32_93 ();
 sg13g2_decap_4 FILLER_32_125 ();
 sg13g2_fill_1 FILLER_32_129 ();
 sg13g2_decap_4 FILLER_32_134 ();
 sg13g2_fill_1 FILLER_32_138 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_fill_2 FILLER_32_154 ();
 sg13g2_fill_1 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_173 ();
 sg13g2_fill_1 FILLER_32_180 ();
 sg13g2_decap_4 FILLER_32_189 ();
 sg13g2_fill_1 FILLER_32_193 ();
 sg13g2_decap_8 FILLER_32_207 ();
 sg13g2_decap_4 FILLER_32_214 ();
 sg13g2_fill_1 FILLER_32_218 ();
 sg13g2_decap_4 FILLER_32_239 ();
 sg13g2_fill_2 FILLER_32_248 ();
 sg13g2_fill_1 FILLER_32_250 ();
 sg13g2_fill_2 FILLER_32_274 ();
 sg13g2_fill_2 FILLER_32_292 ();
 sg13g2_fill_2 FILLER_32_307 ();
 sg13g2_fill_1 FILLER_32_309 ();
 sg13g2_decap_8 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_decap_8 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_fill_2 FILLER_33_49 ();
 sg13g2_fill_2 FILLER_33_90 ();
 sg13g2_fill_2 FILLER_33_104 ();
 sg13g2_fill_1 FILLER_33_106 ();
 sg13g2_fill_1 FILLER_33_137 ();
 sg13g2_fill_1 FILLER_33_150 ();
 sg13g2_fill_2 FILLER_33_166 ();
 sg13g2_fill_1 FILLER_33_168 ();
 sg13g2_decap_4 FILLER_33_174 ();
 sg13g2_fill_2 FILLER_33_178 ();
 sg13g2_decap_8 FILLER_33_194 ();
 sg13g2_fill_2 FILLER_33_211 ();
 sg13g2_fill_2 FILLER_33_223 ();
 sg13g2_fill_2 FILLER_33_237 ();
 sg13g2_fill_1 FILLER_33_239 ();
 sg13g2_fill_2 FILLER_33_258 ();
 sg13g2_fill_1 FILLER_33_260 ();
 sg13g2_fill_2 FILLER_33_277 ();
 sg13g2_fill_1 FILLER_33_279 ();
 sg13g2_fill_1 FILLER_33_312 ();
 sg13g2_decap_8 FILLER_33_379 ();
 sg13g2_decap_8 FILLER_33_386 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_4 FILLER_34_49 ();
 sg13g2_fill_2 FILLER_34_67 ();
 sg13g2_decap_8 FILLER_34_78 ();
 sg13g2_fill_1 FILLER_34_85 ();
 sg13g2_fill_1 FILLER_34_96 ();
 sg13g2_decap_4 FILLER_34_144 ();
 sg13g2_fill_2 FILLER_34_148 ();
 sg13g2_fill_2 FILLER_34_160 ();
 sg13g2_fill_1 FILLER_34_170 ();
 sg13g2_fill_1 FILLER_34_215 ();
 sg13g2_fill_1 FILLER_34_245 ();
 sg13g2_fill_2 FILLER_34_255 ();
 sg13g2_fill_1 FILLER_34_292 ();
 sg13g2_decap_8 FILLER_34_316 ();
 sg13g2_fill_1 FILLER_34_349 ();
 sg13g2_decap_8 FILLER_34_382 ();
 sg13g2_decap_8 FILLER_34_389 ();
 sg13g2_decap_8 FILLER_34_396 ();
 sg13g2_decap_4 FILLER_34_403 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_fill_2 FILLER_35_112 ();
 sg13g2_fill_1 FILLER_35_114 ();
 sg13g2_fill_2 FILLER_35_141 ();
 sg13g2_fill_2 FILLER_35_186 ();
 sg13g2_fill_2 FILLER_35_199 ();
 sg13g2_fill_1 FILLER_35_201 ();
 sg13g2_fill_2 FILLER_35_211 ();
 sg13g2_fill_2 FILLER_35_223 ();
 sg13g2_fill_1 FILLER_35_225 ();
 sg13g2_fill_1 FILLER_35_235 ();
 sg13g2_fill_2 FILLER_35_244 ();
 sg13g2_fill_1 FILLER_35_246 ();
 sg13g2_fill_2 FILLER_35_261 ();
 sg13g2_fill_1 FILLER_35_263 ();
 sg13g2_fill_1 FILLER_35_287 ();
 sg13g2_fill_2 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_390 ();
 sg13g2_decap_8 FILLER_35_397 ();
 sg13g2_decap_4 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_fill_2 FILLER_36_82 ();
 sg13g2_fill_1 FILLER_36_124 ();
 sg13g2_decap_8 FILLER_36_132 ();
 sg13g2_fill_2 FILLER_36_139 ();
 sg13g2_fill_1 FILLER_36_141 ();
 sg13g2_decap_8 FILLER_36_165 ();
 sg13g2_decap_8 FILLER_36_172 ();
 sg13g2_fill_1 FILLER_36_179 ();
 sg13g2_fill_2 FILLER_36_306 ();
 sg13g2_fill_1 FILLER_36_308 ();
 sg13g2_fill_2 FILLER_36_340 ();
 sg13g2_fill_1 FILLER_36_352 ();
 sg13g2_decap_8 FILLER_36_397 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_4 FILLER_37_56 ();
 sg13g2_fill_2 FILLER_37_60 ();
 sg13g2_decap_8 FILLER_37_88 ();
 sg13g2_decap_4 FILLER_37_95 ();
 sg13g2_fill_1 FILLER_37_99 ();
 sg13g2_decap_8 FILLER_37_134 ();
 sg13g2_decap_8 FILLER_37_141 ();
 sg13g2_fill_1 FILLER_37_148 ();
 sg13g2_decap_4 FILLER_37_200 ();
 sg13g2_decap_4 FILLER_37_213 ();
 sg13g2_fill_2 FILLER_37_217 ();
 sg13g2_decap_4 FILLER_37_224 ();
 sg13g2_fill_1 FILLER_37_228 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_fill_2 FILLER_37_245 ();
 sg13g2_fill_1 FILLER_37_247 ();
 sg13g2_fill_2 FILLER_37_253 ();
 sg13g2_fill_1 FILLER_37_255 ();
 sg13g2_fill_2 FILLER_37_274 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_fill_1 FILLER_38_68 ();
 sg13g2_fill_2 FILLER_38_86 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_163 ();
 sg13g2_decap_8 FILLER_38_170 ();
 sg13g2_decap_8 FILLER_38_177 ();
 sg13g2_decap_4 FILLER_38_187 ();
 sg13g2_fill_1 FILLER_38_191 ();
 sg13g2_decap_4 FILLER_38_218 ();
 sg13g2_fill_2 FILLER_38_283 ();
 sg13g2_fill_1 FILLER_38_285 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net8;
 assign uio_oe[1] = net9;
 assign uio_oe[2] = net10;
 assign uio_oe[3] = net11;
 assign uio_oe[4] = net12;
 assign uio_oe[5] = net13;
 assign uio_oe[6] = net14;
 assign uio_oe[7] = net15;
endmodule

module tt_um_toivoh_demo_deluxe (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire advance_frame;
 wire \dtop.detune_counter[10] ;
 wire \dtop.detune_counter[11] ;
 wire \dtop.detune_counter[12] ;
 wire \dtop.detune_counter[13] ;
 wire \dtop.detune_counter[14] ;
 wire \dtop.detune_counter[15] ;
 wire \dtop.detune_counter[16] ;
 wire \dtop.detune_counter[17] ;
 wire \dtop.detune_counter[4] ;
 wire \dtop.detune_counter[5] ;
 wire \dtop.detune_counter[6] ;
 wire \dtop.detune_counter[7] ;
 wire \dtop.detune_counter[8] ;
 wire \dtop.detune_counter[9] ;
 wire \dtop.enable ;
 wire \dtop.ext_control[0] ;
 wire \dtop.ext_control[1] ;
 wire \dtop.ext_control[2] ;
 wire \dtop.ext_control[3] ;
 wire \dtop.ext_control[4] ;
 wire \dtop.ext_control[5] ;
 wire \dtop.ext_control[6] ;
 wire \dtop.oct_counter[0] ;
 wire \dtop.oct_counter[1] ;
 wire \dtop.oct_counter[2] ;
 wire \dtop.oct_counter[3] ;
 wire \dtop.oct_counter[4] ;
 wire \dtop.oct_counter[5] ;
 wire \dtop.oct_counter[6] ;
 wire \dtop.out_sample[0] ;
 wire \dtop.out_sample[1] ;
 wire \dtop.out_sample[2] ;
 wire \dtop.out_sample[3] ;
 wire \dtop.out_sample[4] ;
 wire \dtop.out_sample[5] ;
 wire \dtop.out_sample[6] ;
 wire \dtop.player_inst.program_addr[0] ;
 wire \dtop.player_inst.program_addr[1] ;
 wire \dtop.player_inst.program_addr[2] ;
 wire \dtop.player_inst.program_addr[3] ;
 wire \dtop.player_inst.program_addr[4] ;
 wire \dtop.player_inst.program_addr[5] ;
 wire \dtop.player_inst.program_addr[6] ;
 wire \dtop.player_inst.synth.alu.acc[0] ;
 wire \dtop.player_inst.synth.alu.acc[10] ;
 wire \dtop.player_inst.synth.alu.acc[1] ;
 wire \dtop.player_inst.synth.alu.acc[2] ;
 wire \dtop.player_inst.synth.alu.acc[3] ;
 wire \dtop.player_inst.synth.alu.acc[4] ;
 wire \dtop.player_inst.synth.alu.acc[5] ;
 wire \dtop.player_inst.synth.alu.acc[6] ;
 wire \dtop.player_inst.synth.alu.acc[7] ;
 wire \dtop.player_inst.synth.alu.acc[8] ;
 wire \dtop.player_inst.synth.alu.acc[9] ;
 wire \dtop.player_inst.synth.alu.carry ;
 wire \dtop.player_inst.synth.alu.oct_en ;
 wire \dtop.player_inst.synth.alu.registers[0][0] ;
 wire \dtop.player_inst.synth.alu.registers[0][10] ;
 wire \dtop.player_inst.synth.alu.registers[0][1] ;
 wire \dtop.player_inst.synth.alu.registers[0][2] ;
 wire \dtop.player_inst.synth.alu.registers[0][3] ;
 wire \dtop.player_inst.synth.alu.registers[0][4] ;
 wire \dtop.player_inst.synth.alu.registers[0][5] ;
 wire \dtop.player_inst.synth.alu.registers[0][6] ;
 wire \dtop.player_inst.synth.alu.registers[0][7] ;
 wire \dtop.player_inst.synth.alu.registers[0][8] ;
 wire \dtop.player_inst.synth.alu.registers[0][9] ;
 wire \dtop.player_inst.synth.alu.registers[1][0] ;
 wire \dtop.player_inst.synth.alu.registers[1][10] ;
 wire \dtop.player_inst.synth.alu.registers[1][1] ;
 wire \dtop.player_inst.synth.alu.registers[1][2] ;
 wire \dtop.player_inst.synth.alu.registers[1][3] ;
 wire \dtop.player_inst.synth.alu.registers[1][4] ;
 wire \dtop.player_inst.synth.alu.registers[1][5] ;
 wire \dtop.player_inst.synth.alu.registers[1][6] ;
 wire \dtop.player_inst.synth.alu.registers[1][7] ;
 wire \dtop.player_inst.synth.alu.registers[1][8] ;
 wire \dtop.player_inst.synth.alu.registers[1][9] ;
 wire \dtop.player_inst.synth.alu.registers[2][0] ;
 wire \dtop.player_inst.synth.alu.registers[2][1] ;
 wire \dtop.player_inst.synth.alu.registers[2][2] ;
 wire \dtop.player_inst.synth.alu.registers[2][3] ;
 wire \dtop.player_inst.synth.alu.registers[2][4] ;
 wire \dtop.player_inst.synth.alu.registers[2][5] ;
 wire \dtop.player_inst.synth.alu.registers[2][6] ;
 wire \dtop.player_inst.synth.alu.registers[2][7] ;
 wire \dtop.player_inst.synth.alu.registers[3][0] ;
 wire \dtop.player_inst.synth.alu.registers[3][1] ;
 wire \dtop.player_inst.synth.alu.registers[3][2] ;
 wire \dtop.player_inst.synth.alu.registers[3][3] ;
 wire \dtop.player_inst.synth.alu.registers[3][4] ;
 wire \dtop.player_inst.synth.alu.registers[3][5] ;
 wire \dtop.player_inst.synth.alu.registers[3][6] ;
 wire \dtop.player_inst.synth.alu.registers[3][7] ;
 wire \dtop.player_inst.synth.alu.registers[4][0] ;
 wire \dtop.player_inst.synth.alu.registers[4][10] ;
 wire \dtop.player_inst.synth.alu.registers[4][1] ;
 wire \dtop.player_inst.synth.alu.registers[4][2] ;
 wire \dtop.player_inst.synth.alu.registers[4][3] ;
 wire \dtop.player_inst.synth.alu.registers[4][4] ;
 wire \dtop.player_inst.synth.alu.registers[4][5] ;
 wire \dtop.player_inst.synth.alu.registers[4][6] ;
 wire \dtop.player_inst.synth.alu.registers[4][7] ;
 wire \dtop.player_inst.synth.alu.registers[4][8] ;
 wire \dtop.player_inst.synth.alu.registers[4][9] ;
 wire \dtop.player_inst.synth.alu.registers[5][0] ;
 wire \dtop.player_inst.synth.alu.registers[5][1] ;
 wire \dtop.player_inst.synth.alu.registers[5][2] ;
 wire \dtop.player_inst.synth.alu.registers[5][3] ;
 wire \dtop.player_inst.synth.alu.registers[5][4] ;
 wire \dtop.player_inst.synth.alu.registers[5][5] ;
 wire \dtop.player_inst.synth.alu.registers[5][6] ;
 wire \dtop.vsync ;
 wire \dtop.vtop.color[10] ;
 wire \dtop.vtop.color[11] ;
 wire \dtop.vtop.color[6] ;
 wire \dtop.vtop.color[7] ;
 wire \dtop.vtop.color[8] ;
 wire \dtop.vtop.color[9] ;
 wire \dtop.vtop.dphases[0][0] ;
 wire \dtop.vtop.dphases[0][10] ;
 wire \dtop.vtop.dphases[0][1] ;
 wire \dtop.vtop.dphases[0][2] ;
 wire \dtop.vtop.dphases[0][3] ;
 wire \dtop.vtop.dphases[0][4] ;
 wire \dtop.vtop.dphases[0][5] ;
 wire \dtop.vtop.dphases[0][6] ;
 wire \dtop.vtop.dphases[0][7] ;
 wire \dtop.vtop.dphases[0][8] ;
 wire \dtop.vtop.dphases[0][9] ;
 wire \dtop.vtop.dphases[1][0] ;
 wire \dtop.vtop.dphases[1][10] ;
 wire \dtop.vtop.dphases[1][1] ;
 wire \dtop.vtop.dphases[1][2] ;
 wire \dtop.vtop.dphases[1][3] ;
 wire \dtop.vtop.dphases[1][4] ;
 wire \dtop.vtop.dphases[1][5] ;
 wire \dtop.vtop.dphases[1][6] ;
 wire \dtop.vtop.dphases[1][7] ;
 wire \dtop.vtop.dphases[1][8] ;
 wire \dtop.vtop.dphases[1][9] ;
 wire \dtop.vtop.dphases[2][0] ;
 wire \dtop.vtop.dphases[2][10] ;
 wire \dtop.vtop.dphases[2][1] ;
 wire \dtop.vtop.dphases[2][2] ;
 wire \dtop.vtop.dphases[2][3] ;
 wire \dtop.vtop.dphases[2][4] ;
 wire \dtop.vtop.dphases[2][5] ;
 wire \dtop.vtop.dphases[2][6] ;
 wire \dtop.vtop.dphases[2][7] ;
 wire \dtop.vtop.dphases[2][8] ;
 wire \dtop.vtop.dphases[2][9] ;
 wire \dtop.vtop.force_sat0 ;
 wire \dtop.vtop.logo.addr[10] ;
 wire \dtop.vtop.logo.addr[11] ;
 wire \dtop.vtop.logo.addr[7] ;
 wire \dtop.vtop.logo.addr[8] ;
 wire \dtop.vtop.logo.addr[9] ;
 wire \dtop.vtop.logo_d[1] ;
 wire \dtop.vtop.pipeline.cosappr_acc[0] ;
 wire \dtop.vtop.pipeline.cosappr_acc[1] ;
 wire \dtop.vtop.pipeline.cosappr_acc[2] ;
 wire \dtop.vtop.pipeline.cosappr_acc[3] ;
 wire \dtop.vtop.pipeline.cosappr_acc[4] ;
 wire \dtop.vtop.pipeline.cosappr_acc[5] ;
 wire \dtop.vtop.pipeline.cosappr_acc[6] ;
 wire \dtop.vtop.pipeline.cosappr_acc[7] ;
 wire \dtop.vtop.pipeline.cosappr_acc[8] ;
 wire \dtop.vtop.pipeline.dz[0] ;
 wire \dtop.vtop.pipeline.dz[1] ;
 wire \dtop.vtop.pipeline.dz[2] ;
 wire \dtop.vtop.pipeline.dz[3] ;
 wire \dtop.vtop.pipeline.dz[4] ;
 wire \dtop.vtop.pipeline.dz[5] ;
 wire \dtop.vtop.pipeline.dz[6] ;
 wire \dtop.vtop.pipeline.dz[7] ;
 wire \dtop.vtop.pipeline.dz[8] ;
 wire \dtop.vtop.pipeline.neg_t[0] ;
 wire \dtop.vtop.pipeline.neg_t[1] ;
 wire \dtop.vtop.pipeline.neg_t[2] ;
 wire \dtop.vtop.pipeline.neg_t[3] ;
 wire \dtop.vtop.pipeline.neg_t[4] ;
 wire \dtop.vtop.pipeline.neg_t[5] ;
 wire \dtop.vtop.pipeline.neg_t[6] ;
 wire \dtop.vtop.pipeline.neg_t[7] ;
 wire \dtop.vtop.pipeline.neg_t[8] ;
 wire \dtop.vtop.pipeline.neg_t[9] ;
 wire \dtop.vtop.pipeline.next_nstep_counter[0] ;
 wire \dtop.vtop.pipeline.nstep[0] ;
 wire \dtop.vtop.pipeline.nstep[1] ;
 wire \dtop.vtop.pipeline.nstep_counter[0] ;
 wire \dtop.vtop.pipeline.nstep_counter[1] ;
 wire \dtop.vtop.pipeline.nstep_counter[2] ;
 wire \dtop.vtop.pipeline.nstep_counter[3] ;
 wire \dtop.vtop.pipeline.nstep_counter[4] ;
 wire \dtop.vtop.pipeline.nstep_zg[0] ;
 wire \dtop.vtop.pipeline.nstep_zg[1] ;
 wire \dtop.vtop.pipeline.phases[0][0] ;
 wire \dtop.vtop.pipeline.phases[0][10] ;
 wire \dtop.vtop.pipeline.phases[0][11] ;
 wire \dtop.vtop.pipeline.phases[0][12] ;
 wire \dtop.vtop.pipeline.phases[0][13] ;
 wire \dtop.vtop.pipeline.phases[0][14] ;
 wire \dtop.vtop.pipeline.phases[0][15] ;
 wire \dtop.vtop.pipeline.phases[0][1] ;
 wire \dtop.vtop.pipeline.phases[0][2] ;
 wire \dtop.vtop.pipeline.phases[0][3] ;
 wire \dtop.vtop.pipeline.phases[0][4] ;
 wire \dtop.vtop.pipeline.phases[0][5] ;
 wire \dtop.vtop.pipeline.phases[0][6] ;
 wire \dtop.vtop.pipeline.phases[0][7] ;
 wire \dtop.vtop.pipeline.phases[0][8] ;
 wire \dtop.vtop.pipeline.phases[0][9] ;
 wire \dtop.vtop.pipeline.phases[1][0] ;
 wire \dtop.vtop.pipeline.phases[1][10] ;
 wire \dtop.vtop.pipeline.phases[1][11] ;
 wire \dtop.vtop.pipeline.phases[1][12] ;
 wire \dtop.vtop.pipeline.phases[1][13] ;
 wire \dtop.vtop.pipeline.phases[1][14] ;
 wire \dtop.vtop.pipeline.phases[1][15] ;
 wire \dtop.vtop.pipeline.phases[1][1] ;
 wire \dtop.vtop.pipeline.phases[1][2] ;
 wire \dtop.vtop.pipeline.phases[1][3] ;
 wire \dtop.vtop.pipeline.phases[1][4] ;
 wire \dtop.vtop.pipeline.phases[1][5] ;
 wire \dtop.vtop.pipeline.phases[1][6] ;
 wire \dtop.vtop.pipeline.phases[1][7] ;
 wire \dtop.vtop.pipeline.phases[1][8] ;
 wire \dtop.vtop.pipeline.phases[1][9] ;
 wire \dtop.vtop.pipeline.phases[2][0] ;
 wire \dtop.vtop.pipeline.phases[2][10] ;
 wire \dtop.vtop.pipeline.phases[2][11] ;
 wire \dtop.vtop.pipeline.phases[2][12] ;
 wire \dtop.vtop.pipeline.phases[2][13] ;
 wire \dtop.vtop.pipeline.phases[2][14] ;
 wire \dtop.vtop.pipeline.phases[2][15] ;
 wire \dtop.vtop.pipeline.phases[2][1] ;
 wire \dtop.vtop.pipeline.phases[2][2] ;
 wire \dtop.vtop.pipeline.phases[2][3] ;
 wire \dtop.vtop.pipeline.phases[2][4] ;
 wire \dtop.vtop.pipeline.phases[2][5] ;
 wire \dtop.vtop.pipeline.phases[2][6] ;
 wire \dtop.vtop.pipeline.phases[2][7] ;
 wire \dtop.vtop.pipeline.phases[2][8] ;
 wire \dtop.vtop.pipeline.phases[2][9] ;
 wire \dtop.vtop.pipeline.wave_index[0] ;
 wire \dtop.vtop.pipeline.wave_index[1] ;
 wire \dtop.vtop.pipeline.z[0] ;
 wire \dtop.vtop.pipeline.z[10] ;
 wire \dtop.vtop.pipeline.z[11] ;
 wire \dtop.vtop.pipeline.z[12] ;
 wire \dtop.vtop.pipeline.z[13] ;
 wire \dtop.vtop.pipeline.z[14] ;
 wire \dtop.vtop.pipeline.z[1] ;
 wire \dtop.vtop.pipeline.z[2] ;
 wire \dtop.vtop.pipeline.z[3] ;
 wire \dtop.vtop.pipeline.z[4] ;
 wire \dtop.vtop.pipeline.z[5] ;
 wire \dtop.vtop.pipeline.z[6] ;
 wire \dtop.vtop.pipeline.z[7] ;
 wire \dtop.vtop.pipeline.z[8] ;
 wire \dtop.vtop.pipeline.z[9] ;
 wire \dtop.vtop.pipeline.zg[0] ;
 wire \dtop.vtop.pipeline.zg[1] ;
 wire \dtop.vtop.pipeline.zg[2] ;
 wire \dtop.vtop.pipeline.zg[3] ;
 wire \dtop.vtop.pipeline.zg[4] ;
 wire \dtop.vtop.pipeline.zg[5] ;
 wire \dtop.vtop.pipeline.zg[6] ;
 wire \dtop.vtop.pipeline.zg[7] ;
 wire \dtop.vtop.pipeline.zg[8] ;
 wire \dtop.vtop.pipeline.zg[9] ;
 wire \dtop.vtop.pipeline.zg_acc[0] ;
 wire \dtop.vtop.pipeline.zg_acc[1] ;
 wire \dtop.vtop.pipeline.zg_acc[2] ;
 wire \dtop.vtop.pipeline.zg_acc[3] ;
 wire \dtop.vtop.pipeline.zg_acc[4] ;
 wire \dtop.vtop.pipeline.zg_acc[5] ;
 wire \dtop.vtop.pipeline.zg_acc[6] ;
 wire \dtop.vtop.pipeline.zg_acc[7] ;
 wire \dtop.vtop.pipeline.zg_acc[8] ;
 wire \dtop.vtop.pipeline.zg_acc[9] ;
 wire \dtop.vtop.pipeline.zg_valid ;
 wire \dtop.vtop.rs.saturated ;
 wire \dtop.vtop.rs.scan_y.phase[0] ;
 wire \dtop.vtop.rs.scan_y.phase[1] ;
 wire \dtop.vtop.rs.x_scan.phase[0] ;
 wire \dtop.vtop.rs.x_scan.phase[1] ;
 wire rst_n_reg;
 wire net317;
 wire clknet_leaf_0_clk;
 wire \uio_out0b[5] ;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;

 sg13g2_inv_1 _3863_ (.Y(_3063_),
    .A(net318));
 sg13g2_inv_1 _3864_ (.Y(_3064_),
    .A(\dtop.vtop.pipeline.zg_valid ));
 sg13g2_inv_1 _3865_ (.Y(_3065_),
    .A(\dtop.vtop.pipeline.z[14] ));
 sg13g2_inv_1 _3866_ (.Y(_3066_),
    .A(net629));
 sg13g2_inv_1 _3867_ (.Y(_3067_),
    .A(\dtop.vtop.pipeline.z[12] ));
 sg13g2_inv_1 _3868_ (.Y(_3068_),
    .A(\dtop.vtop.pipeline.z[11] ));
 sg13g2_inv_1 _3869_ (.Y(_3069_),
    .A(\dtop.vtop.pipeline.z[10] ));
 sg13g2_inv_1 _3870_ (.Y(_3070_),
    .A(\dtop.vtop.pipeline.z[9] ));
 sg13g2_inv_1 _3871_ (.Y(_3071_),
    .A(\dtop.vtop.pipeline.z[8] ));
 sg13g2_inv_1 _3872_ (.Y(_3072_),
    .A(\dtop.vtop.pipeline.z[7] ));
 sg13g2_inv_1 _3873_ (.Y(_3073_),
    .A(\dtop.vtop.pipeline.dz[0] ));
 sg13g2_inv_1 _3874_ (.Y(_3074_),
    .A(\dtop.vtop.pipeline.neg_t[6] ));
 sg13g2_inv_1 _3875_ (.Y(_3075_),
    .A(\dtop.vtop.pipeline.neg_t[1] ));
 sg13g2_inv_1 _3876_ (.Y(_3076_),
    .A(net1408));
 sg13g2_inv_1 _3877_ (.Y(_3077_),
    .A(\dtop.player_inst.synth.alu.acc[6] ));
 sg13g2_inv_2 _3878_ (.Y(_3078_),
    .A(\dtop.player_inst.synth.alu.acc[5] ));
 sg13g2_inv_1 _3879_ (.Y(_3079_),
    .A(net1410));
 sg13g2_inv_1 _3880_ (.Y(_3080_),
    .A(net1411));
 sg13g2_inv_1 _3881_ (.Y(_3081_),
    .A(net1412));
 sg13g2_inv_1 _3882_ (.Y(_3082_),
    .A(\dtop.player_inst.synth.alu.acc[1] ));
 sg13g2_inv_1 _3883_ (.Y(_3083_),
    .A(net1414));
 sg13g2_inv_1 _3884_ (.Y(_3084_),
    .A(net383));
 sg13g2_inv_1 _3885_ (.Y(_3085_),
    .A(net430));
 sg13g2_inv_1 _3886_ (.Y(_3086_),
    .A(net402));
 sg13g2_inv_1 _3887_ (.Y(_3087_),
    .A(net404));
 sg13g2_inv_1 _3888_ (.Y(_3088_),
    .A(net437));
 sg13g2_inv_1 _3889_ (.Y(_3089_),
    .A(net427));
 sg13g2_inv_1 _3890_ (.Y(_3090_),
    .A(net368));
 sg13g2_inv_1 _3891_ (.Y(_3091_),
    .A(net447));
 sg13g2_inv_1 _3892_ (.Y(_3092_),
    .A(\dtop.player_inst.synth.alu.acc[9] ));
 sg13g2_inv_1 _3893_ (.Y(_3093_),
    .A(\dtop.player_inst.synth.alu.acc[8] ));
 sg13g2_inv_1 _3894_ (.Y(_3094_),
    .A(net501));
 sg13g2_inv_1 _3895_ (.Y(_3095_),
    .A(net508));
 sg13g2_inv_1 _3896_ (.Y(_3096_),
    .A(net498));
 sg13g2_inv_1 _3897_ (.Y(_3097_),
    .A(net485));
 sg13g2_inv_1 _3898_ (.Y(_3098_),
    .A(net490));
 sg13g2_inv_1 _3899_ (.Y(_3099_),
    .A(net518));
 sg13g2_inv_1 _3900_ (.Y(_3100_),
    .A(net440));
 sg13g2_inv_1 _3901_ (.Y(_3101_),
    .A(net349));
 sg13g2_inv_1 _3902_ (.Y(_3102_),
    .A(net385));
 sg13g2_inv_1 _3903_ (.Y(_3103_),
    .A(net417));
 sg13g2_inv_1 _3904_ (.Y(_3104_),
    .A(net354));
 sg13g2_inv_1 _3905_ (.Y(_3105_),
    .A(net413));
 sg13g2_inv_1 _3906_ (.Y(_3106_),
    .A(net414));
 sg13g2_inv_1 _3907_ (.Y(_3107_),
    .A(net386));
 sg13g2_inv_1 _3908_ (.Y(_3108_),
    .A(net396));
 sg13g2_inv_1 _3909_ (.Y(_3109_),
    .A(net323));
 sg13g2_inv_1 _3910_ (.Y(_3110_),
    .A(net338));
 sg13g2_inv_1 _3911_ (.Y(_3111_),
    .A(net334));
 sg13g2_inv_1 _3912_ (.Y(_3112_),
    .A(net342));
 sg13g2_inv_1 _3913_ (.Y(_3113_),
    .A(net329));
 sg13g2_inv_1 _3914_ (.Y(_3114_),
    .A(net523));
 sg13g2_inv_1 _3915_ (.Y(_3115_),
    .A(net463));
 sg13g2_inv_1 _3916_ (.Y(_3116_),
    .A(net531));
 sg13g2_inv_1 _3917_ (.Y(_3117_),
    .A(net499));
 sg13g2_inv_1 _3918_ (.Y(_3118_),
    .A(net514));
 sg13g2_inv_1 _3919_ (.Y(_3119_),
    .A(net471));
 sg13g2_inv_2 _3920_ (.Y(_3120_),
    .A(net1447));
 sg13g2_inv_2 _3921_ (.Y(_3121_),
    .A(net662));
 sg13g2_inv_1 _3922_ (.Y(_3122_),
    .A(\dtop.vtop.pipeline.zg[7] ));
 sg13g2_inv_2 _3923_ (.Y(_3123_),
    .A(net655));
 sg13g2_inv_1 _3924_ (.Y(_3124_),
    .A(_0075_));
 sg13g2_inv_2 _3925_ (.Y(_3125_),
    .A(net1363));
 sg13g2_inv_2 _3926_ (.Y(_3126_),
    .A(\dtop.detune_counter[14] ));
 sg13g2_inv_1 _3927_ (.Y(_3127_),
    .A(net1397));
 sg13g2_inv_4 _3928_ (.A(net1399),
    .Y(_3128_));
 sg13g2_inv_1 _3929_ (.Y(_3129_),
    .A(net1402));
 sg13g2_inv_2 _3930_ (.Y(_3130_),
    .A(net1405));
 sg13g2_inv_2 _3931_ (.Y(_3131_),
    .A(\dtop.vtop.logo.addr[11] ));
 sg13g2_inv_2 _3932_ (.Y(_3132_),
    .A(\dtop.vtop.logo.addr[10] ));
 sg13g2_inv_2 _3933_ (.Y(_3133_),
    .A(net1415));
 sg13g2_inv_1 _3934_ (.Y(_3134_),
    .A(net1426));
 sg13g2_inv_1 _3935_ (.Y(_3135_),
    .A(\dtop.oct_counter[4] ));
 sg13g2_inv_4 _3936_ (.A(net1392),
    .Y(_3136_));
 sg13g2_inv_2 _3937_ (.Y(_3137_),
    .A(net1378));
 sg13g2_inv_2 _3938_ (.Y(_3138_),
    .A(net1382));
 sg13g2_inv_2 _3939_ (.Y(_3139_),
    .A(net1370));
 sg13g2_inv_2 _3940_ (.Y(_3140_),
    .A(net1376));
 sg13g2_inv_1 _3941_ (.Y(_3141_),
    .A(net1371));
 sg13g2_inv_1 _3942_ (.Y(_3142_),
    .A(net1368));
 sg13g2_inv_1 _3943_ (.Y(_3143_),
    .A(net1357));
 sg13g2_inv_2 _3944_ (.Y(_3144_),
    .A(net1429));
 sg13g2_inv_1 _3945_ (.Y(_3145_),
    .A(\dtop.detune_counter[17] ));
 sg13g2_inv_1 _3946_ (.Y(_3146_),
    .A(net1394));
 sg13g2_inv_1 _3947_ (.Y(_3147_),
    .A(\dtop.vtop.pipeline.wave_index[0] ));
 sg13g2_inv_1 _3948_ (.Y(_3148_),
    .A(net632));
 sg13g2_inv_2 _3949_ (.Y(_3149_),
    .A(\dtop.vtop.rs.x_scan.phase[1] ));
 sg13g2_inv_1 _3950_ (.Y(_3150_),
    .A(_0001_));
 sg13g2_inv_1 _3951_ (.Y(_3151_),
    .A(_0004_));
 sg13g2_inv_1 _3952_ (.Y(_3152_),
    .A(_0003_));
 sg13g2_inv_1 _3953_ (.Y(_3153_),
    .A(_0005_));
 sg13g2_inv_2 _3954_ (.Y(_3154_),
    .A(\dtop.vtop.pipeline.nstep[0] ));
 sg13g2_inv_1 _3955_ (.Y(_3155_),
    .A(net469));
 sg13g2_inv_1 _3956_ (.Y(_3156_),
    .A(net580));
 sg13g2_inv_1 _3957_ (.Y(_3157_),
    .A(_0010_));
 sg13g2_inv_1 _3958_ (.Y(_3158_),
    .A(_0014_));
 sg13g2_inv_1 _3959_ (.Y(_3159_),
    .A(_0020_));
 sg13g2_inv_1 _3960_ (.Y(_3160_),
    .A(_0027_));
 sg13g2_inv_1 _3961_ (.Y(_3161_),
    .A(net496));
 sg13g2_inv_1 _3962_ (.Y(_3162_),
    .A(\dtop.vtop.dphases[1][0] ));
 sg13g2_inv_1 _3963_ (.Y(_3163_),
    .A(net461));
 sg13g2_inv_1 _3964_ (.Y(_3164_),
    .A(\dtop.vtop.dphases[1][1] ));
 sg13g2_inv_1 _3965_ (.Y(_3165_),
    .A(net507));
 sg13g2_inv_1 _3966_ (.Y(_3166_),
    .A(\dtop.vtop.dphases[1][2] ));
 sg13g2_inv_1 _3967_ (.Y(_3167_),
    .A(net474));
 sg13g2_inv_1 _3968_ (.Y(_3168_),
    .A(net475));
 sg13g2_inv_1 _3969_ (.Y(_3169_),
    .A(\dtop.vtop.dphases[1][4] ));
 sg13g2_inv_1 _3970_ (.Y(_3170_),
    .A(\dtop.vtop.dphases[1][5] ));
 sg13g2_inv_1 _3971_ (.Y(_3171_),
    .A(\dtop.vtop.dphases[1][6] ));
 sg13g2_inv_1 _3972_ (.Y(_3172_),
    .A(\dtop.vtop.dphases[1][7] ));
 sg13g2_inv_1 _3973_ (.Y(_3173_),
    .A(net374));
 sg13g2_inv_1 _3974_ (.Y(_3174_),
    .A(\dtop.vtop.dphases[1][9] ));
 sg13g2_inv_1 _3975_ (.Y(_3175_),
    .A(net344));
 sg13g2_inv_1 _3976_ (.Y(_3176_),
    .A(_0058_));
 sg13g2_inv_1 _3977_ (.Y(_3177_),
    .A(_0074_));
 sg13g2_inv_1 _3978_ (.Y(_3178_),
    .A(net614));
 sg13g2_inv_1 _3979_ (.Y(_3179_),
    .A(net615));
 sg13g2_inv_1 _3980_ (.Y(_3180_),
    .A(uio_out[5]));
 sg13g2_inv_1 _3981_ (.Y(_3181_),
    .A(net563));
 sg13g2_inv_1 _3982_ (.Y(_3182_),
    .A(net581));
 sg13g2_inv_1 _3983_ (.Y(_3183_),
    .A(net638));
 sg13g2_and2_2 _3984_ (.A(net1384),
    .B(net1390),
    .X(_3184_));
 sg13g2_nand2_2 _3985_ (.Y(_3185_),
    .A(net1383),
    .B(net1391));
 sg13g2_nor2_2 _3986_ (.A(net1377),
    .B(net1381),
    .Y(_3186_));
 sg13g2_or2_1 _3987_ (.X(_3187_),
    .B(net1381),
    .A(net1377));
 sg13g2_nand2_1 _3988_ (.Y(_3188_),
    .A(_3184_),
    .B(_3186_));
 sg13g2_nand2b_2 _3989_ (.Y(_3189_),
    .B(net1371),
    .A_N(net1375));
 sg13g2_nor4_2 _3990_ (.A(net1367),
    .B(net1349),
    .C(net1347),
    .Y(_3190_),
    .D(net1346));
 sg13g2_nand2_2 _3991_ (.Y(_3191_),
    .A(net692),
    .B(_3190_));
 sg13g2_xor2_1 _3992_ (.B(_3191_),
    .A(net1445),
    .X(_3192_));
 sg13g2_nor2_1 _3993_ (.A(_3144_),
    .B(_3192_),
    .Y(_0100_));
 sg13g2_nor2_1 _3994_ (.A(net669),
    .B(_3191_),
    .Y(_3193_));
 sg13g2_o21ai_1 _3995_ (.B1(net1430),
    .Y(_3194_),
    .A1(net1444),
    .A2(net670));
 sg13g2_a21oi_1 _3996_ (.A1(net1444),
    .A2(net670),
    .Y(_0101_),
    .B1(_3194_));
 sg13g2_nor3_2 _3997_ (.A(_0085_),
    .B(_0084_),
    .C(_3191_),
    .Y(_3195_));
 sg13g2_o21ai_1 _3998_ (.B1(net1430),
    .Y(_3196_),
    .A1(net1442),
    .A2(_3195_));
 sg13g2_a21oi_1 _3999_ (.A1(net574),
    .A2(_3195_),
    .Y(_0102_),
    .B1(_3196_));
 sg13g2_nor2b_2 _4000_ (.A(net1395),
    .B_N(net1396),
    .Y(_3197_));
 sg13g2_and2_1 _4001_ (.A(net1394),
    .B(_3197_),
    .X(_3198_));
 sg13g2_nand2_1 _4002_ (.Y(_3199_),
    .A(net1394),
    .B(_3197_));
 sg13g2_nand2_1 _4003_ (.Y(_3200_),
    .A(net1396),
    .B(net1395));
 sg13g2_nor4_1 _4004_ (.A(net1397),
    .B(net1398),
    .C(_3146_),
    .D(_3200_),
    .Y(_3201_));
 sg13g2_o21ai_1 _4005_ (.B1(_3145_),
    .Y(_3202_),
    .A1(_3198_),
    .A2(_3201_));
 sg13g2_inv_1 _4006_ (.Y(_3203_),
    .A(_3202_));
 sg13g2_nand3b_1 _4007_ (.B(_3154_),
    .C(_3202_),
    .Y(_3204_),
    .A_N(net1352));
 sg13g2_nor2_1 _4008_ (.A(\dtop.vtop.force_sat0 ),
    .B(\dtop.ext_control[6] ),
    .Y(_3205_));
 sg13g2_nand3_1 _4009_ (.B(_3204_),
    .C(_3205_),
    .A(\dtop.vtop.logo_d[1] ),
    .Y(_3206_));
 sg13g2_nor2_2 _4010_ (.A(\dtop.vtop.rs.x_scan.phase[0] ),
    .B(\dtop.vtop.rs.x_scan.phase[1] ),
    .Y(_3207_));
 sg13g2_nor2_2 _4011_ (.A(\dtop.vtop.rs.scan_y.phase[1] ),
    .B(\dtop.vtop.rs.scan_y.phase[0] ),
    .Y(_3208_));
 sg13g2_nand3_1 _4012_ (.B(_3207_),
    .C(_3208_),
    .A(_3206_),
    .Y(_3209_));
 sg13g2_and2_2 _4013_ (.A(\dtop.detune_counter[17] ),
    .B(_3197_),
    .X(_3210_));
 sg13g2_nand3b_1 _4014_ (.B(\dtop.detune_counter[17] ),
    .C(net1396),
    .Y(_3211_),
    .A_N(net1395));
 sg13g2_nor2_1 _4015_ (.A(\dtop.detune_counter[14] ),
    .B(net1397),
    .Y(_3212_));
 sg13g2_nor2_2 _4016_ (.A(net1344),
    .B(_3212_),
    .Y(_3213_));
 sg13g2_nand2_1 _4017_ (.Y(_3214_),
    .A(net1443),
    .B(_0083_));
 sg13g2_a21oi_2 _4018_ (.B1(net1441),
    .Y(_3215_),
    .A2(_0083_),
    .A1(net1443));
 sg13g2_nor2_2 _4019_ (.A(net1445),
    .B(_3215_),
    .Y(_3216_));
 sg13g2_and2_1 _4020_ (.A(net1441),
    .B(net1376),
    .X(_3217_));
 sg13g2_xor2_1 _4021_ (.B(net1376),
    .A(net1441),
    .X(_3218_));
 sg13g2_o21ai_1 _4022_ (.B1(net1382),
    .Y(_3219_),
    .A1(net1445),
    .A2(_3215_));
 sg13g2_o21ai_1 _4023_ (.B1(net1443),
    .Y(_3220_),
    .A1(net1442),
    .A2(_0083_));
 sg13g2_xnor2_1 _4024_ (.Y(_3221_),
    .A(_0093_),
    .B(_3220_));
 sg13g2_nand2b_1 _4025_ (.Y(_3222_),
    .B(net1378),
    .A_N(_3220_));
 sg13g2_o21ai_1 _4026_ (.B1(_3222_),
    .Y(_3223_),
    .A1(_3219_),
    .A2(_3221_));
 sg13g2_a21oi_1 _4027_ (.A1(_3218_),
    .A2(_3223_),
    .Y(_3224_),
    .B1(_3217_));
 sg13g2_xnor2_1 _4028_ (.Y(_3225_),
    .A(_0092_),
    .B(_3216_));
 sg13g2_or2_1 _4029_ (.X(_3226_),
    .B(_3225_),
    .A(_3224_));
 sg13g2_o21ai_1 _4030_ (.B1(_3226_),
    .Y(_3227_),
    .A1(_0092_),
    .A2(_3216_));
 sg13g2_nor2_1 _4031_ (.A(net1444),
    .B(net1446),
    .Y(_3228_));
 sg13g2_xor2_1 _4032_ (.B(net1445),
    .A(net1443),
    .X(_3229_));
 sg13g2_nor2_1 _4033_ (.A(_3215_),
    .B(_3229_),
    .Y(_3230_));
 sg13g2_xnor2_1 _4034_ (.Y(_3231_),
    .A(\dtop.player_inst.program_addr[6] ),
    .B(_3230_));
 sg13g2_nor2_1 _4035_ (.A(net1368),
    .B(_3230_),
    .Y(_3232_));
 sg13g2_a21oi_2 _4036_ (.B1(_3232_),
    .Y(_3233_),
    .A2(_3231_),
    .A1(_3227_));
 sg13g2_a21oi_1 _4037_ (.A1(net1441),
    .A2(net1443),
    .Y(_3234_),
    .B1(net1445));
 sg13g2_a21oi_1 _4038_ (.A1(net1445),
    .A2(_3214_),
    .Y(_3235_),
    .B1(_3234_));
 sg13g2_or2_1 _4039_ (.X(_3236_),
    .B(_3235_),
    .A(_3215_));
 sg13g2_nor2b_1 _4040_ (.A(_3233_),
    .B_N(_3236_),
    .Y(_3237_));
 sg13g2_xor2_1 _4041_ (.B(_3236_),
    .A(_3233_),
    .X(_3238_));
 sg13g2_nor2_1 _4042_ (.A(_0095_),
    .B(_3238_),
    .Y(_3239_));
 sg13g2_xor2_1 _4043_ (.B(_3231_),
    .A(_3227_),
    .X(_3240_));
 sg13g2_xor2_1 _4044_ (.B(_3240_),
    .A(\dtop.vtop.pipeline.dz[6] ),
    .X(_3241_));
 sg13g2_xor2_1 _4045_ (.B(_3238_),
    .A(_0095_),
    .X(_3242_));
 sg13g2_nand2_1 _4046_ (.Y(_3243_),
    .A(_3241_),
    .B(_3242_));
 sg13g2_xor2_1 _4047_ (.B(_3225_),
    .A(_3224_),
    .X(_3244_));
 sg13g2_xor2_1 _4048_ (.B(_3244_),
    .A(\dtop.vtop.pipeline.dz[5] ),
    .X(_3245_));
 sg13g2_xor2_1 _4049_ (.B(_3223_),
    .A(_3218_),
    .X(_3246_));
 sg13g2_xor2_1 _4050_ (.B(_3246_),
    .A(\dtop.vtop.pipeline.dz[4] ),
    .X(_3247_));
 sg13g2_nand4_1 _4051_ (.B(_3242_),
    .C(_3245_),
    .A(_3241_),
    .Y(_3248_),
    .D(_3247_));
 sg13g2_xor2_1 _4052_ (.B(_3221_),
    .A(_3219_),
    .X(_3249_));
 sg13g2_xnor2_1 _4053_ (.Y(_3250_),
    .A(_3219_),
    .B(_3221_));
 sg13g2_nand2_1 _4054_ (.Y(_3251_),
    .A(_0098_),
    .B(_3250_));
 sg13g2_xnor2_1 _4055_ (.Y(_3252_),
    .A(net1382),
    .B(_3216_));
 sg13g2_xnor2_1 _4056_ (.Y(_3253_),
    .A(\dtop.vtop.pipeline.dz[2] ),
    .B(_3252_));
 sg13g2_xnor2_1 _4057_ (.Y(_3254_),
    .A(_0098_),
    .B(_3250_));
 sg13g2_nor2_1 _4058_ (.A(_3253_),
    .B(_3254_),
    .Y(_3255_));
 sg13g2_and2_1 _4059_ (.A(\dtop.vtop.pipeline.dz[1] ),
    .B(net1388),
    .X(_3256_));
 sg13g2_nand2b_1 _4060_ (.Y(_3257_),
    .B(_3252_),
    .A_N(_0099_));
 sg13g2_o21ai_1 _4061_ (.B1(_3257_),
    .Y(_3258_),
    .A1(_0098_),
    .A2(_3250_));
 sg13g2_xor2_1 _4062_ (.B(net1388),
    .A(\dtop.vtop.pipeline.dz[1] ),
    .X(_3259_));
 sg13g2_o21ai_1 _4063_ (.B1(_3259_),
    .Y(_3260_),
    .A1(\dtop.vtop.pipeline.dz[0] ),
    .A2(net1392));
 sg13g2_nor3_1 _4064_ (.A(_3253_),
    .B(_3254_),
    .C(_3260_),
    .Y(_3261_));
 sg13g2_a221oi_1 _4065_ (.B2(_3251_),
    .C1(_3261_),
    .B1(_3258_),
    .A1(_3255_),
    .Y(_3262_),
    .A2(_3256_));
 sg13g2_nand2b_1 _4066_ (.Y(_3263_),
    .B(_3244_),
    .A_N(_0097_));
 sg13g2_nand3_1 _4067_ (.B(_3245_),
    .C(_3246_),
    .A(\dtop.vtop.pipeline.dz[4] ),
    .Y(_3264_));
 sg13g2_a21oi_1 _4068_ (.A1(_3263_),
    .A2(_3264_),
    .Y(_3265_),
    .B1(_3243_));
 sg13g2_nand2b_1 _4069_ (.Y(_3266_),
    .B(_3240_),
    .A_N(_0096_));
 sg13g2_a21oi_1 _4070_ (.A1(_0095_),
    .A2(_3238_),
    .Y(_3267_),
    .B1(_3266_));
 sg13g2_nand3_1 _4071_ (.B(net1443),
    .C(net1445),
    .A(net1441),
    .Y(_3268_));
 sg13g2_o21ai_1 _4072_ (.B1(_3268_),
    .Y(_3269_),
    .A1(net1441),
    .A2(_3214_));
 sg13g2_xor2_1 _4073_ (.B(_3269_),
    .A(_3237_),
    .X(_3270_));
 sg13g2_nor2_1 _4074_ (.A(_0094_),
    .B(_3270_),
    .Y(_3271_));
 sg13g2_nor4_1 _4075_ (.A(_3239_),
    .B(_3265_),
    .C(_3267_),
    .D(_3271_),
    .Y(_3272_));
 sg13g2_o21ai_1 _4076_ (.B1(_3272_),
    .Y(_3273_),
    .A1(_3248_),
    .A2(_3262_));
 sg13g2_nand3_1 _4077_ (.B(_3237_),
    .C(_3268_),
    .A(net1441),
    .Y(_3274_));
 sg13g2_nand2_1 _4078_ (.Y(_3275_),
    .A(_3215_),
    .B(_3233_));
 sg13g2_and4_1 _4079_ (.A(_3207_),
    .B(_3268_),
    .C(_3274_),
    .D(_3275_),
    .X(_3276_));
 sg13g2_nand2_1 _4080_ (.Y(_3277_),
    .A(_0094_),
    .B(_3270_));
 sg13g2_nand3_1 _4081_ (.B(_3276_),
    .C(_3277_),
    .A(_3273_),
    .Y(_3278_));
 sg13g2_o21ai_1 _4082_ (.B1(_3255_),
    .Y(_3279_),
    .A1(_3073_),
    .A2(_3136_));
 sg13g2_nor4_1 _4083_ (.A(_3248_),
    .B(_3260_),
    .C(_3271_),
    .D(_3279_),
    .Y(_3280_));
 sg13g2_or2_1 _4084_ (.X(_3281_),
    .B(net1395),
    .A(\dtop.detune_counter[15] ));
 sg13g2_nor2_1 _4085_ (.A(\dtop.detune_counter[17] ),
    .B(_3281_),
    .Y(_3282_));
 sg13g2_nor2_1 _4086_ (.A(_3210_),
    .B(_3282_),
    .Y(_3283_));
 sg13g2_nor2b_1 _4087_ (.A(_3283_),
    .B_N(_3212_),
    .Y(_3284_));
 sg13g2_nand2_1 _4088_ (.Y(_3285_),
    .A(_0018_),
    .B(net1283));
 sg13g2_a21oi_1 _4089_ (.A1(_0018_),
    .A2(net1283),
    .Y(_3286_),
    .B1(\dtop.vtop.pipeline.neg_t[5] ));
 sg13g2_nand3_1 _4090_ (.B(_0021_),
    .C(net1283),
    .A(\dtop.vtop.pipeline.neg_t[3] ),
    .Y(_3287_));
 sg13g2_nand2_1 _4091_ (.Y(_3288_),
    .A(_0023_),
    .B(net1283));
 sg13g2_a21oi_1 _4092_ (.A1(_0023_),
    .A2(net1283),
    .Y(_3289_),
    .B1(\dtop.vtop.pipeline.neg_t[2] ));
 sg13g2_nand2_1 _4093_ (.Y(_3290_),
    .A(_0077_),
    .B(net1284));
 sg13g2_nand4_1 _4094_ (.B(_3124_),
    .C(_0025_),
    .A(\dtop.vtop.pipeline.neg_t[0] ),
    .Y(_3291_),
    .D(net1283));
 sg13g2_xor2_1 _4095_ (.B(_3290_),
    .A(_0024_),
    .X(_3292_));
 sg13g2_a22oi_1 _4096_ (.Y(_3293_),
    .B1(_3291_),
    .B2(_3292_),
    .A2(_3290_),
    .A1(_3075_));
 sg13g2_xnor2_1 _4097_ (.Y(_3294_),
    .A(_0022_),
    .B(_3288_));
 sg13g2_nor2_1 _4098_ (.A(_3293_),
    .B(_3294_),
    .Y(_3295_));
 sg13g2_o21ai_1 _4099_ (.B1(_3287_),
    .Y(_3296_),
    .A1(_3289_),
    .A2(_3295_));
 sg13g2_nand2_1 _4100_ (.Y(_3297_),
    .A(_0020_),
    .B(net1284));
 sg13g2_a21oi_1 _4101_ (.A1(_0021_),
    .A2(net1284),
    .Y(_3298_),
    .B1(\dtop.vtop.pipeline.neg_t[3] ));
 sg13g2_a21oi_1 _4102_ (.A1(_0019_),
    .A2(_3297_),
    .Y(_3299_),
    .B1(_3298_));
 sg13g2_xor2_1 _4103_ (.B(_3285_),
    .A(_0017_),
    .X(_3300_));
 sg13g2_o21ai_1 _4104_ (.B1(_3300_),
    .Y(_3301_),
    .A1(_0019_),
    .A2(_3297_));
 sg13g2_a21oi_1 _4105_ (.A1(_3296_),
    .A2(_3299_),
    .Y(_3302_),
    .B1(_3301_));
 sg13g2_nand2_1 _4106_ (.Y(_3303_),
    .A(_0016_),
    .B(net1284));
 sg13g2_xor2_1 _4107_ (.B(_3303_),
    .A(_0015_),
    .X(_3304_));
 sg13g2_o21ai_1 _4108_ (.B1(_3304_),
    .Y(_3305_),
    .A1(_3286_),
    .A2(_3302_));
 sg13g2_a21oi_1 _4109_ (.A1(_0000_),
    .A2(net1283),
    .Y(_3306_),
    .B1(\dtop.vtop.pipeline.neg_t[7] ));
 sg13g2_a21oi_1 _4110_ (.A1(_3074_),
    .A2(_3303_),
    .Y(_3307_),
    .B1(_3306_));
 sg13g2_nand2_1 _4111_ (.Y(_3308_),
    .A(_3305_),
    .B(_3307_));
 sg13g2_nand3_1 _4112_ (.B(_0000_),
    .C(net1283),
    .A(\dtop.vtop.pipeline.neg_t[7] ),
    .Y(_3309_));
 sg13g2_nand2_1 _4113_ (.Y(_3310_),
    .A(_0014_),
    .B(net1284));
 sg13g2_o21ai_1 _4114_ (.B1(\dtop.vtop.pipeline.neg_t[9] ),
    .Y(_3311_),
    .A1(_0013_),
    .A2(_3310_));
 sg13g2_nor2b_1 _4115_ (.A(_3311_),
    .B_N(_3309_),
    .Y(_3312_));
 sg13g2_a221oi_1 _4116_ (.B2(_3308_),
    .C1(_0026_),
    .B1(_3312_),
    .A1(_0013_),
    .Y(_3313_),
    .A2(_3310_));
 sg13g2_xnor2_1 _4117_ (.Y(_3314_),
    .A(net1344),
    .B(_3313_));
 sg13g2_nor2_1 _4118_ (.A(_0091_),
    .B(_3314_),
    .Y(_3315_));
 sg13g2_o21ai_1 _4119_ (.B1(_3315_),
    .Y(_3316_),
    .A1(_3278_),
    .A2(_3280_));
 sg13g2_and2_1 _4120_ (.A(_3202_),
    .B(_3276_),
    .X(_3317_));
 sg13g2_a21oi_1 _4121_ (.A1(_3316_),
    .A2(_3317_),
    .Y(_3318_),
    .B1(_3213_));
 sg13g2_o21ai_1 _4122_ (.B1(_3318_),
    .Y(_3319_),
    .A1(_3203_),
    .A2(_3276_));
 sg13g2_nand3b_1 _4123_ (.B(net1395),
    .C(net1396),
    .Y(_3320_),
    .A_N(\dtop.detune_counter[17] ));
 sg13g2_and2_2 _4124_ (.A(net1398),
    .B(net1400),
    .X(_3321_));
 sg13g2_nand2_2 _4125_ (.Y(_3322_),
    .A(net1398),
    .B(net1399));
 sg13g2_nand2_1 _4126_ (.Y(_3323_),
    .A(\dtop.detune_counter[14] ),
    .B(net1397));
 sg13g2_nor2_1 _4127_ (.A(_3322_),
    .B(_3323_),
    .Y(_3324_));
 sg13g2_nor3_2 _4128_ (.A(_3126_),
    .B(net1401),
    .C(net1328),
    .Y(_3325_));
 sg13g2_nor2_2 _4129_ (.A(_3320_),
    .B(_3325_),
    .Y(_3326_));
 sg13g2_or2_2 _4130_ (.X(_3327_),
    .B(_3325_),
    .A(_3320_));
 sg13g2_and2_2 _4131_ (.A(\dtop.vtop.force_sat0 ),
    .B(_3204_),
    .X(_3328_));
 sg13g2_nor2_1 _4132_ (.A(net1282),
    .B(_3328_),
    .Y(_3329_));
 sg13g2_a21o_2 _4133_ (.A2(_3329_),
    .A1(_3319_),
    .B1(_3209_),
    .X(_3330_));
 sg13g2_inv_2 _4134_ (.Y(_3331_),
    .A(_3330_));
 sg13g2_nor2_2 _4135_ (.A(_3120_),
    .B(_3330_),
    .Y(_3332_));
 sg13g2_nand2_1 _4136_ (.Y(_3333_),
    .A(net1447),
    .B(net1358));
 sg13g2_nand2_1 _4137_ (.Y(_3334_),
    .A(net1357),
    .B(_3332_));
 sg13g2_nand2_1 _4138_ (.Y(_3335_),
    .A(_3099_),
    .B(net1385));
 sg13g2_nor2_1 _4139_ (.A(_3100_),
    .B(net1390),
    .Y(_3336_));
 sg13g2_nor2_1 _4140_ (.A(_3099_),
    .B(net1384),
    .Y(_3337_));
 sg13g2_a221oi_1 _4141_ (.B2(_3336_),
    .C1(_3337_),
    .B1(_3335_),
    .A1(\dtop.out_sample[2] ),
    .Y(_3338_),
    .A2(_3138_));
 sg13g2_a221oi_1 _4142_ (.B2(_3098_),
    .C1(_3338_),
    .B1(net1380),
    .A1(_3097_),
    .Y(_3339_),
    .A2(net1377));
 sg13g2_a221oi_1 _4143_ (.B2(\dtop.out_sample[4] ),
    .C1(_3339_),
    .B1(_3140_),
    .A1(\dtop.out_sample[3] ),
    .Y(_3340_),
    .A2(_3137_));
 sg13g2_a221oi_1 _4144_ (.B2(_3095_),
    .C1(_3340_),
    .B1(net1371),
    .A1(_3096_),
    .Y(_3341_),
    .A2(net1374));
 sg13g2_a221oi_1 _4145_ (.B2(\dtop.out_sample[5] ),
    .C1(_3341_),
    .B1(_3141_),
    .A1(\dtop.out_sample[6] ),
    .Y(_3342_),
    .A2(_3139_));
 sg13g2_a21oi_1 _4146_ (.A1(_3094_),
    .A2(net1370),
    .Y(_3343_),
    .B1(_3342_));
 sg13g2_xnor2_1 _4147_ (.Y(_3344_),
    .A(net1445),
    .B(_3343_));
 sg13g2_and2_1 _4148_ (.A(_3326_),
    .B(_3344_),
    .X(_3345_));
 sg13g2_nand2_1 _4149_ (.Y(_3346_),
    .A(_0084_),
    .B(_3345_));
 sg13g2_xor2_1 _4150_ (.B(net1383),
    .A(\dtop.oct_counter[3] ),
    .X(_3347_));
 sg13g2_nand2_2 _4151_ (.Y(_3348_),
    .A(_0006_),
    .B(_3347_));
 sg13g2_nand2_1 _4152_ (.Y(_3349_),
    .A(net1392),
    .B(net1448));
 sg13g2_nor2_1 _4153_ (.A(_0012_),
    .B(_3349_),
    .Y(_3350_));
 sg13g2_nand2_1 _4154_ (.Y(_3351_),
    .A(\dtop.vtop.color[7] ),
    .B(_3350_));
 sg13g2_nand2_2 _4155_ (.Y(_3352_),
    .A(net1448),
    .B(_3347_));
 sg13g2_nand2_1 _4156_ (.Y(_0397_),
    .A(_3351_),
    .B(_3352_));
 sg13g2_o21ai_1 _4157_ (.B1(_0397_),
    .Y(_0398_),
    .A1(\dtop.vtop.color[7] ),
    .A2(_3350_));
 sg13g2_nor2_2 _4158_ (.A(_3136_),
    .B(net1448),
    .Y(_0399_));
 sg13g2_inv_1 _4159_ (.Y(_0400_),
    .A(_0399_));
 sg13g2_xnor2_1 _4160_ (.Y(_0401_),
    .A(_0010_),
    .B(_0399_));
 sg13g2_nand2b_1 _4161_ (.Y(_0402_),
    .B(_0401_),
    .A_N(_0398_));
 sg13g2_nand2_1 _4162_ (.Y(_0403_),
    .A(\dtop.vtop.color[8] ),
    .B(_0399_));
 sg13g2_xnor2_1 _4163_ (.Y(_0404_),
    .A(_3156_),
    .B(_3348_));
 sg13g2_a21o_1 _4164_ (.A2(_0403_),
    .A1(_0402_),
    .B1(_0404_),
    .X(_0405_));
 sg13g2_o21ai_1 _4165_ (.B1(_0405_),
    .Y(_0406_),
    .A1(_3156_),
    .A2(_3348_));
 sg13g2_nand2_1 _4166_ (.Y(_0407_),
    .A(\dtop.vtop.color[10] ),
    .B(_0406_));
 sg13g2_inv_1 _4167_ (.Y(_0408_),
    .A(_0407_));
 sg13g2_nand3_1 _4168_ (.B(_3327_),
    .C(_0408_),
    .A(\dtop.vtop.color[11] ),
    .Y(_0409_));
 sg13g2_nand2b_1 _4169_ (.Y(_0410_),
    .B(_0409_),
    .A_N(_3328_));
 sg13g2_xnor2_1 _4170_ (.Y(_0411_),
    .A(_0009_),
    .B(_0406_));
 sg13g2_a21oi_1 _4171_ (.A1(_3327_),
    .A2(_0411_),
    .Y(_0412_),
    .B1(_0410_));
 sg13g2_nand2_1 _4172_ (.Y(_0413_),
    .A(_3346_),
    .B(_0412_));
 sg13g2_nand3_1 _4173_ (.B(_3332_),
    .C(_0413_),
    .A(net1357),
    .Y(_0414_));
 sg13g2_nand2_1 _4174_ (.Y(_0415_),
    .A(net1448),
    .B(_0410_));
 sg13g2_nand2_1 _4175_ (.Y(_0416_),
    .A(net1448),
    .B(_3327_));
 sg13g2_xnor2_1 _4176_ (.Y(_0417_),
    .A(_0398_),
    .B(_0401_));
 sg13g2_nand2b_1 _4177_ (.Y(_0418_),
    .B(_0417_),
    .A_N(_0416_));
 sg13g2_a21oi_1 _4178_ (.A1(_0415_),
    .A2(_0418_),
    .Y(_0419_),
    .B1(_3334_));
 sg13g2_a21oi_1 _4179_ (.A1(_3143_),
    .A2(uio_out[0]),
    .Y(_0420_),
    .B1(_0419_));
 sg13g2_o21ai_1 _4180_ (.B1(_0420_),
    .Y(_0103_),
    .A1(net469),
    .A2(_0414_));
 sg13g2_nor2_2 _4181_ (.A(_3328_),
    .B(_3345_),
    .Y(_0421_));
 sg13g2_nor2_1 _4182_ (.A(_0083_),
    .B(_3328_),
    .Y(_0422_));
 sg13g2_o21ai_1 _4183_ (.B1(_3327_),
    .Y(_0423_),
    .A1(\dtop.vtop.color[11] ),
    .A2(_0408_));
 sg13g2_o21ai_1 _4184_ (.B1(_0423_),
    .Y(_0424_),
    .A1(_0421_),
    .A2(_0422_));
 sg13g2_nand3_1 _4185_ (.B(_3332_),
    .C(_0424_),
    .A(net1357),
    .Y(_0425_));
 sg13g2_nand2b_1 _4186_ (.Y(_0426_),
    .B(net602),
    .A_N(net1357));
 sg13g2_nand3_1 _4187_ (.B(_0403_),
    .C(_0404_),
    .A(_0402_),
    .Y(_0427_));
 sg13g2_nand2_1 _4188_ (.Y(_0428_),
    .A(_0405_),
    .B(_0427_));
 sg13g2_o21ai_1 _4189_ (.B1(_0415_),
    .Y(_0429_),
    .A1(_0416_),
    .A2(_0428_));
 sg13g2_a21oi_1 _4190_ (.A1(_3155_),
    .A2(_0424_),
    .Y(_0430_),
    .B1(_0429_));
 sg13g2_o21ai_1 _4191_ (.B1(_0426_),
    .Y(_0104_),
    .A1(_3334_),
    .A2(_0430_));
 sg13g2_o21ai_1 _4192_ (.B1(_0414_),
    .Y(_0105_),
    .A1(net1358),
    .A2(_3178_));
 sg13g2_o21ai_1 _4193_ (.B1(_0425_),
    .Y(_0106_),
    .A1(net1358),
    .A2(_3179_));
 sg13g2_nand2b_1 _4194_ (.Y(_0431_),
    .B(net564),
    .A_N(net1360));
 sg13g2_nor2_2 _4195_ (.A(\dtop.vtop.rs.x_scan.phase[0] ),
    .B(_3149_),
    .Y(_0432_));
 sg13g2_o21ai_1 _4196_ (.B1(_0431_),
    .Y(_0107_),
    .A1(_3333_),
    .A2(_0432_));
 sg13g2_nand3_1 _4197_ (.B(net1447),
    .C(net1358),
    .A(net524),
    .Y(_0433_));
 sg13g2_o21ai_1 _4198_ (.B1(net525),
    .Y(_0108_),
    .A1(net1358),
    .A2(_3180_));
 sg13g2_or2_1 _4199_ (.X(_0434_),
    .B(_3323_),
    .A(_3199_));
 sg13g2_nor2b_1 _4200_ (.A(net1396),
    .B_N(net1395),
    .Y(_0435_));
 sg13g2_and2_2 _4201_ (.A(net1394),
    .B(_0435_),
    .X(_0436_));
 sg13g2_nand2_2 _4202_ (.Y(_0437_),
    .A(net1394),
    .B(_0435_));
 sg13g2_nor2_1 _4203_ (.A(net1397),
    .B(_3320_),
    .Y(_0438_));
 sg13g2_a22oi_1 _4204_ (.Y(_0439_),
    .B1(_0438_),
    .B2(net1398),
    .A2(_0436_),
    .A1(_3126_));
 sg13g2_a21o_2 _4205_ (.A2(_0439_),
    .A1(_0434_),
    .B1(_3146_),
    .X(_0440_));
 sg13g2_nor2_1 _4206_ (.A(_3209_),
    .B(_0440_),
    .Y(_0441_));
 sg13g2_a21oi_2 _4207_ (.B1(_3331_),
    .Y(_0442_),
    .A2(_0441_),
    .A1(_3318_));
 sg13g2_nor2_2 _4208_ (.A(net1356),
    .B(\dtop.vtop.pipeline.zg[8] ),
    .Y(_0443_));
 sg13g2_nor2_2 _4209_ (.A(net1355),
    .B(\dtop.vtop.pipeline.zg[7] ),
    .Y(_0444_));
 sg13g2_nor2_1 _4210_ (.A(_0009_),
    .B(_0444_),
    .Y(_0445_));
 sg13g2_or2_1 _4211_ (.X(_0446_),
    .B(\dtop.vtop.pipeline.zg[4] ),
    .A(net1356));
 sg13g2_nor2b_1 _4212_ (.A(_0011_),
    .B_N(_0446_),
    .Y(_0447_));
 sg13g2_nor2_1 _4213_ (.A(net1355),
    .B(\dtop.vtop.pipeline.zg[3] ),
    .Y(_0448_));
 sg13g2_xnor2_1 _4214_ (.Y(_0449_),
    .A(\dtop.vtop.color[7] ),
    .B(_0446_));
 sg13g2_a21oi_1 _4215_ (.A1(_0012_),
    .A2(_0448_),
    .Y(_0450_),
    .B1(_0449_));
 sg13g2_or2_1 _4216_ (.X(_0451_),
    .B(\dtop.vtop.pipeline.zg[5] ),
    .A(net1355));
 sg13g2_xor2_1 _4217_ (.B(_0451_),
    .A(\dtop.vtop.color[8] ),
    .X(_0452_));
 sg13g2_o21ai_1 _4218_ (.B1(_0452_),
    .Y(_0453_),
    .A1(_0447_),
    .A2(_0450_));
 sg13g2_nor2_2 _4219_ (.A(net1355),
    .B(\dtop.vtop.pipeline.zg[6] ),
    .Y(_0454_));
 sg13g2_nor2_1 _4220_ (.A(_0007_),
    .B(_0454_),
    .Y(_0455_));
 sg13g2_a21oi_1 _4221_ (.A1(_3157_),
    .A2(_0451_),
    .Y(_0456_),
    .B1(_0455_));
 sg13g2_xor2_1 _4222_ (.B(_0444_),
    .A(\dtop.vtop.color[10] ),
    .X(_0457_));
 sg13g2_a221oi_1 _4223_ (.B2(_0453_),
    .C1(_0457_),
    .B1(_0456_),
    .A1(_0007_),
    .Y(_0458_),
    .A2(_0454_));
 sg13g2_xor2_1 _4224_ (.B(_0448_),
    .A(\dtop.vtop.color[6] ),
    .X(_0459_));
 sg13g2_xnor2_1 _4225_ (.Y(_0460_),
    .A(_0007_),
    .B(_0454_));
 sg13g2_nor4_1 _4226_ (.A(_0449_),
    .B(_0457_),
    .C(_0459_),
    .D(_0460_),
    .Y(_0461_));
 sg13g2_a22oi_1 _4227_ (.Y(_0462_),
    .B1(_0452_),
    .B2(_0461_),
    .A2(_0443_),
    .A1(_0008_));
 sg13g2_o21ai_1 _4228_ (.B1(_0462_),
    .Y(_0463_),
    .A1(_0445_),
    .A2(_0458_));
 sg13g2_o21ai_1 _4229_ (.B1(_0463_),
    .Y(_0464_),
    .A1(_0008_),
    .A2(_0443_));
 sg13g2_nor2_1 _4230_ (.A(_0007_),
    .B(_0464_),
    .Y(_0465_));
 sg13g2_a21oi_1 _4231_ (.A1(_0454_),
    .A2(_0464_),
    .Y(_0466_),
    .B1(_0465_));
 sg13g2_nor2_1 _4232_ (.A(_3348_),
    .B(_0466_),
    .Y(_0467_));
 sg13g2_mux2_1 _4233_ (.A0(_0010_),
    .A1(_0451_),
    .S(_0464_),
    .X(_0468_));
 sg13g2_xnor2_1 _4234_ (.Y(_0469_),
    .A(_0399_),
    .B(_0468_));
 sg13g2_mux2_1 _4235_ (.A0(_0011_),
    .A1(_0446_),
    .S(_0464_),
    .X(_0470_));
 sg13g2_nand2_1 _4236_ (.Y(_0471_),
    .A(_3352_),
    .B(_0470_));
 sg13g2_mux2_1 _4237_ (.A0(\dtop.vtop.color[6] ),
    .A1(_0448_),
    .S(_0464_),
    .X(_0472_));
 sg13g2_nand2b_1 _4238_ (.Y(_0473_),
    .B(_0472_),
    .A_N(_3349_));
 sg13g2_o21ai_1 _4239_ (.B1(_0473_),
    .Y(_0474_),
    .A1(_3352_),
    .A2(_0470_));
 sg13g2_nand3_1 _4240_ (.B(_0471_),
    .C(_0474_),
    .A(_0469_),
    .Y(_0475_));
 sg13g2_o21ai_1 _4241_ (.B1(_0475_),
    .Y(_0476_),
    .A1(_0400_),
    .A2(_0468_));
 sg13g2_xnor2_1 _4242_ (.Y(_0477_),
    .A(_3348_),
    .B(_0466_));
 sg13g2_nor2b_1 _4243_ (.A(_0477_),
    .B_N(_0476_),
    .Y(_0478_));
 sg13g2_nor2_1 _4244_ (.A(_0467_),
    .B(_0478_),
    .Y(_0479_));
 sg13g2_nor2_1 _4245_ (.A(_0009_),
    .B(_0464_),
    .Y(_0480_));
 sg13g2_a21oi_1 _4246_ (.A1(_0444_),
    .A2(_0464_),
    .Y(_0481_),
    .B1(_0480_));
 sg13g2_or2_1 _4247_ (.X(_0482_),
    .B(_0481_),
    .A(_0479_));
 sg13g2_a21oi_1 _4248_ (.A1(_0479_),
    .A2(_0481_),
    .Y(_0483_),
    .B1(net1282));
 sg13g2_nand3_1 _4249_ (.B(_0482_),
    .C(_0483_),
    .A(_3155_),
    .Y(_0484_));
 sg13g2_and2_1 _4250_ (.A(_3327_),
    .B(_0443_),
    .X(_0485_));
 sg13g2_nand2b_1 _4251_ (.Y(_0486_),
    .B(_0485_),
    .A_N(_0008_));
 sg13g2_o21ai_1 _4252_ (.B1(_0421_),
    .Y(_0487_),
    .A1(_0482_),
    .A2(_0486_));
 sg13g2_a21oi_1 _4253_ (.A1(_0471_),
    .A2(_0474_),
    .Y(_0488_),
    .B1(_0469_));
 sg13g2_nand2b_1 _4254_ (.Y(_0489_),
    .B(_0475_),
    .A_N(_0416_));
 sg13g2_o21ai_1 _4255_ (.B1(net1447),
    .Y(_0490_),
    .A1(_0488_),
    .A2(_0489_));
 sg13g2_nor2_1 _4256_ (.A(_0487_),
    .B(_0490_),
    .Y(_0491_));
 sg13g2_and2_1 _4257_ (.A(_0484_),
    .B(_0491_),
    .X(_0492_));
 sg13g2_and2_1 _4258_ (.A(_0421_),
    .B(_0486_),
    .X(_0493_));
 sg13g2_o21ai_1 _4259_ (.B1(_0493_),
    .Y(_0494_),
    .A1(net1282),
    .A2(_0482_));
 sg13g2_nor2_1 _4260_ (.A(net1447),
    .B(_0494_),
    .Y(_0495_));
 sg13g2_nor3_1 _4261_ (.A(_0442_),
    .B(_0492_),
    .C(_0495_),
    .Y(_0496_));
 sg13g2_mux2_1 _4262_ (.A0(net635),
    .A1(_0496_),
    .S(net1361),
    .X(_0109_));
 sg13g2_nor2_1 _4263_ (.A(net1361),
    .B(net606),
    .Y(_0497_));
 sg13g2_nor2b_1 _4264_ (.A(_0476_),
    .B_N(_0477_),
    .Y(_0498_));
 sg13g2_nor3_1 _4265_ (.A(net1282),
    .B(_0478_),
    .C(_0498_),
    .Y(_0499_));
 sg13g2_nor3_1 _4266_ (.A(_3155_),
    .B(_0487_),
    .C(_0499_),
    .Y(_0500_));
 sg13g2_nor2_1 _4267_ (.A(net1448),
    .B(_0494_),
    .Y(_0501_));
 sg13g2_nor4_1 _4268_ (.A(_3120_),
    .B(_0442_),
    .C(_0500_),
    .D(_0501_),
    .Y(_0502_));
 sg13g2_nor2_1 _4269_ (.A(net1447),
    .B(_3330_),
    .Y(_0503_));
 sg13g2_a21oi_1 _4270_ (.A1(_0424_),
    .A2(_0503_),
    .Y(_0504_),
    .B1(_0502_));
 sg13g2_a21oi_1 _4271_ (.A1(net1362),
    .A2(_0504_),
    .Y(_0110_),
    .B1(_0497_));
 sg13g2_nand2b_1 _4272_ (.Y(_0505_),
    .B(net591),
    .A_N(net1358));
 sg13g2_a21oi_1 _4273_ (.A1(_0482_),
    .A2(_0483_),
    .Y(_0506_),
    .B1(_0487_));
 sg13g2_nor2_1 _4274_ (.A(_0442_),
    .B(_0506_),
    .Y(_0507_));
 sg13g2_nand2_1 _4275_ (.Y(_0508_),
    .A(_3123_),
    .B(_0399_));
 sg13g2_xnor2_1 _4276_ (.Y(_0509_),
    .A(\dtop.vtop.pipeline.zg[6] ),
    .B(_0399_));
 sg13g2_nor2_1 _4277_ (.A(\dtop.vtop.pipeline.zg[4] ),
    .B(_3349_),
    .Y(_0510_));
 sg13g2_or2_1 _4278_ (.X(_0511_),
    .B(_0510_),
    .A(_0028_));
 sg13g2_nand2_1 _4279_ (.Y(_0512_),
    .A(_0028_),
    .B(_0510_));
 sg13g2_nand2_1 _4280_ (.Y(_0513_),
    .A(_3352_),
    .B(_0512_));
 sg13g2_nand3_1 _4281_ (.B(_0511_),
    .C(_0513_),
    .A(_0509_),
    .Y(_0514_));
 sg13g2_xnor2_1 _4282_ (.Y(_0515_),
    .A(_3160_),
    .B(_3348_));
 sg13g2_a21o_1 _4283_ (.A2(_0514_),
    .A1(_0508_),
    .B1(_0515_),
    .X(_0516_));
 sg13g2_o21ai_1 _4284_ (.B1(_0516_),
    .Y(_0517_),
    .A1(_3160_),
    .A2(_3348_));
 sg13g2_nand2_1 _4285_ (.Y(_0518_),
    .A(_3121_),
    .B(_0517_));
 sg13g2_a21o_1 _4286_ (.A2(_0518_),
    .A1(net1355),
    .B1(net1282),
    .X(_0519_));
 sg13g2_o21ai_1 _4287_ (.B1(_0519_),
    .Y(_0520_),
    .A1(_0421_),
    .A2(_0422_));
 sg13g2_nand2_2 _4288_ (.Y(_0521_),
    .A(_3331_),
    .B(_0520_));
 sg13g2_a21oi_1 _4289_ (.A1(_3331_),
    .A2(_0520_),
    .Y(_0522_),
    .B1(net1447));
 sg13g2_o21ai_1 _4290_ (.B1(net1357),
    .Y(_0523_),
    .A1(_3120_),
    .A2(_0507_));
 sg13g2_o21ai_1 _4291_ (.B1(_0505_),
    .Y(_0111_),
    .A1(_0522_),
    .A2(_0523_));
 sg13g2_nand3b_1 _4292_ (.B(_0494_),
    .C(net1447),
    .Y(_0524_),
    .A_N(_0442_));
 sg13g2_nand2_1 _4293_ (.Y(_0525_),
    .A(net524),
    .B(_3120_));
 sg13g2_nand3_1 _4294_ (.B(_0524_),
    .C(_0525_),
    .A(net1358),
    .Y(_0526_));
 sg13g2_o21ai_1 _4295_ (.B1(_0526_),
    .Y(_0527_),
    .A1(net1361),
    .A2(net654));
 sg13g2_inv_1 _4296_ (.Y(_0112_),
    .A(_0527_));
 sg13g2_nor2_1 _4297_ (.A(net1361),
    .B(net609),
    .Y(_0528_));
 sg13g2_a21oi_1 _4298_ (.A1(_3121_),
    .A2(_0517_),
    .Y(_0529_),
    .B1(net1282));
 sg13g2_o21ai_1 _4299_ (.B1(_0529_),
    .Y(_0530_),
    .A1(_3121_),
    .A2(_0517_));
 sg13g2_a21oi_1 _4300_ (.A1(_0485_),
    .A2(_0517_),
    .Y(_0531_),
    .B1(_3328_));
 sg13g2_nand3_1 _4301_ (.B(_0530_),
    .C(_0531_),
    .A(_3346_),
    .Y(_0532_));
 sg13g2_nand2b_1 _4302_ (.Y(_0533_),
    .B(_3155_),
    .A_N(_0532_));
 sg13g2_and2_1 _4303_ (.A(net1448),
    .B(_0531_),
    .X(_0534_));
 sg13g2_a21oi_1 _4304_ (.A1(_0511_),
    .A2(_0513_),
    .Y(_0535_),
    .B1(_0509_));
 sg13g2_nand2_1 _4305_ (.Y(_0536_),
    .A(_3327_),
    .B(_0514_));
 sg13g2_o21ai_1 _4306_ (.B1(_0534_),
    .Y(_0537_),
    .A1(_0535_),
    .A2(_0536_));
 sg13g2_nand3_1 _4307_ (.B(_0533_),
    .C(_0537_),
    .A(_3332_),
    .Y(_0538_));
 sg13g2_nand2_1 _4308_ (.Y(_0539_),
    .A(net1357),
    .B(_0538_));
 sg13g2_a21oi_1 _4309_ (.A1(_3120_),
    .A2(_0507_),
    .Y(_0540_),
    .B1(_0539_));
 sg13g2_nor2_1 _4310_ (.A(_0528_),
    .B(_0540_),
    .Y(_0113_));
 sg13g2_nand3_1 _4311_ (.B(_0514_),
    .C(_0515_),
    .A(_0508_),
    .Y(_0541_));
 sg13g2_nand3_1 _4312_ (.B(_0516_),
    .C(_0541_),
    .A(_3327_),
    .Y(_0542_));
 sg13g2_nand2_1 _4313_ (.Y(_0543_),
    .A(_0534_),
    .B(_0542_));
 sg13g2_and2_1 _4314_ (.A(_3332_),
    .B(_0543_),
    .X(_0544_));
 sg13g2_o21ai_1 _4315_ (.B1(_0544_),
    .Y(_0545_),
    .A1(net1448),
    .A2(_0520_));
 sg13g2_nand2_1 _4316_ (.Y(_0546_),
    .A(_0413_),
    .B(_0503_));
 sg13g2_nand3_1 _4317_ (.B(_0545_),
    .C(_0546_),
    .A(net1359),
    .Y(_0547_));
 sg13g2_o21ai_1 _4318_ (.B1(_0547_),
    .Y(_0548_),
    .A1(net1360),
    .A2(net648));
 sg13g2_inv_1 _4319_ (.Y(_0114_),
    .A(_0548_));
 sg13g2_nand3_1 _4320_ (.B(_3331_),
    .C(_0532_),
    .A(net1357),
    .Y(_0549_));
 sg13g2_o21ai_1 _4321_ (.B1(_0549_),
    .Y(_0115_),
    .A1(net1360),
    .A2(_3181_));
 sg13g2_nor3_1 _4322_ (.A(\dtop.ext_control[5] ),
    .B(\dtop.vtop.rs.x_scan.phase[0] ),
    .C(_3149_),
    .Y(_0550_));
 sg13g2_a21oi_1 _4323_ (.A1(\dtop.ext_control[5] ),
    .A2(_0521_),
    .Y(_0551_),
    .B1(_0550_));
 sg13g2_mux2_1 _4324_ (.A0(net535),
    .A1(_0551_),
    .S(net1361),
    .X(_0116_));
 sg13g2_nand3_1 _4325_ (.B(_0079_),
    .C(_3344_),
    .A(net1362),
    .Y(_0552_));
 sg13g2_o21ai_1 _4326_ (.B1(_0552_),
    .Y(_0553_),
    .A1(net1359),
    .A2(net657));
 sg13g2_inv_1 _4327_ (.Y(_0117_),
    .A(net658));
 sg13g2_o21ai_1 _4328_ (.B1(_0552_),
    .Y(_0118_),
    .A1(net1359),
    .A2(_3182_));
 sg13g2_nor2b_1 _4329_ (.A(_0083_),
    .B_N(_3195_),
    .Y(_0554_));
 sg13g2_nand2b_1 _4330_ (.Y(_0555_),
    .B(_3195_),
    .A_N(_0083_));
 sg13g2_nand2_1 _4331_ (.Y(_0556_),
    .A(net1426),
    .B(net1393));
 sg13g2_nor2_2 _4332_ (.A(net1417),
    .B(net1423),
    .Y(_0557_));
 sg13g2_nor3_1 _4333_ (.A(\dtop.vtop.logo.addr[11] ),
    .B(\dtop.vtop.logo.addr[10] ),
    .C(net1415),
    .Y(_0558_));
 sg13g2_nand3_1 _4334_ (.B(_0557_),
    .C(_0558_),
    .A(\dtop.oct_counter[6] ),
    .Y(_0559_));
 sg13g2_nor4_1 _4335_ (.A(\dtop.oct_counter[4] ),
    .B(\dtop.oct_counter[3] ),
    .C(_0556_),
    .D(_0559_),
    .Y(_0560_));
 sg13g2_a21o_2 _4336_ (.A2(_0560_),
    .A1(_0554_),
    .B1(_0087_),
    .X(_0561_));
 sg13g2_xnor2_1 _4337_ (.Y(_0562_),
    .A(net695),
    .B(_0554_));
 sg13g2_nor2_1 _4338_ (.A(net1242),
    .B(net696),
    .Y(_0119_));
 sg13g2_nor2_1 _4339_ (.A(_0082_),
    .B(_0555_),
    .Y(_0563_));
 sg13g2_xnor2_1 _4340_ (.Y(_0564_),
    .A(net675),
    .B(_0563_));
 sg13g2_nor2_1 _4341_ (.A(net1242),
    .B(net676),
    .Y(_0120_));
 sg13g2_nor3_1 _4342_ (.A(_0082_),
    .B(_0081_),
    .C(_0555_),
    .Y(_0565_));
 sg13g2_nor2_1 _4343_ (.A(net1426),
    .B(_0565_),
    .Y(_0566_));
 sg13g2_and2_1 _4344_ (.A(net1426),
    .B(_0565_),
    .X(_0567_));
 sg13g2_nor3_1 _4345_ (.A(net1242),
    .B(net704),
    .C(_0567_),
    .Y(_0121_));
 sg13g2_nor2b_1 _4346_ (.A(_0046_),
    .B_N(_0565_),
    .Y(_0568_));
 sg13g2_xnor2_1 _4347_ (.Y(_0569_),
    .A(net596),
    .B(_0568_));
 sg13g2_nor2_1 _4348_ (.A(net1242),
    .B(net597),
    .Y(_0122_));
 sg13g2_a21oi_1 _4349_ (.A1(net596),
    .A2(_0567_),
    .Y(_0570_),
    .B1(net1424));
 sg13g2_and3_1 _4350_ (.X(_0571_),
    .A(net1424),
    .B(net1425),
    .C(_0567_));
 sg13g2_nor3_1 _4351_ (.A(net1242),
    .B(_0570_),
    .C(_0571_),
    .Y(_0123_));
 sg13g2_nand3b_1 _4352_ (.B(_0567_),
    .C(net1425),
    .Y(_0572_),
    .A_N(_0051_));
 sg13g2_xor2_1 _4353_ (.B(_0572_),
    .A(net1418),
    .X(_0573_));
 sg13g2_nor2_1 _4354_ (.A(net1242),
    .B(_0573_),
    .Y(_0124_));
 sg13g2_and2_1 _4355_ (.A(net1418),
    .B(_0571_),
    .X(_0574_));
 sg13g2_xnor2_1 _4356_ (.Y(_0575_),
    .A(net1415),
    .B(_0574_));
 sg13g2_nor2_1 _4357_ (.A(net1242),
    .B(_0575_),
    .Y(_0125_));
 sg13g2_nor2b_1 _4358_ (.A(net699),
    .B_N(_0574_),
    .Y(_0576_));
 sg13g2_xnor2_1 _4359_ (.Y(_0577_),
    .A(\dtop.vtop.logo.addr[10] ),
    .B(_0576_));
 sg13g2_nor2_1 _4360_ (.A(net1242),
    .B(net700),
    .Y(_0126_));
 sg13g2_nand3_1 _4361_ (.B(net685),
    .C(_0574_),
    .A(\dtop.vtop.logo.addr[10] ),
    .Y(_0578_));
 sg13g2_xnor2_1 _4362_ (.Y(_0579_),
    .A(_3131_),
    .B(_0578_));
 sg13g2_nor2_1 _4363_ (.A(_0561_),
    .B(net686),
    .Y(_0127_));
 sg13g2_nor2_1 _4364_ (.A(net1369),
    .B(net1346),
    .Y(_0580_));
 sg13g2_nand2b_2 _4365_ (.Y(_0581_),
    .B(_3139_),
    .A_N(_3189_));
 sg13g2_nor2b_2 _4366_ (.A(net1381),
    .B_N(net1378),
    .Y(_0582_));
 sg13g2_nand2b_2 _4367_ (.Y(_0583_),
    .B(net1377),
    .A_N(net1380));
 sg13g2_mux2_1 _4368_ (.A0(_3186_),
    .A1(_0582_),
    .S(_3185_),
    .X(_0584_));
 sg13g2_nand2_1 _4369_ (.Y(_0585_),
    .A(net1327),
    .B(_0584_));
 sg13g2_nor2b_1 _4370_ (.A(net1378),
    .B_N(net1380),
    .Y(_0586_));
 sg13g2_nand2b_2 _4371_ (.Y(_0587_),
    .B(net1380),
    .A_N(net1377));
 sg13g2_nor2_2 _4372_ (.A(net1384),
    .B(net1390),
    .Y(_0588_));
 sg13g2_or2_1 _4373_ (.X(_0589_),
    .B(net1389),
    .A(net1383));
 sg13g2_nor2_1 _4374_ (.A(net1342),
    .B(net1340),
    .Y(_0590_));
 sg13g2_nand2_2 _4375_ (.Y(_0591_),
    .A(net1343),
    .B(_0588_));
 sg13g2_nor2_1 _4376_ (.A(_0581_),
    .B(_0591_),
    .Y(_0592_));
 sg13g2_nor2b_2 _4377_ (.A(net1390),
    .B_N(net1384),
    .Y(_0593_));
 sg13g2_nand2b_1 _4378_ (.Y(_0594_),
    .B(net1383),
    .A_N(net1389));
 sg13g2_nor2_2 _4379_ (.A(net1348),
    .B(net1338),
    .Y(_0595_));
 sg13g2_nor4_1 _4380_ (.A(net1369),
    .B(net1348),
    .C(net1346),
    .D(net1338),
    .Y(_0596_));
 sg13g2_o21ai_1 _4381_ (.B1(net1327),
    .Y(_0597_),
    .A1(_0590_),
    .A2(_0595_));
 sg13g2_and2_1 _4382_ (.A(_0585_),
    .B(_0597_),
    .X(_0598_));
 sg13g2_nor2b_1 _4383_ (.A(net1387),
    .B_N(net1389),
    .Y(_0599_));
 sg13g2_nand2b_1 _4384_ (.Y(_0600_),
    .B(net1389),
    .A_N(net1383));
 sg13g2_nor2_2 _4385_ (.A(net1388),
    .B(net1382),
    .Y(_0601_));
 sg13g2_nor2_1 _4386_ (.A(net1386),
    .B(net1348),
    .Y(_0602_));
 sg13g2_nand2_1 _4387_ (.Y(_0603_),
    .A(net1327),
    .B(_0602_));
 sg13g2_nor4_2 _4388_ (.A(net1369),
    .B(net1348),
    .C(net1346),
    .Y(_0604_),
    .D(net1336));
 sg13g2_nor2_2 _4389_ (.A(_0587_),
    .B(net1337),
    .Y(_0605_));
 sg13g2_nor4_2 _4390_ (.A(net1369),
    .B(net1346),
    .C(net1342),
    .Y(_0606_),
    .D(net1336));
 sg13g2_a21oi_1 _4391_ (.A1(net1327),
    .A2(_0584_),
    .Y(_0607_),
    .B1(_0604_));
 sg13g2_nand3b_1 _4392_ (.B(_0607_),
    .C(_0597_),
    .Y(_0608_),
    .A_N(_0606_));
 sg13g2_nor2b_1 _4393_ (.A(net1372),
    .B_N(net1370),
    .Y(_0609_));
 sg13g2_nand2b_2 _4394_ (.Y(_0610_),
    .B(net1369),
    .A_N(net1371));
 sg13g2_nor2_1 _4395_ (.A(_3140_),
    .B(_0610_),
    .Y(_0611_));
 sg13g2_nand3b_1 _4396_ (.B(net1374),
    .C(net1370),
    .Y(_0612_),
    .A_N(net1372));
 sg13g2_and2_2 _4397_ (.A(net1378),
    .B(net1381),
    .X(_0613_));
 sg13g2_nand2_1 _4398_ (.Y(_0614_),
    .A(net1378),
    .B(net1381));
 sg13g2_nor2_2 _4399_ (.A(net1341),
    .B(net1331),
    .Y(_0615_));
 sg13g2_nor2_2 _4400_ (.A(net1337),
    .B(net1332),
    .Y(_0616_));
 sg13g2_nand2_2 _4401_ (.Y(_0617_),
    .A(_0599_),
    .B(_0613_));
 sg13g2_nor3_1 _4402_ (.A(net1385),
    .B(net1335),
    .C(net1331),
    .Y(_0618_));
 sg13g2_nor4_2 _4403_ (.A(net1367),
    .B(net1347),
    .C(_3189_),
    .Y(_0619_),
    .D(net1336));
 sg13g2_nor3_2 _4404_ (.A(_3190_),
    .B(_0618_),
    .C(_0619_),
    .Y(_0620_));
 sg13g2_nor2b_2 _4405_ (.A(net1370),
    .B_N(net1375),
    .Y(_0621_));
 sg13g2_nand2b_2 _4406_ (.Y(_0622_),
    .B(net1375),
    .A_N(net1369));
 sg13g2_nor2_1 _4407_ (.A(_3141_),
    .B(_0622_),
    .Y(_0623_));
 sg13g2_nand3b_1 _4408_ (.B(net1375),
    .C(net1371),
    .Y(_0624_),
    .A_N(net1370));
 sg13g2_nor2_1 _4409_ (.A(net1372),
    .B(_0622_),
    .Y(_0625_));
 sg13g2_nand2_2 _4410_ (.Y(_0626_),
    .A(_3141_),
    .B(_0621_));
 sg13g2_nor2_1 _4411_ (.A(net1339),
    .B(net1332),
    .Y(_0627_));
 sg13g2_nand2_2 _4412_ (.Y(_0628_),
    .A(_0593_),
    .B(_0613_));
 sg13g2_nor4_2 _4413_ (.A(net1371),
    .B(net1338),
    .C(net1333),
    .Y(_0629_),
    .D(_0622_));
 sg13g2_and2_1 _4414_ (.A(net1385),
    .B(_0582_),
    .X(_0630_));
 sg13g2_nand3b_1 _4415_ (.B(net1377),
    .C(net1383),
    .Y(_0631_),
    .A_N(net1380));
 sg13g2_nor2_1 _4416_ (.A(net1389),
    .B(_0631_),
    .Y(_0632_));
 sg13g2_nand2_1 _4417_ (.Y(_0633_),
    .A(_0582_),
    .B(_0593_));
 sg13g2_nor3_1 _4418_ (.A(net1389),
    .B(net1329),
    .C(_0631_),
    .Y(_0634_));
 sg13g2_nor2_1 _4419_ (.A(_0629_),
    .B(_0634_),
    .Y(_0635_));
 sg13g2_nand2_1 _4420_ (.Y(_0636_),
    .A(_0620_),
    .B(_0635_));
 sg13g2_nor2_2 _4421_ (.A(net1376),
    .B(net1373),
    .Y(_0637_));
 sg13g2_nor2_2 _4422_ (.A(net1374),
    .B(_0610_),
    .Y(_0638_));
 sg13g2_nand2_2 _4423_ (.Y(_0639_),
    .A(_3140_),
    .B(_0609_));
 sg13g2_nor2_2 _4424_ (.A(_0583_),
    .B(net1337),
    .Y(_0640_));
 sg13g2_nor4_2 _4425_ (.A(_3184_),
    .B(_0583_),
    .C(_0588_),
    .Y(_0641_),
    .D(net1319));
 sg13g2_a22oi_1 _4426_ (.Y(_0642_),
    .B1(_0615_),
    .B2(_0638_),
    .A2(net1325),
    .A1(_0590_));
 sg13g2_o21ai_1 _4427_ (.B1(_0642_),
    .Y(_0643_),
    .A1(net1330),
    .A2(_0628_));
 sg13g2_or2_1 _4428_ (.X(_0644_),
    .B(_0643_),
    .A(_0641_));
 sg13g2_nor2_2 _4429_ (.A(_0587_),
    .B(net1339),
    .Y(_0645_));
 sg13g2_nand2_2 _4430_ (.Y(_0646_),
    .A(_0586_),
    .B(_0593_));
 sg13g2_nor4_2 _4431_ (.A(net1371),
    .B(net1342),
    .C(net1339),
    .Y(_0647_),
    .D(_0622_));
 sg13g2_nor2_2 _4432_ (.A(_3185_),
    .B(net1342),
    .Y(_0648_));
 sg13g2_nand2_1 _4433_ (.Y(_0649_),
    .A(_3184_),
    .B(net1343));
 sg13g2_nand2_1 _4434_ (.Y(_0650_),
    .A(_0625_),
    .B(_0648_));
 sg13g2_nand3_1 _4435_ (.B(net1343),
    .C(net1321),
    .A(net1385),
    .Y(_0651_));
 sg13g2_nor2_1 _4436_ (.A(_3188_),
    .B(_0639_),
    .Y(_0652_));
 sg13g2_nor2_1 _4437_ (.A(net1349),
    .B(net1332),
    .Y(_0653_));
 sg13g2_nand4_1 _4438_ (.B(net1390),
    .C(net1377),
    .A(net1384),
    .Y(_0654_),
    .D(net1380));
 sg13g2_a21oi_2 _4439_ (.B1(net1319),
    .Y(_0655_),
    .A2(_0654_),
    .A1(_3188_));
 sg13g2_nand2_1 _4440_ (.Y(_0656_),
    .A(net1343),
    .B(net1323));
 sg13g2_nor2_2 _4441_ (.A(net1330),
    .B(_0646_),
    .Y(_0657_));
 sg13g2_nand2_1 _4442_ (.Y(_0658_),
    .A(net1322),
    .B(_0645_));
 sg13g2_nand4_1 _4443_ (.B(_3184_),
    .C(net1343),
    .A(net1371),
    .Y(_0659_),
    .D(_0621_));
 sg13g2_nor2_2 _4444_ (.A(_3136_),
    .B(_0631_),
    .Y(_0660_));
 sg13g2_nand2_2 _4445_ (.Y(_0661_),
    .A(_3184_),
    .B(_0582_));
 sg13g2_nor3_2 _4446_ (.A(net1374),
    .B(_0610_),
    .C(_0631_),
    .Y(_0662_));
 sg13g2_nor3_2 _4447_ (.A(net1386),
    .B(net1348),
    .C(net1329),
    .Y(_0663_));
 sg13g2_nor2_2 _4448_ (.A(net1384),
    .B(_0583_),
    .Y(_0664_));
 sg13g2_nor2_1 _4449_ (.A(_0591_),
    .B(net1319),
    .Y(_0665_));
 sg13g2_nor2_1 _4450_ (.A(_0617_),
    .B(_0626_),
    .Y(_0666_));
 sg13g2_nor4_2 _4451_ (.A(net1387),
    .B(net1372),
    .C(net1331),
    .Y(_0667_),
    .D(_0622_));
 sg13g2_nor2_1 _4452_ (.A(net1329),
    .B(_0654_),
    .Y(_0668_));
 sg13g2_nor4_2 _4453_ (.A(net1386),
    .B(net1389),
    .C(net1377),
    .Y(_0669_),
    .D(net1380));
 sg13g2_nor4_2 _4454_ (.A(net1374),
    .B(net1347),
    .C(net1340),
    .Y(_0670_),
    .D(_0610_));
 sg13g2_nor2_1 _4455_ (.A(_0668_),
    .B(_0670_),
    .Y(_0671_));
 sg13g2_nand2_1 _4456_ (.Y(_0672_),
    .A(net1321),
    .B(net1318));
 sg13g2_nor4_2 _4457_ (.A(net1384),
    .B(net1374),
    .C(_0583_),
    .Y(_0673_),
    .D(_0610_));
 sg13g2_nand2_1 _4458_ (.Y(_0674_),
    .A(_3136_),
    .B(_0673_));
 sg13g2_o21ai_1 _4459_ (.B1(net1326),
    .Y(_0675_),
    .A1(_0630_),
    .A2(net1318));
 sg13g2_and2_1 _4460_ (.A(net1367),
    .B(_0637_),
    .X(_0676_));
 sg13g2_nand2_1 _4461_ (.Y(_0677_),
    .A(net1367),
    .B(_0637_));
 sg13g2_nor2_2 _4462_ (.A(net1319),
    .B(_0646_),
    .Y(_0678_));
 sg13g2_and2_1 _4463_ (.A(_0605_),
    .B(_0638_),
    .X(_0679_));
 sg13g2_nor2_1 _4464_ (.A(_0628_),
    .B(_0639_),
    .Y(_0680_));
 sg13g2_a21oi_1 _4465_ (.A1(_0628_),
    .A2(_0649_),
    .Y(_0681_),
    .B1(net1319));
 sg13g2_o21ai_1 _4466_ (.B1(net1326),
    .Y(_0682_),
    .A1(_0616_),
    .A2(_0645_));
 sg13g2_nand2_1 _4467_ (.Y(_0683_),
    .A(net1320),
    .B(_0630_));
 sg13g2_a22oi_1 _4468_ (.Y(_0684_),
    .B1(_0660_),
    .B2(net1327),
    .A2(_0632_),
    .A1(net1321));
 sg13g2_nor3_2 _4469_ (.A(net1340),
    .B(net1331),
    .C(net1329),
    .Y(_0685_));
 sg13g2_nand2_1 _4470_ (.Y(_0686_),
    .A(net1322),
    .B(_0660_));
 sg13g2_nand2_1 _4471_ (.Y(_0687_),
    .A(_0605_),
    .B(net1320));
 sg13g2_nand3_1 _4472_ (.B(net1340),
    .C(_0613_),
    .A(net1327),
    .Y(_0688_));
 sg13g2_a221oi_1 _4473_ (.B2(net1322),
    .C1(_0685_),
    .B1(_0660_),
    .A1(_0605_),
    .Y(_0689_),
    .A2(net1321));
 sg13g2_nand3_1 _4474_ (.B(_0688_),
    .C(_0689_),
    .A(_0684_),
    .Y(_0690_));
 sg13g2_nor4_2 _4475_ (.A(net1367),
    .B(net1347),
    .C(_3189_),
    .Y(_0691_),
    .D(net1340));
 sg13g2_nor2_1 _4476_ (.A(net1334),
    .B(_0654_),
    .Y(_0692_));
 sg13g2_nor3_2 _4477_ (.A(net1348),
    .B(net1339),
    .C(net1329),
    .Y(_0693_));
 sg13g2_nor4_2 _4478_ (.A(net1368),
    .B(_3187_),
    .C(net1346),
    .Y(_0694_),
    .D(net1338));
 sg13g2_or2_1 _4479_ (.X(_0695_),
    .B(_0694_),
    .A(_0693_));
 sg13g2_a221oi_1 _4480_ (.B2(_0638_),
    .C1(_0695_),
    .B1(_0616_),
    .A1(_0605_),
    .Y(_0696_),
    .A2(net1325));
 sg13g2_nor4_2 _4481_ (.A(net1374),
    .B(net1347),
    .C(net1336),
    .Y(_0697_),
    .D(_0610_));
 sg13g2_nor3_1 _4482_ (.A(net1342),
    .B(net1341),
    .C(net1330),
    .Y(_0698_));
 sg13g2_or2_1 _4483_ (.X(_0699_),
    .B(_0698_),
    .A(_0697_));
 sg13g2_nor4_2 _4484_ (.A(net1374),
    .B(net1347),
    .C(net1338),
    .Y(_0700_),
    .D(_0610_));
 sg13g2_nor3_2 _4485_ (.A(net1342),
    .B(net1336),
    .C(net1329),
    .Y(_0701_));
 sg13g2_inv_1 _4486_ (.Y(_0702_),
    .A(_0701_));
 sg13g2_nor2_1 _4487_ (.A(_0697_),
    .B(_0700_),
    .Y(_0703_));
 sg13g2_nor4_1 _4488_ (.A(_0697_),
    .B(_0698_),
    .C(_0700_),
    .D(_0701_),
    .Y(_0704_));
 sg13g2_o21ai_1 _4489_ (.B1(net1326),
    .Y(_0705_),
    .A1(_0648_),
    .A2(_0669_));
 sg13g2_a21oi_1 _4490_ (.A1(_0591_),
    .A2(_0661_),
    .Y(_0706_),
    .B1(net1319));
 sg13g2_a22oi_1 _4491_ (.Y(_0707_),
    .B1(_0664_),
    .B2(_0621_),
    .A2(net1323),
    .A1(_0616_));
 sg13g2_nand2_1 _4492_ (.Y(_0708_),
    .A(_0651_),
    .B(_0675_));
 sg13g2_a21oi_1 _4493_ (.A1(_3186_),
    .A2(net1321),
    .Y(_0709_),
    .B1(_0663_));
 sg13g2_nand4_1 _4494_ (.B(_0674_),
    .C(_0677_),
    .A(net1335),
    .Y(_0710_),
    .D(_0707_));
 sg13g2_nor4_1 _4495_ (.A(_0655_),
    .B(_0678_),
    .C(_0679_),
    .D(_0710_),
    .Y(_0711_));
 sg13g2_nand4_1 _4496_ (.B(_0696_),
    .C(_0709_),
    .A(_0603_),
    .Y(_0712_),
    .D(_0711_));
 sg13g2_nor3_1 _4497_ (.A(_0667_),
    .B(_0706_),
    .C(_0708_),
    .Y(_0713_));
 sg13g2_nor3_1 _4498_ (.A(_0681_),
    .B(_0691_),
    .C(_0692_),
    .Y(_0714_));
 sg13g2_nand4_1 _4499_ (.B(_0703_),
    .C(_0713_),
    .A(_0672_),
    .Y(_0715_),
    .D(_0714_));
 sg13g2_nand4_1 _4500_ (.B(_0671_),
    .C(_0682_),
    .A(_0656_),
    .Y(_0716_),
    .D(_0705_));
 sg13g2_nor4_1 _4501_ (.A(_0690_),
    .B(_0712_),
    .C(_0715_),
    .D(_0716_),
    .Y(_0717_));
 sg13g2_nor3_1 _4502_ (.A(_0608_),
    .B(_0636_),
    .C(_0644_),
    .Y(_0718_));
 sg13g2_nand2_1 _4503_ (.Y(_0719_),
    .A(_0717_),
    .B(_0718_));
 sg13g2_nor3_2 _4504_ (.A(net1338),
    .B(net1334),
    .C(net1331),
    .Y(_0720_));
 sg13g2_nor2_2 _4505_ (.A(net1334),
    .B(_0646_),
    .Y(_0721_));
 sg13g2_nand2_1 _4506_ (.Y(_0722_),
    .A(net1324),
    .B(_0645_));
 sg13g2_nor4_1 _4507_ (.A(_0644_),
    .B(_0694_),
    .C(_0720_),
    .D(_0721_),
    .Y(_0723_));
 sg13g2_and2_1 _4508_ (.A(_0719_),
    .B(_0723_),
    .X(_0724_));
 sg13g2_o21ai_1 _4509_ (.B1(_3320_),
    .Y(_0725_),
    .A1(_3145_),
    .A2(_3281_));
 sg13g2_and2_1 _4510_ (.A(_3324_),
    .B(_0725_),
    .X(_0726_));
 sg13g2_nand2_1 _4511_ (.Y(_0727_),
    .A(net1328),
    .B(_0725_));
 sg13g2_nor3_2 _4512_ (.A(net1396),
    .B(net1395),
    .C(net1394),
    .Y(_0728_));
 sg13g2_or3_2 _4513_ (.A(net1396),
    .B(net1395),
    .C(net1394),
    .X(_0729_));
 sg13g2_and2_2 _4514_ (.A(net1345),
    .B(_0729_),
    .X(_0730_));
 sg13g2_or4_2 _4515_ (.A(_3146_),
    .B(_3320_),
    .C(_3322_),
    .D(_3323_),
    .X(_0731_));
 sg13g2_and2_1 _4516_ (.A(_0730_),
    .B(_0731_),
    .X(_0732_));
 sg13g2_nand2_2 _4517_ (.Y(_0733_),
    .A(_0730_),
    .B(_0731_));
 sg13g2_a22oi_1 _4518_ (.Y(_0734_),
    .B1(_0730_),
    .B2(_0731_),
    .A2(_0725_),
    .A1(net1328));
 sg13g2_and2_2 _4519_ (.A(net1401),
    .B(net1402),
    .X(_0735_));
 sg13g2_nand2_2 _4520_ (.Y(_0736_),
    .A(net1401),
    .B(net1402));
 sg13g2_nand3_1 _4521_ (.B(net1300),
    .C(_0735_),
    .A(_3322_),
    .Y(_0737_));
 sg13g2_nand2_1 _4522_ (.Y(_0738_),
    .A(_0000_),
    .B(_3210_));
 sg13g2_xnor2_1 _4523_ (.Y(_0739_),
    .A(_0090_),
    .B(_0735_));
 sg13g2_o21ai_1 _4524_ (.B1(_3321_),
    .Y(_0740_),
    .A1(net1397),
    .A2(_0728_));
 sg13g2_inv_1 _4525_ (.Y(_0741_),
    .A(_0740_));
 sg13g2_nand3_1 _4526_ (.B(net1322),
    .C(_0627_),
    .A(net1282),
    .Y(_0742_));
 sg13g2_nand3_1 _4527_ (.B(_0728_),
    .C(_0739_),
    .A(_0641_),
    .Y(_0743_));
 sg13g2_a22oi_1 _4528_ (.Y(_0744_),
    .B1(_0741_),
    .B2(_0720_),
    .A2(_0721_),
    .A1(_0436_));
 sg13g2_nand3_1 _4529_ (.B(_0743_),
    .C(_0744_),
    .A(_0742_),
    .Y(_0745_));
 sg13g2_a21oi_1 _4530_ (.A1(net1344),
    .A2(_0737_),
    .Y(_0746_),
    .B1(_0642_));
 sg13g2_a221oi_1 _4531_ (.B2(_0746_),
    .C1(_0745_),
    .B1(_0738_),
    .A1(net1446),
    .Y(_0747_),
    .A2(_0694_));
 sg13g2_o21ai_1 _4532_ (.B1(_0747_),
    .Y(_0748_),
    .A1(_0436_),
    .A2(_0719_));
 sg13g2_o21ai_1 _4533_ (.B1(net1362),
    .Y(_0749_),
    .A1(_0724_),
    .A2(_0748_));
 sg13g2_nor2_2 _4534_ (.A(_0087_),
    .B(_0749_),
    .Y(_0750_));
 sg13g2_nand4_1 _4535_ (.B(net1343),
    .C(_0593_),
    .A(net1367),
    .Y(_0751_),
    .D(_0637_));
 sg13g2_nor3_1 _4536_ (.A(net1347),
    .B(net1336),
    .C(net1335),
    .Y(_0752_));
 sg13g2_nor3_1 _4537_ (.A(_0629_),
    .B(_0634_),
    .C(_0752_),
    .Y(_0753_));
 sg13g2_o21ai_1 _4538_ (.B1(_0753_),
    .Y(_0754_),
    .A1(net1319),
    .A2(_0649_));
 sg13g2_nand2b_1 _4539_ (.Y(_0755_),
    .B(_0751_),
    .A_N(_0754_));
 sg13g2_nand2_2 _4540_ (.Y(_0756_),
    .A(_0750_),
    .B(_0755_));
 sg13g2_o21ai_1 _4541_ (.B1(net1436),
    .Y(_0757_),
    .A1(\dtop.player_inst.synth.alu.acc[0] ),
    .A2(net1139));
 sg13g2_a21oi_1 _4542_ (.A1(_3119_),
    .A2(net1139),
    .Y(_0128_),
    .B1(_0757_));
 sg13g2_o21ai_1 _4543_ (.B1(net1434),
    .Y(_0758_),
    .A1(\dtop.player_inst.synth.alu.acc[1] ),
    .A2(net1140));
 sg13g2_a21oi_1 _4544_ (.A1(_3118_),
    .A2(net1140),
    .Y(_0129_),
    .B1(_0758_));
 sg13g2_o21ai_1 _4545_ (.B1(net1434),
    .Y(_0759_),
    .A1(\dtop.player_inst.synth.alu.acc[2] ),
    .A2(net1140));
 sg13g2_a21oi_1 _4546_ (.A1(_3117_),
    .A2(net1141),
    .Y(_0130_),
    .B1(_0759_));
 sg13g2_o21ai_1 _4547_ (.B1(net1434),
    .Y(_0760_),
    .A1(\dtop.player_inst.synth.alu.acc[3] ),
    .A2(net1140));
 sg13g2_a21oi_1 _4548_ (.A1(_3116_),
    .A2(net1140),
    .Y(_0131_),
    .B1(_0760_));
 sg13g2_o21ai_1 _4549_ (.B1(net1436),
    .Y(_0761_),
    .A1(\dtop.player_inst.synth.alu.acc[4] ),
    .A2(net1139));
 sg13g2_a21oi_1 _4550_ (.A1(_3115_),
    .A2(net1142),
    .Y(_0132_),
    .B1(_0761_));
 sg13g2_o21ai_1 _4551_ (.B1(net1434),
    .Y(_0762_),
    .A1(\dtop.player_inst.synth.alu.acc[5] ),
    .A2(net1140));
 sg13g2_a21oi_1 _4552_ (.A1(_3114_),
    .A2(net1140),
    .Y(_0133_),
    .B1(_0762_));
 sg13g2_o21ai_1 _4553_ (.B1(net1436),
    .Y(_0763_),
    .A1(\dtop.player_inst.synth.alu.acc[6] ),
    .A2(net1139));
 sg13g2_a21oi_1 _4554_ (.A1(_3113_),
    .A2(net1139),
    .Y(_0134_),
    .B1(_0763_));
 sg13g2_o21ai_1 _4555_ (.B1(net1434),
    .Y(_0764_),
    .A1(net1408),
    .A2(net1141));
 sg13g2_a21oi_1 _4556_ (.A1(_3112_),
    .A2(net1141),
    .Y(_0135_),
    .B1(_0764_));
 sg13g2_o21ai_1 _4557_ (.B1(net1436),
    .Y(_0765_),
    .A1(\dtop.player_inst.synth.alu.acc[8] ),
    .A2(net1142));
 sg13g2_a21oi_1 _4558_ (.A1(_3111_),
    .A2(net1139),
    .Y(_0136_),
    .B1(_0765_));
 sg13g2_o21ai_1 _4559_ (.B1(net1434),
    .Y(_0766_),
    .A1(\dtop.player_inst.synth.alu.acc[9] ),
    .A2(net1140));
 sg13g2_a21oi_1 _4560_ (.A1(_3110_),
    .A2(net1141),
    .Y(_0137_),
    .B1(_0766_));
 sg13g2_o21ai_1 _4561_ (.B1(net1436),
    .Y(_0767_),
    .A1(net1407),
    .A2(net1139));
 sg13g2_a21oi_1 _4562_ (.A1(_3109_),
    .A2(net1139),
    .Y(_0138_),
    .B1(_0767_));
 sg13g2_nor3_2 _4563_ (.A(_0583_),
    .B(net1336),
    .C(net1329),
    .Y(_0768_));
 sg13g2_nand2_1 _4564_ (.Y(_0769_),
    .A(_0750_),
    .B(_0768_));
 sg13g2_o21ai_1 _4565_ (.B1(net1427),
    .Y(_0770_),
    .A1(net1414),
    .A2(net1137));
 sg13g2_a21oi_1 _4566_ (.A1(_3108_),
    .A2(net1137),
    .Y(_0139_),
    .B1(_0770_));
 sg13g2_o21ai_1 _4567_ (.B1(net1428),
    .Y(_0771_),
    .A1(net1413),
    .A2(net1137));
 sg13g2_a21oi_1 _4568_ (.A1(_3107_),
    .A2(net1137),
    .Y(_0140_),
    .B1(_0771_));
 sg13g2_o21ai_1 _4569_ (.B1(net1427),
    .Y(_0772_),
    .A1(net1412),
    .A2(net1136));
 sg13g2_a21oi_1 _4570_ (.A1(_3106_),
    .A2(net1136),
    .Y(_0141_),
    .B1(_0772_));
 sg13g2_o21ai_1 _4571_ (.B1(net1429),
    .Y(_0773_),
    .A1(net1411),
    .A2(net1136));
 sg13g2_a21oi_1 _4572_ (.A1(_3105_),
    .A2(net1136),
    .Y(_0142_),
    .B1(_0773_));
 sg13g2_o21ai_1 _4573_ (.B1(net1429),
    .Y(_0774_),
    .A1(net1410),
    .A2(net1136));
 sg13g2_a21oi_1 _4574_ (.A1(_3104_),
    .A2(net1136),
    .Y(_0143_),
    .B1(_0774_));
 sg13g2_o21ai_1 _4575_ (.B1(net1433),
    .Y(_0775_),
    .A1(\dtop.player_inst.synth.alu.acc[5] ),
    .A2(net1138));
 sg13g2_a21oi_1 _4576_ (.A1(_3103_),
    .A2(net1138),
    .Y(_0144_),
    .B1(_0775_));
 sg13g2_o21ai_1 _4577_ (.B1(net1429),
    .Y(_0776_),
    .A1(net1409),
    .A2(net1136));
 sg13g2_a21oi_1 _4578_ (.A1(_3102_),
    .A2(net1136),
    .Y(_0145_),
    .B1(_0776_));
 sg13g2_o21ai_1 _4579_ (.B1(net1433),
    .Y(_0777_),
    .A1(net1408),
    .A2(net1138));
 sg13g2_a21oi_1 _4580_ (.A1(_3101_),
    .A2(net1138),
    .Y(_0146_),
    .B1(_0777_));
 sg13g2_nor2_2 _4581_ (.A(_3144_),
    .B(_0749_),
    .Y(_0778_));
 sg13g2_nand3_1 _4582_ (.B(_0616_),
    .C(_0778_),
    .A(net1324),
    .Y(_0779_));
 sg13g2_nand3_1 _4583_ (.B(net1437),
    .C(net1134),
    .A(net436),
    .Y(_0780_));
 sg13g2_o21ai_1 _4584_ (.B1(_0780_),
    .Y(_0147_),
    .A1(_3083_),
    .A2(net1134));
 sg13g2_nand3_1 _4585_ (.B(net1437),
    .C(net1134),
    .A(net408),
    .Y(_0781_));
 sg13g2_o21ai_1 _4586_ (.B1(_0781_),
    .Y(_0148_),
    .A1(_3082_),
    .A2(net1134));
 sg13g2_nand3_1 _4587_ (.B(net1427),
    .C(net1132),
    .A(net420),
    .Y(_0782_));
 sg13g2_o21ai_1 _4588_ (.B1(_0782_),
    .Y(_0149_),
    .A1(_3081_),
    .A2(net1132));
 sg13g2_nand3_1 _4589_ (.B(net1433),
    .C(net1135),
    .A(net423),
    .Y(_0783_));
 sg13g2_o21ai_1 _4590_ (.B1(_0783_),
    .Y(_0150_),
    .A1(_3080_),
    .A2(net1135));
 sg13g2_nand3_1 _4591_ (.B(net1427),
    .C(net1132),
    .A(net406),
    .Y(_0784_));
 sg13g2_o21ai_1 _4592_ (.B1(_0784_),
    .Y(_0151_),
    .A1(_3079_),
    .A2(net1132));
 sg13g2_nand3_1 _4593_ (.B(net1438),
    .C(net1133),
    .A(net505),
    .Y(_0785_));
 sg13g2_o21ai_1 _4594_ (.B1(_0785_),
    .Y(_0152_),
    .A1(_3078_),
    .A2(net1133));
 sg13g2_nand3_1 _4595_ (.B(net1433),
    .C(net1132),
    .A(net380),
    .Y(_0786_));
 sg13g2_o21ai_1 _4596_ (.B1(_0786_),
    .Y(_0153_),
    .A1(_3077_),
    .A2(net1132));
 sg13g2_nand3_1 _4597_ (.B(net1431),
    .C(net1132),
    .A(net444),
    .Y(_0787_));
 sg13g2_o21ai_1 _4598_ (.B1(_0787_),
    .Y(_0154_),
    .A1(_3076_),
    .A2(net1132));
 sg13g2_nand3_1 _4599_ (.B(net1435),
    .C(net1133),
    .A(net434),
    .Y(_0788_));
 sg13g2_o21ai_1 _4600_ (.B1(_0788_),
    .Y(_0155_),
    .A1(_3093_),
    .A2(net1133));
 sg13g2_nand3_1 _4601_ (.B(net1435),
    .C(net1133),
    .A(net480),
    .Y(_0789_));
 sg13g2_o21ai_1 _4602_ (.B1(_0789_),
    .Y(_0156_),
    .A1(_3092_),
    .A2(net1133));
 sg13g2_nand3_1 _4603_ (.B(net1434),
    .C(net1133),
    .A(net442),
    .Y(_0790_));
 sg13g2_o21ai_1 _4604_ (.B1(_0790_),
    .Y(_0157_),
    .A1(_3091_),
    .A2(net1133));
 sg13g2_nand2_1 _4605_ (.Y(_0791_),
    .A(_0595_),
    .B(net1324));
 sg13g2_a221oi_1 _4606_ (.B2(_0653_),
    .C1(_0673_),
    .B1(_0638_),
    .A1(_0615_),
    .Y(_0792_),
    .A2(net1320));
 sg13g2_and2_1 _4607_ (.A(_0791_),
    .B(_0792_),
    .X(_0793_));
 sg13g2_o21ai_1 _4608_ (.B1(net1321),
    .Y(_0794_),
    .A1(_0595_),
    .A2(_0601_));
 sg13g2_o21ai_1 _4609_ (.B1(_0631_),
    .Y(_0795_),
    .A1(net1340),
    .A2(net1331));
 sg13g2_nand2_1 _4610_ (.Y(_0796_),
    .A(net1317),
    .B(_0795_));
 sg13g2_nand2_1 _4611_ (.Y(_0797_),
    .A(_0794_),
    .B(_0796_));
 sg13g2_nor2_1 _4612_ (.A(_3188_),
    .B(_0626_),
    .Y(_0798_));
 sg13g2_nor3_2 _4613_ (.A(net1349),
    .B(net1348),
    .C(net1334),
    .Y(_0799_));
 sg13g2_nand2b_2 _4614_ (.Y(_0800_),
    .B(_0669_),
    .A_N(net1334));
 sg13g2_o21ai_1 _4615_ (.B1(_0800_),
    .Y(_0801_),
    .A1(_0617_),
    .A2(_0626_));
 sg13g2_nand2_1 _4616_ (.Y(_0802_),
    .A(_0627_),
    .B(net1316));
 sg13g2_o21ai_1 _4617_ (.B1(_0802_),
    .Y(_0803_),
    .A1(_0581_),
    .A2(_0646_));
 sg13g2_a22oi_1 _4618_ (.Y(_0804_),
    .B1(net1318),
    .B2(net1316),
    .A2(_0648_),
    .A1(net1326));
 sg13g2_inv_1 _4619_ (.Y(_0805_),
    .A(_0804_));
 sg13g2_nor2_1 _4620_ (.A(_0803_),
    .B(_0805_),
    .Y(_0806_));
 sg13g2_a21oi_1 _4621_ (.A1(_0617_),
    .A2(_0628_),
    .Y(_0807_),
    .B1(net1330));
 sg13g2_nor3_1 _4622_ (.A(net1386),
    .B(net1342),
    .C(net1334),
    .Y(_0808_));
 sg13g2_nor2_1 _4623_ (.A(_0807_),
    .B(_0808_),
    .Y(_0809_));
 sg13g2_nor2_1 _4624_ (.A(_0797_),
    .B(_0801_),
    .Y(_0810_));
 sg13g2_a21oi_1 _4625_ (.A1(_0621_),
    .A2(net1318),
    .Y(_0811_),
    .B1(_0697_));
 sg13g2_nand4_1 _4626_ (.B(_0651_),
    .C(_0810_),
    .A(_0598_),
    .Y(_0812_),
    .D(_0811_));
 sg13g2_nor2_1 _4627_ (.A(_0798_),
    .B(_0799_),
    .Y(_0813_));
 sg13g2_and2_1 _4628_ (.A(_0603_),
    .B(_0813_),
    .X(_0814_));
 sg13g2_nand4_1 _4629_ (.B(_0806_),
    .C(_0809_),
    .A(_0793_),
    .Y(_0815_),
    .D(_0814_));
 sg13g2_nor3_2 _4630_ (.A(_0690_),
    .B(_0812_),
    .C(_0815_),
    .Y(_0816_));
 sg13g2_nor4_2 _4631_ (.A(_0691_),
    .B(_0692_),
    .C(_0694_),
    .Y(_0817_),
    .D(_0720_));
 sg13g2_a21oi_1 _4632_ (.A1(net1349),
    .A2(net1341),
    .Y(_0818_),
    .B1(net1342));
 sg13g2_o21ai_1 _4633_ (.B1(net1316),
    .Y(_0819_),
    .A1(_0664_),
    .A2(_0818_));
 sg13g2_nor2_1 _4634_ (.A(_0662_),
    .B(_0663_),
    .Y(_0820_));
 sg13g2_nor3_1 _4635_ (.A(net1384),
    .B(net1332),
    .C(_0639_),
    .Y(_0821_));
 sg13g2_nor3_1 _4636_ (.A(_0693_),
    .B(_0698_),
    .C(_0821_),
    .Y(_0822_));
 sg13g2_nand4_1 _4637_ (.B(_0819_),
    .C(_0820_),
    .A(_0817_),
    .Y(_0823_),
    .D(_0822_));
 sg13g2_nor3_1 _4638_ (.A(_0583_),
    .B(net1337),
    .C(net1334),
    .Y(_0824_));
 sg13g2_a221oi_1 _4639_ (.B2(net1323),
    .C1(_0700_),
    .B1(_0664_),
    .A1(net1324),
    .Y(_0825_),
    .A2(_0640_));
 sg13g2_a221oi_1 _4640_ (.B2(_3186_),
    .C1(_3190_),
    .B1(net1317),
    .A1(net1343),
    .Y(_0826_),
    .A2(net1323));
 sg13g2_nor2b_1 _4641_ (.A(_0618_),
    .B_N(_0826_),
    .Y(_0827_));
 sg13g2_nand3b_1 _4642_ (.B(_0825_),
    .C(_0827_),
    .Y(_0828_),
    .A_N(_0755_));
 sg13g2_nor3_1 _4643_ (.A(net1349),
    .B(net1348),
    .C(net1329),
    .Y(_0829_));
 sg13g2_nor4_2 _4644_ (.A(net1369),
    .B(net1346),
    .C(net1340),
    .Y(_0830_),
    .D(net1331));
 sg13g2_nor4_2 _4645_ (.A(_0606_),
    .B(_0670_),
    .C(_0829_),
    .Y(_0831_),
    .D(_0830_));
 sg13g2_a21oi_1 _4646_ (.A1(_0591_),
    .A2(_0661_),
    .Y(_0832_),
    .B1(_0626_));
 sg13g2_nor2_1 _4647_ (.A(_0619_),
    .B(_0680_),
    .Y(_0833_));
 sg13g2_nand2_1 _4648_ (.Y(_0834_),
    .A(_0722_),
    .B(_0831_));
 sg13g2_a21oi_1 _4649_ (.A1(_0616_),
    .A2(net1317),
    .Y(_0835_),
    .B1(_0832_));
 sg13g2_nand4_1 _4650_ (.B(_0831_),
    .C(_0833_),
    .A(_0722_),
    .Y(_0836_),
    .D(_0835_));
 sg13g2_nor2_1 _4651_ (.A(net1335),
    .B(_0649_),
    .Y(_0837_));
 sg13g2_nor2_2 _4652_ (.A(_0583_),
    .B(net1341),
    .Y(_0838_));
 sg13g2_nor3_1 _4653_ (.A(_0583_),
    .B(net1341),
    .C(net1335),
    .Y(_0839_));
 sg13g2_a221oi_1 _4654_ (.B2(_0645_),
    .C1(_0652_),
    .B1(_0638_),
    .A1(net1324),
    .Y(_0840_),
    .A2(_0630_));
 sg13g2_nor4_1 _4655_ (.A(_0665_),
    .B(_0679_),
    .C(_0837_),
    .D(_0839_),
    .Y(_0841_));
 sg13g2_nand2_1 _4656_ (.Y(_0842_),
    .A(_0840_),
    .B(_0841_));
 sg13g2_nor4_1 _4657_ (.A(_0823_),
    .B(_0828_),
    .C(_0836_),
    .D(_0842_),
    .Y(_0843_));
 sg13g2_and3_1 _4658_ (.X(_0844_),
    .A(_0778_),
    .B(_0816_),
    .C(_0843_));
 sg13g2_o21ai_1 _4659_ (.B1(net1437),
    .Y(_0845_),
    .A1(net546),
    .A2(net1130));
 sg13g2_a21oi_1 _4660_ (.A1(_3083_),
    .A2(net1130),
    .Y(_0158_),
    .B1(_0845_));
 sg13g2_o21ai_1 _4661_ (.B1(net1437),
    .Y(_0846_),
    .A1(net542),
    .A2(net1130));
 sg13g2_a21oi_1 _4662_ (.A1(_3082_),
    .A2(net1129),
    .Y(_0159_),
    .B1(_0846_));
 sg13g2_o21ai_1 _4663_ (.B1(net1433),
    .Y(_0847_),
    .A1(net548),
    .A2(net1128));
 sg13g2_a21oi_1 _4664_ (.A1(_3081_),
    .A2(net1128),
    .Y(_0160_),
    .B1(_0847_));
 sg13g2_o21ai_1 _4665_ (.B1(net1431),
    .Y(_0848_),
    .A1(net585),
    .A2(net1131));
 sg13g2_a21oi_1 _4666_ (.A1(_3080_),
    .A2(net1131),
    .Y(_0161_),
    .B1(_0848_));
 sg13g2_o21ai_1 _4667_ (.B1(net1428),
    .Y(_0849_),
    .A1(net588),
    .A2(net1128));
 sg13g2_a21oi_1 _4668_ (.A1(_3079_),
    .A2(net1128),
    .Y(_0162_),
    .B1(_0849_));
 sg13g2_o21ai_1 _4669_ (.B1(net1438),
    .Y(_0850_),
    .A1(net584),
    .A2(net1129));
 sg13g2_a21oi_1 _4670_ (.A1(_3078_),
    .A2(net1130),
    .Y(_0163_),
    .B1(_0850_));
 sg13g2_o21ai_1 _4671_ (.B1(net1433),
    .Y(_0851_),
    .A1(net549),
    .A2(net1128));
 sg13g2_a21oi_1 _4672_ (.A1(_3077_),
    .A2(net1128),
    .Y(_0164_),
    .B1(_0851_));
 sg13g2_o21ai_1 _4673_ (.B1(net1431),
    .Y(_0852_),
    .A1(net560),
    .A2(net1128));
 sg13g2_a21oi_1 _4674_ (.A1(_3076_),
    .A2(net1128),
    .Y(_0165_),
    .B1(_0852_));
 sg13g2_o21ai_1 _4675_ (.B1(net1435),
    .Y(_0853_),
    .A1(net540),
    .A2(net1129));
 sg13g2_a21oi_1 _4676_ (.A1(_3093_),
    .A2(net1129),
    .Y(_0166_),
    .B1(_0853_));
 sg13g2_o21ai_1 _4677_ (.B1(net1434),
    .Y(_0854_),
    .A1(net586),
    .A2(net1129));
 sg13g2_a21oi_1 _4678_ (.A1(_3092_),
    .A2(net1129),
    .Y(_0167_),
    .B1(_0854_));
 sg13g2_o21ai_1 _4679_ (.B1(net1438),
    .Y(_0855_),
    .A1(net534),
    .A2(net1129));
 sg13g2_a21oi_1 _4680_ (.A1(_3091_),
    .A2(net1129),
    .Y(_0168_),
    .B1(_0855_));
 sg13g2_nand2_1 _4681_ (.Y(_0856_),
    .A(_3190_),
    .B(_0750_));
 sg13g2_o21ai_1 _4682_ (.B1(net1429),
    .Y(_0857_),
    .A1(net1414),
    .A2(net1127));
 sg13g2_a21oi_1 _4683_ (.A1(_3100_),
    .A2(net1127),
    .Y(_0169_),
    .B1(_0857_));
 sg13g2_o21ai_1 _4684_ (.B1(net1428),
    .Y(_0858_),
    .A1(net1413),
    .A2(net1127));
 sg13g2_a21oi_1 _4685_ (.A1(_3099_),
    .A2(net1127),
    .Y(_0170_),
    .B1(_0858_));
 sg13g2_o21ai_1 _4686_ (.B1(net1429),
    .Y(_0859_),
    .A1(net1412),
    .A2(net1127));
 sg13g2_a21oi_1 _4687_ (.A1(_3098_),
    .A2(net1126),
    .Y(_0171_),
    .B1(_0859_));
 sg13g2_o21ai_1 _4688_ (.B1(net1429),
    .Y(_0860_),
    .A1(net1411),
    .A2(net1127));
 sg13g2_a21oi_1 _4689_ (.A1(_3097_),
    .A2(net1126),
    .Y(_0172_),
    .B1(_0860_));
 sg13g2_o21ai_1 _4690_ (.B1(net1429),
    .Y(_0861_),
    .A1(net1410),
    .A2(net1126));
 sg13g2_a21oi_1 _4691_ (.A1(_3096_),
    .A2(net1126),
    .Y(_0173_),
    .B1(_0861_));
 sg13g2_o21ai_1 _4692_ (.B1(net1430),
    .Y(_0862_),
    .A1(\dtop.player_inst.synth.alu.acc[5] ),
    .A2(net1126));
 sg13g2_a21oi_1 _4693_ (.A1(_3095_),
    .A2(net1126),
    .Y(_0174_),
    .B1(_0862_));
 sg13g2_o21ai_1 _4694_ (.B1(net1430),
    .Y(_0863_),
    .A1(net1409),
    .A2(net1126));
 sg13g2_a21oi_1 _4695_ (.A1(_3094_),
    .A2(net1126),
    .Y(_0175_),
    .B1(_0863_));
 sg13g2_a22oi_1 _4696_ (.Y(_0864_),
    .B1(net1322),
    .B2(_0838_),
    .A2(_0615_),
    .A1(net1324));
 sg13g2_nand2b_1 _4697_ (.Y(_0865_),
    .B(_0864_),
    .A_N(_0679_));
 sg13g2_a22oi_1 _4698_ (.Y(_0866_),
    .B1(net1317),
    .B2(_3186_),
    .A2(net1325),
    .A1(_0582_));
 sg13g2_nor2_1 _4699_ (.A(net1340),
    .B(_0866_),
    .Y(_0867_));
 sg13g2_and2_1 _4700_ (.A(_0595_),
    .B(net1317),
    .X(_0868_));
 sg13g2_nor2_1 _4701_ (.A(net1335),
    .B(_0633_),
    .Y(_0869_));
 sg13g2_nor4_2 _4702_ (.A(_0652_),
    .B(net1301),
    .C(_0868_),
    .Y(_0870_),
    .D(_0869_));
 sg13g2_o21ai_1 _4703_ (.B1(_0870_),
    .Y(_0871_),
    .A1(net1341),
    .A2(_0866_));
 sg13g2_nor3_1 _4704_ (.A(_0823_),
    .B(_0865_),
    .C(_0871_),
    .Y(_0872_));
 sg13g2_nand2_1 _4705_ (.Y(_0873_),
    .A(_0816_),
    .B(_0872_));
 sg13g2_nand2_1 _4706_ (.Y(_0874_),
    .A(_0778_),
    .B(_0873_));
 sg13g2_inv_1 _4707_ (.Y(_0875_),
    .A(net1125));
 sg13g2_nand2_1 _4708_ (.Y(_0876_),
    .A(net1320),
    .B(_0669_));
 sg13g2_a21oi_1 _4709_ (.A1(net1389),
    .A2(_0662_),
    .Y(_0877_),
    .B1(_0799_));
 sg13g2_a22oi_1 _4710_ (.Y(_0878_),
    .B1(net1318),
    .B2(net1326),
    .A2(_0648_),
    .A1(net1320));
 sg13g2_o21ai_1 _4711_ (.B1(_0650_),
    .Y(_0879_),
    .A1(_0581_),
    .A2(_0654_));
 sg13g2_a221oi_1 _4712_ (.B2(net1316),
    .C1(_0604_),
    .B1(_0640_),
    .A1(_0616_),
    .Y(_0880_),
    .A2(net1322));
 sg13g2_a21oi_1 _4713_ (.A1(net1327),
    .A2(_0838_),
    .Y(_0881_),
    .B1(_0691_));
 sg13g2_and2_1 _4714_ (.A(_0880_),
    .B(_0881_),
    .X(_0882_));
 sg13g2_nand4_1 _4715_ (.B(_0877_),
    .C(_0878_),
    .A(_0876_),
    .Y(_0883_),
    .D(_0882_));
 sg13g2_a21oi_1 _4716_ (.A1(net1322),
    .A2(_0648_),
    .Y(_0884_),
    .B1(_0665_));
 sg13g2_o21ai_1 _4717_ (.B1(_0884_),
    .Y(_0885_),
    .A1(net1349),
    .A2(_0866_));
 sg13g2_nor4_2 _4718_ (.A(_0699_),
    .B(_0867_),
    .C(_0883_),
    .Y(_0886_),
    .D(_0885_));
 sg13g2_a22oi_1 _4719_ (.Y(_0887_),
    .B1(net1316),
    .B2(_0838_),
    .A2(_0669_),
    .A1(net1326));
 sg13g2_nand2_1 _4720_ (.Y(_0888_),
    .A(_0804_),
    .B(_0887_));
 sg13g2_and4_1 _4721_ (.A(_0804_),
    .B(_0825_),
    .C(_0831_),
    .D(_0887_),
    .X(_0889_));
 sg13g2_nor4_2 _4722_ (.A(net1369),
    .B(net1346),
    .C(net1338),
    .Y(_0890_),
    .D(net1331));
 sg13g2_a21oi_1 _4723_ (.A1(_0602_),
    .A2(net1325),
    .Y(_0891_),
    .B1(_0720_));
 sg13g2_nor4_1 _4724_ (.A(_0647_),
    .B(_0666_),
    .C(_0701_),
    .D(_0721_),
    .Y(_0892_));
 sg13g2_nand3b_1 _4725_ (.B(_0891_),
    .C(_0892_),
    .Y(_0893_),
    .A_N(_0890_));
 sg13g2_nand4_1 _4726_ (.B(net1343),
    .C(_0588_),
    .A(net1367),
    .Y(_0894_),
    .D(_0637_));
 sg13g2_nand4_1 _4727_ (.B(net1368),
    .C(_0599_),
    .A(net1380),
    .Y(_0895_),
    .D(_0637_));
 sg13g2_nand3_1 _4728_ (.B(_0894_),
    .C(_0895_),
    .A(_0751_),
    .Y(_0896_));
 sg13g2_or4_1 _4729_ (.A(_0678_),
    .B(_0679_),
    .C(_0837_),
    .D(_0896_),
    .X(_0897_));
 sg13g2_nor3_1 _4730_ (.A(net1347),
    .B(net1336),
    .C(_0677_),
    .Y(_0898_));
 sg13g2_or4_1 _4731_ (.A(_0668_),
    .B(_0681_),
    .C(_0832_),
    .D(_0898_),
    .X(_0899_));
 sg13g2_nor4_2 _4732_ (.A(_0636_),
    .B(_0893_),
    .C(_0897_),
    .Y(_0900_),
    .D(_0899_));
 sg13g2_nand3_1 _4733_ (.B(_0889_),
    .C(_0900_),
    .A(_0886_),
    .Y(_0901_));
 sg13g2_nand3_1 _4734_ (.B(_0686_),
    .C(_0793_),
    .A(_0682_),
    .Y(_0902_));
 sg13g2_nor2_1 _4735_ (.A(_0685_),
    .B(_0692_),
    .Y(_0903_));
 sg13g2_a221oi_1 _4736_ (.B2(_3136_),
    .C1(_0685_),
    .B1(_0662_),
    .A1(net1325),
    .Y(_0904_),
    .A2(net1318));
 sg13g2_o21ai_1 _4737_ (.B1(_0903_),
    .Y(_0905_),
    .A1(_0633_),
    .A2(net1319));
 sg13g2_a22oi_1 _4738_ (.Y(_0906_),
    .B1(net1316),
    .B2(_0648_),
    .A2(net1318),
    .A1(net1320));
 sg13g2_nand4_1 _4739_ (.B(_0802_),
    .C(_0870_),
    .A(_0687_),
    .Y(_0907_),
    .D(_0906_));
 sg13g2_nor3_1 _4740_ (.A(_0902_),
    .B(_0905_),
    .C(_0907_),
    .Y(_0908_));
 sg13g2_nand2_1 _4741_ (.Y(_0909_),
    .A(_0886_),
    .B(_0908_));
 sg13g2_nor2_2 _4742_ (.A(_0694_),
    .B(_0885_),
    .Y(_0910_));
 sg13g2_nand4_1 _4743_ (.B(_0900_),
    .C(_0909_),
    .A(_0889_),
    .Y(_0911_),
    .D(_0910_));
 sg13g2_nand2_1 _4744_ (.Y(_0912_),
    .A(_0901_),
    .B(_0911_));
 sg13g2_nor2b_1 _4745_ (.A(_0694_),
    .B_N(_0908_),
    .Y(_0913_));
 sg13g2_nor2b_1 _4746_ (.A(_0901_),
    .B_N(_0913_),
    .Y(_0914_));
 sg13g2_nor4_2 _4747_ (.A(_0883_),
    .B(_0885_),
    .C(_0905_),
    .Y(_0915_),
    .D(net1224));
 sg13g2_nor2b_1 _4748_ (.A(_0912_),
    .B_N(_0915_),
    .Y(_0916_));
 sg13g2_nor2_2 _4749_ (.A(_0912_),
    .B(_0915_),
    .Y(_0917_));
 sg13g2_nand2_1 _4750_ (.Y(_0918_),
    .A(net1406),
    .B(_0917_));
 sg13g2_nor2_1 _4751_ (.A(_0886_),
    .B(_0911_),
    .Y(_0919_));
 sg13g2_or2_1 _4752_ (.X(_0920_),
    .B(_0915_),
    .A(net1409));
 sg13g2_nand2_1 _4753_ (.Y(_0921_),
    .A(_0919_),
    .B(_0920_));
 sg13g2_a22oi_1 _4754_ (.Y(_0922_),
    .B1(net1152),
    .B2(net1414),
    .A2(_0914_),
    .A1(net1413));
 sg13g2_nand3_1 _4755_ (.B(_0921_),
    .C(_0922_),
    .A(_0918_),
    .Y(_0923_));
 sg13g2_inv_1 _4756_ (.Y(_0924_),
    .A(_0923_));
 sg13g2_a221oi_1 _4757_ (.B2(_0725_),
    .C1(_0014_),
    .B1(net1328),
    .A1(\dtop.detune_counter[17] ),
    .Y(_0925_),
    .A2(_3197_));
 sg13g2_nand3_1 _4758_ (.B(net1345),
    .C(_0727_),
    .A(_3158_),
    .Y(_0926_));
 sg13g2_nor2_2 _4759_ (.A(_3128_),
    .B(_3210_),
    .Y(_0927_));
 sg13g2_nand2_2 _4760_ (.Y(_0928_),
    .A(net1400),
    .B(net1345));
 sg13g2_a21o_1 _4761_ (.A2(_0725_),
    .A1(net1328),
    .B1(_0928_),
    .X(_0929_));
 sg13g2_nor2_1 _4762_ (.A(_0014_),
    .B(_0929_),
    .Y(_0930_));
 sg13g2_nor2_2 _4763_ (.A(_0647_),
    .B(_0890_),
    .Y(_0931_));
 sg13g2_inv_1 _4764_ (.Y(_0932_),
    .A(_0931_));
 sg13g2_nor4_1 _4765_ (.A(_0663_),
    .B(_0693_),
    .C(_0829_),
    .D(_0830_),
    .Y(_0933_));
 sg13g2_nand4_1 _4766_ (.B(_0675_),
    .C(_0817_),
    .A(_0620_),
    .Y(_0934_),
    .D(_0933_));
 sg13g2_nor2_1 _4767_ (.A(_0608_),
    .B(_0934_),
    .Y(_0935_));
 sg13g2_o21ai_1 _4768_ (.B1(net1317),
    .Y(_0936_),
    .A1(_0640_),
    .A2(_0795_));
 sg13g2_o21ai_1 _4769_ (.B1(_3186_),
    .Y(_0937_),
    .A1(net1321),
    .A2(net1317));
 sg13g2_nand3b_1 _4770_ (.B(_0936_),
    .C(_0937_),
    .Y(_0938_),
    .A_N(_0896_));
 sg13g2_o21ai_1 _4771_ (.B1(net1320),
    .Y(_0939_),
    .A1(_0664_),
    .A2(_0818_));
 sg13g2_nor3_1 _4772_ (.A(_0609_),
    .B(_0629_),
    .C(_0667_),
    .Y(_0940_));
 sg13g2_nand4_1 _4773_ (.B(_0683_),
    .C(_0939_),
    .A(net1330),
    .Y(_0941_),
    .D(_0940_));
 sg13g2_nor4_2 _4774_ (.A(_0608_),
    .B(_0934_),
    .C(_0938_),
    .Y(_0942_),
    .D(_0941_));
 sg13g2_or4_2 _4775_ (.A(_0608_),
    .B(_0934_),
    .C(_0938_),
    .D(_0941_),
    .X(_0943_));
 sg13g2_nor3_1 _4776_ (.A(_0888_),
    .B(_0932_),
    .C(_0943_),
    .Y(_0944_));
 sg13g2_nor2_2 _4777_ (.A(net1399),
    .B(_0926_),
    .Y(_0945_));
 sg13g2_nand2_2 _4778_ (.Y(_0946_),
    .A(_3128_),
    .B(_0925_));
 sg13g2_a22oi_1 _4779_ (.Y(_0947_),
    .B1(net1320),
    .B2(_0605_),
    .A2(_0616_),
    .A1(net1326));
 sg13g2_and3_1 _4780_ (.X(_0948_),
    .A(_0931_),
    .B(_0942_),
    .C(_0947_));
 sg13g2_and4_1 _4781_ (.A(_0806_),
    .B(_0931_),
    .C(_0942_),
    .D(_0947_),
    .X(_0949_));
 sg13g2_nor2_1 _4782_ (.A(_0943_),
    .B(_0949_),
    .Y(_0950_));
 sg13g2_and2_1 _4783_ (.A(_0803_),
    .B(_0942_),
    .X(_0951_));
 sg13g2_nand2_1 _4784_ (.Y(_0952_),
    .A(_0803_),
    .B(_0942_));
 sg13g2_a22oi_1 _4785_ (.Y(_0953_),
    .B1(_0945_),
    .B2(_0951_),
    .A2(_0944_),
    .A1(net1281));
 sg13g2_nor2_2 _4786_ (.A(_0925_),
    .B(_0927_),
    .Y(_0954_));
 sg13g2_nand2_2 _4787_ (.Y(_0955_),
    .A(_0926_),
    .B(_0928_));
 sg13g2_nor2_1 _4788_ (.A(_0436_),
    .B(_0943_),
    .Y(_0956_));
 sg13g2_nand2_1 _4789_ (.Y(_0957_),
    .A(_0437_),
    .B(_0942_));
 sg13g2_nor3_1 _4790_ (.A(_0953_),
    .B(_0954_),
    .C(_0957_),
    .Y(_0958_));
 sg13g2_or2_1 _4791_ (.X(_0959_),
    .B(_0958_),
    .A(_0801_));
 sg13g2_inv_2 _4792_ (.Y(_0960_),
    .A(net1171));
 sg13g2_nand4_1 _4793_ (.B(_0686_),
    .C(_0791_),
    .A(_0674_),
    .Y(_0961_),
    .D(_0931_));
 sg13g2_or3_1 _4794_ (.A(_0700_),
    .B(_0805_),
    .C(_0961_),
    .X(_0962_));
 sg13g2_nand4_1 _4795_ (.B(_0887_),
    .C(_0906_),
    .A(_0702_),
    .Y(_0963_),
    .D(_0947_));
 sg13g2_nor2_1 _4796_ (.A(_0962_),
    .B(_0963_),
    .Y(_0964_));
 sg13g2_a221oi_1 _4797_ (.B2(_0627_),
    .C1(_0824_),
    .B1(net1316),
    .A1(net1326),
    .Y(_0965_),
    .A2(_0645_));
 sg13g2_nor2b_1 _4798_ (.A(_0962_),
    .B_N(_0800_),
    .Y(_0966_));
 sg13g2_nor2b_1 _4799_ (.A(_0699_),
    .B_N(_0965_),
    .Y(_0967_));
 sg13g2_nand4_1 _4800_ (.B(_0877_),
    .C(_0939_),
    .A(_0809_),
    .Y(_0968_),
    .D(_0967_));
 sg13g2_nor4_1 _4801_ (.A(_0842_),
    .B(_0938_),
    .C(_0963_),
    .D(_0968_),
    .Y(_0969_));
 sg13g2_a221oi_1 _4802_ (.B2(net1318),
    .C1(_0680_),
    .B1(_0638_),
    .A1(_0615_),
    .Y(_0970_),
    .A2(_0621_));
 sg13g2_nand2_1 _4803_ (.Y(_0971_),
    .A(_0683_),
    .B(_0970_));
 sg13g2_a221oi_1 _4804_ (.B2(net1322),
    .C1(_0821_),
    .B1(_0664_),
    .A1(net1325),
    .Y(_0972_),
    .A2(_0645_));
 sg13g2_nand4_1 _4805_ (.B(_0659_),
    .C(_0671_),
    .A(_0658_),
    .Y(_0973_),
    .D(_0972_));
 sg13g2_nor4_2 _4806_ (.A(_0641_),
    .B(_0754_),
    .C(_0971_),
    .Y(_0974_),
    .D(_0973_));
 sg13g2_nand4_1 _4807_ (.B(_0966_),
    .C(_0969_),
    .A(_0935_),
    .Y(_0975_),
    .D(_0974_));
 sg13g2_nand2_1 _4808_ (.Y(_0976_),
    .A(_0964_),
    .B(_0975_));
 sg13g2_nor3_1 _4809_ (.A(net1349),
    .B(_0943_),
    .C(_0949_),
    .Y(_0977_));
 sg13g2_a21oi_1 _4810_ (.A1(_0804_),
    .A2(_0931_),
    .Y(_0978_),
    .B1(_0943_));
 sg13g2_a22oi_1 _4811_ (.Y(_0979_),
    .B1(_0978_),
    .B2(net1281),
    .A2(_0952_),
    .A1(_0945_));
 sg13g2_o21ai_1 _4812_ (.B1(_0979_),
    .Y(_0980_),
    .A1(_0925_),
    .A2(_0977_));
 sg13g2_a22oi_1 _4813_ (.Y(_0981_),
    .B1(_0980_),
    .B2(_0956_),
    .A2(_0976_),
    .A1(_0943_));
 sg13g2_inv_2 _4814_ (.Y(_0982_),
    .A(_0981_));
 sg13g2_a21oi_2 _4815_ (.B1(_0928_),
    .Y(_0983_),
    .A2(_0727_),
    .A1(_3158_));
 sg13g2_o21ai_1 _4816_ (.B1(_0927_),
    .Y(_0984_),
    .A1(_0014_),
    .A2(_0726_));
 sg13g2_nor2_1 _4817_ (.A(_0978_),
    .B(_0984_),
    .Y(_0985_));
 sg13g2_a21oi_1 _4818_ (.A1(_0947_),
    .A2(_0950_),
    .Y(_0986_),
    .B1(_0946_));
 sg13g2_nor3_1 _4819_ (.A(_0932_),
    .B(_0949_),
    .C(_0955_),
    .Y(_0987_));
 sg13g2_nand3_1 _4820_ (.B(net1281),
    .C(_0942_),
    .A(_0806_),
    .Y(_0988_));
 sg13g2_nor3_1 _4821_ (.A(_0944_),
    .B(_0948_),
    .C(_0988_),
    .Y(_0989_));
 sg13g2_or4_1 _4822_ (.A(_0957_),
    .B(_0985_),
    .C(_0987_),
    .D(_0989_),
    .X(_0990_));
 sg13g2_nand3_1 _4823_ (.B(_0965_),
    .C(_0966_),
    .A(_0943_),
    .Y(_0991_));
 sg13g2_o21ai_1 _4824_ (.B1(_0991_),
    .Y(_0992_),
    .A1(_0986_),
    .A2(_0990_));
 sg13g2_nand3b_1 _4825_ (.B(_0864_),
    .C(_0894_),
    .Y(_0993_),
    .A_N(_0679_));
 sg13g2_a21o_1 _4826_ (.A2(_0673_),
    .A1(net1390),
    .B1(_0665_),
    .X(_0994_));
 sg13g2_nor4_2 _4827_ (.A(_0655_),
    .B(net1301),
    .C(_0993_),
    .Y(_0995_),
    .D(_0994_));
 sg13g2_nor2_2 _4828_ (.A(net1335),
    .B(_0661_),
    .Y(_0996_));
 sg13g2_nand2_1 _4829_ (.Y(_0997_),
    .A(_0659_),
    .B(_0800_));
 sg13g2_nor4_1 _4830_ (.A(_0667_),
    .B(_0868_),
    .C(_0996_),
    .D(_0997_),
    .Y(_0998_));
 sg13g2_o21ai_1 _4831_ (.B1(_0704_),
    .Y(_0999_),
    .A1(net1386),
    .A2(_0866_));
 sg13g2_nand4_1 _4832_ (.B(_0687_),
    .C(_0802_),
    .A(_0682_),
    .Y(_1000_),
    .D(_0906_));
 sg13g2_nor4_2 _4833_ (.A(_0888_),
    .B(_0961_),
    .C(net1279),
    .Y(_1001_),
    .D(_1000_));
 sg13g2_a22oi_1 _4834_ (.Y(_1002_),
    .B1(net1316),
    .B2(_0605_),
    .A2(_0648_),
    .A1(net1324));
 sg13g2_a21oi_1 _4835_ (.A1(net1324),
    .A2(_0616_),
    .Y(_1003_),
    .B1(_0768_));
 sg13g2_nand2_1 _4836_ (.Y(_1004_),
    .A(_1002_),
    .B(_1003_));
 sg13g2_or4_1 _4837_ (.A(_3190_),
    .B(_0619_),
    .C(_0678_),
    .D(_0680_),
    .X(_1005_));
 sg13g2_nor4_2 _4838_ (.A(_0754_),
    .B(_0834_),
    .C(_1004_),
    .Y(_1006_),
    .D(_1005_));
 sg13g2_and2_1 _4839_ (.A(_0751_),
    .B(_0835_),
    .X(_1007_));
 sg13g2_and3_1 _4840_ (.X(_1008_),
    .A(_0751_),
    .B(_0835_),
    .C(_0998_));
 sg13g2_and4_1 _4841_ (.A(_0995_),
    .B(_1001_),
    .C(_1006_),
    .D(_1008_),
    .X(_1009_));
 sg13g2_nand4_1 _4842_ (.B(_1001_),
    .C(_1006_),
    .A(_0995_),
    .Y(_1010_),
    .D(_1008_));
 sg13g2_nor4_1 _4843_ (.A(_0596_),
    .B(_0662_),
    .C(_0663_),
    .D(_0799_),
    .Y(_1011_));
 sg13g2_nand4_1 _4844_ (.B(_0903_),
    .C(_0936_),
    .A(_0607_),
    .Y(_1012_),
    .D(_1011_));
 sg13g2_nand2_1 _4845_ (.Y(_1013_),
    .A(_0642_),
    .B(_0794_));
 sg13g2_nor4_2 _4846_ (.A(_0807_),
    .B(_0879_),
    .C(_1012_),
    .Y(_1014_),
    .D(_1013_));
 sg13g2_nor4_1 _4847_ (.A(_0592_),
    .B(_0668_),
    .C(_0691_),
    .D(_0798_),
    .Y(_1015_));
 sg13g2_and3_1 _4848_ (.X(_1016_),
    .A(_0684_),
    .B(_0696_),
    .C(_1015_));
 sg13g2_nor3_2 _4849_ (.A(_3137_),
    .B(net1338),
    .C(net1334),
    .Y(_1017_));
 sg13g2_inv_1 _4850_ (.Y(_1018_),
    .A(net1314));
 sg13g2_and3_1 _4851_ (.X(_1019_),
    .A(_1014_),
    .B(_1016_),
    .C(_1018_));
 sg13g2_nand3_1 _4852_ (.B(_1016_),
    .C(_1018_),
    .A(_1014_),
    .Y(_1020_));
 sg13g2_nand2b_1 _4853_ (.Y(_1021_),
    .B(_0659_),
    .A_N(net1279));
 sg13g2_nor3_1 _4854_ (.A(_0655_),
    .B(_0993_),
    .C(_1021_),
    .Y(_1022_));
 sg13g2_nand3_1 _4855_ (.B(_1019_),
    .C(_1022_),
    .A(_1010_),
    .Y(_1023_));
 sg13g2_and2_2 _4856_ (.A(_0995_),
    .B(_1014_),
    .X(_1024_));
 sg13g2_nand4_1 _4857_ (.B(_1019_),
    .C(_1022_),
    .A(_1010_),
    .Y(_1025_),
    .D(_1024_));
 sg13g2_a21oi_1 _4858_ (.A1(_0638_),
    .A2(_0640_),
    .Y(_1026_),
    .B1(_0801_));
 sg13g2_nand2_1 _4859_ (.Y(_1027_),
    .A(_0884_),
    .B(_1026_));
 sg13g2_nor4_1 _4860_ (.A(_0993_),
    .B(_0996_),
    .C(net1279),
    .D(_1027_),
    .Y(_1028_));
 sg13g2_nand2_2 _4861_ (.Y(_1029_),
    .A(_1014_),
    .B(_1028_));
 sg13g2_nand4_1 _4862_ (.B(_1014_),
    .C(_1016_),
    .A(_1001_),
    .Y(_1030_),
    .D(_1026_));
 sg13g2_a21oi_2 _4863_ (.B1(_1030_),
    .Y(_1031_),
    .A2(_1019_),
    .A1(_1009_));
 sg13g2_a21o_2 _4864_ (.A2(_1019_),
    .A1(_1009_),
    .B1(_1030_),
    .X(_1032_));
 sg13g2_nand2b_1 _4865_ (.Y(_1033_),
    .B(_1032_),
    .A_N(_1029_));
 sg13g2_nor3_1 _4866_ (.A(_1025_),
    .B(_1029_),
    .C(_1031_),
    .Y(_1034_));
 sg13g2_nor2_1 _4867_ (.A(_0077_),
    .B(net1223),
    .Y(_1035_));
 sg13g2_nor2_1 _4868_ (.A(_0025_),
    .B(net1223),
    .Y(_1036_));
 sg13g2_mux2_1 _4869_ (.A0(_1036_),
    .A1(_1035_),
    .S(net1168),
    .X(_1037_));
 sg13g2_mux2_1 _4870_ (.A0(net1405),
    .A1(\dtop.player_inst.synth.alu.registers[4][0] ),
    .S(net1222),
    .X(_1038_));
 sg13g2_nor2_1 _4871_ (.A(_0023_),
    .B(net1222),
    .Y(_1039_));
 sg13g2_mux2_1 _4872_ (.A0(_1039_),
    .A1(_1038_),
    .S(net1168),
    .X(_1040_));
 sg13g2_mux2_1 _4873_ (.A0(_1037_),
    .A1(_1040_),
    .S(net1170),
    .X(_1041_));
 sg13g2_or2_1 _4874_ (.X(_1042_),
    .B(_1041_),
    .A(net1172));
 sg13g2_nor2b_2 _4875_ (.A(net1170),
    .B_N(net1168),
    .Y(_1043_));
 sg13g2_nor3_2 _4876_ (.A(_3133_),
    .B(\dtop.vtop.rs.saturated ),
    .C(net1223),
    .Y(_1044_));
 sg13g2_nor3_2 _4877_ (.A(_3131_),
    .B(\dtop.vtop.rs.saturated ),
    .C(net1223),
    .Y(_1045_));
 sg13g2_nor3_2 _4878_ (.A(_3132_),
    .B(net1393),
    .C(net1223),
    .Y(_1046_));
 sg13g2_mux2_1 _4879_ (.A0(_1046_),
    .A1(_1045_),
    .S(net1168),
    .X(_1047_));
 sg13g2_a22oi_1 _4880_ (.Y(_1048_),
    .B1(_1047_),
    .B2(net1170),
    .A2(_1044_),
    .A1(_1043_));
 sg13g2_nand2b_1 _4881_ (.Y(_1049_),
    .B(_1030_),
    .A_N(_1025_));
 sg13g2_inv_2 _4882_ (.Y(_1050_),
    .A(net1220));
 sg13g2_a21oi_1 _4883_ (.A1(net1172),
    .A2(_1048_),
    .Y(_1051_),
    .B1(net1219));
 sg13g2_o21ai_1 _4884_ (.B1(_1024_),
    .Y(_1052_),
    .A1(_1010_),
    .A2(_1020_));
 sg13g2_nand2_1 _4885_ (.Y(_1053_),
    .A(_1023_),
    .B(_1052_));
 sg13g2_nand3_1 _4886_ (.B(_1029_),
    .C(_1031_),
    .A(\dtop.player_inst.synth.alu.oct_en ),
    .Y(_1054_));
 sg13g2_or2_1 _4887_ (.X(_1055_),
    .B(_1054_),
    .A(_1053_));
 sg13g2_nor2b_1 _4888_ (.A(net1414),
    .B_N(\dtop.player_inst.synth.alu.carry ),
    .Y(_1056_));
 sg13g2_or2_1 _4889_ (.X(_1057_),
    .B(_1056_),
    .A(_1055_));
 sg13g2_nor3_2 _4890_ (.A(_1029_),
    .B(_1032_),
    .C(_1053_),
    .Y(_1058_));
 sg13g2_nor3_2 _4891_ (.A(net1393),
    .B(net1335),
    .C(_0661_),
    .Y(_1059_));
 sg13g2_nand2_1 _4892_ (.Y(_1060_),
    .A(\dtop.oct_counter[5] ),
    .B(_1059_));
 sg13g2_a22oi_1 _4893_ (.Y(_1061_),
    .B1(net1279),
    .B2(net1446),
    .A2(net1301),
    .A1(\dtop.player_inst.synth.alu.registers[2][0] ));
 sg13g2_nand2b_2 _4894_ (.Y(_1062_),
    .B(_1023_),
    .A_N(_1052_));
 sg13g2_nor2_2 _4895_ (.A(_1033_),
    .B(_1062_),
    .Y(_1063_));
 sg13g2_nor3_2 _4896_ (.A(_1025_),
    .B(_1029_),
    .C(_1032_),
    .Y(_1064_));
 sg13g2_a22oi_1 _4897_ (.Y(_1065_),
    .B1(_1063_),
    .B2(\dtop.player_inst.synth.alu.registers[5][0] ),
    .A2(_1058_),
    .A1(\dtop.player_inst.synth.alu.registers[3][0] ));
 sg13g2_a22oi_1 _4898_ (.Y(_1066_),
    .B1(_1064_),
    .B2(\dtop.player_inst.synth.alu.registers[0][0] ),
    .A2(net1315),
    .A1(\dtop.player_inst.synth.alu.registers[1][0] ));
 sg13g2_and2_1 _4899_ (.A(_1065_),
    .B(_1066_),
    .X(_1067_));
 sg13g2_nand4_1 _4900_ (.B(_1060_),
    .C(_1061_),
    .A(_1057_),
    .Y(_1068_),
    .D(_1067_));
 sg13g2_a21oi_2 _4901_ (.B1(_1068_),
    .Y(_1069_),
    .A2(_1051_),
    .A1(_1042_));
 sg13g2_xnor2_1 _4902_ (.Y(_1070_),
    .A(_0924_),
    .B(_1069_));
 sg13g2_nand3_1 _4903_ (.B(net1431),
    .C(net1125),
    .A(net1414),
    .Y(_1071_));
 sg13g2_o21ai_1 _4904_ (.B1(_1071_),
    .Y(_0176_),
    .A1(net1125),
    .A2(_1070_));
 sg13g2_nand3_1 _4905_ (.B(net1437),
    .C(net1125),
    .A(net1413),
    .Y(_1072_));
 sg13g2_xor2_1 _4906_ (.B(net1406),
    .A(net1414),
    .X(_1073_));
 sg13g2_nand2_1 _4907_ (.Y(_1074_),
    .A(_0905_),
    .B(_1073_));
 sg13g2_nor3_2 _4908_ (.A(_0886_),
    .B(_0911_),
    .C(_0915_),
    .Y(_1075_));
 sg13g2_a22oi_1 _4909_ (.Y(_1076_),
    .B1(_1075_),
    .B2(\dtop.player_inst.synth.alu.acc[7] ),
    .A2(net1224),
    .A1(\dtop.player_inst.synth.alu.acc[2] ));
 sg13g2_a22oi_1 _4910_ (.Y(_1077_),
    .B1(_0917_),
    .B2(\dtop.player_inst.synth.alu.acc[9] ),
    .A2(net1152),
    .A1(net1413));
 sg13g2_nand3_1 _4911_ (.B(_1076_),
    .C(_1077_),
    .A(_1074_),
    .Y(_1078_));
 sg13g2_inv_1 _4912_ (.Y(_1079_),
    .A(_1078_));
 sg13g2_nand3b_1 _4913_ (.B(net1281),
    .C(_0956_),
    .Y(_1080_),
    .A_N(_0887_));
 sg13g2_o21ai_1 _4914_ (.B1(_1080_),
    .Y(_1081_),
    .A1(_0087_),
    .A2(_0910_));
 sg13g2_inv_1 _4915_ (.Y(_1082_),
    .A(net1217));
 sg13g2_mux2_1 _4916_ (.A0(_1035_),
    .A1(_1039_),
    .S(net1168),
    .X(_1083_));
 sg13g2_mux2_1 _4917_ (.A0(net1404),
    .A1(\dtop.player_inst.synth.alu.registers[4][1] ),
    .S(net1222),
    .X(_1084_));
 sg13g2_mux2_1 _4918_ (.A0(_1038_),
    .A1(_1084_),
    .S(net1167),
    .X(_1085_));
 sg13g2_mux4_1 _4919_ (.S0(net1169),
    .A0(_1035_),
    .A1(_1038_),
    .A2(_1039_),
    .A3(_1084_),
    .S1(net1167),
    .X(_1086_));
 sg13g2_mux2_1 _4920_ (.A0(_1045_),
    .A1(_1036_),
    .S(net1168),
    .X(_1087_));
 sg13g2_a221oi_1 _4921_ (.B2(net1170),
    .C1(_0960_),
    .B1(_1087_),
    .A1(_1043_),
    .Y(_1088_),
    .A2(_1046_));
 sg13g2_o21ai_1 _4922_ (.B1(_1050_),
    .Y(_1089_),
    .A1(net1171),
    .A2(_1086_));
 sg13g2_nand2b_1 _4923_ (.Y(_1090_),
    .B(_1056_),
    .A_N(_1055_));
 sg13g2_and2_1 _4924_ (.A(net1425),
    .B(_1059_),
    .X(_1091_));
 sg13g2_a221oi_1 _4925_ (.B2(\dtop.oct_counter[1] ),
    .C1(_1091_),
    .B1(net1279),
    .A1(\dtop.player_inst.synth.alu.registers[2][1] ),
    .Y(_1092_),
    .A2(net1301));
 sg13g2_a22oi_1 _4926_ (.Y(_1093_),
    .B1(_1063_),
    .B2(\dtop.player_inst.synth.alu.registers[5][1] ),
    .A2(_1058_),
    .A1(\dtop.player_inst.synth.alu.registers[3][1] ));
 sg13g2_a22oi_1 _4927_ (.Y(_1094_),
    .B1(_1064_),
    .B2(\dtop.player_inst.synth.alu.registers[0][1] ),
    .A2(net1315),
    .A1(\dtop.player_inst.synth.alu.registers[1][1] ));
 sg13g2_and4_1 _4928_ (.A(_1090_),
    .B(_1092_),
    .C(_1093_),
    .D(_1094_),
    .X(_1095_));
 sg13g2_o21ai_1 _4929_ (.B1(_1095_),
    .Y(_1096_),
    .A1(_1088_),
    .A2(_1089_));
 sg13g2_xnor2_1 _4930_ (.Y(_1097_),
    .A(net1217),
    .B(_1096_));
 sg13g2_nand2b_1 _4931_ (.Y(_1098_),
    .B(_1078_),
    .A_N(_1097_));
 sg13g2_xnor2_1 _4932_ (.Y(_1099_),
    .A(_1079_),
    .B(_1097_));
 sg13g2_mux2_1 _4933_ (.A0(_0924_),
    .A1(_1082_),
    .S(_1069_),
    .X(_1100_));
 sg13g2_a21oi_1 _4934_ (.A1(_1099_),
    .A2(_1100_),
    .Y(_1101_),
    .B1(net1125));
 sg13g2_o21ai_1 _4935_ (.B1(_1101_),
    .Y(_1102_),
    .A1(_1099_),
    .A2(_1100_));
 sg13g2_nand2_1 _4936_ (.Y(_0177_),
    .A(_1072_),
    .B(_1102_));
 sg13g2_nand3_1 _4937_ (.B(net1437),
    .C(net1124),
    .A(net1412),
    .Y(_1103_));
 sg13g2_o21ai_1 _4938_ (.B1(_1098_),
    .Y(_1104_),
    .A1(_1099_),
    .A2(_1100_));
 sg13g2_nand2_1 _4939_ (.Y(_1105_),
    .A(\dtop.player_inst.synth.alu.acc[8] ),
    .B(_0901_));
 sg13g2_xnor2_1 _4940_ (.Y(_1106_),
    .A(net1413),
    .B(net1407));
 sg13g2_nor2_1 _4941_ (.A(_0904_),
    .B(_1106_),
    .Y(_1107_));
 sg13g2_a221oi_1 _4942_ (.B2(net1412),
    .C1(_1107_),
    .B1(net1152),
    .A1(net1411),
    .Y(_1108_),
    .A2(net1224));
 sg13g2_o21ai_1 _4943_ (.B1(_1108_),
    .Y(_1109_),
    .A1(_0915_),
    .A2(_1105_));
 sg13g2_nand2_1 _4944_ (.Y(_1110_),
    .A(net1170),
    .B(_1037_));
 sg13g2_nand2_1 _4945_ (.Y(_1111_),
    .A(_0982_),
    .B(_1047_));
 sg13g2_nand3_1 _4946_ (.B(_1110_),
    .C(_1111_),
    .A(net1172),
    .Y(_1112_));
 sg13g2_mux2_1 _4947_ (.A0(net1402),
    .A1(\dtop.player_inst.synth.alu.registers[4][2] ),
    .S(net1222),
    .X(_1113_));
 sg13g2_mux2_1 _4948_ (.A0(_1084_),
    .A1(_1113_),
    .S(net1166),
    .X(_1114_));
 sg13g2_mux4_1 _4949_ (.S0(net1169),
    .A0(_1039_),
    .A1(_1084_),
    .A2(_1038_),
    .A3(_1113_),
    .S1(net1167),
    .X(_1115_));
 sg13g2_nor2_1 _4950_ (.A(net1172),
    .B(_1115_),
    .Y(_1116_));
 sg13g2_nor2_1 _4951_ (.A(net1219),
    .B(_1116_),
    .Y(_1117_));
 sg13g2_a22oi_1 _4952_ (.Y(_1118_),
    .B1(_1063_),
    .B2(\dtop.player_inst.synth.alu.registers[5][2] ),
    .A2(net1314),
    .A1(\dtop.player_inst.synth.alu.registers[1][2] ));
 sg13g2_a22oi_1 _4953_ (.Y(_1119_),
    .B1(net1218),
    .B2(\dtop.player_inst.synth.alu.registers[0][2] ),
    .A2(_1058_),
    .A1(\dtop.player_inst.synth.alu.registers[3][2] ));
 sg13g2_a22oi_1 _4954_ (.Y(_1120_),
    .B1(net1279),
    .B2(\dtop.oct_counter[2] ),
    .A2(net1301),
    .A1(\dtop.player_inst.synth.alu.registers[2][2] ));
 sg13g2_nand3_1 _4955_ (.B(_1119_),
    .C(_1120_),
    .A(_1118_),
    .Y(_1121_));
 sg13g2_a221oi_1 _4956_ (.B2(_1117_),
    .C1(_1121_),
    .B1(_1112_),
    .A1(net1424),
    .Y(_1122_),
    .A2(_1059_));
 sg13g2_xnor2_1 _4957_ (.Y(_1123_),
    .A(net1217),
    .B(_1122_));
 sg13g2_and2_1 _4958_ (.A(_1109_),
    .B(_1123_),
    .X(_1124_));
 sg13g2_xor2_1 _4959_ (.B(_1123_),
    .A(_1109_),
    .X(_1125_));
 sg13g2_and2_1 _4960_ (.A(_1104_),
    .B(_1125_),
    .X(_1126_));
 sg13g2_o21ai_1 _4961_ (.B1(net1111),
    .Y(_1127_),
    .A1(_1104_),
    .A2(_1125_));
 sg13g2_o21ai_1 _4962_ (.B1(_1103_),
    .Y(_0178_),
    .A1(_1126_),
    .A2(_1127_));
 sg13g2_nand3_1 _4963_ (.B(net1437),
    .C(net1124),
    .A(net1411),
    .Y(_1128_));
 sg13g2_a21oi_1 _4964_ (.A1(_1104_),
    .A2(_1125_),
    .Y(_1129_),
    .B1(_1124_));
 sg13g2_nand2_1 _4965_ (.Y(_1130_),
    .A(\dtop.player_inst.synth.alu.acc[9] ),
    .B(_1075_));
 sg13g2_xor2_1 _4966_ (.B(net1406),
    .A(net1412),
    .X(_1131_));
 sg13g2_a22oi_1 _4967_ (.Y(_1132_),
    .B1(_1131_),
    .B2(_0905_),
    .A2(net1224),
    .A1(\dtop.player_inst.synth.alu.acc[4] ));
 sg13g2_a22oi_1 _4968_ (.Y(_1133_),
    .B1(_0917_),
    .B2(net1408),
    .A2(net1152),
    .A1(net1411));
 sg13g2_nand3_1 _4969_ (.B(_1132_),
    .C(_1133_),
    .A(_1130_),
    .Y(_1134_));
 sg13g2_nor2_2 _4970_ (.A(_1023_),
    .B(_1024_),
    .Y(_1135_));
 sg13g2_a221oi_1 _4971_ (.B2(_3126_),
    .C1(_3213_),
    .B1(net1300),
    .A1(_3158_),
    .Y(_1136_),
    .A2(_3210_));
 sg13g2_inv_1 _4972_ (.Y(_1137_),
    .A(_1136_));
 sg13g2_nor3_2 _4973_ (.A(_1023_),
    .B(_1024_),
    .C(_1137_),
    .Y(_1138_));
 sg13g2_a221oi_1 _4974_ (.B2(_0731_),
    .C1(_0736_),
    .B1(_0730_),
    .A1(net1328),
    .Y(_1139_),
    .A2(_0725_));
 sg13g2_and3_1 _4975_ (.X(_1140_),
    .A(net1399),
    .B(_0925_),
    .C(_1139_));
 sg13g2_and2_1 _4976_ (.A(_3159_),
    .B(_1140_),
    .X(_1141_));
 sg13g2_nor2_1 _4977_ (.A(net1404),
    .B(\dtop.detune_counter[7] ),
    .Y(_1142_));
 sg13g2_and2_1 _4978_ (.A(_1139_),
    .B(_1142_),
    .X(_1143_));
 sg13g2_nand2b_1 _4979_ (.Y(_1144_),
    .B(net1345),
    .A_N(_0016_));
 sg13g2_nor3_1 _4980_ (.A(_0018_),
    .B(_0020_),
    .C(_1144_),
    .Y(_1145_));
 sg13g2_o21ai_1 _4981_ (.B1(_1145_),
    .Y(_1146_),
    .A1(_0733_),
    .A2(_0929_));
 sg13g2_nand3b_1 _4982_ (.B(_0020_),
    .C(net1345),
    .Y(_1147_),
    .A_N(_0018_));
 sg13g2_nor2_1 _4983_ (.A(_0016_),
    .B(_1147_),
    .Y(_1148_));
 sg13g2_a221oi_1 _4984_ (.B2(\dtop.detune_counter[17] ),
    .C1(_0016_),
    .B1(_3197_),
    .A1(_0018_),
    .Y(_1149_),
    .A2(_3159_));
 sg13g2_a21oi_1 _4985_ (.A1(_1144_),
    .A2(_1147_),
    .Y(_1150_),
    .B1(_1149_));
 sg13g2_a21oi_1 _4986_ (.A1(_0734_),
    .A2(_1148_),
    .Y(_1151_),
    .B1(_1150_));
 sg13g2_a221oi_1 _4987_ (.B2(_1151_),
    .C1(_1143_),
    .B1(_1146_),
    .A1(net1280),
    .Y(_1152_),
    .A2(_1139_));
 sg13g2_nor2_1 _4988_ (.A(_1141_),
    .B(_1152_),
    .Y(_1153_));
 sg13g2_or2_1 _4989_ (.X(_1154_),
    .B(_1152_),
    .A(_1141_));
 sg13g2_and2_1 _4990_ (.A(_0954_),
    .B(_1143_),
    .X(_1155_));
 sg13g2_nand2_1 _4991_ (.Y(_1156_),
    .A(_0954_),
    .B(_1143_));
 sg13g2_or3_1 _4992_ (.A(_1140_),
    .B(_1143_),
    .C(_1148_),
    .X(_1157_));
 sg13g2_nand2_1 _4993_ (.Y(_1158_),
    .A(_0732_),
    .B(net1280));
 sg13g2_nand4_1 _4994_ (.B(_0732_),
    .C(_0927_),
    .A(_0727_),
    .Y(_1159_),
    .D(_1145_));
 sg13g2_and4_1 _4995_ (.A(_0016_),
    .B(_0018_),
    .C(_3159_),
    .D(net1344),
    .X(_1160_));
 sg13g2_o21ai_1 _4996_ (.B1(_0018_),
    .Y(_1161_),
    .A1(_1149_),
    .A2(_1160_));
 sg13g2_nand2_1 _4997_ (.Y(_1162_),
    .A(_1159_),
    .B(_1161_));
 sg13g2_a21oi_2 _4998_ (.B1(_1162_),
    .Y(_1163_),
    .A2(_1158_),
    .A1(_1157_));
 sg13g2_a21o_1 _4999_ (.A2(_1158_),
    .A1(_1157_),
    .B1(_1162_),
    .X(_1164_));
 sg13g2_nor2_1 _5000_ (.A(_1155_),
    .B(_1163_),
    .Y(_1165_));
 sg13g2_nand2_1 _5001_ (.Y(_1166_),
    .A(_1156_),
    .B(_1164_));
 sg13g2_a21oi_1 _5002_ (.A1(_1156_),
    .A2(_1164_),
    .Y(_1167_),
    .B1(_1154_));
 sg13g2_o21ai_1 _5003_ (.B1(_1153_),
    .Y(_1168_),
    .A1(_1155_),
    .A2(_1163_));
 sg13g2_nor2_1 _5004_ (.A(_0733_),
    .B(_1168_),
    .Y(_1169_));
 sg13g2_o21ai_1 _5005_ (.B1(_1154_),
    .Y(_1170_),
    .A1(_1155_),
    .A2(_1163_));
 sg13g2_nand3_1 _5006_ (.B(_1156_),
    .C(_1164_),
    .A(_1154_),
    .Y(_1171_));
 sg13g2_a22oi_1 _5007_ (.Y(_1172_),
    .B1(_1171_),
    .B2(net1280),
    .A2(_1170_),
    .A1(_0945_));
 sg13g2_nor2_1 _5008_ (.A(_0955_),
    .B(_1153_),
    .Y(_1173_));
 sg13g2_nor2_1 _5009_ (.A(net1300),
    .B(_0955_),
    .Y(_1174_));
 sg13g2_nand2_1 _5010_ (.Y(_1175_),
    .A(_0733_),
    .B(_0954_));
 sg13g2_nor2b_2 _5011_ (.A(net1402),
    .B_N(net1401),
    .Y(_1176_));
 sg13g2_nand2_1 _5012_ (.Y(_1177_),
    .A(_0726_),
    .B(_1176_));
 sg13g2_nand3_1 _5013_ (.B(_0733_),
    .C(_1176_),
    .A(_0726_),
    .Y(_1178_));
 sg13g2_a21oi_1 _5014_ (.A1(_1153_),
    .A2(_1178_),
    .Y(_1179_),
    .B1(_0984_));
 sg13g2_a221oi_1 _5015_ (.B2(_1168_),
    .C1(_1173_),
    .B1(_1179_),
    .A1(_1166_),
    .Y(_1180_),
    .A2(_1174_));
 sg13g2_o21ai_1 _5016_ (.B1(_1180_),
    .Y(_1181_),
    .A1(_1169_),
    .A2(_1172_));
 sg13g2_o21ai_1 _5017_ (.B1(net1403),
    .Y(_1182_),
    .A1(net1401),
    .A2(net1402));
 sg13g2_o21ai_1 _5018_ (.B1(_3130_),
    .Y(_1183_),
    .A1(_0735_),
    .A2(_1182_));
 sg13g2_nor3_1 _5019_ (.A(\dtop.detune_counter[10] ),
    .B(net1404),
    .C(\dtop.detune_counter[9] ),
    .Y(_1184_));
 sg13g2_nand2b_1 _5020_ (.Y(_1185_),
    .B(net1405),
    .A_N(_1184_));
 sg13g2_and2_1 _5021_ (.A(_1183_),
    .B(_1185_),
    .X(_1186_));
 sg13g2_nor2_1 _5022_ (.A(net1403),
    .B(_3130_),
    .Y(_1187_));
 sg13g2_a21oi_2 _5023_ (.B1(_1186_),
    .Y(_1188_),
    .A2(_1187_),
    .A1(_0735_));
 sg13g2_a21oi_1 _5024_ (.A1(_3128_),
    .A2(_0730_),
    .Y(_1189_),
    .B1(_0983_));
 sg13g2_nand2b_1 _5025_ (.Y(_1190_),
    .B(_1188_),
    .A_N(_1189_));
 sg13g2_nor3_2 _5026_ (.A(\dtop.detune_counter[14] ),
    .B(\dtop.detune_counter[17] ),
    .C(_3281_),
    .Y(_1191_));
 sg13g2_nand2_2 _5027_ (.Y(_1192_),
    .A(_3126_),
    .B(_3282_));
 sg13g2_nand2_1 _5028_ (.Y(_1193_),
    .A(_1183_),
    .B(_1188_));
 sg13g2_a21oi_1 _5029_ (.A1(_1183_),
    .A2(_1188_),
    .Y(_1194_),
    .B1(_1192_));
 sg13g2_nor3_1 _5030_ (.A(_0014_),
    .B(_0929_),
    .C(_1186_),
    .Y(_1195_));
 sg13g2_nand2_1 _5031_ (.Y(_1196_),
    .A(_3129_),
    .B(net1405));
 sg13g2_and2_1 _5032_ (.A(_1182_),
    .B(_1196_),
    .X(_1197_));
 sg13g2_nand2_2 _5033_ (.Y(_1198_),
    .A(net1403),
    .B(_3130_));
 sg13g2_nor3_1 _5034_ (.A(_3128_),
    .B(_0736_),
    .C(_1198_),
    .Y(_1199_));
 sg13g2_nor3_1 _5035_ (.A(net1280),
    .B(_1197_),
    .C(_1199_),
    .Y(_1200_));
 sg13g2_nor3_1 _5036_ (.A(_3321_),
    .B(_1195_),
    .C(_1200_),
    .Y(_1201_));
 sg13g2_a21oi_1 _5037_ (.A1(net1403),
    .A2(_3130_),
    .Y(_1202_),
    .B1(_3322_));
 sg13g2_nor3_1 _5038_ (.A(_3321_),
    .B(_1193_),
    .C(_1197_),
    .Y(_1203_));
 sg13g2_nor2_1 _5039_ (.A(_3130_),
    .B(_1176_),
    .Y(_1204_));
 sg13g2_nor2_1 _5040_ (.A(net1403),
    .B(_1204_),
    .Y(_1205_));
 sg13g2_nand2_1 _5041_ (.Y(_1206_),
    .A(_1189_),
    .B(_1205_));
 sg13g2_nor4_1 _5042_ (.A(_3321_),
    .B(_1189_),
    .C(_1195_),
    .D(_1200_),
    .Y(_1207_));
 sg13g2_o21ai_1 _5043_ (.B1(_1206_),
    .Y(_1208_),
    .A1(_1202_),
    .A2(_1207_));
 sg13g2_nor2_1 _5044_ (.A(_1191_),
    .B(_1203_),
    .Y(_1209_));
 sg13g2_a22oi_1 _5045_ (.Y(_1210_),
    .B1(_1208_),
    .B2(_1209_),
    .A2(_1194_),
    .A1(_1190_));
 sg13g2_nor2_1 _5046_ (.A(_1062_),
    .B(_1210_),
    .Y(_1211_));
 sg13g2_nor2_1 _5047_ (.A(\dtop.detune_counter[12] ),
    .B(net1400),
    .Y(_1212_));
 sg13g2_o21ai_1 _5048_ (.B1(_1184_),
    .Y(_1213_),
    .A1(net1344),
    .A2(_1212_));
 sg13g2_nand2b_1 _5049_ (.Y(_1214_),
    .B(_1213_),
    .A_N(_3213_));
 sg13g2_inv_1 _5050_ (.Y(_1215_),
    .A(_1214_));
 sg13g2_o21ai_1 _5051_ (.B1(_1215_),
    .Y(_1216_),
    .A1(_1023_),
    .A2(_1024_));
 sg13g2_nor2b_2 _5052_ (.A(_1216_),
    .B_N(_1062_),
    .Y(_1217_));
 sg13g2_nor2_1 _5053_ (.A(_0945_),
    .B(_0983_),
    .Y(_1218_));
 sg13g2_nand2_1 _5054_ (.Y(_1219_),
    .A(_0436_),
    .B(net1280));
 sg13g2_nand3_1 _5055_ (.B(_1218_),
    .C(_1219_),
    .A(_1175_),
    .Y(_1220_));
 sg13g2_a22oi_1 _5056_ (.Y(_1221_),
    .B1(_1217_),
    .B2(_1220_),
    .A2(_1181_),
    .A1(_1138_));
 sg13g2_a221oi_1 _5057_ (.B2(_1220_),
    .C1(_1211_),
    .B1(_1217_),
    .A1(_1138_),
    .Y(_1222_),
    .A2(_1181_));
 sg13g2_nand2b_1 _5058_ (.Y(_1223_),
    .B(_1221_),
    .A_N(_1211_));
 sg13g2_nor2_1 _5059_ (.A(_0946_),
    .B(_1168_),
    .Y(_1224_));
 sg13g2_nor3_2 _5060_ (.A(_1154_),
    .B(_1155_),
    .C(_1163_),
    .Y(_1225_));
 sg13g2_or2_1 _5061_ (.X(_1226_),
    .B(_1225_),
    .A(_1218_));
 sg13g2_a21oi_1 _5062_ (.A1(_0925_),
    .A2(_1165_),
    .Y(_1227_),
    .B1(_1173_));
 sg13g2_a21o_1 _5063_ (.A2(_1227_),
    .A1(_1226_),
    .B1(_1224_),
    .X(_1228_));
 sg13g2_nand2_1 _5064_ (.Y(_1229_),
    .A(_0955_),
    .B(_1219_));
 sg13g2_a21oi_1 _5065_ (.A1(net1280),
    .A2(_1198_),
    .Y(_1230_),
    .B1(_3322_));
 sg13g2_o21ai_1 _5066_ (.B1(_1230_),
    .Y(_1231_),
    .A1(net1280),
    .A2(_1205_));
 sg13g2_nor2_1 _5067_ (.A(_1191_),
    .B(_1201_),
    .Y(_1232_));
 sg13g2_mux2_1 _5068_ (.A0(_1183_),
    .A1(_1188_),
    .S(net1280),
    .X(_1233_));
 sg13g2_a221oi_1 _5069_ (.B2(_1191_),
    .C1(_1062_),
    .B1(_1233_),
    .A1(_1231_),
    .Y(_1234_),
    .A2(_1232_));
 sg13g2_a221oi_1 _5070_ (.B2(_1217_),
    .C1(_1234_),
    .B1(_1229_),
    .A1(_1138_),
    .Y(_1235_),
    .A2(_1228_));
 sg13g2_a221oi_1 _5071_ (.B2(_1225_),
    .C1(_0984_),
    .B1(_1177_),
    .A1(_0726_),
    .Y(_1236_),
    .A2(_1167_));
 sg13g2_o21ai_1 _5072_ (.B1(_0925_),
    .Y(_1237_),
    .A1(net1399),
    .A2(_1164_));
 sg13g2_nor2_1 _5073_ (.A(_1225_),
    .B(_1237_),
    .Y(_1238_));
 sg13g2_and2_1 _5074_ (.A(_0954_),
    .B(_1171_),
    .X(_1239_));
 sg13g2_or4_1 _5075_ (.A(_1224_),
    .B(_1236_),
    .C(_1238_),
    .D(_1239_),
    .X(_1240_));
 sg13g2_nand2_1 _5076_ (.Y(_1241_),
    .A(_0925_),
    .B(_1219_));
 sg13g2_a21oi_1 _5077_ (.A1(_3210_),
    .A2(_1205_),
    .Y(_1242_),
    .B1(_3322_));
 sg13g2_o21ai_1 _5078_ (.B1(_1242_),
    .Y(_1243_),
    .A1(_0945_),
    .A2(_1198_));
 sg13g2_nand2_1 _5079_ (.Y(_1244_),
    .A(_0928_),
    .B(_1197_));
 sg13g2_nand2_1 _5080_ (.Y(_1245_),
    .A(_3322_),
    .B(_1244_));
 sg13g2_a21oi_1 _5081_ (.A1(net1399),
    .A2(_1186_),
    .Y(_1246_),
    .B1(_1245_));
 sg13g2_a21oi_1 _5082_ (.A1(_0955_),
    .A2(_1246_),
    .Y(_1247_),
    .B1(_1203_));
 sg13g2_nand2_1 _5083_ (.Y(_1248_),
    .A(_1243_),
    .B(_1247_));
 sg13g2_nor2_1 _5084_ (.A(_0927_),
    .B(_1183_),
    .Y(_1249_));
 sg13g2_nor2_1 _5085_ (.A(_1192_),
    .B(_1249_),
    .Y(_1250_));
 sg13g2_or2_1 _5086_ (.X(_1251_),
    .B(_1188_),
    .A(_0945_));
 sg13g2_a221oi_1 _5087_ (.B2(_1251_),
    .C1(_1062_),
    .B1(_1250_),
    .A1(_1192_),
    .Y(_1252_),
    .A2(_1248_));
 sg13g2_a221oi_1 _5088_ (.B2(_1217_),
    .C1(_1252_),
    .B1(_1241_),
    .A1(_1138_),
    .Y(_1253_),
    .A2(_1240_));
 sg13g2_or3_2 _5089_ (.A(net1300),
    .B(_1235_),
    .C(_1253_),
    .X(_1254_));
 sg13g2_o21ai_1 _5090_ (.B1(_1253_),
    .Y(_1255_),
    .A1(net1300),
    .A2(_1235_));
 sg13g2_and2_1 _5091_ (.A(_1254_),
    .B(_1255_),
    .X(_1256_));
 sg13g2_nand2_1 _5092_ (.Y(_1257_),
    .A(_1254_),
    .B(_1255_));
 sg13g2_nand3_1 _5093_ (.B(_1254_),
    .C(_1255_),
    .A(_1222_),
    .Y(_1258_));
 sg13g2_xnor2_1 _5094_ (.Y(_1259_),
    .A(_0733_),
    .B(_1235_));
 sg13g2_a21oi_2 _5095_ (.B1(_1259_),
    .Y(_1260_),
    .A2(_1255_),
    .A1(_1254_));
 sg13g2_nor4_2 _5096_ (.A(net1300),
    .B(_1222_),
    .C(_1235_),
    .Y(_1261_),
    .D(_1253_));
 sg13g2_xnor2_1 _5097_ (.Y(_1262_),
    .A(_1223_),
    .B(_1254_));
 sg13g2_nand2_1 _5098_ (.Y(_1263_),
    .A(_1260_),
    .B(_1262_));
 sg13g2_nor2b_1 _5099_ (.A(_1177_),
    .B_N(_1225_),
    .Y(_1264_));
 sg13g2_nor2_1 _5100_ (.A(_1167_),
    .B(_1264_),
    .Y(_1265_));
 sg13g2_o21ai_1 _5101_ (.B1(_1265_),
    .Y(_1266_),
    .A1(_0946_),
    .A2(_1165_));
 sg13g2_nor3_1 _5102_ (.A(_0000_),
    .B(_0736_),
    .C(_1198_),
    .Y(_1267_));
 sg13g2_a21oi_1 _5103_ (.A1(_0928_),
    .A2(_1267_),
    .Y(_1268_),
    .B1(_1245_));
 sg13g2_nor2_1 _5104_ (.A(_1242_),
    .B(_1268_),
    .Y(_1269_));
 sg13g2_nor2_1 _5105_ (.A(_1191_),
    .B(_1269_),
    .Y(_1270_));
 sg13g2_nor3_1 _5106_ (.A(_1062_),
    .B(_1250_),
    .C(_1270_),
    .Y(_1271_));
 sg13g2_a221oi_1 _5107_ (.B2(_1138_),
    .C1(_1271_),
    .B1(_1266_),
    .A1(_0954_),
    .Y(_1272_),
    .A2(_1217_));
 sg13g2_xor2_1 _5108_ (.B(_1272_),
    .A(_1261_),
    .X(_1273_));
 sg13g2_xnor2_1 _5109_ (.Y(_1274_),
    .A(_1261_),
    .B(_1272_));
 sg13g2_a221oi_1 _5110_ (.B2(_1262_),
    .C1(_1274_),
    .B1(_1260_),
    .A1(_1222_),
    .Y(_1275_),
    .A2(_1256_));
 sg13g2_nand3_1 _5111_ (.B(_1031_),
    .C(_1135_),
    .A(_1029_),
    .Y(_1276_));
 sg13g2_o21ai_1 _5112_ (.B1(_0659_),
    .Y(_1277_),
    .A1(_1033_),
    .A2(_1053_));
 sg13g2_nand2b_2 _5113_ (.Y(_1278_),
    .B(_1276_),
    .A_N(_1277_));
 sg13g2_o21ai_1 _5114_ (.B1(_1278_),
    .Y(_1279_),
    .A1(_1260_),
    .A2(_1273_));
 sg13g2_nand2_1 _5115_ (.Y(_1280_),
    .A(\dtop.oct_counter[3] ),
    .B(_0999_));
 sg13g2_nand2_1 _5116_ (.Y(_1281_),
    .A(\dtop.player_inst.synth.alu.registers[1][3] ),
    .B(net1314));
 sg13g2_a22oi_1 _5117_ (.Y(_1282_),
    .B1(_1059_),
    .B2(net1418),
    .A2(net1301),
    .A1(\dtop.player_inst.synth.alu.registers[2][3] ));
 sg13g2_nand4_1 _5118_ (.B(_1280_),
    .C(_1281_),
    .A(net1220),
    .Y(_1283_),
    .D(_1282_));
 sg13g2_a21o_1 _5119_ (.A2(_1063_),
    .A1(\dtop.player_inst.synth.alu.registers[5][3] ),
    .B1(_1283_),
    .X(_1284_));
 sg13g2_a221oi_1 _5120_ (.B2(\dtop.player_inst.synth.alu.registers[0][3] ),
    .C1(_1284_),
    .B1(net1218),
    .A1(\dtop.player_inst.synth.alu.registers[3][3] ),
    .Y(_1285_),
    .A2(_1058_));
 sg13g2_o21ai_1 _5121_ (.B1(_1285_),
    .Y(_1286_),
    .A1(_1275_),
    .A2(_1279_));
 sg13g2_nor2_1 _5122_ (.A(\dtop.detune_counter[10] ),
    .B(net1222),
    .Y(_1287_));
 sg13g2_a21oi_1 _5123_ (.A1(_3116_),
    .A2(net1222),
    .Y(_1288_),
    .B1(_1287_));
 sg13g2_mux2_1 _5124_ (.A0(_1113_),
    .A1(_1288_),
    .S(net1166),
    .X(_1289_));
 sg13g2_mux4_1 _5125_ (.S0(_0982_),
    .A0(_1083_),
    .A1(_1087_),
    .A2(_1289_),
    .A3(_1085_),
    .S1(_0960_),
    .X(_1290_));
 sg13g2_nand2b_1 _5126_ (.Y(_1291_),
    .B(_1050_),
    .A_N(_1290_));
 sg13g2_nand2_1 _5127_ (.Y(_1292_),
    .A(_1286_),
    .B(_1291_));
 sg13g2_nand3_1 _5128_ (.B(_1286_),
    .C(_1291_),
    .A(net1217),
    .Y(_1293_));
 sg13g2_a21o_1 _5129_ (.A2(_1291_),
    .A1(_1286_),
    .B1(net1217),
    .X(_1294_));
 sg13g2_nand2_1 _5130_ (.Y(_1295_),
    .A(_1293_),
    .B(_1294_));
 sg13g2_nand3_1 _5131_ (.B(_1293_),
    .C(_1294_),
    .A(_1134_),
    .Y(_1296_));
 sg13g2_a21oi_1 _5132_ (.A1(_1293_),
    .A2(_1294_),
    .Y(_1297_),
    .B1(_1134_));
 sg13g2_xor2_1 _5133_ (.B(_1295_),
    .A(_1134_),
    .X(_1298_));
 sg13g2_nor2_1 _5134_ (.A(_1129_),
    .B(_1298_),
    .Y(_1299_));
 sg13g2_a21o_1 _5135_ (.A2(_1298_),
    .A1(_1129_),
    .B1(net1125),
    .X(_1300_));
 sg13g2_o21ai_1 _5136_ (.B1(_1128_),
    .Y(_0179_),
    .A1(_1299_),
    .A2(_1300_));
 sg13g2_nand3_1 _5137_ (.B(net1437),
    .C(net1124),
    .A(net1410),
    .Y(_1301_));
 sg13g2_o21ai_1 _5138_ (.B1(_1296_),
    .Y(_1302_),
    .A1(_1129_),
    .A2(_1297_));
 sg13g2_xor2_1 _5139_ (.B(net1406),
    .A(net1411),
    .X(_1303_));
 sg13g2_nand2_1 _5140_ (.Y(_1304_),
    .A(\dtop.player_inst.synth.alu.acc[5] ),
    .B(net1224));
 sg13g2_a22oi_1 _5141_ (.Y(_1305_),
    .B1(_1303_),
    .B2(_0905_),
    .A2(_0917_),
    .A1(net1409));
 sg13g2_a22oi_1 _5142_ (.Y(_1306_),
    .B1(_1075_),
    .B2(_0063_),
    .A2(net1152),
    .A1(net1410));
 sg13g2_nand3_1 _5143_ (.B(_1305_),
    .C(_1306_),
    .A(_1304_),
    .Y(_1307_));
 sg13g2_nand2_1 _5144_ (.Y(_1308_),
    .A(net1172),
    .B(_1041_));
 sg13g2_nand2_1 _5145_ (.Y(_1309_),
    .A(\dtop.player_inst.synth.alu.registers[4][4] ),
    .B(net1221));
 sg13g2_o21ai_1 _5146_ (.B1(_1309_),
    .Y(_1310_),
    .A1(_3128_),
    .A2(net1222));
 sg13g2_mux2_1 _5147_ (.A0(_1288_),
    .A1(_1310_),
    .S(net1167),
    .X(_1311_));
 sg13g2_mux2_1 _5148_ (.A0(_1114_),
    .A1(_1311_),
    .S(net1169),
    .X(_1312_));
 sg13g2_a21oi_1 _5149_ (.A1(_0960_),
    .A2(_1312_),
    .Y(_1313_),
    .B1(net1220));
 sg13g2_nand3_1 _5150_ (.B(_1259_),
    .C(_1273_),
    .A(_1258_),
    .Y(_1314_));
 sg13g2_nand2_1 _5151_ (.Y(_1315_),
    .A(_1278_),
    .B(_1314_));
 sg13g2_nand2_1 _5152_ (.Y(_1316_),
    .A(\dtop.player_inst.synth.alu.registers[5][4] ),
    .B(_1063_));
 sg13g2_a22oi_1 _5153_ (.Y(_1317_),
    .B1(net1314),
    .B2(\dtop.player_inst.synth.alu.registers[1][4] ),
    .A2(net1301),
    .A1(\dtop.player_inst.synth.alu.registers[2][4] ));
 sg13g2_inv_1 _5154_ (.Y(_1318_),
    .A(_1317_));
 sg13g2_a221oi_1 _5155_ (.B2(\dtop.vtop.logo.addr[9] ),
    .C1(_1318_),
    .B1(_1059_),
    .A1(\dtop.oct_counter[4] ),
    .Y(_1319_),
    .A2(_0999_));
 sg13g2_nand3_1 _5156_ (.B(_1316_),
    .C(_1319_),
    .A(net1220),
    .Y(_1320_));
 sg13g2_a221oi_1 _5157_ (.B2(\dtop.player_inst.synth.alu.registers[0][4] ),
    .C1(_1320_),
    .B1(net1218),
    .A1(\dtop.player_inst.synth.alu.registers[3][4] ),
    .Y(_1321_),
    .A2(_1058_));
 sg13g2_a22oi_1 _5158_ (.Y(_1322_),
    .B1(_1315_),
    .B2(_1321_),
    .A2(_1313_),
    .A1(_1308_));
 sg13g2_xnor2_1 _5159_ (.Y(_1323_),
    .A(net1217),
    .B(_1322_));
 sg13g2_nor2b_1 _5160_ (.A(_1323_),
    .B_N(_1307_),
    .Y(_1324_));
 sg13g2_xnor2_1 _5161_ (.Y(_1325_),
    .A(_1307_),
    .B(_1323_));
 sg13g2_o21ai_1 _5162_ (.B1(net1111),
    .Y(_1326_),
    .A1(_1302_),
    .A2(_1325_));
 sg13g2_a21o_1 _5163_ (.A2(_1325_),
    .A1(_1302_),
    .B1(_1326_),
    .X(_1327_));
 sg13g2_nand2_1 _5164_ (.Y(_0180_),
    .A(_1301_),
    .B(_1327_));
 sg13g2_nand3_1 _5165_ (.B(net1438),
    .C(net1124),
    .A(net709),
    .Y(_1328_));
 sg13g2_a21oi_2 _5166_ (.B1(_1324_),
    .Y(_1329_),
    .A2(_1325_),
    .A1(_1302_));
 sg13g2_nor2_1 _5167_ (.A(_3078_),
    .B(_0912_),
    .Y(_1330_));
 sg13g2_a21oi_2 _5168_ (.B1(_0901_),
    .Y(_1331_),
    .A2(_0910_),
    .A1(_0909_));
 sg13g2_xor2_1 _5169_ (.B(net1406),
    .A(net1410),
    .X(_1332_));
 sg13g2_a221oi_1 _5170_ (.B2(_0905_),
    .C1(_1330_),
    .B1(_1332_),
    .A1(_0920_),
    .Y(_1333_),
    .A2(_1331_));
 sg13g2_nor2_1 _5171_ (.A(\dtop.detune_counter[12] ),
    .B(net1221),
    .Y(_1334_));
 sg13g2_a21oi_1 _5172_ (.A1(_3114_),
    .A2(net1221),
    .Y(_1335_),
    .B1(_1334_));
 sg13g2_mux2_1 _5173_ (.A0(_1310_),
    .A1(_1335_),
    .S(net1167),
    .X(_1336_));
 sg13g2_mux2_1 _5174_ (.A0(_1289_),
    .A1(_1336_),
    .S(net1169),
    .X(_1337_));
 sg13g2_nand2_1 _5175_ (.Y(_1338_),
    .A(_0960_),
    .B(_1337_));
 sg13g2_a21oi_1 _5176_ (.A1(net1172),
    .A2(_1086_),
    .Y(_1339_),
    .B1(net1219));
 sg13g2_nor2_1 _5177_ (.A(_1259_),
    .B(_1262_),
    .Y(_1340_));
 sg13g2_and2_1 _5178_ (.A(_1273_),
    .B(_1278_),
    .X(_1341_));
 sg13g2_xnor2_1 _5179_ (.Y(_1342_),
    .A(_1257_),
    .B(_1340_));
 sg13g2_nand2_1 _5180_ (.Y(_1343_),
    .A(_1341_),
    .B(_1342_));
 sg13g2_nand3b_1 _5181_ (.B(_0996_),
    .C(\dtop.vtop.logo.addr[10] ),
    .Y(_1344_),
    .A_N(net1393));
 sg13g2_a22oi_1 _5182_ (.Y(_1345_),
    .B1(_1058_),
    .B2(\dtop.player_inst.synth.alu.registers[3][5] ),
    .A2(net1279),
    .A1(net1426));
 sg13g2_a22oi_1 _5183_ (.Y(_1346_),
    .B1(_1063_),
    .B2(\dtop.player_inst.synth.alu.registers[5][5] ),
    .A2(_0657_),
    .A1(\dtop.player_inst.synth.alu.registers[2][5] ));
 sg13g2_nand4_1 _5184_ (.B(_1344_),
    .C(_1345_),
    .A(net1220),
    .Y(_1347_),
    .D(_1346_));
 sg13g2_a221oi_1 _5185_ (.B2(\dtop.player_inst.synth.alu.registers[0][5] ),
    .C1(_1347_),
    .B1(_1064_),
    .A1(\dtop.player_inst.synth.alu.registers[1][5] ),
    .Y(_1348_),
    .A2(net1315));
 sg13g2_a22oi_1 _5186_ (.Y(_1349_),
    .B1(_1343_),
    .B2(_1348_),
    .A2(_1339_),
    .A1(_1338_));
 sg13g2_xnor2_1 _5187_ (.Y(_1350_),
    .A(_1081_),
    .B(_1349_));
 sg13g2_or2_1 _5188_ (.X(_1351_),
    .B(_1350_),
    .A(_1333_));
 sg13g2_xnor2_1 _5189_ (.Y(_1352_),
    .A(_1333_),
    .B(_1350_));
 sg13g2_nor2_1 _5190_ (.A(_1329_),
    .B(_1352_),
    .Y(_1353_));
 sg13g2_a21o_1 _5191_ (.A2(_1352_),
    .A1(_1329_),
    .B1(net1124),
    .X(_1354_));
 sg13g2_o21ai_1 _5192_ (.B1(_1328_),
    .Y(_0181_),
    .A1(_1353_),
    .A2(_1354_));
 sg13g2_nand3_1 _5193_ (.B(net1438),
    .C(net1124),
    .A(net1409),
    .Y(_1355_));
 sg13g2_o21ai_1 _5194_ (.B1(_1351_),
    .Y(_1356_),
    .A1(_1329_),
    .A2(_1352_));
 sg13g2_xnor2_1 _5195_ (.Y(_1357_),
    .A(\dtop.player_inst.synth.alu.acc[5] ),
    .B(net1407));
 sg13g2_o21ai_1 _5196_ (.B1(_1331_),
    .Y(_1358_),
    .A1(net1408),
    .A2(_0915_));
 sg13g2_o21ai_1 _5197_ (.B1(_1358_),
    .Y(_1359_),
    .A1(_0904_),
    .A2(_1357_));
 sg13g2_a221oi_1 _5198_ (.B2(net1410),
    .C1(_1359_),
    .B1(_0917_),
    .A1(net1409),
    .Y(_1360_),
    .A2(_0916_));
 sg13g2_mux2_1 _5199_ (.A0(_0059_),
    .A1(_0067_),
    .S(net1221),
    .X(_1361_));
 sg13g2_nand2_1 _5200_ (.Y(_1362_),
    .A(net1166),
    .B(_1361_));
 sg13g2_o21ai_1 _5201_ (.B1(_1362_),
    .Y(_1363_),
    .A1(net1166),
    .A2(_1335_));
 sg13g2_nor2_1 _5202_ (.A(net1169),
    .B(_1311_),
    .Y(_1364_));
 sg13g2_a21oi_1 _5203_ (.A1(net1169),
    .A2(_1363_),
    .Y(_1365_),
    .B1(_1364_));
 sg13g2_a21o_1 _5204_ (.A2(_1115_),
    .A1(net1172),
    .B1(net1219),
    .X(_1366_));
 sg13g2_a21o_1 _5205_ (.A2(_1365_),
    .A1(_0960_),
    .B1(_1366_),
    .X(_1367_));
 sg13g2_nand2_1 _5206_ (.Y(_1368_),
    .A(_1223_),
    .B(_1259_));
 sg13g2_o21ai_1 _5207_ (.B1(_1278_),
    .Y(_1369_),
    .A1(_1257_),
    .A2(_1368_));
 sg13g2_a21o_1 _5208_ (.A2(_1273_),
    .A1(_1260_),
    .B1(_1369_),
    .X(_1370_));
 sg13g2_a21oi_1 _5209_ (.A1(_1259_),
    .A2(_1274_),
    .Y(_1371_),
    .B1(_1370_));
 sg13g2_nand2_1 _5210_ (.Y(_1372_),
    .A(net1425),
    .B(net1279));
 sg13g2_nand2_1 _5211_ (.Y(_1373_),
    .A(\dtop.player_inst.synth.alu.registers[1][6] ),
    .B(net1314));
 sg13g2_a22oi_1 _5212_ (.Y(_1374_),
    .B1(_1059_),
    .B2(\dtop.vtop.logo.addr[11] ),
    .A2(net1301),
    .A1(\dtop.player_inst.synth.alu.registers[2][6] ));
 sg13g2_nand4_1 _5213_ (.B(_1372_),
    .C(_1373_),
    .A(net1220),
    .Y(_1375_),
    .D(_1374_));
 sg13g2_a21oi_1 _5214_ (.A1(\dtop.player_inst.synth.alu.registers[0][6] ),
    .A2(net1218),
    .Y(_1376_),
    .B1(_1375_));
 sg13g2_a22oi_1 _5215_ (.Y(_1377_),
    .B1(_1063_),
    .B2(\dtop.player_inst.synth.alu.registers[5][6] ),
    .A2(_1058_),
    .A1(\dtop.player_inst.synth.alu.registers[3][6] ));
 sg13g2_nand2_1 _5216_ (.Y(_1378_),
    .A(_1376_),
    .B(_1377_));
 sg13g2_o21ai_1 _5217_ (.B1(_1367_),
    .Y(_1379_),
    .A1(_1371_),
    .A2(_1378_));
 sg13g2_xnor2_1 _5218_ (.Y(_1380_),
    .A(_1082_),
    .B(_1379_));
 sg13g2_nor2_1 _5219_ (.A(_1360_),
    .B(_1380_),
    .Y(_1381_));
 sg13g2_xnor2_1 _5220_ (.Y(_1382_),
    .A(_1360_),
    .B(_1380_));
 sg13g2_inv_1 _5221_ (.Y(_1383_),
    .A(_1382_));
 sg13g2_and2_1 _5222_ (.A(_1356_),
    .B(_1383_),
    .X(_1384_));
 sg13g2_o21ai_1 _5223_ (.B1(net1111),
    .Y(_1385_),
    .A1(_1356_),
    .A2(_1383_));
 sg13g2_o21ai_1 _5224_ (.B1(_1355_),
    .Y(_0182_),
    .A1(_1384_),
    .A2(_1385_));
 sg13g2_a21oi_1 _5225_ (.A1(net1408),
    .A2(net1438),
    .Y(_1386_),
    .B1(_0875_));
 sg13g2_a21oi_1 _5226_ (.A1(_1356_),
    .A2(_1383_),
    .Y(_1387_),
    .B1(_1381_));
 sg13g2_xor2_1 _5227_ (.B(net1406),
    .A(net1409),
    .X(_1388_));
 sg13g2_a22oi_1 _5228_ (.Y(_1389_),
    .B1(_1388_),
    .B2(_0905_),
    .A2(_0917_),
    .A1(net1411));
 sg13g2_a22oi_1 _5229_ (.Y(_1390_),
    .B1(_0916_),
    .B2(net1408),
    .A2(net1224),
    .A1(\dtop.player_inst.synth.alu.acc[8] ));
 sg13g2_nand2_1 _5230_ (.Y(_1391_),
    .A(_1389_),
    .B(_1390_));
 sg13g2_mux2_1 _5231_ (.A0(_0090_),
    .A1(_0068_),
    .S(net1221),
    .X(_1392_));
 sg13g2_mux2_1 _5232_ (.A0(_1361_),
    .A1(_1392_),
    .S(net1166),
    .X(_1393_));
 sg13g2_inv_1 _5233_ (.Y(_1394_),
    .A(_1393_));
 sg13g2_mux4_1 _5234_ (.S0(net1169),
    .A0(_1085_),
    .A1(_1289_),
    .A2(_1336_),
    .A3(_1394_),
    .S1(_0960_),
    .X(_1395_));
 sg13g2_nor2_1 _5235_ (.A(net1219),
    .B(_1395_),
    .Y(_1396_));
 sg13g2_nand2_1 _5236_ (.Y(_1397_),
    .A(_1273_),
    .B(_1368_));
 sg13g2_nand3_1 _5237_ (.B(_1278_),
    .C(_1397_),
    .A(_1257_),
    .Y(_1398_));
 sg13g2_a21oi_1 _5238_ (.A1(\dtop.player_inst.synth.alu.registers[3][7] ),
    .A2(_1058_),
    .Y(_1399_),
    .B1(_1050_));
 sg13g2_a22oi_1 _5239_ (.Y(_1400_),
    .B1(net1218),
    .B2(\dtop.player_inst.synth.alu.registers[0][7] ),
    .A2(_0657_),
    .A1(\dtop.player_inst.synth.alu.registers[2][7] ));
 sg13g2_a22oi_1 _5240_ (.Y(_1401_),
    .B1(net1314),
    .B2(\dtop.player_inst.synth.alu.registers[1][7] ),
    .A2(_0996_),
    .A1(\dtop.detune_counter[4] ));
 sg13g2_nand3_1 _5241_ (.B(_1400_),
    .C(_1401_),
    .A(_1399_),
    .Y(_1402_));
 sg13g2_a21oi_1 _5242_ (.A1(_1340_),
    .A2(_1341_),
    .Y(_1403_),
    .B1(_1402_));
 sg13g2_a21oi_1 _5243_ (.A1(_1398_),
    .A2(_1403_),
    .Y(_1404_),
    .B1(_1396_));
 sg13g2_xnor2_1 _5244_ (.Y(_1405_),
    .A(_1082_),
    .B(_1404_));
 sg13g2_nor2_1 _5245_ (.A(_1391_),
    .B(_1405_),
    .Y(_1406_));
 sg13g2_nand2_1 _5246_ (.Y(_1407_),
    .A(_1391_),
    .B(_1405_));
 sg13g2_nor2b_1 _5247_ (.A(_1406_),
    .B_N(_1407_),
    .Y(_1408_));
 sg13g2_xor2_1 _5248_ (.B(_1408_),
    .A(_1387_),
    .X(_1409_));
 sg13g2_a21oi_1 _5249_ (.A1(net1111),
    .A2(_1409_),
    .Y(_0183_),
    .B1(_1386_));
 sg13g2_nand3_1 _5250_ (.B(net1435),
    .C(net1124),
    .A(net653),
    .Y(_1410_));
 sg13g2_xor2_1 _5251_ (.B(net1407),
    .A(net1408),
    .X(_1411_));
 sg13g2_a22oi_1 _5252_ (.Y(_1412_),
    .B1(_1411_),
    .B2(_0905_),
    .A2(net1224),
    .A1(\dtop.player_inst.synth.alu.acc[9] ));
 sg13g2_a22oi_1 _5253_ (.Y(_1413_),
    .B1(_0917_),
    .B2(net1412),
    .A2(net1152),
    .A1(\dtop.player_inst.synth.alu.acc[8] ));
 sg13g2_nand2_1 _5254_ (.Y(_1414_),
    .A(_1412_),
    .B(_1413_));
 sg13g2_nand3_1 _5255_ (.B(_1263_),
    .C(_1341_),
    .A(_1258_),
    .Y(_1415_));
 sg13g2_a22oi_1 _5256_ (.Y(_1416_),
    .B1(net1314),
    .B2(\dtop.player_inst.synth.alu.registers[1][8] ),
    .A2(_0996_),
    .A1(\dtop.detune_counter[5] ));
 sg13g2_nand2_1 _5257_ (.Y(_1417_),
    .A(net1219),
    .B(_1416_));
 sg13g2_a21oi_1 _5258_ (.A1(\dtop.player_inst.synth.alu.registers[0][8] ),
    .A2(net1218),
    .Y(_1418_),
    .B1(_1417_));
 sg13g2_mux2_1 _5259_ (.A0(_0062_),
    .A1(_0069_),
    .S(net1221),
    .X(_1419_));
 sg13g2_mux2_1 _5260_ (.A0(_1392_),
    .A1(_1419_),
    .S(net1166),
    .X(_1420_));
 sg13g2_nand2_1 _5261_ (.Y(_1421_),
    .A(net1169),
    .B(_1420_));
 sg13g2_a21oi_1 _5262_ (.A1(_0982_),
    .A2(_1363_),
    .Y(_1422_),
    .B1(net1171));
 sg13g2_a221oi_1 _5263_ (.B2(_1422_),
    .C1(net1219),
    .B1(_1421_),
    .A1(net1171),
    .Y(_1423_),
    .A2(_1312_));
 sg13g2_a21oi_1 _5264_ (.A1(_1415_),
    .A2(_1418_),
    .Y(_1424_),
    .B1(_1423_));
 sg13g2_xnor2_1 _5265_ (.Y(_1425_),
    .A(net1217),
    .B(_1424_));
 sg13g2_inv_1 _5266_ (.Y(_1426_),
    .A(_1425_));
 sg13g2_nand2_1 _5267_ (.Y(_1427_),
    .A(_1414_),
    .B(_1426_));
 sg13g2_xnor2_1 _5268_ (.Y(_1428_),
    .A(_1414_),
    .B(_1425_));
 sg13g2_a21oi_1 _5269_ (.A1(_1387_),
    .A2(_1407_),
    .Y(_1429_),
    .B1(_1406_));
 sg13g2_nand2_1 _5270_ (.Y(_1430_),
    .A(_1428_),
    .B(_1429_));
 sg13g2_o21ai_1 _5271_ (.B1(net1111),
    .Y(_1431_),
    .A1(_1428_),
    .A2(_1429_));
 sg13g2_nand2b_1 _5272_ (.Y(_1432_),
    .B(_1430_),
    .A_N(_1431_));
 sg13g2_nand2_1 _5273_ (.Y(_0184_),
    .A(_1410_),
    .B(_1432_));
 sg13g2_a21oi_1 _5274_ (.A1(net668),
    .A2(net1435),
    .Y(_1433_),
    .B1(net1111));
 sg13g2_nand2_1 _5275_ (.Y(_1434_),
    .A(net1406),
    .B(net1224));
 sg13g2_xnor2_1 _5276_ (.Y(_1435_),
    .A(net1407),
    .B(\dtop.player_inst.synth.alu.acc[8] ));
 sg13g2_o21ai_1 _5277_ (.B1(_1434_),
    .Y(_1436_),
    .A1(_0904_),
    .A2(_1435_));
 sg13g2_a221oi_1 _5278_ (.B2(net1413),
    .C1(_1436_),
    .B1(_0917_),
    .A1(\dtop.player_inst.synth.alu.acc[9] ),
    .Y(_1437_),
    .A2(net1152));
 sg13g2_nand2b_1 _5279_ (.Y(_1438_),
    .B(_1262_),
    .A_N(_1260_));
 sg13g2_and2_1 _5280_ (.A(net1171),
    .B(_1337_),
    .X(_1439_));
 sg13g2_and2_1 _5281_ (.A(_0981_),
    .B(net1166),
    .X(_1440_));
 sg13g2_mux2_1 _5282_ (.A0(_0089_),
    .A1(_0070_),
    .S(net1221),
    .X(_1441_));
 sg13g2_nor2_1 _5283_ (.A(_0982_),
    .B(net1166),
    .Y(_1442_));
 sg13g2_a22oi_1 _5284_ (.Y(_1443_),
    .B1(_1442_),
    .B2(_1419_),
    .A2(_1441_),
    .A1(_1440_));
 sg13g2_a21oi_1 _5285_ (.A1(_0982_),
    .A2(_1393_),
    .Y(_1444_),
    .B1(net1171));
 sg13g2_and2_1 _5286_ (.A(_1443_),
    .B(_1444_),
    .X(_1445_));
 sg13g2_o21ai_1 _5287_ (.B1(_1050_),
    .Y(_1446_),
    .A1(_1439_),
    .A2(_1445_));
 sg13g2_nand2_1 _5288_ (.Y(_1447_),
    .A(\dtop.player_inst.synth.alu.registers[0][9] ),
    .B(net1218));
 sg13g2_a22oi_1 _5289_ (.Y(_1448_),
    .B1(net1314),
    .B2(\dtop.player_inst.synth.alu.registers[1][9] ),
    .A2(_0996_),
    .A1(\dtop.detune_counter[6] ));
 sg13g2_nand3_1 _5290_ (.B(_1447_),
    .C(_1448_),
    .A(_1446_),
    .Y(_1449_));
 sg13g2_a21oi_1 _5291_ (.A1(_1341_),
    .A2(_1438_),
    .Y(_1450_),
    .B1(_1449_));
 sg13g2_xnor2_1 _5292_ (.Y(_1451_),
    .A(net1217),
    .B(_1450_));
 sg13g2_inv_1 _5293_ (.Y(_1452_),
    .A(_1451_));
 sg13g2_nor2_1 _5294_ (.A(_1437_),
    .B(_1452_),
    .Y(_1453_));
 sg13g2_xor2_1 _5295_ (.B(_1451_),
    .A(_1437_),
    .X(_1454_));
 sg13g2_and2_1 _5296_ (.A(_1427_),
    .B(_1430_),
    .X(_1455_));
 sg13g2_xnor2_1 _5297_ (.Y(_1456_),
    .A(_1454_),
    .B(_1455_));
 sg13g2_a21oi_1 _5298_ (.A1(net1111),
    .A2(_1456_),
    .Y(_0185_),
    .B1(_1433_));
 sg13g2_nand3_1 _5299_ (.B(net1435),
    .C(net1124),
    .A(net447),
    .Y(_1457_));
 sg13g2_xor2_1 _5300_ (.B(\dtop.player_inst.synth.alu.acc[9] ),
    .A(net1407),
    .X(_1458_));
 sg13g2_o21ai_1 _5301_ (.B1(_1434_),
    .Y(_1459_),
    .A1(_0904_),
    .A2(_1458_));
 sg13g2_a21oi_1 _5302_ (.A1(net1406),
    .A2(net1152),
    .Y(_1460_),
    .B1(_1459_));
 sg13g2_mux2_1 _5303_ (.A0(_0088_),
    .A1(_0071_),
    .S(net1221),
    .X(_1461_));
 sg13g2_a22oi_1 _5304_ (.Y(_1462_),
    .B1(_1461_),
    .B2(_1440_),
    .A2(_1442_),
    .A1(_1441_));
 sg13g2_a21oi_1 _5305_ (.A1(_0982_),
    .A2(_1420_),
    .Y(_1463_),
    .B1(net1171));
 sg13g2_a221oi_1 _5306_ (.B2(_1463_),
    .C1(net1219),
    .B1(_1462_),
    .A1(net1171),
    .Y(_1464_),
    .A2(_1365_));
 sg13g2_a21oi_1 _5307_ (.A1(\dtop.player_inst.synth.alu.registers[1][10] ),
    .A2(net1315),
    .Y(_1465_),
    .B1(_1050_));
 sg13g2_nand2_1 _5308_ (.Y(_1466_),
    .A(_1029_),
    .B(_1032_));
 sg13g2_nor2_1 _5309_ (.A(_0063_),
    .B(_1466_),
    .Y(_1467_));
 sg13g2_a22oi_1 _5310_ (.Y(_1468_),
    .B1(_1135_),
    .B2(_1467_),
    .A2(net1218),
    .A1(\dtop.player_inst.synth.alu.registers[0][10] ));
 sg13g2_a21oi_1 _5311_ (.A1(_1465_),
    .A2(_1468_),
    .Y(_1469_),
    .B1(_1464_));
 sg13g2_xnor2_1 _5312_ (.Y(_1470_),
    .A(_1081_),
    .B(_1469_));
 sg13g2_xor2_1 _5313_ (.B(_1470_),
    .A(_1460_),
    .X(_1471_));
 sg13g2_a21oi_1 _5314_ (.A1(_1414_),
    .A2(_1426_),
    .Y(_1472_),
    .B1(_1453_));
 sg13g2_a22oi_1 _5315_ (.Y(_1473_),
    .B1(_1472_),
    .B2(_1430_),
    .A2(_1452_),
    .A1(_1437_));
 sg13g2_o21ai_1 _5316_ (.B1(net1111),
    .Y(_1474_),
    .A1(_1471_),
    .A2(_1473_));
 sg13g2_a21o_1 _5317_ (.A2(_1473_),
    .A1(_1471_),
    .B1(_1474_),
    .X(_1475_));
 sg13g2_nand2_1 _5318_ (.Y(_0186_),
    .A(_1457_),
    .B(_1475_));
 sg13g2_nor2_1 _5319_ (.A(_0873_),
    .B(_0885_),
    .Y(_1476_));
 sg13g2_nor3_2 _5320_ (.A(_0087_),
    .B(_0749_),
    .C(_1476_),
    .Y(_1477_));
 sg13g2_o21ai_1 _5321_ (.B1(_1477_),
    .Y(_1478_),
    .A1(_1460_),
    .A2(_1470_));
 sg13g2_a21oi_1 _5322_ (.A1(_1471_),
    .A2(_1473_),
    .Y(_1479_),
    .B1(_1478_));
 sg13g2_o21ai_1 _5323_ (.B1(net1438),
    .Y(_1480_),
    .A1(net600),
    .A2(_1477_));
 sg13g2_nor2_1 _5324_ (.A(_1479_),
    .B(_1480_),
    .Y(_0187_));
 sg13g2_nand2_1 _5325_ (.Y(_1481_),
    .A(_0750_),
    .B(_0836_));
 sg13g2_o21ai_1 _5326_ (.B1(net1432),
    .Y(_1482_),
    .A1(net1414),
    .A2(net1123));
 sg13g2_a21oi_1 _5327_ (.A1(_3090_),
    .A2(net1123),
    .Y(_0188_),
    .B1(_1482_));
 sg13g2_o21ai_1 _5328_ (.B1(net1432),
    .Y(_1483_),
    .A1(net1413),
    .A2(net1122));
 sg13g2_a21oi_1 _5329_ (.A1(_3089_),
    .A2(net1123),
    .Y(_0189_),
    .B1(_1483_));
 sg13g2_o21ai_1 _5330_ (.B1(net1427),
    .Y(_1484_),
    .A1(net1412),
    .A2(net1122));
 sg13g2_a21oi_1 _5331_ (.A1(_3088_),
    .A2(net1122),
    .Y(_0190_),
    .B1(_1484_));
 sg13g2_o21ai_1 _5332_ (.B1(net1433),
    .Y(_1485_),
    .A1(\dtop.player_inst.synth.alu.acc[3] ),
    .A2(net1123));
 sg13g2_a21oi_1 _5333_ (.A1(_3087_),
    .A2(net1123),
    .Y(_0191_),
    .B1(_1485_));
 sg13g2_o21ai_1 _5334_ (.B1(net1427),
    .Y(_1486_),
    .A1(net1410),
    .A2(net1122));
 sg13g2_a21oi_1 _5335_ (.A1(_3086_),
    .A2(net1122),
    .Y(_0192_),
    .B1(_1486_));
 sg13g2_o21ai_1 _5336_ (.B1(net1433),
    .Y(_1487_),
    .A1(\dtop.player_inst.synth.alu.acc[5] ),
    .A2(net1122));
 sg13g2_a21oi_1 _5337_ (.A1(_3085_),
    .A2(net1122),
    .Y(_0193_),
    .B1(_1487_));
 sg13g2_o21ai_1 _5338_ (.B1(net1432),
    .Y(_1488_),
    .A1(net1409),
    .A2(net1123));
 sg13g2_a21oi_1 _5339_ (.A1(_3084_),
    .A2(net1122),
    .Y(_0194_),
    .B1(_1488_));
 sg13g2_nand2_1 _5340_ (.Y(_1489_),
    .A(_0678_),
    .B(_0778_));
 sg13g2_nand3_1 _5341_ (.B(net1432),
    .C(net1120),
    .A(net356),
    .Y(_1490_));
 sg13g2_o21ai_1 _5342_ (.B1(_1490_),
    .Y(_0195_),
    .A1(_3083_),
    .A2(net1120));
 sg13g2_nand3_1 _5343_ (.B(net1431),
    .C(net1119),
    .A(net410),
    .Y(_1491_));
 sg13g2_o21ai_1 _5344_ (.B1(_1491_),
    .Y(_0196_),
    .A1(_3082_),
    .A2(net1119));
 sg13g2_nand3_1 _5345_ (.B(net1427),
    .C(net1121),
    .A(net428),
    .Y(_1492_));
 sg13g2_o21ai_1 _5346_ (.B1(_1492_),
    .Y(_0197_),
    .A1(_3081_),
    .A2(net1121));
 sg13g2_nand3_1 _5347_ (.B(net1431),
    .C(net1120),
    .A(net398),
    .Y(_1493_));
 sg13g2_o21ai_1 _5348_ (.B1(_1493_),
    .Y(_0198_),
    .A1(_3080_),
    .A2(net1120));
 sg13g2_nand3_1 _5349_ (.B(net1427),
    .C(net1121),
    .A(net391),
    .Y(_1494_));
 sg13g2_o21ai_1 _5350_ (.B1(_1494_),
    .Y(_0199_),
    .A1(_3079_),
    .A2(net1121));
 sg13g2_nand3_1 _5351_ (.B(net1431),
    .C(net1119),
    .A(net512),
    .Y(_1495_));
 sg13g2_o21ai_1 _5352_ (.B1(_1495_),
    .Y(_0200_),
    .A1(_3078_),
    .A2(net1119));
 sg13g2_nand3_1 _5353_ (.B(net1432),
    .C(net1119),
    .A(net351),
    .Y(_1496_));
 sg13g2_o21ai_1 _5354_ (.B1(_1496_),
    .Y(_0201_),
    .A1(_3077_),
    .A2(net1119));
 sg13g2_nand3_1 _5355_ (.B(net1431),
    .C(net1119),
    .A(net359),
    .Y(_1497_));
 sg13g2_o21ai_1 _5356_ (.B1(_1497_),
    .Y(_0202_),
    .A1(_3076_),
    .A2(net1119));
 sg13g2_nor2_1 _5357_ (.A(_0080_),
    .B(_0578_),
    .Y(_1498_));
 sg13g2_nand3b_1 _5358_ (.B(_0079_),
    .C(_1498_),
    .Y(_1499_),
    .A_N(net1393));
 sg13g2_nor2_2 _5359_ (.A(_0561_),
    .B(_1499_),
    .Y(_1500_));
 sg13g2_nor2b_1 _5360_ (.A(_1500_),
    .B_N(net663),
    .Y(_1501_));
 sg13g2_nand2b_2 _5361_ (.Y(_1502_),
    .B(\dtop.detune_counter[4] ),
    .A_N(_1501_));
 sg13g2_nor2_1 _5362_ (.A(_0077_),
    .B(_1502_),
    .Y(_1503_));
 sg13g2_and2_1 _5363_ (.A(net646),
    .B(_1503_),
    .X(_1504_));
 sg13g2_and3_1 _5364_ (.X(_1505_),
    .A(net1404),
    .B(net1405),
    .C(_1504_));
 sg13g2_and2_2 _5365_ (.A(_0735_),
    .B(_1505_),
    .X(_1506_));
 sg13g2_nand2_1 _5366_ (.Y(_1507_),
    .A(net1399),
    .B(_1506_));
 sg13g2_nand3_1 _5367_ (.B(net1328),
    .C(_1506_),
    .A(net1396),
    .Y(_1508_));
 sg13g2_xor2_1 _5368_ (.B(_1508_),
    .A(net636),
    .X(_1509_));
 sg13g2_nor2_1 _5369_ (.A(net661),
    .B(_1508_),
    .Y(_1510_));
 sg13g2_xnor2_1 _5370_ (.Y(_1511_),
    .A(_3146_),
    .B(_1510_));
 sg13g2_o21ai_1 _5371_ (.B1(net1440),
    .Y(_1512_),
    .A1(_1509_),
    .A2(_1511_));
 sg13g2_and2_1 _5372_ (.A(_0078_),
    .B(_1512_),
    .X(_1513_));
 sg13g2_xnor2_1 _5373_ (.Y(_1514_),
    .A(net665),
    .B(_1501_));
 sg13g2_nor2_1 _5374_ (.A(net1095),
    .B(_1514_),
    .Y(_0203_));
 sg13g2_xor2_1 _5375_ (.B(_1502_),
    .A(net656),
    .X(_1515_));
 sg13g2_nor2_1 _5376_ (.A(net1095),
    .B(_1515_),
    .Y(_0204_));
 sg13g2_nor2_1 _5377_ (.A(net646),
    .B(_1503_),
    .Y(_1516_));
 sg13g2_nor3_1 _5378_ (.A(_1504_),
    .B(net1096),
    .C(net647),
    .Y(_0205_));
 sg13g2_nor3_1 _5379_ (.A(_0077_),
    .B(_0023_),
    .C(_1502_),
    .Y(_1517_));
 sg13g2_xnor2_1 _5380_ (.Y(_1518_),
    .A(net1405),
    .B(_1517_));
 sg13g2_nor2_1 _5381_ (.A(net1095),
    .B(net688),
    .Y(_0206_));
 sg13g2_a21oi_1 _5382_ (.A1(net1405),
    .A2(_1504_),
    .Y(_1519_),
    .B1(net1404));
 sg13g2_nor3_1 _5383_ (.A(_1505_),
    .B(net1096),
    .C(net667),
    .Y(_0207_));
 sg13g2_and3_1 _5384_ (.X(_1520_),
    .A(net1405),
    .B(_3159_),
    .C(_1504_));
 sg13g2_xnor2_1 _5385_ (.Y(_1521_),
    .A(net1402),
    .B(_1520_));
 sg13g2_nor2_1 _5386_ (.A(net1096),
    .B(_1521_),
    .Y(_0208_));
 sg13g2_a21oi_1 _5387_ (.A1(net571),
    .A2(_1505_),
    .Y(_1522_),
    .B1(net1401));
 sg13g2_nor3_1 _5388_ (.A(_1506_),
    .B(net1096),
    .C(net572),
    .Y(_0209_));
 sg13g2_nand3b_1 _5389_ (.B(_1505_),
    .C(net571),
    .Y(_1523_),
    .A_N(_0016_));
 sg13g2_xnor2_1 _5390_ (.Y(_1524_),
    .A(net1399),
    .B(_1523_));
 sg13g2_nor2b_1 _5391_ (.A(net1096),
    .B_N(_1524_),
    .Y(_0210_));
 sg13g2_xnor2_1 _5392_ (.Y(_1525_),
    .A(net698),
    .B(_1507_));
 sg13g2_nor2_1 _5393_ (.A(net1096),
    .B(_1525_),
    .Y(_0211_));
 sg13g2_nand3_1 _5394_ (.B(_3321_),
    .C(_1506_),
    .A(net568),
    .Y(_1526_));
 sg13g2_a21oi_1 _5395_ (.A1(_3321_),
    .A2(_1506_),
    .Y(_1527_),
    .B1(net1397));
 sg13g2_nor2_1 _5396_ (.A(net1095),
    .B(_1527_),
    .Y(_1528_));
 sg13g2_and2_1 _5397_ (.A(_1526_),
    .B(_1528_),
    .X(_0212_));
 sg13g2_a221oi_1 _5398_ (.B2(_3126_),
    .C1(net1095),
    .B1(_1526_),
    .A1(net1328),
    .Y(_0213_),
    .A2(_1506_));
 sg13g2_nor2_1 _5399_ (.A(_0090_),
    .B(_1526_),
    .Y(_1529_));
 sg13g2_xnor2_1 _5400_ (.Y(_1530_),
    .A(net583),
    .B(_1529_));
 sg13g2_nor2_1 _5401_ (.A(net1095),
    .B(_1530_),
    .Y(_0214_));
 sg13g2_nor2_1 _5402_ (.A(_1509_),
    .B(net1095),
    .Y(_0215_));
 sg13g2_nor2_1 _5403_ (.A(_1511_),
    .B(net1095),
    .Y(_0216_));
 sg13g2_and3_2 _5404_ (.X(_1531_),
    .A(_0083_),
    .B(_3228_),
    .C(_0676_));
 sg13g2_nand4_1 _5405_ (.B(_0083_),
    .C(_3228_),
    .A(net1367),
    .Y(_1532_),
    .D(_0637_));
 sg13g2_nand2_1 _5406_ (.Y(_1533_),
    .A(_0093_),
    .B(net1299));
 sg13g2_nand3_1 _5407_ (.B(_0601_),
    .C(net1296),
    .A(_0093_),
    .Y(_1534_));
 sg13g2_nand2_1 _5408_ (.Y(_1535_),
    .A(_3147_),
    .B(\dtop.vtop.pipeline.wave_index[1] ));
 sg13g2_nand2_1 _5409_ (.Y(_1536_),
    .A(_0001_),
    .B(net1295));
 sg13g2_o21ai_1 _5410_ (.B1(_1536_),
    .Y(_1537_),
    .A1(net1295),
    .A2(_1535_));
 sg13g2_nand2_1 _5411_ (.Y(_1538_),
    .A(net1388),
    .B(net1295));
 sg13g2_nor2_1 _5412_ (.A(_3147_),
    .B(_3148_),
    .Y(_1539_));
 sg13g2_and2_1 _5413_ (.A(_3202_),
    .B(_1539_),
    .X(_1540_));
 sg13g2_o21ai_1 _5414_ (.B1(net1307),
    .Y(_1541_),
    .A1(_0004_),
    .A2(_1539_));
 sg13g2_o21ai_1 _5415_ (.B1(_1538_),
    .Y(_1542_),
    .A1(_1540_),
    .A2(_1541_));
 sg13g2_inv_4 _5416_ (.A(net1252),
    .Y(_1543_));
 sg13g2_mux2_2 _5417_ (.A0(_3150_),
    .A1(_3153_),
    .S(net1308),
    .X(_1544_));
 sg13g2_mux2_1 _5418_ (.A0(_0001_),
    .A1(_0005_),
    .S(net1311),
    .X(_1545_));
 sg13g2_mux2_2 _5419_ (.A0(_0003_),
    .A1(_0004_),
    .S(net1309),
    .X(_1546_));
 sg13g2_mux2_1 _5420_ (.A0(_3152_),
    .A1(_3151_),
    .S(net1309),
    .X(_1547_));
 sg13g2_nor2_1 _5421_ (.A(_1544_),
    .B(net1285),
    .Y(_1548_));
 sg13g2_nand2_1 _5422_ (.Y(_1549_),
    .A(_0002_),
    .B(net1274));
 sg13g2_nor2_2 _5423_ (.A(net1291),
    .B(net1285),
    .Y(_1550_));
 sg13g2_nand2_2 _5424_ (.Y(_1551_),
    .A(_1544_),
    .B(net1288));
 sg13g2_o21ai_1 _5425_ (.B1(net1287),
    .Y(_1552_),
    .A1(\dtop.vtop.pipeline.phases[2][15] ),
    .A2(net1290));
 sg13g2_nor2_1 _5426_ (.A(net1290),
    .B(net1287),
    .Y(_1553_));
 sg13g2_nand3_1 _5427_ (.B(_1544_),
    .C(net1285),
    .A(\dtop.vtop.pipeline.zg_acc[8] ),
    .Y(_1554_));
 sg13g2_nand2_1 _5428_ (.Y(_1555_),
    .A(\dtop.vtop.pipeline.phases[1][15] ),
    .B(net1290));
 sg13g2_nor2_1 _5429_ (.A(_1544_),
    .B(net1288),
    .Y(_1556_));
 sg13g2_nand3_1 _5430_ (.B(_1554_),
    .C(_1555_),
    .A(_1552_),
    .Y(_1557_));
 sg13g2_nand2_2 _5431_ (.Y(_1558_),
    .A(_1549_),
    .B(_1557_));
 sg13g2_a21oi_2 _5432_ (.B1(_0440_),
    .Y(_1559_),
    .A2(net1299),
    .A1(_0434_));
 sg13g2_or2_1 _5433_ (.X(_1560_),
    .B(_1559_),
    .A(net1241));
 sg13g2_nand3_1 _5434_ (.B(_1557_),
    .C(_1559_),
    .A(_1549_),
    .Y(_1561_));
 sg13g2_nand2b_1 _5435_ (.Y(_1562_),
    .B(_1553_),
    .A_N(_0061_));
 sg13g2_a221oi_1 _5436_ (.B2(\dtop.vtop.pipeline.phases[1][14] ),
    .C1(net1274),
    .B1(net1272),
    .A1(\dtop.vtop.pipeline.phases[2][14] ),
    .Y(_1563_),
    .A2(_1550_));
 sg13g2_a22oi_1 _5437_ (.Y(_1564_),
    .B1(_1562_),
    .B2(_1563_),
    .A2(net1274),
    .A1(_0060_));
 sg13g2_xnor2_1 _5438_ (.Y(_1565_),
    .A(_1561_),
    .B(_1564_));
 sg13g2_o21ai_1 _5439_ (.B1(net1287),
    .Y(_1566_),
    .A1(\dtop.vtop.pipeline.phases[2][12] ),
    .A2(net1290));
 sg13g2_a22oi_1 _5440_ (.Y(_1567_),
    .B1(net1270),
    .B2(\dtop.vtop.pipeline.phases[1][12] ),
    .A2(net1273),
    .A1(\dtop.vtop.pipeline.zg_acc[5] ));
 sg13g2_and2_1 _5441_ (.A(_1566_),
    .B(_1567_),
    .X(_1568_));
 sg13g2_a21o_1 _5442_ (.A2(net1274),
    .A1(_0056_),
    .B1(_1568_),
    .X(_1569_));
 sg13g2_xor2_1 _5443_ (.B(_1569_),
    .A(net1237),
    .X(_1570_));
 sg13g2_o21ai_1 _5444_ (.B1(net1287),
    .Y(_1571_),
    .A1(\dtop.vtop.pipeline.phases[2][10] ),
    .A2(net1289));
 sg13g2_a22oi_1 _5445_ (.Y(_1572_),
    .B1(net1272),
    .B2(\dtop.vtop.pipeline.phases[1][10] ),
    .A2(_1553_),
    .A1(\dtop.vtop.pipeline.zg_acc[3] ));
 sg13g2_and2_1 _5446_ (.A(_1571_),
    .B(_1572_),
    .X(_1573_));
 sg13g2_a21o_2 _5447_ (.A2(net1274),
    .A1(_0052_),
    .B1(_1573_),
    .X(_1574_));
 sg13g2_xnor2_1 _5448_ (.Y(_1575_),
    .A(net1236),
    .B(_1574_));
 sg13g2_xor2_1 _5449_ (.B(_1574_),
    .A(net1235),
    .X(_1576_));
 sg13g2_o21ai_1 _5450_ (.B1(net1287),
    .Y(_1577_),
    .A1(\dtop.vtop.pipeline.phases[2][8] ),
    .A2(net1289));
 sg13g2_a22oi_1 _5451_ (.Y(_1578_),
    .B1(net1272),
    .B2(\dtop.vtop.pipeline.phases[1][8] ),
    .A2(net1273),
    .A1(\dtop.vtop.pipeline.zg_acc[1] ));
 sg13g2_a22oi_1 _5452_ (.Y(_1579_),
    .B1(_1577_),
    .B2(_1578_),
    .A2(net1274),
    .A1(_0047_));
 sg13g2_xor2_1 _5453_ (.B(_1579_),
    .A(net1235),
    .X(_1580_));
 sg13g2_xnor2_1 _5454_ (.Y(_1581_),
    .A(net1235),
    .B(_1579_));
 sg13g2_a22oi_1 _5455_ (.Y(_1582_),
    .B1(net1272),
    .B2(\dtop.vtop.pipeline.phases[1][7] ),
    .A2(net1273),
    .A1(\dtop.vtop.pipeline.zg_acc[0] ));
 sg13g2_o21ai_1 _5456_ (.B1(_1546_),
    .Y(_1583_),
    .A1(\dtop.vtop.pipeline.phases[2][7] ),
    .A2(net1291));
 sg13g2_a22oi_1 _5457_ (.Y(_1584_),
    .B1(_1582_),
    .B2(_1583_),
    .A2(net1275),
    .A1(_0044_));
 sg13g2_xor2_1 _5458_ (.B(_1584_),
    .A(net1235),
    .X(_1585_));
 sg13g2_xnor2_1 _5459_ (.Y(_1586_),
    .A(net1235),
    .B(_1584_));
 sg13g2_nand2_1 _5460_ (.Y(_1587_),
    .A(\dtop.vtop.pipeline.phases[1][6] ),
    .B(net1291));
 sg13g2_o21ai_1 _5461_ (.B1(net1288),
    .Y(_1588_),
    .A1(\dtop.vtop.pipeline.phases[2][6] ),
    .A2(net1291));
 sg13g2_a22oi_1 _5462_ (.Y(_1589_),
    .B1(_1587_),
    .B2(_1588_),
    .A2(net1275),
    .A1(_0042_));
 sg13g2_xor2_1 _5463_ (.B(_1589_),
    .A(net1235),
    .X(_1590_));
 sg13g2_xnor2_1 _5464_ (.Y(_1591_),
    .A(net1235),
    .B(_1589_));
 sg13g2_a21oi_1 _5465_ (.A1(net1197),
    .A2(net1196),
    .Y(_1592_),
    .B1(net1202));
 sg13g2_o21ai_1 _5466_ (.B1(net1204),
    .Y(_1593_),
    .A1(net1199),
    .A2(_1591_));
 sg13g2_o21ai_1 _5467_ (.B1(net1287),
    .Y(_1594_),
    .A1(\dtop.vtop.pipeline.phases[2][9] ),
    .A2(net1289));
 sg13g2_a22oi_1 _5468_ (.Y(_1595_),
    .B1(net1271),
    .B2(\dtop.vtop.pipeline.phases[1][9] ),
    .A2(net1273),
    .A1(\dtop.vtop.pipeline.zg_acc[2] ));
 sg13g2_a22oi_1 _5469_ (.Y(_1596_),
    .B1(_1594_),
    .B2(_1595_),
    .A2(net1274),
    .A1(_0049_));
 sg13g2_xor2_1 _5470_ (.B(_1596_),
    .A(net1236),
    .X(_1597_));
 sg13g2_xnor2_1 _5471_ (.Y(_1598_),
    .A(net1235),
    .B(_1596_));
 sg13g2_nand2_2 _5472_ (.Y(_1599_),
    .A(net1197),
    .B(net1195));
 sg13g2_xor2_1 _5473_ (.B(_1589_),
    .A(_1584_),
    .X(_1600_));
 sg13g2_xnor2_1 _5474_ (.Y(_1601_),
    .A(_1584_),
    .B(_1589_));
 sg13g2_a21oi_1 _5475_ (.A1(net1199),
    .A2(net1196),
    .Y(_1602_),
    .B1(net1203));
 sg13g2_o21ai_1 _5476_ (.B1(net1200),
    .Y(_1603_),
    .A1(net1198),
    .A2(net1195));
 sg13g2_o21ai_1 _5477_ (.B1(net1189),
    .Y(_1604_),
    .A1(net1204),
    .A2(_1601_));
 sg13g2_nor3_1 _5478_ (.A(net1208),
    .B(_1592_),
    .C(_1604_),
    .Y(_1605_));
 sg13g2_nand3_1 _5479_ (.B(net1199),
    .C(net1195),
    .A(net1202),
    .Y(_1606_));
 sg13g2_nand2_1 _5480_ (.Y(_1607_),
    .A(net1194),
    .B(_1606_));
 sg13g2_o21ai_1 _5481_ (.B1(net1204),
    .Y(_1608_),
    .A1(net1197),
    .A2(net1196));
 sg13g2_nand2_1 _5482_ (.Y(_1609_),
    .A(net1208),
    .B(_1608_));
 sg13g2_nor2b_1 _5483_ (.A(_1604_),
    .B_N(_1608_),
    .Y(_1610_));
 sg13g2_a21oi_1 _5484_ (.A1(_1604_),
    .A2(_1607_),
    .Y(_1611_),
    .B1(_1609_));
 sg13g2_nand2_2 _5485_ (.Y(_1612_),
    .A(net1202),
    .B(_1590_));
 sg13g2_nor2_2 _5486_ (.A(net1208),
    .B(net1189),
    .Y(_1613_));
 sg13g2_nand2_2 _5487_ (.Y(_1614_),
    .A(net1209),
    .B(net1191));
 sg13g2_nor2_1 _5488_ (.A(net1200),
    .B(net1198),
    .Y(_1615_));
 sg13g2_nand2_1 _5489_ (.Y(_1616_),
    .A(net1203),
    .B(net1199));
 sg13g2_a21oi_1 _5490_ (.A1(net1196),
    .A2(_1616_),
    .Y(_1617_),
    .B1(_1614_));
 sg13g2_o21ai_1 _5491_ (.B1(net1292),
    .Y(_1618_),
    .A1(\dtop.vtop.pipeline.phases[1][11] ),
    .A2(net1288));
 sg13g2_a22oi_1 _5492_ (.Y(_1619_),
    .B1(net1273),
    .B2(\dtop.vtop.pipeline.zg_acc[4] ),
    .A2(_1550_),
    .A1(\dtop.vtop.pipeline.phases[2][11] ));
 sg13g2_a22oi_1 _5493_ (.Y(_1620_),
    .B1(_1618_),
    .B2(_1619_),
    .A2(net1275),
    .A1(_0054_));
 sg13g2_inv_1 _5494_ (.Y(_1621_),
    .A(_1620_));
 sg13g2_xnor2_1 _5495_ (.Y(_1622_),
    .A(net1237),
    .B(_1621_));
 sg13g2_xnor2_1 _5496_ (.Y(_1623_),
    .A(net1236),
    .B(_1620_));
 sg13g2_nor4_1 _5497_ (.A(net1215),
    .B(_1605_),
    .C(_1611_),
    .D(_1617_),
    .Y(_1624_));
 sg13g2_and2_1 _5498_ (.A(net1215),
    .B(_1585_),
    .X(_1625_));
 sg13g2_o21ai_1 _5499_ (.B1(net1184),
    .Y(_1626_),
    .A1(_1624_),
    .A2(_1625_));
 sg13g2_o21ai_1 _5500_ (.B1(net1288),
    .Y(_1627_),
    .A1(\dtop.vtop.pipeline.phases[2][13] ),
    .A2(net1290));
 sg13g2_a22oi_1 _5501_ (.Y(_1628_),
    .B1(net1273),
    .B2(_3176_),
    .A2(net1290),
    .A1(\dtop.vtop.pipeline.phases[1][13] ));
 sg13g2_a22oi_1 _5502_ (.Y(_1629_),
    .B1(_1627_),
    .B2(_1628_),
    .A2(net1274),
    .A1(_0057_));
 sg13g2_xnor2_1 _5503_ (.Y(_1630_),
    .A(net1237),
    .B(_1629_));
 sg13g2_inv_1 _5504_ (.Y(_1631_),
    .A(net1179));
 sg13g2_a21oi_1 _5505_ (.A1(net1197),
    .A2(_1612_),
    .Y(_1632_),
    .B1(net1190));
 sg13g2_nand2_2 _5506_ (.Y(_1633_),
    .A(net1202),
    .B(net1197));
 sg13g2_o21ai_1 _5507_ (.B1(net1203),
    .Y(_1634_),
    .A1(net1197),
    .A2(net1195));
 sg13g2_nand2_1 _5508_ (.Y(_1635_),
    .A(net1204),
    .B(_1600_));
 sg13g2_nand2_1 _5509_ (.Y(_1636_),
    .A(net1204),
    .B(_1601_));
 sg13g2_a21oi_1 _5510_ (.A1(_1633_),
    .A2(_1635_),
    .Y(_1637_),
    .B1(net1194));
 sg13g2_nor2_1 _5511_ (.A(net1211),
    .B(_1637_),
    .Y(_1638_));
 sg13g2_or3_1 _5512_ (.A(net1211),
    .B(_1632_),
    .C(_1637_),
    .X(_1639_));
 sg13g2_nand3_1 _5513_ (.B(net1199),
    .C(net1196),
    .A(_1581_),
    .Y(_1640_));
 sg13g2_and3_1 _5514_ (.X(_1641_),
    .A(net1193),
    .B(_1599_),
    .C(_1640_));
 sg13g2_o21ai_1 _5515_ (.B1(net1211),
    .Y(_1642_),
    .A1(_1637_),
    .A2(_1641_));
 sg13g2_nand3_1 _5516_ (.B(_1639_),
    .C(_1642_),
    .A(net1214),
    .Y(_1643_));
 sg13g2_nand3_1 _5517_ (.B(net1197),
    .C(_1590_),
    .A(net1202),
    .Y(_1644_));
 sg13g2_and3_1 _5518_ (.X(_1645_),
    .A(_1593_),
    .B(net1193),
    .C(_1644_));
 sg13g2_a21oi_1 _5519_ (.A1(_1636_),
    .A2(_1644_),
    .Y(_1646_),
    .B1(net1193));
 sg13g2_or3_1 _5520_ (.A(net1208),
    .B(_1645_),
    .C(_1646_),
    .X(_1647_));
 sg13g2_a21oi_2 _5521_ (.B1(net1190),
    .Y(_1648_),
    .A2(_1586_),
    .A1(net1202));
 sg13g2_o21ai_1 _5522_ (.B1(net1193),
    .Y(_1649_),
    .A1(net1203),
    .A2(net1199));
 sg13g2_a221oi_1 _5523_ (.B2(_1648_),
    .C1(net1211),
    .B1(_1636_),
    .A1(net1190),
    .Y(_1650_),
    .A2(_1601_));
 sg13g2_nor2_1 _5524_ (.A(net1214),
    .B(_1650_),
    .Y(_1651_));
 sg13g2_a21oi_1 _5525_ (.A1(_1647_),
    .A2(_1651_),
    .Y(_1652_),
    .B1(net1185));
 sg13g2_a21oi_1 _5526_ (.A1(_1643_),
    .A2(_1652_),
    .Y(_1653_),
    .B1(_1631_));
 sg13g2_nor2_1 _5527_ (.A(net1214),
    .B(net1178),
    .Y(_1654_));
 sg13g2_or2_1 _5528_ (.X(_1655_),
    .B(net1180),
    .A(net1213));
 sg13g2_o21ai_1 _5529_ (.B1(net1187),
    .Y(_1656_),
    .A1(net1200),
    .A2(net1198));
 sg13g2_a21o_1 _5530_ (.A2(_1600_),
    .A1(net1200),
    .B1(_1656_),
    .X(_1657_));
 sg13g2_o21ai_1 _5531_ (.B1(net1191),
    .Y(_1658_),
    .A1(_1602_),
    .A2(_1615_));
 sg13g2_nand3_1 _5532_ (.B(_1657_),
    .C(_1658_),
    .A(net1209),
    .Y(_1659_));
 sg13g2_nand2_2 _5533_ (.Y(_1660_),
    .A(net1201),
    .B(net1187));
 sg13g2_nand3_1 _5534_ (.B(net1198),
    .C(net1187),
    .A(net1200),
    .Y(_1661_));
 sg13g2_nand3_1 _5535_ (.B(_1600_),
    .C(_1661_),
    .A(net1205),
    .Y(_1662_));
 sg13g2_nand3_1 _5536_ (.B(_1659_),
    .C(_1662_),
    .A(net1181),
    .Y(_1663_));
 sg13g2_nor3_2 _5537_ (.A(net1202),
    .B(net1197),
    .C(net1188),
    .Y(_1664_));
 sg13g2_nor2_1 _5538_ (.A(net1209),
    .B(_1664_),
    .Y(_1665_));
 sg13g2_nand3_1 _5539_ (.B(net1188),
    .C(_1599_),
    .A(net1203),
    .Y(_1666_));
 sg13g2_nand3_1 _5540_ (.B(net1198),
    .C(net1195),
    .A(net1200),
    .Y(_1667_));
 sg13g2_nand3_1 _5541_ (.B(_1666_),
    .C(_1667_),
    .A(_1665_),
    .Y(_1668_));
 sg13g2_nand2_1 _5542_ (.Y(_1669_),
    .A(net1209),
    .B(_1656_));
 sg13g2_nand3_1 _5543_ (.B(_1668_),
    .C(_1669_),
    .A(net1183),
    .Y(_1670_));
 sg13g2_a21oi_1 _5544_ (.A1(_1663_),
    .A2(_1670_),
    .Y(_1671_),
    .B1(_1655_));
 sg13g2_nand4_1 _5545_ (.B(_1612_),
    .C(_1613_),
    .A(_1593_),
    .Y(_1672_),
    .D(_1633_));
 sg13g2_nand2_1 _5546_ (.Y(_1673_),
    .A(net1184),
    .B(_1672_));
 sg13g2_nor2_1 _5547_ (.A(net1195),
    .B(_1616_),
    .Y(_1674_));
 sg13g2_nand3_1 _5548_ (.B(net1199),
    .C(net1196),
    .A(net1203),
    .Y(_1675_));
 sg13g2_nand2_1 _5549_ (.Y(_1676_),
    .A(net1188),
    .B(_1675_));
 sg13g2_nor2_1 _5550_ (.A(net1211),
    .B(_1676_),
    .Y(_1677_));
 sg13g2_nand3_1 _5551_ (.B(net1188),
    .C(_1675_),
    .A(net1207),
    .Y(_1678_));
 sg13g2_a21oi_1 _5552_ (.A1(net1195),
    .A2(_1616_),
    .Y(_1679_),
    .B1(_1676_));
 sg13g2_or3_1 _5553_ (.A(net1212),
    .B(_1645_),
    .C(_1679_),
    .X(_1680_));
 sg13g2_a21oi_1 _5554_ (.A1(net1212),
    .A2(_1646_),
    .Y(_1681_),
    .B1(_1673_));
 sg13g2_nor2b_2 _5555_ (.A(net1178),
    .B_N(net1214),
    .Y(_1682_));
 sg13g2_nand2_2 _5556_ (.Y(_1683_),
    .A(net1207),
    .B(_1664_));
 sg13g2_nor2_1 _5557_ (.A(net1195),
    .B(_1683_),
    .Y(_1684_));
 sg13g2_nor2_1 _5558_ (.A(net1205),
    .B(_1661_),
    .Y(_1685_));
 sg13g2_xnor2_1 _5559_ (.Y(_1686_),
    .A(net1196),
    .B(_1683_));
 sg13g2_nor3_1 _5560_ (.A(net1184),
    .B(_1685_),
    .C(_1686_),
    .Y(_1687_));
 sg13g2_a21oi_1 _5561_ (.A1(_1680_),
    .A2(_1681_),
    .Y(_1688_),
    .B1(_1687_));
 sg13g2_a221oi_1 _5562_ (.B2(_1688_),
    .C1(_1671_),
    .B1(_1682_),
    .A1(_1626_),
    .Y(_1689_),
    .A2(_1653_));
 sg13g2_xor2_1 _5563_ (.B(_1689_),
    .A(net1238),
    .X(_1690_));
 sg13g2_xnor2_1 _5564_ (.Y(_1691_),
    .A(net1239),
    .B(_1689_));
 sg13g2_a21o_1 _5565_ (.A2(_1612_),
    .A1(_1593_),
    .B1(net1189),
    .X(_1692_));
 sg13g2_nand3_1 _5566_ (.B(_1606_),
    .C(_1608_),
    .A(net1189),
    .Y(_1693_));
 sg13g2_nand3_1 _5567_ (.B(_1692_),
    .C(_1693_),
    .A(net1208),
    .Y(_1694_));
 sg13g2_nand2_1 _5568_ (.Y(_1695_),
    .A(_1600_),
    .B(_1612_));
 sg13g2_a22oi_1 _5569_ (.Y(_1696_),
    .B1(_1613_),
    .B2(_1695_),
    .A2(_1610_),
    .A1(net1212));
 sg13g2_a21o_1 _5570_ (.A2(_1696_),
    .A1(_1694_),
    .B1(net1185),
    .X(_1697_));
 sg13g2_nor2_2 _5571_ (.A(_1576_),
    .B(net1182),
    .Y(_1698_));
 sg13g2_a22oi_1 _5572_ (.Y(_1699_),
    .B1(_1695_),
    .B2(net1189),
    .A2(_1648_),
    .A1(_1608_));
 sg13g2_nand2b_1 _5573_ (.Y(_1700_),
    .B(net1179),
    .A_N(net1215));
 sg13g2_a21oi_1 _5574_ (.A1(_1698_),
    .A2(_1699_),
    .Y(_1701_),
    .B1(_1700_));
 sg13g2_nor2_2 _5575_ (.A(net1211),
    .B(net1181),
    .Y(_1702_));
 sg13g2_nand4_1 _5576_ (.B(net1189),
    .C(_1612_),
    .A(_1593_),
    .Y(_1703_),
    .D(_1633_));
 sg13g2_o21ai_1 _5577_ (.B1(_1703_),
    .Y(_1704_),
    .A1(net1190),
    .A2(_1600_));
 sg13g2_o21ai_1 _5578_ (.B1(_1702_),
    .Y(_1705_),
    .A1(_1664_),
    .A2(_1704_));
 sg13g2_nand3_1 _5579_ (.B(_1701_),
    .C(_1705_),
    .A(_1697_),
    .Y(_1706_));
 sg13g2_a21oi_1 _5580_ (.A1(_1633_),
    .A2(_1634_),
    .Y(_1707_),
    .B1(net1193));
 sg13g2_inv_1 _5581_ (.Y(_1708_),
    .A(_1707_));
 sg13g2_o21ai_1 _5582_ (.B1(_1702_),
    .Y(_1709_),
    .A1(_1632_),
    .A2(_1707_));
 sg13g2_o21ai_1 _5583_ (.B1(net1203),
    .Y(_1710_),
    .A1(net1199),
    .A2(net1196));
 sg13g2_and2_1 _5584_ (.A(_1648_),
    .B(_1710_),
    .X(_1711_));
 sg13g2_a21oi_1 _5585_ (.A1(_1599_),
    .A2(_1634_),
    .Y(_1712_),
    .B1(net1193));
 sg13g2_o21ai_1 _5586_ (.B1(_1698_),
    .Y(_1713_),
    .A1(_1711_),
    .A2(_1712_));
 sg13g2_nand2_1 _5587_ (.Y(_1714_),
    .A(net1187),
    .B(_1602_));
 sg13g2_a21oi_1 _5588_ (.A1(_1600_),
    .A2(_1683_),
    .Y(_1715_),
    .B1(net1184));
 sg13g2_o21ai_1 _5589_ (.B1(_1715_),
    .Y(_1716_),
    .A1(net1207),
    .A2(_1714_));
 sg13g2_nand4_1 _5590_ (.B(_1709_),
    .C(_1713_),
    .A(_1682_),
    .Y(_1717_),
    .D(_1716_));
 sg13g2_nor2_1 _5591_ (.A(net1209),
    .B(_1675_),
    .Y(_1718_));
 sg13g2_nor2b_2 _5592_ (.A(_1664_),
    .B_N(_1702_),
    .Y(_1719_));
 sg13g2_nand2_1 _5593_ (.Y(_1720_),
    .A(net1188),
    .B(_1710_));
 sg13g2_nand2_1 _5594_ (.Y(_1721_),
    .A(_1719_),
    .B(_1720_));
 sg13g2_o21ai_1 _5595_ (.B1(_1603_),
    .Y(_1722_),
    .A1(_1614_),
    .A2(_1615_));
 sg13g2_o21ai_1 _5596_ (.B1(net1181),
    .Y(_1723_),
    .A1(_1718_),
    .A2(_1722_));
 sg13g2_nand3_1 _5597_ (.B(_1721_),
    .C(_1723_),
    .A(_1654_),
    .Y(_1724_));
 sg13g2_xnor2_1 _5598_ (.Y(_1725_),
    .A(_1579_),
    .B(_1589_));
 sg13g2_a21oi_1 _5599_ (.A1(net1194),
    .A2(_1725_),
    .Y(_1726_),
    .B1(net1211));
 sg13g2_o21ai_1 _5600_ (.B1(_1726_),
    .Y(_1727_),
    .A1(_1592_),
    .A2(_1604_));
 sg13g2_a21oi_1 _5601_ (.A1(net1189),
    .A2(_1725_),
    .Y(_1728_),
    .B1(net1208));
 sg13g2_nand3_1 _5602_ (.B(_1608_),
    .C(_1728_),
    .A(_1606_),
    .Y(_1729_));
 sg13g2_nand3_1 _5603_ (.B(_1727_),
    .C(_1729_),
    .A(net1182),
    .Y(_1730_));
 sg13g2_a21oi_1 _5604_ (.A1(net1202),
    .A2(_1601_),
    .Y(_1731_),
    .B1(net1182));
 sg13g2_nand2_1 _5605_ (.Y(_1732_),
    .A(_1635_),
    .B(_1731_));
 sg13g2_and2_1 _5606_ (.A(net1215),
    .B(net1178),
    .X(_1733_));
 sg13g2_nand3_1 _5607_ (.B(_1732_),
    .C(_1733_),
    .A(_1730_),
    .Y(_1734_));
 sg13g2_nand4_1 _5608_ (.B(_1717_),
    .C(_1724_),
    .A(_1706_),
    .Y(_1735_),
    .D(_1734_));
 sg13g2_xnor2_1 _5609_ (.Y(_1736_),
    .A(net1239),
    .B(_1735_));
 sg13g2_xor2_1 _5610_ (.B(_1735_),
    .A(net1239),
    .X(_1737_));
 sg13g2_nand2_1 _5611_ (.Y(_1738_),
    .A(_1543_),
    .B(_1737_));
 sg13g2_nand2_1 _5612_ (.Y(_1739_),
    .A(net1252),
    .B(_1690_));
 sg13g2_nand3_1 _5613_ (.B(_1738_),
    .C(_1739_),
    .A(net1254),
    .Y(_1740_));
 sg13g2_nand2_1 _5614_ (.Y(_1741_),
    .A(net337),
    .B(_1534_));
 sg13g2_o21ai_1 _5615_ (.B1(_1741_),
    .Y(_0217_),
    .A1(net1278),
    .A2(_1740_));
 sg13g2_nand2_1 _5616_ (.Y(_1742_),
    .A(net1252),
    .B(_1736_));
 sg13g2_nand3_1 _5617_ (.B(_1599_),
    .C(_1634_),
    .A(net1193),
    .Y(_1743_));
 sg13g2_nor2b_1 _5618_ (.A(_1712_),
    .B_N(_1743_),
    .Y(_1744_));
 sg13g2_nor2_1 _5619_ (.A(net1182),
    .B(_1744_),
    .Y(_1745_));
 sg13g2_nand2b_1 _5620_ (.Y(_1746_),
    .B(net1189),
    .A_N(_1725_));
 sg13g2_nand3_1 _5621_ (.B(_1635_),
    .C(_1746_),
    .A(_1633_),
    .Y(_1747_));
 sg13g2_a21oi_1 _5622_ (.A1(_1634_),
    .A2(_1648_),
    .Y(_1748_),
    .B1(net1208));
 sg13g2_a221oi_1 _5623_ (.B2(_1708_),
    .C1(net1185),
    .B1(_1748_),
    .A1(_1638_),
    .Y(_1749_),
    .A2(_1747_));
 sg13g2_o21ai_1 _5624_ (.B1(_1733_),
    .Y(_1750_),
    .A1(_1745_),
    .A2(_1749_));
 sg13g2_nand2_1 _5625_ (.Y(_1751_),
    .A(net1191),
    .B(_1667_));
 sg13g2_nand2_1 _5626_ (.Y(_1752_),
    .A(_1660_),
    .B(_1751_));
 sg13g2_nand3_1 _5627_ (.B(_1675_),
    .C(_1683_),
    .A(_1603_),
    .Y(_1753_));
 sg13g2_nand3_1 _5628_ (.B(_1660_),
    .C(_1698_),
    .A(_1649_),
    .Y(_1754_));
 sg13g2_nand2_1 _5629_ (.Y(_1755_),
    .A(net1214),
    .B(_1754_));
 sg13g2_a221oi_1 _5630_ (.B2(net1181),
    .C1(_1755_),
    .B1(_1753_),
    .A1(_1719_),
    .Y(_1756_),
    .A2(_1752_));
 sg13g2_nor2_2 _5631_ (.A(net1213),
    .B(net1183),
    .Y(_1757_));
 sg13g2_o21ai_1 _5632_ (.B1(_1757_),
    .Y(_1758_),
    .A1(net1191),
    .A2(_1718_));
 sg13g2_nor2_1 _5633_ (.A(_1684_),
    .B(_1758_),
    .Y(_1759_));
 sg13g2_o21ai_1 _5634_ (.B1(_1631_),
    .Y(_1760_),
    .A1(_1756_),
    .A2(_1759_));
 sg13g2_nand3_1 _5635_ (.B(_1633_),
    .C(_1710_),
    .A(net1187),
    .Y(_1761_));
 sg13g2_nand3_1 _5636_ (.B(_1658_),
    .C(_1761_),
    .A(net1205),
    .Y(_1762_));
 sg13g2_or2_1 _5637_ (.X(_1763_),
    .B(_1761_),
    .A(net1205));
 sg13g2_nand2b_1 _5638_ (.Y(_1764_),
    .B(net1184),
    .A_N(net1214));
 sg13g2_a21oi_1 _5639_ (.A1(_1613_),
    .A2(_1634_),
    .Y(_1765_),
    .B1(_1764_));
 sg13g2_and3_1 _5640_ (.X(_1766_),
    .A(_1762_),
    .B(_1763_),
    .C(_1765_));
 sg13g2_nor3_1 _5641_ (.A(net1211),
    .B(_1707_),
    .C(_1711_),
    .Y(_1767_));
 sg13g2_a21oi_1 _5642_ (.A1(_1603_),
    .A2(_1675_),
    .Y(_1768_),
    .B1(_1614_));
 sg13g2_nand2_1 _5643_ (.Y(_1769_),
    .A(net1209),
    .B(_1603_));
 sg13g2_o21ai_1 _5644_ (.B1(_1757_),
    .Y(_1770_),
    .A1(_1656_),
    .A2(_1769_));
 sg13g2_nor3_1 _5645_ (.A(_1767_),
    .B(_1768_),
    .C(_1770_),
    .Y(_1771_));
 sg13g2_o21ai_1 _5646_ (.B1(net1178),
    .Y(_1772_),
    .A1(_1766_),
    .A2(_1771_));
 sg13g2_nand4_1 _5647_ (.B(_1654_),
    .C(_1702_),
    .A(net1188),
    .Y(_1773_),
    .D(_1710_));
 sg13g2_nand4_1 _5648_ (.B(_1760_),
    .C(_1772_),
    .A(_1750_),
    .Y(_1774_),
    .D(_1773_));
 sg13g2_xor2_1 _5649_ (.B(_1774_),
    .A(net1238),
    .X(_1775_));
 sg13g2_xnor2_1 _5650_ (.Y(_1776_),
    .A(net1238),
    .B(_1774_));
 sg13g2_o21ai_1 _5651_ (.B1(_1742_),
    .Y(_1777_),
    .A1(net1252),
    .A2(_1776_));
 sg13g2_nor2_1 _5652_ (.A(net1254),
    .B(net1252),
    .Y(_1778_));
 sg13g2_a22oi_1 _5653_ (.Y(_1779_),
    .B1(_1778_),
    .B2(_1691_),
    .A2(_1777_),
    .A1(net1254));
 sg13g2_nand2_1 _5654_ (.Y(_1780_),
    .A(net325),
    .B(net1278));
 sg13g2_o21ai_1 _5655_ (.B1(_1780_),
    .Y(_0218_),
    .A1(net1278),
    .A2(_1779_));
 sg13g2_a22oi_1 _5656_ (.Y(_1781_),
    .B1(_1710_),
    .B2(net1187),
    .A2(_1675_),
    .A1(_1648_));
 sg13g2_o21ai_1 _5657_ (.B1(net1209),
    .Y(_1782_),
    .A1(net1200),
    .A2(net1191));
 sg13g2_a21oi_1 _5658_ (.A1(net1205),
    .A2(_1781_),
    .Y(_1783_),
    .B1(net1183));
 sg13g2_o21ai_1 _5659_ (.B1(_1783_),
    .Y(_1784_),
    .A1(_1781_),
    .A2(_1782_));
 sg13g2_a21oi_1 _5660_ (.A1(_1675_),
    .A2(_1752_),
    .Y(_1785_),
    .B1(_1698_));
 sg13g2_a221oi_1 _5661_ (.B2(_1751_),
    .C1(_1674_),
    .B1(_1660_),
    .A1(net1207),
    .Y(_1786_),
    .A2(net1184));
 sg13g2_o21ai_1 _5662_ (.B1(_1784_),
    .Y(_1787_),
    .A1(_1785_),
    .A2(_1786_));
 sg13g2_nor4_1 _5663_ (.A(net1214),
    .B(_1613_),
    .C(net1184),
    .D(net1178),
    .Y(_1788_));
 sg13g2_a21oi_1 _5664_ (.A1(net1191),
    .A2(_1603_),
    .Y(_1789_),
    .B1(net1183));
 sg13g2_a22oi_1 _5665_ (.Y(_1790_),
    .B1(_1789_),
    .B2(_1714_),
    .A2(_1719_),
    .A1(_1660_));
 sg13g2_a22oi_1 _5666_ (.Y(_1791_),
    .B1(_1790_),
    .B2(_1682_),
    .A2(_1788_),
    .A1(_1678_));
 sg13g2_a21oi_1 _5667_ (.A1(_1648_),
    .A2(_1698_),
    .Y(_1792_),
    .B1(_1791_));
 sg13g2_a21oi_1 _5668_ (.A1(net1203),
    .A2(net1193),
    .Y(_1793_),
    .B1(net1205));
 sg13g2_o21ai_1 _5669_ (.B1(_1633_),
    .Y(_1794_),
    .A1(net1187),
    .A2(_1615_));
 sg13g2_a221oi_1 _5670_ (.B2(net1205),
    .C1(_1764_),
    .B1(_1794_),
    .A1(_1720_),
    .Y(_1795_),
    .A2(_1793_));
 sg13g2_a21oi_1 _5671_ (.A1(_1649_),
    .A2(_1660_),
    .Y(_1796_),
    .B1(net1209));
 sg13g2_a21oi_1 _5672_ (.A1(net1191),
    .A2(_1603_),
    .Y(_1797_),
    .B1(_1669_));
 sg13g2_o21ai_1 _5673_ (.B1(_1757_),
    .Y(_1798_),
    .A1(_1796_),
    .A2(_1797_));
 sg13g2_nand2b_1 _5674_ (.Y(_1799_),
    .B(_1798_),
    .A_N(_1795_));
 sg13g2_a221oi_1 _5675_ (.B2(net1178),
    .C1(_1792_),
    .B1(_1799_),
    .A1(_1733_),
    .Y(_1800_),
    .A2(_1787_));
 sg13g2_xnor2_1 _5676_ (.Y(_1801_),
    .A(net1238),
    .B(_1800_));
 sg13g2_xor2_1 _5677_ (.B(_1800_),
    .A(net1239),
    .X(_1802_));
 sg13g2_mux2_1 _5678_ (.A0(_1775_),
    .A1(_1801_),
    .S(_1543_),
    .X(_1803_));
 sg13g2_mux4_1 _5679_ (.S0(_1543_),
    .A0(_1690_),
    .A1(_1737_),
    .A2(_1776_),
    .A3(_1802_),
    .S1(net1254),
    .X(_1804_));
 sg13g2_nand2_1 _5680_ (.Y(_1805_),
    .A(net332),
    .B(net1278));
 sg13g2_o21ai_1 _5681_ (.B1(_1805_),
    .Y(_0219_),
    .A1(net1276),
    .A2(_1804_));
 sg13g2_a21oi_1 _5682_ (.A1(net1210),
    .A2(_1656_),
    .Y(_1806_),
    .B1(net1183));
 sg13g2_nor2_1 _5683_ (.A(net1213),
    .B(_1806_),
    .Y(_1807_));
 sg13g2_o21ai_1 _5684_ (.B1(net1180),
    .Y(_1808_),
    .A1(net1213),
    .A2(_1806_));
 sg13g2_nor3_1 _5685_ (.A(net1214),
    .B(net1210),
    .C(_1648_),
    .Y(_1809_));
 sg13g2_nor2_1 _5686_ (.A(net1181),
    .B(_1793_),
    .Y(_1810_));
 sg13g2_nand4_1 _5687_ (.B(_1661_),
    .C(_1683_),
    .A(net1178),
    .Y(_1811_),
    .D(_1810_));
 sg13g2_o21ai_1 _5688_ (.B1(_1811_),
    .Y(_1812_),
    .A1(_1808_),
    .A2(_1809_));
 sg13g2_or2_1 _5689_ (.X(_1813_),
    .B(_1675_),
    .A(_1614_));
 sg13g2_a21oi_1 _5690_ (.A1(net1200),
    .A2(net1187),
    .Y(_1814_),
    .B1(net1206));
 sg13g2_a21o_1 _5691_ (.A2(_1649_),
    .A1(net1206),
    .B1(_1814_),
    .X(_1815_));
 sg13g2_nand3_1 _5692_ (.B(net1192),
    .C(_1667_),
    .A(net1206),
    .Y(_1816_));
 sg13g2_nand4_1 _5693_ (.B(_1813_),
    .C(_1815_),
    .A(net1183),
    .Y(_1817_),
    .D(_1816_));
 sg13g2_a21o_1 _5694_ (.A2(_1815_),
    .A1(_1813_),
    .B1(net1183),
    .X(_1818_));
 sg13g2_nand3_1 _5695_ (.B(_1817_),
    .C(_1818_),
    .A(net1213),
    .Y(_1819_));
 sg13g2_nand2_1 _5696_ (.Y(_1820_),
    .A(net1205),
    .B(_1789_));
 sg13g2_nor3_1 _5697_ (.A(_1602_),
    .B(_1614_),
    .C(net1184),
    .Y(_1821_));
 sg13g2_nor2_1 _5698_ (.A(_1719_),
    .B(_1821_),
    .Y(_1822_));
 sg13g2_nand3_1 _5699_ (.B(_1820_),
    .C(_1822_),
    .A(net1213),
    .Y(_1823_));
 sg13g2_a21oi_1 _5700_ (.A1(_1677_),
    .A2(_1757_),
    .Y(_1824_),
    .B1(net1178));
 sg13g2_a22oi_1 _5701_ (.Y(_1825_),
    .B1(_1823_),
    .B2(_1824_),
    .A2(_1819_),
    .A1(_1812_));
 sg13g2_xor2_1 _5702_ (.B(_1825_),
    .A(net1238),
    .X(_1826_));
 sg13g2_and2_1 _5703_ (.A(_1543_),
    .B(_1826_),
    .X(_1827_));
 sg13g2_a21oi_1 _5704_ (.A1(net1252),
    .A2(_1801_),
    .Y(_1828_),
    .B1(_1827_));
 sg13g2_nand2_1 _5705_ (.Y(_1829_),
    .A(net1253),
    .B(_1828_));
 sg13g2_o21ai_1 _5706_ (.B1(_1829_),
    .Y(_1830_),
    .A1(net1254),
    .A2(_1777_));
 sg13g2_mux4_1 _5707_ (.S0(_1543_),
    .A0(_1736_),
    .A1(_1775_),
    .A2(_1801_),
    .A3(_1826_),
    .S1(net1253),
    .X(_1831_));
 sg13g2_nand2_1 _5708_ (.Y(_1832_),
    .A(net328),
    .B(net1278));
 sg13g2_o21ai_1 _5709_ (.B1(_1832_),
    .Y(_0220_),
    .A1(_1534_),
    .A2(_1830_));
 sg13g2_a21oi_1 _5710_ (.A1(net1191),
    .A2(_1667_),
    .Y(_1833_),
    .B1(net1210));
 sg13g2_a221oi_1 _5711_ (.B2(net1206),
    .C1(net1181),
    .B1(_1751_),
    .A1(_1613_),
    .Y(_1834_),
    .A2(_1674_));
 sg13g2_nor2_1 _5712_ (.A(net1183),
    .B(_1814_),
    .Y(_1835_));
 sg13g2_o21ai_1 _5713_ (.B1(_1733_),
    .Y(_1836_),
    .A1(_1834_),
    .A2(_1835_));
 sg13g2_a21oi_1 _5714_ (.A1(net1213),
    .A2(_1820_),
    .Y(_1837_),
    .B1(net1179));
 sg13g2_o21ai_1 _5715_ (.B1(_1808_),
    .Y(_1838_),
    .A1(net1181),
    .A2(_1665_));
 sg13g2_o21ai_1 _5716_ (.B1(_1836_),
    .Y(_1839_),
    .A1(_1837_),
    .A2(_1838_));
 sg13g2_xor2_1 _5717_ (.B(_1839_),
    .A(net1238),
    .X(_1840_));
 sg13g2_mux2_1 _5718_ (.A0(_1826_),
    .A1(_1840_),
    .S(_1543_),
    .X(_1841_));
 sg13g2_nand2b_1 _5719_ (.Y(_1842_),
    .B(net1253),
    .A_N(_1841_));
 sg13g2_o21ai_1 _5720_ (.B1(_1842_),
    .Y(_1843_),
    .A1(net1253),
    .A2(_1803_));
 sg13g2_nand2_1 _5721_ (.Y(_1844_),
    .A(net327),
    .B(net1276));
 sg13g2_o21ai_1 _5722_ (.B1(_1844_),
    .Y(_0221_),
    .A1(net1276),
    .A2(_1843_));
 sg13g2_nor2_1 _5723_ (.A(net1253),
    .B(_1828_),
    .Y(_1845_));
 sg13g2_o21ai_1 _5724_ (.B1(net1213),
    .Y(_1846_),
    .A1(net1181),
    .A2(_1833_));
 sg13g2_a21oi_1 _5725_ (.A1(_1631_),
    .A2(_1820_),
    .Y(_1847_),
    .B1(_1846_));
 sg13g2_o21ai_1 _5726_ (.B1(_1655_),
    .Y(_1848_),
    .A1(_1807_),
    .A2(_1847_));
 sg13g2_xnor2_1 _5727_ (.Y(_1849_),
    .A(net1238),
    .B(_1848_));
 sg13g2_mux2_1 _5728_ (.A0(_1840_),
    .A1(_1849_),
    .S(_1543_),
    .X(_1850_));
 sg13g2_a21oi_2 _5729_ (.B1(_1845_),
    .Y(_1851_),
    .A2(_1850_),
    .A1(net1253));
 sg13g2_nand2_1 _5730_ (.Y(_1852_),
    .A(net326),
    .B(net1276));
 sg13g2_o21ai_1 _5731_ (.B1(_1852_),
    .Y(_0222_),
    .A1(net1276),
    .A2(_1851_));
 sg13g2_xor2_1 _5732_ (.B(_1808_),
    .A(net1238),
    .X(_1853_));
 sg13g2_nor2_1 _5733_ (.A(net1252),
    .B(_1853_),
    .Y(_1854_));
 sg13g2_a21oi_2 _5734_ (.B1(_1854_),
    .Y(_1855_),
    .A2(_1849_),
    .A1(net1252));
 sg13g2_nand2_1 _5735_ (.Y(_1856_),
    .A(net1253),
    .B(_1855_));
 sg13g2_o21ai_1 _5736_ (.B1(_1856_),
    .Y(_1857_),
    .A1(net1253),
    .A2(_1841_));
 sg13g2_nand2_1 _5737_ (.Y(_1858_),
    .A(net340),
    .B(net1277));
 sg13g2_o21ai_1 _5738_ (.B1(_1858_),
    .Y(_0223_),
    .A1(net1276),
    .A2(_1857_));
 sg13g2_mux2_1 _5739_ (.A0(net1241),
    .A1(_1853_),
    .S(_1542_),
    .X(_1859_));
 sg13g2_nand2_1 _5740_ (.Y(_1860_),
    .A(net1255),
    .B(_1859_));
 sg13g2_o21ai_1 _5741_ (.B1(_1860_),
    .Y(_1861_),
    .A1(net1255),
    .A2(_1850_));
 sg13g2_nand2_1 _5742_ (.Y(_1862_),
    .A(net331),
    .B(net1277));
 sg13g2_o21ai_1 _5743_ (.B1(_1862_),
    .Y(_0224_),
    .A1(net1277),
    .A2(_1861_));
 sg13g2_mux2_2 _5744_ (.A0(_1855_),
    .A1(net1241),
    .S(net1255),
    .X(_1863_));
 sg13g2_nand2_1 _5745_ (.Y(_1864_),
    .A(net333),
    .B(net1277));
 sg13g2_o21ai_1 _5746_ (.B1(_1864_),
    .Y(_0225_),
    .A1(net1277),
    .A2(_1863_));
 sg13g2_a21oi_1 _5747_ (.A1(_1549_),
    .A2(_1557_),
    .Y(_1865_),
    .B1(net1278));
 sg13g2_a21oi_1 _5748_ (.A1(_3173_),
    .A2(net1276),
    .Y(_0226_),
    .B1(_1865_));
 sg13g2_a21oi_1 _5749_ (.A1(_3175_),
    .A2(net1276),
    .Y(_0227_),
    .B1(_1865_));
 sg13g2_nand4_1 _5750_ (.B(_3138_),
    .C(_0093_),
    .A(net1388),
    .Y(_1866_),
    .D(net1296));
 sg13g2_nand2_1 _5751_ (.Y(_1867_),
    .A(net341),
    .B(net1269));
 sg13g2_o21ai_1 _5752_ (.B1(_1867_),
    .Y(_0228_),
    .A1(_1740_),
    .A2(net1269));
 sg13g2_nand2_1 _5753_ (.Y(_1868_),
    .A(net348),
    .B(net1269));
 sg13g2_o21ai_1 _5754_ (.B1(_1868_),
    .Y(_0229_),
    .A1(_1779_),
    .A2(net1269));
 sg13g2_nand2_1 _5755_ (.Y(_1869_),
    .A(net395),
    .B(net1269));
 sg13g2_o21ai_1 _5756_ (.B1(_1869_),
    .Y(_0230_),
    .A1(_1804_),
    .A2(net1268));
 sg13g2_nor2_1 _5757_ (.A(_1831_),
    .B(net1268),
    .Y(_1870_));
 sg13g2_a21oi_1 _5758_ (.A1(_3168_),
    .A2(net1269),
    .Y(_0231_),
    .B1(_1870_));
 sg13g2_nand2_1 _5759_ (.Y(_1871_),
    .A(net353),
    .B(net1268));
 sg13g2_o21ai_1 _5760_ (.B1(_1871_),
    .Y(_0232_),
    .A1(_1843_),
    .A2(net1268));
 sg13g2_nand2_1 _5761_ (.Y(_1872_),
    .A(net346),
    .B(net1268));
 sg13g2_o21ai_1 _5762_ (.B1(_1872_),
    .Y(_0233_),
    .A1(_1851_),
    .A2(net1268));
 sg13g2_nand2_1 _5763_ (.Y(_1873_),
    .A(net422),
    .B(net1267));
 sg13g2_o21ai_1 _5764_ (.B1(_1873_),
    .Y(_0234_),
    .A1(_1857_),
    .A2(net1267));
 sg13g2_nand2_1 _5765_ (.Y(_1874_),
    .A(net388),
    .B(net1267));
 sg13g2_o21ai_1 _5766_ (.B1(_1874_),
    .Y(_0235_),
    .A1(_1861_),
    .A2(net1267));
 sg13g2_nand2_1 _5767_ (.Y(_1875_),
    .A(net367),
    .B(net1267));
 sg13g2_o21ai_1 _5768_ (.B1(_1875_),
    .Y(_0236_),
    .A1(_1863_),
    .A2(net1267));
 sg13g2_mux2_1 _5769_ (.A0(_1859_),
    .A1(net1241),
    .S(net1255),
    .X(_1876_));
 sg13g2_nand2_1 _5770_ (.Y(_1877_),
    .A(net357),
    .B(net1267));
 sg13g2_o21ai_1 _5771_ (.B1(_1877_),
    .Y(_0237_),
    .A1(net1267),
    .A2(_1876_));
 sg13g2_nand2_1 _5772_ (.Y(_1878_),
    .A(net399),
    .B(net1269));
 sg13g2_o21ai_1 _5773_ (.B1(_1878_),
    .Y(_0238_),
    .A1(_1558_),
    .A2(net1268));
 sg13g2_nor2b_2 _5774_ (.A(net1388),
    .B_N(net1382),
    .Y(_1879_));
 sg13g2_nand2_1 _5775_ (.Y(_1880_),
    .A(net1296),
    .B(_1879_));
 sg13g2_nand3_1 _5776_ (.B(net1296),
    .C(_1879_),
    .A(_0093_),
    .Y(_1881_));
 sg13g2_inv_1 _5777_ (.Y(_1882_),
    .A(net1265));
 sg13g2_nand2_1 _5778_ (.Y(_1883_),
    .A(net429),
    .B(net1266));
 sg13g2_o21ai_1 _5779_ (.B1(_1883_),
    .Y(_0239_),
    .A1(_1740_),
    .A2(net1266));
 sg13g2_nand2_1 _5780_ (.Y(_1884_),
    .A(net373),
    .B(net1266));
 sg13g2_o21ai_1 _5781_ (.B1(_1884_),
    .Y(_0240_),
    .A1(_1779_),
    .A2(net1266));
 sg13g2_nand2_1 _5782_ (.Y(_1885_),
    .A(net363),
    .B(net1266));
 sg13g2_o21ai_1 _5783_ (.B1(_1885_),
    .Y(_0241_),
    .A1(_1804_),
    .A2(_1881_));
 sg13g2_nand2_1 _5784_ (.Y(_1886_),
    .A(net433),
    .B(net1266));
 sg13g2_o21ai_1 _5785_ (.B1(_1886_),
    .Y(_0242_),
    .A1(_1830_),
    .A2(net1266));
 sg13g2_nand2_1 _5786_ (.Y(_1887_),
    .A(net358),
    .B(net1265));
 sg13g2_o21ai_1 _5787_ (.B1(_1887_),
    .Y(_0243_),
    .A1(_1843_),
    .A2(net1265));
 sg13g2_nand2_1 _5788_ (.Y(_1888_),
    .A(net362),
    .B(net1265));
 sg13g2_o21ai_1 _5789_ (.B1(_1888_),
    .Y(_0244_),
    .A1(_1851_),
    .A2(net1265));
 sg13g2_nand2_1 _5790_ (.Y(_1889_),
    .A(net379),
    .B(net1264));
 sg13g2_o21ai_1 _5791_ (.B1(_1889_),
    .Y(_0245_),
    .A1(_1857_),
    .A2(net1264));
 sg13g2_nand2_1 _5792_ (.Y(_1890_),
    .A(net382),
    .B(net1264));
 sg13g2_o21ai_1 _5793_ (.B1(_1890_),
    .Y(_0246_),
    .A1(_1861_),
    .A2(net1264));
 sg13g2_nand2_1 _5794_ (.Y(_1891_),
    .A(net361),
    .B(net1264));
 sg13g2_o21ai_1 _5795_ (.B1(_1891_),
    .Y(_0247_),
    .A1(_1863_),
    .A2(net1264));
 sg13g2_nand2_1 _5796_ (.Y(_1892_),
    .A(net364),
    .B(net1264));
 sg13g2_o21ai_1 _5797_ (.B1(_1892_),
    .Y(_0248_),
    .A1(net1241),
    .A2(net1264));
 sg13g2_nor2_1 _5798_ (.A(net502),
    .B(_1882_),
    .Y(_1893_));
 sg13g2_a21oi_1 _5799_ (.A1(_1558_),
    .A2(_1882_),
    .Y(_0249_),
    .B1(_1893_));
 sg13g2_and2_1 _5800_ (.A(_1215_),
    .B(_1440_),
    .X(_1894_));
 sg13g2_nor2_1 _5801_ (.A(net1170),
    .B(net1168),
    .Y(_1895_));
 sg13g2_nor2_1 _5802_ (.A(net1403),
    .B(\dtop.ext_control[1] ),
    .Y(_1896_));
 sg13g2_o21ai_1 _5803_ (.B1(net1344),
    .Y(_1897_),
    .A1(_3327_),
    .A2(_1896_));
 sg13g2_a221oi_1 _5804_ (.B2(net1170),
    .C1(_1440_),
    .B1(_1897_),
    .A1(_1137_),
    .Y(_1898_),
    .A2(_1895_));
 sg13g2_a21oi_1 _5805_ (.A1(net1300),
    .A2(_1264_),
    .Y(_1899_),
    .B1(_1167_));
 sg13g2_nor2_1 _5806_ (.A(_0983_),
    .B(_1169_),
    .Y(_1900_));
 sg13g2_nor2_1 _5807_ (.A(_1899_),
    .B(_1900_),
    .Y(_1901_));
 sg13g2_a21oi_1 _5808_ (.A1(_1192_),
    .A2(_1244_),
    .Y(_1902_),
    .B1(_0733_));
 sg13g2_o21ai_1 _5809_ (.B1(_1902_),
    .Y(_1903_),
    .A1(_1192_),
    .A2(_1249_));
 sg13g2_inv_1 _5810_ (.Y(_1904_),
    .A(_1903_));
 sg13g2_nand2_2 _5811_ (.Y(_1905_),
    .A(\dtop.ext_control[0] ),
    .B(net1282));
 sg13g2_nand2b_1 _5812_ (.Y(_1906_),
    .B(_3326_),
    .A_N(\dtop.ext_control[2] ));
 sg13g2_nand2_1 _5813_ (.Y(_1907_),
    .A(_1905_),
    .B(_1906_));
 sg13g2_o21ai_1 _5814_ (.B1(_1043_),
    .Y(_1908_),
    .A1(_1903_),
    .A2(_1907_));
 sg13g2_o21ai_1 _5815_ (.B1(_1908_),
    .Y(_1909_),
    .A1(_0020_),
    .A2(_0982_));
 sg13g2_a21oi_1 _5816_ (.A1(_1895_),
    .A2(_1901_),
    .Y(_1910_),
    .B1(_1909_));
 sg13g2_a22oi_1 _5817_ (.Y(_1911_),
    .B1(_1898_),
    .B2(_1910_),
    .A2(_1894_),
    .A1(_1174_));
 sg13g2_nand2_1 _5818_ (.Y(_1912_),
    .A(net1300),
    .B(_1249_));
 sg13g2_or2_1 _5819_ (.X(_1913_),
    .B(_1244_),
    .A(_0733_));
 sg13g2_o21ai_1 _5820_ (.B1(_1913_),
    .Y(_1914_),
    .A1(_1193_),
    .A2(_1197_));
 sg13g2_nand2_1 _5821_ (.Y(_1915_),
    .A(_3321_),
    .B(_1187_));
 sg13g2_xor2_1 _5822_ (.B(_1915_),
    .A(_1914_),
    .X(_1916_));
 sg13g2_a22oi_1 _5823_ (.Y(_1917_),
    .B1(_1916_),
    .B2(_1192_),
    .A2(_1912_),
    .A1(_1194_));
 sg13g2_nor3_1 _5824_ (.A(_1904_),
    .B(_1906_),
    .C(_1917_),
    .Y(_1918_));
 sg13g2_a21oi_1 _5825_ (.A1(_1905_),
    .A2(_1918_),
    .Y(_1919_),
    .B1(_1908_));
 sg13g2_nand2b_1 _5826_ (.Y(_1920_),
    .B(_1895_),
    .A_N(_1901_));
 sg13g2_nand2b_1 _5827_ (.Y(_1921_),
    .B(net1170),
    .A_N(_0021_));
 sg13g2_nand3_1 _5828_ (.B(_1920_),
    .C(_1921_),
    .A(_1898_),
    .Y(_1922_));
 sg13g2_nand2_1 _5829_ (.Y(_1923_),
    .A(_1175_),
    .B(_1894_));
 sg13g2_o21ai_1 _5830_ (.B1(_1923_),
    .Y(_1924_),
    .A1(_1919_),
    .A2(_1922_));
 sg13g2_and2_1 _5831_ (.A(_1292_),
    .B(_1924_),
    .X(_1925_));
 sg13g2_o21ai_1 _5832_ (.B1(_1917_),
    .Y(_1926_),
    .A1(_1903_),
    .A2(_1906_));
 sg13g2_nand2_1 _5833_ (.Y(_1927_),
    .A(_1905_),
    .B(_1926_));
 sg13g2_nand2_1 _5834_ (.Y(_1928_),
    .A(net1168),
    .B(_1927_));
 sg13g2_a21oi_2 _5835_ (.B1(_1894_),
    .Y(_1929_),
    .A2(_1928_),
    .A1(_1898_));
 sg13g2_nand4_1 _5836_ (.B(_1006_),
    .C(_1007_),
    .A(_0778_),
    .Y(_1930_),
    .D(_1476_));
 sg13g2_a21oi_1 _5837_ (.A1(_0923_),
    .A2(_1069_),
    .Y(_1931_),
    .B1(_1924_));
 sg13g2_nor2_1 _5838_ (.A(_1911_),
    .B(_1931_),
    .Y(_1932_));
 sg13g2_a21oi_1 _5839_ (.A1(_1109_),
    .A2(_1122_),
    .Y(_1933_),
    .B1(_1924_));
 sg13g2_o21ai_1 _5840_ (.B1(_1924_),
    .Y(_1934_),
    .A1(_1079_),
    .A2(_1096_));
 sg13g2_nand2_1 _5841_ (.Y(_1935_),
    .A(_1911_),
    .B(_1934_));
 sg13g2_nor2_1 _5842_ (.A(_1933_),
    .B(_1935_),
    .Y(_1936_));
 sg13g2_nor3_1 _5843_ (.A(_1929_),
    .B(_1932_),
    .C(_1936_),
    .Y(_1937_));
 sg13g2_nor2_1 _5844_ (.A(_1322_),
    .B(_1924_),
    .Y(_1938_));
 sg13g2_a22oi_1 _5845_ (.Y(_1939_),
    .B1(_1938_),
    .B2(_1307_),
    .A2(_1925_),
    .A1(_1134_));
 sg13g2_o21ai_1 _5846_ (.B1(_1929_),
    .Y(_1940_),
    .A1(_1911_),
    .A2(_1939_));
 sg13g2_nor2_1 _5847_ (.A(_1930_),
    .B(_1937_),
    .Y(_1941_));
 sg13g2_a22oi_1 _5848_ (.Y(_1942_),
    .B1(_1940_),
    .B2(_1941_),
    .A2(_1930_),
    .A1(net439));
 sg13g2_inv_1 _5849_ (.Y(_0250_),
    .A(_1942_));
 sg13g2_xnor2_1 _5850_ (.Y(_1943_),
    .A(net1393),
    .B(_1498_));
 sg13g2_nor3_1 _5851_ (.A(_3144_),
    .B(_0561_),
    .C(net707),
    .Y(_0251_));
 sg13g2_nor3_1 _5852_ (.A(_0085_),
    .B(\dtop.vtop.rs.x_scan.phase[0] ),
    .C(_3149_),
    .Y(_1944_));
 sg13g2_o21ai_1 _5853_ (.B1(_3140_),
    .Y(_1945_),
    .A1(net1368),
    .A2(\dtop.vtop.rs.x_scan.phase[0] ));
 sg13g2_nand4_1 _5854_ (.B(net1443),
    .C(_3142_),
    .A(net1442),
    .Y(_1946_),
    .D(_0093_));
 sg13g2_o21ai_1 _5855_ (.B1(\dtop.vtop.rs.x_scan.phase[0] ),
    .Y(_1947_),
    .A1(net1368),
    .A2(_3149_));
 sg13g2_a22oi_1 _5856_ (.Y(_1948_),
    .B1(_1947_),
    .B2(net1376),
    .A2(_1946_),
    .A1(_3149_));
 sg13g2_nor3_1 _5857_ (.A(net1441),
    .B(net1443),
    .C(_0093_),
    .Y(_1949_));
 sg13g2_nor3_1 _5858_ (.A(net1373),
    .B(_3353_),
    .C(net1349),
    .Y(_1950_));
 sg13g2_a21oi_1 _5859_ (.A1(_0085_),
    .A2(_0001_),
    .Y(_1951_),
    .B1(_1944_));
 sg13g2_o21ai_1 _5860_ (.B1(_1951_),
    .Y(_1952_),
    .A1(_0001_),
    .A2(_0432_));
 sg13g2_nand2_1 _5861_ (.Y(_1953_),
    .A(_1945_),
    .B(_1950_));
 sg13g2_o21ai_1 _5862_ (.B1(_1948_),
    .Y(_1954_),
    .A1(_3149_),
    .A2(_1949_));
 sg13g2_nor3_2 _5863_ (.A(_1952_),
    .B(_1953_),
    .C(_1954_),
    .Y(_1955_));
 sg13g2_a21oi_1 _5864_ (.A1(_0432_),
    .A2(_1955_),
    .Y(_1956_),
    .B1(_0087_));
 sg13g2_nand2_1 _5865_ (.Y(_1957_),
    .A(net320),
    .B(_1956_));
 sg13g2_nand2b_1 _5866_ (.Y(_1958_),
    .B(\dtop.vtop.rs.scan_y.phase[1] ),
    .A_N(\dtop.vtop.rs.scan_y.phase[0] ));
 sg13g2_o21ai_1 _5867_ (.B1(net321),
    .Y(_0252_),
    .A1(_1956_),
    .A2(_1958_));
 sg13g2_o21ai_1 _5868_ (.B1(_3333_),
    .Y(_0253_),
    .A1(net1358),
    .A2(_3183_));
 sg13g2_and2_1 _5869_ (.A(\dtop.vtop.rs.scan_y.phase[1] ),
    .B(\dtop.vtop.rs.scan_y.phase[0] ),
    .X(_1959_));
 sg13g2_nor3_1 _5870_ (.A(_0082_),
    .B(_0080_),
    .C(_1959_),
    .Y(_1960_));
 sg13g2_nor3_1 _5871_ (.A(net1393),
    .B(_0055_),
    .C(_0064_),
    .Y(_1961_));
 sg13g2_nand3_1 _5872_ (.B(_0055_),
    .C(_0064_),
    .A(net1393),
    .Y(_1962_));
 sg13g2_nand3_1 _5873_ (.B(_0080_),
    .C(_1959_),
    .A(net1426),
    .Y(_1963_));
 sg13g2_nor2_1 _5874_ (.A(_1962_),
    .B(_1963_),
    .Y(_1964_));
 sg13g2_a21oi_1 _5875_ (.A1(_1960_),
    .A2(_1961_),
    .Y(_1965_),
    .B1(_1964_));
 sg13g2_xnor2_1 _5876_ (.Y(_1966_),
    .A(_0081_),
    .B(\dtop.vtop.rs.scan_y.phase[0] ));
 sg13g2_o21ai_1 _5877_ (.B1(net1423),
    .Y(_1967_),
    .A1(\dtop.vtop.rs.scan_y.phase[1] ),
    .A2(\dtop.vtop.rs.scan_y.phase[0] ));
 sg13g2_nand3_1 _5878_ (.B(_1966_),
    .C(_1967_),
    .A(net1425),
    .Y(_1968_));
 sg13g2_nor2b_1 _5879_ (.A(_3208_),
    .B_N(net1417),
    .Y(_1969_));
 sg13g2_nand2b_1 _5880_ (.Y(_1970_),
    .B(_0082_),
    .A_N(net1418));
 sg13g2_nand2b_2 _5881_ (.Y(_1971_),
    .B(net1423),
    .A_N(net1417));
 sg13g2_nand3_1 _5882_ (.B(_1970_),
    .C(_1971_),
    .A(net1426),
    .Y(_1972_));
 sg13g2_o21ai_1 _5883_ (.B1(_1972_),
    .Y(_1973_),
    .A1(net1426),
    .A2(_1969_));
 sg13g2_nor4_1 _5884_ (.A(_0555_),
    .B(_1965_),
    .C(_1968_),
    .D(_1973_),
    .Y(_1974_));
 sg13g2_nor2_1 _5885_ (.A(net650),
    .B(_1974_),
    .Y(_1975_));
 sg13g2_and2_1 _5886_ (.A(net650),
    .B(_1974_),
    .X(_1976_));
 sg13g2_nor3_1 _5887_ (.A(_3144_),
    .B(net651),
    .C(_1976_),
    .Y(_0254_));
 sg13g2_o21ai_1 _5888_ (.B1(net1430),
    .Y(_1977_),
    .A1(net604),
    .A2(_1976_));
 sg13g2_a21oi_1 _5889_ (.A1(net604),
    .A2(_1976_),
    .Y(_0255_),
    .B1(_1977_));
 sg13g2_or2_1 _5890_ (.X(_1978_),
    .B(_1955_),
    .A(\dtop.vtop.rs.x_scan.phase[0] ));
 sg13g2_nand2_1 _5891_ (.Y(_1979_),
    .A(\dtop.vtop.rs.x_scan.phase[0] ),
    .B(_1955_));
 sg13g2_and3_1 _5892_ (.X(_0256_),
    .A(net1430),
    .B(_1978_),
    .C(_1979_));
 sg13g2_o21ai_1 _5893_ (.B1(net1430),
    .Y(_1980_),
    .A1(net634),
    .A2(_1979_));
 sg13g2_a21o_1 _5894_ (.A2(_1979_),
    .A1(net634),
    .B1(_1980_),
    .X(_0257_));
 sg13g2_nand2b_2 _5895_ (.Y(_1981_),
    .B(_3191_),
    .A_N(_0087_));
 sg13g2_nand2_2 _5896_ (.Y(_1982_),
    .A(net1391),
    .B(net1362));
 sg13g2_xnor2_1 _5897_ (.Y(_1983_),
    .A(net1392),
    .B(net1362));
 sg13g2_nor2_1 _5898_ (.A(_1981_),
    .B(net678),
    .Y(_0258_));
 sg13g2_xor2_1 _5899_ (.B(_1982_),
    .A(net1388),
    .X(_1984_));
 sg13g2_nor2_1 _5900_ (.A(_1981_),
    .B(_1984_),
    .Y(_0259_));
 sg13g2_nor2_2 _5901_ (.A(_0003_),
    .B(_1982_),
    .Y(_1985_));
 sg13g2_xnor2_1 _5902_ (.Y(_1986_),
    .A(net1382),
    .B(_1985_));
 sg13g2_nor2_1 _5903_ (.A(_1981_),
    .B(_1986_),
    .Y(_0260_));
 sg13g2_nor4_1 _5904_ (.A(_3137_),
    .B(_0001_),
    .C(_0003_),
    .D(_1982_),
    .Y(_1987_));
 sg13g2_a21oi_1 _5905_ (.A1(_3150_),
    .A2(_1985_),
    .Y(_1988_),
    .B1(net1379));
 sg13g2_nor3_1 _5906_ (.A(_1981_),
    .B(_1987_),
    .C(_1988_),
    .Y(_0261_));
 sg13g2_nor4_2 _5907_ (.A(_3140_),
    .B(_0003_),
    .C(net1333),
    .Y(_1989_),
    .D(_1982_));
 sg13g2_a21oi_1 _5908_ (.A1(_0613_),
    .A2(_1985_),
    .Y(_1990_),
    .B1(net1376));
 sg13g2_nor3_1 _5909_ (.A(_1981_),
    .B(_1989_),
    .C(_1990_),
    .Y(_0262_));
 sg13g2_nand2_1 _5910_ (.Y(_1991_),
    .A(net1373),
    .B(_1989_));
 sg13g2_xnor2_1 _5911_ (.Y(_1992_),
    .A(net1373),
    .B(_1989_));
 sg13g2_nor2_1 _5912_ (.A(_1981_),
    .B(_1992_),
    .Y(_0263_));
 sg13g2_xnor2_1 _5913_ (.Y(_1993_),
    .A(_3139_),
    .B(_1991_));
 sg13g2_nor2_1 _5914_ (.A(_1981_),
    .B(_1993_),
    .Y(_0264_));
 sg13g2_nor2_1 _5915_ (.A(_3065_),
    .B(net1355),
    .Y(_1994_));
 sg13g2_nand2b_1 _5916_ (.Y(_1995_),
    .B(\dtop.vtop.pipeline.z[14] ),
    .A_N(net1355));
 sg13g2_nand2b_1 _5917_ (.Y(_1996_),
    .B(\dtop.vtop.pipeline.z[9] ),
    .A_N(\dtop.vtop.pipeline.zg[4] ));
 sg13g2_nand2b_1 _5918_ (.Y(_1997_),
    .B(\dtop.vtop.pipeline.z[6] ),
    .A_N(\dtop.vtop.pipeline.zg[1] ));
 sg13g2_nor2b_1 _5919_ (.A(\dtop.vtop.pipeline.z[5] ),
    .B_N(\dtop.vtop.pipeline.zg[0] ),
    .Y(_1998_));
 sg13g2_nor2b_1 _5920_ (.A(\dtop.vtop.pipeline.z[6] ),
    .B_N(\dtop.vtop.pipeline.zg[1] ),
    .Y(_1999_));
 sg13g2_a221oi_1 _5921_ (.B2(_1998_),
    .C1(_1999_),
    .B1(_1997_),
    .A1(_3072_),
    .Y(_2000_),
    .A2(\dtop.vtop.pipeline.zg[2] ));
 sg13g2_nand2b_1 _5922_ (.Y(_2001_),
    .B(\dtop.vtop.pipeline.z[8] ),
    .A_N(\dtop.vtop.pipeline.zg[3] ));
 sg13g2_o21ai_1 _5923_ (.B1(_2001_),
    .Y(_2002_),
    .A1(_3072_),
    .A2(\dtop.vtop.pipeline.zg[2] ));
 sg13g2_a22oi_1 _5924_ (.Y(_2003_),
    .B1(\dtop.vtop.pipeline.zg[3] ),
    .B2(_3071_),
    .A2(\dtop.vtop.pipeline.zg[4] ),
    .A1(_3070_));
 sg13g2_o21ai_1 _5925_ (.B1(_2003_),
    .Y(_2004_),
    .A1(_2000_),
    .A2(_2002_));
 sg13g2_a22oi_1 _5926_ (.Y(_2005_),
    .B1(_1996_),
    .B2(_2004_),
    .A2(\dtop.vtop.pipeline.zg[5] ),
    .A1(_3069_));
 sg13g2_nand2_1 _5927_ (.Y(_2006_),
    .A(\dtop.vtop.pipeline.z[11] ),
    .B(_3123_));
 sg13g2_o21ai_1 _5928_ (.B1(_2006_),
    .Y(_2007_),
    .A1(_3069_),
    .A2(\dtop.vtop.pipeline.zg[5] ));
 sg13g2_a22oi_1 _5929_ (.Y(_2008_),
    .B1(\dtop.vtop.pipeline.zg[6] ),
    .B2(_3068_),
    .A2(\dtop.vtop.pipeline.zg[7] ),
    .A1(_3067_));
 sg13g2_o21ai_1 _5930_ (.B1(_2008_),
    .Y(_2009_),
    .A1(_2005_),
    .A2(_2007_));
 sg13g2_a22oi_1 _5931_ (.Y(_2010_),
    .B1(_3122_),
    .B2(\dtop.vtop.pipeline.z[12] ),
    .A2(_3121_),
    .A1(\dtop.vtop.pipeline.z[13] ));
 sg13g2_a22oi_1 _5932_ (.Y(_2011_),
    .B1(\dtop.vtop.pipeline.zg[8] ),
    .B2(_3066_),
    .A2(net1355),
    .A1(_3065_));
 sg13g2_inv_1 _5933_ (.Y(_2012_),
    .A(_2011_));
 sg13g2_a21oi_2 _5934_ (.B1(_2012_),
    .Y(_2013_),
    .A2(_2010_),
    .A1(_2009_));
 sg13g2_a21o_1 _5935_ (.A2(_2010_),
    .A1(_2009_),
    .B1(_2012_),
    .X(_2014_));
 sg13g2_nor2_1 _5936_ (.A(_1994_),
    .B(_2013_),
    .Y(_2015_));
 sg13g2_inv_2 _5937_ (.Y(_2016_),
    .A(net1231));
 sg13g2_nand3_1 _5938_ (.B(_3202_),
    .C(_2016_),
    .A(net645),
    .Y(_2017_));
 sg13g2_nand3_1 _5939_ (.B(_3127_),
    .C(_3198_),
    .A(\dtop.detune_counter[14] ),
    .Y(_2018_));
 sg13g2_o21ai_1 _5940_ (.B1(_2018_),
    .Y(_2019_),
    .A1(_0090_),
    .A2(_0437_));
 sg13g2_nor3_1 _5941_ (.A(_3127_),
    .B(net1398),
    .C(_3320_),
    .Y(_2020_));
 sg13g2_o21ai_1 _5942_ (.B1(net1394),
    .Y(_2021_),
    .A1(_2019_),
    .A2(_2020_));
 sg13g2_nand2b_1 _5943_ (.Y(_2022_),
    .B(net632),
    .A_N(_2021_));
 sg13g2_nand2_1 _5944_ (.Y(_2023_),
    .A(_1535_),
    .B(_2022_));
 sg13g2_nor2_1 _5945_ (.A(\dtop.vtop.pipeline.wave_index[0] ),
    .B(_2021_),
    .Y(_2024_));
 sg13g2_a21oi_1 _5946_ (.A1(_1535_),
    .A2(_2022_),
    .Y(_2025_),
    .B1(_2024_));
 sg13g2_inv_1 _5947_ (.Y(_2026_),
    .A(net1228));
 sg13g2_and2_1 _5948_ (.A(_2017_),
    .B(net1229),
    .X(_2027_));
 sg13g2_nand2_2 _5949_ (.Y(_2028_),
    .A(_2017_),
    .B(net1229));
 sg13g2_nor2_2 _5950_ (.A(net1293),
    .B(_2028_),
    .Y(_2029_));
 sg13g2_mux2_1 _5951_ (.A0(net1366),
    .A1(net689),
    .S(_2029_),
    .X(_0265_));
 sg13g2_mux2_1 _5952_ (.A0(net1364),
    .A1(net1354),
    .S(_2029_),
    .X(_0266_));
 sg13g2_nor2_1 _5953_ (.A(_0091_),
    .B(_2016_),
    .Y(_2030_));
 sg13g2_o21ai_1 _5954_ (.B1(net1230),
    .Y(_2031_),
    .A1(net1365),
    .A2(net1363));
 sg13g2_nor2_1 _5955_ (.A(_0076_),
    .B(net1230),
    .Y(_2032_));
 sg13g2_a21oi_1 _5956_ (.A1(_3124_),
    .A2(net1234),
    .Y(_2033_),
    .B1(_2032_));
 sg13g2_nand2_1 _5957_ (.Y(_2034_),
    .A(_2031_),
    .B(_2033_));
 sg13g2_xor2_1 _5958_ (.B(_2033_),
    .A(_2031_),
    .X(_2035_));
 sg13g2_o21ai_1 _5959_ (.B1(net1306),
    .Y(_2036_),
    .A1(net610),
    .A2(net1165));
 sg13g2_a21oi_1 _5960_ (.A1(net1165),
    .A2(_2035_),
    .Y(_0267_),
    .B1(_2036_));
 sg13g2_nand3_1 _5961_ (.B(_3125_),
    .C(net1230),
    .A(net1365),
    .Y(_2037_));
 sg13g2_mux2_1 _5962_ (.A0(_0065_),
    .A1(_0024_),
    .S(net1230),
    .X(_2038_));
 sg13g2_xnor2_1 _5963_ (.Y(_2039_),
    .A(_2037_),
    .B(_2038_));
 sg13g2_xnor2_1 _5964_ (.Y(_2040_),
    .A(_2034_),
    .B(_2039_));
 sg13g2_o21ai_1 _5965_ (.B1(net1312),
    .Y(_2041_),
    .A1(net567),
    .A2(net1163));
 sg13g2_a21oi_1 _5966_ (.A1(net1163),
    .A2(_2040_),
    .Y(_0268_),
    .B1(_2041_));
 sg13g2_nand2b_1 _5967_ (.Y(_2042_),
    .B(_2038_),
    .A_N(_2040_));
 sg13g2_nor3_2 _5968_ (.A(net1365),
    .B(_3125_),
    .C(_2016_),
    .Y(_2043_));
 sg13g2_mux2_1 _5969_ (.A0(_0099_),
    .A1(_0022_),
    .S(net1234),
    .X(_2044_));
 sg13g2_nor2_1 _5970_ (.A(_2043_),
    .B(_2044_),
    .Y(_2045_));
 sg13g2_xor2_1 _5971_ (.B(_2044_),
    .A(_2043_),
    .X(_2046_));
 sg13g2_xnor2_1 _5972_ (.Y(_2047_),
    .A(_2042_),
    .B(_2046_));
 sg13g2_o21ai_1 _5973_ (.B1(net1312),
    .Y(_2048_),
    .A1(net545),
    .A2(net1163));
 sg13g2_a21oi_1 _5974_ (.A1(net1163),
    .A2(_2047_),
    .Y(_0269_),
    .B1(_2048_));
 sg13g2_nor2_1 _5975_ (.A(_2045_),
    .B(_2047_),
    .Y(_2049_));
 sg13g2_mux2_1 _5976_ (.A0(_0098_),
    .A1(_0066_),
    .S(net1232),
    .X(_2050_));
 sg13g2_nand3_1 _5977_ (.B(net1363),
    .C(net1232),
    .A(\dtop.vtop.pipeline.nstep_zg[0] ),
    .Y(_2051_));
 sg13g2_xnor2_1 _5978_ (.Y(_2052_),
    .A(_2050_),
    .B(_2051_));
 sg13g2_xnor2_1 _5979_ (.Y(_2053_),
    .A(_2049_),
    .B(_2052_));
 sg13g2_inv_1 _5980_ (.Y(_2054_),
    .A(_2053_));
 sg13g2_o21ai_1 _5981_ (.B1(net1306),
    .Y(_2055_),
    .A1(net625),
    .A2(net1165));
 sg13g2_a21oi_1 _5982_ (.A1(net1165),
    .A2(_2054_),
    .Y(_0270_),
    .B1(_2055_));
 sg13g2_nand2_2 _5983_ (.Y(_2056_),
    .A(_2050_),
    .B(_2053_));
 sg13g2_mux2_1 _5984_ (.A0(\dtop.vtop.pipeline.dz[4] ),
    .A1(\dtop.vtop.pipeline.neg_t[4] ),
    .S(net1232),
    .X(_2057_));
 sg13g2_xor2_1 _5985_ (.B(_2057_),
    .A(_2056_),
    .X(_2058_));
 sg13g2_o21ai_1 _5986_ (.B1(net1312),
    .Y(_2059_),
    .A1(net566),
    .A2(net1163));
 sg13g2_a21oi_1 _5987_ (.A1(net1163),
    .A2(_2058_),
    .Y(_0271_),
    .B1(_2059_));
 sg13g2_mux2_1 _5988_ (.A0(\dtop.vtop.pipeline.dz[5] ),
    .A1(\dtop.vtop.pipeline.neg_t[5] ),
    .S(net1233),
    .X(_2060_));
 sg13g2_nor3_2 _5989_ (.A(_2056_),
    .B(_2057_),
    .C(_2060_),
    .Y(_2061_));
 sg13g2_o21ai_1 _5990_ (.B1(_2060_),
    .Y(_2062_),
    .A1(_2056_),
    .A2(_2057_));
 sg13g2_nand2b_1 _5991_ (.Y(_2063_),
    .B(_2062_),
    .A_N(_2061_));
 sg13g2_inv_1 _5992_ (.Y(_2064_),
    .A(_2063_));
 sg13g2_o21ai_1 _5993_ (.B1(net1312),
    .Y(_2065_),
    .A1(net601),
    .A2(net1164));
 sg13g2_a21oi_1 _5994_ (.A1(net1164),
    .A2(_2064_),
    .Y(_0272_),
    .B1(_2065_));
 sg13g2_mux2_1 _5995_ (.A0(_0096_),
    .A1(_0015_),
    .S(net1233),
    .X(_2066_));
 sg13g2_nand2_1 _5996_ (.Y(_2067_),
    .A(_2061_),
    .B(_2066_));
 sg13g2_xnor2_1 _5997_ (.Y(_2068_),
    .A(_2061_),
    .B(_2066_));
 sg13g2_inv_1 _5998_ (.Y(_2069_),
    .A(_2068_));
 sg13g2_o21ai_1 _5999_ (.B1(net1312),
    .Y(_2070_),
    .A1(net557),
    .A2(net1164));
 sg13g2_a21oi_1 _6000_ (.A1(net1164),
    .A2(_2069_),
    .Y(_0273_),
    .B1(_2070_));
 sg13g2_mux2_1 _6001_ (.A0(\dtop.vtop.pipeline.dz[7] ),
    .A1(\dtop.vtop.pipeline.neg_t[7] ),
    .S(net1233),
    .X(_2071_));
 sg13g2_nor2_1 _6002_ (.A(_2067_),
    .B(_2071_),
    .Y(_2072_));
 sg13g2_xor2_1 _6003_ (.B(_2071_),
    .A(_2067_),
    .X(_2073_));
 sg13g2_o21ai_1 _6004_ (.B1(net1312),
    .Y(_2074_),
    .A1(net627),
    .A2(net1163));
 sg13g2_a21oi_1 _6005_ (.A1(net1163),
    .A2(_2073_),
    .Y(_0274_),
    .B1(_2074_));
 sg13g2_mux2_1 _6006_ (.A0(_0094_),
    .A1(_0013_),
    .S(net1232),
    .X(_2075_));
 sg13g2_nand2_1 _6007_ (.Y(_2076_),
    .A(_2072_),
    .B(_2075_));
 sg13g2_xnor2_1 _6008_ (.Y(_2077_),
    .A(_2072_),
    .B(_2075_));
 sg13g2_inv_1 _6009_ (.Y(_2078_),
    .A(_2077_));
 sg13g2_o21ai_1 _6010_ (.B1(net1306),
    .Y(_2079_),
    .A1(net529),
    .A2(net1165));
 sg13g2_a21oi_1 _6011_ (.A1(net1165),
    .A2(_2078_),
    .Y(_0275_),
    .B1(_2079_));
 sg13g2_xnor2_1 _6012_ (.Y(_2080_),
    .A(_0026_),
    .B(_2076_));
 sg13g2_o21ai_1 _6013_ (.B1(net1312),
    .Y(_2081_),
    .A1(net577),
    .A2(net1164));
 sg13g2_a21oi_1 _6014_ (.A1(net1164),
    .A2(_2080_),
    .Y(_0276_),
    .B1(_2081_));
 sg13g2_or4_1 _6015_ (.A(_3064_),
    .B(_0091_),
    .C(_3278_),
    .D(net1230),
    .X(_2082_));
 sg13g2_a21oi_1 _6016_ (.A1(net599),
    .A2(net1101),
    .Y(_2083_),
    .B1(net1293));
 sg13g2_o21ai_1 _6017_ (.B1(_2083_),
    .Y(_0277_),
    .A1(_2035_),
    .A2(net1101));
 sg13g2_a21oi_1 _6018_ (.A1(net621),
    .A2(net1101),
    .Y(_2084_),
    .B1(net1293));
 sg13g2_o21ai_1 _6019_ (.B1(_2084_),
    .Y(_0278_),
    .A1(_2040_),
    .A2(net1101));
 sg13g2_a21oi_1 _6020_ (.A1(net559),
    .A2(net1101),
    .Y(_2085_),
    .B1(net1293));
 sg13g2_o21ai_1 _6021_ (.B1(_2085_),
    .Y(_0279_),
    .A1(_2047_),
    .A2(net1101));
 sg13g2_a21oi_1 _6022_ (.A1(net520),
    .A2(net1102),
    .Y(_2086_),
    .B1(net1294));
 sg13g2_o21ai_1 _6023_ (.B1(_2086_),
    .Y(_0280_),
    .A1(_2054_),
    .A2(net1103));
 sg13g2_a21oi_1 _6024_ (.A1(net617),
    .A2(net1102),
    .Y(_2087_),
    .B1(net1293));
 sg13g2_o21ai_1 _6025_ (.B1(_2087_),
    .Y(_0281_),
    .A1(_2058_),
    .A2(net1103));
 sg13g2_a21oi_1 _6026_ (.A1(net644),
    .A2(net1102),
    .Y(_2088_),
    .B1(net1299));
 sg13g2_o21ai_1 _6027_ (.B1(_2088_),
    .Y(_0282_),
    .A1(_2064_),
    .A2(net1102));
 sg13g2_a21oi_1 _6028_ (.A1(net576),
    .A2(net1102),
    .Y(_2089_),
    .B1(net1293));
 sg13g2_o21ai_1 _6029_ (.B1(_2089_),
    .Y(_0283_),
    .A1(_2069_),
    .A2(net1102));
 sg13g2_a21oi_1 _6030_ (.A1(net516),
    .A2(net1102),
    .Y(_2090_),
    .B1(net1293));
 sg13g2_o21ai_1 _6031_ (.B1(_2090_),
    .Y(_0284_),
    .A1(_2073_),
    .A2(net1102));
 sg13g2_a21oi_1 _6032_ (.A1(net595),
    .A2(net1101),
    .Y(_2091_),
    .B1(net1293));
 sg13g2_o21ai_1 _6033_ (.B1(_2091_),
    .Y(_0285_),
    .A1(_2078_),
    .A2(net1101));
 sg13g2_a21oi_1 _6034_ (.A1(_3278_),
    .A2(_2016_),
    .Y(_2092_),
    .B1(_3064_));
 sg13g2_nor2_1 _6035_ (.A(_3073_),
    .B(net1365),
    .Y(_2093_));
 sg13g2_nand2_1 _6036_ (.Y(_2094_),
    .A(_3125_),
    .B(_2093_));
 sg13g2_o21ai_1 _6037_ (.B1(_0075_),
    .Y(_2095_),
    .A1(_1994_),
    .A2(_2013_));
 sg13g2_nand3_1 _6038_ (.B(_2014_),
    .C(_2094_),
    .A(_1995_),
    .Y(_2096_));
 sg13g2_and2_1 _6039_ (.A(_2095_),
    .B(_2096_),
    .X(_2097_));
 sg13g2_a21oi_1 _6040_ (.A1(net1099),
    .A2(_2097_),
    .Y(_2098_),
    .B1(net487));
 sg13g2_nand3_1 _6041_ (.B(_2095_),
    .C(_2096_),
    .A(net487),
    .Y(_2099_));
 sg13g2_and3_1 _6042_ (.X(_2100_),
    .A(net487),
    .B(net1099),
    .C(_2097_));
 sg13g2_nor3_1 _6043_ (.A(net1294),
    .B(net488),
    .C(_2100_),
    .Y(_0286_));
 sg13g2_mux2_1 _6044_ (.A0(_0065_),
    .A1(_0076_),
    .S(net1365),
    .X(_2101_));
 sg13g2_a21oi_2 _6045_ (.B1(_0024_),
    .Y(_2102_),
    .A2(_2014_),
    .A1(_1995_));
 sg13g2_nor4_2 _6046_ (.A(net1363),
    .B(_1994_),
    .C(_2013_),
    .Y(_2103_),
    .D(_2101_));
 sg13g2_nor2_1 _6047_ (.A(_2102_),
    .B(_2103_),
    .Y(_2104_));
 sg13g2_o21ai_1 _6048_ (.B1(net712),
    .Y(_2105_),
    .A1(_2102_),
    .A2(_2103_));
 sg13g2_nor3_1 _6049_ (.A(\dtop.vtop.pipeline.z[1] ),
    .B(_2102_),
    .C(_2103_),
    .Y(_2106_));
 sg13g2_xor2_1 _6050_ (.B(_2104_),
    .A(net642),
    .X(_2107_));
 sg13g2_xnor2_1 _6051_ (.Y(_2108_),
    .A(_2099_),
    .B(_2107_));
 sg13g2_o21ai_1 _6052_ (.B1(net1305),
    .Y(_2109_),
    .A1(net642),
    .A2(net1098));
 sg13g2_a21oi_1 _6053_ (.A1(net1098),
    .A2(_2108_),
    .Y(_0287_),
    .B1(_2109_));
 sg13g2_mux2_1 _6054_ (.A0(_0099_),
    .A1(_0065_),
    .S(net1365),
    .X(_2110_));
 sg13g2_nor2_1 _6055_ (.A(net1363),
    .B(_2110_),
    .Y(_2111_));
 sg13g2_a21oi_1 _6056_ (.A1(net1363),
    .A2(_2093_),
    .Y(_2112_),
    .B1(_2111_));
 sg13g2_mux2_2 _6057_ (.A0(_0022_),
    .A1(_2112_),
    .S(net1231),
    .X(_2113_));
 sg13g2_nor2b_1 _6058_ (.A(_2113_),
    .B_N(\dtop.vtop.pipeline.z[2] ),
    .Y(_2114_));
 sg13g2_xnor2_1 _6059_ (.Y(_2115_),
    .A(net623),
    .B(_2113_));
 sg13g2_o21ai_1 _6060_ (.B1(_2105_),
    .Y(_2116_),
    .A1(_2099_),
    .A2(_2106_));
 sg13g2_xnor2_1 _6061_ (.Y(_2117_),
    .A(_2115_),
    .B(_2116_));
 sg13g2_o21ai_1 _6062_ (.B1(net1305),
    .Y(_2118_),
    .A1(net623),
    .A2(net1098));
 sg13g2_a21oi_1 _6063_ (.A1(net1098),
    .A2(_2117_),
    .Y(_0288_),
    .B1(_2118_));
 sg13g2_mux2_1 _6064_ (.A0(_0098_),
    .A1(_0099_),
    .S(net1365),
    .X(_2119_));
 sg13g2_mux2_1 _6065_ (.A0(_2101_),
    .A1(_2119_),
    .S(_3125_),
    .X(_2120_));
 sg13g2_mux2_1 _6066_ (.A0(_0066_),
    .A1(_2120_),
    .S(net1230),
    .X(_2121_));
 sg13g2_nand2b_1 _6067_ (.Y(_2122_),
    .B(net711),
    .A_N(_2121_));
 sg13g2_xor2_1 _6068_ (.B(_2121_),
    .A(net641),
    .X(_2123_));
 sg13g2_a21oi_1 _6069_ (.A1(_2115_),
    .A2(_2116_),
    .Y(_2124_),
    .B1(_2114_));
 sg13g2_xnor2_1 _6070_ (.Y(_2125_),
    .A(_2123_),
    .B(_2124_));
 sg13g2_o21ai_1 _6071_ (.B1(net1305),
    .Y(_2126_),
    .A1(net641),
    .A2(net1098));
 sg13g2_a21oi_1 _6072_ (.A1(net1098),
    .A2(_2125_),
    .Y(_0289_),
    .B1(_2126_));
 sg13g2_nor2_1 _6073_ (.A(_0019_),
    .B(net1233),
    .Y(_2127_));
 sg13g2_nand2b_1 _6074_ (.Y(_2128_),
    .B(net1364),
    .A_N(_2110_));
 sg13g2_mux2_1 _6075_ (.A0(_0072_),
    .A1(_0098_),
    .S(net1366),
    .X(_2129_));
 sg13g2_o21ai_1 _6076_ (.B1(_2128_),
    .Y(_2130_),
    .A1(net1364),
    .A2(_2129_));
 sg13g2_a21oi_2 _6077_ (.B1(_2127_),
    .Y(_2131_),
    .A2(_2130_),
    .A1(net1232));
 sg13g2_nor2b_1 _6078_ (.A(_2131_),
    .B_N(\dtop.vtop.pipeline.z[4] ),
    .Y(_2132_));
 sg13g2_xnor2_1 _6079_ (.Y(_2133_),
    .A(net608),
    .B(_2131_));
 sg13g2_o21ai_1 _6080_ (.B1(_2122_),
    .Y(_2134_),
    .A1(_2123_),
    .A2(_2124_));
 sg13g2_xnor2_1 _6081_ (.Y(_2135_),
    .A(_2133_),
    .B(_2134_));
 sg13g2_o21ai_1 _6082_ (.B1(net1304),
    .Y(_2136_),
    .A1(net608),
    .A2(net1098));
 sg13g2_a21oi_1 _6083_ (.A1(net1098),
    .A2(_2135_),
    .Y(_0290_),
    .B1(_2136_));
 sg13g2_a21oi_1 _6084_ (.A1(_2133_),
    .A2(_2134_),
    .Y(_2137_),
    .B1(_2132_));
 sg13g2_mux2_1 _6085_ (.A0(_0097_),
    .A1(_0072_),
    .S(\dtop.vtop.pipeline.nstep_zg[0] ),
    .X(_2138_));
 sg13g2_mux2_1 _6086_ (.A0(_2119_),
    .A1(_2138_),
    .S(_3125_),
    .X(_2139_));
 sg13g2_mux2_2 _6087_ (.A0(_0017_),
    .A1(_2139_),
    .S(net1230),
    .X(_2140_));
 sg13g2_nand2b_1 _6088_ (.Y(_2141_),
    .B(\dtop.vtop.pipeline.z[5] ),
    .A_N(_2140_));
 sg13g2_nor2b_1 _6089_ (.A(\dtop.vtop.pipeline.z[5] ),
    .B_N(_2140_),
    .Y(_2142_));
 sg13g2_xor2_1 _6090_ (.B(_2140_),
    .A(net664),
    .X(_2143_));
 sg13g2_xnor2_1 _6091_ (.Y(_2144_),
    .A(_2137_),
    .B(_2143_));
 sg13g2_o21ai_1 _6092_ (.B1(net1304),
    .Y(_2145_),
    .A1(net664),
    .A2(net1097));
 sg13g2_a21oi_1 _6093_ (.A1(net1097),
    .A2(_2144_),
    .Y(_0291_),
    .B1(_2145_));
 sg13g2_mux2_1 _6094_ (.A0(_0096_),
    .A1(_0097_),
    .S(net1365),
    .X(_2146_));
 sg13g2_mux2_1 _6095_ (.A0(_2129_),
    .A1(_2146_),
    .S(_3125_),
    .X(_2147_));
 sg13g2_mux2_2 _6096_ (.A0(_0015_),
    .A1(_2147_),
    .S(net1232),
    .X(_2148_));
 sg13g2_nor2b_1 _6097_ (.A(_2148_),
    .B_N(\dtop.vtop.pipeline.z[6] ),
    .Y(_2149_));
 sg13g2_xor2_1 _6098_ (.B(_2148_),
    .A(\dtop.vtop.pipeline.z[6] ),
    .X(_2150_));
 sg13g2_inv_1 _6099_ (.Y(_2151_),
    .A(_2150_));
 sg13g2_o21ai_1 _6100_ (.B1(_2141_),
    .Y(_2152_),
    .A1(_2137_),
    .A2(_2142_));
 sg13g2_xnor2_1 _6101_ (.Y(_2153_),
    .A(_2151_),
    .B(_2152_));
 sg13g2_o21ai_1 _6102_ (.B1(net1304),
    .Y(_2154_),
    .A1(net652),
    .A2(net1097));
 sg13g2_a21oi_1 _6103_ (.A1(net1097),
    .A2(_2153_),
    .Y(_0292_),
    .B1(_2154_));
 sg13g2_mux2_1 _6104_ (.A0(_0095_),
    .A1(_0096_),
    .S(net1366),
    .X(_2155_));
 sg13g2_mux2_1 _6105_ (.A0(_2138_),
    .A1(_2155_),
    .S(_3125_),
    .X(_2156_));
 sg13g2_mux2_2 _6106_ (.A0(_0073_),
    .A1(_2156_),
    .S(net1232),
    .X(_2157_));
 sg13g2_nor2_1 _6107_ (.A(_3072_),
    .B(_2157_),
    .Y(_2158_));
 sg13g2_xnor2_1 _6108_ (.Y(_2159_),
    .A(\dtop.vtop.pipeline.z[7] ),
    .B(_2157_));
 sg13g2_a21o_1 _6109_ (.A2(_2152_),
    .A1(_2151_),
    .B1(_2149_),
    .X(_2160_));
 sg13g2_xnor2_1 _6110_ (.Y(_2161_),
    .A(_2159_),
    .B(_2160_));
 sg13g2_o21ai_1 _6111_ (.B1(net1304),
    .Y(_2162_),
    .A1(net622),
    .A2(net1097));
 sg13g2_a21oi_1 _6112_ (.A1(net1097),
    .A2(_2161_),
    .Y(_0293_),
    .B1(_2162_));
 sg13g2_nand2b_1 _6113_ (.Y(_2163_),
    .B(net1366),
    .A_N(_0095_));
 sg13g2_o21ai_1 _6114_ (.B1(_2163_),
    .Y(_2164_),
    .A1(net1366),
    .A2(_0094_));
 sg13g2_nand2_1 _6115_ (.Y(_2165_),
    .A(net1364),
    .B(_2146_));
 sg13g2_o21ai_1 _6116_ (.B1(_2165_),
    .Y(_2166_),
    .A1(net1364),
    .A2(_2164_));
 sg13g2_mux2_1 _6117_ (.A0(_0013_),
    .A1(_2166_),
    .S(net1230),
    .X(_2167_));
 sg13g2_nor2_1 _6118_ (.A(_3071_),
    .B(_2167_),
    .Y(_2168_));
 sg13g2_xnor2_1 _6119_ (.Y(_2169_),
    .A(\dtop.vtop.pipeline.z[8] ),
    .B(_2167_));
 sg13g2_a21o_1 _6120_ (.A2(_2160_),
    .A1(_2159_),
    .B1(_2158_),
    .X(_2170_));
 sg13g2_xor2_1 _6121_ (.B(_2170_),
    .A(_2169_),
    .X(_2171_));
 sg13g2_nand2b_1 _6122_ (.Y(_2172_),
    .B(net1099),
    .A_N(_2171_));
 sg13g2_o21ai_1 _6123_ (.B1(_2172_),
    .Y(_2173_),
    .A1(net630),
    .A2(net1099));
 sg13g2_nor2_1 _6124_ (.A(net1294),
    .B(_2173_),
    .Y(_0294_));
 sg13g2_nor2_1 _6125_ (.A(_0026_),
    .B(net1233),
    .Y(_2174_));
 sg13g2_a21oi_1 _6126_ (.A1(\dtop.vtop.pipeline.dz[8] ),
    .A2(net1366),
    .Y(_2175_),
    .B1(net1364));
 sg13g2_a21oi_1 _6127_ (.A1(net1364),
    .A2(_2155_),
    .Y(_2176_),
    .B1(_2175_));
 sg13g2_a21oi_2 _6128_ (.B1(_2174_),
    .Y(_2177_),
    .A2(_2176_),
    .A1(net1232));
 sg13g2_nand2_1 _6129_ (.Y(_2178_),
    .A(_3070_),
    .B(_2177_));
 sg13g2_nor2_1 _6130_ (.A(_3070_),
    .B(_2177_),
    .Y(_2179_));
 sg13g2_xnor2_1 _6131_ (.Y(_2180_),
    .A(net637),
    .B(_2177_));
 sg13g2_a21o_1 _6132_ (.A2(_2170_),
    .A1(_2169_),
    .B1(_2168_),
    .X(_2181_));
 sg13g2_xnor2_1 _6133_ (.Y(_2182_),
    .A(_2180_),
    .B(_2181_));
 sg13g2_o21ai_1 _6134_ (.B1(net1304),
    .Y(_2183_),
    .A1(net637),
    .A2(net1097));
 sg13g2_a21oi_1 _6135_ (.A1(net1097),
    .A2(_2182_),
    .Y(_0295_),
    .B1(_2183_));
 sg13g2_a21oi_1 _6136_ (.A1(net1363),
    .A2(_2164_),
    .Y(_2184_),
    .B1(_2016_));
 sg13g2_nand2b_1 _6137_ (.Y(_2185_),
    .B(\dtop.vtop.pipeline.z[10] ),
    .A_N(_2184_));
 sg13g2_xnor2_1 _6138_ (.Y(_2186_),
    .A(\dtop.vtop.pipeline.z[10] ),
    .B(_2184_));
 sg13g2_and2_1 _6139_ (.A(_2178_),
    .B(_2181_),
    .X(_2187_));
 sg13g2_nor3_1 _6140_ (.A(_2179_),
    .B(_2186_),
    .C(_2187_),
    .Y(_2188_));
 sg13g2_o21ai_1 _6141_ (.B1(_2186_),
    .Y(_2189_),
    .A1(_2179_),
    .A2(_2187_));
 sg13g2_nor2b_1 _6142_ (.A(_2188_),
    .B_N(_2189_),
    .Y(_2190_));
 sg13g2_nand2b_1 _6143_ (.Y(_2191_),
    .B(net1099),
    .A_N(_2190_));
 sg13g2_o21ai_1 _6144_ (.B1(_2191_),
    .Y(_2192_),
    .A1(net640),
    .A2(net1099));
 sg13g2_nor2_1 _6145_ (.A(net1294),
    .B(_2192_),
    .Y(_0296_));
 sg13g2_nand3_1 _6146_ (.B(net1366),
    .C(net1363),
    .A(\dtop.vtop.pipeline.dz[8] ),
    .Y(_2193_));
 sg13g2_nand3_1 _6147_ (.B(net1231),
    .C(_2193_),
    .A(_3068_),
    .Y(_2194_));
 sg13g2_a21o_1 _6148_ (.A2(_2193_),
    .A1(net1231),
    .B1(_3068_),
    .X(_2195_));
 sg13g2_nand2_1 _6149_ (.Y(_2196_),
    .A(_2194_),
    .B(_2195_));
 sg13g2_and2_1 _6150_ (.A(_2185_),
    .B(_2189_),
    .X(_2197_));
 sg13g2_xnor2_1 _6151_ (.Y(_2198_),
    .A(_2196_),
    .B(_2197_));
 sg13g2_o21ai_1 _6152_ (.B1(net1304),
    .Y(_2199_),
    .A1(net579),
    .A2(net1099));
 sg13g2_a21oi_1 _6153_ (.A1(net1099),
    .A2(_2198_),
    .Y(_0297_),
    .B1(_2199_));
 sg13g2_xnor2_1 _6154_ (.Y(_2200_),
    .A(_3067_),
    .B(net1231));
 sg13g2_nand2_1 _6155_ (.Y(_2201_),
    .A(_2195_),
    .B(_2197_));
 sg13g2_nand2_1 _6156_ (.Y(_2202_),
    .A(_2194_),
    .B(_2201_));
 sg13g2_xnor2_1 _6157_ (.Y(_2203_),
    .A(_2200_),
    .B(_2202_));
 sg13g2_o21ai_1 _6158_ (.B1(net1305),
    .Y(_2204_),
    .A1(net619),
    .A2(net1100));
 sg13g2_a21oi_1 _6159_ (.A1(net1100),
    .A2(_2203_),
    .Y(_0298_),
    .B1(_2204_));
 sg13g2_nor3_1 _6160_ (.A(_3067_),
    .B(_2016_),
    .C(_2202_),
    .Y(_2205_));
 sg13g2_nor3_1 _6161_ (.A(\dtop.vtop.pipeline.z[12] ),
    .B(net1231),
    .C(_2201_),
    .Y(_2206_));
 sg13g2_o21ai_1 _6162_ (.B1(net1100),
    .Y(_2207_),
    .A1(_2205_),
    .A2(_2206_));
 sg13g2_o21ai_1 _6163_ (.B1(net1304),
    .Y(_2208_),
    .A1(_3066_),
    .A2(_2207_));
 sg13g2_nand2_1 _6164_ (.Y(_2209_),
    .A(_3066_),
    .B(net1231));
 sg13g2_a21oi_1 _6165_ (.A1(_3066_),
    .A2(_2207_),
    .Y(_0299_),
    .B1(_2208_));
 sg13g2_o21ai_1 _6166_ (.B1(_2209_),
    .Y(_2210_),
    .A1(_3066_),
    .A2(_2205_));
 sg13g2_nor2_1 _6167_ (.A(_2207_),
    .B(_2210_),
    .Y(_2211_));
 sg13g2_o21ai_1 _6168_ (.B1(net1304),
    .Y(_2212_),
    .A1(net426),
    .A2(_2211_));
 sg13g2_a21oi_1 _6169_ (.A1(net426),
    .A2(_2211_),
    .Y(_0300_),
    .B1(_2212_));
 sg13g2_nand3_1 _6170_ (.B(_3148_),
    .C(net1307),
    .A(\dtop.vtop.pipeline.wave_index[0] ),
    .Y(_2213_));
 sg13g2_o21ai_1 _6171_ (.B1(_2213_),
    .Y(_2214_),
    .A1(net1382),
    .A2(_1538_));
 sg13g2_nand2_1 _6172_ (.Y(_2215_),
    .A(_0029_),
    .B(net1275));
 sg13g2_nand2_1 _6173_ (.Y(_2216_),
    .A(\dtop.vtop.pipeline.phases[1][0] ),
    .B(net1291));
 sg13g2_a22oi_1 _6174_ (.Y(_2217_),
    .B1(net1286),
    .B2(_2216_),
    .A2(_1544_),
    .A1(_3161_));
 sg13g2_xnor2_1 _6175_ (.Y(_2218_),
    .A(net1289),
    .B(net1287));
 sg13g2_nor3_1 _6176_ (.A(\dtop.vtop.dphases[2][0] ),
    .B(net1289),
    .C(net1285),
    .Y(_2219_));
 sg13g2_a221oi_1 _6177_ (.B2(_0031_),
    .C1(_2219_),
    .B1(net1263),
    .A1(_3162_),
    .Y(_2220_),
    .A2(net1271));
 sg13g2_and2_1 _6178_ (.A(net1351),
    .B(_2220_),
    .X(_2221_));
 sg13g2_a22oi_1 _6179_ (.Y(_2222_),
    .B1(_2221_),
    .B2(_0030_),
    .A2(_2217_),
    .A1(_2215_));
 sg13g2_nand4_1 _6180_ (.B(_2215_),
    .C(_2217_),
    .A(_0030_),
    .Y(_2223_),
    .D(_2221_));
 sg13g2_nand2_1 _6181_ (.Y(_2224_),
    .A(net1310),
    .B(_2223_));
 sg13g2_nor2_1 _6182_ (.A(_2222_),
    .B(_2224_),
    .Y(_2225_));
 sg13g2_mux2_1 _6183_ (.A0(net448),
    .A1(_2225_),
    .S(net1251),
    .X(_0301_));
 sg13g2_a21oi_1 _6184_ (.A1(\dtop.vtop.pipeline.phases[2][1] ),
    .A2(_1546_),
    .Y(_2226_),
    .B1(net1291));
 sg13g2_a221oi_1 _6185_ (.B2(_0032_),
    .C1(_2226_),
    .B1(net1275),
    .A1(_3163_),
    .Y(_2227_),
    .A2(net1286));
 sg13g2_nor3_1 _6186_ (.A(\dtop.vtop.dphases[2][1] ),
    .B(net1289),
    .C(net1285),
    .Y(_2228_));
 sg13g2_a221oi_1 _6187_ (.B2(_0033_),
    .C1(_2228_),
    .B1(_2218_),
    .A1(_3164_),
    .Y(_2229_),
    .A2(net1271));
 sg13g2_mux2_2 _6188_ (.A0(_2220_),
    .A1(_2229_),
    .S(net1351),
    .X(_2230_));
 sg13g2_nand3_1 _6189_ (.B(_2227_),
    .C(_2230_),
    .A(_0030_),
    .Y(_2231_));
 sg13g2_a21oi_1 _6190_ (.A1(_0030_),
    .A2(_2230_),
    .Y(_2232_),
    .B1(_2227_));
 sg13g2_a21o_1 _6191_ (.A2(_2230_),
    .A1(_0030_),
    .B1(_2227_),
    .X(_2233_));
 sg13g2_nand2_1 _6192_ (.Y(_2234_),
    .A(_2231_),
    .B(_2233_));
 sg13g2_xnor2_1 _6193_ (.Y(_2235_),
    .A(_2223_),
    .B(_2234_));
 sg13g2_nor2_2 _6194_ (.A(_0093_),
    .B(net1313),
    .Y(_2236_));
 sg13g2_xor2_1 _6195_ (.B(\dtop.player_inst.program_addr[2] ),
    .A(net1398),
    .X(_2237_));
 sg13g2_xor2_1 _6196_ (.B(\dtop.player_inst.program_addr[1] ),
    .A(net1400),
    .X(_2238_));
 sg13g2_or2_1 _6197_ (.X(_2239_),
    .B(_2238_),
    .A(_2237_));
 sg13g2_nor2_1 _6198_ (.A(_0729_),
    .B(_2239_),
    .Y(_2240_));
 sg13g2_nor2b_1 _6199_ (.A(_2240_),
    .B_N(_2236_),
    .Y(_2241_));
 sg13g2_nand2b_2 _6200_ (.Y(_2242_),
    .B(_2236_),
    .A_N(_2240_));
 sg13g2_nor2_1 _6201_ (.A(net1309),
    .B(net1261),
    .Y(_2243_));
 sg13g2_nand2_1 _6202_ (.Y(_2244_),
    .A(net1379),
    .B(_0728_));
 sg13g2_nand4_1 _6203_ (.B(_3321_),
    .C(_0728_),
    .A(net1379),
    .Y(_2245_),
    .D(_1879_));
 sg13g2_a21o_1 _6204_ (.A2(_2245_),
    .A1(_2238_),
    .B1(_2244_),
    .X(_2246_));
 sg13g2_a21oi_1 _6205_ (.A1(_3152_),
    .A2(_2244_),
    .Y(_2247_),
    .B1(net1309));
 sg13g2_and2_1 _6206_ (.A(_2246_),
    .B(_2247_),
    .X(_2248_));
 sg13g2_nor3_2 _6207_ (.A(net1311),
    .B(net1261),
    .C(_2248_),
    .Y(_2249_));
 sg13g2_nand3_1 _6208_ (.B(_2238_),
    .C(_2245_),
    .A(_2237_),
    .Y(_2250_));
 sg13g2_nand4_1 _6209_ (.B(_0728_),
    .C(_2239_),
    .A(net1379),
    .Y(_2251_),
    .D(_2250_));
 sg13g2_a21oi_1 _6210_ (.A1(_3138_),
    .A2(_2244_),
    .Y(_2252_),
    .B1(net1309));
 sg13g2_nand2_1 _6211_ (.Y(_2253_),
    .A(_2251_),
    .B(_2252_));
 sg13g2_nand2_1 _6212_ (.Y(_2254_),
    .A(_2249_),
    .B(_2253_));
 sg13g2_o21ai_1 _6213_ (.B1(_2254_),
    .Y(_2255_),
    .A1(net1298),
    .A2(_2235_));
 sg13g2_nand2_1 _6214_ (.Y(_2256_),
    .A(net1250),
    .B(_2255_));
 sg13g2_o21ai_1 _6215_ (.B1(_2256_),
    .Y(_0302_),
    .A1(_3163_),
    .A2(net1250));
 sg13g2_o21ai_1 _6216_ (.B1(_2231_),
    .Y(_2257_),
    .A1(_2223_),
    .A2(_2232_));
 sg13g2_a21oi_1 _6217_ (.A1(\dtop.vtop.pipeline.phases[2][2] ),
    .A2(net1288),
    .Y(_2258_),
    .B1(net1291));
 sg13g2_a221oi_1 _6218_ (.B2(_0034_),
    .C1(_2258_),
    .B1(net1275),
    .A1(_3165_),
    .Y(_2259_),
    .A2(net1286));
 sg13g2_nor3_1 _6219_ (.A(\dtop.vtop.dphases[2][2] ),
    .B(net1289),
    .C(net1285),
    .Y(_2260_));
 sg13g2_a221oi_1 _6220_ (.B2(_0035_),
    .C1(_2260_),
    .B1(_2218_),
    .A1(_3166_),
    .Y(_2261_),
    .A2(net1271));
 sg13g2_mux2_1 _6221_ (.A0(_2229_),
    .A1(_2261_),
    .S(net1351),
    .X(_2262_));
 sg13g2_mux2_1 _6222_ (.A0(_2262_),
    .A1(_2221_),
    .S(net1353),
    .X(_2263_));
 sg13g2_and2_1 _6223_ (.A(_2259_),
    .B(_2263_),
    .X(_2264_));
 sg13g2_or2_1 _6224_ (.X(_2265_),
    .B(_2263_),
    .A(_2259_));
 sg13g2_nand2b_1 _6225_ (.Y(_2266_),
    .B(_2265_),
    .A_N(_2264_));
 sg13g2_xor2_1 _6226_ (.B(_2266_),
    .A(_2257_),
    .X(_2267_));
 sg13g2_o21ai_1 _6227_ (.B1(_2254_),
    .Y(_2268_),
    .A1(net1298),
    .A2(_2267_));
 sg13g2_nand2_1 _6228_ (.Y(_2269_),
    .A(net1250),
    .B(_2268_));
 sg13g2_o21ai_1 _6229_ (.B1(_2269_),
    .Y(_0303_),
    .A1(_3165_),
    .A2(net1250));
 sg13g2_a21oi_1 _6230_ (.A1(_2257_),
    .A2(_2265_),
    .Y(_2270_),
    .B1(_2264_));
 sg13g2_a21oi_1 _6231_ (.A1(\dtop.vtop.pipeline.phases[1][3] ),
    .A2(net1291),
    .Y(_2271_),
    .B1(net1288));
 sg13g2_a221oi_1 _6232_ (.B2(_0036_),
    .C1(_2271_),
    .B1(net1275),
    .A1(_3167_),
    .Y(_2272_),
    .A2(_1544_));
 sg13g2_nor3_1 _6233_ (.A(\dtop.vtop.dphases[2][3] ),
    .B(net1289),
    .C(net1285),
    .Y(_2273_));
 sg13g2_a221oi_1 _6234_ (.B2(_0037_),
    .C1(_2273_),
    .B1(_2218_),
    .A1(_3168_),
    .Y(_2274_),
    .A2(net1271));
 sg13g2_mux2_1 _6235_ (.A0(_2261_),
    .A1(_2274_),
    .S(net1351),
    .X(_2275_));
 sg13g2_mux2_1 _6236_ (.A0(_2275_),
    .A1(_2230_),
    .S(net1353),
    .X(_2276_));
 sg13g2_and2_1 _6237_ (.A(_2272_),
    .B(_2276_),
    .X(_2277_));
 sg13g2_inv_1 _6238_ (.Y(_2278_),
    .A(_2277_));
 sg13g2_xnor2_1 _6239_ (.Y(_2279_),
    .A(_2272_),
    .B(_2276_));
 sg13g2_xor2_1 _6240_ (.B(_2279_),
    .A(_2270_),
    .X(_2280_));
 sg13g2_a21o_1 _6241_ (.A2(_2280_),
    .A1(net1310),
    .B1(_2249_),
    .X(_2281_));
 sg13g2_mux2_1 _6242_ (.A0(net478),
    .A1(_2281_),
    .S(net1251),
    .X(_0304_));
 sg13g2_nor2_1 _6243_ (.A(net467),
    .B(net1251),
    .Y(_2282_));
 sg13g2_nor2_1 _6244_ (.A(_3250_),
    .B(net1299),
    .Y(_2283_));
 sg13g2_a22oi_1 _6245_ (.Y(_2284_),
    .B1(_2246_),
    .B2(_2247_),
    .A2(net1309),
    .A1(_3249_));
 sg13g2_or2_1 _6246_ (.X(_2285_),
    .B(_2283_),
    .A(_2248_));
 sg13g2_nor2_1 _6247_ (.A(\dtop.detune_counter[4] ),
    .B(net1259),
    .Y(_2286_));
 sg13g2_a21o_1 _6248_ (.A2(_2252_),
    .A1(_2251_),
    .B1(_2283_),
    .X(_2287_));
 sg13g2_a21oi_1 _6249_ (.A1(net1248),
    .A2(net1246),
    .Y(_2288_),
    .B1(_2286_));
 sg13g2_o21ai_1 _6250_ (.B1(_2278_),
    .Y(_2289_),
    .A1(_2270_),
    .A2(_2279_));
 sg13g2_nor3_1 _6251_ (.A(_0038_),
    .B(_1544_),
    .C(net1286),
    .Y(_2290_));
 sg13g2_a221oi_1 _6252_ (.B2(\dtop.vtop.pipeline.phases[1][4] ),
    .C1(_2290_),
    .B1(net1271),
    .A1(\dtop.vtop.pipeline.phases[2][4] ),
    .Y(_2291_),
    .A2(_1550_));
 sg13g2_a22oi_1 _6253_ (.Y(_2292_),
    .B1(net1263),
    .B2(_0039_),
    .A2(net1270),
    .A1(_3169_));
 sg13g2_o21ai_1 _6254_ (.B1(_2292_),
    .Y(_2293_),
    .A1(\dtop.vtop.dphases[2][4] ),
    .A2(_1551_));
 sg13g2_nor2_1 _6255_ (.A(net1351),
    .B(_2274_),
    .Y(_2294_));
 sg13g2_a21o_1 _6256_ (.A2(_2293_),
    .A1(net1350),
    .B1(_2294_),
    .X(_2295_));
 sg13g2_nor2_1 _6257_ (.A(net1353),
    .B(_2295_),
    .Y(_2296_));
 sg13g2_a21oi_2 _6258_ (.B1(_2296_),
    .Y(_2297_),
    .A2(_2262_),
    .A1(net1353));
 sg13g2_nor2_1 _6259_ (.A(_2291_),
    .B(_2297_),
    .Y(_2298_));
 sg13g2_xor2_1 _6260_ (.B(_2297_),
    .A(_2291_),
    .X(_2299_));
 sg13g2_xor2_1 _6261_ (.B(_2299_),
    .A(_2289_),
    .X(_2300_));
 sg13g2_a22oi_1 _6262_ (.Y(_2301_),
    .B1(_2300_),
    .B2(net1309),
    .A2(_2288_),
    .A1(_2243_));
 sg13g2_a21oi_1 _6263_ (.A1(net1251),
    .A2(_2301_),
    .Y(_0305_),
    .B1(_2282_));
 sg13g2_nand2b_1 _6264_ (.Y(_2302_),
    .B(_3198_),
    .A_N(_3212_));
 sg13g2_nand2_1 _6265_ (.Y(_2303_),
    .A(_3126_),
    .B(net1397));
 sg13g2_nor3_1 _6266_ (.A(_3199_),
    .B(_1533_),
    .C(_2303_),
    .Y(_2304_));
 sg13g2_a21oi_2 _6267_ (.B1(_2304_),
    .Y(_2305_),
    .A2(_2302_),
    .A1(_2236_));
 sg13g2_a21o_1 _6268_ (.A2(_2302_),
    .A1(_2236_),
    .B1(_2304_),
    .X(_2306_));
 sg13g2_nor2_1 _6269_ (.A(_0082_),
    .B(net1240),
    .Y(_2307_));
 sg13g2_a21oi_1 _6270_ (.A1(_2253_),
    .A2(net1259),
    .Y(_2308_),
    .B1(_2242_));
 sg13g2_mux2_1 _6271_ (.A0(_0077_),
    .A1(\dtop.detune_counter[4] ),
    .S(net1259),
    .X(_2309_));
 sg13g2_mux2_1 _6272_ (.A0(_2309_),
    .A1(net1248),
    .S(net1247),
    .X(_2310_));
 sg13g2_a21oi_1 _6273_ (.A1(_2242_),
    .A2(_2310_),
    .Y(_2311_),
    .B1(_2308_));
 sg13g2_nand2_1 _6274_ (.Y(_2312_),
    .A(_2307_),
    .B(_2311_));
 sg13g2_xor2_1 _6275_ (.B(_2311_),
    .A(_2307_),
    .X(_2313_));
 sg13g2_a21oi_1 _6276_ (.A1(_2289_),
    .A2(_2299_),
    .Y(_2314_),
    .B1(_2298_));
 sg13g2_nor3_1 _6277_ (.A(_0040_),
    .B(_1544_),
    .C(net1285),
    .Y(_2315_));
 sg13g2_a221oi_1 _6278_ (.B2(\dtop.vtop.pipeline.phases[1][5] ),
    .C1(_2315_),
    .B1(net1271),
    .A1(\dtop.vtop.pipeline.phases[2][5] ),
    .Y(_2316_),
    .A2(_1550_));
 sg13g2_a22oi_1 _6279_ (.Y(_2317_),
    .B1(net1263),
    .B2(_0041_),
    .A2(net1270),
    .A1(_3170_));
 sg13g2_o21ai_1 _6280_ (.B1(_2317_),
    .Y(_2318_),
    .A1(\dtop.vtop.dphases[2][5] ),
    .A2(_1551_));
 sg13g2_mux2_1 _6281_ (.A0(_2293_),
    .A1(_2318_),
    .S(net1350),
    .X(_2319_));
 sg13g2_nor2_1 _6282_ (.A(net1354),
    .B(_2319_),
    .Y(_2320_));
 sg13g2_a21oi_2 _6283_ (.B1(_2320_),
    .Y(_2321_),
    .A2(_2275_),
    .A1(net1353));
 sg13g2_nor2_1 _6284_ (.A(_2316_),
    .B(_2321_),
    .Y(_2322_));
 sg13g2_inv_1 _6285_ (.Y(_2323_),
    .A(_2322_));
 sg13g2_xnor2_1 _6286_ (.Y(_2324_),
    .A(_2316_),
    .B(_2321_));
 sg13g2_o21ai_1 _6287_ (.B1(net1310),
    .Y(_2325_),
    .A1(_2314_),
    .A2(_2324_));
 sg13g2_a21oi_1 _6288_ (.A1(_2314_),
    .A2(_2324_),
    .Y(_2326_),
    .B1(_2325_));
 sg13g2_a21o_1 _6289_ (.A2(_2313_),
    .A1(net1298),
    .B1(_2326_),
    .X(_2327_));
 sg13g2_mux2_1 _6290_ (.A0(net511),
    .A1(_2327_),
    .S(net1251),
    .X(_0306_));
 sg13g2_nor2_1 _6291_ (.A(_0081_),
    .B(net1240),
    .Y(_2328_));
 sg13g2_mux2_1 _6292_ (.A0(_0023_),
    .A1(\dtop.detune_counter[5] ),
    .S(net1259),
    .X(_2329_));
 sg13g2_mux2_1 _6293_ (.A0(_2329_),
    .A1(_2286_),
    .S(net1247),
    .X(_2330_));
 sg13g2_a21oi_1 _6294_ (.A1(_2242_),
    .A2(_2330_),
    .Y(_2331_),
    .B1(_2308_));
 sg13g2_and2_1 _6295_ (.A(_2328_),
    .B(_2331_),
    .X(_2332_));
 sg13g2_xnor2_1 _6296_ (.Y(_2333_),
    .A(_2328_),
    .B(_2331_));
 sg13g2_nor2_1 _6297_ (.A(_2312_),
    .B(_2333_),
    .Y(_2334_));
 sg13g2_a21oi_1 _6298_ (.A1(_2312_),
    .A2(_2333_),
    .Y(_2335_),
    .B1(net1309));
 sg13g2_nand2b_1 _6299_ (.Y(_2336_),
    .B(_2335_),
    .A_N(_2334_));
 sg13g2_o21ai_1 _6300_ (.B1(_2323_),
    .Y(_2337_),
    .A1(_2314_),
    .A2(_2324_));
 sg13g2_a22oi_1 _6301_ (.Y(_2338_),
    .B1(net1263),
    .B2(_0043_),
    .A2(net1270),
    .A1(_3171_));
 sg13g2_o21ai_1 _6302_ (.B1(_2338_),
    .Y(_2339_),
    .A1(\dtop.vtop.dphases[2][6] ),
    .A2(_1551_));
 sg13g2_mux2_1 _6303_ (.A0(_2318_),
    .A1(_2339_),
    .S(net1350),
    .X(_2340_));
 sg13g2_mux2_1 _6304_ (.A0(_2340_),
    .A1(_2295_),
    .S(net1353),
    .X(_2341_));
 sg13g2_nor2b_1 _6305_ (.A(_2341_),
    .B_N(_1589_),
    .Y(_2342_));
 sg13g2_xnor2_1 _6306_ (.Y(_2343_),
    .A(_1589_),
    .B(_2341_));
 sg13g2_xnor2_1 _6307_ (.Y(_2344_),
    .A(_2337_),
    .B(_2343_));
 sg13g2_o21ai_1 _6308_ (.B1(_2336_),
    .Y(_2345_),
    .A1(net1298),
    .A2(_2344_));
 sg13g2_mux2_1 _6309_ (.A0(net506),
    .A1(_2345_),
    .S(net1250),
    .X(_0307_));
 sg13g2_nor2_1 _6310_ (.A(_0046_),
    .B(net1240),
    .Y(_2346_));
 sg13g2_mux2_1 _6311_ (.A0(_0021_),
    .A1(\dtop.detune_counter[6] ),
    .S(net1259),
    .X(_2347_));
 sg13g2_mux2_1 _6312_ (.A0(_2347_),
    .A1(_2309_),
    .S(net1247),
    .X(_2348_));
 sg13g2_nor2_1 _6313_ (.A(net1262),
    .B(_2348_),
    .Y(_2349_));
 sg13g2_a21oi_1 _6314_ (.A1(net1261),
    .A2(net1259),
    .Y(_2350_),
    .B1(_2349_));
 sg13g2_nand2b_1 _6315_ (.Y(_2351_),
    .B(_2346_),
    .A_N(_2350_));
 sg13g2_xnor2_1 _6316_ (.Y(_2352_),
    .A(_2346_),
    .B(_2350_));
 sg13g2_or3_1 _6317_ (.A(_2332_),
    .B(_2334_),
    .C(_2352_),
    .X(_2353_));
 sg13g2_o21ai_1 _6318_ (.B1(_2352_),
    .Y(_2354_),
    .A1(_2332_),
    .A2(_2334_));
 sg13g2_nand3_1 _6319_ (.B(_2353_),
    .C(_2354_),
    .A(net1298),
    .Y(_2355_));
 sg13g2_a21oi_1 _6320_ (.A1(_2337_),
    .A2(_2343_),
    .Y(_2356_),
    .B1(_2342_));
 sg13g2_a22oi_1 _6321_ (.Y(_2357_),
    .B1(net1263),
    .B2(_0045_),
    .A2(net1270),
    .A1(_3172_));
 sg13g2_o21ai_1 _6322_ (.B1(_2357_),
    .Y(_2358_),
    .A1(\dtop.vtop.dphases[2][7] ),
    .A2(_1551_));
 sg13g2_mux2_1 _6323_ (.A0(_2339_),
    .A1(_2358_),
    .S(net1350),
    .X(_2359_));
 sg13g2_nand2b_1 _6324_ (.Y(_2360_),
    .B(net1353),
    .A_N(_2319_));
 sg13g2_o21ai_1 _6325_ (.B1(_2360_),
    .Y(_2361_),
    .A1(net1353),
    .A2(_2359_));
 sg13g2_nand2_1 _6326_ (.Y(_2362_),
    .A(_1584_),
    .B(_2361_));
 sg13g2_xnor2_1 _6327_ (.Y(_2363_),
    .A(_1584_),
    .B(_2361_));
 sg13g2_nor2_1 _6328_ (.A(_2356_),
    .B(_2363_),
    .Y(_2364_));
 sg13g2_a21o_1 _6329_ (.A2(_2363_),
    .A1(_2356_),
    .B1(net1298),
    .X(_2365_));
 sg13g2_o21ai_1 _6330_ (.B1(_2355_),
    .Y(_2366_),
    .A1(_2364_),
    .A2(_2365_));
 sg13g2_mux2_1 _6331_ (.A0(net479),
    .A1(_2366_),
    .S(net1250),
    .X(_0308_));
 sg13g2_nand2_2 _6332_ (.Y(_2367_),
    .A(net1425),
    .B(_2305_));
 sg13g2_nor2_1 _6333_ (.A(_0020_),
    .B(net1260),
    .Y(_2368_));
 sg13g2_a21oi_1 _6334_ (.A1(_3130_),
    .A2(net1260),
    .Y(_2369_),
    .B1(_2368_));
 sg13g2_mux2_1 _6335_ (.A0(_2369_),
    .A1(_2329_),
    .S(net1246),
    .X(_2370_));
 sg13g2_nand2_1 _6336_ (.Y(_2371_),
    .A(net1261),
    .B(_2288_));
 sg13g2_o21ai_1 _6337_ (.B1(_2371_),
    .Y(_2372_),
    .A1(net1261),
    .A2(_2370_));
 sg13g2_nor2b_1 _6338_ (.A(_2367_),
    .B_N(_2372_),
    .Y(_2373_));
 sg13g2_xor2_1 _6339_ (.B(_2372_),
    .A(_2367_),
    .X(_2374_));
 sg13g2_nand3_1 _6340_ (.B(_2354_),
    .C(_2374_),
    .A(_2351_),
    .Y(_2375_));
 sg13g2_a21oi_1 _6341_ (.A1(_2351_),
    .A2(_2354_),
    .Y(_2376_),
    .B1(_2374_));
 sg13g2_nand2_1 _6342_ (.Y(_2377_),
    .A(net1298),
    .B(_2375_));
 sg13g2_o21ai_1 _6343_ (.B1(_2362_),
    .Y(_2378_),
    .A1(_2356_),
    .A2(_2363_));
 sg13g2_nand2b_1 _6344_ (.Y(_2379_),
    .B(net1270),
    .A_N(\dtop.vtop.dphases[1][8] ));
 sg13g2_o21ai_1 _6345_ (.B1(_2379_),
    .Y(_2380_),
    .A1(\dtop.vtop.dphases[2][8] ),
    .A2(_1551_));
 sg13g2_a21oi_2 _6346_ (.B1(_2380_),
    .Y(_2381_),
    .A2(net1263),
    .A1(_0048_));
 sg13g2_nor2_1 _6347_ (.A(net1350),
    .B(_2358_),
    .Y(_2382_));
 sg13g2_a21oi_1 _6348_ (.A1(net1350),
    .A2(_2381_),
    .Y(_2383_),
    .B1(_2382_));
 sg13g2_mux2_1 _6349_ (.A0(_2383_),
    .A1(_2340_),
    .S(net1352),
    .X(_2384_));
 sg13g2_nor2b_1 _6350_ (.A(_2384_),
    .B_N(_1579_),
    .Y(_2385_));
 sg13g2_xnor2_1 _6351_ (.Y(_2386_),
    .A(_1579_),
    .B(_2384_));
 sg13g2_o21ai_1 _6352_ (.B1(net1310),
    .Y(_2387_),
    .A1(_2378_),
    .A2(_2386_));
 sg13g2_a21o_1 _6353_ (.A2(_2386_),
    .A1(_2378_),
    .B1(_2387_),
    .X(_2388_));
 sg13g2_o21ai_1 _6354_ (.B1(_2388_),
    .Y(_2389_),
    .A1(_2376_),
    .A2(_2377_));
 sg13g2_mux2_1 _6355_ (.A0(net473),
    .A1(_2389_),
    .S(net1249),
    .X(_0309_));
 sg13g2_a21oi_1 _6356_ (.A1(_2378_),
    .A2(_2386_),
    .Y(_2390_),
    .B1(_2385_));
 sg13g2_a22oi_1 _6357_ (.Y(_2391_),
    .B1(net1263),
    .B2(_0050_),
    .A2(net1270),
    .A1(_3174_));
 sg13g2_o21ai_1 _6358_ (.B1(_2391_),
    .Y(_2392_),
    .A1(\dtop.vtop.dphases[2][9] ),
    .A2(_1551_));
 sg13g2_nor2_1 _6359_ (.A(\dtop.vtop.pipeline.nstep[0] ),
    .B(_2392_),
    .Y(_2393_));
 sg13g2_a21oi_1 _6360_ (.A1(\dtop.vtop.pipeline.nstep[0] ),
    .A2(_2381_),
    .Y(_2394_),
    .B1(_2393_));
 sg13g2_nor2_1 _6361_ (.A(net1352),
    .B(_2394_),
    .Y(_2395_));
 sg13g2_nor2b_1 _6362_ (.A(_2359_),
    .B_N(net1352),
    .Y(_2396_));
 sg13g2_nor3_1 _6363_ (.A(_1596_),
    .B(_2395_),
    .C(_2396_),
    .Y(_2397_));
 sg13g2_o21ai_1 _6364_ (.B1(_1596_),
    .Y(_2398_),
    .A1(_2395_),
    .A2(_2396_));
 sg13g2_nor2b_1 _6365_ (.A(_2397_),
    .B_N(_2398_),
    .Y(_2399_));
 sg13g2_nand2_1 _6366_ (.Y(_2400_),
    .A(net1262),
    .B(_2310_));
 sg13g2_mux2_1 _6367_ (.A0(_0018_),
    .A1(net1403),
    .S(net1259),
    .X(_2401_));
 sg13g2_nor2b_1 _6368_ (.A(net1247),
    .B_N(_2401_),
    .Y(_2402_));
 sg13g2_a21oi_1 _6369_ (.A1(net1247),
    .A2(_2347_),
    .Y(_2403_),
    .B1(_2402_));
 sg13g2_o21ai_1 _6370_ (.B1(_2400_),
    .Y(_2404_),
    .A1(net1262),
    .A2(_2403_));
 sg13g2_or3_1 _6371_ (.A(_0051_),
    .B(net1240),
    .C(_2404_),
    .X(_2405_));
 sg13g2_o21ai_1 _6372_ (.B1(_2404_),
    .Y(_2406_),
    .A1(_0051_),
    .A2(net1240));
 sg13g2_and2_1 _6373_ (.A(_2405_),
    .B(_2406_),
    .X(_2407_));
 sg13g2_o21ai_1 _6374_ (.B1(_2407_),
    .Y(_2408_),
    .A1(_2373_),
    .A2(_2376_));
 sg13g2_or3_1 _6375_ (.A(_2373_),
    .B(_2376_),
    .C(_2407_),
    .X(_2409_));
 sg13g2_a21o_1 _6376_ (.A2(_2409_),
    .A1(_2408_),
    .B1(net1310),
    .X(_2410_));
 sg13g2_xnor2_1 _6377_ (.Y(_2411_),
    .A(_2390_),
    .B(_2399_));
 sg13g2_o21ai_1 _6378_ (.B1(_2410_),
    .Y(_2412_),
    .A1(net1297),
    .A2(_2411_));
 sg13g2_nor2_1 _6379_ (.A(net466),
    .B(net1249),
    .Y(_2413_));
 sg13g2_a21oi_1 _6380_ (.A1(net1249),
    .A2(_2412_),
    .Y(_0310_),
    .B1(_2413_));
 sg13g2_nor2_1 _6381_ (.A(net476),
    .B(net1249),
    .Y(_2414_));
 sg13g2_nand2_1 _6382_ (.Y(_2415_),
    .A(net1418),
    .B(_2305_));
 sg13g2_nor2_1 _6383_ (.A(_0016_),
    .B(net1260),
    .Y(_2416_));
 sg13g2_a21oi_1 _6384_ (.A1(_3129_),
    .A2(net1260),
    .Y(_2417_),
    .B1(_2416_));
 sg13g2_mux2_1 _6385_ (.A0(_2417_),
    .A1(_2369_),
    .S(net1246),
    .X(_2418_));
 sg13g2_mux2_1 _6386_ (.A0(_2330_),
    .A1(_2418_),
    .S(_2242_),
    .X(_2419_));
 sg13g2_nor2_1 _6387_ (.A(_2415_),
    .B(_2419_),
    .Y(_2420_));
 sg13g2_xnor2_1 _6388_ (.Y(_2421_),
    .A(_2415_),
    .B(_2419_));
 sg13g2_nand3_1 _6389_ (.B(_2408_),
    .C(_2421_),
    .A(_2405_),
    .Y(_2422_));
 sg13g2_a21oi_1 _6390_ (.A1(_2405_),
    .A2(_2408_),
    .Y(_2423_),
    .B1(_2421_));
 sg13g2_nor2_1 _6391_ (.A(net1310),
    .B(_2423_),
    .Y(_2424_));
 sg13g2_nand2b_1 _6392_ (.Y(_2425_),
    .B(net1270),
    .A_N(\dtop.vtop.dphases[1][10] ));
 sg13g2_o21ai_1 _6393_ (.B1(_2425_),
    .Y(_2426_),
    .A1(\dtop.vtop.dphases[2][10] ),
    .A2(_1551_));
 sg13g2_a21oi_2 _6394_ (.B1(_2426_),
    .Y(_2427_),
    .A2(net1263),
    .A1(_0053_));
 sg13g2_nor2_1 _6395_ (.A(net1350),
    .B(_2392_),
    .Y(_2428_));
 sg13g2_a21oi_1 _6396_ (.A1(net1350),
    .A2(_2427_),
    .Y(_2429_),
    .B1(_2428_));
 sg13g2_mux2_1 _6397_ (.A0(_2429_),
    .A1(_2383_),
    .S(net1352),
    .X(_2430_));
 sg13g2_nor2_1 _6398_ (.A(_1574_),
    .B(_2430_),
    .Y(_2431_));
 sg13g2_xor2_1 _6399_ (.B(_2430_),
    .A(_1574_),
    .X(_2432_));
 sg13g2_o21ai_1 _6400_ (.B1(_2398_),
    .Y(_2433_),
    .A1(_2390_),
    .A2(_2397_));
 sg13g2_o21ai_1 _6401_ (.B1(net1308),
    .Y(_2434_),
    .A1(_2432_),
    .A2(_2433_));
 sg13g2_a21oi_1 _6402_ (.A1(_2432_),
    .A2(_2433_),
    .Y(_2435_),
    .B1(_2434_));
 sg13g2_a21oi_2 _6403_ (.B1(_2435_),
    .Y(_2436_),
    .A2(_2424_),
    .A1(_2422_));
 sg13g2_a21oi_1 _6404_ (.A1(net1249),
    .A2(_2436_),
    .Y(_0311_),
    .B1(_2414_));
 sg13g2_nor2_1 _6405_ (.A(net468),
    .B(net1250),
    .Y(_2437_));
 sg13g2_mux2_1 _6406_ (.A0(_0000_),
    .A1(net1401),
    .S(net1259),
    .X(_2438_));
 sg13g2_mux2_1 _6407_ (.A0(_2438_),
    .A1(_2401_),
    .S(net1247),
    .X(_2439_));
 sg13g2_mux2_1 _6408_ (.A0(_2348_),
    .A1(_2439_),
    .S(_2242_),
    .X(_2440_));
 sg13g2_nor3_1 _6409_ (.A(_0055_),
    .B(net1240),
    .C(_2440_),
    .Y(_2441_));
 sg13g2_o21ai_1 _6410_ (.B1(_2440_),
    .Y(_2442_),
    .A1(_0055_),
    .A2(net1240));
 sg13g2_nor2b_1 _6411_ (.A(_2441_),
    .B_N(_2442_),
    .Y(_2443_));
 sg13g2_o21ai_1 _6412_ (.B1(_2443_),
    .Y(_2444_),
    .A1(_2420_),
    .A2(_2423_));
 sg13g2_nor3_1 _6413_ (.A(_2420_),
    .B(_2423_),
    .C(_2443_),
    .Y(_2445_));
 sg13g2_nor2_1 _6414_ (.A(net1310),
    .B(_2445_),
    .Y(_2446_));
 sg13g2_a21oi_2 _6415_ (.B1(_2431_),
    .Y(_2447_),
    .A2(_2433_),
    .A1(_2432_));
 sg13g2_nor2_1 _6416_ (.A(net1352),
    .B(_2427_),
    .Y(_2448_));
 sg13g2_a21o_1 _6417_ (.A2(_2394_),
    .A1(net1352),
    .B1(_2448_),
    .X(_2449_));
 sg13g2_nor2_1 _6418_ (.A(_1621_),
    .B(_2449_),
    .Y(_2450_));
 sg13g2_and2_1 _6419_ (.A(_1621_),
    .B(_2449_),
    .X(_2451_));
 sg13g2_or2_1 _6420_ (.X(_2452_),
    .B(_2451_),
    .A(_2450_));
 sg13g2_nor2_1 _6421_ (.A(_2447_),
    .B(_2451_),
    .Y(_2453_));
 sg13g2_or2_1 _6422_ (.X(_2454_),
    .B(_2452_),
    .A(_2447_));
 sg13g2_a21oi_1 _6423_ (.A1(_2447_),
    .A2(_2452_),
    .Y(_2455_),
    .B1(net1297));
 sg13g2_a22oi_1 _6424_ (.Y(_2456_),
    .B1(_2454_),
    .B2(_2455_),
    .A2(_2446_),
    .A1(_2444_));
 sg13g2_a21oi_1 _6425_ (.A1(net1250),
    .A2(_2456_),
    .Y(_0312_),
    .B1(_2437_));
 sg13g2_nor2b_1 _6426_ (.A(_2441_),
    .B_N(_2444_),
    .Y(_2457_));
 sg13g2_nand2_2 _6427_ (.Y(_2458_),
    .A(\dtop.vtop.logo.addr[10] ),
    .B(_2305_));
 sg13g2_nor2_1 _6428_ (.A(_3128_),
    .B(net1248),
    .Y(_2459_));
 sg13g2_a21oi_1 _6429_ (.A1(_0014_),
    .A2(_2285_),
    .Y(_2460_),
    .B1(_2459_));
 sg13g2_nand2_1 _6430_ (.Y(_2461_),
    .A(net1246),
    .B(_2417_));
 sg13g2_o21ai_1 _6431_ (.B1(_2461_),
    .Y(_2462_),
    .A1(_2287_),
    .A2(_2460_));
 sg13g2_mux2_1 _6432_ (.A0(_2370_),
    .A1(_2462_),
    .S(_2242_),
    .X(_2463_));
 sg13g2_or2_1 _6433_ (.X(_2464_),
    .B(_2463_),
    .A(_2458_));
 sg13g2_and2_1 _6434_ (.A(_2458_),
    .B(_2463_),
    .X(_2465_));
 sg13g2_xor2_1 _6435_ (.B(_2463_),
    .A(_2458_),
    .X(_2466_));
 sg13g2_xnor2_1 _6436_ (.Y(_2467_),
    .A(_2457_),
    .B(_2466_));
 sg13g2_nand2_1 _6437_ (.Y(_2468_),
    .A(net1296),
    .B(_2467_));
 sg13g2_a21o_1 _6438_ (.A2(_2429_),
    .A1(net1352),
    .B1(_2448_),
    .X(_2469_));
 sg13g2_xor2_1 _6439_ (.B(_2469_),
    .A(_1569_),
    .X(_2470_));
 sg13g2_nor3_1 _6440_ (.A(_2450_),
    .B(_2453_),
    .C(_2470_),
    .Y(_2471_));
 sg13g2_o21ai_1 _6441_ (.B1(_2470_),
    .Y(_2472_),
    .A1(_2450_),
    .A2(_2453_));
 sg13g2_nand2_1 _6442_ (.Y(_2473_),
    .A(net1308),
    .B(_2472_));
 sg13g2_o21ai_1 _6443_ (.B1(_2468_),
    .Y(_2474_),
    .A1(_2471_),
    .A2(_2473_));
 sg13g2_mux2_1 _6444_ (.A0(net455),
    .A1(_2474_),
    .S(net1249),
    .X(_0313_));
 sg13g2_o21ai_1 _6445_ (.B1(_2464_),
    .Y(_2475_),
    .A1(_2457_),
    .A2(_2465_));
 sg13g2_or2_1 _6446_ (.X(_2476_),
    .B(net1260),
    .A(_0059_));
 sg13g2_o21ai_1 _6447_ (.B1(_2476_),
    .Y(_2477_),
    .A1(net1398),
    .A2(net1248));
 sg13g2_o21ai_1 _6448_ (.B1(_2242_),
    .Y(_2478_),
    .A1(net1247),
    .A2(_2477_));
 sg13g2_a21oi_1 _6449_ (.A1(net1247),
    .A2(_2438_),
    .Y(_2479_),
    .B1(_2478_));
 sg13g2_a21oi_1 _6450_ (.A1(net1262),
    .A2(_2403_),
    .Y(_2480_),
    .B1(_2479_));
 sg13g2_nor3_1 _6451_ (.A(_0080_),
    .B(_2306_),
    .C(_2480_),
    .Y(_2481_));
 sg13g2_o21ai_1 _6452_ (.B1(_2480_),
    .Y(_2482_),
    .A1(_0080_),
    .A2(net1240));
 sg13g2_nand2b_1 _6453_ (.Y(_2483_),
    .B(_2482_),
    .A_N(_2481_));
 sg13g2_inv_1 _6454_ (.Y(_2484_),
    .A(_2483_));
 sg13g2_xnor2_1 _6455_ (.Y(_2485_),
    .A(_2475_),
    .B(_2483_));
 sg13g2_o21ai_1 _6456_ (.B1(_2472_),
    .Y(_2486_),
    .A1(_1569_),
    .A2(_2469_));
 sg13g2_or2_1 _6457_ (.X(_2487_),
    .B(_2427_),
    .A(_1629_));
 sg13g2_nand2_1 _6458_ (.Y(_2488_),
    .A(_1629_),
    .B(_2427_));
 sg13g2_nand2_1 _6459_ (.Y(_2489_),
    .A(_2487_),
    .B(_2488_));
 sg13g2_nor2_1 _6460_ (.A(net1308),
    .B(_2485_),
    .Y(_2490_));
 sg13g2_xor2_1 _6461_ (.B(_2489_),
    .A(_2486_),
    .X(_2491_));
 sg13g2_a21oi_2 _6462_ (.B1(_2490_),
    .Y(_2492_),
    .A2(_2491_),
    .A1(net1308));
 sg13g2_mux2_1 _6463_ (.A0(net451),
    .A1(_2492_),
    .S(net1249),
    .X(_0314_));
 sg13g2_a21oi_1 _6464_ (.A1(_2475_),
    .A2(_2484_),
    .Y(_2493_),
    .B1(_2481_));
 sg13g2_nor3_1 _6465_ (.A(_0003_),
    .B(_1533_),
    .C(_2306_),
    .Y(_2494_));
 sg13g2_nand2_1 _6466_ (.Y(_2495_),
    .A(_0090_),
    .B(net1248));
 sg13g2_o21ai_1 _6467_ (.B1(_2495_),
    .Y(_2496_),
    .A1(_3127_),
    .A2(net1248));
 sg13g2_a21oi_1 _6468_ (.A1(net1246),
    .A2(_2460_),
    .Y(_2497_),
    .B1(net1262));
 sg13g2_o21ai_1 _6469_ (.B1(_2497_),
    .Y(_2498_),
    .A1(net1246),
    .A2(_2496_));
 sg13g2_nand2_1 _6470_ (.Y(_2499_),
    .A(_2245_),
    .B(_2498_));
 sg13g2_a21oi_1 _6471_ (.A1(net1261),
    .A2(_2418_),
    .Y(_2500_),
    .B1(_2499_));
 sg13g2_nand2_1 _6472_ (.Y(_2501_),
    .A(_2494_),
    .B(_2500_));
 sg13g2_xnor2_1 _6473_ (.Y(_2502_),
    .A(_2494_),
    .B(_2500_));
 sg13g2_xor2_1 _6474_ (.B(_2502_),
    .A(_2493_),
    .X(_2503_));
 sg13g2_nand2_1 _6475_ (.Y(_2504_),
    .A(net1296),
    .B(_2503_));
 sg13g2_xnor2_1 _6476_ (.Y(_2505_),
    .A(_1564_),
    .B(_2427_));
 sg13g2_nand2_1 _6477_ (.Y(_2506_),
    .A(_2486_),
    .B(_2487_));
 sg13g2_a21oi_1 _6478_ (.A1(_2488_),
    .A2(_2506_),
    .Y(_2507_),
    .B1(_2505_));
 sg13g2_nand3_1 _6479_ (.B(_2505_),
    .C(_2506_),
    .A(_2488_),
    .Y(_2508_));
 sg13g2_nand2_1 _6480_ (.Y(_2509_),
    .A(net1308),
    .B(_2508_));
 sg13g2_o21ai_1 _6481_ (.B1(_2504_),
    .Y(_2510_),
    .A1(_2507_),
    .A2(_2509_));
 sg13g2_mux2_1 _6482_ (.A0(net482),
    .A1(_2510_),
    .S(_2214_),
    .X(_0315_));
 sg13g2_nand2_1 _6483_ (.Y(_2511_),
    .A(_0062_),
    .B(net1248));
 sg13g2_o21ai_1 _6484_ (.B1(_2511_),
    .Y(_2512_),
    .A1(_3126_),
    .A2(net1248));
 sg13g2_a21oi_1 _6485_ (.A1(net1246),
    .A2(_2477_),
    .Y(_2513_),
    .B1(net1261));
 sg13g2_o21ai_1 _6486_ (.B1(_2513_),
    .Y(_2514_),
    .A1(net1246),
    .A2(_2512_));
 sg13g2_nand2_1 _6487_ (.Y(_2515_),
    .A(_2245_),
    .B(_2514_));
 sg13g2_a21oi_1 _6488_ (.A1(net1261),
    .A2(_2439_),
    .Y(_2516_),
    .B1(_2515_));
 sg13g2_o21ai_1 _6489_ (.B1(_2501_),
    .Y(_2517_),
    .A1(_2493_),
    .A2(_2502_));
 sg13g2_xnor2_1 _6490_ (.Y(_2518_),
    .A(_2516_),
    .B(_2517_));
 sg13g2_nand2b_1 _6491_ (.Y(_2519_),
    .B(net1296),
    .A_N(_2518_));
 sg13g2_a21oi_1 _6492_ (.A1(_1564_),
    .A2(_2427_),
    .Y(_2520_),
    .B1(_2507_));
 sg13g2_xor2_1 _6493_ (.B(_2427_),
    .A(_1558_),
    .X(_2521_));
 sg13g2_xnor2_1 _6494_ (.Y(_2522_),
    .A(_2520_),
    .B(_2521_));
 sg13g2_o21ai_1 _6495_ (.B1(_2519_),
    .Y(_2523_),
    .A1(net1296),
    .A2(_2522_));
 sg13g2_mux2_1 _6496_ (.A0(net465),
    .A1(_2523_),
    .S(net1249),
    .X(_0316_));
 sg13g2_nand4_1 _6497_ (.B(\dtop.vtop.pipeline.wave_index[1] ),
    .C(net1307),
    .A(_3147_),
    .Y(_2524_),
    .D(_2017_));
 sg13g2_nand2_1 _6498_ (.Y(_2525_),
    .A(_1880_),
    .B(_2524_));
 sg13g2_nand2_1 _6499_ (.Y(_2526_),
    .A(_2225_),
    .B(net1147));
 sg13g2_o21ai_1 _6500_ (.B1(_2526_),
    .Y(_0317_),
    .A1(_3161_),
    .A2(net1147));
 sg13g2_mux2_1 _6501_ (.A0(net477),
    .A1(_2255_),
    .S(net1147),
    .X(_0318_));
 sg13g2_mux2_1 _6502_ (.A0(net457),
    .A1(_2268_),
    .S(net1147),
    .X(_0319_));
 sg13g2_nand2_1 _6503_ (.Y(_2527_),
    .A(_2281_),
    .B(net1148));
 sg13g2_o21ai_1 _6504_ (.B1(_2527_),
    .Y(_0320_),
    .A1(_3167_),
    .A2(net1148));
 sg13g2_nor2_1 _6505_ (.A(net495),
    .B(net1148),
    .Y(_2528_));
 sg13g2_a21oi_1 _6506_ (.A1(_2301_),
    .A2(net1147),
    .Y(_0321_),
    .B1(_2528_));
 sg13g2_mux2_1 _6507_ (.A0(net522),
    .A1(_2327_),
    .S(net1147),
    .X(_0322_));
 sg13g2_mux2_1 _6508_ (.A0(net454),
    .A1(_2345_),
    .S(net1147),
    .X(_0323_));
 sg13g2_mux2_1 _6509_ (.A0(net458),
    .A1(_2366_),
    .S(net1147),
    .X(_0324_));
 sg13g2_mux2_1 _6510_ (.A0(net486),
    .A1(_2389_),
    .S(net1146),
    .X(_0325_));
 sg13g2_nor2_1 _6511_ (.A(net510),
    .B(net1146),
    .Y(_2529_));
 sg13g2_a21oi_1 _6512_ (.A1(_2412_),
    .A2(net1146),
    .Y(_0326_),
    .B1(_2529_));
 sg13g2_nor2_1 _6513_ (.A(net459),
    .B(net1146),
    .Y(_2530_));
 sg13g2_a21oi_1 _6514_ (.A1(_2436_),
    .A2(net1146),
    .Y(_0327_),
    .B1(_2530_));
 sg13g2_nor2_1 _6515_ (.A(net431),
    .B(net1148),
    .Y(_2531_));
 sg13g2_a21oi_1 _6516_ (.A1(_2456_),
    .A2(net1148),
    .Y(_0328_),
    .B1(_2531_));
 sg13g2_mux2_1 _6517_ (.A0(net504),
    .A1(_2474_),
    .S(net1148),
    .X(_0329_));
 sg13g2_mux2_1 _6518_ (.A0(net483),
    .A1(_2492_),
    .S(net1146),
    .X(_0330_));
 sg13g2_mux2_1 _6519_ (.A0(net453),
    .A1(_2510_),
    .S(net1146),
    .X(_0331_));
 sg13g2_mux2_1 _6520_ (.A0(net509),
    .A1(_2523_),
    .S(net1146),
    .X(_0332_));
 sg13g2_and2_1 _6521_ (.A(net1430),
    .B(net336),
    .X(_0333_));
 sg13g2_nand2_1 _6522_ (.Y(_2532_),
    .A(_3147_),
    .B(_3148_));
 sg13g2_nand2_1 _6523_ (.Y(_2533_),
    .A(\dtop.vtop.pipeline.cosappr_acc[3] ),
    .B(net1302));
 sg13g2_nor2_1 _6524_ (.A(net1210),
    .B(_2533_),
    .Y(_2534_));
 sg13g2_xnor2_1 _6525_ (.Y(_2535_),
    .A(net1210),
    .B(_2533_));
 sg13g2_nand2_1 _6526_ (.Y(_2536_),
    .A(\dtop.vtop.pipeline.cosappr_acc[2] ),
    .B(net1302));
 sg13g2_nor2_1 _6527_ (.A(net1192),
    .B(_2536_),
    .Y(_2537_));
 sg13g2_nand2_1 _6528_ (.Y(_2538_),
    .A(net376),
    .B(net1302));
 sg13g2_nand2b_1 _6529_ (.Y(_2539_),
    .B(net1201),
    .A_N(_2538_));
 sg13g2_and3_1 _6530_ (.X(_2540_),
    .A(\dtop.vtop.pipeline.cosappr_acc[0] ),
    .B(net1198),
    .C(net1302));
 sg13g2_xnor2_1 _6531_ (.Y(_2541_),
    .A(net1201),
    .B(_2538_));
 sg13g2_nand2_1 _6532_ (.Y(_2542_),
    .A(_2540_),
    .B(_2541_));
 sg13g2_xnor2_1 _6533_ (.Y(_2543_),
    .A(net1192),
    .B(_2536_));
 sg13g2_a21oi_1 _6534_ (.A1(_2539_),
    .A2(_2542_),
    .Y(_2544_),
    .B1(_2543_));
 sg13g2_nor2_1 _6535_ (.A(_2537_),
    .B(_2544_),
    .Y(_2545_));
 sg13g2_nor2_1 _6536_ (.A(_2535_),
    .B(_2545_),
    .Y(_2546_));
 sg13g2_xor2_1 _6537_ (.B(_2545_),
    .A(_2535_),
    .X(_2547_));
 sg13g2_mux2_1 _6538_ (.A0(net570),
    .A1(_2547_),
    .S(_2027_),
    .X(_0334_));
 sg13g2_nand2_1 _6539_ (.Y(_2548_),
    .A(\dtop.vtop.pipeline.cosappr_acc[4] ),
    .B(net1302));
 sg13g2_nor2_1 _6540_ (.A(net1186),
    .B(_2548_),
    .Y(_2549_));
 sg13g2_xnor2_1 _6541_ (.Y(_2550_),
    .A(net1186),
    .B(_2548_));
 sg13g2_nor2_1 _6542_ (.A(_2534_),
    .B(_2546_),
    .Y(_2551_));
 sg13g2_nor2_1 _6543_ (.A(_2550_),
    .B(_2551_),
    .Y(_2552_));
 sg13g2_xor2_1 _6544_ (.B(_2551_),
    .A(_2550_),
    .X(_2553_));
 sg13g2_mux2_1 _6545_ (.A0(net598),
    .A1(_2553_),
    .S(net1151),
    .X(_0335_));
 sg13g2_and2_1 _6546_ (.A(\dtop.vtop.pipeline.cosappr_acc[5] ),
    .B(net1303),
    .X(_2554_));
 sg13g2_xnor2_1 _6547_ (.Y(_2555_),
    .A(net1216),
    .B(_2554_));
 sg13g2_nor2_1 _6548_ (.A(_2549_),
    .B(_2552_),
    .Y(_2556_));
 sg13g2_nor2_1 _6549_ (.A(_2555_),
    .B(_2556_),
    .Y(_2557_));
 sg13g2_xor2_1 _6550_ (.B(_2556_),
    .A(_2555_),
    .X(_2558_));
 sg13g2_mux2_1 _6551_ (.A0(net544),
    .A1(_2558_),
    .S(net1151),
    .X(_0336_));
 sg13g2_nand2_1 _6552_ (.Y(_2559_),
    .A(\dtop.vtop.pipeline.cosappr_acc[6] ),
    .B(net1303));
 sg13g2_inv_1 _6553_ (.Y(_2560_),
    .A(_2559_));
 sg13g2_xnor2_1 _6554_ (.Y(_2561_),
    .A(net1180),
    .B(_2560_));
 sg13g2_a21oi_1 _6555_ (.A1(net1216),
    .A2(_2554_),
    .Y(_2562_),
    .B1(_2557_));
 sg13g2_nor2_1 _6556_ (.A(_2561_),
    .B(_2562_),
    .Y(_2563_));
 sg13g2_xor2_1 _6557_ (.B(_2562_),
    .A(_2561_),
    .X(_2564_));
 sg13g2_nor2_1 _6558_ (.A(net1149),
    .B(_2564_),
    .Y(_2565_));
 sg13g2_a21oi_1 _6559_ (.A1(_3156_),
    .A2(net1149),
    .Y(_0337_),
    .B1(_2565_));
 sg13g2_nor2_1 _6560_ (.A(net562),
    .B(net1151),
    .Y(_2566_));
 sg13g2_nand2_1 _6561_ (.Y(_2567_),
    .A(net424),
    .B(net1302));
 sg13g2_a21oi_1 _6562_ (.A1(net1180),
    .A2(_2560_),
    .Y(_2568_),
    .B1(_2563_));
 sg13g2_nor2_1 _6563_ (.A(_2567_),
    .B(_2568_),
    .Y(_2569_));
 sg13g2_xnor2_1 _6564_ (.Y(_2570_),
    .A(_2567_),
    .B(_2568_));
 sg13g2_a21oi_1 _6565_ (.A1(net1151),
    .A2(_2570_),
    .Y(_0338_),
    .B1(_2566_));
 sg13g2_nand2_1 _6566_ (.Y(_2571_),
    .A(net452),
    .B(net1302));
 sg13g2_mux2_2 _6567_ (.A0(_2571_),
    .A1(net452),
    .S(_2569_),
    .X(_2572_));
 sg13g2_nor2_1 _6568_ (.A(net528),
    .B(net1151),
    .Y(_2573_));
 sg13g2_a21oi_1 _6569_ (.A1(net1151),
    .A2(_2572_),
    .Y(_0339_),
    .B1(_2573_));
 sg13g2_nor2b_2 _6570_ (.A(net1273),
    .B_N(net1303),
    .Y(_2574_));
 sg13g2_o21ai_1 _6571_ (.B1(net1303),
    .Y(_2575_),
    .A1(net1290),
    .A2(net1287));
 sg13g2_nand2_1 _6572_ (.Y(_2576_),
    .A(\dtop.vtop.pipeline.zg_acc[0] ),
    .B(_2574_));
 sg13g2_nor2_1 _6573_ (.A(_1804_),
    .B(_2576_),
    .Y(_2577_));
 sg13g2_xor2_1 _6574_ (.B(_2576_),
    .A(_1804_),
    .X(_2578_));
 sg13g2_mux2_1 _6575_ (.A0(net484),
    .A1(_2578_),
    .S(net1150),
    .X(_0340_));
 sg13g2_nand2_1 _6576_ (.Y(_2579_),
    .A(\dtop.vtop.pipeline.zg_acc[1] ),
    .B(_2574_));
 sg13g2_nor2b_1 _6577_ (.A(_2579_),
    .B_N(_1831_),
    .Y(_2580_));
 sg13g2_xnor2_1 _6578_ (.Y(_2581_),
    .A(_1831_),
    .B(_2579_));
 sg13g2_xnor2_1 _6579_ (.Y(_2582_),
    .A(_2577_),
    .B(_2581_));
 sg13g2_nor2_1 _6580_ (.A(net517),
    .B(net1150),
    .Y(_2583_));
 sg13g2_a21oi_1 _6581_ (.A1(net1150),
    .A2(_2582_),
    .Y(_0341_),
    .B1(_2583_));
 sg13g2_a21oi_1 _6582_ (.A1(_2577_),
    .A2(_2581_),
    .Y(_2584_),
    .B1(_2580_));
 sg13g2_nand2_1 _6583_ (.Y(_2585_),
    .A(\dtop.vtop.pipeline.zg_acc[2] ),
    .B(_2574_));
 sg13g2_or2_1 _6584_ (.X(_2586_),
    .B(_2585_),
    .A(_1843_));
 sg13g2_xnor2_1 _6585_ (.Y(_2587_),
    .A(_1843_),
    .B(_2585_));
 sg13g2_xor2_1 _6586_ (.B(_2587_),
    .A(_2584_),
    .X(_2588_));
 sg13g2_mux2_1 _6587_ (.A0(net533),
    .A1(_2588_),
    .S(net1150),
    .X(_0342_));
 sg13g2_nand2_1 _6588_ (.Y(_2589_),
    .A(\dtop.vtop.pipeline.zg_acc[3] ),
    .B(_2574_));
 sg13g2_nor2_1 _6589_ (.A(_1851_),
    .B(_2589_),
    .Y(_2590_));
 sg13g2_nand2_1 _6590_ (.Y(_2591_),
    .A(_1851_),
    .B(_2589_));
 sg13g2_nand2b_1 _6591_ (.Y(_2592_),
    .B(_2591_),
    .A_N(_2590_));
 sg13g2_o21ai_1 _6592_ (.B1(_2586_),
    .Y(_2593_),
    .A1(_2584_),
    .A2(_2587_));
 sg13g2_xnor2_1 _6593_ (.Y(_2594_),
    .A(_2592_),
    .B(_2593_));
 sg13g2_mux2_1 _6594_ (.A0(net612),
    .A1(_2594_),
    .S(net1150),
    .X(_0343_));
 sg13g2_a21oi_1 _6595_ (.A1(_2591_),
    .A2(_2593_),
    .Y(_2595_),
    .B1(_2590_));
 sg13g2_nand2_1 _6596_ (.Y(_2596_),
    .A(\dtop.vtop.pipeline.zg_acc[4] ),
    .B(_2574_));
 sg13g2_or2_1 _6597_ (.X(_2597_),
    .B(_2596_),
    .A(_1857_));
 sg13g2_and2_1 _6598_ (.A(_1857_),
    .B(_2596_),
    .X(_2598_));
 sg13g2_xor2_1 _6599_ (.B(_2596_),
    .A(_1857_),
    .X(_2599_));
 sg13g2_xnor2_1 _6600_ (.Y(_2600_),
    .A(_2595_),
    .B(_2599_));
 sg13g2_mux2_1 _6601_ (.A0(net649),
    .A1(_2600_),
    .S(net1150),
    .X(_0344_));
 sg13g2_o21ai_1 _6602_ (.B1(_2597_),
    .Y(_2601_),
    .A1(_2595_),
    .A2(_2598_));
 sg13g2_nand2_1 _6603_ (.Y(_2602_),
    .A(\dtop.vtop.pipeline.zg_acc[5] ),
    .B(_2574_));
 sg13g2_nand2_1 _6604_ (.Y(_2603_),
    .A(_1861_),
    .B(_2602_));
 sg13g2_nor2_1 _6605_ (.A(_1861_),
    .B(_2602_),
    .Y(_2604_));
 sg13g2_xnor2_1 _6606_ (.Y(_2605_),
    .A(_1861_),
    .B(_2602_));
 sg13g2_xnor2_1 _6607_ (.Y(_2606_),
    .A(_2601_),
    .B(_2605_));
 sg13g2_mux2_1 _6608_ (.A0(net616),
    .A1(_2606_),
    .S(net1150),
    .X(_0345_));
 sg13g2_nor2_1 _6609_ (.A(_0058_),
    .B(_2575_),
    .Y(_2607_));
 sg13g2_nor2b_1 _6610_ (.A(_1863_),
    .B_N(_2607_),
    .Y(_2608_));
 sg13g2_xnor2_1 _6611_ (.Y(_2609_),
    .A(_1863_),
    .B(_2607_));
 sg13g2_o21ai_1 _6612_ (.B1(_2603_),
    .Y(_2610_),
    .A1(_2601_),
    .A2(_2604_));
 sg13g2_inv_1 _6613_ (.Y(_2611_),
    .A(_2610_));
 sg13g2_xnor2_1 _6614_ (.Y(_2612_),
    .A(_2609_),
    .B(_2610_));
 sg13g2_nor2_1 _6615_ (.A(net1149),
    .B(_2612_),
    .Y(_2613_));
 sg13g2_a21oi_1 _6616_ (.A1(_3123_),
    .A2(net1149),
    .Y(_0346_),
    .B1(_2613_));
 sg13g2_nor3_1 _6617_ (.A(_0061_),
    .B(_1876_),
    .C(_2575_),
    .Y(_2614_));
 sg13g2_o21ai_1 _6618_ (.B1(_1876_),
    .Y(_2615_),
    .A1(_0061_),
    .A2(_2575_));
 sg13g2_nor2b_1 _6619_ (.A(_2614_),
    .B_N(_2615_),
    .Y(_2616_));
 sg13g2_a21oi_1 _6620_ (.A1(_2609_),
    .A2(_2611_),
    .Y(_2617_),
    .B1(_2608_));
 sg13g2_xnor2_1 _6621_ (.Y(_2618_),
    .A(_2616_),
    .B(_2617_));
 sg13g2_mux2_1 _6622_ (.A0(net631),
    .A1(_2618_),
    .S(net1151),
    .X(_0347_));
 sg13g2_a22oi_1 _6623_ (.Y(_2619_),
    .B1(_2574_),
    .B2(_3177_),
    .A2(net1273),
    .A1(_1540_));
 sg13g2_nor2_1 _6624_ (.A(net1241),
    .B(_2619_),
    .Y(_2620_));
 sg13g2_xnor2_1 _6625_ (.Y(_2621_),
    .A(net1241),
    .B(_2619_));
 sg13g2_inv_1 _6626_ (.Y(_2622_),
    .A(_2621_));
 sg13g2_nand2_1 _6627_ (.Y(_2623_),
    .A(_2609_),
    .B(_2616_));
 sg13g2_a21oi_1 _6628_ (.A1(_2608_),
    .A2(_2615_),
    .Y(_2624_),
    .B1(_2614_));
 sg13g2_o21ai_1 _6629_ (.B1(_2624_),
    .Y(_2625_),
    .A1(_2610_),
    .A2(_2623_));
 sg13g2_xnor2_1 _6630_ (.Y(_2626_),
    .A(_2621_),
    .B(_2625_));
 sg13g2_nor2_1 _6631_ (.A(net1149),
    .B(_2626_),
    .Y(_2627_));
 sg13g2_a21oi_1 _6632_ (.A1(_3121_),
    .A2(net1149),
    .Y(_0348_),
    .B1(_2627_));
 sg13g2_a21oi_1 _6633_ (.A1(_2622_),
    .A2(_2625_),
    .Y(_2628_),
    .B1(_2620_));
 sg13g2_nor2_1 _6634_ (.A(\dtop.vtop.pipeline.zg_acc[9] ),
    .B(_2575_),
    .Y(_2629_));
 sg13g2_xor2_1 _6635_ (.B(_2629_),
    .A(net1241),
    .X(_2630_));
 sg13g2_xnor2_1 _6636_ (.Y(_2631_),
    .A(_2628_),
    .B(_2630_));
 sg13g2_mux2_1 _6637_ (.A0(net1356),
    .A1(_2631_),
    .S(net1150),
    .X(_0349_));
 sg13g2_a21oi_1 _6638_ (.A1(net527),
    .A2(net1302),
    .Y(_2632_),
    .B1(net1198));
 sg13g2_nor3_1 _6639_ (.A(net1228),
    .B(_2540_),
    .C(_2632_),
    .Y(_2633_));
 sg13g2_a21o_1 _6640_ (.A2(net1228),
    .A1(net527),
    .B1(_2633_),
    .X(_0350_));
 sg13g2_nand2_1 _6641_ (.Y(_2634_),
    .A(net376),
    .B(net1228));
 sg13g2_xnor2_1 _6642_ (.Y(_2635_),
    .A(_2540_),
    .B(_2541_));
 sg13g2_o21ai_1 _6643_ (.B1(_2634_),
    .Y(_0351_),
    .A1(net1228),
    .A2(_2635_));
 sg13g2_and3_1 _6644_ (.X(_2636_),
    .A(_2539_),
    .B(_2542_),
    .C(_2543_));
 sg13g2_nor3_1 _6645_ (.A(net1228),
    .B(_2544_),
    .C(_2636_),
    .Y(_2637_));
 sg13g2_a21o_1 _6646_ (.A2(net1228),
    .A1(net494),
    .B1(_2637_),
    .X(_0352_));
 sg13g2_mux2_1 _6647_ (.A0(net446),
    .A1(_2547_),
    .S(net1176),
    .X(_0353_));
 sg13g2_mux2_1 _6648_ (.A0(net450),
    .A1(_2553_),
    .S(net1176),
    .X(_0354_));
 sg13g2_mux2_1 _6649_ (.A0(net460),
    .A1(_2558_),
    .S(net1176),
    .X(_0355_));
 sg13g2_mux2_1 _6650_ (.A0(net456),
    .A1(_2564_),
    .S(net1177),
    .X(_0356_));
 sg13g2_nand2_1 _6651_ (.Y(_2638_),
    .A(net424),
    .B(net1229));
 sg13g2_o21ai_1 _6652_ (.B1(_2638_),
    .Y(_0357_),
    .A1(net1229),
    .A2(_2570_));
 sg13g2_nand2_1 _6653_ (.Y(_2639_),
    .A(net452),
    .B(net1229));
 sg13g2_o21ai_1 _6654_ (.B1(_2639_),
    .Y(_0358_),
    .A1(net1229),
    .A2(_2572_));
 sg13g2_mux2_1 _6655_ (.A0(net628),
    .A1(_2578_),
    .S(net1176),
    .X(_0359_));
 sg13g2_nand2_1 _6656_ (.Y(_2640_),
    .A(net573),
    .B(net1229));
 sg13g2_o21ai_1 _6657_ (.B1(_2640_),
    .Y(_0360_),
    .A1(net1228),
    .A2(_2582_));
 sg13g2_mux2_1 _6658_ (.A0(net590),
    .A1(_2588_),
    .S(net1176),
    .X(_0361_));
 sg13g2_mux2_1 _6659_ (.A0(net613),
    .A1(_2594_),
    .S(net1176),
    .X(_0362_));
 sg13g2_mux2_1 _6660_ (.A0(net624),
    .A1(_2600_),
    .S(net1176),
    .X(_0363_));
 sg13g2_mux2_1 _6661_ (.A0(net551),
    .A1(_2606_),
    .S(net1177),
    .X(_0364_));
 sg13g2_mux2_1 _6662_ (.A0(net418),
    .A1(_2612_),
    .S(net1176),
    .X(_0365_));
 sg13g2_mux2_1 _6663_ (.A0(net425),
    .A1(_2618_),
    .S(net1177),
    .X(_0366_));
 sg13g2_mux2_1 _6664_ (.A0(net513),
    .A1(_2626_),
    .S(net1177),
    .X(_0367_));
 sg13g2_mux2_1 _6665_ (.A0(net491),
    .A1(_2631_),
    .S(net1177),
    .X(_0368_));
 sg13g2_a21oi_1 _6666_ (.A1(_2017_),
    .A2(net1177),
    .Y(_0369_),
    .B1(net1294));
 sg13g2_nand2_1 _6667_ (.Y(_2641_),
    .A(net1307),
    .B(_2028_));
 sg13g2_nand2_1 _6668_ (.Y(_2642_),
    .A(_3148_),
    .B(_0004_));
 sg13g2_a21oi_1 _6669_ (.A1(_2022_),
    .A2(_2642_),
    .Y(_0370_),
    .B1(_2641_));
 sg13g2_a21oi_1 _6670_ (.A1(net552),
    .A2(_3148_),
    .Y(_2643_),
    .B1(_2023_));
 sg13g2_nor2_1 _6671_ (.A(_2641_),
    .B(net553),
    .Y(_0371_));
 sg13g2_or3_1 _6672_ (.A(net554),
    .B(\dtop.vtop.pipeline.nstep_counter[0] ),
    .C(net1149),
    .X(_2644_));
 sg13g2_or2_1 _6673_ (.X(_2645_),
    .B(_2644_),
    .A(net593));
 sg13g2_or2_1 _6674_ (.X(_2646_),
    .B(_2645_),
    .A(net537));
 sg13g2_nor2_1 _6675_ (.A(net1398),
    .B(_3202_),
    .Y(_2647_));
 sg13g2_xor2_1 _6676_ (.B(_2647_),
    .A(_0030_),
    .X(_2648_));
 sg13g2_nor2_1 _6677_ (.A(net1400),
    .B(_3202_),
    .Y(_2649_));
 sg13g2_xnor2_1 _6678_ (.Y(_2650_),
    .A(\dtop.vtop.pipeline.nstep[0] ),
    .B(_2649_));
 sg13g2_nor2_1 _6679_ (.A(_2648_),
    .B(_2650_),
    .Y(_2651_));
 sg13g2_nor3_1 _6680_ (.A(net492),
    .B(_2646_),
    .C(_2651_),
    .Y(_2652_));
 sg13g2_or2_1 _6681_ (.X(_2653_),
    .B(_2652_),
    .A(\dtop.vtop.pipeline.nstep[0] ));
 sg13g2_nand2_1 _6682_ (.Y(_2654_),
    .A(\dtop.vtop.pipeline.nstep[0] ),
    .B(_2652_));
 sg13g2_nand3_1 _6683_ (.B(net690),
    .C(_2654_),
    .A(net1311),
    .Y(_2655_));
 sg13g2_inv_1 _6684_ (.Y(_0372_),
    .A(_2655_));
 sg13g2_xor2_1 _6685_ (.B(_2654_),
    .A(net1354),
    .X(_2656_));
 sg13g2_nor2_1 _6686_ (.A(net1297),
    .B(_2656_),
    .Y(_0373_));
 sg13g2_nor2_1 _6687_ (.A(\dtop.vtop.pipeline.nstep_counter[0] ),
    .B(_2641_),
    .Y(_2657_));
 sg13g2_a21oi_1 _6688_ (.A1(_3063_),
    .A2(_2029_),
    .Y(_0374_),
    .B1(_2657_));
 sg13g2_o21ai_1 _6689_ (.B1(net554),
    .Y(_2658_),
    .A1(\dtop.vtop.pipeline.nstep_counter[0] ),
    .A2(net1149));
 sg13g2_nand3_1 _6690_ (.B(_2644_),
    .C(net555),
    .A(net1312),
    .Y(_0375_));
 sg13g2_a21oi_1 _6691_ (.A1(net593),
    .A2(_2644_),
    .Y(_2659_),
    .B1(net1299));
 sg13g2_nand2_1 _6692_ (.Y(_0376_),
    .A(_2645_),
    .B(_2659_));
 sg13g2_a21oi_1 _6693_ (.A1(net537),
    .A2(_2645_),
    .Y(_2660_),
    .B1(net1299));
 sg13g2_nand2_1 _6694_ (.Y(_0377_),
    .A(_2646_),
    .B(net538));
 sg13g2_a21o_1 _6695_ (.A2(_2646_),
    .A1(net492),
    .B1(net1299),
    .X(_0378_));
 sg13g2_nor2_1 _6696_ (.A(_0601_),
    .B(net1308),
    .Y(_2661_));
 sg13g2_a21oi_1 _6697_ (.A1(net1308),
    .A2(net1303),
    .Y(_2662_),
    .B1(_2661_));
 sg13g2_mux2_1 _6698_ (.A0(net370),
    .A1(_2225_),
    .S(net1257),
    .X(_0379_));
 sg13g2_mux2_1 _6699_ (.A0(net393),
    .A1(_2255_),
    .S(net1257),
    .X(_0380_));
 sg13g2_mux2_1 _6700_ (.A0(net389),
    .A1(_2268_),
    .S(net1257),
    .X(_0381_));
 sg13g2_mux2_1 _6701_ (.A0(net365),
    .A1(_2281_),
    .S(net1258),
    .X(_0382_));
 sg13g2_nor2_1 _6702_ (.A(net432),
    .B(net1257),
    .Y(_2663_));
 sg13g2_a21oi_1 _6703_ (.A1(_2301_),
    .A2(net1257),
    .Y(_0383_),
    .B1(_2663_));
 sg13g2_mux2_1 _6704_ (.A0(net401),
    .A1(_2327_),
    .S(net1257),
    .X(_0384_));
 sg13g2_mux2_1 _6705_ (.A0(net394),
    .A1(_2345_),
    .S(net1257),
    .X(_0385_));
 sg13g2_mux2_1 _6706_ (.A0(net416),
    .A1(_2366_),
    .S(net1257),
    .X(_0386_));
 sg13g2_mux2_1 _6707_ (.A0(net412),
    .A1(_2389_),
    .S(net1256),
    .X(_0387_));
 sg13g2_nor2_1 _6708_ (.A(net419),
    .B(net1256),
    .Y(_2664_));
 sg13g2_a21oi_1 _6709_ (.A1(_2412_),
    .A2(net1256),
    .Y(_0388_),
    .B1(_2664_));
 sg13g2_nor2_1 _6710_ (.A(net347),
    .B(net1256),
    .Y(_2665_));
 sg13g2_a21oi_1 _6711_ (.A1(_2436_),
    .A2(net1256),
    .Y(_0389_),
    .B1(_2665_));
 sg13g2_nor2_1 _6712_ (.A(net372),
    .B(net1258),
    .Y(_2666_));
 sg13g2_a21oi_1 _6713_ (.A1(_2456_),
    .A2(net1258),
    .Y(_0390_),
    .B1(_2666_));
 sg13g2_mux2_1 _6714_ (.A0(net378),
    .A1(_2474_),
    .S(net1258),
    .X(_0391_));
 sg13g2_mux2_1 _6715_ (.A0(net366),
    .A1(_2492_),
    .S(net1256),
    .X(_0392_));
 sg13g2_mux2_1 _6716_ (.A0(net384),
    .A1(_2510_),
    .S(net1256),
    .X(_0393_));
 sg13g2_mux2_1 _6717_ (.A0(net390),
    .A1(_2523_),
    .S(net1256),
    .X(_0394_));
 sg13g2_nor2_1 _6718_ (.A(_3213_),
    .B(_1191_),
    .Y(_2667_));
 sg13g2_o21ai_1 _6719_ (.B1(_3249_),
    .Y(_2668_),
    .A1(_2467_),
    .A2(_2485_));
 sg13g2_nand2_1 _6720_ (.Y(_2669_),
    .A(_2503_),
    .B(_2668_));
 sg13g2_o21ai_1 _6721_ (.B1(_2669_),
    .Y(_2670_),
    .A1(_3250_),
    .A2(_2503_));
 sg13g2_xor2_1 _6722_ (.B(_2670_),
    .A(_2518_),
    .X(_2671_));
 sg13g2_nor2_1 _6723_ (.A(_3283_),
    .B(_2303_),
    .Y(_2672_));
 sg13g2_o21ai_1 _6724_ (.B1(_2672_),
    .Y(_2673_),
    .A1(net1344),
    .A2(_2671_));
 sg13g2_a21oi_1 _6725_ (.A1(net1344),
    .A2(_2671_),
    .Y(_2674_),
    .B1(_2673_));
 sg13g2_nor2_2 _6726_ (.A(_2667_),
    .B(_2674_),
    .Y(_2675_));
 sg13g2_a21oi_1 _6727_ (.A1(\dtop.enable ),
    .A2(_3249_),
    .Y(_2676_),
    .B1(_3246_));
 sg13g2_a21o_1 _6728_ (.A2(_3246_),
    .A1(_3353_),
    .B1(_2676_),
    .X(_2677_));
 sg13g2_nor2b_2 _6729_ (.A(_2677_),
    .B_N(_3244_),
    .Y(_2678_));
 sg13g2_nand2_1 _6730_ (.Y(_2679_),
    .A(_3240_),
    .B(_2678_));
 sg13g2_or2_1 _6731_ (.X(_2680_),
    .B(_2679_),
    .A(_3238_));
 sg13g2_nor2_1 _6732_ (.A(_3269_),
    .B(_2680_),
    .Y(_2681_));
 sg13g2_and2_1 _6733_ (.A(_3270_),
    .B(_2680_),
    .X(_2682_));
 sg13g2_xor2_1 _6734_ (.B(_2679_),
    .A(_3238_),
    .X(_2683_));
 sg13g2_xnor2_1 _6735_ (.Y(_2684_),
    .A(_3238_),
    .B(_2679_));
 sg13g2_xor2_1 _6736_ (.B(_2678_),
    .A(_3240_),
    .X(_2685_));
 sg13g2_xnor2_1 _6737_ (.Y(_2686_),
    .A(_3240_),
    .B(_2678_));
 sg13g2_xnor2_1 _6738_ (.Y(_2687_),
    .A(_3244_),
    .B(_2677_));
 sg13g2_xor2_1 _6739_ (.B(_2677_),
    .A(_3244_),
    .X(_2688_));
 sg13g2_nor2_2 _6740_ (.A(_2686_),
    .B(net1227),
    .Y(_2689_));
 sg13g2_nand2_2 _6741_ (.Y(_2690_),
    .A(_2685_),
    .B(net1225));
 sg13g2_nand2_1 _6742_ (.Y(_2691_),
    .A(net1361),
    .B(_3250_));
 sg13g2_xor2_1 _6743_ (.B(_2691_),
    .A(_3246_),
    .X(_2692_));
 sg13g2_xnor2_1 _6744_ (.Y(_2693_),
    .A(_3246_),
    .B(_2691_));
 sg13g2_nor2_2 _6745_ (.A(net1227),
    .B(net1243),
    .Y(_2694_));
 sg13g2_nand2_2 _6746_ (.Y(_2695_),
    .A(net1225),
    .B(net1245));
 sg13g2_nor2_2 _6747_ (.A(net1403),
    .B(_0740_),
    .Y(_2696_));
 sg13g2_nand2_1 _6748_ (.Y(_2697_),
    .A(net1401),
    .B(_0051_));
 sg13g2_a22oi_1 _6749_ (.Y(_2698_),
    .B1(_2697_),
    .B2(net1402),
    .A2(_2692_),
    .A1(_1176_));
 sg13g2_xor2_1 _6750_ (.B(_2698_),
    .A(_0023_),
    .X(_2699_));
 sg13g2_nand2_1 _6751_ (.Y(_2700_),
    .A(_2696_),
    .B(_2699_));
 sg13g2_xnor2_1 _6752_ (.Y(_2701_),
    .A(net1362),
    .B(_3249_));
 sg13g2_and2_1 _6753_ (.A(net1425),
    .B(_2701_),
    .X(_2702_));
 sg13g2_xnor2_1 _6754_ (.Y(_2703_),
    .A(\dtop.oct_counter[4] ),
    .B(net1383));
 sg13g2_o21ai_1 _6755_ (.B1(_2703_),
    .Y(_2704_),
    .A1(\dtop.oct_counter[3] ),
    .A2(_3136_));
 sg13g2_o21ai_1 _6756_ (.B1(_2704_),
    .Y(_2705_),
    .A1(_3135_),
    .A2(net1383));
 sg13g2_xnor2_1 _6757_ (.Y(_2706_),
    .A(_0046_),
    .B(_3252_));
 sg13g2_nand2b_1 _6758_ (.Y(_2707_),
    .B(_2705_),
    .A_N(_2706_));
 sg13g2_o21ai_1 _6759_ (.B1(_2707_),
    .Y(_2708_),
    .A1(_3134_),
    .A2(_3252_));
 sg13g2_xor2_1 _6760_ (.B(_2701_),
    .A(net1425),
    .X(_2709_));
 sg13g2_a21oi_1 _6761_ (.A1(_2708_),
    .A2(_2709_),
    .Y(_2710_),
    .B1(_2702_));
 sg13g2_nor2_1 _6762_ (.A(_2700_),
    .B(_2710_),
    .Y(_2711_));
 sg13g2_nand2_1 _6763_ (.Y(_2712_),
    .A(_2700_),
    .B(_2710_));
 sg13g2_nand2b_1 _6764_ (.Y(_2713_),
    .B(_2712_),
    .A_N(_2711_));
 sg13g2_xor2_1 _6765_ (.B(_2698_),
    .A(_0077_),
    .X(_2714_));
 sg13g2_xor2_1 _6766_ (.B(_2709_),
    .A(_2708_),
    .X(_2715_));
 sg13g2_nand3_1 _6767_ (.B(_2714_),
    .C(_2715_),
    .A(_2696_),
    .Y(_2716_));
 sg13g2_a21oi_1 _6768_ (.A1(_2696_),
    .A2(_2714_),
    .Y(_2717_),
    .B1(_2715_));
 sg13g2_nand2_1 _6769_ (.Y(_2718_),
    .A(_0025_),
    .B(_2698_));
 sg13g2_nand2b_1 _6770_ (.Y(_2719_),
    .B(_2706_),
    .A_N(_2705_));
 sg13g2_a221oi_1 _6771_ (.B2(_2706_),
    .C1(_2704_),
    .B1(_0025_),
    .A1(\dtop.oct_counter[3] ),
    .Y(_2720_),
    .A2(_3136_));
 sg13g2_nand2b_1 _6772_ (.Y(_2721_),
    .B(_2720_),
    .A_N(_2698_));
 sg13g2_a21o_1 _6773_ (.A2(_2719_),
    .A1(_2707_),
    .B1(_0025_),
    .X(_2722_));
 sg13g2_nand4_1 _6774_ (.B(_2718_),
    .C(_2721_),
    .A(_2696_),
    .Y(_2723_),
    .D(_2722_));
 sg13g2_a21oi_2 _6775_ (.B1(_2717_),
    .Y(_2724_),
    .A2(_2723_),
    .A1(_2716_));
 sg13g2_xor2_1 _6776_ (.B(_2724_),
    .A(_2713_),
    .X(_2725_));
 sg13g2_nand2_1 _6777_ (.Y(_2726_),
    .A(net1243),
    .B(net1143));
 sg13g2_nor2_2 _6778_ (.A(net1243),
    .B(net1143),
    .Y(_2727_));
 sg13g2_or2_1 _6779_ (.X(_2728_),
    .B(net1144),
    .A(net1243));
 sg13g2_and2_1 _6780_ (.A(net1118),
    .B(net1117),
    .X(_2729_));
 sg13g2_nand2_1 _6781_ (.Y(_2730_),
    .A(net1118),
    .B(_2728_));
 sg13g2_nor2_2 _6782_ (.A(net1225),
    .B(_2727_),
    .Y(_2731_));
 sg13g2_nand2_2 _6783_ (.Y(_2732_),
    .A(net1227),
    .B(net1109));
 sg13g2_nor2_2 _6784_ (.A(_2685_),
    .B(_2694_),
    .Y(_2733_));
 sg13g2_nand2_1 _6785_ (.Y(_2734_),
    .A(net1174),
    .B(_2695_));
 sg13g2_nand2_2 _6786_ (.Y(_2735_),
    .A(_2732_),
    .B(_2733_));
 sg13g2_nand3_1 _6787_ (.B(_2690_),
    .C(_2735_),
    .A(net1155),
    .Y(_2736_));
 sg13g2_a21oi_2 _6788_ (.B1(_2711_),
    .Y(_2737_),
    .A2(_2724_),
    .A1(_2712_));
 sg13g2_nor2_1 _6789_ (.A(_0729_),
    .B(_2737_),
    .Y(_2738_));
 sg13g2_nor2_1 _6790_ (.A(_0059_),
    .B(_0736_),
    .Y(_2739_));
 sg13g2_xnor2_1 _6791_ (.Y(_2740_),
    .A(_0090_),
    .B(_2739_));
 sg13g2_nor2_1 _6792_ (.A(_0020_),
    .B(_3322_),
    .Y(_2741_));
 sg13g2_nor2b_1 _6793_ (.A(_2740_),
    .B_N(_2741_),
    .Y(_2742_));
 sg13g2_nor2b_1 _6794_ (.A(_2741_),
    .B_N(_0090_),
    .Y(_2743_));
 sg13g2_nor3_1 _6795_ (.A(_0729_),
    .B(_2742_),
    .C(_2743_),
    .Y(_2744_));
 sg13g2_a22oi_1 _6796_ (.Y(_2745_),
    .B1(_2744_),
    .B2(_2737_),
    .A2(_2740_),
    .A1(_2738_));
 sg13g2_inv_2 _6797_ (.Y(_2746_),
    .A(net1113));
 sg13g2_xnor2_1 _6798_ (.Y(_2747_),
    .A(_0059_),
    .B(_0735_));
 sg13g2_nor2b_1 _6799_ (.A(_2747_),
    .B_N(_2741_),
    .Y(_2748_));
 sg13g2_nor2b_1 _6800_ (.A(_2741_),
    .B_N(_0059_),
    .Y(_2749_));
 sg13g2_nor3_1 _6801_ (.A(_0729_),
    .B(_2748_),
    .C(_2749_),
    .Y(_2750_));
 sg13g2_a22oi_1 _6802_ (.Y(_2751_),
    .B1(_2750_),
    .B2(_2737_),
    .A2(_2747_),
    .A1(_2738_));
 sg13g2_inv_4 _6803_ (.A(net1112),
    .Y(_2752_));
 sg13g2_nor2_2 _6804_ (.A(_2746_),
    .B(_2752_),
    .Y(_2753_));
 sg13g2_nand2_1 _6805_ (.Y(_2754_),
    .A(net1116),
    .B(_2751_));
 sg13g2_nor2_2 _6806_ (.A(_2690_),
    .B(net1244),
    .Y(_2755_));
 sg13g2_nor2_1 _6807_ (.A(_3240_),
    .B(net1226),
    .Y(_2756_));
 sg13g2_nand2_1 _6808_ (.Y(_2757_),
    .A(net1118),
    .B(_2756_));
 sg13g2_nand2_1 _6809_ (.Y(_2758_),
    .A(net1110),
    .B(net1173));
 sg13g2_a21oi_1 _6810_ (.A1(net1110),
    .A2(net1173),
    .Y(_2759_),
    .B1(_2755_));
 sg13g2_a21oi_1 _6811_ (.A1(net1160),
    .A2(_2759_),
    .Y(_2760_),
    .B1(net1106));
 sg13g2_nor2_1 _6812_ (.A(net1156),
    .B(_2752_),
    .Y(_2761_));
 sg13g2_nand2_2 _6813_ (.Y(_2762_),
    .A(net1159),
    .B(net1112));
 sg13g2_nor2_2 _6814_ (.A(_2686_),
    .B(net1226),
    .Y(_2763_));
 sg13g2_nor2_1 _6815_ (.A(_2694_),
    .B(_2763_),
    .Y(_2764_));
 sg13g2_nor3_2 _6816_ (.A(net1159),
    .B(net1175),
    .C(_2695_),
    .Y(_2765_));
 sg13g2_nand2_2 _6817_ (.Y(_2766_),
    .A(net1161),
    .B(_2752_));
 sg13g2_nor2_1 _6818_ (.A(net1227),
    .B(net1143),
    .Y(_2767_));
 sg13g2_nor2_1 _6819_ (.A(_2685_),
    .B(_2767_),
    .Y(_2768_));
 sg13g2_nor2b_1 _6820_ (.A(_2766_),
    .B_N(_2768_),
    .Y(_2769_));
 sg13g2_nor2_2 _6821_ (.A(net1156),
    .B(_2685_),
    .Y(_2770_));
 sg13g2_nand2_1 _6822_ (.Y(_2771_),
    .A(net1161),
    .B(net1174));
 sg13g2_nand2_2 _6823_ (.Y(_2772_),
    .A(_2752_),
    .B(_2770_));
 sg13g2_nand2_2 _6824_ (.Y(_2773_),
    .A(net1225),
    .B(net1144));
 sg13g2_a221oi_1 _6825_ (.B2(_2732_),
    .C1(_2765_),
    .B1(_2769_),
    .A1(net1104),
    .Y(_2774_),
    .A2(_2764_));
 sg13g2_nor2_2 _6826_ (.A(_2746_),
    .B(net1112),
    .Y(_2775_));
 sg13g2_nand2_2 _6827_ (.Y(_2776_),
    .A(net1245),
    .B(net1144));
 sg13g2_nand3_1 _6828_ (.B(net1245),
    .C(net1145),
    .A(_2689_),
    .Y(_2777_));
 sg13g2_nand2_2 _6829_ (.Y(_2778_),
    .A(_2757_),
    .B(_2777_));
 sg13g2_a21o_1 _6830_ (.A2(_2778_),
    .A1(net1160),
    .B1(_2765_),
    .X(_2779_));
 sg13g2_a221oi_1 _6831_ (.B2(_2779_),
    .C1(net1419),
    .B1(_2775_),
    .A1(_2736_),
    .Y(_2780_),
    .A2(_2760_));
 sg13g2_o21ai_1 _6832_ (.B1(_2780_),
    .Y(_2781_),
    .A1(net1114),
    .A2(_2774_));
 sg13g2_nand2_2 _6833_ (.Y(_2782_),
    .A(_2687_),
    .B(net1244));
 sg13g2_nand2_1 _6834_ (.Y(_2783_),
    .A(net1225),
    .B(net1117));
 sg13g2_nand3_1 _6835_ (.B(net1118),
    .C(_2783_),
    .A(net1174),
    .Y(_2784_));
 sg13g2_a21oi_1 _6836_ (.A1(_2777_),
    .A2(_2784_),
    .Y(_2785_),
    .B1(net1160));
 sg13g2_nor2_2 _6837_ (.A(net1154),
    .B(net1118),
    .Y(_2786_));
 sg13g2_nand2_2 _6838_ (.Y(_2787_),
    .A(net1227),
    .B(net1243));
 sg13g2_nand2b_2 _6839_ (.Y(_2788_),
    .B(net1143),
    .A_N(_2787_));
 sg13g2_nor2_1 _6840_ (.A(_2685_),
    .B(_2788_),
    .Y(_2789_));
 sg13g2_nand2b_1 _6841_ (.Y(_2790_),
    .B(net1174),
    .A_N(_2788_));
 sg13g2_o21ai_1 _6842_ (.B1(net1104),
    .Y(_2791_),
    .A1(_2786_),
    .A2(_2789_));
 sg13g2_o21ai_1 _6843_ (.B1(_2791_),
    .Y(_2792_),
    .A1(_2772_),
    .A2(_2782_));
 sg13g2_o21ai_1 _6844_ (.B1(_2746_),
    .Y(_2793_),
    .A1(_2785_),
    .A2(_2792_));
 sg13g2_nor2_2 _6845_ (.A(net1154),
    .B(_2727_),
    .Y(_2794_));
 sg13g2_nand2_2 _6846_ (.Y(_2795_),
    .A(net1108),
    .B(net1153));
 sg13g2_nand3_1 _6847_ (.B(net1226),
    .C(_2693_),
    .A(net1175),
    .Y(_2796_));
 sg13g2_o21ai_1 _6848_ (.B1(net1153),
    .Y(_2797_),
    .A1(net1225),
    .A2(net1108));
 sg13g2_nand2b_1 _6849_ (.Y(_2798_),
    .B(_2797_),
    .A_N(_2794_));
 sg13g2_nand2_1 _6850_ (.Y(_2799_),
    .A(_2695_),
    .B(_2768_));
 sg13g2_a21oi_1 _6851_ (.A1(net1244),
    .A2(net1143),
    .Y(_2800_),
    .B1(net1154));
 sg13g2_nor2_1 _6852_ (.A(net1156),
    .B(_2800_),
    .Y(_2801_));
 sg13g2_a21oi_1 _6853_ (.A1(_2799_),
    .A2(_2801_),
    .Y(_2802_),
    .B1(net1106));
 sg13g2_o21ai_1 _6854_ (.B1(_2802_),
    .Y(_2803_),
    .A1(net1159),
    .A2(_2798_));
 sg13g2_nand2_2 _6855_ (.Y(_2804_),
    .A(net1243),
    .B(net1173));
 sg13g2_nor2_1 _6856_ (.A(_3238_),
    .B(_2804_),
    .Y(_2805_));
 sg13g2_o21ai_1 _6857_ (.B1(_2775_),
    .Y(_2806_),
    .A1(_2785_),
    .A2(_2805_));
 sg13g2_nand4_1 _6858_ (.B(_2793_),
    .C(_2803_),
    .A(net1422),
    .Y(_2807_),
    .D(_2806_));
 sg13g2_nand3_1 _6859_ (.B(_2781_),
    .C(_2807_),
    .A(net1416),
    .Y(_2808_));
 sg13g2_nor2_1 _6860_ (.A(net1154),
    .B(net1143),
    .Y(_2809_));
 sg13g2_nor2_2 _6861_ (.A(_2690_),
    .B(_2728_),
    .Y(_2810_));
 sg13g2_nand2_1 _6862_ (.Y(_2811_),
    .A(_2689_),
    .B(_2727_));
 sg13g2_a21oi_1 _6863_ (.A1(_2732_),
    .A2(net1153),
    .Y(_2812_),
    .B1(_2810_));
 sg13g2_nor2_1 _6864_ (.A(_2766_),
    .B(_2812_),
    .Y(_2813_));
 sg13g2_nand2_2 _6865_ (.Y(_2814_),
    .A(net1156),
    .B(net1112));
 sg13g2_nand2_2 _6866_ (.Y(_2815_),
    .A(_2689_),
    .B(net1108));
 sg13g2_a21oi_1 _6867_ (.A1(_2758_),
    .A2(_2815_),
    .Y(_2816_),
    .B1(_2814_));
 sg13g2_o21ai_1 _6868_ (.B1(net1116),
    .Y(_2817_),
    .A1(_2813_),
    .A2(_2816_));
 sg13g2_nor2_1 _6869_ (.A(net1115),
    .B(net1112),
    .Y(_2818_));
 sg13g2_nor2_1 _6870_ (.A(net1244),
    .B(net1143),
    .Y(_2819_));
 sg13g2_nand4_1 _6871_ (.B(_2770_),
    .C(_2782_),
    .A(net1118),
    .Y(_2820_),
    .D(net1105));
 sg13g2_o21ai_1 _6872_ (.B1(net1155),
    .Y(_2821_),
    .A1(_2789_),
    .A2(_2810_));
 sg13g2_or2_1 _6873_ (.X(_2822_),
    .B(_2821_),
    .A(_2753_));
 sg13g2_nor2_1 _6874_ (.A(net1108),
    .B(_2734_),
    .Y(_2823_));
 sg13g2_nand2_2 _6875_ (.Y(_2824_),
    .A(_2730_),
    .B(net1153));
 sg13g2_a21o_1 _6876_ (.A2(_2824_),
    .A1(_2815_),
    .B1(_2762_),
    .X(_2825_));
 sg13g2_nand4_1 _6877_ (.B(_2820_),
    .C(_2822_),
    .A(_2817_),
    .Y(_2826_),
    .D(_2825_));
 sg13g2_nor2b_1 _6878_ (.A(_1971_),
    .B_N(_2826_),
    .Y(_2827_));
 sg13g2_nand2_1 _6879_ (.Y(_2828_),
    .A(net1155),
    .B(_2778_));
 sg13g2_nand3_1 _6880_ (.B(net1117),
    .C(_2778_),
    .A(_2684_),
    .Y(_2829_));
 sg13g2_nor2_1 _6881_ (.A(net1153),
    .B(_2809_),
    .Y(_2830_));
 sg13g2_nor2_1 _6882_ (.A(_2819_),
    .B(_2830_),
    .Y(_2831_));
 sg13g2_nand2_1 _6883_ (.Y(_2832_),
    .A(_2776_),
    .B(_2831_));
 sg13g2_nor2_1 _6884_ (.A(net1154),
    .B(net1108),
    .Y(_2833_));
 sg13g2_nand2_1 _6885_ (.Y(_2834_),
    .A(net1104),
    .B(_2833_));
 sg13g2_nand2_2 _6886_ (.Y(_2835_),
    .A(net1117),
    .B(_2773_));
 sg13g2_nand3_1 _6887_ (.B(net1117),
    .C(_2773_),
    .A(net1174),
    .Y(_2836_));
 sg13g2_o21ai_1 _6888_ (.B1(_2834_),
    .Y(_2837_),
    .A1(_2814_),
    .A2(_2832_));
 sg13g2_o21ai_1 _6889_ (.B1(_2829_),
    .Y(_2838_),
    .A1(net1155),
    .A2(_2836_));
 sg13g2_a22oi_1 _6890_ (.Y(_2839_),
    .B1(_2838_),
    .B2(_2775_),
    .A2(_2837_),
    .A1(net1114));
 sg13g2_or3_1 _6891_ (.A(net1245),
    .B(_2772_),
    .C(_2773_),
    .X(_2840_));
 sg13g2_a21o_1 _6892_ (.A2(_2840_),
    .A1(_2829_),
    .B1(net1113),
    .X(_2841_));
 sg13g2_nand2_1 _6893_ (.Y(_2842_),
    .A(net1243),
    .B(_2767_));
 sg13g2_or2_1 _6894_ (.X(_2843_),
    .B(_2796_),
    .A(net1145));
 sg13g2_nor2_1 _6895_ (.A(_2762_),
    .B(_2843_),
    .Y(_2844_));
 sg13g2_o21ai_1 _6896_ (.B1(_2804_),
    .Y(_2845_),
    .A1(net1115),
    .A2(_2811_));
 sg13g2_a21oi_1 _6897_ (.A1(_2761_),
    .A2(_2845_),
    .Y(_2846_),
    .B1(_2844_));
 sg13g2_nand3_1 _6898_ (.B(_2841_),
    .C(_2846_),
    .A(_2839_),
    .Y(_2847_));
 sg13g2_a21oi_1 _6899_ (.A1(_0557_),
    .A2(_2847_),
    .Y(_2848_),
    .B1(_2827_));
 sg13g2_nand3_1 _6900_ (.B(_2808_),
    .C(_2848_),
    .A(_3133_),
    .Y(_2849_));
 sg13g2_nand3_1 _6901_ (.B(_2770_),
    .C(_2819_),
    .A(net1227),
    .Y(_2850_));
 sg13g2_nor2_2 _6902_ (.A(net1113),
    .B(_2752_),
    .Y(_2851_));
 sg13g2_nor2_1 _6903_ (.A(_2753_),
    .B(net1105),
    .Y(_2852_));
 sg13g2_nand3_1 _6904_ (.B(_2727_),
    .C(net1173),
    .A(net1161),
    .Y(_2853_));
 sg13g2_a22oi_1 _6905_ (.Y(_2854_),
    .B1(_2853_),
    .B2(net1105),
    .A2(_2852_),
    .A1(_2850_));
 sg13g2_nand2_1 _6906_ (.Y(_2855_),
    .A(net1225),
    .B(_2727_));
 sg13g2_nand3_1 _6907_ (.B(net1118),
    .C(_2855_),
    .A(net1175),
    .Y(_2856_));
 sg13g2_nand2b_1 _6908_ (.Y(_2857_),
    .B(_2856_),
    .A_N(_2786_));
 sg13g2_a21oi_1 _6909_ (.A1(net1158),
    .A2(_2857_),
    .Y(_2858_),
    .B1(_2854_));
 sg13g2_nor2_2 _6910_ (.A(net1157),
    .B(_2755_),
    .Y(_2859_));
 sg13g2_nand2_1 _6911_ (.Y(_2860_),
    .A(_2795_),
    .B(_2859_));
 sg13g2_nor2_1 _6912_ (.A(net1110),
    .B(_2763_),
    .Y(_2861_));
 sg13g2_o21ai_1 _6913_ (.B1(net1158),
    .Y(_2862_),
    .A1(net1109),
    .A2(_2763_));
 sg13g2_a21oi_1 _6914_ (.A1(_2860_),
    .A2(_2862_),
    .Y(_2863_),
    .B1(net1107));
 sg13g2_nor3_1 _6915_ (.A(net1420),
    .B(_2858_),
    .C(_2863_),
    .Y(_2864_));
 sg13g2_o21ai_1 _6916_ (.B1(_2852_),
    .Y(_2865_),
    .A1(net1156),
    .A2(_2790_));
 sg13g2_nand2_1 _6917_ (.Y(_2866_),
    .A(net1143),
    .B(_2770_));
 sg13g2_o21ai_1 _6918_ (.B1(net1105),
    .Y(_2867_),
    .A1(_2782_),
    .A2(_2866_));
 sg13g2_a22oi_1 _6919_ (.Y(_2868_),
    .B1(_2865_),
    .B2(_2867_),
    .A2(_2831_),
    .A1(net1156));
 sg13g2_a21oi_1 _6920_ (.A1(net1225),
    .A2(net1108),
    .Y(_2869_),
    .B1(net1174));
 sg13g2_nor2_1 _6921_ (.A(net1161),
    .B(_2869_),
    .Y(_2870_));
 sg13g2_o21ai_1 _6922_ (.B1(net1161),
    .Y(_2871_),
    .A1(_2800_),
    .A2(_2823_));
 sg13g2_a21oi_1 _6923_ (.A1(_2824_),
    .A2(_2870_),
    .Y(_2872_),
    .B1(net1107));
 sg13g2_nand2b_1 _6924_ (.Y(_2873_),
    .B(net1419),
    .A_N(_2868_));
 sg13g2_a21oi_1 _6925_ (.A1(_2871_),
    .A2(_2872_),
    .Y(_2874_),
    .B1(_2873_));
 sg13g2_o21ai_1 _6926_ (.B1(net1416),
    .Y(_2875_),
    .A1(_2864_),
    .A2(_2874_));
 sg13g2_a21oi_1 _6927_ (.A1(_2695_),
    .A2(_2776_),
    .Y(_2876_),
    .B1(_2772_));
 sg13g2_and2_1 _6928_ (.A(net1155),
    .B(net1173),
    .X(_2877_));
 sg13g2_a22oi_1 _6929_ (.Y(_2878_),
    .B1(_2877_),
    .B2(net1144),
    .A2(_2810_),
    .A1(net1155));
 sg13g2_inv_1 _6930_ (.Y(_2879_),
    .A(_2878_));
 sg13g2_nand2_1 _6931_ (.Y(_2880_),
    .A(net1174),
    .B(_2694_));
 sg13g2_o21ai_1 _6932_ (.B1(_2878_),
    .Y(_2881_),
    .A1(net1159),
    .A2(_2880_));
 sg13g2_a21oi_1 _6933_ (.A1(_2773_),
    .A2(_2876_),
    .Y(_2882_),
    .B1(_2881_));
 sg13g2_nor2b_1 _6934_ (.A(_2844_),
    .B_N(_2882_),
    .Y(_2883_));
 sg13g2_nor2_1 _6935_ (.A(net1157),
    .B(_2786_),
    .Y(_2884_));
 sg13g2_a221oi_1 _6936_ (.B2(_2795_),
    .C1(net1107),
    .B1(_2884_),
    .A1(net1157),
    .Y(_2885_),
    .A2(_2812_));
 sg13g2_a21oi_1 _6937_ (.A1(_2788_),
    .A2(_2842_),
    .Y(_2886_),
    .B1(_2771_));
 sg13g2_o21ai_1 _6938_ (.B1(_2775_),
    .Y(_2887_),
    .A1(_2881_),
    .A2(_2886_));
 sg13g2_o21ai_1 _6939_ (.B1(_2887_),
    .Y(_2888_),
    .A1(net1113),
    .A2(_2883_));
 sg13g2_o21ai_1 _6940_ (.B1(_0557_),
    .Y(_2889_),
    .A1(_2885_),
    .A2(_2888_));
 sg13g2_nor4_1 _6941_ (.A(net1161),
    .B(net1153),
    .C(net1112),
    .D(_2869_),
    .Y(_2890_));
 sg13g2_o21ai_1 _6942_ (.B1(net1104),
    .Y(_2891_),
    .A1(_2809_),
    .A2(_2823_));
 sg13g2_nand3_1 _6943_ (.B(_2840_),
    .C(_2891_),
    .A(net1115),
    .Y(_2892_));
 sg13g2_nand2_1 _6944_ (.Y(_2893_),
    .A(_2795_),
    .B(_2815_));
 sg13g2_a21oi_1 _6945_ (.A1(_2797_),
    .A2(_2815_),
    .Y(_2894_),
    .B1(_2814_));
 sg13g2_nor3_1 _6946_ (.A(_2890_),
    .B(_2892_),
    .C(_2894_),
    .Y(_2895_));
 sg13g2_o21ai_1 _6947_ (.B1(net1112),
    .Y(_2896_),
    .A1(net1227),
    .A2(net1244));
 sg13g2_nor2_1 _6948_ (.A(_2694_),
    .B(net1112),
    .Y(_2897_));
 sg13g2_nor2_1 _6949_ (.A(_2866_),
    .B(_2897_),
    .Y(_2898_));
 sg13g2_a221oi_1 _6950_ (.B2(_2898_),
    .C1(net1115),
    .B1(_2896_),
    .A1(_2734_),
    .Y(_2899_),
    .A2(_2870_));
 sg13g2_or3_1 _6951_ (.A(_1971_),
    .B(_2895_),
    .C(_2899_),
    .X(_2900_));
 sg13g2_nand4_1 _6952_ (.B(_2875_),
    .C(_2889_),
    .A(net1415),
    .Y(_2901_),
    .D(_2900_));
 sg13g2_nand3_1 _6953_ (.B(_2849_),
    .C(_2901_),
    .A(\dtop.vtop.logo.addr[11] ),
    .Y(_2902_));
 sg13g2_nand3_1 _6954_ (.B(net1109),
    .C(_2787_),
    .A(_2685_),
    .Y(_2903_));
 sg13g2_a21oi_1 _6955_ (.A1(_2735_),
    .A2(_2903_),
    .Y(_2904_),
    .B1(_2762_));
 sg13g2_a22oi_1 _6956_ (.Y(_2905_),
    .B1(_2763_),
    .B2(net1244),
    .A2(_2733_),
    .A1(net1109));
 sg13g2_nor2_2 _6957_ (.A(_2731_),
    .B(_2771_),
    .Y(_2906_));
 sg13g2_a21oi_1 _6958_ (.A1(_2897_),
    .A2(_2906_),
    .Y(_2907_),
    .B1(net1419));
 sg13g2_o21ai_1 _6959_ (.B1(_2907_),
    .Y(_2908_),
    .A1(_2814_),
    .A2(_2905_));
 sg13g2_nand2_1 _6960_ (.Y(_2909_),
    .A(_2768_),
    .B(_2776_));
 sg13g2_nand2_1 _6961_ (.Y(_2910_),
    .A(net1156),
    .B(_2909_));
 sg13g2_nand2_1 _6962_ (.Y(_2911_),
    .A(_2787_),
    .B(_2869_));
 sg13g2_nand2b_1 _6963_ (.Y(_2912_),
    .B(_2911_),
    .A_N(_2910_));
 sg13g2_a21oi_1 _6964_ (.A1(_2797_),
    .A2(_2859_),
    .Y(_2913_),
    .B1(_2752_));
 sg13g2_or2_1 _6965_ (.X(_2914_),
    .B(_2797_),
    .A(_2767_));
 sg13g2_o21ai_1 _6966_ (.B1(net1419),
    .Y(_2915_),
    .A1(_2766_),
    .A2(_2914_));
 sg13g2_a21oi_1 _6967_ (.A1(_2912_),
    .A2(_2913_),
    .Y(_2916_),
    .B1(_2915_));
 sg13g2_o21ai_1 _6968_ (.B1(net1116),
    .Y(_2917_),
    .A1(_2904_),
    .A2(_2908_));
 sg13g2_nor2_1 _6969_ (.A(_2916_),
    .B(_2917_),
    .Y(_2918_));
 sg13g2_nand3_1 _6970_ (.B(_2763_),
    .C(_2851_),
    .A(net1243),
    .Y(_2919_));
 sg13g2_nand2_1 _6971_ (.Y(_2920_),
    .A(net1421),
    .B(net1158));
 sg13g2_nor3_1 _6972_ (.A(net1145),
    .B(_2919_),
    .C(_2920_),
    .Y(_2921_));
 sg13g2_o21ai_1 _6973_ (.B1(net1416),
    .Y(_2922_),
    .A1(_2918_),
    .A2(_2921_));
 sg13g2_a21oi_1 _6974_ (.A1(net1244),
    .A2(_2763_),
    .Y(_2923_),
    .B1(net1420));
 sg13g2_nand2_1 _6975_ (.Y(_2924_),
    .A(_2914_),
    .B(_2923_));
 sg13g2_nand3_1 _6976_ (.B(_2804_),
    .C(_2911_),
    .A(net1420),
    .Y(_2925_));
 sg13g2_a21oi_1 _6977_ (.A1(_2924_),
    .A2(_2925_),
    .Y(_2926_),
    .B1(net1158));
 sg13g2_or2_1 _6978_ (.X(_2927_),
    .B(net1107),
    .A(net1416));
 sg13g2_nand2_2 _6979_ (.Y(_2928_),
    .A(net1226),
    .B(net1118));
 sg13g2_nor2_2 _6980_ (.A(net1175),
    .B(_2928_),
    .Y(_2929_));
 sg13g2_nor2_1 _6981_ (.A(net1420),
    .B(_2929_),
    .Y(_2930_));
 sg13g2_nand2_1 _6982_ (.Y(_2931_),
    .A(_2685_),
    .B(_2835_));
 sg13g2_and2_1 _6983_ (.A(net1420),
    .B(_2931_),
    .X(_2932_));
 sg13g2_a22oi_1 _6984_ (.Y(_2933_),
    .B1(_2932_),
    .B2(_2824_),
    .A2(_2930_),
    .A1(_2795_));
 sg13g2_nor2_1 _6985_ (.A(_2926_),
    .B(_2927_),
    .Y(_2934_));
 sg13g2_o21ai_1 _6986_ (.B1(_2934_),
    .Y(_2935_),
    .A1(net1162),
    .A2(_2933_));
 sg13g2_nand3_1 _6987_ (.B(_2746_),
    .C(_2928_),
    .A(net1420),
    .Y(_2936_));
 sg13g2_nor2_1 _6988_ (.A(net1421),
    .B(net1158),
    .Y(_2937_));
 sg13g2_nand2_1 _6989_ (.Y(_2938_),
    .A(net1226),
    .B(_2730_));
 sg13g2_nand3_1 _6990_ (.B(_2937_),
    .C(_2938_),
    .A(_2818_),
    .Y(_2939_));
 sg13g2_o21ai_1 _6991_ (.B1(_2939_),
    .Y(_2940_),
    .A1(_2766_),
    .A2(_2936_));
 sg13g2_nand3_1 _6992_ (.B(_2787_),
    .C(_2940_),
    .A(net1175),
    .Y(_2941_));
 sg13g2_nand4_1 _6993_ (.B(_2922_),
    .C(_2935_),
    .A(net1415),
    .Y(_2942_),
    .D(_2941_));
 sg13g2_nand3_1 _6994_ (.B(_2735_),
    .C(_2931_),
    .A(net1162),
    .Y(_2943_));
 sg13g2_nor2_2 _6995_ (.A(_2731_),
    .B(_2799_),
    .Y(_2944_));
 sg13g2_or3_1 _6996_ (.A(_2683_),
    .B(_2810_),
    .C(_2944_),
    .X(_2945_));
 sg13g2_nand3_1 _6997_ (.B(_2943_),
    .C(_2945_),
    .A(_2753_),
    .Y(_2946_));
 sg13g2_nand3_1 _6998_ (.B(_2906_),
    .C(_2928_),
    .A(net1105),
    .Y(_2947_));
 sg13g2_nand3_1 _6999_ (.B(_2946_),
    .C(_2947_),
    .A(net1420),
    .Y(_2948_));
 sg13g2_nand2_1 _7000_ (.Y(_2949_),
    .A(net1153),
    .B(_2788_));
 sg13g2_a21oi_1 _7001_ (.A1(net1153),
    .A2(_2788_),
    .Y(_2950_),
    .B1(net1160));
 sg13g2_nor2_1 _7002_ (.A(net1158),
    .B(_2929_),
    .Y(_2951_));
 sg13g2_a221oi_1 _7003_ (.B2(_2795_),
    .C1(net1107),
    .B1(_2951_),
    .A1(net1157),
    .Y(_2952_),
    .A2(_2949_));
 sg13g2_nor3_1 _7004_ (.A(net1116),
    .B(_2772_),
    .C(_2928_),
    .Y(_2953_));
 sg13g2_nor3_1 _7005_ (.A(net1421),
    .B(_2952_),
    .C(_2953_),
    .Y(_2954_));
 sg13g2_nor2b_1 _7006_ (.A(_2954_),
    .B_N(net1416),
    .Y(_2955_));
 sg13g2_o21ai_1 _7007_ (.B1(net1160),
    .Y(_2956_),
    .A1(_2810_),
    .A2(_2944_));
 sg13g2_or3_1 _7008_ (.A(net1161),
    .B(_2731_),
    .C(_2734_),
    .X(_2957_));
 sg13g2_nand3_1 _7009_ (.B(_2956_),
    .C(_2957_),
    .A(net1419),
    .Y(_2958_));
 sg13g2_nor2_1 _7010_ (.A(net1421),
    .B(net1162),
    .Y(_2959_));
 sg13g2_nand2b_1 _7011_ (.Y(_2960_),
    .B(net1157),
    .A_N(net1422));
 sg13g2_a221oi_1 _7012_ (.B2(_2843_),
    .C1(_2927_),
    .B1(_2959_),
    .A1(_2937_),
    .Y(_2961_),
    .A2(_2949_));
 sg13g2_a22oi_1 _7013_ (.Y(_2962_),
    .B1(_2958_),
    .B2(_2961_),
    .A2(_2955_),
    .A1(_2948_));
 sg13g2_a21oi_1 _7014_ (.A1(_3133_),
    .A2(_2962_),
    .Y(_2963_),
    .B1(\dtop.vtop.logo.addr[11] ));
 sg13g2_nand3_1 _7015_ (.B(net1154),
    .C(_2735_),
    .A(net1160),
    .Y(_2964_));
 sg13g2_a21oi_1 _7016_ (.A1(_2815_),
    .A2(_2950_),
    .Y(_2965_),
    .B1(net1106));
 sg13g2_and2_1 _7017_ (.A(_2770_),
    .B(_2787_),
    .X(_2966_));
 sg13g2_nor3_1 _7018_ (.A(net1159),
    .B(net1174),
    .C(_2788_),
    .Y(_2967_));
 sg13g2_a21o_1 _7019_ (.A2(_2966_),
    .A1(_2776_),
    .B1(_2967_),
    .X(_2968_));
 sg13g2_nand3_1 _7020_ (.B(net1105),
    .C(_2966_),
    .A(net1110),
    .Y(_2969_));
 sg13g2_o21ai_1 _7021_ (.B1(_2969_),
    .Y(_2970_),
    .A1(net1113),
    .A2(_2878_));
 sg13g2_a21oi_1 _7022_ (.A1(_2851_),
    .A2(_2968_),
    .Y(_2971_),
    .B1(_2970_));
 sg13g2_o21ai_1 _7023_ (.B1(_2878_),
    .Y(_2972_),
    .A1(net1155),
    .A2(_2797_));
 sg13g2_a22oi_1 _7024_ (.Y(_2973_),
    .B1(_2972_),
    .B2(_2775_),
    .A2(_2965_),
    .A1(_2964_));
 sg13g2_a21oi_1 _7025_ (.A1(_2971_),
    .A2(_2973_),
    .Y(_2974_),
    .B1(net1419));
 sg13g2_nor2_1 _7026_ (.A(net1108),
    .B(_2896_),
    .Y(_2975_));
 sg13g2_a21oi_1 _7027_ (.A1(_2776_),
    .A2(_2835_),
    .Y(_2976_),
    .B1(_2751_));
 sg13g2_nor3_1 _7028_ (.A(_2771_),
    .B(_2975_),
    .C(_2976_),
    .Y(_2977_));
 sg13g2_nor3_1 _7029_ (.A(net1154),
    .B(_2726_),
    .C(_2814_),
    .Y(_2978_));
 sg13g2_nor2_1 _7030_ (.A(_2766_),
    .B(_2909_),
    .Y(_2979_));
 sg13g2_nor2_1 _7031_ (.A(_2746_),
    .B(_2978_),
    .Y(_2980_));
 sg13g2_a221oi_1 _7032_ (.B2(net1104),
    .C1(_2979_),
    .B1(_2798_),
    .A1(_2752_),
    .Y(_2981_),
    .A2(_2765_));
 sg13g2_or2_1 _7033_ (.X(_2982_),
    .B(_2765_),
    .A(net1113));
 sg13g2_o21ai_1 _7034_ (.B1(net1422),
    .Y(_2983_),
    .A1(_2977_),
    .A2(_2982_));
 sg13g2_a21oi_1 _7035_ (.A1(_2980_),
    .A2(_2981_),
    .Y(_2984_),
    .B1(_2983_));
 sg13g2_o21ai_1 _7036_ (.B1(net1416),
    .Y(_2985_),
    .A1(_2974_),
    .A2(_2984_));
 sg13g2_a21oi_1 _7037_ (.A1(_2836_),
    .A2(_2903_),
    .Y(_2986_),
    .B1(_2814_));
 sg13g2_a21oi_1 _7038_ (.A1(net1227),
    .A2(_2819_),
    .Y(_2987_),
    .B1(_2734_));
 sg13g2_o21ai_1 _7039_ (.B1(net1104),
    .Y(_2988_),
    .A1(_2833_),
    .A2(_2987_));
 sg13g2_o21ai_1 _7040_ (.B1(_2988_),
    .Y(_2989_),
    .A1(_2766_),
    .A2(_2804_));
 sg13g2_o21ai_1 _7041_ (.B1(net1116),
    .Y(_2990_),
    .A1(_2986_),
    .A2(_2989_));
 sg13g2_o21ai_1 _7042_ (.B1(_2990_),
    .Y(_2991_),
    .A1(net1162),
    .A2(_2919_));
 sg13g2_or2_1 _7043_ (.X(_2992_),
    .B(_2991_),
    .A(_2953_));
 sg13g2_nor2b_1 _7044_ (.A(_2735_),
    .B_N(_2775_),
    .Y(_2993_));
 sg13g2_nand3_1 _7045_ (.B(_2818_),
    .C(_2835_),
    .A(net1175),
    .Y(_2994_));
 sg13g2_a21oi_1 _7046_ (.A1(_2758_),
    .A2(_2815_),
    .Y(_2995_),
    .B1(net1107));
 sg13g2_nor3_1 _7047_ (.A(net1157),
    .B(_2993_),
    .C(_2995_),
    .Y(_2996_));
 sg13g2_nand2b_1 _7048_ (.Y(_2997_),
    .B(net1106),
    .A_N(_2757_));
 sg13g2_nand3_1 _7049_ (.B(_2861_),
    .C(_2880_),
    .A(_2753_),
    .Y(_2998_));
 sg13g2_nand4_1 _7050_ (.B(_2919_),
    .C(_2997_),
    .A(net1157),
    .Y(_2999_),
    .D(_2998_));
 sg13g2_a21oi_1 _7051_ (.A1(_2994_),
    .A2(_2996_),
    .Y(_3000_),
    .B1(_1971_));
 sg13g2_a221oi_1 _7052_ (.B2(_3000_),
    .C1(net1415),
    .B1(_2999_),
    .A1(_0557_),
    .Y(_3001_),
    .A2(_2992_));
 sg13g2_a21oi_1 _7053_ (.A1(_2815_),
    .A2(_2914_),
    .Y(_3002_),
    .B1(_2762_));
 sg13g2_nor2b_1 _7054_ (.A(_2814_),
    .B_N(_2798_),
    .Y(_3003_));
 sg13g2_or3_1 _7055_ (.A(_2979_),
    .B(_3002_),
    .C(_3003_),
    .X(_3004_));
 sg13g2_nand3_1 _7056_ (.B(net1117),
    .C(net1173),
    .A(net1159),
    .Y(_3005_));
 sg13g2_nand4_1 _7057_ (.B(net1117),
    .C(net1173),
    .A(net1159),
    .Y(_3006_),
    .D(_2851_));
 sg13g2_nand4_1 _7058_ (.B(_2822_),
    .C(_2969_),
    .A(net1419),
    .Y(_3007_),
    .D(_3006_));
 sg13g2_a21oi_1 _7059_ (.A1(net1113),
    .A2(_3004_),
    .Y(_3008_),
    .B1(_3007_));
 sg13g2_nand3_1 _7060_ (.B(net1110),
    .C(_2735_),
    .A(net1160),
    .Y(_3009_));
 sg13g2_a21oi_1 _7061_ (.A1(net1154),
    .A2(_2735_),
    .Y(_3010_),
    .B1(net1106));
 sg13g2_nand2_1 _7062_ (.Y(_3011_),
    .A(net1104),
    .B(_2944_));
 sg13g2_a21oi_1 _7063_ (.A1(_2829_),
    .A2(_3011_),
    .Y(_3012_),
    .B1(net1113));
 sg13g2_and3_1 _7064_ (.X(_3013_),
    .A(_2783_),
    .B(net1105),
    .C(_2966_));
 sg13g2_nor3_1 _7065_ (.A(net1422),
    .B(_3012_),
    .C(_3013_),
    .Y(_3014_));
 sg13g2_o21ai_1 _7066_ (.B1(_2829_),
    .Y(_3015_),
    .A1(net1155),
    .A2(_2797_));
 sg13g2_a22oi_1 _7067_ (.Y(_3016_),
    .B1(_3015_),
    .B2(_2775_),
    .A2(_3010_),
    .A1(_3009_));
 sg13g2_a21oi_1 _7068_ (.A1(_3014_),
    .A2(_3016_),
    .Y(_3017_),
    .B1(_3008_));
 sg13g2_a22oi_1 _7069_ (.Y(_3018_),
    .B1(_2897_),
    .B2(_2906_),
    .A2(_2893_),
    .A1(net1104));
 sg13g2_o21ai_1 _7070_ (.B1(_3018_),
    .Y(_3019_),
    .A1(_2759_),
    .A2(_2814_));
 sg13g2_a21oi_1 _7071_ (.A1(net1244),
    .A2(_2877_),
    .Y(_3020_),
    .B1(_2879_));
 sg13g2_o21ai_1 _7072_ (.B1(_3020_),
    .Y(_3021_),
    .A1(_2762_),
    .A2(_2836_));
 sg13g2_and3_1 _7073_ (.X(_3022_),
    .A(net1105),
    .B(_2855_),
    .C(_2906_));
 sg13g2_a221oi_1 _7074_ (.B2(net1106),
    .C1(_3022_),
    .B1(_3021_),
    .A1(net1114),
    .Y(_3023_),
    .A2(_3019_));
 sg13g2_nor2_1 _7075_ (.A(_1971_),
    .B(_3023_),
    .Y(_3024_));
 sg13g2_o21ai_1 _7076_ (.B1(_2828_),
    .Y(_3025_),
    .A1(_2762_),
    .A2(_2909_));
 sg13g2_o21ai_1 _7077_ (.B1(_2746_),
    .Y(_3026_),
    .A1(_2876_),
    .A2(_3025_));
 sg13g2_nand2_1 _7078_ (.Y(_3027_),
    .A(_2828_),
    .B(_3005_));
 sg13g2_nor2_1 _7079_ (.A(net1162),
    .B(_2929_),
    .Y(_3028_));
 sg13g2_a221oi_1 _7080_ (.B2(_2799_),
    .C1(net1106),
    .B1(_3028_),
    .A1(net1159),
    .Y(_3029_),
    .A2(_2832_));
 sg13g2_a21oi_1 _7081_ (.A1(_2775_),
    .A2(_3027_),
    .Y(_3030_),
    .B1(_3029_));
 sg13g2_nand2_1 _7082_ (.Y(_3031_),
    .A(_3026_),
    .B(_3030_));
 sg13g2_a221oi_1 _7083_ (.B2(_0557_),
    .C1(_3024_),
    .B1(_3031_),
    .A1(net1416),
    .Y(_3032_),
    .A2(_3017_));
 sg13g2_a22oi_1 _7084_ (.Y(_3033_),
    .B1(_3032_),
    .B2(net1415),
    .A2(_3001_),
    .A1(_2985_));
 sg13g2_or2_1 _7085_ (.X(_3034_),
    .B(_3033_),
    .A(\dtop.vtop.logo.addr[11] ));
 sg13g2_nor3_1 _7086_ (.A(net1106),
    .B(_2833_),
    .C(_2910_),
    .Y(_3035_));
 sg13g2_a21oi_1 _7087_ (.A1(_2859_),
    .A2(_2949_),
    .Y(_3036_),
    .B1(_3035_));
 sg13g2_o21ai_1 _7088_ (.B1(net1107),
    .Y(_3037_),
    .A1(_2777_),
    .A2(_2960_));
 sg13g2_a21oi_1 _7089_ (.A1(net1117),
    .A2(net1173),
    .Y(_3038_),
    .B1(net1162));
 sg13g2_a21oi_1 _7090_ (.A1(_2815_),
    .A2(_3038_),
    .Y(_3039_),
    .B1(_2884_));
 sg13g2_nor2b_1 _7091_ (.A(_3039_),
    .B_N(net1421),
    .Y(_3040_));
 sg13g2_o21ai_1 _7092_ (.B1(_3037_),
    .Y(_3041_),
    .A1(net1421),
    .A2(_3036_));
 sg13g2_o21ai_1 _7093_ (.B1(net1416),
    .Y(_3042_),
    .A1(_3040_),
    .A2(_3041_));
 sg13g2_nand3_1 _7094_ (.B(_2782_),
    .C(_2870_),
    .A(net1108),
    .Y(_3043_));
 sg13g2_nand3_1 _7095_ (.B(_2871_),
    .C(_3043_),
    .A(net1420),
    .Y(_3044_));
 sg13g2_nor2b_1 _7096_ (.A(_2794_),
    .B_N(_2937_),
    .Y(_3045_));
 sg13g2_a221oi_1 _7097_ (.B2(net1175),
    .C1(_2960_),
    .B1(_2732_),
    .A1(_2689_),
    .Y(_3046_),
    .A2(_2730_));
 sg13g2_a21oi_1 _7098_ (.A1(_2795_),
    .A2(_3045_),
    .Y(_3047_),
    .B1(_3046_));
 sg13g2_a21oi_1 _7099_ (.A1(_3044_),
    .A2(_3047_),
    .Y(_3048_),
    .B1(_2927_));
 sg13g2_a22oi_1 _7100_ (.Y(_3049_),
    .B1(_2829_),
    .B2(_0557_),
    .A2(_2821_),
    .A1(net1419));
 sg13g2_o21ai_1 _7101_ (.B1(_3133_),
    .Y(_3050_),
    .A1(_2753_),
    .A2(_3049_));
 sg13g2_nor2_1 _7102_ (.A(_3048_),
    .B(_3050_),
    .Y(_3051_));
 sg13g2_nand2_1 _7103_ (.Y(_3052_),
    .A(_3042_),
    .B(_3051_));
 sg13g2_and3_1 _7104_ (.X(_3053_),
    .A(net1422),
    .B(_2796_),
    .C(_2884_));
 sg13g2_nor4_1 _7105_ (.A(net1421),
    .B(net1157),
    .C(_2733_),
    .D(_2929_),
    .Y(_3054_));
 sg13g2_o21ai_1 _7106_ (.B1(net1415),
    .Y(_3055_),
    .A1(_2755_),
    .A2(_2960_));
 sg13g2_o21ai_1 _7107_ (.B1(_2753_),
    .Y(_3056_),
    .A1(_2794_),
    .A2(_2920_));
 sg13g2_or4_1 _7108_ (.A(_3053_),
    .B(_3054_),
    .C(_3055_),
    .D(_3056_),
    .X(_3057_));
 sg13g2_nand3_1 _7109_ (.B(_3052_),
    .C(_3057_),
    .A(\dtop.vtop.logo.addr[11] ),
    .Y(_3058_));
 sg13g2_a21oi_1 _7110_ (.A1(_3034_),
    .A2(_3058_),
    .Y(_3059_),
    .B1(_3132_));
 sg13g2_a21oi_1 _7111_ (.A1(_2942_),
    .A2(_2963_),
    .Y(_3060_),
    .B1(\dtop.vtop.logo.addr[10] ));
 sg13g2_a21o_1 _7112_ (.A2(_3060_),
    .A1(_2902_),
    .B1(_3059_),
    .X(_3061_));
 sg13g2_nor4_1 _7113_ (.A(_2675_),
    .B(_2681_),
    .C(_2682_),
    .D(_3061_),
    .Y(_3062_));
 sg13g2_mux2_1 _7114_ (.A0(net462),
    .A1(_3062_),
    .S(net1361),
    .X(_0395_));
 sg13g2_mux2_1 _7115_ (.A0(_3062_),
    .A1(net558),
    .S(net1361),
    .X(_0396_));
 sg13g2_dfrbp_1 _7116_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net12),
    .D(net2),
    .Q_N(_3551_),
    .Q(\dtop.ext_control[0] ));
 sg13g2_dfrbp_1 _7117_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net13),
    .D(net3),
    .Q_N(_3552_),
    .Q(\dtop.ext_control[1] ));
 sg13g2_dfrbp_1 _7118_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net14),
    .D(net4),
    .Q_N(_3553_),
    .Q(\dtop.ext_control[2] ));
 sg13g2_dfrbp_1 _7119_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net15),
    .D(net5),
    .Q_N(_0079_),
    .Q(\dtop.ext_control[3] ));
 sg13g2_dfrbp_1 _7120_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net16),
    .D(net6),
    .Q_N(_0006_),
    .Q(\dtop.ext_control[4] ));
 sg13g2_dfrbp_1 _7121_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net17),
    .D(net7),
    .Q_N(_3554_),
    .Q(\dtop.ext_control[5] ));
 sg13g2_dfrbp_1 _7122_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net35),
    .D(net8),
    .Q_N(_3555_),
    .Q(\dtop.ext_control[6] ));
 sg13g2_dfrbp_1 _7123_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net11),
    .D(net9),
    .Q_N(_0078_),
    .Q(advance_frame));
 sg13g2_dfrbp_1 _7124_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net258),
    .D(_0100_),
    .Q_N(_0085_),
    .Q(\dtop.oct_counter[0] ));
 sg13g2_dfrbp_1 _7125_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net257),
    .D(net671),
    .Q_N(_0084_),
    .Q(\dtop.oct_counter[1] ));
 sg13g2_dfrbp_1 _7126_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net256),
    .D(net575),
    .Q_N(_0083_),
    .Q(\dtop.oct_counter[2] ));
 sg13g2_dfrbp_1 _7127_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net255),
    .D(net470),
    .Q_N(_3550_),
    .Q(uio_out[0]));
 sg13g2_dfrbp_1 _7128_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net253),
    .D(_0104_),
    .Q_N(_3549_),
    .Q(uio_out[1]));
 sg13g2_dfrbp_1 _7129_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net251),
    .D(_0105_),
    .Q_N(_3548_),
    .Q(uio_out[2]));
 sg13g2_dfrbp_1 _7130_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net249),
    .D(_0106_),
    .Q_N(_3547_),
    .Q(uio_out[3]));
 sg13g2_dfrbp_1 _7131_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net247),
    .D(net565),
    .Q_N(_3546_),
    .Q(uio_out[4]));
 sg13g2_dfrbp_1 _7132_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net245),
    .D(net526),
    .Q_N(_3545_),
    .Q(uio_out[5]));
 sg13g2_dfrbp_1 _7133_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net243),
    .D(_0109_),
    .Q_N(_3544_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _7134_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net242),
    .D(net607),
    .Q_N(_3543_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _7135_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net241),
    .D(net592),
    .Q_N(_3542_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _7136_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net240),
    .D(_0112_),
    .Q_N(_3541_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _7137_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net239),
    .D(_0113_),
    .Q_N(_3540_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _7138_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net238),
    .D(_0114_),
    .Q_N(_3539_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _7139_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net237),
    .D(_0115_),
    .Q_N(_3538_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _7140_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net267),
    .D(net536),
    .Q_N(_3556_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _7141_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net236),
    .D(net1),
    .Q_N(_0087_),
    .Q(rst_n_reg));
 sg13g2_dfrbp_1 _7142_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net235),
    .D(_0117_),
    .Q_N(_3537_),
    .Q(uio_out[6]));
 sg13g2_dfrbp_1 _7143_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net234),
    .D(net582),
    .Q_N(_3536_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _7144_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net233),
    .D(_0119_),
    .Q_N(_0082_),
    .Q(\dtop.oct_counter[3] ));
 sg13g2_dfrbp_1 _7145_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net232),
    .D(_0120_),
    .Q_N(_0081_),
    .Q(\dtop.oct_counter[4] ));
 sg13g2_dfrbp_1 _7146_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net231),
    .D(_0121_),
    .Q_N(_0046_),
    .Q(\dtop.oct_counter[5] ));
 sg13g2_dfrbp_1 _7147_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net230),
    .D(_0122_),
    .Q_N(_3535_),
    .Q(\dtop.oct_counter[6] ));
 sg13g2_dfrbp_1 _7148_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net229),
    .D(_0123_),
    .Q_N(_0051_),
    .Q(\dtop.vtop.logo.addr[7] ));
 sg13g2_dfrbp_1 _7149_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net228),
    .D(_0124_),
    .Q_N(_3534_),
    .Q(\dtop.vtop.logo.addr[8] ));
 sg13g2_dfrbp_1 _7150_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net227),
    .D(_0125_),
    .Q_N(_0055_),
    .Q(\dtop.vtop.logo.addr[9] ));
 sg13g2_dfrbp_1 _7151_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net226),
    .D(_0126_),
    .Q_N(_0064_),
    .Q(\dtop.vtop.logo.addr[10] ));
 sg13g2_dfrbp_1 _7152_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net225),
    .D(_0127_),
    .Q_N(_0080_),
    .Q(\dtop.vtop.logo.addr[11] ));
 sg13g2_dfrbp_1 _7153_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net224),
    .D(net472),
    .Q_N(_3533_),
    .Q(\dtop.player_inst.synth.alu.registers[4][0] ));
 sg13g2_dfrbp_1 _7154_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net222),
    .D(net515),
    .Q_N(_3532_),
    .Q(\dtop.player_inst.synth.alu.registers[4][1] ));
 sg13g2_dfrbp_1 _7155_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net220),
    .D(net500),
    .Q_N(_3531_),
    .Q(\dtop.player_inst.synth.alu.registers[4][2] ));
 sg13g2_dfrbp_1 _7156_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net218),
    .D(net532),
    .Q_N(_3530_),
    .Q(\dtop.player_inst.synth.alu.registers[4][3] ));
 sg13g2_dfrbp_1 _7157_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net216),
    .D(net464),
    .Q_N(_3529_),
    .Q(\dtop.player_inst.synth.alu.registers[4][4] ));
 sg13g2_dfrbp_1 _7158_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net214),
    .D(_0133_),
    .Q_N(_3528_),
    .Q(\dtop.player_inst.synth.alu.registers[4][5] ));
 sg13g2_dfrbp_1 _7159_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net212),
    .D(net330),
    .Q_N(_0067_),
    .Q(\dtop.player_inst.synth.alu.registers[4][6] ));
 sg13g2_dfrbp_1 _7160_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net210),
    .D(net343),
    .Q_N(_0068_),
    .Q(\dtop.player_inst.synth.alu.registers[4][7] ));
 sg13g2_dfrbp_1 _7161_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net208),
    .D(net335),
    .Q_N(_0069_),
    .Q(\dtop.player_inst.synth.alu.registers[4][8] ));
 sg13g2_dfrbp_1 _7162_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net206),
    .D(net339),
    .Q_N(_0070_),
    .Q(\dtop.player_inst.synth.alu.registers[4][9] ));
 sg13g2_dfrbp_1 _7163_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net204),
    .D(net324),
    .Q_N(_0071_),
    .Q(\dtop.player_inst.synth.alu.registers[4][10] ));
 sg13g2_dfrbp_1 _7164_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net202),
    .D(net397),
    .Q_N(_3527_),
    .Q(\dtop.player_inst.synth.alu.registers[2][0] ));
 sg13g2_dfrbp_1 _7165_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net200),
    .D(net387),
    .Q_N(_3526_),
    .Q(\dtop.player_inst.synth.alu.registers[2][1] ));
 sg13g2_dfrbp_1 _7166_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net198),
    .D(net415),
    .Q_N(_3525_),
    .Q(\dtop.player_inst.synth.alu.registers[2][2] ));
 sg13g2_dfrbp_1 _7167_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net196),
    .D(_0142_),
    .Q_N(_3524_),
    .Q(\dtop.player_inst.synth.alu.registers[2][3] ));
 sg13g2_dfrbp_1 _7168_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net194),
    .D(net355),
    .Q_N(_3523_),
    .Q(\dtop.player_inst.synth.alu.registers[2][4] ));
 sg13g2_dfrbp_1 _7169_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net192),
    .D(_0144_),
    .Q_N(_3522_),
    .Q(\dtop.player_inst.synth.alu.registers[2][5] ));
 sg13g2_dfrbp_1 _7170_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net190),
    .D(_0145_),
    .Q_N(_3521_),
    .Q(\dtop.player_inst.synth.alu.registers[2][6] ));
 sg13g2_dfrbp_1 _7171_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net188),
    .D(net350),
    .Q_N(_3520_),
    .Q(\dtop.player_inst.synth.alu.registers[2][7] ));
 sg13g2_dfrbp_1 _7172_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net186),
    .D(_0147_),
    .Q_N(_3519_),
    .Q(\dtop.player_inst.synth.alu.registers[1][0] ));
 sg13g2_dfrbp_1 _7173_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net184),
    .D(net409),
    .Q_N(_3518_),
    .Q(\dtop.player_inst.synth.alu.registers[1][1] ));
 sg13g2_dfrbp_1 _7174_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net182),
    .D(net421),
    .Q_N(_3517_),
    .Q(\dtop.player_inst.synth.alu.registers[1][2] ));
 sg13g2_dfrbp_1 _7175_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net180),
    .D(_0150_),
    .Q_N(_3516_),
    .Q(\dtop.player_inst.synth.alu.registers[1][3] ));
 sg13g2_dfrbp_1 _7176_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net178),
    .D(net407),
    .Q_N(_3515_),
    .Q(\dtop.player_inst.synth.alu.registers[1][4] ));
 sg13g2_dfrbp_1 _7177_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net176),
    .D(_0152_),
    .Q_N(_3514_),
    .Q(\dtop.player_inst.synth.alu.registers[1][5] ));
 sg13g2_dfrbp_1 _7178_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net174),
    .D(net381),
    .Q_N(_3513_),
    .Q(\dtop.player_inst.synth.alu.registers[1][6] ));
 sg13g2_dfrbp_1 _7179_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net172),
    .D(net445),
    .Q_N(_3512_),
    .Q(\dtop.player_inst.synth.alu.registers[1][7] ));
 sg13g2_dfrbp_1 _7180_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net170),
    .D(net435),
    .Q_N(_3511_),
    .Q(\dtop.player_inst.synth.alu.registers[1][8] ));
 sg13g2_dfrbp_1 _7181_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net168),
    .D(net481),
    .Q_N(_3510_),
    .Q(\dtop.player_inst.synth.alu.registers[1][9] ));
 sg13g2_dfrbp_1 _7182_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net166),
    .D(net443),
    .Q_N(_3509_),
    .Q(\dtop.player_inst.synth.alu.registers[1][10] ));
 sg13g2_dfrbp_1 _7183_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net164),
    .D(net547),
    .Q_N(_3508_),
    .Q(\dtop.player_inst.synth.alu.registers[0][0] ));
 sg13g2_dfrbp_1 _7184_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net162),
    .D(net543),
    .Q_N(_3507_),
    .Q(\dtop.player_inst.synth.alu.registers[0][1] ));
 sg13g2_dfrbp_1 _7185_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net160),
    .D(_0160_),
    .Q_N(_3506_),
    .Q(\dtop.player_inst.synth.alu.registers[0][2] ));
 sg13g2_dfrbp_1 _7186_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net158),
    .D(_0161_),
    .Q_N(_3505_),
    .Q(\dtop.player_inst.synth.alu.registers[0][3] ));
 sg13g2_dfrbp_1 _7187_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net156),
    .D(net589),
    .Q_N(_3504_),
    .Q(\dtop.player_inst.synth.alu.registers[0][4] ));
 sg13g2_dfrbp_1 _7188_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net154),
    .D(_0163_),
    .Q_N(_3503_),
    .Q(\dtop.player_inst.synth.alu.registers[0][5] ));
 sg13g2_dfrbp_1 _7189_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net152),
    .D(net550),
    .Q_N(_3502_),
    .Q(\dtop.player_inst.synth.alu.registers[0][6] ));
 sg13g2_dfrbp_1 _7190_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net150),
    .D(net561),
    .Q_N(_3501_),
    .Q(\dtop.player_inst.synth.alu.registers[0][7] ));
 sg13g2_dfrbp_1 _7191_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net148),
    .D(net541),
    .Q_N(_3500_),
    .Q(\dtop.player_inst.synth.alu.registers[0][8] ));
 sg13g2_dfrbp_1 _7192_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net146),
    .D(net587),
    .Q_N(_3499_),
    .Q(\dtop.player_inst.synth.alu.registers[0][9] ));
 sg13g2_dfrbp_1 _7193_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net144),
    .D(_0168_),
    .Q_N(_3498_),
    .Q(\dtop.player_inst.synth.alu.registers[0][10] ));
 sg13g2_dfrbp_1 _7194_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net142),
    .D(net441),
    .Q_N(_3497_),
    .Q(\dtop.out_sample[0] ));
 sg13g2_dfrbp_1 _7195_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net140),
    .D(net519),
    .Q_N(_3496_),
    .Q(\dtop.out_sample[1] ));
 sg13g2_dfrbp_1 _7196_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net138),
    .D(_0171_),
    .Q_N(_3495_),
    .Q(\dtop.out_sample[2] ));
 sg13g2_dfrbp_1 _7197_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net136),
    .D(_0172_),
    .Q_N(_3494_),
    .Q(\dtop.out_sample[3] ));
 sg13g2_dfrbp_1 _7198_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net134),
    .D(_0173_),
    .Q_N(_3493_),
    .Q(\dtop.out_sample[4] ));
 sg13g2_dfrbp_1 _7199_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net132),
    .D(_0174_),
    .Q_N(_3492_),
    .Q(\dtop.out_sample[5] ));
 sg13g2_dfrbp_1 _7200_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net130),
    .D(_0175_),
    .Q_N(_3491_),
    .Q(\dtop.out_sample[6] ));
 sg13g2_dfrbp_1 _7201_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net128),
    .D(_0176_),
    .Q_N(_3490_),
    .Q(\dtop.player_inst.synth.alu.acc[0] ));
 sg13g2_dfrbp_1 _7202_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net126),
    .D(_0177_),
    .Q_N(_3489_),
    .Q(\dtop.player_inst.synth.alu.acc[1] ));
 sg13g2_dfrbp_1 _7203_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net124),
    .D(_0178_),
    .Q_N(_3488_),
    .Q(\dtop.player_inst.synth.alu.acc[2] ));
 sg13g2_dfrbp_1 _7204_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net122),
    .D(_0179_),
    .Q_N(_3487_),
    .Q(\dtop.player_inst.synth.alu.acc[3] ));
 sg13g2_dfrbp_1 _7205_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net120),
    .D(_0180_),
    .Q_N(_3486_),
    .Q(\dtop.player_inst.synth.alu.acc[4] ));
 sg13g2_dfrbp_1 _7206_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net118),
    .D(_0181_),
    .Q_N(_3485_),
    .Q(\dtop.player_inst.synth.alu.acc[5] ));
 sg13g2_dfrbp_1 _7207_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net116),
    .D(_0182_),
    .Q_N(_3484_),
    .Q(\dtop.player_inst.synth.alu.acc[6] ));
 sg13g2_dfrbp_1 _7208_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net114),
    .D(_0183_),
    .Q_N(_3483_),
    .Q(\dtop.player_inst.synth.alu.acc[7] ));
 sg13g2_dfrbp_1 _7209_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net112),
    .D(_0184_),
    .Q_N(_3482_),
    .Q(\dtop.player_inst.synth.alu.acc[8] ));
 sg13g2_dfrbp_1 _7210_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net110),
    .D(_0185_),
    .Q_N(_3481_),
    .Q(\dtop.player_inst.synth.alu.acc[9] ));
 sg13g2_dfrbp_1 _7211_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net108),
    .D(_0186_),
    .Q_N(_0063_),
    .Q(\dtop.player_inst.synth.alu.acc[10] ));
 sg13g2_dfrbp_1 _7212_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net106),
    .D(_0187_),
    .Q_N(_3480_),
    .Q(\dtop.player_inst.synth.alu.carry ));
 sg13g2_dfrbp_1 _7213_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net104),
    .D(net369),
    .Q_N(_3479_),
    .Q(\dtop.player_inst.synth.alu.registers[5][0] ));
 sg13g2_dfrbp_1 _7214_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net102),
    .D(_0189_),
    .Q_N(_3478_),
    .Q(\dtop.player_inst.synth.alu.registers[5][1] ));
 sg13g2_dfrbp_1 _7215_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net100),
    .D(net438),
    .Q_N(_3477_),
    .Q(\dtop.player_inst.synth.alu.registers[5][2] ));
 sg13g2_dfrbp_1 _7216_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net98),
    .D(net405),
    .Q_N(_3476_),
    .Q(\dtop.player_inst.synth.alu.registers[5][3] ));
 sg13g2_dfrbp_1 _7217_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net96),
    .D(net403),
    .Q_N(_3475_),
    .Q(\dtop.player_inst.synth.alu.registers[5][4] ));
 sg13g2_dfrbp_1 _7218_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net94),
    .D(_0193_),
    .Q_N(_3474_),
    .Q(\dtop.player_inst.synth.alu.registers[5][5] ));
 sg13g2_dfrbp_1 _7219_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net92),
    .D(_0194_),
    .Q_N(_3473_),
    .Q(\dtop.player_inst.synth.alu.registers[5][6] ));
 sg13g2_dfrbp_1 _7220_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net90),
    .D(_0195_),
    .Q_N(_3472_),
    .Q(\dtop.player_inst.synth.alu.registers[3][0] ));
 sg13g2_dfrbp_1 _7221_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net88),
    .D(net411),
    .Q_N(_3471_),
    .Q(\dtop.player_inst.synth.alu.registers[3][1] ));
 sg13g2_dfrbp_1 _7222_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net86),
    .D(_0197_),
    .Q_N(_3470_),
    .Q(\dtop.player_inst.synth.alu.registers[3][2] ));
 sg13g2_dfrbp_1 _7223_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net84),
    .D(_0198_),
    .Q_N(_3469_),
    .Q(\dtop.player_inst.synth.alu.registers[3][3] ));
 sg13g2_dfrbp_1 _7224_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net82),
    .D(net392),
    .Q_N(_3468_),
    .Q(\dtop.player_inst.synth.alu.registers[3][4] ));
 sg13g2_dfrbp_1 _7225_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net80),
    .D(_0200_),
    .Q_N(_3467_),
    .Q(\dtop.player_inst.synth.alu.registers[3][5] ));
 sg13g2_dfrbp_1 _7226_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net78),
    .D(net352),
    .Q_N(_3466_),
    .Q(\dtop.player_inst.synth.alu.registers[3][6] ));
 sg13g2_dfrbp_1 _7227_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net76),
    .D(net360),
    .Q_N(_3465_),
    .Q(\dtop.player_inst.synth.alu.registers[3][7] ));
 sg13g2_dfrbp_1 _7228_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net74),
    .D(_0203_),
    .Q_N(_0025_),
    .Q(\dtop.detune_counter[4] ));
 sg13g2_dfrbp_1 _7229_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net73),
    .D(_0204_),
    .Q_N(_0077_),
    .Q(\dtop.detune_counter[5] ));
 sg13g2_dfrbp_1 _7230_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net72),
    .D(_0205_),
    .Q_N(_0023_),
    .Q(\dtop.detune_counter[6] ));
 sg13g2_dfrbp_1 _7231_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net71),
    .D(_0206_),
    .Q_N(_0021_),
    .Q(\dtop.detune_counter[7] ));
 sg13g2_dfrbp_1 _7232_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net70),
    .D(_0207_),
    .Q_N(_0020_),
    .Q(\dtop.detune_counter[8] ));
 sg13g2_dfrbp_1 _7233_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net69),
    .D(_0208_),
    .Q_N(_0018_),
    .Q(\dtop.detune_counter[9] ));
 sg13g2_dfrbp_1 _7234_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net68),
    .D(_0209_),
    .Q_N(_0016_),
    .Q(\dtop.detune_counter[10] ));
 sg13g2_dfrbp_1 _7235_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net67),
    .D(_0210_),
    .Q_N(_0000_),
    .Q(\dtop.detune_counter[11] ));
 sg13g2_dfrbp_1 _7236_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net66),
    .D(_0211_),
    .Q_N(_0014_),
    .Q(\dtop.detune_counter[12] ));
 sg13g2_dfrbp_1 _7237_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net65),
    .D(_0212_),
    .Q_N(_0059_),
    .Q(\dtop.detune_counter[13] ));
 sg13g2_dfrbp_1 _7238_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net64),
    .D(net569),
    .Q_N(_0090_),
    .Q(\dtop.detune_counter[14] ));
 sg13g2_dfrbp_1 _7239_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net63),
    .D(_0214_),
    .Q_N(_0062_),
    .Q(\dtop.detune_counter[15] ));
 sg13g2_dfrbp_1 _7240_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net62),
    .D(_0215_),
    .Q_N(_0089_),
    .Q(\dtop.detune_counter[16] ));
 sg13g2_dfrbp_1 _7241_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net61),
    .D(_0216_),
    .Q_N(_0088_),
    .Q(\dtop.detune_counter[17] ));
 sg13g2_dfrbp_1 _7242_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net60),
    .D(_0217_),
    .Q_N(_0031_),
    .Q(\dtop.vtop.dphases[0][0] ));
 sg13g2_dfrbp_1 _7243_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net59),
    .D(_0218_),
    .Q_N(_0033_),
    .Q(\dtop.vtop.dphases[0][1] ));
 sg13g2_dfrbp_1 _7244_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net58),
    .D(_0219_),
    .Q_N(_0035_),
    .Q(\dtop.vtop.dphases[0][2] ));
 sg13g2_dfrbp_1 _7245_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net57),
    .D(_0220_),
    .Q_N(_0037_),
    .Q(\dtop.vtop.dphases[0][3] ));
 sg13g2_dfrbp_1 _7246_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net56),
    .D(_0221_),
    .Q_N(_0039_),
    .Q(\dtop.vtop.dphases[0][4] ));
 sg13g2_dfrbp_1 _7247_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net55),
    .D(_0222_),
    .Q_N(_0041_),
    .Q(\dtop.vtop.dphases[0][5] ));
 sg13g2_dfrbp_1 _7248_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net54),
    .D(_0223_),
    .Q_N(_0043_),
    .Q(\dtop.vtop.dphases[0][6] ));
 sg13g2_dfrbp_1 _7249_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net53),
    .D(_0224_),
    .Q_N(_0045_),
    .Q(\dtop.vtop.dphases[0][7] ));
 sg13g2_dfrbp_1 _7250_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net52),
    .D(_0225_),
    .Q_N(_0048_),
    .Q(\dtop.vtop.dphases[0][8] ));
 sg13g2_dfrbp_1 _7251_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net51),
    .D(net375),
    .Q_N(_0050_),
    .Q(\dtop.vtop.dphases[0][9] ));
 sg13g2_dfrbp_1 _7252_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net50),
    .D(net345),
    .Q_N(_0053_),
    .Q(\dtop.vtop.dphases[0][10] ));
 sg13g2_dfrbp_1 _7253_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net49),
    .D(_0228_),
    .Q_N(_3464_),
    .Q(\dtop.vtop.dphases[1][0] ));
 sg13g2_dfrbp_1 _7254_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net48),
    .D(_0229_),
    .Q_N(_3463_),
    .Q(\dtop.vtop.dphases[1][1] ));
 sg13g2_dfrbp_1 _7255_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net47),
    .D(_0230_),
    .Q_N(_3462_),
    .Q(\dtop.vtop.dphases[1][2] ));
 sg13g2_dfrbp_1 _7256_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net46),
    .D(_0231_),
    .Q_N(_3461_),
    .Q(\dtop.vtop.dphases[1][3] ));
 sg13g2_dfrbp_1 _7257_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net45),
    .D(_0232_),
    .Q_N(_3460_),
    .Q(\dtop.vtop.dphases[1][4] ));
 sg13g2_dfrbp_1 _7258_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net44),
    .D(_0233_),
    .Q_N(_3459_),
    .Q(\dtop.vtop.dphases[1][5] ));
 sg13g2_dfrbp_1 _7259_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net43),
    .D(_0234_),
    .Q_N(_3458_),
    .Q(\dtop.vtop.dphases[1][6] ));
 sg13g2_dfrbp_1 _7260_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net42),
    .D(_0235_),
    .Q_N(_3457_),
    .Q(\dtop.vtop.dphases[1][7] ));
 sg13g2_dfrbp_1 _7261_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net41),
    .D(_0236_),
    .Q_N(_3456_),
    .Q(\dtop.vtop.dphases[1][8] ));
 sg13g2_dfrbp_1 _7262_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net40),
    .D(_0237_),
    .Q_N(_3455_),
    .Q(\dtop.vtop.dphases[1][9] ));
 sg13g2_dfrbp_1 _7263_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net39),
    .D(net400),
    .Q_N(_3454_),
    .Q(\dtop.vtop.dphases[1][10] ));
 sg13g2_dfrbp_1 _7264_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net38),
    .D(_0239_),
    .Q_N(_3453_),
    .Q(\dtop.vtop.dphases[2][0] ));
 sg13g2_dfrbp_1 _7265_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net37),
    .D(_0240_),
    .Q_N(_3452_),
    .Q(\dtop.vtop.dphases[2][1] ));
 sg13g2_dfrbp_1 _7266_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net36),
    .D(_0241_),
    .Q_N(_3451_),
    .Q(\dtop.vtop.dphases[2][2] ));
 sg13g2_dfrbp_1 _7267_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net34),
    .D(_0242_),
    .Q_N(_3450_),
    .Q(\dtop.vtop.dphases[2][3] ));
 sg13g2_dfrbp_1 _7268_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net33),
    .D(_0243_),
    .Q_N(_3449_),
    .Q(\dtop.vtop.dphases[2][4] ));
 sg13g2_dfrbp_1 _7269_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net32),
    .D(_0244_),
    .Q_N(_3448_),
    .Q(\dtop.vtop.dphases[2][5] ));
 sg13g2_dfrbp_1 _7270_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net31),
    .D(_0245_),
    .Q_N(_3447_),
    .Q(\dtop.vtop.dphases[2][6] ));
 sg13g2_dfrbp_1 _7271_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net30),
    .D(_0246_),
    .Q_N(_3446_),
    .Q(\dtop.vtop.dphases[2][7] ));
 sg13g2_dfrbp_1 _7272_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net29),
    .D(_0247_),
    .Q_N(_3445_),
    .Q(\dtop.vtop.dphases[2][8] ));
 sg13g2_dfrbp_1 _7273_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net28),
    .D(_0248_),
    .Q_N(_3444_),
    .Q(\dtop.vtop.dphases[2][9] ));
 sg13g2_dfrbp_1 _7274_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net27),
    .D(net503),
    .Q_N(_3443_),
    .Q(\dtop.vtop.dphases[2][10] ));
 sg13g2_dfrbp_1 _7275_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net26),
    .D(_0250_),
    .Q_N(_3442_),
    .Q(\dtop.player_inst.synth.alu.oct_en ));
 sg13g2_dfrbp_1 _7276_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net25),
    .D(_0251_),
    .Q_N(_3441_),
    .Q(\dtop.vtop.rs.saturated ));
 sg13g2_dfrbp_1 _7277_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net24),
    .D(net322),
    .Q_N(\uio_out0b[5] ),
    .Q(\dtop.vsync ));
 sg13g2_dfrbp_1 _7278_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net23),
    .D(net639),
    .Q_N(_3440_),
    .Q(uio_oe[5]));
 sg13g2_dfrbp_1 _7279_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net22),
    .D(_0254_),
    .Q_N(_3439_),
    .Q(\dtop.vtop.rs.scan_y.phase[0] ));
 sg13g2_dfrbp_1 _7280_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net21),
    .D(net605),
    .Q_N(_3438_),
    .Q(\dtop.vtop.rs.scan_y.phase[1] ));
 sg13g2_dfrbp_1 _7281_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net20),
    .D(_0256_),
    .Q_N(_3437_),
    .Q(\dtop.vtop.rs.x_scan.phase[0] ));
 sg13g2_dfrbp_1 _7282_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net19),
    .D(_0257_),
    .Q_N(_3436_),
    .Q(\dtop.vtop.rs.x_scan.phase[1] ));
 sg13g2_dfrbp_1 _7283_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net18),
    .D(net679),
    .Q_N(_3435_),
    .Q(\dtop.player_inst.program_addr[0] ));
 sg13g2_dfrbp_1 _7284_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net10),
    .D(_0259_),
    .Q_N(_0003_),
    .Q(\dtop.player_inst.program_addr[1] ));
 sg13g2_dfrbp_1 _7285_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net315),
    .D(_0260_),
    .Q_N(_0001_),
    .Q(\dtop.player_inst.program_addr[2] ));
 sg13g2_dfrbp_1 _7286_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net314),
    .D(net660),
    .Q_N(_0093_),
    .Q(\dtop.player_inst.program_addr[3] ));
 sg13g2_dfrbp_1 _7287_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net313),
    .D(net673),
    .Q_N(_3434_),
    .Q(\dtop.player_inst.program_addr[4] ));
 sg13g2_dfrbp_1 _7288_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net312),
    .D(net684),
    .Q_N(_0092_),
    .Q(\dtop.player_inst.program_addr[5] ));
 sg13g2_dfrbp_1 _7289_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net311),
    .D(_0264_),
    .Q_N(_0086_),
    .Q(\dtop.player_inst.program_addr[6] ));
 sg13g2_dfrbp_1 _7290_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net310),
    .D(_0265_),
    .Q_N(_3433_),
    .Q(\dtop.vtop.pipeline.nstep_zg[0] ));
 sg13g2_dfrbp_1 _7291_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net309),
    .D(net682),
    .Q_N(_3432_),
    .Q(\dtop.vtop.pipeline.nstep_zg[1] ));
 sg13g2_dfrbp_1 _7292_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net308),
    .D(net611),
    .Q_N(_0075_),
    .Q(\dtop.vtop.pipeline.neg_t[0] ));
 sg13g2_dfrbp_1 _7293_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net306),
    .D(_0268_),
    .Q_N(_0024_),
    .Q(\dtop.vtop.pipeline.neg_t[1] ));
 sg13g2_dfrbp_1 _7294_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net304),
    .D(_0269_),
    .Q_N(_0022_),
    .Q(\dtop.vtop.pipeline.neg_t[2] ));
 sg13g2_dfrbp_1 _7295_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net302),
    .D(net626),
    .Q_N(_0066_),
    .Q(\dtop.vtop.pipeline.neg_t[3] ));
 sg13g2_dfrbp_1 _7296_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net300),
    .D(_0271_),
    .Q_N(_0019_),
    .Q(\dtop.vtop.pipeline.neg_t[4] ));
 sg13g2_dfrbp_1 _7297_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net298),
    .D(_0272_),
    .Q_N(_0017_),
    .Q(\dtop.vtop.pipeline.neg_t[5] ));
 sg13g2_dfrbp_1 _7298_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net296),
    .D(_0273_),
    .Q_N(_0015_),
    .Q(\dtop.vtop.pipeline.neg_t[6] ));
 sg13g2_dfrbp_1 _7299_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net294),
    .D(_0274_),
    .Q_N(_0073_),
    .Q(\dtop.vtop.pipeline.neg_t[7] ));
 sg13g2_dfrbp_1 _7300_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net292),
    .D(net530),
    .Q_N(_0013_),
    .Q(\dtop.vtop.pipeline.neg_t[8] ));
 sg13g2_dfrbp_1 _7301_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net290),
    .D(net578),
    .Q_N(_0026_),
    .Q(\dtop.vtop.pipeline.neg_t[9] ));
 sg13g2_dfrbp_1 _7302_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net288),
    .D(_0277_),
    .Q_N(_0076_),
    .Q(\dtop.vtop.pipeline.dz[0] ));
 sg13g2_dfrbp_1 _7303_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net286),
    .D(_0278_),
    .Q_N(_0065_),
    .Q(\dtop.vtop.pipeline.dz[1] ));
 sg13g2_dfrbp_1 _7304_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net284),
    .D(_0279_),
    .Q_N(_0099_),
    .Q(\dtop.vtop.pipeline.dz[2] ));
 sg13g2_dfrbp_1 _7305_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net282),
    .D(net521),
    .Q_N(_0098_),
    .Q(\dtop.vtop.pipeline.dz[3] ));
 sg13g2_dfrbp_1 _7306_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net280),
    .D(net618),
    .Q_N(_0072_),
    .Q(\dtop.vtop.pipeline.dz[4] ));
 sg13g2_dfrbp_1 _7307_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net278),
    .D(_0282_),
    .Q_N(_0097_),
    .Q(\dtop.vtop.pipeline.dz[5] ));
 sg13g2_dfrbp_1 _7308_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net276),
    .D(_0283_),
    .Q_N(_0096_),
    .Q(\dtop.vtop.pipeline.dz[6] ));
 sg13g2_dfrbp_1 _7309_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net274),
    .D(_0284_),
    .Q_N(_0095_),
    .Q(\dtop.vtop.pipeline.dz[7] ));
 sg13g2_dfrbp_1 _7310_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net272),
    .D(_0285_),
    .Q_N(_0094_),
    .Q(\dtop.vtop.pipeline.dz[8] ));
 sg13g2_dfrbp_1 _7311_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net270),
    .D(net489),
    .Q_N(_3431_),
    .Q(\dtop.vtop.pipeline.z[0] ));
 sg13g2_dfrbp_1 _7312_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net268),
    .D(net643),
    .Q_N(_3430_),
    .Q(\dtop.vtop.pipeline.z[1] ));
 sg13g2_dfrbp_1 _7313_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net266),
    .D(_0288_),
    .Q_N(_3429_),
    .Q(\dtop.vtop.pipeline.z[2] ));
 sg13g2_dfrbp_1 _7314_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net264),
    .D(_0289_),
    .Q_N(_3428_),
    .Q(\dtop.vtop.pipeline.z[3] ));
 sg13g2_dfrbp_1 _7315_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net262),
    .D(_0290_),
    .Q_N(_3427_),
    .Q(\dtop.vtop.pipeline.z[4] ));
 sg13g2_dfrbp_1 _7316_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net260),
    .D(_0291_),
    .Q_N(_3426_),
    .Q(\dtop.vtop.pipeline.z[5] ));
 sg13g2_dfrbp_1 _7317_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net254),
    .D(_0292_),
    .Q_N(_3425_),
    .Q(\dtop.vtop.pipeline.z[6] ));
 sg13g2_dfrbp_1 _7318_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net250),
    .D(_0293_),
    .Q_N(_3424_),
    .Q(\dtop.vtop.pipeline.z[7] ));
 sg13g2_dfrbp_1 _7319_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net246),
    .D(_0294_),
    .Q_N(_3423_),
    .Q(\dtop.vtop.pipeline.z[8] ));
 sg13g2_dfrbp_1 _7320_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net223),
    .D(_0295_),
    .Q_N(_3422_),
    .Q(\dtop.vtop.pipeline.z[9] ));
 sg13g2_dfrbp_1 _7321_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net219),
    .D(_0296_),
    .Q_N(_3421_),
    .Q(\dtop.vtop.pipeline.z[10] ));
 sg13g2_dfrbp_1 _7322_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net215),
    .D(_0297_),
    .Q_N(_3420_),
    .Q(\dtop.vtop.pipeline.z[11] ));
 sg13g2_dfrbp_1 _7323_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net211),
    .D(net620),
    .Q_N(_3419_),
    .Q(\dtop.vtop.pipeline.z[12] ));
 sg13g2_dfrbp_1 _7324_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net207),
    .D(_0299_),
    .Q_N(_3418_),
    .Q(\dtop.vtop.pipeline.z[13] ));
 sg13g2_dfrbp_1 _7325_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net203),
    .D(_0300_),
    .Q_N(_3417_),
    .Q(\dtop.vtop.pipeline.z[14] ));
 sg13g2_dfrbp_1 _7326_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net199),
    .D(net449),
    .Q_N(_3416_),
    .Q(\dtop.vtop.pipeline.phases[1][0] ));
 sg13g2_dfrbp_1 _7327_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net197),
    .D(_0302_),
    .Q_N(_3415_),
    .Q(\dtop.vtop.pipeline.phases[1][1] ));
 sg13g2_dfrbp_1 _7328_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net195),
    .D(_0303_),
    .Q_N(_3414_),
    .Q(\dtop.vtop.pipeline.phases[1][2] ));
 sg13g2_dfrbp_1 _7329_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net193),
    .D(_0304_),
    .Q_N(_3413_),
    .Q(\dtop.vtop.pipeline.phases[1][3] ));
 sg13g2_dfrbp_1 _7330_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net191),
    .D(_0305_),
    .Q_N(_3412_),
    .Q(\dtop.vtop.pipeline.phases[1][4] ));
 sg13g2_dfrbp_1 _7331_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net189),
    .D(_0306_),
    .Q_N(_3411_),
    .Q(\dtop.vtop.pipeline.phases[1][5] ));
 sg13g2_dfrbp_1 _7332_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net187),
    .D(_0307_),
    .Q_N(_3410_),
    .Q(\dtop.vtop.pipeline.phases[1][6] ));
 sg13g2_dfrbp_1 _7333_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net185),
    .D(_0308_),
    .Q_N(_3409_),
    .Q(\dtop.vtop.pipeline.phases[1][7] ));
 sg13g2_dfrbp_1 _7334_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net183),
    .D(_0309_),
    .Q_N(_3408_),
    .Q(\dtop.vtop.pipeline.phases[1][8] ));
 sg13g2_dfrbp_1 _7335_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net181),
    .D(_0310_),
    .Q_N(_3407_),
    .Q(\dtop.vtop.pipeline.phases[1][9] ));
 sg13g2_dfrbp_1 _7336_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net179),
    .D(_0311_),
    .Q_N(_3406_),
    .Q(\dtop.vtop.pipeline.phases[1][10] ));
 sg13g2_dfrbp_1 _7337_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net177),
    .D(_0312_),
    .Q_N(_3405_),
    .Q(\dtop.vtop.pipeline.phases[1][11] ));
 sg13g2_dfrbp_1 _7338_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net175),
    .D(_0313_),
    .Q_N(_3404_),
    .Q(\dtop.vtop.pipeline.phases[1][12] ));
 sg13g2_dfrbp_1 _7339_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net173),
    .D(_0314_),
    .Q_N(_3403_),
    .Q(\dtop.vtop.pipeline.phases[1][13] ));
 sg13g2_dfrbp_1 _7340_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net171),
    .D(_0315_),
    .Q_N(_3402_),
    .Q(\dtop.vtop.pipeline.phases[1][14] ));
 sg13g2_dfrbp_1 _7341_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net169),
    .D(_0316_),
    .Q_N(_3401_),
    .Q(\dtop.vtop.pipeline.phases[1][15] ));
 sg13g2_dfrbp_1 _7342_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net167),
    .D(net497),
    .Q_N(_3400_),
    .Q(\dtop.vtop.pipeline.phases[2][0] ));
 sg13g2_dfrbp_1 _7343_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net165),
    .D(_0318_),
    .Q_N(_3399_),
    .Q(\dtop.vtop.pipeline.phases[2][1] ));
 sg13g2_dfrbp_1 _7344_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net163),
    .D(_0319_),
    .Q_N(_3398_),
    .Q(\dtop.vtop.pipeline.phases[2][2] ));
 sg13g2_dfrbp_1 _7345_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net161),
    .D(_0320_),
    .Q_N(_3397_),
    .Q(\dtop.vtop.pipeline.phases[2][3] ));
 sg13g2_dfrbp_1 _7346_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net159),
    .D(_0321_),
    .Q_N(_3396_),
    .Q(\dtop.vtop.pipeline.phases[2][4] ));
 sg13g2_dfrbp_1 _7347_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net157),
    .D(_0322_),
    .Q_N(_3395_),
    .Q(\dtop.vtop.pipeline.phases[2][5] ));
 sg13g2_dfrbp_1 _7348_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net155),
    .D(_0323_),
    .Q_N(_3394_),
    .Q(\dtop.vtop.pipeline.phases[2][6] ));
 sg13g2_dfrbp_1 _7349_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net153),
    .D(_0324_),
    .Q_N(_3393_),
    .Q(\dtop.vtop.pipeline.phases[2][7] ));
 sg13g2_dfrbp_1 _7350_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net151),
    .D(_0325_),
    .Q_N(_3392_),
    .Q(\dtop.vtop.pipeline.phases[2][8] ));
 sg13g2_dfrbp_1 _7351_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net149),
    .D(_0326_),
    .Q_N(_3391_),
    .Q(\dtop.vtop.pipeline.phases[2][9] ));
 sg13g2_dfrbp_1 _7352_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net147),
    .D(_0327_),
    .Q_N(_3390_),
    .Q(\dtop.vtop.pipeline.phases[2][10] ));
 sg13g2_dfrbp_1 _7353_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net145),
    .D(_0328_),
    .Q_N(_3389_),
    .Q(\dtop.vtop.pipeline.phases[2][11] ));
 sg13g2_dfrbp_1 _7354_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net143),
    .D(_0329_),
    .Q_N(_3388_),
    .Q(\dtop.vtop.pipeline.phases[2][12] ));
 sg13g2_dfrbp_1 _7355_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net141),
    .D(_0330_),
    .Q_N(_3387_),
    .Q(\dtop.vtop.pipeline.phases[2][13] ));
 sg13g2_dfrbp_1 _7356_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net139),
    .D(_0331_),
    .Q_N(_3386_),
    .Q(\dtop.vtop.pipeline.phases[2][14] ));
 sg13g2_dfrbp_1 _7357_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net137),
    .D(_0332_),
    .Q_N(_3385_),
    .Q(\dtop.vtop.pipeline.phases[2][15] ));
 sg13g2_dfrbp_1 _7358_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net135),
    .D(_0333_),
    .Q_N(_3353_),
    .Q(\dtop.enable ));
 sg13g2_dfrbp_1 _7359_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net133),
    .D(_0334_),
    .Q_N(_0012_),
    .Q(\dtop.vtop.color[6] ));
 sg13g2_dfrbp_1 _7360_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net131),
    .D(_0335_),
    .Q_N(_0011_),
    .Q(\dtop.vtop.color[7] ));
 sg13g2_dfrbp_1 _7361_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net129),
    .D(_0336_),
    .Q_N(_0010_),
    .Q(\dtop.vtop.color[8] ));
 sg13g2_dfrbp_1 _7362_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net127),
    .D(_0337_),
    .Q_N(_0007_),
    .Q(\dtop.vtop.color[9] ));
 sg13g2_dfrbp_1 _7363_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net125),
    .D(_0338_),
    .Q_N(_0009_),
    .Q(\dtop.vtop.color[10] ));
 sg13g2_dfrbp_1 _7364_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net123),
    .D(_0339_),
    .Q_N(_0008_),
    .Q(\dtop.vtop.color[11] ));
 sg13g2_dfrbp_1 _7365_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net121),
    .D(_0340_),
    .Q_N(_3384_),
    .Q(\dtop.vtop.pipeline.zg[0] ));
 sg13g2_dfrbp_1 _7366_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net119),
    .D(_0341_),
    .Q_N(_3383_),
    .Q(\dtop.vtop.pipeline.zg[1] ));
 sg13g2_dfrbp_1 _7367_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net117),
    .D(_0342_),
    .Q_N(_3382_),
    .Q(\dtop.vtop.pipeline.zg[2] ));
 sg13g2_dfrbp_1 _7368_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net115),
    .D(_0343_),
    .Q_N(_3381_),
    .Q(\dtop.vtop.pipeline.zg[3] ));
 sg13g2_dfrbp_1 _7369_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net113),
    .D(_0344_),
    .Q_N(_3380_),
    .Q(\dtop.vtop.pipeline.zg[4] ));
 sg13g2_dfrbp_1 _7370_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net111),
    .D(_0345_),
    .Q_N(_0028_),
    .Q(\dtop.vtop.pipeline.zg[5] ));
 sg13g2_dfrbp_1 _7371_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net109),
    .D(_0346_),
    .Q_N(_3379_),
    .Q(\dtop.vtop.pipeline.zg[6] ));
 sg13g2_dfrbp_1 _7372_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net107),
    .D(_0347_),
    .Q_N(_0027_),
    .Q(\dtop.vtop.pipeline.zg[7] ));
 sg13g2_dfrbp_1 _7373_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net105),
    .D(_0348_),
    .Q_N(_3378_),
    .Q(\dtop.vtop.pipeline.zg[8] ));
 sg13g2_dfrbp_1 _7374_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net103),
    .D(_0349_),
    .Q_N(_3377_),
    .Q(\dtop.vtop.pipeline.zg[9] ));
 sg13g2_dfrbp_1 _7375_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net101),
    .D(_0350_),
    .Q_N(_3376_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[0] ));
 sg13g2_dfrbp_1 _7376_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net99),
    .D(net377),
    .Q_N(_3375_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[1] ));
 sg13g2_dfrbp_1 _7377_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net97),
    .D(_0352_),
    .Q_N(_3374_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[2] ));
 sg13g2_dfrbp_1 _7378_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net95),
    .D(_0353_),
    .Q_N(_3373_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[3] ));
 sg13g2_dfrbp_1 _7379_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net93),
    .D(_0354_),
    .Q_N(_3372_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[4] ));
 sg13g2_dfrbp_1 _7380_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net91),
    .D(_0355_),
    .Q_N(_3371_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[5] ));
 sg13g2_dfrbp_1 _7381_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net89),
    .D(_0356_),
    .Q_N(_3370_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[6] ));
 sg13g2_dfrbp_1 _7382_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net87),
    .D(_0357_),
    .Q_N(_3369_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[7] ));
 sg13g2_dfrbp_1 _7383_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net85),
    .D(_0358_),
    .Q_N(_3368_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[8] ));
 sg13g2_dfrbp_1 _7384_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net83),
    .D(_0359_),
    .Q_N(_3367_),
    .Q(\dtop.vtop.pipeline.zg_acc[0] ));
 sg13g2_dfrbp_1 _7385_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net81),
    .D(_0360_),
    .Q_N(_3366_),
    .Q(\dtop.vtop.pipeline.zg_acc[1] ));
 sg13g2_dfrbp_1 _7386_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net79),
    .D(_0361_),
    .Q_N(_3365_),
    .Q(\dtop.vtop.pipeline.zg_acc[2] ));
 sg13g2_dfrbp_1 _7387_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net77),
    .D(_0362_),
    .Q_N(_3364_),
    .Q(\dtop.vtop.pipeline.zg_acc[3] ));
 sg13g2_dfrbp_1 _7388_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net75),
    .D(_0363_),
    .Q_N(_3363_),
    .Q(\dtop.vtop.pipeline.zg_acc[4] ));
 sg13g2_dfrbp_1 _7389_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net307),
    .D(_0364_),
    .Q_N(_3362_),
    .Q(\dtop.vtop.pipeline.zg_acc[5] ));
 sg13g2_dfrbp_1 _7390_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net305),
    .D(_0365_),
    .Q_N(_0058_),
    .Q(\dtop.vtop.pipeline.zg_acc[6] ));
 sg13g2_dfrbp_1 _7391_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net303),
    .D(_0366_),
    .Q_N(_0061_),
    .Q(\dtop.vtop.pipeline.zg_acc[7] ));
 sg13g2_dfrbp_1 _7392_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net301),
    .D(_0367_),
    .Q_N(_0074_),
    .Q(\dtop.vtop.pipeline.zg_acc[8] ));
 sg13g2_dfrbp_1 _7393_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net299),
    .D(_0368_),
    .Q_N(_3361_),
    .Q(\dtop.vtop.pipeline.zg_acc[9] ));
 sg13g2_dfrbp_1 _7394_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net297),
    .D(_0369_),
    .Q_N(_0091_),
    .Q(\dtop.vtop.pipeline.zg_valid ));
 sg13g2_dfrbp_1 _7395_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net293),
    .D(net633),
    .Q_N(_0004_),
    .Q(\dtop.vtop.pipeline.wave_index[0] ));
 sg13g2_dfrbp_1 _7396_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net291),
    .D(_0371_),
    .Q_N(_0005_),
    .Q(\dtop.vtop.pipeline.wave_index[1] ));
 sg13g2_dfrbp_1 _7397_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net289),
    .D(_0372_),
    .Q_N(_3360_),
    .Q(\dtop.vtop.pipeline.nstep[0] ));
 sg13g2_dfrbp_1 _7398_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net287),
    .D(_0373_),
    .Q_N(_0030_),
    .Q(\dtop.vtop.pipeline.nstep[1] ));
 sg13g2_dfrbp_1 _7399_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net285),
    .D(net319),
    .Q_N(\dtop.vtop.pipeline.next_nstep_counter[0] ),
    .Q(\dtop.vtop.pipeline.nstep_counter[0] ));
 sg13g2_dfrbp_1 _7400_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net281),
    .D(net556),
    .Q_N(_3359_),
    .Q(\dtop.vtop.pipeline.nstep_counter[1] ));
 sg13g2_dfrbp_1 _7401_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net277),
    .D(net594),
    .Q_N(_3358_),
    .Q(\dtop.vtop.pipeline.nstep_counter[2] ));
 sg13g2_dfrbp_1 _7402_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net273),
    .D(net539),
    .Q_N(_3357_),
    .Q(\dtop.vtop.pipeline.nstep_counter[3] ));
 sg13g2_dfrbp_1 _7403_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net269),
    .D(net493),
    .Q_N(_3356_),
    .Q(\dtop.vtop.pipeline.nstep_counter[4] ));
 sg13g2_dfrbp_1 _7404_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net265),
    .D(net371),
    .Q_N(_0029_),
    .Q(\dtop.vtop.pipeline.phases[0][0] ));
 sg13g2_dfrbp_1 _7405_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net263),
    .D(_0380_),
    .Q_N(_0032_),
    .Q(\dtop.vtop.pipeline.phases[0][1] ));
 sg13g2_dfrbp_1 _7406_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net261),
    .D(_0381_),
    .Q_N(_0034_),
    .Q(\dtop.vtop.pipeline.phases[0][2] ));
 sg13g2_dfrbp_1 _7407_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net259),
    .D(_0382_),
    .Q_N(_0036_),
    .Q(\dtop.vtop.pipeline.phases[0][3] ));
 sg13g2_dfrbp_1 _7408_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net252),
    .D(_0383_),
    .Q_N(_0038_),
    .Q(\dtop.vtop.pipeline.phases[0][4] ));
 sg13g2_dfrbp_1 _7409_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net248),
    .D(_0384_),
    .Q_N(_0040_),
    .Q(\dtop.vtop.pipeline.phases[0][5] ));
 sg13g2_dfrbp_1 _7410_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net244),
    .D(_0385_),
    .Q_N(_0042_),
    .Q(\dtop.vtop.pipeline.phases[0][6] ));
 sg13g2_dfrbp_1 _7411_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net221),
    .D(_0386_),
    .Q_N(_0044_),
    .Q(\dtop.vtop.pipeline.phases[0][7] ));
 sg13g2_dfrbp_1 _7412_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net217),
    .D(_0387_),
    .Q_N(_0047_),
    .Q(\dtop.vtop.pipeline.phases[0][8] ));
 sg13g2_dfrbp_1 _7413_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net213),
    .D(_0388_),
    .Q_N(_0049_),
    .Q(\dtop.vtop.pipeline.phases[0][9] ));
 sg13g2_dfrbp_1 _7414_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net209),
    .D(_0389_),
    .Q_N(_0052_),
    .Q(\dtop.vtop.pipeline.phases[0][10] ));
 sg13g2_dfrbp_1 _7415_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net205),
    .D(_0390_),
    .Q_N(_0054_),
    .Q(\dtop.vtop.pipeline.phases[0][11] ));
 sg13g2_dfrbp_1 _7416_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net201),
    .D(_0391_),
    .Q_N(_0056_),
    .Q(\dtop.vtop.pipeline.phases[0][12] ));
 sg13g2_dfrbp_1 _7417_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net295),
    .D(_0392_),
    .Q_N(_0057_),
    .Q(\dtop.vtop.pipeline.phases[0][13] ));
 sg13g2_dfrbp_1 _7418_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net283),
    .D(_0393_),
    .Q_N(_0060_),
    .Q(\dtop.vtop.pipeline.phases[0][14] ));
 sg13g2_dfrbp_1 _7419_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net279),
    .D(_0394_),
    .Q_N(_0002_),
    .Q(\dtop.vtop.pipeline.phases[0][15] ));
 sg13g2_dfrbp_1 _7420_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net275),
    .D(_0395_),
    .Q_N(_3355_),
    .Q(\dtop.vtop.logo_d[1] ));
 sg13g2_dfrbp_1 _7421_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net271),
    .D(_0396_),
    .Q_N(_3354_),
    .Q(\dtop.vtop.force_sat0 ));
 sg13g2_tiehi _7123__11 (.L_HI(net11));
 sg13g2_tiehi _7116__12 (.L_HI(net12));
 sg13g2_tiehi _7117__13 (.L_HI(net13));
 sg13g2_tiehi _7118__14 (.L_HI(net14));
 sg13g2_tiehi _7119__15 (.L_HI(net15));
 sg13g2_tiehi _7120__16 (.L_HI(net16));
 sg13g2_tiehi _7121__17 (.L_HI(net17));
 sg13g2_tiehi _7283__18 (.L_HI(net18));
 sg13g2_tiehi _7282__19 (.L_HI(net19));
 sg13g2_tiehi _7281__20 (.L_HI(net20));
 sg13g2_tiehi _7280__21 (.L_HI(net21));
 sg13g2_tiehi _7279__22 (.L_HI(net22));
 sg13g2_tiehi _7278__23 (.L_HI(net23));
 sg13g2_tiehi _7277__24 (.L_HI(net24));
 sg13g2_tiehi _7276__25 (.L_HI(net25));
 sg13g2_tiehi _7275__26 (.L_HI(net26));
 sg13g2_tiehi _7274__27 (.L_HI(net27));
 sg13g2_tiehi _7273__28 (.L_HI(net28));
 sg13g2_tiehi _7272__29 (.L_HI(net29));
 sg13g2_tiehi _7271__30 (.L_HI(net30));
 sg13g2_tiehi _7270__31 (.L_HI(net31));
 sg13g2_tiehi _7269__32 (.L_HI(net32));
 sg13g2_tiehi _7268__33 (.L_HI(net33));
 sg13g2_tiehi _7267__34 (.L_HI(net34));
 sg13g2_tiehi _7122__35 (.L_HI(net35));
 sg13g2_tiehi _7266__36 (.L_HI(net36));
 sg13g2_tiehi _7265__37 (.L_HI(net37));
 sg13g2_tiehi _7264__38 (.L_HI(net38));
 sg13g2_tiehi _7263__39 (.L_HI(net39));
 sg13g2_tiehi _7262__40 (.L_HI(net40));
 sg13g2_tiehi _7261__41 (.L_HI(net41));
 sg13g2_tiehi _7260__42 (.L_HI(net42));
 sg13g2_tiehi _7259__43 (.L_HI(net43));
 sg13g2_tiehi _7258__44 (.L_HI(net44));
 sg13g2_tiehi _7257__45 (.L_HI(net45));
 sg13g2_tiehi _7256__46 (.L_HI(net46));
 sg13g2_tiehi _7255__47 (.L_HI(net47));
 sg13g2_tiehi _7254__48 (.L_HI(net48));
 sg13g2_tiehi _7253__49 (.L_HI(net49));
 sg13g2_tiehi _7252__50 (.L_HI(net50));
 sg13g2_tiehi _7251__51 (.L_HI(net51));
 sg13g2_tiehi _7250__52 (.L_HI(net52));
 sg13g2_tiehi _7249__53 (.L_HI(net53));
 sg13g2_tiehi _7248__54 (.L_HI(net54));
 sg13g2_tiehi _7247__55 (.L_HI(net55));
 sg13g2_tiehi _7246__56 (.L_HI(net56));
 sg13g2_tiehi _7245__57 (.L_HI(net57));
 sg13g2_tiehi _7244__58 (.L_HI(net58));
 sg13g2_tiehi _7243__59 (.L_HI(net59));
 sg13g2_tiehi _7242__60 (.L_HI(net60));
 sg13g2_tiehi _7241__61 (.L_HI(net61));
 sg13g2_tiehi _7240__62 (.L_HI(net62));
 sg13g2_tiehi _7239__63 (.L_HI(net63));
 sg13g2_tiehi _7238__64 (.L_HI(net64));
 sg13g2_tiehi _7237__65 (.L_HI(net65));
 sg13g2_tiehi _7236__66 (.L_HI(net66));
 sg13g2_tiehi _7235__67 (.L_HI(net67));
 sg13g2_tiehi _7234__68 (.L_HI(net68));
 sg13g2_tiehi _7233__69 (.L_HI(net69));
 sg13g2_tiehi _7232__70 (.L_HI(net70));
 sg13g2_tiehi _7231__71 (.L_HI(net71));
 sg13g2_tiehi _7230__72 (.L_HI(net72));
 sg13g2_tiehi _7229__73 (.L_HI(net73));
 sg13g2_tiehi _7228__74 (.L_HI(net74));
 sg13g2_tiehi _7388__75 (.L_HI(net75));
 sg13g2_tiehi _7227__76 (.L_HI(net76));
 sg13g2_tiehi _7387__77 (.L_HI(net77));
 sg13g2_tiehi _7226__78 (.L_HI(net78));
 sg13g2_tiehi _7386__79 (.L_HI(net79));
 sg13g2_tiehi _7225__80 (.L_HI(net80));
 sg13g2_tiehi _7385__81 (.L_HI(net81));
 sg13g2_tiehi _7224__82 (.L_HI(net82));
 sg13g2_tiehi _7384__83 (.L_HI(net83));
 sg13g2_tiehi _7223__84 (.L_HI(net84));
 sg13g2_tiehi _7383__85 (.L_HI(net85));
 sg13g2_tiehi _7222__86 (.L_HI(net86));
 sg13g2_tiehi _7382__87 (.L_HI(net87));
 sg13g2_tiehi _7221__88 (.L_HI(net88));
 sg13g2_tiehi _7381__89 (.L_HI(net89));
 sg13g2_tiehi _7220__90 (.L_HI(net90));
 sg13g2_tiehi _7380__91 (.L_HI(net91));
 sg13g2_tiehi _7219__92 (.L_HI(net92));
 sg13g2_tiehi _7379__93 (.L_HI(net93));
 sg13g2_tiehi _7218__94 (.L_HI(net94));
 sg13g2_tiehi _7378__95 (.L_HI(net95));
 sg13g2_tiehi _7217__96 (.L_HI(net96));
 sg13g2_tiehi _7377__97 (.L_HI(net97));
 sg13g2_tiehi _7216__98 (.L_HI(net98));
 sg13g2_tiehi _7376__99 (.L_HI(net99));
 sg13g2_tiehi _7215__100 (.L_HI(net100));
 sg13g2_tiehi _7375__101 (.L_HI(net101));
 sg13g2_tiehi _7214__102 (.L_HI(net102));
 sg13g2_tiehi _7374__103 (.L_HI(net103));
 sg13g2_tiehi _7213__104 (.L_HI(net104));
 sg13g2_tiehi _7373__105 (.L_HI(net105));
 sg13g2_tiehi _7212__106 (.L_HI(net106));
 sg13g2_tiehi _7372__107 (.L_HI(net107));
 sg13g2_tiehi _7211__108 (.L_HI(net108));
 sg13g2_tiehi _7371__109 (.L_HI(net109));
 sg13g2_tiehi _7210__110 (.L_HI(net110));
 sg13g2_tiehi _7370__111 (.L_HI(net111));
 sg13g2_tiehi _7209__112 (.L_HI(net112));
 sg13g2_tiehi _7369__113 (.L_HI(net113));
 sg13g2_tiehi _7208__114 (.L_HI(net114));
 sg13g2_tiehi _7368__115 (.L_HI(net115));
 sg13g2_tiehi _7207__116 (.L_HI(net116));
 sg13g2_tiehi _7367__117 (.L_HI(net117));
 sg13g2_tiehi _7206__118 (.L_HI(net118));
 sg13g2_tiehi _7366__119 (.L_HI(net119));
 sg13g2_tiehi _7205__120 (.L_HI(net120));
 sg13g2_tiehi _7365__121 (.L_HI(net121));
 sg13g2_tiehi _7204__122 (.L_HI(net122));
 sg13g2_tiehi _7364__123 (.L_HI(net123));
 sg13g2_tiehi _7203__124 (.L_HI(net124));
 sg13g2_tiehi _7363__125 (.L_HI(net125));
 sg13g2_tiehi _7202__126 (.L_HI(net126));
 sg13g2_tiehi _7362__127 (.L_HI(net127));
 sg13g2_tiehi _7201__128 (.L_HI(net128));
 sg13g2_tiehi _7361__129 (.L_HI(net129));
 sg13g2_tiehi _7200__130 (.L_HI(net130));
 sg13g2_tiehi _7360__131 (.L_HI(net131));
 sg13g2_tiehi _7199__132 (.L_HI(net132));
 sg13g2_tiehi _7359__133 (.L_HI(net133));
 sg13g2_tiehi _7198__134 (.L_HI(net134));
 sg13g2_tiehi _7358__135 (.L_HI(net135));
 sg13g2_tiehi _7197__136 (.L_HI(net136));
 sg13g2_tiehi _7357__137 (.L_HI(net137));
 sg13g2_tiehi _7196__138 (.L_HI(net138));
 sg13g2_tiehi _7356__139 (.L_HI(net139));
 sg13g2_tiehi _7195__140 (.L_HI(net140));
 sg13g2_tiehi _7355__141 (.L_HI(net141));
 sg13g2_tiehi _7194__142 (.L_HI(net142));
 sg13g2_tiehi _7354__143 (.L_HI(net143));
 sg13g2_tiehi _7193__144 (.L_HI(net144));
 sg13g2_tiehi _7353__145 (.L_HI(net145));
 sg13g2_tiehi _7192__146 (.L_HI(net146));
 sg13g2_tiehi _7352__147 (.L_HI(net147));
 sg13g2_tiehi _7191__148 (.L_HI(net148));
 sg13g2_tiehi _7351__149 (.L_HI(net149));
 sg13g2_tiehi _7190__150 (.L_HI(net150));
 sg13g2_tiehi _7350__151 (.L_HI(net151));
 sg13g2_tiehi _7189__152 (.L_HI(net152));
 sg13g2_tiehi _7349__153 (.L_HI(net153));
 sg13g2_tiehi _7188__154 (.L_HI(net154));
 sg13g2_tiehi _7348__155 (.L_HI(net155));
 sg13g2_tiehi _7187__156 (.L_HI(net156));
 sg13g2_tiehi _7347__157 (.L_HI(net157));
 sg13g2_tiehi _7186__158 (.L_HI(net158));
 sg13g2_tiehi _7346__159 (.L_HI(net159));
 sg13g2_tiehi _7185__160 (.L_HI(net160));
 sg13g2_tiehi _7345__161 (.L_HI(net161));
 sg13g2_tiehi _7184__162 (.L_HI(net162));
 sg13g2_tiehi _7344__163 (.L_HI(net163));
 sg13g2_tiehi _7183__164 (.L_HI(net164));
 sg13g2_tiehi _7343__165 (.L_HI(net165));
 sg13g2_tiehi _7182__166 (.L_HI(net166));
 sg13g2_tiehi _7342__167 (.L_HI(net167));
 sg13g2_tiehi _7181__168 (.L_HI(net168));
 sg13g2_tiehi _7341__169 (.L_HI(net169));
 sg13g2_tiehi _7180__170 (.L_HI(net170));
 sg13g2_tiehi _7340__171 (.L_HI(net171));
 sg13g2_tiehi _7179__172 (.L_HI(net172));
 sg13g2_tiehi _7339__173 (.L_HI(net173));
 sg13g2_tiehi _7178__174 (.L_HI(net174));
 sg13g2_tiehi _7338__175 (.L_HI(net175));
 sg13g2_tiehi _7177__176 (.L_HI(net176));
 sg13g2_tiehi _7337__177 (.L_HI(net177));
 sg13g2_tiehi _7176__178 (.L_HI(net178));
 sg13g2_tiehi _7336__179 (.L_HI(net179));
 sg13g2_tiehi _7175__180 (.L_HI(net180));
 sg13g2_tiehi _7335__181 (.L_HI(net181));
 sg13g2_tiehi _7174__182 (.L_HI(net182));
 sg13g2_tiehi _7334__183 (.L_HI(net183));
 sg13g2_tiehi _7173__184 (.L_HI(net184));
 sg13g2_tiehi _7333__185 (.L_HI(net185));
 sg13g2_tiehi _7172__186 (.L_HI(net186));
 sg13g2_tiehi _7332__187 (.L_HI(net187));
 sg13g2_tiehi _7171__188 (.L_HI(net188));
 sg13g2_tiehi _7331__189 (.L_HI(net189));
 sg13g2_tiehi _7170__190 (.L_HI(net190));
 sg13g2_tiehi _7330__191 (.L_HI(net191));
 sg13g2_tiehi _7169__192 (.L_HI(net192));
 sg13g2_tiehi _7329__193 (.L_HI(net193));
 sg13g2_tiehi _7168__194 (.L_HI(net194));
 sg13g2_tiehi _7328__195 (.L_HI(net195));
 sg13g2_tiehi _7167__196 (.L_HI(net196));
 sg13g2_tiehi _7327__197 (.L_HI(net197));
 sg13g2_tiehi _7166__198 (.L_HI(net198));
 sg13g2_tiehi _7326__199 (.L_HI(net199));
 sg13g2_tiehi _7165__200 (.L_HI(net200));
 sg13g2_tiehi _7416__201 (.L_HI(net201));
 sg13g2_tiehi _7164__202 (.L_HI(net202));
 sg13g2_tiehi _7325__203 (.L_HI(net203));
 sg13g2_tiehi _7163__204 (.L_HI(net204));
 sg13g2_tiehi _7415__205 (.L_HI(net205));
 sg13g2_tiehi _7162__206 (.L_HI(net206));
 sg13g2_tiehi _7324__207 (.L_HI(net207));
 sg13g2_tiehi _7161__208 (.L_HI(net208));
 sg13g2_tiehi _7414__209 (.L_HI(net209));
 sg13g2_tiehi _7160__210 (.L_HI(net210));
 sg13g2_tiehi _7323__211 (.L_HI(net211));
 sg13g2_tiehi _7159__212 (.L_HI(net212));
 sg13g2_tiehi _7413__213 (.L_HI(net213));
 sg13g2_tiehi _7158__214 (.L_HI(net214));
 sg13g2_tiehi _7322__215 (.L_HI(net215));
 sg13g2_tiehi _7157__216 (.L_HI(net216));
 sg13g2_tiehi _7412__217 (.L_HI(net217));
 sg13g2_tiehi _7156__218 (.L_HI(net218));
 sg13g2_tiehi _7321__219 (.L_HI(net219));
 sg13g2_tiehi _7155__220 (.L_HI(net220));
 sg13g2_tiehi _7411__221 (.L_HI(net221));
 sg13g2_tiehi _7154__222 (.L_HI(net222));
 sg13g2_tiehi _7320__223 (.L_HI(net223));
 sg13g2_tiehi _7153__224 (.L_HI(net224));
 sg13g2_tiehi _7152__225 (.L_HI(net225));
 sg13g2_tiehi _7151__226 (.L_HI(net226));
 sg13g2_tiehi _7150__227 (.L_HI(net227));
 sg13g2_tiehi _7149__228 (.L_HI(net228));
 sg13g2_tiehi _7148__229 (.L_HI(net229));
 sg13g2_tiehi _7147__230 (.L_HI(net230));
 sg13g2_tiehi _7146__231 (.L_HI(net231));
 sg13g2_tiehi _7145__232 (.L_HI(net232));
 sg13g2_tiehi _7144__233 (.L_HI(net233));
 sg13g2_tiehi _7143__234 (.L_HI(net234));
 sg13g2_tiehi _7142__235 (.L_HI(net235));
 sg13g2_tiehi _7141__236 (.L_HI(net236));
 sg13g2_tiehi _7139__237 (.L_HI(net237));
 sg13g2_tiehi _7138__238 (.L_HI(net238));
 sg13g2_tiehi _7137__239 (.L_HI(net239));
 sg13g2_tiehi _7136__240 (.L_HI(net240));
 sg13g2_tiehi _7135__241 (.L_HI(net241));
 sg13g2_tiehi _7134__242 (.L_HI(net242));
 sg13g2_tiehi _7133__243 (.L_HI(net243));
 sg13g2_tiehi _7410__244 (.L_HI(net244));
 sg13g2_tiehi _7132__245 (.L_HI(net245));
 sg13g2_tiehi _7319__246 (.L_HI(net246));
 sg13g2_tiehi _7131__247 (.L_HI(net247));
 sg13g2_tiehi _7409__248 (.L_HI(net248));
 sg13g2_tiehi _7130__249 (.L_HI(net249));
 sg13g2_tiehi _7318__250 (.L_HI(net250));
 sg13g2_tiehi _7129__251 (.L_HI(net251));
 sg13g2_tiehi _7408__252 (.L_HI(net252));
 sg13g2_tiehi _7128__253 (.L_HI(net253));
 sg13g2_tiehi _7317__254 (.L_HI(net254));
 sg13g2_tiehi _7127__255 (.L_HI(net255));
 sg13g2_tiehi _7126__256 (.L_HI(net256));
 sg13g2_tiehi _7125__257 (.L_HI(net257));
 sg13g2_tiehi _7124__258 (.L_HI(net258));
 sg13g2_tiehi _7407__259 (.L_HI(net259));
 sg13g2_tiehi _7316__260 (.L_HI(net260));
 sg13g2_tiehi _7406__261 (.L_HI(net261));
 sg13g2_tiehi _7315__262 (.L_HI(net262));
 sg13g2_tiehi _7405__263 (.L_HI(net263));
 sg13g2_tiehi _7314__264 (.L_HI(net264));
 sg13g2_tiehi _7404__265 (.L_HI(net265));
 sg13g2_tiehi _7313__266 (.L_HI(net266));
 sg13g2_tiehi _7140__267 (.L_HI(net267));
 sg13g2_tiehi _7312__268 (.L_HI(net268));
 sg13g2_tiehi _7403__269 (.L_HI(net269));
 sg13g2_tiehi _7311__270 (.L_HI(net270));
 sg13g2_tiehi _7421__271 (.L_HI(net271));
 sg13g2_tiehi _7310__272 (.L_HI(net272));
 sg13g2_tiehi _7402__273 (.L_HI(net273));
 sg13g2_tiehi _7309__274 (.L_HI(net274));
 sg13g2_tiehi _7420__275 (.L_HI(net275));
 sg13g2_tiehi _7308__276 (.L_HI(net276));
 sg13g2_tiehi _7401__277 (.L_HI(net277));
 sg13g2_tiehi _7307__278 (.L_HI(net278));
 sg13g2_tiehi _7419__279 (.L_HI(net279));
 sg13g2_tiehi _7306__280 (.L_HI(net280));
 sg13g2_tiehi _7400__281 (.L_HI(net281));
 sg13g2_tiehi _7305__282 (.L_HI(net282));
 sg13g2_tiehi _7418__283 (.L_HI(net283));
 sg13g2_tiehi _7304__284 (.L_HI(net284));
 sg13g2_tiehi _7399__285 (.L_HI(net285));
 sg13g2_tiehi _7303__286 (.L_HI(net286));
 sg13g2_tiehi _7398__287 (.L_HI(net287));
 sg13g2_tiehi _7302__288 (.L_HI(net288));
 sg13g2_tiehi _7397__289 (.L_HI(net289));
 sg13g2_tiehi _7301__290 (.L_HI(net290));
 sg13g2_tiehi _7396__291 (.L_HI(net291));
 sg13g2_tiehi _7300__292 (.L_HI(net292));
 sg13g2_tiehi _7395__293 (.L_HI(net293));
 sg13g2_tiehi _7299__294 (.L_HI(net294));
 sg13g2_tiehi _7417__295 (.L_HI(net295));
 sg13g2_tiehi _7298__296 (.L_HI(net296));
 sg13g2_tiehi _7394__297 (.L_HI(net297));
 sg13g2_tiehi _7297__298 (.L_HI(net298));
 sg13g2_tiehi _7393__299 (.L_HI(net299));
 sg13g2_tiehi _7296__300 (.L_HI(net300));
 sg13g2_tiehi _7392__301 (.L_HI(net301));
 sg13g2_tiehi _7295__302 (.L_HI(net302));
 sg13g2_tiehi _7391__303 (.L_HI(net303));
 sg13g2_tiehi _7294__304 (.L_HI(net304));
 sg13g2_tiehi _7390__305 (.L_HI(net305));
 sg13g2_tiehi _7293__306 (.L_HI(net306));
 sg13g2_tiehi _7389__307 (.L_HI(net307));
 sg13g2_tiehi _7292__308 (.L_HI(net308));
 sg13g2_tiehi _7291__309 (.L_HI(net309));
 sg13g2_tiehi _7290__310 (.L_HI(net310));
 sg13g2_tiehi _7289__311 (.L_HI(net311));
 sg13g2_tiehi _7288__312 (.L_HI(net312));
 sg13g2_tiehi _7287__313 (.L_HI(net313));
 sg13g2_tiehi _7286__314 (.L_HI(net314));
 sg13g2_tiehi _7285__315 (.L_HI(net315));
 sg13g2_tiehi tt_um_toivoh_demo_deluxe_316 (.L_HI(net316));
 sg13g2_tiehi tt_um_toivoh_demo_deluxe_317 (.L_HI(net317));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _7730_ (.A(uio_oe[5]),
    .X(uio_oe[0]));
 sg13g2_buf_1 _7731_ (.A(uio_oe[5]),
    .X(uio_oe[1]));
 sg13g2_buf_1 _7732_ (.A(uio_oe[5]),
    .X(uio_oe[2]));
 sg13g2_buf_1 _7733_ (.A(uio_oe[5]),
    .X(uio_oe[3]));
 sg13g2_buf_1 _7734_ (.A(uio_oe[5]),
    .X(uio_oe[4]));
 sg13g2_buf_2 fanout1095 (.A(_1513_),
    .X(net1095));
 sg13g2_buf_2 fanout1096 (.A(_1513_),
    .X(net1096));
 sg13g2_buf_2 fanout1097 (.A(net1100),
    .X(net1097));
 sg13g2_buf_2 fanout1098 (.A(net1100),
    .X(net1098));
 sg13g2_buf_2 fanout1099 (.A(net1100),
    .X(net1099));
 sg13g2_buf_2 fanout1100 (.A(_2092_),
    .X(net1100));
 sg13g2_buf_2 fanout1101 (.A(net1103),
    .X(net1101));
 sg13g2_buf_2 fanout1102 (.A(net1103),
    .X(net1102));
 sg13g2_buf_1 fanout1103 (.A(_2082_),
    .X(net1103));
 sg13g2_buf_2 fanout1104 (.A(_2761_),
    .X(net1104));
 sg13g2_buf_2 fanout1105 (.A(_2818_),
    .X(net1105));
 sg13g2_buf_2 fanout1106 (.A(_2754_),
    .X(net1106));
 sg13g2_buf_2 fanout1107 (.A(_2754_),
    .X(net1107));
 sg13g2_buf_2 fanout1108 (.A(net1110),
    .X(net1108));
 sg13g2_buf_1 fanout1109 (.A(net1110),
    .X(net1109));
 sg13g2_buf_2 fanout1110 (.A(_2729_),
    .X(net1110));
 sg13g2_buf_2 fanout1111 (.A(_0875_),
    .X(net1111));
 sg13g2_buf_4 fanout1112 (.X(net1112),
    .A(_2751_));
 sg13g2_buf_2 fanout1113 (.A(net1114),
    .X(net1113));
 sg13g2_buf_1 fanout1114 (.A(net1115),
    .X(net1114));
 sg13g2_buf_2 fanout1115 (.A(net1116),
    .X(net1115));
 sg13g2_buf_4 fanout1116 (.X(net1116),
    .A(_2745_));
 sg13g2_buf_4 fanout1117 (.X(net1117),
    .A(_2728_));
 sg13g2_buf_4 fanout1118 (.X(net1118),
    .A(_2726_));
 sg13g2_buf_2 fanout1119 (.A(net1121),
    .X(net1119));
 sg13g2_buf_1 fanout1120 (.A(net1121),
    .X(net1120));
 sg13g2_buf_2 fanout1121 (.A(_1489_),
    .X(net1121));
 sg13g2_buf_2 fanout1122 (.A(_1481_),
    .X(net1122));
 sg13g2_buf_2 fanout1123 (.A(_1481_),
    .X(net1123));
 sg13g2_buf_2 fanout1124 (.A(net1125),
    .X(net1124));
 sg13g2_buf_2 fanout1125 (.A(_0874_),
    .X(net1125));
 sg13g2_buf_2 fanout1126 (.A(_0856_),
    .X(net1126));
 sg13g2_buf_2 fanout1127 (.A(_0856_),
    .X(net1127));
 sg13g2_buf_2 fanout1128 (.A(net1131),
    .X(net1128));
 sg13g2_buf_4 fanout1129 (.X(net1129),
    .A(net1131));
 sg13g2_buf_1 fanout1130 (.A(net1131),
    .X(net1130));
 sg13g2_buf_2 fanout1131 (.A(_0844_),
    .X(net1131));
 sg13g2_buf_2 fanout1132 (.A(net1135),
    .X(net1132));
 sg13g2_buf_2 fanout1133 (.A(net1135),
    .X(net1133));
 sg13g2_buf_1 fanout1134 (.A(net1135),
    .X(net1134));
 sg13g2_buf_2 fanout1135 (.A(_0779_),
    .X(net1135));
 sg13g2_buf_2 fanout1136 (.A(net1138),
    .X(net1136));
 sg13g2_buf_1 fanout1137 (.A(net1138),
    .X(net1137));
 sg13g2_buf_2 fanout1138 (.A(_0769_),
    .X(net1138));
 sg13g2_buf_2 fanout1139 (.A(net1142),
    .X(net1139));
 sg13g2_buf_2 fanout1140 (.A(net1141),
    .X(net1140));
 sg13g2_buf_1 fanout1141 (.A(net1142),
    .X(net1141));
 sg13g2_buf_1 fanout1142 (.A(_0756_),
    .X(net1142));
 sg13g2_buf_2 fanout1143 (.A(net1145),
    .X(net1143));
 sg13g2_buf_2 fanout1144 (.A(net1145),
    .X(net1144));
 sg13g2_buf_4 fanout1145 (.X(net1145),
    .A(_2725_));
 sg13g2_buf_4 fanout1146 (.X(net1146),
    .A(net1148));
 sg13g2_buf_4 fanout1147 (.X(net1147),
    .A(net1148));
 sg13g2_buf_4 fanout1148 (.X(net1148),
    .A(_2525_));
 sg13g2_buf_4 fanout1149 (.X(net1149),
    .A(_2028_));
 sg13g2_buf_4 fanout1150 (.X(net1150),
    .A(net1151));
 sg13g2_buf_4 fanout1151 (.X(net1151),
    .A(_2027_));
 sg13g2_buf_2 fanout1152 (.A(_0916_),
    .X(net1152));
 sg13g2_buf_4 fanout1153 (.X(net1153),
    .A(_2733_));
 sg13g2_buf_4 fanout1154 (.X(net1154),
    .A(_2690_));
 sg13g2_buf_2 fanout1155 (.A(net1156),
    .X(net1155));
 sg13g2_buf_4 fanout1156 (.X(net1156),
    .A(_2684_));
 sg13g2_buf_2 fanout1157 (.A(net1158),
    .X(net1157));
 sg13g2_buf_2 fanout1158 (.A(_2684_),
    .X(net1158));
 sg13g2_buf_2 fanout1159 (.A(net1162),
    .X(net1159));
 sg13g2_buf_2 fanout1160 (.A(net1161),
    .X(net1160));
 sg13g2_buf_2 fanout1161 (.A(net1162),
    .X(net1161));
 sg13g2_buf_4 fanout1162 (.X(net1162),
    .A(_2683_));
 sg13g2_buf_2 fanout1163 (.A(net1165),
    .X(net1163));
 sg13g2_buf_2 fanout1164 (.A(net1165),
    .X(net1164));
 sg13g2_buf_2 fanout1165 (.A(_2030_),
    .X(net1165));
 sg13g2_buf_2 fanout1166 (.A(net1167),
    .X(net1166));
 sg13g2_buf_2 fanout1167 (.A(_0992_),
    .X(net1167));
 sg13g2_buf_2 fanout1168 (.A(_0992_),
    .X(net1168));
 sg13g2_buf_4 fanout1169 (.X(net1169),
    .A(_0981_));
 sg13g2_buf_2 fanout1170 (.A(_0981_),
    .X(net1170));
 sg13g2_buf_2 fanout1171 (.A(net1172),
    .X(net1171));
 sg13g2_buf_2 fanout1172 (.A(_0959_),
    .X(net1172));
 sg13g2_buf_4 fanout1173 (.X(net1173),
    .A(_2756_));
 sg13g2_buf_2 fanout1174 (.A(net1175),
    .X(net1174));
 sg13g2_buf_4 fanout1175 (.X(net1175),
    .A(_2686_));
 sg13g2_buf_4 fanout1176 (.X(net1176),
    .A(_2026_));
 sg13g2_buf_4 fanout1177 (.X(net1177),
    .A(_2026_));
 sg13g2_buf_2 fanout1178 (.A(net1179),
    .X(net1178));
 sg13g2_buf_1 fanout1179 (.A(net1180),
    .X(net1179));
 sg13g2_buf_2 fanout1180 (.A(_1630_),
    .X(net1180));
 sg13g2_buf_4 fanout1181 (.X(net1181),
    .A(_1623_));
 sg13g2_buf_1 fanout1182 (.A(_1623_),
    .X(net1182));
 sg13g2_buf_2 fanout1183 (.A(net1186),
    .X(net1183));
 sg13g2_buf_2 fanout1184 (.A(net1185),
    .X(net1184));
 sg13g2_buf_1 fanout1185 (.A(net1186),
    .X(net1185));
 sg13g2_buf_2 fanout1186 (.A(_1622_),
    .X(net1186));
 sg13g2_buf_4 fanout1187 (.X(net1187),
    .A(_1598_));
 sg13g2_buf_2 fanout1188 (.A(_1598_),
    .X(net1188));
 sg13g2_buf_2 fanout1189 (.A(net1190),
    .X(net1189));
 sg13g2_buf_2 fanout1190 (.A(_1598_),
    .X(net1190));
 sg13g2_buf_2 fanout1191 (.A(net1192),
    .X(net1191));
 sg13g2_buf_2 fanout1192 (.A(net1194),
    .X(net1192));
 sg13g2_buf_2 fanout1193 (.A(net1194),
    .X(net1193));
 sg13g2_buf_2 fanout1194 (.A(_1597_),
    .X(net1194));
 sg13g2_buf_4 fanout1195 (.X(net1195),
    .A(_1591_));
 sg13g2_buf_2 fanout1196 (.A(_1590_),
    .X(net1196));
 sg13g2_buf_2 fanout1197 (.A(net1198),
    .X(net1197));
 sg13g2_buf_4 fanout1198 (.X(net1198),
    .A(_1586_));
 sg13g2_buf_4 fanout1199 (.X(net1199),
    .A(_1585_));
 sg13g2_buf_2 fanout1200 (.A(net1201),
    .X(net1200));
 sg13g2_buf_2 fanout1201 (.A(_1581_),
    .X(net1201));
 sg13g2_buf_4 fanout1202 (.X(net1202),
    .A(_1581_));
 sg13g2_buf_2 fanout1203 (.A(_1580_),
    .X(net1203));
 sg13g2_buf_2 fanout1204 (.A(_1580_),
    .X(net1204));
 sg13g2_buf_2 fanout1205 (.A(net1207),
    .X(net1205));
 sg13g2_buf_1 fanout1206 (.A(net1207),
    .X(net1206));
 sg13g2_buf_2 fanout1207 (.A(net1208),
    .X(net1207));
 sg13g2_buf_2 fanout1208 (.A(_1576_),
    .X(net1208));
 sg13g2_buf_2 fanout1209 (.A(net1210),
    .X(net1209));
 sg13g2_buf_2 fanout1210 (.A(net1212),
    .X(net1210));
 sg13g2_buf_2 fanout1211 (.A(net1212),
    .X(net1211));
 sg13g2_buf_2 fanout1212 (.A(_1575_),
    .X(net1212));
 sg13g2_buf_2 fanout1213 (.A(net1216),
    .X(net1213));
 sg13g2_buf_2 fanout1214 (.A(net1216),
    .X(net1214));
 sg13g2_buf_1 fanout1215 (.A(net1216),
    .X(net1215));
 sg13g2_buf_4 fanout1216 (.X(net1216),
    .A(_1570_));
 sg13g2_buf_4 fanout1217 (.X(net1217),
    .A(_1081_));
 sg13g2_buf_4 fanout1218 (.X(net1218),
    .A(_1064_));
 sg13g2_buf_2 fanout1219 (.A(net1220),
    .X(net1219));
 sg13g2_buf_2 fanout1220 (.A(_1049_),
    .X(net1220));
 sg13g2_buf_2 fanout1221 (.A(net1222),
    .X(net1221));
 sg13g2_buf_2 fanout1222 (.A(net1223),
    .X(net1222));
 sg13g2_buf_4 fanout1223 (.X(net1223),
    .A(_1034_));
 sg13g2_buf_2 fanout1224 (.A(_0914_),
    .X(net1224));
 sg13g2_buf_4 fanout1225 (.X(net1225),
    .A(_2688_));
 sg13g2_buf_2 fanout1226 (.A(_2688_),
    .X(net1226));
 sg13g2_buf_4 fanout1227 (.X(net1227),
    .A(_2687_));
 sg13g2_buf_2 fanout1228 (.A(net1229),
    .X(net1228));
 sg13g2_buf_4 fanout1229 (.X(net1229),
    .A(_2025_));
 sg13g2_buf_2 fanout1230 (.A(net1231),
    .X(net1230));
 sg13g2_buf_2 fanout1231 (.A(net1234),
    .X(net1231));
 sg13g2_buf_4 fanout1232 (.X(net1232),
    .A(net1234));
 sg13g2_buf_2 fanout1233 (.A(net1234),
    .X(net1233));
 sg13g2_buf_2 fanout1234 (.A(_2015_),
    .X(net1234));
 sg13g2_buf_4 fanout1235 (.X(net1235),
    .A(net1236));
 sg13g2_buf_2 fanout1236 (.A(net1237),
    .X(net1236));
 sg13g2_buf_2 fanout1237 (.A(_1565_),
    .X(net1237));
 sg13g2_buf_4 fanout1238 (.X(net1238),
    .A(_1560_));
 sg13g2_buf_2 fanout1239 (.A(_1560_),
    .X(net1239));
 sg13g2_buf_2 fanout1240 (.A(_2306_),
    .X(net1240));
 sg13g2_buf_2 fanout1241 (.A(_1558_),
    .X(net1241));
 sg13g2_buf_2 fanout1242 (.A(_0561_),
    .X(net1242));
 sg13g2_buf_4 fanout1243 (.X(net1243),
    .A(_2693_));
 sg13g2_buf_4 fanout1244 (.X(net1244),
    .A(_2692_));
 sg13g2_buf_2 fanout1245 (.A(_2692_),
    .X(net1245));
 sg13g2_buf_2 fanout1246 (.A(_2287_),
    .X(net1246));
 sg13g2_buf_2 fanout1247 (.A(_2287_),
    .X(net1247));
 sg13g2_buf_2 fanout1248 (.A(_2285_),
    .X(net1248));
 sg13g2_buf_4 fanout1249 (.X(net1249),
    .A(_2214_));
 sg13g2_buf_4 fanout1250 (.X(net1250),
    .A(net1251));
 sg13g2_buf_2 fanout1251 (.A(_2214_),
    .X(net1251));
 sg13g2_buf_4 fanout1252 (.X(net1252),
    .A(_1542_));
 sg13g2_buf_2 fanout1253 (.A(net1255),
    .X(net1253));
 sg13g2_buf_1 fanout1254 (.A(net1255),
    .X(net1254));
 sg13g2_buf_2 fanout1255 (.A(_1537_),
    .X(net1255));
 sg13g2_buf_4 fanout1256 (.X(net1256),
    .A(net1258));
 sg13g2_buf_4 fanout1257 (.X(net1257),
    .A(net1258));
 sg13g2_buf_2 fanout1258 (.A(_2662_),
    .X(net1258));
 sg13g2_buf_4 fanout1259 (.X(net1259),
    .A(_2284_));
 sg13g2_buf_1 fanout1260 (.A(_2284_),
    .X(net1260));
 sg13g2_buf_2 fanout1261 (.A(_2241_),
    .X(net1261));
 sg13g2_buf_1 fanout1262 (.A(_2241_),
    .X(net1262));
 sg13g2_buf_4 fanout1263 (.X(net1263),
    .A(_2218_));
 sg13g2_buf_2 fanout1264 (.A(net1265),
    .X(net1264));
 sg13g2_buf_2 fanout1265 (.A(net1266),
    .X(net1265));
 sg13g2_buf_2 fanout1266 (.A(_1881_),
    .X(net1266));
 sg13g2_buf_2 fanout1267 (.A(net1268),
    .X(net1267));
 sg13g2_buf_2 fanout1268 (.A(net1269),
    .X(net1268));
 sg13g2_buf_4 fanout1269 (.X(net1269),
    .A(_1866_));
 sg13g2_buf_4 fanout1270 (.X(net1270),
    .A(net1271));
 sg13g2_buf_4 fanout1271 (.X(net1271),
    .A(_1556_));
 sg13g2_buf_2 fanout1272 (.A(_1556_),
    .X(net1272));
 sg13g2_buf_4 fanout1273 (.X(net1273),
    .A(_1553_));
 sg13g2_buf_4 fanout1274 (.X(net1274),
    .A(_1548_));
 sg13g2_buf_2 fanout1275 (.A(_1548_),
    .X(net1275));
 sg13g2_buf_2 fanout1276 (.A(net1278),
    .X(net1276));
 sg13g2_buf_1 fanout1277 (.A(net1278),
    .X(net1277));
 sg13g2_buf_2 fanout1278 (.A(_1534_),
    .X(net1278));
 sg13g2_buf_4 fanout1279 (.X(net1279),
    .A(_0999_));
 sg13g2_buf_2 fanout1280 (.A(_0930_),
    .X(net1280));
 sg13g2_buf_1 fanout1281 (.A(_0930_),
    .X(net1281));
 sg13g2_buf_4 fanout1282 (.X(net1282),
    .A(_3326_));
 sg13g2_buf_2 fanout1283 (.A(_3284_),
    .X(net1283));
 sg13g2_buf_1 fanout1284 (.A(_3284_),
    .X(net1284));
 sg13g2_buf_4 fanout1285 (.X(net1285),
    .A(_1547_));
 sg13g2_buf_2 fanout1286 (.A(_1547_),
    .X(net1286));
 sg13g2_buf_4 fanout1287 (.X(net1287),
    .A(net1288));
 sg13g2_buf_4 fanout1288 (.X(net1288),
    .A(_1546_));
 sg13g2_buf_4 fanout1289 (.X(net1289),
    .A(net1292));
 sg13g2_buf_2 fanout1290 (.A(net1292),
    .X(net1290));
 sg13g2_buf_4 fanout1291 (.X(net1291),
    .A(net1292));
 sg13g2_buf_2 fanout1292 (.A(_1545_),
    .X(net1292));
 sg13g2_buf_4 fanout1293 (.X(net1293),
    .A(net1294));
 sg13g2_buf_2 fanout1294 (.A(net1295),
    .X(net1294));
 sg13g2_buf_2 fanout1295 (.A(_1531_),
    .X(net1295));
 sg13g2_buf_2 fanout1296 (.A(net1297),
    .X(net1296));
 sg13g2_buf_2 fanout1297 (.A(net1298),
    .X(net1297));
 sg13g2_buf_2 fanout1298 (.A(net1299),
    .X(net1298));
 sg13g2_buf_2 fanout1299 (.A(_1531_),
    .X(net1299));
 sg13g2_buf_4 fanout1300 (.X(net1300),
    .A(_0732_));
 sg13g2_buf_4 fanout1301 (.X(net1301),
    .A(_0657_));
 sg13g2_buf_2 fanout1302 (.A(net1303),
    .X(net1302));
 sg13g2_buf_2 fanout1303 (.A(_2532_),
    .X(net1303));
 sg13g2_buf_4 fanout1304 (.X(net1304),
    .A(net1306));
 sg13g2_buf_1 fanout1305 (.A(net1306),
    .X(net1305));
 sg13g2_buf_2 fanout1306 (.A(net1307),
    .X(net1306));
 sg13g2_buf_2 fanout1307 (.A(net1313),
    .X(net1307));
 sg13g2_buf_2 fanout1308 (.A(net1311),
    .X(net1308));
 sg13g2_buf_2 fanout1309 (.A(net1310),
    .X(net1309));
 sg13g2_buf_2 fanout1310 (.A(net1311),
    .X(net1310));
 sg13g2_buf_2 fanout1311 (.A(net1313),
    .X(net1311));
 sg13g2_buf_2 fanout1312 (.A(net1313),
    .X(net1312));
 sg13g2_buf_2 fanout1313 (.A(_1532_),
    .X(net1313));
 sg13g2_buf_4 fanout1314 (.X(net1314),
    .A(_1017_));
 sg13g2_buf_2 fanout1315 (.A(_1017_),
    .X(net1315));
 sg13g2_buf_2 fanout1316 (.A(net1317),
    .X(net1316));
 sg13g2_buf_4 fanout1317 (.X(net1317),
    .A(_0676_));
 sg13g2_buf_2 fanout1318 (.A(_0653_),
    .X(net1318));
 sg13g2_buf_2 fanout1319 (.A(_0639_),
    .X(net1319));
 sg13g2_buf_2 fanout1320 (.A(net1321),
    .X(net1320));
 sg13g2_buf_2 fanout1321 (.A(_0625_),
    .X(net1321));
 sg13g2_buf_4 fanout1322 (.X(net1322),
    .A(_0623_));
 sg13g2_buf_1 fanout1323 (.A(_0623_),
    .X(net1323));
 sg13g2_buf_2 fanout1324 (.A(net1325),
    .X(net1324));
 sg13g2_buf_2 fanout1325 (.A(_0611_),
    .X(net1325));
 sg13g2_buf_2 fanout1326 (.A(net1327),
    .X(net1326));
 sg13g2_buf_2 fanout1327 (.A(_0580_),
    .X(net1327));
 sg13g2_buf_2 fanout1328 (.A(_3324_),
    .X(net1328));
 sg13g2_buf_4 fanout1329 (.X(net1329),
    .A(_0624_));
 sg13g2_buf_2 fanout1330 (.A(_0624_),
    .X(net1330));
 sg13g2_buf_4 fanout1331 (.X(net1331),
    .A(net1333));
 sg13g2_buf_2 fanout1332 (.A(net1333),
    .X(net1332));
 sg13g2_buf_2 fanout1333 (.A(_0614_),
    .X(net1333));
 sg13g2_buf_4 fanout1334 (.X(net1334),
    .A(_0612_));
 sg13g2_buf_2 fanout1335 (.A(_0612_),
    .X(net1335));
 sg13g2_buf_4 fanout1336 (.X(net1336),
    .A(_0600_));
 sg13g2_buf_2 fanout1337 (.A(_0600_),
    .X(net1337));
 sg13g2_buf_4 fanout1338 (.X(net1338),
    .A(net1339));
 sg13g2_buf_2 fanout1339 (.A(_0594_),
    .X(net1339));
 sg13g2_buf_4 fanout1340 (.X(net1340),
    .A(_0589_));
 sg13g2_buf_2 fanout1341 (.A(_0589_),
    .X(net1341));
 sg13g2_buf_4 fanout1342 (.X(net1342),
    .A(_0587_));
 sg13g2_buf_2 fanout1343 (.A(_0586_),
    .X(net1343));
 sg13g2_buf_4 fanout1344 (.X(net1344),
    .A(_3211_));
 sg13g2_buf_2 fanout1345 (.A(_3211_),
    .X(net1345));
 sg13g2_buf_4 fanout1346 (.X(net1346),
    .A(_3189_));
 sg13g2_buf_4 fanout1347 (.X(net1347),
    .A(_3187_));
 sg13g2_buf_4 fanout1348 (.X(net1348),
    .A(_3187_));
 sg13g2_buf_4 fanout1349 (.X(net1349),
    .A(_3185_));
 sg13g2_buf_2 fanout1350 (.A(_3154_),
    .X(net1350));
 sg13g2_buf_2 fanout1351 (.A(_3154_),
    .X(net1351));
 sg13g2_buf_2 fanout1352 (.A(net1354),
    .X(net1352));
 sg13g2_buf_2 fanout1353 (.A(net1354),
    .X(net1353));
 sg13g2_buf_2 fanout1354 (.A(net691),
    .X(net1354));
 sg13g2_buf_2 fanout1355 (.A(net1356),
    .X(net1355));
 sg13g2_buf_2 fanout1356 (.A(net674),
    .X(net1356));
 sg13g2_buf_2 fanout1357 (.A(net1359),
    .X(net1357));
 sg13g2_buf_2 fanout1358 (.A(net1359),
    .X(net1358));
 sg13g2_buf_2 fanout1359 (.A(net1360),
    .X(net1359));
 sg13g2_buf_1 fanout1360 (.A(net1362),
    .X(net1360));
 sg13g2_buf_4 fanout1361 (.X(net1361),
    .A(net1362));
 sg13g2_buf_4 fanout1362 (.X(net1362),
    .A(\dtop.enable ));
 sg13g2_buf_4 fanout1363 (.X(net1363),
    .A(\dtop.vtop.pipeline.nstep_zg[1] ));
 sg13g2_buf_2 fanout1364 (.A(net681),
    .X(net1364));
 sg13g2_buf_4 fanout1365 (.X(net1365),
    .A(net1366));
 sg13g2_buf_2 fanout1366 (.A(net701),
    .X(net1366));
 sg13g2_buf_2 fanout1367 (.A(net1368),
    .X(net1367));
 sg13g2_buf_2 fanout1368 (.A(_0086_),
    .X(net1368));
 sg13g2_buf_4 fanout1369 (.X(net1369),
    .A(\dtop.player_inst.program_addr[6] ));
 sg13g2_buf_2 fanout1370 (.A(\dtop.player_inst.program_addr[6] ),
    .X(net1370));
 sg13g2_buf_4 fanout1371 (.X(net1371),
    .A(net1373));
 sg13g2_buf_1 fanout1372 (.A(net1373),
    .X(net1372));
 sg13g2_buf_2 fanout1373 (.A(net683),
    .X(net1373));
 sg13g2_buf_4 fanout1374 (.X(net1374),
    .A(net1375));
 sg13g2_buf_2 fanout1375 (.A(net1376),
    .X(net1375));
 sg13g2_buf_2 fanout1376 (.A(net672),
    .X(net1376));
 sg13g2_buf_4 fanout1377 (.X(net1377),
    .A(net1378));
 sg13g2_buf_2 fanout1378 (.A(net1379),
    .X(net1378));
 sg13g2_buf_2 fanout1379 (.A(net659),
    .X(net1379));
 sg13g2_buf_4 fanout1380 (.X(net1380),
    .A(net1381));
 sg13g2_buf_2 fanout1381 (.A(net1382),
    .X(net1381));
 sg13g2_buf_4 fanout1382 (.X(net1382),
    .A(net705));
 sg13g2_buf_2 fanout1383 (.A(net1387),
    .X(net1383));
 sg13g2_buf_2 fanout1384 (.A(net1386),
    .X(net1384));
 sg13g2_buf_1 fanout1385 (.A(net1386),
    .X(net1385));
 sg13g2_buf_4 fanout1386 (.X(net1386),
    .A(net1387));
 sg13g2_buf_1 fanout1387 (.A(net1388),
    .X(net1387));
 sg13g2_buf_4 fanout1388 (.X(net1388),
    .A(net710));
 sg13g2_buf_2 fanout1389 (.A(net1391),
    .X(net1389));
 sg13g2_buf_2 fanout1390 (.A(net1391),
    .X(net1390));
 sg13g2_buf_2 fanout1391 (.A(net1392),
    .X(net1391));
 sg13g2_buf_2 fanout1392 (.A(net677),
    .X(net1392));
 sg13g2_buf_4 fanout1393 (.X(net1393),
    .A(net706));
 sg13g2_buf_2 fanout1394 (.A(_0088_),
    .X(net1394));
 sg13g2_buf_2 fanout1395 (.A(\dtop.detune_counter[16] ),
    .X(net1395));
 sg13g2_buf_2 fanout1396 (.A(net583),
    .X(net1396));
 sg13g2_buf_2 fanout1397 (.A(net568),
    .X(net1397));
 sg13g2_buf_4 fanout1398 (.X(net1398),
    .A(\dtop.detune_counter[12] ));
 sg13g2_buf_4 fanout1399 (.X(net1399),
    .A(net1400));
 sg13g2_buf_2 fanout1400 (.A(\dtop.detune_counter[11] ),
    .X(net1400));
 sg13g2_buf_4 fanout1401 (.X(net1401),
    .A(\dtop.detune_counter[10] ));
 sg13g2_buf_4 fanout1402 (.X(net1402),
    .A(net571));
 sg13g2_buf_4 fanout1403 (.X(net1403),
    .A(\dtop.detune_counter[8] ));
 sg13g2_buf_2 fanout1404 (.A(net666),
    .X(net1404));
 sg13g2_buf_4 fanout1405 (.X(net1405),
    .A(net687));
 sg13g2_buf_4 fanout1406 (.X(net1406),
    .A(net1407));
 sg13g2_buf_4 fanout1407 (.X(net1407),
    .A(\dtop.player_inst.synth.alu.acc[10] ));
 sg13g2_buf_4 fanout1408 (.X(net1408),
    .A(net693));
 sg13g2_buf_4 fanout1409 (.X(net1409),
    .A(\dtop.player_inst.synth.alu.acc[6] ));
 sg13g2_buf_4 fanout1410 (.X(net1410),
    .A(net697));
 sg13g2_buf_4 fanout1411 (.X(net1411),
    .A(\dtop.player_inst.synth.alu.acc[3] ));
 sg13g2_buf_4 fanout1412 (.X(net1412),
    .A(net702));
 sg13g2_buf_4 fanout1413 (.X(net1413),
    .A(net708));
 sg13g2_buf_4 fanout1414 (.X(net1414),
    .A(net694));
 sg13g2_buf_4 fanout1415 (.X(net1415),
    .A(net685));
 sg13g2_buf_2 fanout1416 (.A(net1417),
    .X(net1416));
 sg13g2_buf_1 fanout1417 (.A(net1418),
    .X(net1417));
 sg13g2_buf_4 fanout1418 (.X(net1418),
    .A(net680));
 sg13g2_buf_2 fanout1419 (.A(net1422),
    .X(net1419));
 sg13g2_buf_2 fanout1420 (.A(net1421),
    .X(net1420));
 sg13g2_buf_2 fanout1421 (.A(net1422),
    .X(net1421));
 sg13g2_buf_2 fanout1422 (.A(net1423),
    .X(net1422));
 sg13g2_buf_2 fanout1423 (.A(net1424),
    .X(net1423));
 sg13g2_buf_2 fanout1424 (.A(net603),
    .X(net1424));
 sg13g2_buf_4 fanout1425 (.X(net1425),
    .A(\dtop.oct_counter[6] ));
 sg13g2_buf_4 fanout1426 (.X(net1426),
    .A(net703));
 sg13g2_buf_2 fanout1427 (.A(net1428),
    .X(net1427));
 sg13g2_buf_1 fanout1428 (.A(net1440),
    .X(net1428));
 sg13g2_buf_2 fanout1429 (.A(net1440),
    .X(net1429));
 sg13g2_buf_4 fanout1430 (.X(net1430),
    .A(net1440));
 sg13g2_buf_2 fanout1431 (.A(net1439),
    .X(net1431));
 sg13g2_buf_2 fanout1432 (.A(net1439),
    .X(net1432));
 sg13g2_buf_2 fanout1433 (.A(net1439),
    .X(net1433));
 sg13g2_buf_2 fanout1434 (.A(net1436),
    .X(net1434));
 sg13g2_buf_2 fanout1435 (.A(net1436),
    .X(net1435));
 sg13g2_buf_2 fanout1436 (.A(net1439),
    .X(net1436));
 sg13g2_buf_2 fanout1437 (.A(net1438),
    .X(net1437));
 sg13g2_buf_2 fanout1438 (.A(net1439),
    .X(net1438));
 sg13g2_buf_2 fanout1439 (.A(net1440),
    .X(net1439));
 sg13g2_buf_2 fanout1440 (.A(rst_n_reg),
    .X(net1440));
 sg13g2_buf_2 fanout1441 (.A(net1442),
    .X(net1441));
 sg13g2_buf_1 fanout1442 (.A(\dtop.oct_counter[2] ),
    .X(net1442));
 sg13g2_buf_2 fanout1443 (.A(net1444),
    .X(net1443));
 sg13g2_buf_1 fanout1444 (.A(\dtop.oct_counter[1] ),
    .X(net1444));
 sg13g2_buf_4 fanout1445 (.X(net1445),
    .A(net1446));
 sg13g2_buf_4 fanout1446 (.X(net1446),
    .A(\dtop.oct_counter[0] ));
 sg13g2_buf_4 fanout1447 (.X(net1447),
    .A(\dtop.ext_control[5] ));
 sg13g2_buf_4 fanout1448 (.X(net1448),
    .A(\dtop.ext_control[4] ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_tiehi _7284__10 (.L_HI(net10));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_8 clkload7 (.A(clknet_leaf_45_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_46_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_7_clk));
 sg13g2_inv_2 clkload10 (.A(clknet_leaf_14_clk));
 sg13g2_inv_8 clkload11 (.A(clknet_leaf_15_clk));
 sg13g2_inv_2 clkload12 (.A(clknet_leaf_9_clk));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_10_clk));
 sg13g2_inv_8 clkload14 (.A(clknet_leaf_16_clk));
 sg13g2_inv_1 clkload15 (.A(clknet_leaf_8_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_20_clk));
 sg13g2_inv_4 clkload17 (.A(clknet_leaf_21_clk));
 sg13g2_inv_4 clkload18 (.A(clknet_leaf_32_clk));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_33_clk));
 sg13g2_inv_4 clkload20 (.A(clknet_leaf_34_clk));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_35_clk));
 sg13g2_inv_4 clkload22 (.A(clknet_leaf_18_clk));
 sg13g2_inv_1 clkload23 (.A(clknet_leaf_19_clk));
 sg13g2_inv_4 clkload24 (.A(clknet_leaf_27_clk));
 sg13g2_inv_1 clkload25 (.A(clknet_leaf_29_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\dtop.vtop.pipeline.next_nstep_counter[0] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0374_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold3 (.A(\dtop.vsync ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold4 (.A(_1957_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0252_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold6 (.A(\dtop.player_inst.synth.alu.registers[4][10] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0138_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold8 (.A(\dtop.vtop.dphases[0][1] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold9 (.A(\dtop.vtop.dphases[0][5] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold10 (.A(\dtop.vtop.dphases[0][4] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold11 (.A(\dtop.vtop.dphases[0][3] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold12 (.A(\dtop.player_inst.synth.alu.registers[4][6] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0134_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold14 (.A(\dtop.vtop.dphases[0][7] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold15 (.A(\dtop.vtop.dphases[0][2] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold16 (.A(\dtop.vtop.dphases[0][8] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold17 (.A(\dtop.player_inst.synth.alu.registers[4][8] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0136_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold19 (.A(_3353_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold20 (.A(\dtop.vtop.dphases[0][0] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold21 (.A(\dtop.player_inst.synth.alu.registers[4][9] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0137_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold23 (.A(\dtop.vtop.dphases[0][6] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold24 (.A(\dtop.vtop.dphases[1][0] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold25 (.A(\dtop.player_inst.synth.alu.registers[4][7] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0135_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold27 (.A(\dtop.vtop.dphases[0][10] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0227_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold29 (.A(\dtop.vtop.dphases[1][5] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold30 (.A(\dtop.vtop.pipeline.phases[0][10] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold31 (.A(\dtop.vtop.dphases[1][1] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold32 (.A(\dtop.player_inst.synth.alu.registers[2][7] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0146_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold34 (.A(\dtop.player_inst.synth.alu.registers[3][6] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0201_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold36 (.A(\dtop.vtop.dphases[1][4] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold37 (.A(\dtop.player_inst.synth.alu.registers[2][4] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0143_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold39 (.A(\dtop.player_inst.synth.alu.registers[3][0] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold40 (.A(\dtop.vtop.dphases[1][9] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold41 (.A(\dtop.vtop.dphases[2][4] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold42 (.A(\dtop.player_inst.synth.alu.registers[3][7] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0202_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold44 (.A(\dtop.vtop.dphases[2][8] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold45 (.A(\dtop.vtop.dphases[2][5] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold46 (.A(\dtop.vtop.dphases[2][2] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold47 (.A(\dtop.vtop.dphases[2][9] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold48 (.A(\dtop.vtop.pipeline.phases[0][3] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold49 (.A(\dtop.vtop.pipeline.phases[0][13] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold50 (.A(\dtop.vtop.dphases[1][8] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold51 (.A(\dtop.player_inst.synth.alu.registers[5][0] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0188_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold53 (.A(\dtop.vtop.pipeline.phases[0][0] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0379_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold55 (.A(\dtop.vtop.pipeline.phases[0][11] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold56 (.A(\dtop.vtop.dphases[2][1] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold57 (.A(\dtop.vtop.dphases[0][9] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0226_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold59 (.A(\dtop.vtop.pipeline.cosappr_acc[1] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0351_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold61 (.A(\dtop.vtop.pipeline.phases[0][12] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold62 (.A(\dtop.vtop.dphases[2][6] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold63 (.A(\dtop.player_inst.synth.alu.registers[1][6] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0153_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold65 (.A(\dtop.vtop.dphases[2][7] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold66 (.A(\dtop.player_inst.synth.alu.registers[5][6] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold67 (.A(\dtop.vtop.pipeline.phases[0][14] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold68 (.A(\dtop.player_inst.synth.alu.registers[2][6] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold69 (.A(\dtop.player_inst.synth.alu.registers[2][1] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0140_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold71 (.A(\dtop.vtop.dphases[1][7] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold72 (.A(\dtop.vtop.pipeline.phases[0][2] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold73 (.A(\dtop.vtop.pipeline.phases[0][15] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold74 (.A(\dtop.player_inst.synth.alu.registers[3][4] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0199_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold76 (.A(\dtop.vtop.pipeline.phases[0][1] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold77 (.A(\dtop.vtop.pipeline.phases[0][6] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold78 (.A(\dtop.vtop.dphases[1][2] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold79 (.A(\dtop.player_inst.synth.alu.registers[2][0] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0139_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold81 (.A(\dtop.player_inst.synth.alu.registers[3][3] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold82 (.A(\dtop.vtop.dphases[1][10] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0238_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold84 (.A(\dtop.vtop.pipeline.phases[0][5] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold85 (.A(\dtop.player_inst.synth.alu.registers[5][4] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0192_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold87 (.A(\dtop.player_inst.synth.alu.registers[5][3] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0191_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold89 (.A(\dtop.player_inst.synth.alu.registers[1][4] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0151_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold91 (.A(\dtop.player_inst.synth.alu.registers[1][1] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0148_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold93 (.A(\dtop.player_inst.synth.alu.registers[3][1] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0196_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold95 (.A(\dtop.vtop.pipeline.phases[0][8] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold96 (.A(\dtop.player_inst.synth.alu.registers[2][3] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold97 (.A(\dtop.player_inst.synth.alu.registers[2][2] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0141_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold99 (.A(\dtop.vtop.pipeline.phases[0][7] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold100 (.A(\dtop.player_inst.synth.alu.registers[2][5] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold101 (.A(\dtop.vtop.pipeline.zg_acc[6] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold102 (.A(\dtop.vtop.pipeline.phases[0][9] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold103 (.A(\dtop.player_inst.synth.alu.registers[1][2] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0149_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold105 (.A(\dtop.vtop.dphases[1][6] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold106 (.A(\dtop.player_inst.synth.alu.registers[1][3] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold107 (.A(\dtop.vtop.pipeline.cosappr_acc[7] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold108 (.A(\dtop.vtop.pipeline.zg_acc[7] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold109 (.A(\dtop.vtop.pipeline.z[14] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold110 (.A(\dtop.player_inst.synth.alu.registers[5][1] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold111 (.A(\dtop.player_inst.synth.alu.registers[3][2] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold112 (.A(\dtop.vtop.dphases[2][0] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold113 (.A(\dtop.player_inst.synth.alu.registers[5][5] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold114 (.A(\dtop.vtop.pipeline.phases[2][11] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold115 (.A(\dtop.vtop.pipeline.phases[0][4] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold116 (.A(\dtop.vtop.dphases[2][3] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold117 (.A(\dtop.player_inst.synth.alu.registers[1][8] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0155_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold119 (.A(\dtop.player_inst.synth.alu.registers[1][0] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold120 (.A(\dtop.player_inst.synth.alu.registers[5][2] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0190_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold122 (.A(\dtop.player_inst.synth.alu.oct_en ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold123 (.A(\dtop.out_sample[0] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0169_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold125 (.A(\dtop.player_inst.synth.alu.registers[1][10] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0157_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold127 (.A(\dtop.player_inst.synth.alu.registers[1][7] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0154_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold129 (.A(\dtop.vtop.pipeline.cosappr_acc[3] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold130 (.A(\dtop.player_inst.synth.alu.acc[10] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold131 (.A(\dtop.vtop.pipeline.phases[1][0] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0301_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold133 (.A(\dtop.vtop.pipeline.cosappr_acc[4] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold134 (.A(\dtop.vtop.pipeline.phases[1][13] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold135 (.A(\dtop.vtop.pipeline.cosappr_acc[8] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold136 (.A(\dtop.vtop.pipeline.phases[2][14] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold137 (.A(\dtop.vtop.pipeline.phases[2][6] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold138 (.A(\dtop.vtop.pipeline.phases[1][12] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold139 (.A(\dtop.vtop.pipeline.cosappr_acc[6] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold140 (.A(\dtop.vtop.pipeline.phases[2][2] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold141 (.A(\dtop.vtop.pipeline.phases[2][7] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold142 (.A(\dtop.vtop.pipeline.phases[2][10] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold143 (.A(\dtop.vtop.pipeline.cosappr_acc[5] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold144 (.A(\dtop.vtop.pipeline.phases[1][1] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold145 (.A(\dtop.vtop.logo_d[1] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold146 (.A(\dtop.player_inst.synth.alu.registers[4][4] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0132_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold148 (.A(\dtop.vtop.pipeline.phases[1][15] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold149 (.A(\dtop.vtop.pipeline.phases[1][9] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold150 (.A(\dtop.vtop.pipeline.phases[1][4] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold151 (.A(\dtop.vtop.pipeline.phases[1][11] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold152 (.A(\dtop.ext_control[4] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0103_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold154 (.A(\dtop.player_inst.synth.alu.registers[4][0] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0128_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold156 (.A(\dtop.vtop.pipeline.phases[1][8] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold157 (.A(\dtop.vtop.pipeline.phases[2][3] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold158 (.A(\dtop.vtop.dphases[1][3] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold159 (.A(\dtop.vtop.pipeline.phases[1][10] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold160 (.A(\dtop.vtop.pipeline.phases[2][1] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold161 (.A(\dtop.vtop.pipeline.phases[1][3] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold162 (.A(\dtop.vtop.pipeline.phases[1][7] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold163 (.A(\dtop.player_inst.synth.alu.registers[1][9] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0156_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold165 (.A(\dtop.vtop.pipeline.phases[1][14] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold166 (.A(\dtop.vtop.pipeline.phases[2][13] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold167 (.A(\dtop.vtop.pipeline.zg[0] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold168 (.A(\dtop.out_sample[3] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold169 (.A(\dtop.vtop.pipeline.phases[2][8] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold170 (.A(\dtop.vtop.pipeline.z[0] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold171 (.A(_2098_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0286_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold173 (.A(\dtop.out_sample[2] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold174 (.A(\dtop.vtop.pipeline.zg_acc[9] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold175 (.A(\dtop.vtop.pipeline.nstep_counter[4] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0378_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold177 (.A(\dtop.vtop.pipeline.cosappr_acc[2] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold178 (.A(\dtop.vtop.pipeline.phases[2][4] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold179 (.A(\dtop.vtop.pipeline.phases[2][0] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0317_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold181 (.A(\dtop.out_sample[4] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold182 (.A(\dtop.player_inst.synth.alu.registers[4][2] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0130_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold184 (.A(\dtop.out_sample[6] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold185 (.A(\dtop.vtop.dphases[2][10] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0249_),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold187 (.A(\dtop.vtop.pipeline.phases[2][12] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold188 (.A(\dtop.player_inst.synth.alu.registers[1][5] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold189 (.A(\dtop.vtop.pipeline.phases[1][6] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold190 (.A(\dtop.vtop.pipeline.phases[1][2] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold191 (.A(\dtop.out_sample[5] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold192 (.A(\dtop.vtop.pipeline.phases[2][15] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold193 (.A(\dtop.vtop.pipeline.phases[2][9] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold194 (.A(\dtop.vtop.pipeline.phases[1][5] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold195 (.A(\dtop.player_inst.synth.alu.registers[3][5] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold196 (.A(\dtop.vtop.pipeline.zg_acc[8] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold197 (.A(\dtop.player_inst.synth.alu.registers[4][1] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0129_),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold199 (.A(\dtop.vtop.pipeline.dz[7] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold200 (.A(\dtop.vtop.pipeline.zg[1] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold201 (.A(\dtop.out_sample[1] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0170_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold203 (.A(\dtop.vtop.pipeline.dz[3] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0280_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold205 (.A(\dtop.vtop.pipeline.phases[2][5] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold206 (.A(\dtop.player_inst.synth.alu.registers[4][5] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold207 (.A(\uio_out0b[5] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0433_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0108_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold210 (.A(\dtop.vtop.pipeline.cosappr_acc[0] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold211 (.A(\dtop.vtop.color[11] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold212 (.A(\dtop.vtop.pipeline.neg_t[8] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0275_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold214 (.A(\dtop.player_inst.synth.alu.registers[4][3] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0131_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold216 (.A(\dtop.vtop.pipeline.zg[2] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold217 (.A(\dtop.player_inst.synth.alu.registers[0][10] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold218 (.A(uo_out[7]),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0116_),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold220 (.A(\dtop.vtop.pipeline.nstep_counter[3] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold221 (.A(_2660_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0377_),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold223 (.A(\dtop.player_inst.synth.alu.registers[0][8] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0166_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold225 (.A(\dtop.player_inst.synth.alu.registers[0][1] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0159_),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold227 (.A(\dtop.vtop.color[8] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold228 (.A(\dtop.vtop.pipeline.neg_t[2] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold229 (.A(\dtop.player_inst.synth.alu.registers[0][0] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0158_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold231 (.A(\dtop.player_inst.synth.alu.registers[0][2] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold232 (.A(\dtop.player_inst.synth.alu.registers[0][6] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0164_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold234 (.A(\dtop.vtop.pipeline.zg_acc[5] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold235 (.A(\dtop.vtop.pipeline.wave_index[0] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold236 (.A(_2643_),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold237 (.A(\dtop.vtop.pipeline.nstep_counter[1] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold238 (.A(_2658_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0375_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold240 (.A(\dtop.vtop.pipeline.neg_t[6] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold241 (.A(\dtop.vtop.force_sat0 ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold242 (.A(\dtop.vtop.pipeline.dz[2] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold243 (.A(\dtop.player_inst.synth.alu.registers[0][7] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0165_),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold245 (.A(\dtop.vtop.color[10] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold246 (.A(uo_out[6]),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold247 (.A(uio_out[4]),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0107_),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold249 (.A(\dtop.vtop.pipeline.neg_t[4] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold250 (.A(\dtop.vtop.pipeline.neg_t[1] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold251 (.A(\dtop.detune_counter[13] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0213_),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold253 (.A(\dtop.vtop.color[6] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold254 (.A(\dtop.detune_counter[9] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold255 (.A(_1522_),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold256 (.A(\dtop.vtop.pipeline.zg_acc[1] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold257 (.A(\dtop.oct_counter[2] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0102_),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold259 (.A(\dtop.vtop.pipeline.dz[6] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold260 (.A(\dtop.vtop.pipeline.neg_t[9] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold261 (.A(_0276_),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold262 (.A(\dtop.vtop.pipeline.z[11] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold263 (.A(\dtop.vtop.color[9] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold264 (.A(uio_out[7]),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold265 (.A(_0118_),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold266 (.A(\dtop.detune_counter[15] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold267 (.A(\dtop.player_inst.synth.alu.registers[0][5] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold268 (.A(\dtop.player_inst.synth.alu.registers[0][3] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold269 (.A(\dtop.player_inst.synth.alu.registers[0][9] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0167_),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold271 (.A(\dtop.player_inst.synth.alu.registers[0][4] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold272 (.A(_0162_),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold273 (.A(\dtop.vtop.pipeline.zg_acc[2] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold274 (.A(uo_out[2]),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0111_),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold276 (.A(\dtop.vtop.pipeline.nstep_counter[2] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0376_),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold278 (.A(\dtop.vtop.pipeline.dz[8] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold279 (.A(\dtop.oct_counter[6] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0569_),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold281 (.A(\dtop.vtop.color[7] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold282 (.A(\dtop.vtop.pipeline.dz[0] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold283 (.A(\dtop.player_inst.synth.alu.carry ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold284 (.A(\dtop.vtop.pipeline.neg_t[5] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold285 (.A(uio_out[1]),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold286 (.A(\dtop.vtop.logo.addr[7] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold287 (.A(\dtop.vtop.rs.scan_y.phase[1] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0255_),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold289 (.A(uo_out[1]),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0110_),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold291 (.A(\dtop.vtop.pipeline.z[4] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold292 (.A(uo_out[4]),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold293 (.A(\dtop.vtop.pipeline.neg_t[0] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold294 (.A(_0267_),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold295 (.A(\dtop.vtop.pipeline.zg[3] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold296 (.A(\dtop.vtop.pipeline.zg_acc[3] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold297 (.A(uio_out[2]),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold298 (.A(uio_out[3]),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold299 (.A(\dtop.vtop.pipeline.zg[5] ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold300 (.A(\dtop.vtop.pipeline.dz[4] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0281_),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold302 (.A(\dtop.vtop.pipeline.z[12] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0298_),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold304 (.A(\dtop.vtop.pipeline.dz[1] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold305 (.A(\dtop.vtop.pipeline.z[7] ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold306 (.A(\dtop.vtop.pipeline.z[2] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold307 (.A(\dtop.vtop.pipeline.zg_acc[4] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold308 (.A(\dtop.vtop.pipeline.neg_t[3] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0270_),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold310 (.A(\dtop.vtop.pipeline.neg_t[7] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold311 (.A(\dtop.vtop.pipeline.zg_acc[0] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold312 (.A(\dtop.vtop.pipeline.z[13] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold313 (.A(\dtop.vtop.pipeline.z[8] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold314 (.A(\dtop.vtop.pipeline.zg[7] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold315 (.A(\dtop.vtop.pipeline.wave_index[1] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold316 (.A(_0370_),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold317 (.A(\dtop.vtop.rs.x_scan.phase[1] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold318 (.A(uo_out[0]),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold319 (.A(\dtop.detune_counter[16] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold320 (.A(\dtop.vtop.pipeline.z[9] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold321 (.A(uio_oe[5]),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold322 (.A(_0253_),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold323 (.A(\dtop.vtop.pipeline.z[10] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold324 (.A(\dtop.vtop.pipeline.z[3] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold325 (.A(\dtop.vtop.pipeline.z[1] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0287_),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold327 (.A(\dtop.vtop.pipeline.dz[5] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold328 (.A(\dtop.vtop.pipeline.zg_valid ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold329 (.A(\dtop.detune_counter[6] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold330 (.A(_1516_),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold331 (.A(uo_out[5]),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold332 (.A(\dtop.vtop.pipeline.zg[4] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold333 (.A(\dtop.vtop.rs.scan_y.phase[0] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold334 (.A(_1975_),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold335 (.A(\dtop.vtop.pipeline.z[6] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold336 (.A(\dtop.player_inst.synth.alu.acc[8] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold337 (.A(uo_out[3]),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold338 (.A(\dtop.vtop.pipeline.zg[6] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold339 (.A(\dtop.detune_counter[5] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold340 (.A(uio_out[6]),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold341 (.A(_0553_),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold342 (.A(\dtop.player_inst.program_addr[3] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold343 (.A(_0261_),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold344 (.A(_0089_),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold345 (.A(\dtop.vtop.pipeline.zg[8] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold346 (.A(_0078_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold347 (.A(\dtop.vtop.pipeline.z[5] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0025_),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold349 (.A(\dtop.detune_counter[8] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold350 (.A(_1519_),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold351 (.A(\dtop.player_inst.synth.alu.acc[9] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0085_),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold353 (.A(_3193_),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold354 (.A(_0101_),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold355 (.A(\dtop.player_inst.program_addr[4] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold356 (.A(_0262_),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold357 (.A(\dtop.vtop.pipeline.zg[9] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold358 (.A(\dtop.oct_counter[4] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0564_),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold360 (.A(\dtop.player_inst.program_addr[0] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold361 (.A(_1983_),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0258_),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold363 (.A(\dtop.vtop.logo.addr[8] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold364 (.A(\dtop.vtop.pipeline.nstep_zg[1] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold365 (.A(_0266_),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold366 (.A(\dtop.player_inst.program_addr[5] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0263_),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold368 (.A(\dtop.vtop.logo.addr[9] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold369 (.A(_0579_),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold370 (.A(\dtop.detune_counter[7] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold371 (.A(_1518_),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold372 (.A(\dtop.vtop.pipeline.nstep[0] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold373 (.A(_2653_),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold374 (.A(\dtop.vtop.pipeline.nstep[1] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold375 (.A(\dtop.enable ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold376 (.A(\dtop.player_inst.synth.alu.acc[7] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold377 (.A(\dtop.player_inst.synth.alu.acc[0] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold378 (.A(\dtop.oct_counter[3] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold379 (.A(_0562_),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold380 (.A(\dtop.player_inst.synth.alu.acc[4] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold381 (.A(_0014_),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0055_),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold383 (.A(_0577_),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold384 (.A(\dtop.vtop.pipeline.nstep_zg[0] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold385 (.A(\dtop.player_inst.synth.alu.acc[2] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold386 (.A(\dtop.oct_counter[5] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold387 (.A(_0566_),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold388 (.A(\dtop.player_inst.program_addr[2] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold389 (.A(\dtop.vtop.rs.saturated ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold390 (.A(_1943_),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold391 (.A(\dtop.player_inst.synth.alu.acc[1] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold392 (.A(\dtop.player_inst.synth.alu.acc[5] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold393 (.A(\dtop.player_inst.program_addr[1] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold394 (.A(\dtop.vtop.pipeline.z[3] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold395 (.A(\dtop.vtop.pipeline.z[1] ),
    .X(net712));
 sg13g2_antennanp ANTENNA_1 (.A(uio_out[1]));
 sg13g2_antennanp ANTENNA_2 (.A(uio_out[2]));
 sg13g2_antennanp ANTENNA_3 (.A(uio_out[3]));
 sg13g2_antennanp ANTENNA_4 (.A(uo_out[1]));
 sg13g2_antennanp ANTENNA_5 (.A(uo_out[3]));
 sg13g2_antennanp ANTENNA_6 (.A(uio_out[1]));
 sg13g2_antennanp ANTENNA_7 (.A(uio_out[3]));
 sg13g2_antennanp ANTENNA_8 (.A(uo_out[0]));
 sg13g2_antennanp ANTENNA_9 (.A(uo_out[1]));
 sg13g2_antennanp ANTENNA_10 (.A(uo_out[3]));
 sg13g2_antennanp ANTENNA_11 (.A(uio_out[1]));
 sg13g2_antennanp ANTENNA_12 (.A(uio_out[1]));
 sg13g2_antennanp ANTENNA_13 (.A(uio_out[3]));
 sg13g2_antennanp ANTENNA_14 (.A(uo_out[0]));
 sg13g2_antennanp ANTENNA_15 (.A(uo_out[0]));
 sg13g2_antennanp ANTENNA_16 (.A(uo_out[1]));
 sg13g2_antennanp ANTENNA_17 (.A(uo_out[3]));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_decap_8 FILLER_13_588 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_decap_8 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_637 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_8 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_decap_8 FILLER_13_798 ();
 sg13g2_decap_8 FILLER_13_805 ();
 sg13g2_decap_8 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_833 ();
 sg13g2_decap_8 FILLER_13_840 ();
 sg13g2_decap_8 FILLER_13_847 ();
 sg13g2_decap_8 FILLER_13_854 ();
 sg13g2_fill_1 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_8 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_511 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_574 ();
 sg13g2_decap_8 FILLER_14_581 ();
 sg13g2_decap_8 FILLER_14_588 ();
 sg13g2_decap_8 FILLER_14_595 ();
 sg13g2_decap_8 FILLER_14_602 ();
 sg13g2_decap_8 FILLER_14_609 ();
 sg13g2_decap_8 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_623 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_decap_8 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_decap_8 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_658 ();
 sg13g2_decap_8 FILLER_14_665 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_decap_8 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_decap_8 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_14_840 ();
 sg13g2_decap_8 FILLER_14_847 ();
 sg13g2_decap_8 FILLER_14_854 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_4 FILLER_15_70 ();
 sg13g2_fill_1 FILLER_15_74 ();
 sg13g2_fill_2 FILLER_15_80 ();
 sg13g2_fill_1 FILLER_15_82 ();
 sg13g2_decap_4 FILLER_15_91 ();
 sg13g2_fill_1 FILLER_15_100 ();
 sg13g2_decap_8 FILLER_15_113 ();
 sg13g2_fill_2 FILLER_15_120 ();
 sg13g2_decap_8 FILLER_15_127 ();
 sg13g2_decap_4 FILLER_15_134 ();
 sg13g2_fill_1 FILLER_15_138 ();
 sg13g2_decap_8 FILLER_15_144 ();
 sg13g2_decap_8 FILLER_15_151 ();
 sg13g2_fill_2 FILLER_15_158 ();
 sg13g2_fill_1 FILLER_15_167 ();
 sg13g2_decap_8 FILLER_15_178 ();
 sg13g2_fill_2 FILLER_15_185 ();
 sg13g2_decap_8 FILLER_15_192 ();
 sg13g2_decap_8 FILLER_15_199 ();
 sg13g2_decap_8 FILLER_15_206 ();
 sg13g2_decap_8 FILLER_15_213 ();
 sg13g2_decap_8 FILLER_15_220 ();
 sg13g2_decap_8 FILLER_15_227 ();
 sg13g2_decap_8 FILLER_15_234 ();
 sg13g2_decap_8 FILLER_15_241 ();
 sg13g2_decap_8 FILLER_15_248 ();
 sg13g2_decap_8 FILLER_15_255 ();
 sg13g2_decap_8 FILLER_15_262 ();
 sg13g2_decap_8 FILLER_15_269 ();
 sg13g2_decap_8 FILLER_15_276 ();
 sg13g2_decap_8 FILLER_15_283 ();
 sg13g2_decap_8 FILLER_15_290 ();
 sg13g2_decap_8 FILLER_15_297 ();
 sg13g2_decap_8 FILLER_15_304 ();
 sg13g2_decap_8 FILLER_15_311 ();
 sg13g2_decap_8 FILLER_15_318 ();
 sg13g2_decap_8 FILLER_15_325 ();
 sg13g2_decap_8 FILLER_15_332 ();
 sg13g2_decap_8 FILLER_15_339 ();
 sg13g2_decap_8 FILLER_15_346 ();
 sg13g2_decap_8 FILLER_15_353 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_decap_8 FILLER_15_367 ();
 sg13g2_decap_8 FILLER_15_374 ();
 sg13g2_decap_8 FILLER_15_381 ();
 sg13g2_decap_8 FILLER_15_388 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_15_409 ();
 sg13g2_decap_8 FILLER_15_416 ();
 sg13g2_decap_8 FILLER_15_423 ();
 sg13g2_decap_8 FILLER_15_430 ();
 sg13g2_decap_8 FILLER_15_437 ();
 sg13g2_decap_8 FILLER_15_444 ();
 sg13g2_decap_8 FILLER_15_451 ();
 sg13g2_decap_8 FILLER_15_458 ();
 sg13g2_decap_8 FILLER_15_465 ();
 sg13g2_decap_8 FILLER_15_472 ();
 sg13g2_decap_8 FILLER_15_479 ();
 sg13g2_decap_8 FILLER_15_486 ();
 sg13g2_decap_8 FILLER_15_493 ();
 sg13g2_decap_8 FILLER_15_500 ();
 sg13g2_decap_8 FILLER_15_507 ();
 sg13g2_decap_8 FILLER_15_514 ();
 sg13g2_decap_8 FILLER_15_521 ();
 sg13g2_decap_8 FILLER_15_528 ();
 sg13g2_decap_8 FILLER_15_535 ();
 sg13g2_decap_8 FILLER_15_542 ();
 sg13g2_decap_8 FILLER_15_549 ();
 sg13g2_decap_8 FILLER_15_556 ();
 sg13g2_decap_8 FILLER_15_563 ();
 sg13g2_decap_8 FILLER_15_570 ();
 sg13g2_decap_8 FILLER_15_577 ();
 sg13g2_decap_8 FILLER_15_584 ();
 sg13g2_decap_8 FILLER_15_591 ();
 sg13g2_decap_8 FILLER_15_598 ();
 sg13g2_decap_8 FILLER_15_605 ();
 sg13g2_decap_8 FILLER_15_612 ();
 sg13g2_decap_8 FILLER_15_619 ();
 sg13g2_decap_8 FILLER_15_626 ();
 sg13g2_decap_8 FILLER_15_633 ();
 sg13g2_decap_8 FILLER_15_640 ();
 sg13g2_decap_8 FILLER_15_647 ();
 sg13g2_decap_8 FILLER_15_654 ();
 sg13g2_decap_8 FILLER_15_661 ();
 sg13g2_decap_8 FILLER_15_668 ();
 sg13g2_decap_8 FILLER_15_675 ();
 sg13g2_decap_8 FILLER_15_682 ();
 sg13g2_decap_8 FILLER_15_689 ();
 sg13g2_decap_8 FILLER_15_696 ();
 sg13g2_decap_8 FILLER_15_703 ();
 sg13g2_decap_8 FILLER_15_710 ();
 sg13g2_decap_8 FILLER_15_717 ();
 sg13g2_decap_8 FILLER_15_724 ();
 sg13g2_decap_8 FILLER_15_731 ();
 sg13g2_decap_8 FILLER_15_738 ();
 sg13g2_decap_8 FILLER_15_745 ();
 sg13g2_decap_8 FILLER_15_752 ();
 sg13g2_decap_8 FILLER_15_759 ();
 sg13g2_decap_8 FILLER_15_766 ();
 sg13g2_decap_8 FILLER_15_773 ();
 sg13g2_decap_8 FILLER_15_780 ();
 sg13g2_decap_8 FILLER_15_787 ();
 sg13g2_decap_8 FILLER_15_794 ();
 sg13g2_decap_8 FILLER_15_801 ();
 sg13g2_decap_8 FILLER_15_808 ();
 sg13g2_decap_8 FILLER_15_815 ();
 sg13g2_decap_8 FILLER_15_822 ();
 sg13g2_decap_8 FILLER_15_829 ();
 sg13g2_decap_8 FILLER_15_836 ();
 sg13g2_decap_8 FILLER_15_843 ();
 sg13g2_decap_8 FILLER_15_850 ();
 sg13g2_decap_4 FILLER_15_857 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_4 FILLER_16_49 ();
 sg13g2_fill_2 FILLER_16_53 ();
 sg13g2_fill_2 FILLER_16_63 ();
 sg13g2_fill_2 FILLER_16_75 ();
 sg13g2_fill_1 FILLER_16_77 ();
 sg13g2_fill_2 FILLER_16_91 ();
 sg13g2_fill_1 FILLER_16_113 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_fill_2 FILLER_16_141 ();
 sg13g2_fill_1 FILLER_16_143 ();
 sg13g2_fill_1 FILLER_16_149 ();
 sg13g2_fill_2 FILLER_16_192 ();
 sg13g2_decap_8 FILLER_16_199 ();
 sg13g2_decap_4 FILLER_16_206 ();
 sg13g2_fill_2 FILLER_16_210 ();
 sg13g2_decap_4 FILLER_16_220 ();
 sg13g2_fill_1 FILLER_16_224 ();
 sg13g2_fill_2 FILLER_16_233 ();
 sg13g2_decap_8 FILLER_16_240 ();
 sg13g2_decap_8 FILLER_16_247 ();
 sg13g2_decap_8 FILLER_16_254 ();
 sg13g2_decap_8 FILLER_16_261 ();
 sg13g2_decap_8 FILLER_16_268 ();
 sg13g2_decap_8 FILLER_16_275 ();
 sg13g2_decap_8 FILLER_16_282 ();
 sg13g2_decap_8 FILLER_16_289 ();
 sg13g2_decap_8 FILLER_16_296 ();
 sg13g2_decap_8 FILLER_16_303 ();
 sg13g2_decap_8 FILLER_16_310 ();
 sg13g2_decap_8 FILLER_16_317 ();
 sg13g2_decap_8 FILLER_16_324 ();
 sg13g2_decap_8 FILLER_16_331 ();
 sg13g2_decap_8 FILLER_16_338 ();
 sg13g2_decap_8 FILLER_16_345 ();
 sg13g2_decap_8 FILLER_16_352 ();
 sg13g2_decap_8 FILLER_16_359 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_decap_8 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_16_415 ();
 sg13g2_decap_8 FILLER_16_422 ();
 sg13g2_decap_8 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_16_436 ();
 sg13g2_decap_8 FILLER_16_443 ();
 sg13g2_decap_8 FILLER_16_450 ();
 sg13g2_decap_8 FILLER_16_457 ();
 sg13g2_decap_8 FILLER_16_464 ();
 sg13g2_decap_8 FILLER_16_471 ();
 sg13g2_decap_8 FILLER_16_478 ();
 sg13g2_decap_8 FILLER_16_485 ();
 sg13g2_decap_8 FILLER_16_492 ();
 sg13g2_decap_8 FILLER_16_499 ();
 sg13g2_decap_8 FILLER_16_506 ();
 sg13g2_decap_8 FILLER_16_513 ();
 sg13g2_decap_8 FILLER_16_520 ();
 sg13g2_decap_8 FILLER_16_527 ();
 sg13g2_decap_8 FILLER_16_534 ();
 sg13g2_decap_8 FILLER_16_541 ();
 sg13g2_decap_8 FILLER_16_548 ();
 sg13g2_decap_8 FILLER_16_555 ();
 sg13g2_decap_8 FILLER_16_562 ();
 sg13g2_decap_8 FILLER_16_569 ();
 sg13g2_decap_8 FILLER_16_576 ();
 sg13g2_decap_8 FILLER_16_583 ();
 sg13g2_decap_8 FILLER_16_590 ();
 sg13g2_decap_8 FILLER_16_597 ();
 sg13g2_decap_8 FILLER_16_604 ();
 sg13g2_decap_8 FILLER_16_611 ();
 sg13g2_decap_8 FILLER_16_618 ();
 sg13g2_decap_8 FILLER_16_625 ();
 sg13g2_decap_8 FILLER_16_632 ();
 sg13g2_decap_8 FILLER_16_639 ();
 sg13g2_decap_8 FILLER_16_646 ();
 sg13g2_decap_8 FILLER_16_653 ();
 sg13g2_decap_8 FILLER_16_660 ();
 sg13g2_decap_8 FILLER_16_667 ();
 sg13g2_decap_8 FILLER_16_674 ();
 sg13g2_decap_8 FILLER_16_681 ();
 sg13g2_decap_8 FILLER_16_688 ();
 sg13g2_decap_8 FILLER_16_695 ();
 sg13g2_decap_8 FILLER_16_702 ();
 sg13g2_decap_8 FILLER_16_709 ();
 sg13g2_decap_8 FILLER_16_716 ();
 sg13g2_decap_8 FILLER_16_723 ();
 sg13g2_decap_8 FILLER_16_730 ();
 sg13g2_decap_8 FILLER_16_737 ();
 sg13g2_decap_8 FILLER_16_744 ();
 sg13g2_decap_8 FILLER_16_751 ();
 sg13g2_decap_8 FILLER_16_758 ();
 sg13g2_decap_8 FILLER_16_765 ();
 sg13g2_decap_8 FILLER_16_772 ();
 sg13g2_decap_8 FILLER_16_779 ();
 sg13g2_decap_8 FILLER_16_786 ();
 sg13g2_decap_8 FILLER_16_793 ();
 sg13g2_decap_8 FILLER_16_800 ();
 sg13g2_decap_8 FILLER_16_807 ();
 sg13g2_decap_8 FILLER_16_814 ();
 sg13g2_decap_8 FILLER_16_821 ();
 sg13g2_decap_8 FILLER_16_828 ();
 sg13g2_decap_8 FILLER_16_835 ();
 sg13g2_decap_8 FILLER_16_842 ();
 sg13g2_decap_8 FILLER_16_849 ();
 sg13g2_decap_4 FILLER_16_856 ();
 sg13g2_fill_2 FILLER_16_860 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_fill_1 FILLER_17_42 ();
 sg13g2_fill_1 FILLER_17_65 ();
 sg13g2_fill_2 FILLER_17_87 ();
 sg13g2_fill_2 FILLER_17_94 ();
 sg13g2_fill_1 FILLER_17_96 ();
 sg13g2_fill_1 FILLER_17_110 ();
 sg13g2_fill_2 FILLER_17_132 ();
 sg13g2_fill_1 FILLER_17_144 ();
 sg13g2_fill_1 FILLER_17_154 ();
 sg13g2_fill_1 FILLER_17_169 ();
 sg13g2_fill_2 FILLER_17_199 ();
 sg13g2_fill_2 FILLER_17_222 ();
 sg13g2_fill_1 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_249 ();
 sg13g2_decap_8 FILLER_17_256 ();
 sg13g2_decap_8 FILLER_17_263 ();
 sg13g2_decap_8 FILLER_17_270 ();
 sg13g2_decap_8 FILLER_17_277 ();
 sg13g2_decap_8 FILLER_17_284 ();
 sg13g2_decap_8 FILLER_17_291 ();
 sg13g2_decap_8 FILLER_17_298 ();
 sg13g2_decap_8 FILLER_17_305 ();
 sg13g2_decap_8 FILLER_17_312 ();
 sg13g2_decap_8 FILLER_17_319 ();
 sg13g2_decap_8 FILLER_17_326 ();
 sg13g2_decap_8 FILLER_17_333 ();
 sg13g2_decap_8 FILLER_17_340 ();
 sg13g2_decap_8 FILLER_17_347 ();
 sg13g2_decap_8 FILLER_17_354 ();
 sg13g2_decap_8 FILLER_17_361 ();
 sg13g2_decap_8 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_8 FILLER_17_403 ();
 sg13g2_decap_8 FILLER_17_410 ();
 sg13g2_decap_8 FILLER_17_417 ();
 sg13g2_decap_8 FILLER_17_424 ();
 sg13g2_decap_8 FILLER_17_431 ();
 sg13g2_decap_8 FILLER_17_438 ();
 sg13g2_decap_8 FILLER_17_445 ();
 sg13g2_decap_8 FILLER_17_452 ();
 sg13g2_decap_8 FILLER_17_459 ();
 sg13g2_decap_8 FILLER_17_466 ();
 sg13g2_decap_8 FILLER_17_473 ();
 sg13g2_decap_8 FILLER_17_480 ();
 sg13g2_decap_8 FILLER_17_487 ();
 sg13g2_decap_8 FILLER_17_494 ();
 sg13g2_decap_8 FILLER_17_501 ();
 sg13g2_decap_8 FILLER_17_508 ();
 sg13g2_decap_8 FILLER_17_515 ();
 sg13g2_decap_8 FILLER_17_522 ();
 sg13g2_decap_8 FILLER_17_529 ();
 sg13g2_decap_8 FILLER_17_536 ();
 sg13g2_decap_8 FILLER_17_543 ();
 sg13g2_decap_8 FILLER_17_550 ();
 sg13g2_decap_8 FILLER_17_557 ();
 sg13g2_decap_8 FILLER_17_564 ();
 sg13g2_decap_8 FILLER_17_571 ();
 sg13g2_decap_8 FILLER_17_578 ();
 sg13g2_decap_8 FILLER_17_585 ();
 sg13g2_decap_8 FILLER_17_592 ();
 sg13g2_decap_8 FILLER_17_599 ();
 sg13g2_decap_8 FILLER_17_606 ();
 sg13g2_decap_8 FILLER_17_613 ();
 sg13g2_decap_8 FILLER_17_620 ();
 sg13g2_decap_8 FILLER_17_627 ();
 sg13g2_decap_8 FILLER_17_634 ();
 sg13g2_decap_8 FILLER_17_641 ();
 sg13g2_decap_8 FILLER_17_648 ();
 sg13g2_decap_8 FILLER_17_655 ();
 sg13g2_decap_8 FILLER_17_662 ();
 sg13g2_decap_8 FILLER_17_669 ();
 sg13g2_decap_8 FILLER_17_676 ();
 sg13g2_decap_8 FILLER_17_683 ();
 sg13g2_decap_8 FILLER_17_690 ();
 sg13g2_decap_8 FILLER_17_697 ();
 sg13g2_decap_8 FILLER_17_704 ();
 sg13g2_decap_8 FILLER_17_711 ();
 sg13g2_decap_8 FILLER_17_718 ();
 sg13g2_decap_8 FILLER_17_725 ();
 sg13g2_decap_8 FILLER_17_732 ();
 sg13g2_decap_8 FILLER_17_739 ();
 sg13g2_decap_8 FILLER_17_746 ();
 sg13g2_decap_8 FILLER_17_753 ();
 sg13g2_decap_8 FILLER_17_760 ();
 sg13g2_decap_8 FILLER_17_767 ();
 sg13g2_decap_8 FILLER_17_774 ();
 sg13g2_decap_8 FILLER_17_781 ();
 sg13g2_decap_8 FILLER_17_788 ();
 sg13g2_decap_8 FILLER_17_795 ();
 sg13g2_decap_8 FILLER_17_802 ();
 sg13g2_decap_8 FILLER_17_809 ();
 sg13g2_decap_8 FILLER_17_816 ();
 sg13g2_decap_8 FILLER_17_823 ();
 sg13g2_decap_8 FILLER_17_830 ();
 sg13g2_decap_8 FILLER_17_837 ();
 sg13g2_decap_8 FILLER_17_844 ();
 sg13g2_decap_8 FILLER_17_851 ();
 sg13g2_decap_4 FILLER_17_858 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_4 FILLER_18_35 ();
 sg13g2_fill_1 FILLER_18_49 ();
 sg13g2_fill_2 FILLER_18_55 ();
 sg13g2_fill_2 FILLER_18_67 ();
 sg13g2_fill_1 FILLER_18_69 ();
 sg13g2_decap_4 FILLER_18_102 ();
 sg13g2_decap_4 FILLER_18_126 ();
 sg13g2_fill_2 FILLER_18_130 ();
 sg13g2_fill_2 FILLER_18_138 ();
 sg13g2_fill_1 FILLER_18_143 ();
 sg13g2_decap_4 FILLER_18_149 ();
 sg13g2_fill_1 FILLER_18_153 ();
 sg13g2_decap_4 FILLER_18_159 ();
 sg13g2_fill_2 FILLER_18_167 ();
 sg13g2_fill_1 FILLER_18_175 ();
 sg13g2_fill_1 FILLER_18_187 ();
 sg13g2_fill_2 FILLER_18_208 ();
 sg13g2_fill_1 FILLER_18_210 ();
 sg13g2_decap_4 FILLER_18_222 ();
 sg13g2_fill_2 FILLER_18_226 ();
 sg13g2_decap_8 FILLER_18_241 ();
 sg13g2_decap_8 FILLER_18_248 ();
 sg13g2_decap_8 FILLER_18_255 ();
 sg13g2_decap_8 FILLER_18_262 ();
 sg13g2_decap_8 FILLER_18_269 ();
 sg13g2_decap_8 FILLER_18_276 ();
 sg13g2_decap_8 FILLER_18_283 ();
 sg13g2_decap_8 FILLER_18_290 ();
 sg13g2_decap_8 FILLER_18_297 ();
 sg13g2_decap_8 FILLER_18_304 ();
 sg13g2_decap_8 FILLER_18_311 ();
 sg13g2_decap_8 FILLER_18_318 ();
 sg13g2_decap_8 FILLER_18_325 ();
 sg13g2_decap_8 FILLER_18_332 ();
 sg13g2_decap_8 FILLER_18_339 ();
 sg13g2_decap_8 FILLER_18_346 ();
 sg13g2_decap_8 FILLER_18_353 ();
 sg13g2_decap_8 FILLER_18_360 ();
 sg13g2_decap_8 FILLER_18_367 ();
 sg13g2_decap_8 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_18_409 ();
 sg13g2_decap_8 FILLER_18_416 ();
 sg13g2_decap_8 FILLER_18_423 ();
 sg13g2_decap_8 FILLER_18_430 ();
 sg13g2_decap_8 FILLER_18_437 ();
 sg13g2_decap_8 FILLER_18_444 ();
 sg13g2_decap_8 FILLER_18_451 ();
 sg13g2_decap_8 FILLER_18_458 ();
 sg13g2_decap_8 FILLER_18_465 ();
 sg13g2_decap_8 FILLER_18_472 ();
 sg13g2_decap_8 FILLER_18_479 ();
 sg13g2_decap_8 FILLER_18_486 ();
 sg13g2_decap_8 FILLER_18_493 ();
 sg13g2_decap_8 FILLER_18_500 ();
 sg13g2_decap_8 FILLER_18_507 ();
 sg13g2_decap_8 FILLER_18_514 ();
 sg13g2_decap_8 FILLER_18_521 ();
 sg13g2_decap_8 FILLER_18_528 ();
 sg13g2_decap_8 FILLER_18_535 ();
 sg13g2_decap_8 FILLER_18_542 ();
 sg13g2_decap_8 FILLER_18_549 ();
 sg13g2_decap_8 FILLER_18_556 ();
 sg13g2_decap_8 FILLER_18_563 ();
 sg13g2_decap_8 FILLER_18_570 ();
 sg13g2_decap_8 FILLER_18_577 ();
 sg13g2_decap_8 FILLER_18_584 ();
 sg13g2_decap_8 FILLER_18_591 ();
 sg13g2_decap_8 FILLER_18_598 ();
 sg13g2_decap_8 FILLER_18_605 ();
 sg13g2_decap_8 FILLER_18_612 ();
 sg13g2_decap_8 FILLER_18_619 ();
 sg13g2_decap_8 FILLER_18_626 ();
 sg13g2_decap_8 FILLER_18_633 ();
 sg13g2_decap_8 FILLER_18_640 ();
 sg13g2_decap_8 FILLER_18_647 ();
 sg13g2_decap_8 FILLER_18_654 ();
 sg13g2_decap_8 FILLER_18_661 ();
 sg13g2_decap_8 FILLER_18_668 ();
 sg13g2_decap_8 FILLER_18_675 ();
 sg13g2_decap_8 FILLER_18_682 ();
 sg13g2_decap_8 FILLER_18_689 ();
 sg13g2_decap_8 FILLER_18_696 ();
 sg13g2_decap_8 FILLER_18_703 ();
 sg13g2_decap_8 FILLER_18_710 ();
 sg13g2_decap_8 FILLER_18_717 ();
 sg13g2_decap_8 FILLER_18_724 ();
 sg13g2_decap_8 FILLER_18_731 ();
 sg13g2_decap_8 FILLER_18_738 ();
 sg13g2_decap_8 FILLER_18_745 ();
 sg13g2_decap_8 FILLER_18_752 ();
 sg13g2_decap_8 FILLER_18_759 ();
 sg13g2_decap_8 FILLER_18_766 ();
 sg13g2_decap_8 FILLER_18_773 ();
 sg13g2_decap_8 FILLER_18_780 ();
 sg13g2_decap_8 FILLER_18_787 ();
 sg13g2_decap_8 FILLER_18_794 ();
 sg13g2_decap_8 FILLER_18_801 ();
 sg13g2_decap_8 FILLER_18_808 ();
 sg13g2_decap_8 FILLER_18_815 ();
 sg13g2_decap_8 FILLER_18_822 ();
 sg13g2_decap_8 FILLER_18_829 ();
 sg13g2_decap_8 FILLER_18_836 ();
 sg13g2_decap_8 FILLER_18_843 ();
 sg13g2_decap_8 FILLER_18_850 ();
 sg13g2_decap_4 FILLER_18_857 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_fill_2 FILLER_19_58 ();
 sg13g2_fill_1 FILLER_19_74 ();
 sg13g2_fill_2 FILLER_19_85 ();
 sg13g2_fill_1 FILLER_19_87 ();
 sg13g2_fill_2 FILLER_19_103 ();
 sg13g2_fill_1 FILLER_19_105 ();
 sg13g2_decap_4 FILLER_19_133 ();
 sg13g2_fill_1 FILLER_19_137 ();
 sg13g2_decap_4 FILLER_19_157 ();
 sg13g2_fill_2 FILLER_19_161 ();
 sg13g2_fill_2 FILLER_19_179 ();
 sg13g2_fill_1 FILLER_19_181 ();
 sg13g2_fill_2 FILLER_19_197 ();
 sg13g2_fill_1 FILLER_19_199 ();
 sg13g2_fill_2 FILLER_19_205 ();
 sg13g2_decap_8 FILLER_19_240 ();
 sg13g2_decap_8 FILLER_19_247 ();
 sg13g2_decap_8 FILLER_19_254 ();
 sg13g2_decap_8 FILLER_19_261 ();
 sg13g2_decap_8 FILLER_19_268 ();
 sg13g2_decap_8 FILLER_19_275 ();
 sg13g2_decap_8 FILLER_19_282 ();
 sg13g2_decap_8 FILLER_19_289 ();
 sg13g2_decap_8 FILLER_19_296 ();
 sg13g2_decap_8 FILLER_19_303 ();
 sg13g2_decap_8 FILLER_19_310 ();
 sg13g2_decap_8 FILLER_19_317 ();
 sg13g2_decap_8 FILLER_19_324 ();
 sg13g2_decap_8 FILLER_19_331 ();
 sg13g2_decap_8 FILLER_19_338 ();
 sg13g2_decap_8 FILLER_19_345 ();
 sg13g2_decap_8 FILLER_19_352 ();
 sg13g2_decap_8 FILLER_19_359 ();
 sg13g2_decap_8 FILLER_19_366 ();
 sg13g2_decap_8 FILLER_19_373 ();
 sg13g2_decap_8 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_decap_8 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_19_415 ();
 sg13g2_decap_8 FILLER_19_422 ();
 sg13g2_decap_8 FILLER_19_429 ();
 sg13g2_decap_8 FILLER_19_436 ();
 sg13g2_decap_8 FILLER_19_443 ();
 sg13g2_decap_8 FILLER_19_450 ();
 sg13g2_decap_8 FILLER_19_457 ();
 sg13g2_decap_8 FILLER_19_464 ();
 sg13g2_decap_8 FILLER_19_471 ();
 sg13g2_decap_8 FILLER_19_478 ();
 sg13g2_decap_8 FILLER_19_485 ();
 sg13g2_decap_8 FILLER_19_492 ();
 sg13g2_decap_8 FILLER_19_499 ();
 sg13g2_decap_8 FILLER_19_506 ();
 sg13g2_decap_8 FILLER_19_513 ();
 sg13g2_decap_8 FILLER_19_520 ();
 sg13g2_decap_8 FILLER_19_527 ();
 sg13g2_decap_8 FILLER_19_534 ();
 sg13g2_decap_8 FILLER_19_541 ();
 sg13g2_decap_8 FILLER_19_548 ();
 sg13g2_decap_8 FILLER_19_555 ();
 sg13g2_decap_8 FILLER_19_562 ();
 sg13g2_decap_8 FILLER_19_569 ();
 sg13g2_decap_8 FILLER_19_576 ();
 sg13g2_decap_8 FILLER_19_583 ();
 sg13g2_decap_8 FILLER_19_590 ();
 sg13g2_decap_8 FILLER_19_597 ();
 sg13g2_decap_8 FILLER_19_604 ();
 sg13g2_decap_8 FILLER_19_611 ();
 sg13g2_decap_8 FILLER_19_618 ();
 sg13g2_decap_8 FILLER_19_625 ();
 sg13g2_decap_8 FILLER_19_632 ();
 sg13g2_decap_8 FILLER_19_639 ();
 sg13g2_decap_8 FILLER_19_646 ();
 sg13g2_decap_8 FILLER_19_653 ();
 sg13g2_decap_8 FILLER_19_660 ();
 sg13g2_decap_8 FILLER_19_667 ();
 sg13g2_decap_8 FILLER_19_674 ();
 sg13g2_decap_8 FILLER_19_681 ();
 sg13g2_decap_8 FILLER_19_688 ();
 sg13g2_decap_8 FILLER_19_695 ();
 sg13g2_decap_8 FILLER_19_702 ();
 sg13g2_decap_8 FILLER_19_709 ();
 sg13g2_decap_8 FILLER_19_716 ();
 sg13g2_decap_8 FILLER_19_723 ();
 sg13g2_decap_8 FILLER_19_730 ();
 sg13g2_decap_8 FILLER_19_737 ();
 sg13g2_decap_8 FILLER_19_744 ();
 sg13g2_decap_8 FILLER_19_751 ();
 sg13g2_decap_8 FILLER_19_758 ();
 sg13g2_decap_8 FILLER_19_765 ();
 sg13g2_decap_8 FILLER_19_772 ();
 sg13g2_decap_8 FILLER_19_779 ();
 sg13g2_decap_8 FILLER_19_786 ();
 sg13g2_decap_8 FILLER_19_793 ();
 sg13g2_decap_8 FILLER_19_800 ();
 sg13g2_decap_8 FILLER_19_807 ();
 sg13g2_decap_8 FILLER_19_814 ();
 sg13g2_decap_8 FILLER_19_821 ();
 sg13g2_decap_8 FILLER_19_828 ();
 sg13g2_decap_8 FILLER_19_835 ();
 sg13g2_decap_8 FILLER_19_842 ();
 sg13g2_decap_8 FILLER_19_849 ();
 sg13g2_decap_4 FILLER_19_856 ();
 sg13g2_fill_2 FILLER_19_860 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_fill_2 FILLER_20_42 ();
 sg13g2_fill_2 FILLER_20_60 ();
 sg13g2_fill_1 FILLER_20_62 ();
 sg13g2_fill_2 FILLER_20_73 ();
 sg13g2_fill_1 FILLER_20_75 ();
 sg13g2_fill_1 FILLER_20_81 ();
 sg13g2_fill_2 FILLER_20_88 ();
 sg13g2_fill_2 FILLER_20_98 ();
 sg13g2_fill_1 FILLER_20_100 ();
 sg13g2_decap_4 FILLER_20_120 ();
 sg13g2_decap_8 FILLER_20_132 ();
 sg13g2_fill_2 FILLER_20_165 ();
 sg13g2_fill_2 FILLER_20_187 ();
 sg13g2_decap_4 FILLER_20_215 ();
 sg13g2_fill_2 FILLER_20_219 ();
 sg13g2_fill_1 FILLER_20_234 ();
 sg13g2_decap_8 FILLER_20_243 ();
 sg13g2_decap_8 FILLER_20_250 ();
 sg13g2_decap_8 FILLER_20_257 ();
 sg13g2_decap_8 FILLER_20_264 ();
 sg13g2_decap_8 FILLER_20_271 ();
 sg13g2_decap_8 FILLER_20_278 ();
 sg13g2_decap_8 FILLER_20_285 ();
 sg13g2_decap_8 FILLER_20_292 ();
 sg13g2_decap_8 FILLER_20_299 ();
 sg13g2_decap_8 FILLER_20_306 ();
 sg13g2_decap_8 FILLER_20_313 ();
 sg13g2_decap_8 FILLER_20_320 ();
 sg13g2_decap_8 FILLER_20_327 ();
 sg13g2_decap_8 FILLER_20_334 ();
 sg13g2_decap_8 FILLER_20_341 ();
 sg13g2_decap_8 FILLER_20_348 ();
 sg13g2_decap_8 FILLER_20_355 ();
 sg13g2_decap_8 FILLER_20_362 ();
 sg13g2_decap_8 FILLER_20_369 ();
 sg13g2_decap_8 FILLER_20_376 ();
 sg13g2_decap_8 FILLER_20_383 ();
 sg13g2_decap_8 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_397 ();
 sg13g2_decap_8 FILLER_20_404 ();
 sg13g2_decap_8 FILLER_20_411 ();
 sg13g2_decap_8 FILLER_20_418 ();
 sg13g2_decap_8 FILLER_20_425 ();
 sg13g2_decap_8 FILLER_20_432 ();
 sg13g2_decap_8 FILLER_20_439 ();
 sg13g2_decap_8 FILLER_20_446 ();
 sg13g2_decap_8 FILLER_20_453 ();
 sg13g2_decap_8 FILLER_20_460 ();
 sg13g2_decap_8 FILLER_20_467 ();
 sg13g2_decap_8 FILLER_20_474 ();
 sg13g2_decap_8 FILLER_20_481 ();
 sg13g2_decap_8 FILLER_20_488 ();
 sg13g2_decap_8 FILLER_20_495 ();
 sg13g2_decap_8 FILLER_20_502 ();
 sg13g2_decap_8 FILLER_20_509 ();
 sg13g2_decap_8 FILLER_20_516 ();
 sg13g2_decap_8 FILLER_20_523 ();
 sg13g2_decap_8 FILLER_20_530 ();
 sg13g2_decap_8 FILLER_20_537 ();
 sg13g2_decap_8 FILLER_20_544 ();
 sg13g2_decap_8 FILLER_20_551 ();
 sg13g2_decap_8 FILLER_20_558 ();
 sg13g2_decap_8 FILLER_20_565 ();
 sg13g2_decap_8 FILLER_20_572 ();
 sg13g2_decap_8 FILLER_20_579 ();
 sg13g2_decap_8 FILLER_20_586 ();
 sg13g2_decap_8 FILLER_20_593 ();
 sg13g2_decap_8 FILLER_20_600 ();
 sg13g2_decap_8 FILLER_20_607 ();
 sg13g2_decap_8 FILLER_20_614 ();
 sg13g2_decap_8 FILLER_20_621 ();
 sg13g2_decap_8 FILLER_20_628 ();
 sg13g2_decap_8 FILLER_20_635 ();
 sg13g2_decap_8 FILLER_20_642 ();
 sg13g2_decap_8 FILLER_20_649 ();
 sg13g2_decap_8 FILLER_20_656 ();
 sg13g2_decap_8 FILLER_20_663 ();
 sg13g2_decap_8 FILLER_20_670 ();
 sg13g2_decap_8 FILLER_20_677 ();
 sg13g2_decap_8 FILLER_20_684 ();
 sg13g2_decap_8 FILLER_20_691 ();
 sg13g2_decap_8 FILLER_20_698 ();
 sg13g2_decap_8 FILLER_20_705 ();
 sg13g2_decap_8 FILLER_20_712 ();
 sg13g2_decap_8 FILLER_20_719 ();
 sg13g2_decap_8 FILLER_20_726 ();
 sg13g2_decap_8 FILLER_20_733 ();
 sg13g2_decap_8 FILLER_20_740 ();
 sg13g2_decap_8 FILLER_20_747 ();
 sg13g2_decap_8 FILLER_20_754 ();
 sg13g2_decap_8 FILLER_20_761 ();
 sg13g2_decap_8 FILLER_20_768 ();
 sg13g2_decap_8 FILLER_20_775 ();
 sg13g2_decap_8 FILLER_20_782 ();
 sg13g2_decap_8 FILLER_20_789 ();
 sg13g2_decap_8 FILLER_20_796 ();
 sg13g2_decap_8 FILLER_20_803 ();
 sg13g2_decap_8 FILLER_20_810 ();
 sg13g2_decap_8 FILLER_20_817 ();
 sg13g2_decap_8 FILLER_20_824 ();
 sg13g2_decap_8 FILLER_20_831 ();
 sg13g2_decap_8 FILLER_20_838 ();
 sg13g2_decap_8 FILLER_20_845 ();
 sg13g2_decap_8 FILLER_20_852 ();
 sg13g2_fill_2 FILLER_20_859 ();
 sg13g2_fill_1 FILLER_20_861 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_4 FILLER_21_28 ();
 sg13g2_fill_2 FILLER_21_32 ();
 sg13g2_fill_1 FILLER_21_61 ();
 sg13g2_fill_2 FILLER_21_76 ();
 sg13g2_fill_1 FILLER_21_78 ();
 sg13g2_fill_1 FILLER_21_87 ();
 sg13g2_fill_2 FILLER_21_105 ();
 sg13g2_fill_2 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_139 ();
 sg13g2_fill_1 FILLER_21_166 ();
 sg13g2_fill_2 FILLER_21_193 ();
 sg13g2_fill_1 FILLER_21_195 ();
 sg13g2_decap_8 FILLER_21_239 ();
 sg13g2_decap_8 FILLER_21_246 ();
 sg13g2_decap_8 FILLER_21_279 ();
 sg13g2_decap_4 FILLER_21_286 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_fill_1 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_316 ();
 sg13g2_decap_8 FILLER_21_323 ();
 sg13g2_fill_1 FILLER_21_330 ();
 sg13g2_decap_8 FILLER_21_335 ();
 sg13g2_decap_8 FILLER_21_342 ();
 sg13g2_decap_8 FILLER_21_349 ();
 sg13g2_decap_8 FILLER_21_356 ();
 sg13g2_decap_8 FILLER_21_363 ();
 sg13g2_decap_8 FILLER_21_370 ();
 sg13g2_decap_8 FILLER_21_377 ();
 sg13g2_decap_8 FILLER_21_384 ();
 sg13g2_decap_8 FILLER_21_391 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_decap_8 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_21_412 ();
 sg13g2_decap_8 FILLER_21_419 ();
 sg13g2_decap_8 FILLER_21_426 ();
 sg13g2_decap_8 FILLER_21_433 ();
 sg13g2_decap_8 FILLER_21_440 ();
 sg13g2_decap_8 FILLER_21_447 ();
 sg13g2_decap_8 FILLER_21_454 ();
 sg13g2_decap_8 FILLER_21_461 ();
 sg13g2_decap_8 FILLER_21_468 ();
 sg13g2_decap_8 FILLER_21_475 ();
 sg13g2_decap_8 FILLER_21_482 ();
 sg13g2_decap_8 FILLER_21_489 ();
 sg13g2_decap_8 FILLER_21_496 ();
 sg13g2_decap_8 FILLER_21_503 ();
 sg13g2_decap_8 FILLER_21_510 ();
 sg13g2_decap_8 FILLER_21_517 ();
 sg13g2_decap_8 FILLER_21_524 ();
 sg13g2_decap_8 FILLER_21_531 ();
 sg13g2_decap_8 FILLER_21_538 ();
 sg13g2_decap_8 FILLER_21_545 ();
 sg13g2_decap_8 FILLER_21_552 ();
 sg13g2_decap_8 FILLER_21_559 ();
 sg13g2_decap_8 FILLER_21_566 ();
 sg13g2_decap_8 FILLER_21_573 ();
 sg13g2_decap_8 FILLER_21_580 ();
 sg13g2_decap_8 FILLER_21_587 ();
 sg13g2_decap_8 FILLER_21_594 ();
 sg13g2_decap_8 FILLER_21_601 ();
 sg13g2_decap_8 FILLER_21_608 ();
 sg13g2_decap_8 FILLER_21_615 ();
 sg13g2_decap_8 FILLER_21_622 ();
 sg13g2_decap_8 FILLER_21_629 ();
 sg13g2_decap_8 FILLER_21_636 ();
 sg13g2_decap_8 FILLER_21_643 ();
 sg13g2_decap_8 FILLER_21_650 ();
 sg13g2_decap_8 FILLER_21_657 ();
 sg13g2_decap_8 FILLER_21_664 ();
 sg13g2_decap_8 FILLER_21_671 ();
 sg13g2_decap_8 FILLER_21_678 ();
 sg13g2_decap_8 FILLER_21_685 ();
 sg13g2_decap_8 FILLER_21_692 ();
 sg13g2_decap_8 FILLER_21_699 ();
 sg13g2_decap_8 FILLER_21_706 ();
 sg13g2_decap_8 FILLER_21_713 ();
 sg13g2_decap_8 FILLER_21_720 ();
 sg13g2_decap_8 FILLER_21_727 ();
 sg13g2_decap_8 FILLER_21_734 ();
 sg13g2_decap_8 FILLER_21_741 ();
 sg13g2_decap_8 FILLER_21_748 ();
 sg13g2_decap_8 FILLER_21_755 ();
 sg13g2_decap_8 FILLER_21_762 ();
 sg13g2_decap_8 FILLER_21_769 ();
 sg13g2_decap_8 FILLER_21_776 ();
 sg13g2_decap_8 FILLER_21_783 ();
 sg13g2_decap_8 FILLER_21_790 ();
 sg13g2_decap_8 FILLER_21_797 ();
 sg13g2_decap_8 FILLER_21_804 ();
 sg13g2_decap_8 FILLER_21_811 ();
 sg13g2_decap_8 FILLER_21_818 ();
 sg13g2_decap_8 FILLER_21_825 ();
 sg13g2_decap_8 FILLER_21_832 ();
 sg13g2_decap_8 FILLER_21_839 ();
 sg13g2_decap_8 FILLER_21_846 ();
 sg13g2_decap_8 FILLER_21_853 ();
 sg13g2_fill_2 FILLER_21_860 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_fill_2 FILLER_22_62 ();
 sg13g2_fill_2 FILLER_22_69 ();
 sg13g2_fill_1 FILLER_22_81 ();
 sg13g2_fill_2 FILLER_22_95 ();
 sg13g2_fill_2 FILLER_22_115 ();
 sg13g2_fill_1 FILLER_22_117 ();
 sg13g2_decap_8 FILLER_22_128 ();
 sg13g2_fill_2 FILLER_22_135 ();
 sg13g2_fill_2 FILLER_22_144 ();
 sg13g2_fill_1 FILLER_22_146 ();
 sg13g2_decap_4 FILLER_22_152 ();
 sg13g2_decap_4 FILLER_22_171 ();
 sg13g2_fill_1 FILLER_22_175 ();
 sg13g2_decap_4 FILLER_22_181 ();
 sg13g2_fill_2 FILLER_22_185 ();
 sg13g2_decap_4 FILLER_22_192 ();
 sg13g2_fill_2 FILLER_22_202 ();
 sg13g2_decap_8 FILLER_22_249 ();
 sg13g2_decap_8 FILLER_22_256 ();
 sg13g2_decap_4 FILLER_22_263 ();
 sg13g2_decap_8 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_decap_8 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_370 ();
 sg13g2_decap_8 FILLER_22_377 ();
 sg13g2_decap_4 FILLER_22_384 ();
 sg13g2_fill_2 FILLER_22_388 ();
 sg13g2_decap_8 FILLER_22_403 ();
 sg13g2_decap_8 FILLER_22_410 ();
 sg13g2_decap_8 FILLER_22_417 ();
 sg13g2_decap_8 FILLER_22_424 ();
 sg13g2_decap_8 FILLER_22_431 ();
 sg13g2_decap_8 FILLER_22_438 ();
 sg13g2_decap_8 FILLER_22_445 ();
 sg13g2_decap_8 FILLER_22_452 ();
 sg13g2_decap_8 FILLER_22_459 ();
 sg13g2_decap_8 FILLER_22_466 ();
 sg13g2_decap_8 FILLER_22_473 ();
 sg13g2_decap_8 FILLER_22_480 ();
 sg13g2_decap_8 FILLER_22_487 ();
 sg13g2_decap_8 FILLER_22_494 ();
 sg13g2_decap_8 FILLER_22_501 ();
 sg13g2_decap_8 FILLER_22_508 ();
 sg13g2_decap_8 FILLER_22_515 ();
 sg13g2_decap_8 FILLER_22_522 ();
 sg13g2_decap_8 FILLER_22_529 ();
 sg13g2_decap_8 FILLER_22_536 ();
 sg13g2_decap_8 FILLER_22_543 ();
 sg13g2_decap_8 FILLER_22_550 ();
 sg13g2_decap_8 FILLER_22_557 ();
 sg13g2_decap_8 FILLER_22_564 ();
 sg13g2_decap_8 FILLER_22_571 ();
 sg13g2_decap_8 FILLER_22_578 ();
 sg13g2_decap_8 FILLER_22_585 ();
 sg13g2_decap_8 FILLER_22_592 ();
 sg13g2_decap_8 FILLER_22_599 ();
 sg13g2_decap_8 FILLER_22_606 ();
 sg13g2_decap_8 FILLER_22_613 ();
 sg13g2_decap_8 FILLER_22_620 ();
 sg13g2_decap_8 FILLER_22_627 ();
 sg13g2_decap_8 FILLER_22_634 ();
 sg13g2_decap_8 FILLER_22_641 ();
 sg13g2_decap_8 FILLER_22_648 ();
 sg13g2_decap_8 FILLER_22_655 ();
 sg13g2_decap_8 FILLER_22_662 ();
 sg13g2_decap_8 FILLER_22_669 ();
 sg13g2_decap_8 FILLER_22_676 ();
 sg13g2_decap_8 FILLER_22_683 ();
 sg13g2_decap_8 FILLER_22_690 ();
 sg13g2_decap_8 FILLER_22_697 ();
 sg13g2_decap_8 FILLER_22_704 ();
 sg13g2_decap_8 FILLER_22_711 ();
 sg13g2_decap_8 FILLER_22_718 ();
 sg13g2_decap_8 FILLER_22_725 ();
 sg13g2_decap_8 FILLER_22_732 ();
 sg13g2_decap_8 FILLER_22_739 ();
 sg13g2_decap_8 FILLER_22_746 ();
 sg13g2_decap_8 FILLER_22_753 ();
 sg13g2_decap_8 FILLER_22_760 ();
 sg13g2_decap_8 FILLER_22_767 ();
 sg13g2_decap_8 FILLER_22_774 ();
 sg13g2_decap_8 FILLER_22_781 ();
 sg13g2_decap_8 FILLER_22_788 ();
 sg13g2_decap_8 FILLER_22_795 ();
 sg13g2_decap_8 FILLER_22_802 ();
 sg13g2_decap_8 FILLER_22_809 ();
 sg13g2_decap_8 FILLER_22_816 ();
 sg13g2_decap_8 FILLER_22_823 ();
 sg13g2_decap_8 FILLER_22_830 ();
 sg13g2_decap_8 FILLER_22_837 ();
 sg13g2_decap_8 FILLER_22_844 ();
 sg13g2_decap_8 FILLER_22_851 ();
 sg13g2_decap_4 FILLER_22_858 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_4 FILLER_23_35 ();
 sg13g2_fill_2 FILLER_23_49 ();
 sg13g2_fill_1 FILLER_23_57 ();
 sg13g2_fill_1 FILLER_23_89 ();
 sg13g2_decap_8 FILLER_23_95 ();
 sg13g2_decap_8 FILLER_23_102 ();
 sg13g2_decap_4 FILLER_23_109 ();
 sg13g2_decap_8 FILLER_23_118 ();
 sg13g2_decap_8 FILLER_23_125 ();
 sg13g2_fill_2 FILLER_23_132 ();
 sg13g2_fill_1 FILLER_23_134 ();
 sg13g2_decap_8 FILLER_23_152 ();
 sg13g2_fill_2 FILLER_23_159 ();
 sg13g2_fill_1 FILLER_23_161 ();
 sg13g2_fill_1 FILLER_23_166 ();
 sg13g2_decap_4 FILLER_23_172 ();
 sg13g2_decap_4 FILLER_23_197 ();
 sg13g2_decap_4 FILLER_23_206 ();
 sg13g2_decap_8 FILLER_23_214 ();
 sg13g2_fill_2 FILLER_23_221 ();
 sg13g2_fill_2 FILLER_23_232 ();
 sg13g2_fill_2 FILLER_23_288 ();
 sg13g2_fill_2 FILLER_23_308 ();
 sg13g2_fill_2 FILLER_23_332 ();
 sg13g2_fill_1 FILLER_23_334 ();
 sg13g2_fill_1 FILLER_23_340 ();
 sg13g2_decap_4 FILLER_23_367 ();
 sg13g2_fill_2 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_377 ();
 sg13g2_fill_2 FILLER_23_384 ();
 sg13g2_decap_8 FILLER_23_412 ();
 sg13g2_decap_8 FILLER_23_419 ();
 sg13g2_decap_8 FILLER_23_426 ();
 sg13g2_decap_8 FILLER_23_433 ();
 sg13g2_decap_8 FILLER_23_440 ();
 sg13g2_decap_8 FILLER_23_447 ();
 sg13g2_decap_8 FILLER_23_454 ();
 sg13g2_decap_8 FILLER_23_461 ();
 sg13g2_decap_8 FILLER_23_468 ();
 sg13g2_decap_8 FILLER_23_475 ();
 sg13g2_decap_8 FILLER_23_482 ();
 sg13g2_decap_8 FILLER_23_489 ();
 sg13g2_decap_8 FILLER_23_496 ();
 sg13g2_decap_8 FILLER_23_503 ();
 sg13g2_decap_8 FILLER_23_510 ();
 sg13g2_decap_8 FILLER_23_517 ();
 sg13g2_decap_8 FILLER_23_524 ();
 sg13g2_decap_8 FILLER_23_531 ();
 sg13g2_decap_8 FILLER_23_538 ();
 sg13g2_decap_8 FILLER_23_545 ();
 sg13g2_decap_8 FILLER_23_552 ();
 sg13g2_decap_8 FILLER_23_559 ();
 sg13g2_decap_8 FILLER_23_566 ();
 sg13g2_decap_8 FILLER_23_573 ();
 sg13g2_decap_8 FILLER_23_580 ();
 sg13g2_decap_8 FILLER_23_587 ();
 sg13g2_decap_8 FILLER_23_594 ();
 sg13g2_decap_8 FILLER_23_601 ();
 sg13g2_decap_8 FILLER_23_608 ();
 sg13g2_decap_8 FILLER_23_615 ();
 sg13g2_decap_8 FILLER_23_622 ();
 sg13g2_decap_8 FILLER_23_629 ();
 sg13g2_decap_8 FILLER_23_636 ();
 sg13g2_decap_8 FILLER_23_643 ();
 sg13g2_decap_8 FILLER_23_650 ();
 sg13g2_decap_8 FILLER_23_657 ();
 sg13g2_decap_8 FILLER_23_664 ();
 sg13g2_decap_8 FILLER_23_671 ();
 sg13g2_decap_8 FILLER_23_678 ();
 sg13g2_decap_8 FILLER_23_685 ();
 sg13g2_decap_8 FILLER_23_692 ();
 sg13g2_decap_8 FILLER_23_699 ();
 sg13g2_decap_8 FILLER_23_706 ();
 sg13g2_decap_8 FILLER_23_713 ();
 sg13g2_decap_8 FILLER_23_720 ();
 sg13g2_decap_8 FILLER_23_727 ();
 sg13g2_decap_8 FILLER_23_734 ();
 sg13g2_decap_8 FILLER_23_741 ();
 sg13g2_decap_8 FILLER_23_748 ();
 sg13g2_decap_8 FILLER_23_755 ();
 sg13g2_decap_8 FILLER_23_762 ();
 sg13g2_decap_8 FILLER_23_769 ();
 sg13g2_decap_8 FILLER_23_776 ();
 sg13g2_decap_8 FILLER_23_783 ();
 sg13g2_decap_8 FILLER_23_790 ();
 sg13g2_decap_8 FILLER_23_797 ();
 sg13g2_decap_8 FILLER_23_804 ();
 sg13g2_decap_8 FILLER_23_811 ();
 sg13g2_decap_8 FILLER_23_818 ();
 sg13g2_decap_8 FILLER_23_825 ();
 sg13g2_decap_8 FILLER_23_832 ();
 sg13g2_decap_8 FILLER_23_839 ();
 sg13g2_decap_8 FILLER_23_846 ();
 sg13g2_decap_8 FILLER_23_853 ();
 sg13g2_fill_2 FILLER_23_860 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_21 ();
 sg13g2_fill_1 FILLER_24_23 ();
 sg13g2_decap_4 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_32 ();
 sg13g2_fill_2 FILLER_24_46 ();
 sg13g2_decap_4 FILLER_24_53 ();
 sg13g2_fill_1 FILLER_24_66 ();
 sg13g2_decap_4 FILLER_24_77 ();
 sg13g2_fill_1 FILLER_24_81 ();
 sg13g2_decap_8 FILLER_24_87 ();
 sg13g2_decap_8 FILLER_24_94 ();
 sg13g2_decap_4 FILLER_24_117 ();
 sg13g2_decap_4 FILLER_24_129 ();
 sg13g2_fill_1 FILLER_24_133 ();
 sg13g2_fill_2 FILLER_24_150 ();
 sg13g2_fill_2 FILLER_24_174 ();
 sg13g2_fill_1 FILLER_24_176 ();
 sg13g2_decap_4 FILLER_24_181 ();
 sg13g2_fill_2 FILLER_24_224 ();
 sg13g2_fill_1 FILLER_24_251 ();
 sg13g2_fill_1 FILLER_24_292 ();
 sg13g2_fill_1 FILLER_24_315 ();
 sg13g2_fill_2 FILLER_24_321 ();
 sg13g2_fill_2 FILLER_24_344 ();
 sg13g2_fill_2 FILLER_24_359 ();
 sg13g2_fill_1 FILLER_24_361 ();
 sg13g2_fill_2 FILLER_24_404 ();
 sg13g2_decap_4 FILLER_24_441 ();
 sg13g2_fill_1 FILLER_24_445 ();
 sg13g2_decap_8 FILLER_24_450 ();
 sg13g2_decap_8 FILLER_24_457 ();
 sg13g2_decap_8 FILLER_24_464 ();
 sg13g2_decap_8 FILLER_24_471 ();
 sg13g2_decap_8 FILLER_24_478 ();
 sg13g2_decap_8 FILLER_24_485 ();
 sg13g2_decap_8 FILLER_24_492 ();
 sg13g2_decap_8 FILLER_24_499 ();
 sg13g2_decap_8 FILLER_24_506 ();
 sg13g2_decap_8 FILLER_24_513 ();
 sg13g2_decap_8 FILLER_24_520 ();
 sg13g2_decap_8 FILLER_24_527 ();
 sg13g2_decap_8 FILLER_24_534 ();
 sg13g2_decap_8 FILLER_24_541 ();
 sg13g2_decap_8 FILLER_24_548 ();
 sg13g2_decap_8 FILLER_24_555 ();
 sg13g2_decap_8 FILLER_24_562 ();
 sg13g2_decap_8 FILLER_24_569 ();
 sg13g2_decap_8 FILLER_24_576 ();
 sg13g2_decap_8 FILLER_24_583 ();
 sg13g2_decap_8 FILLER_24_590 ();
 sg13g2_decap_8 FILLER_24_597 ();
 sg13g2_decap_8 FILLER_24_604 ();
 sg13g2_decap_8 FILLER_24_611 ();
 sg13g2_decap_8 FILLER_24_618 ();
 sg13g2_decap_8 FILLER_24_625 ();
 sg13g2_decap_8 FILLER_24_632 ();
 sg13g2_decap_8 FILLER_24_639 ();
 sg13g2_decap_8 FILLER_24_646 ();
 sg13g2_decap_8 FILLER_24_653 ();
 sg13g2_decap_8 FILLER_24_660 ();
 sg13g2_decap_8 FILLER_24_667 ();
 sg13g2_decap_8 FILLER_24_674 ();
 sg13g2_decap_8 FILLER_24_681 ();
 sg13g2_decap_8 FILLER_24_688 ();
 sg13g2_decap_8 FILLER_24_695 ();
 sg13g2_decap_8 FILLER_24_702 ();
 sg13g2_decap_8 FILLER_24_709 ();
 sg13g2_decap_8 FILLER_24_716 ();
 sg13g2_decap_8 FILLER_24_723 ();
 sg13g2_decap_8 FILLER_24_730 ();
 sg13g2_decap_8 FILLER_24_737 ();
 sg13g2_decap_8 FILLER_24_744 ();
 sg13g2_decap_8 FILLER_24_751 ();
 sg13g2_decap_8 FILLER_24_758 ();
 sg13g2_decap_8 FILLER_24_765 ();
 sg13g2_decap_8 FILLER_24_772 ();
 sg13g2_decap_8 FILLER_24_779 ();
 sg13g2_decap_8 FILLER_24_786 ();
 sg13g2_decap_8 FILLER_24_793 ();
 sg13g2_decap_8 FILLER_24_800 ();
 sg13g2_decap_8 FILLER_24_807 ();
 sg13g2_decap_8 FILLER_24_814 ();
 sg13g2_decap_8 FILLER_24_821 ();
 sg13g2_decap_8 FILLER_24_828 ();
 sg13g2_decap_8 FILLER_24_835 ();
 sg13g2_decap_8 FILLER_24_842 ();
 sg13g2_decap_8 FILLER_24_849 ();
 sg13g2_decap_4 FILLER_24_856 ();
 sg13g2_fill_2 FILLER_24_860 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_fill_2 FILLER_25_11 ();
 sg13g2_decap_8 FILLER_25_60 ();
 sg13g2_decap_4 FILLER_25_91 ();
 sg13g2_fill_1 FILLER_25_95 ();
 sg13g2_fill_1 FILLER_25_122 ();
 sg13g2_fill_2 FILLER_25_164 ();
 sg13g2_fill_1 FILLER_25_166 ();
 sg13g2_fill_2 FILLER_25_177 ();
 sg13g2_fill_2 FILLER_25_205 ();
 sg13g2_fill_2 FILLER_25_217 ();
 sg13g2_decap_4 FILLER_25_250 ();
 sg13g2_fill_1 FILLER_25_254 ();
 sg13g2_fill_2 FILLER_25_269 ();
 sg13g2_fill_2 FILLER_25_279 ();
 sg13g2_fill_1 FILLER_25_316 ();
 sg13g2_fill_1 FILLER_25_343 ();
 sg13g2_fill_2 FILLER_25_373 ();
 sg13g2_fill_2 FILLER_25_399 ();
 sg13g2_fill_1 FILLER_25_434 ();
 sg13g2_decap_4 FILLER_25_461 ();
 sg13g2_fill_1 FILLER_25_465 ();
 sg13g2_decap_8 FILLER_25_469 ();
 sg13g2_decap_8 FILLER_25_476 ();
 sg13g2_decap_8 FILLER_25_483 ();
 sg13g2_decap_8 FILLER_25_490 ();
 sg13g2_decap_8 FILLER_25_497 ();
 sg13g2_decap_8 FILLER_25_504 ();
 sg13g2_decap_8 FILLER_25_511 ();
 sg13g2_decap_8 FILLER_25_518 ();
 sg13g2_decap_8 FILLER_25_525 ();
 sg13g2_decap_8 FILLER_25_532 ();
 sg13g2_decap_8 FILLER_25_539 ();
 sg13g2_decap_8 FILLER_25_546 ();
 sg13g2_decap_8 FILLER_25_553 ();
 sg13g2_decap_8 FILLER_25_560 ();
 sg13g2_decap_8 FILLER_25_567 ();
 sg13g2_decap_8 FILLER_25_574 ();
 sg13g2_decap_8 FILLER_25_581 ();
 sg13g2_decap_8 FILLER_25_588 ();
 sg13g2_decap_8 FILLER_25_595 ();
 sg13g2_decap_8 FILLER_25_602 ();
 sg13g2_decap_8 FILLER_25_609 ();
 sg13g2_decap_8 FILLER_25_616 ();
 sg13g2_decap_8 FILLER_25_623 ();
 sg13g2_decap_8 FILLER_25_630 ();
 sg13g2_decap_8 FILLER_25_637 ();
 sg13g2_decap_8 FILLER_25_644 ();
 sg13g2_decap_8 FILLER_25_651 ();
 sg13g2_decap_8 FILLER_25_658 ();
 sg13g2_decap_8 FILLER_25_665 ();
 sg13g2_decap_8 FILLER_25_672 ();
 sg13g2_decap_8 FILLER_25_679 ();
 sg13g2_decap_8 FILLER_25_686 ();
 sg13g2_decap_8 FILLER_25_693 ();
 sg13g2_decap_8 FILLER_25_700 ();
 sg13g2_decap_8 FILLER_25_707 ();
 sg13g2_decap_8 FILLER_25_714 ();
 sg13g2_decap_8 FILLER_25_721 ();
 sg13g2_decap_8 FILLER_25_728 ();
 sg13g2_decap_8 FILLER_25_735 ();
 sg13g2_decap_8 FILLER_25_742 ();
 sg13g2_decap_8 FILLER_25_749 ();
 sg13g2_decap_8 FILLER_25_756 ();
 sg13g2_decap_8 FILLER_25_763 ();
 sg13g2_decap_8 FILLER_25_770 ();
 sg13g2_decap_8 FILLER_25_777 ();
 sg13g2_decap_8 FILLER_25_784 ();
 sg13g2_decap_8 FILLER_25_791 ();
 sg13g2_decap_8 FILLER_25_798 ();
 sg13g2_decap_8 FILLER_25_805 ();
 sg13g2_decap_8 FILLER_25_812 ();
 sg13g2_decap_8 FILLER_25_819 ();
 sg13g2_decap_8 FILLER_25_826 ();
 sg13g2_decap_8 FILLER_25_833 ();
 sg13g2_decap_8 FILLER_25_840 ();
 sg13g2_decap_8 FILLER_25_847 ();
 sg13g2_decap_8 FILLER_25_854 ();
 sg13g2_fill_1 FILLER_25_861 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_4 ();
 sg13g2_fill_1 FILLER_26_32 ();
 sg13g2_fill_2 FILLER_26_63 ();
 sg13g2_fill_1 FILLER_26_65 ();
 sg13g2_decap_4 FILLER_26_94 ();
 sg13g2_fill_1 FILLER_26_98 ();
 sg13g2_fill_1 FILLER_26_123 ();
 sg13g2_fill_2 FILLER_26_128 ();
 sg13g2_fill_1 FILLER_26_136 ();
 sg13g2_fill_2 FILLER_26_142 ();
 sg13g2_fill_1 FILLER_26_144 ();
 sg13g2_fill_1 FILLER_26_154 ();
 sg13g2_fill_1 FILLER_26_159 ();
 sg13g2_fill_1 FILLER_26_173 ();
 sg13g2_fill_2 FILLER_26_179 ();
 sg13g2_fill_2 FILLER_26_186 ();
 sg13g2_fill_1 FILLER_26_188 ();
 sg13g2_fill_1 FILLER_26_203 ();
 sg13g2_decap_4 FILLER_26_235 ();
 sg13g2_fill_2 FILLER_26_239 ();
 sg13g2_decap_8 FILLER_26_275 ();
 sg13g2_decap_4 FILLER_26_282 ();
 sg13g2_fill_2 FILLER_26_286 ();
 sg13g2_fill_2 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_fill_2 FILLER_26_329 ();
 sg13g2_decap_8 FILLER_26_345 ();
 sg13g2_fill_1 FILLER_26_380 ();
 sg13g2_decap_4 FILLER_26_417 ();
 sg13g2_fill_1 FILLER_26_421 ();
 sg13g2_fill_1 FILLER_26_466 ();
 sg13g2_decap_8 FILLER_26_476 ();
 sg13g2_decap_8 FILLER_26_483 ();
 sg13g2_decap_8 FILLER_26_490 ();
 sg13g2_decap_8 FILLER_26_497 ();
 sg13g2_decap_8 FILLER_26_504 ();
 sg13g2_decap_8 FILLER_26_511 ();
 sg13g2_decap_8 FILLER_26_518 ();
 sg13g2_decap_8 FILLER_26_525 ();
 sg13g2_decap_8 FILLER_26_532 ();
 sg13g2_decap_8 FILLER_26_539 ();
 sg13g2_decap_8 FILLER_26_546 ();
 sg13g2_decap_8 FILLER_26_553 ();
 sg13g2_decap_8 FILLER_26_560 ();
 sg13g2_decap_8 FILLER_26_567 ();
 sg13g2_decap_8 FILLER_26_574 ();
 sg13g2_decap_8 FILLER_26_581 ();
 sg13g2_decap_8 FILLER_26_588 ();
 sg13g2_decap_8 FILLER_26_595 ();
 sg13g2_decap_8 FILLER_26_602 ();
 sg13g2_decap_8 FILLER_26_609 ();
 sg13g2_decap_8 FILLER_26_616 ();
 sg13g2_decap_8 FILLER_26_623 ();
 sg13g2_decap_8 FILLER_26_630 ();
 sg13g2_decap_8 FILLER_26_637 ();
 sg13g2_decap_8 FILLER_26_644 ();
 sg13g2_decap_8 FILLER_26_651 ();
 sg13g2_decap_8 FILLER_26_658 ();
 sg13g2_decap_8 FILLER_26_665 ();
 sg13g2_decap_8 FILLER_26_672 ();
 sg13g2_decap_8 FILLER_26_679 ();
 sg13g2_decap_8 FILLER_26_686 ();
 sg13g2_decap_8 FILLER_26_693 ();
 sg13g2_decap_8 FILLER_26_700 ();
 sg13g2_decap_8 FILLER_26_707 ();
 sg13g2_decap_8 FILLER_26_714 ();
 sg13g2_decap_8 FILLER_26_721 ();
 sg13g2_decap_8 FILLER_26_728 ();
 sg13g2_decap_8 FILLER_26_735 ();
 sg13g2_decap_8 FILLER_26_742 ();
 sg13g2_decap_8 FILLER_26_749 ();
 sg13g2_decap_8 FILLER_26_756 ();
 sg13g2_decap_8 FILLER_26_763 ();
 sg13g2_decap_8 FILLER_26_770 ();
 sg13g2_decap_8 FILLER_26_777 ();
 sg13g2_decap_8 FILLER_26_784 ();
 sg13g2_decap_8 FILLER_26_791 ();
 sg13g2_decap_8 FILLER_26_798 ();
 sg13g2_decap_8 FILLER_26_805 ();
 sg13g2_decap_8 FILLER_26_812 ();
 sg13g2_decap_8 FILLER_26_819 ();
 sg13g2_decap_8 FILLER_26_826 ();
 sg13g2_decap_8 FILLER_26_833 ();
 sg13g2_decap_8 FILLER_26_840 ();
 sg13g2_decap_8 FILLER_26_847 ();
 sg13g2_decap_8 FILLER_26_854 ();
 sg13g2_fill_1 FILLER_26_861 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_31 ();
 sg13g2_fill_2 FILLER_27_47 ();
 sg13g2_decap_8 FILLER_27_57 ();
 sg13g2_decap_8 FILLER_27_64 ();
 sg13g2_decap_8 FILLER_27_71 ();
 sg13g2_fill_1 FILLER_27_78 ();
 sg13g2_fill_2 FILLER_27_91 ();
 sg13g2_decap_4 FILLER_27_120 ();
 sg13g2_fill_1 FILLER_27_124 ();
 sg13g2_fill_2 FILLER_27_130 ();
 sg13g2_fill_2 FILLER_27_136 ();
 sg13g2_fill_1 FILLER_27_138 ();
 sg13g2_fill_2 FILLER_27_177 ();
 sg13g2_fill_1 FILLER_27_248 ();
 sg13g2_decap_4 FILLER_27_282 ();
 sg13g2_decap_8 FILLER_27_291 ();
 sg13g2_decap_4 FILLER_27_298 ();
 sg13g2_fill_2 FILLER_27_302 ();
 sg13g2_fill_2 FILLER_27_314 ();
 sg13g2_decap_4 FILLER_27_342 ();
 sg13g2_fill_1 FILLER_27_346 ();
 sg13g2_fill_1 FILLER_27_405 ();
 sg13g2_decap_4 FILLER_27_442 ();
 sg13g2_fill_2 FILLER_27_446 ();
 sg13g2_fill_2 FILLER_27_456 ();
 sg13g2_fill_1 FILLER_27_458 ();
 sg13g2_fill_1 FILLER_27_464 ();
 sg13g2_decap_8 FILLER_27_482 ();
 sg13g2_decap_4 FILLER_27_489 ();
 sg13g2_decap_8 FILLER_27_496 ();
 sg13g2_decap_8 FILLER_27_503 ();
 sg13g2_decap_8 FILLER_27_510 ();
 sg13g2_decap_8 FILLER_27_517 ();
 sg13g2_decap_8 FILLER_27_524 ();
 sg13g2_decap_8 FILLER_27_531 ();
 sg13g2_decap_8 FILLER_27_538 ();
 sg13g2_decap_8 FILLER_27_545 ();
 sg13g2_decap_8 FILLER_27_552 ();
 sg13g2_decap_8 FILLER_27_559 ();
 sg13g2_decap_8 FILLER_27_566 ();
 sg13g2_decap_8 FILLER_27_573 ();
 sg13g2_decap_8 FILLER_27_580 ();
 sg13g2_decap_8 FILLER_27_587 ();
 sg13g2_decap_8 FILLER_27_594 ();
 sg13g2_decap_8 FILLER_27_601 ();
 sg13g2_decap_8 FILLER_27_608 ();
 sg13g2_decap_8 FILLER_27_615 ();
 sg13g2_decap_8 FILLER_27_622 ();
 sg13g2_decap_8 FILLER_27_629 ();
 sg13g2_decap_8 FILLER_27_636 ();
 sg13g2_decap_8 FILLER_27_643 ();
 sg13g2_decap_8 FILLER_27_650 ();
 sg13g2_decap_8 FILLER_27_657 ();
 sg13g2_decap_8 FILLER_27_664 ();
 sg13g2_decap_8 FILLER_27_671 ();
 sg13g2_decap_8 FILLER_27_678 ();
 sg13g2_decap_8 FILLER_27_685 ();
 sg13g2_decap_8 FILLER_27_692 ();
 sg13g2_decap_8 FILLER_27_699 ();
 sg13g2_decap_8 FILLER_27_706 ();
 sg13g2_decap_8 FILLER_27_713 ();
 sg13g2_decap_8 FILLER_27_720 ();
 sg13g2_decap_8 FILLER_27_727 ();
 sg13g2_decap_8 FILLER_27_734 ();
 sg13g2_decap_8 FILLER_27_741 ();
 sg13g2_decap_8 FILLER_27_748 ();
 sg13g2_decap_8 FILLER_27_755 ();
 sg13g2_decap_8 FILLER_27_762 ();
 sg13g2_decap_8 FILLER_27_769 ();
 sg13g2_decap_8 FILLER_27_776 ();
 sg13g2_decap_8 FILLER_27_783 ();
 sg13g2_decap_8 FILLER_27_790 ();
 sg13g2_decap_8 FILLER_27_797 ();
 sg13g2_decap_8 FILLER_27_804 ();
 sg13g2_decap_8 FILLER_27_811 ();
 sg13g2_decap_8 FILLER_27_818 ();
 sg13g2_decap_8 FILLER_27_825 ();
 sg13g2_decap_8 FILLER_27_832 ();
 sg13g2_decap_8 FILLER_27_839 ();
 sg13g2_decap_8 FILLER_27_846 ();
 sg13g2_decap_8 FILLER_27_853 ();
 sg13g2_fill_2 FILLER_27_860 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_14 ();
 sg13g2_fill_2 FILLER_28_81 ();
 sg13g2_fill_1 FILLER_28_83 ();
 sg13g2_decap_8 FILLER_28_92 ();
 sg13g2_fill_2 FILLER_28_99 ();
 sg13g2_decap_4 FILLER_28_113 ();
 sg13g2_fill_1 FILLER_28_152 ();
 sg13g2_fill_1 FILLER_28_157 ();
 sg13g2_fill_2 FILLER_28_178 ();
 sg13g2_fill_1 FILLER_28_180 ();
 sg13g2_fill_2 FILLER_28_186 ();
 sg13g2_fill_1 FILLER_28_207 ();
 sg13g2_fill_1 FILLER_28_227 ();
 sg13g2_decap_4 FILLER_28_254 ();
 sg13g2_fill_2 FILLER_28_355 ();
 sg13g2_fill_2 FILLER_28_378 ();
 sg13g2_fill_2 FILLER_28_460 ();
 sg13g2_fill_1 FILLER_28_493 ();
 sg13g2_decap_8 FILLER_28_503 ();
 sg13g2_decap_8 FILLER_28_510 ();
 sg13g2_decap_8 FILLER_28_517 ();
 sg13g2_decap_8 FILLER_28_524 ();
 sg13g2_decap_8 FILLER_28_531 ();
 sg13g2_decap_8 FILLER_28_538 ();
 sg13g2_decap_8 FILLER_28_545 ();
 sg13g2_decap_8 FILLER_28_552 ();
 sg13g2_decap_8 FILLER_28_559 ();
 sg13g2_decap_8 FILLER_28_566 ();
 sg13g2_decap_8 FILLER_28_573 ();
 sg13g2_decap_8 FILLER_28_580 ();
 sg13g2_decap_8 FILLER_28_587 ();
 sg13g2_decap_8 FILLER_28_594 ();
 sg13g2_decap_8 FILLER_28_601 ();
 sg13g2_decap_8 FILLER_28_608 ();
 sg13g2_decap_8 FILLER_28_615 ();
 sg13g2_decap_8 FILLER_28_622 ();
 sg13g2_decap_8 FILLER_28_629 ();
 sg13g2_decap_8 FILLER_28_636 ();
 sg13g2_decap_8 FILLER_28_643 ();
 sg13g2_decap_8 FILLER_28_650 ();
 sg13g2_decap_8 FILLER_28_657 ();
 sg13g2_decap_8 FILLER_28_664 ();
 sg13g2_decap_8 FILLER_28_671 ();
 sg13g2_decap_8 FILLER_28_678 ();
 sg13g2_decap_8 FILLER_28_685 ();
 sg13g2_decap_8 FILLER_28_692 ();
 sg13g2_decap_8 FILLER_28_699 ();
 sg13g2_decap_8 FILLER_28_706 ();
 sg13g2_decap_8 FILLER_28_713 ();
 sg13g2_decap_8 FILLER_28_720 ();
 sg13g2_decap_8 FILLER_28_727 ();
 sg13g2_decap_8 FILLER_28_734 ();
 sg13g2_decap_8 FILLER_28_741 ();
 sg13g2_decap_8 FILLER_28_748 ();
 sg13g2_decap_8 FILLER_28_755 ();
 sg13g2_decap_8 FILLER_28_762 ();
 sg13g2_decap_8 FILLER_28_769 ();
 sg13g2_decap_8 FILLER_28_776 ();
 sg13g2_decap_8 FILLER_28_783 ();
 sg13g2_decap_8 FILLER_28_790 ();
 sg13g2_decap_8 FILLER_28_797 ();
 sg13g2_decap_8 FILLER_28_804 ();
 sg13g2_decap_8 FILLER_28_811 ();
 sg13g2_decap_8 FILLER_28_818 ();
 sg13g2_decap_8 FILLER_28_825 ();
 sg13g2_decap_8 FILLER_28_832 ();
 sg13g2_decap_8 FILLER_28_839 ();
 sg13g2_decap_8 FILLER_28_846 ();
 sg13g2_decap_8 FILLER_28_853 ();
 sg13g2_fill_2 FILLER_28_860 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_9 ();
 sg13g2_fill_1 FILLER_29_36 ();
 sg13g2_fill_2 FILLER_29_41 ();
 sg13g2_fill_1 FILLER_29_43 ();
 sg13g2_fill_1 FILLER_29_53 ();
 sg13g2_fill_2 FILLER_29_64 ();
 sg13g2_fill_2 FILLER_29_79 ();
 sg13g2_decap_8 FILLER_29_104 ();
 sg13g2_fill_2 FILLER_29_111 ();
 sg13g2_fill_1 FILLER_29_127 ();
 sg13g2_decap_8 FILLER_29_135 ();
 sg13g2_fill_2 FILLER_29_264 ();
 sg13g2_fill_1 FILLER_29_266 ();
 sg13g2_fill_2 FILLER_29_272 ();
 sg13g2_fill_2 FILLER_29_292 ();
 sg13g2_fill_1 FILLER_29_294 ();
 sg13g2_decap_4 FILLER_29_299 ();
 sg13g2_fill_2 FILLER_29_335 ();
 sg13g2_decap_4 FILLER_29_347 ();
 sg13g2_fill_1 FILLER_29_361 ();
 sg13g2_decap_8 FILLER_29_383 ();
 sg13g2_fill_1 FILLER_29_390 ();
 sg13g2_decap_8 FILLER_29_395 ();
 sg13g2_fill_2 FILLER_29_413 ();
 sg13g2_decap_8 FILLER_29_503 ();
 sg13g2_decap_8 FILLER_29_510 ();
 sg13g2_decap_8 FILLER_29_517 ();
 sg13g2_decap_8 FILLER_29_524 ();
 sg13g2_decap_8 FILLER_29_531 ();
 sg13g2_decap_8 FILLER_29_538 ();
 sg13g2_decap_8 FILLER_29_545 ();
 sg13g2_decap_8 FILLER_29_552 ();
 sg13g2_decap_8 FILLER_29_559 ();
 sg13g2_decap_8 FILLER_29_566 ();
 sg13g2_decap_8 FILLER_29_573 ();
 sg13g2_decap_8 FILLER_29_580 ();
 sg13g2_decap_8 FILLER_29_587 ();
 sg13g2_decap_8 FILLER_29_594 ();
 sg13g2_decap_8 FILLER_29_601 ();
 sg13g2_decap_8 FILLER_29_608 ();
 sg13g2_decap_8 FILLER_29_615 ();
 sg13g2_decap_8 FILLER_29_622 ();
 sg13g2_decap_8 FILLER_29_629 ();
 sg13g2_decap_8 FILLER_29_636 ();
 sg13g2_decap_8 FILLER_29_643 ();
 sg13g2_decap_8 FILLER_29_650 ();
 sg13g2_decap_8 FILLER_29_657 ();
 sg13g2_decap_8 FILLER_29_664 ();
 sg13g2_decap_8 FILLER_29_671 ();
 sg13g2_decap_8 FILLER_29_678 ();
 sg13g2_decap_8 FILLER_29_685 ();
 sg13g2_decap_8 FILLER_29_692 ();
 sg13g2_decap_8 FILLER_29_699 ();
 sg13g2_decap_8 FILLER_29_706 ();
 sg13g2_decap_8 FILLER_29_713 ();
 sg13g2_decap_8 FILLER_29_720 ();
 sg13g2_decap_8 FILLER_29_727 ();
 sg13g2_decap_8 FILLER_29_734 ();
 sg13g2_decap_8 FILLER_29_741 ();
 sg13g2_decap_8 FILLER_29_748 ();
 sg13g2_decap_8 FILLER_29_755 ();
 sg13g2_decap_8 FILLER_29_762 ();
 sg13g2_decap_8 FILLER_29_769 ();
 sg13g2_decap_8 FILLER_29_776 ();
 sg13g2_decap_8 FILLER_29_783 ();
 sg13g2_decap_8 FILLER_29_790 ();
 sg13g2_decap_8 FILLER_29_797 ();
 sg13g2_decap_8 FILLER_29_804 ();
 sg13g2_decap_8 FILLER_29_811 ();
 sg13g2_decap_8 FILLER_29_818 ();
 sg13g2_decap_8 FILLER_29_825 ();
 sg13g2_decap_8 FILLER_29_832 ();
 sg13g2_decap_8 FILLER_29_839 ();
 sg13g2_decap_8 FILLER_29_846 ();
 sg13g2_decap_8 FILLER_29_853 ();
 sg13g2_fill_2 FILLER_29_860 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_fill_1 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_47 ();
 sg13g2_decap_4 FILLER_30_54 ();
 sg13g2_fill_1 FILLER_30_85 ();
 sg13g2_fill_2 FILLER_30_102 ();
 sg13g2_fill_1 FILLER_30_104 ();
 sg13g2_fill_2 FILLER_30_131 ();
 sg13g2_fill_1 FILLER_30_159 ();
 sg13g2_fill_1 FILLER_30_182 ();
 sg13g2_fill_1 FILLER_30_196 ();
 sg13g2_fill_2 FILLER_30_219 ();
 sg13g2_fill_1 FILLER_30_235 ();
 sg13g2_fill_2 FILLER_30_245 ();
 sg13g2_fill_1 FILLER_30_247 ();
 sg13g2_fill_1 FILLER_30_254 ();
 sg13g2_fill_2 FILLER_30_264 ();
 sg13g2_decap_8 FILLER_30_288 ();
 sg13g2_decap_8 FILLER_30_295 ();
 sg13g2_fill_2 FILLER_30_348 ();
 sg13g2_fill_1 FILLER_30_350 ();
 sg13g2_fill_2 FILLER_30_361 ();
 sg13g2_fill_1 FILLER_30_363 ();
 sg13g2_decap_8 FILLER_30_396 ();
 sg13g2_fill_2 FILLER_30_403 ();
 sg13g2_fill_1 FILLER_30_423 ();
 sg13g2_decap_4 FILLER_30_442 ();
 sg13g2_fill_1 FILLER_30_446 ();
 sg13g2_decap_4 FILLER_30_456 ();
 sg13g2_decap_8 FILLER_30_501 ();
 sg13g2_decap_8 FILLER_30_508 ();
 sg13g2_decap_8 FILLER_30_515 ();
 sg13g2_decap_8 FILLER_30_522 ();
 sg13g2_decap_8 FILLER_30_529 ();
 sg13g2_decap_8 FILLER_30_536 ();
 sg13g2_decap_8 FILLER_30_543 ();
 sg13g2_decap_8 FILLER_30_550 ();
 sg13g2_decap_8 FILLER_30_557 ();
 sg13g2_decap_8 FILLER_30_564 ();
 sg13g2_decap_8 FILLER_30_571 ();
 sg13g2_decap_8 FILLER_30_578 ();
 sg13g2_decap_8 FILLER_30_585 ();
 sg13g2_decap_8 FILLER_30_592 ();
 sg13g2_decap_8 FILLER_30_599 ();
 sg13g2_decap_8 FILLER_30_606 ();
 sg13g2_decap_8 FILLER_30_613 ();
 sg13g2_decap_8 FILLER_30_620 ();
 sg13g2_decap_8 FILLER_30_627 ();
 sg13g2_decap_8 FILLER_30_634 ();
 sg13g2_decap_8 FILLER_30_641 ();
 sg13g2_decap_8 FILLER_30_648 ();
 sg13g2_decap_8 FILLER_30_655 ();
 sg13g2_decap_8 FILLER_30_662 ();
 sg13g2_decap_8 FILLER_30_669 ();
 sg13g2_decap_8 FILLER_30_676 ();
 sg13g2_decap_8 FILLER_30_683 ();
 sg13g2_decap_8 FILLER_30_690 ();
 sg13g2_decap_8 FILLER_30_697 ();
 sg13g2_decap_8 FILLER_30_704 ();
 sg13g2_decap_8 FILLER_30_711 ();
 sg13g2_decap_8 FILLER_30_718 ();
 sg13g2_decap_8 FILLER_30_725 ();
 sg13g2_decap_8 FILLER_30_732 ();
 sg13g2_decap_8 FILLER_30_739 ();
 sg13g2_decap_8 FILLER_30_746 ();
 sg13g2_decap_8 FILLER_30_753 ();
 sg13g2_decap_8 FILLER_30_760 ();
 sg13g2_decap_8 FILLER_30_767 ();
 sg13g2_decap_8 FILLER_30_774 ();
 sg13g2_decap_8 FILLER_30_781 ();
 sg13g2_decap_8 FILLER_30_788 ();
 sg13g2_decap_8 FILLER_30_795 ();
 sg13g2_decap_8 FILLER_30_802 ();
 sg13g2_decap_8 FILLER_30_809 ();
 sg13g2_decap_8 FILLER_30_816 ();
 sg13g2_decap_8 FILLER_30_823 ();
 sg13g2_decap_8 FILLER_30_830 ();
 sg13g2_decap_8 FILLER_30_837 ();
 sg13g2_decap_8 FILLER_30_844 ();
 sg13g2_decap_8 FILLER_30_851 ();
 sg13g2_decap_4 FILLER_30_858 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_fill_1 FILLER_31_21 ();
 sg13g2_fill_1 FILLER_31_26 ();
 sg13g2_fill_2 FILLER_31_36 ();
 sg13g2_fill_2 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_51 ();
 sg13g2_fill_1 FILLER_31_103 ();
 sg13g2_fill_1 FILLER_31_113 ();
 sg13g2_fill_1 FILLER_31_123 ();
 sg13g2_fill_2 FILLER_31_142 ();
 sg13g2_fill_1 FILLER_31_154 ();
 sg13g2_fill_1 FILLER_31_170 ();
 sg13g2_fill_1 FILLER_31_226 ();
 sg13g2_fill_2 FILLER_31_288 ();
 sg13g2_fill_1 FILLER_31_290 ();
 sg13g2_fill_2 FILLER_31_323 ();
 sg13g2_fill_1 FILLER_31_325 ();
 sg13g2_decap_4 FILLER_31_362 ();
 sg13g2_fill_1 FILLER_31_371 ();
 sg13g2_fill_2 FILLER_31_395 ();
 sg13g2_decap_8 FILLER_31_425 ();
 sg13g2_fill_1 FILLER_31_458 ();
 sg13g2_fill_2 FILLER_31_464 ();
 sg13g2_decap_8 FILLER_31_500 ();
 sg13g2_decap_8 FILLER_31_507 ();
 sg13g2_decap_8 FILLER_31_514 ();
 sg13g2_decap_8 FILLER_31_521 ();
 sg13g2_decap_8 FILLER_31_528 ();
 sg13g2_decap_8 FILLER_31_535 ();
 sg13g2_decap_8 FILLER_31_542 ();
 sg13g2_decap_8 FILLER_31_549 ();
 sg13g2_decap_8 FILLER_31_556 ();
 sg13g2_decap_8 FILLER_31_563 ();
 sg13g2_decap_8 FILLER_31_570 ();
 sg13g2_decap_8 FILLER_31_577 ();
 sg13g2_decap_8 FILLER_31_584 ();
 sg13g2_decap_8 FILLER_31_591 ();
 sg13g2_decap_8 FILLER_31_598 ();
 sg13g2_decap_8 FILLER_31_605 ();
 sg13g2_decap_8 FILLER_31_612 ();
 sg13g2_decap_8 FILLER_31_619 ();
 sg13g2_decap_8 FILLER_31_626 ();
 sg13g2_decap_8 FILLER_31_633 ();
 sg13g2_decap_8 FILLER_31_640 ();
 sg13g2_decap_8 FILLER_31_647 ();
 sg13g2_decap_8 FILLER_31_654 ();
 sg13g2_decap_8 FILLER_31_661 ();
 sg13g2_decap_8 FILLER_31_668 ();
 sg13g2_decap_8 FILLER_31_675 ();
 sg13g2_decap_8 FILLER_31_682 ();
 sg13g2_decap_8 FILLER_31_689 ();
 sg13g2_decap_8 FILLER_31_696 ();
 sg13g2_decap_8 FILLER_31_703 ();
 sg13g2_decap_8 FILLER_31_710 ();
 sg13g2_decap_8 FILLER_31_717 ();
 sg13g2_decap_8 FILLER_31_724 ();
 sg13g2_decap_8 FILLER_31_731 ();
 sg13g2_decap_8 FILLER_31_738 ();
 sg13g2_decap_8 FILLER_31_745 ();
 sg13g2_decap_8 FILLER_31_752 ();
 sg13g2_decap_8 FILLER_31_759 ();
 sg13g2_decap_8 FILLER_31_766 ();
 sg13g2_decap_8 FILLER_31_773 ();
 sg13g2_decap_8 FILLER_31_780 ();
 sg13g2_decap_8 FILLER_31_787 ();
 sg13g2_decap_8 FILLER_31_794 ();
 sg13g2_decap_8 FILLER_31_801 ();
 sg13g2_decap_8 FILLER_31_808 ();
 sg13g2_decap_8 FILLER_31_815 ();
 sg13g2_decap_8 FILLER_31_822 ();
 sg13g2_decap_8 FILLER_31_829 ();
 sg13g2_decap_8 FILLER_31_836 ();
 sg13g2_decap_8 FILLER_31_843 ();
 sg13g2_decap_8 FILLER_31_850 ();
 sg13g2_decap_4 FILLER_31_857 ();
 sg13g2_fill_1 FILLER_31_861 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_52 ();
 sg13g2_fill_2 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_88 ();
 sg13g2_fill_2 FILLER_32_95 ();
 sg13g2_fill_1 FILLER_32_97 ();
 sg13g2_fill_2 FILLER_32_128 ();
 sg13g2_fill_2 FILLER_32_160 ();
 sg13g2_decap_4 FILLER_32_195 ();
 sg13g2_fill_2 FILLER_32_209 ();
 sg13g2_fill_2 FILLER_32_215 ();
 sg13g2_fill_2 FILLER_32_242 ();
 sg13g2_fill_2 FILLER_32_264 ();
 sg13g2_fill_1 FILLER_32_285 ();
 sg13g2_fill_1 FILLER_32_296 ();
 sg13g2_fill_2 FILLER_32_310 ();
 sg13g2_fill_2 FILLER_32_322 ();
 sg13g2_decap_8 FILLER_32_345 ();
 sg13g2_fill_1 FILLER_32_352 ();
 sg13g2_decap_4 FILLER_32_376 ();
 sg13g2_decap_8 FILLER_32_398 ();
 sg13g2_decap_4 FILLER_32_405 ();
 sg13g2_fill_2 FILLER_32_409 ();
 sg13g2_decap_4 FILLER_32_416 ();
 sg13g2_fill_1 FILLER_32_420 ();
 sg13g2_decap_4 FILLER_32_433 ();
 sg13g2_fill_1 FILLER_32_437 ();
 sg13g2_fill_2 FILLER_32_455 ();
 sg13g2_fill_2 FILLER_32_488 ();
 sg13g2_decap_8 FILLER_32_506 ();
 sg13g2_decap_8 FILLER_32_513 ();
 sg13g2_decap_8 FILLER_32_520 ();
 sg13g2_decap_8 FILLER_32_527 ();
 sg13g2_decap_8 FILLER_32_534 ();
 sg13g2_decap_8 FILLER_32_541 ();
 sg13g2_decap_8 FILLER_32_548 ();
 sg13g2_decap_8 FILLER_32_555 ();
 sg13g2_decap_8 FILLER_32_562 ();
 sg13g2_decap_8 FILLER_32_569 ();
 sg13g2_decap_8 FILLER_32_576 ();
 sg13g2_decap_8 FILLER_32_583 ();
 sg13g2_decap_8 FILLER_32_590 ();
 sg13g2_decap_8 FILLER_32_597 ();
 sg13g2_decap_8 FILLER_32_604 ();
 sg13g2_decap_8 FILLER_32_611 ();
 sg13g2_decap_8 FILLER_32_618 ();
 sg13g2_decap_8 FILLER_32_625 ();
 sg13g2_decap_8 FILLER_32_632 ();
 sg13g2_decap_8 FILLER_32_639 ();
 sg13g2_decap_8 FILLER_32_646 ();
 sg13g2_decap_8 FILLER_32_653 ();
 sg13g2_decap_8 FILLER_32_660 ();
 sg13g2_decap_8 FILLER_32_667 ();
 sg13g2_decap_8 FILLER_32_674 ();
 sg13g2_decap_8 FILLER_32_681 ();
 sg13g2_decap_8 FILLER_32_688 ();
 sg13g2_decap_8 FILLER_32_695 ();
 sg13g2_decap_8 FILLER_32_702 ();
 sg13g2_decap_8 FILLER_32_709 ();
 sg13g2_decap_8 FILLER_32_716 ();
 sg13g2_decap_8 FILLER_32_723 ();
 sg13g2_decap_8 FILLER_32_730 ();
 sg13g2_decap_8 FILLER_32_737 ();
 sg13g2_decap_8 FILLER_32_744 ();
 sg13g2_decap_8 FILLER_32_751 ();
 sg13g2_decap_8 FILLER_32_758 ();
 sg13g2_decap_8 FILLER_32_765 ();
 sg13g2_decap_8 FILLER_32_772 ();
 sg13g2_decap_8 FILLER_32_779 ();
 sg13g2_decap_8 FILLER_32_786 ();
 sg13g2_decap_8 FILLER_32_793 ();
 sg13g2_decap_8 FILLER_32_800 ();
 sg13g2_decap_8 FILLER_32_807 ();
 sg13g2_decap_8 FILLER_32_814 ();
 sg13g2_decap_8 FILLER_32_821 ();
 sg13g2_decap_8 FILLER_32_828 ();
 sg13g2_decap_8 FILLER_32_835 ();
 sg13g2_decap_8 FILLER_32_842 ();
 sg13g2_decap_8 FILLER_32_849 ();
 sg13g2_decap_4 FILLER_32_856 ();
 sg13g2_fill_2 FILLER_32_860 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_15 ();
 sg13g2_fill_2 FILLER_33_25 ();
 sg13g2_fill_2 FILLER_33_74 ();
 sg13g2_fill_1 FILLER_33_76 ();
 sg13g2_fill_2 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_110 ();
 sg13g2_decap_4 FILLER_33_121 ();
 sg13g2_fill_2 FILLER_33_125 ();
 sg13g2_fill_2 FILLER_33_130 ();
 sg13g2_fill_2 FILLER_33_158 ();
 sg13g2_fill_1 FILLER_33_160 ();
 sg13g2_fill_1 FILLER_33_201 ();
 sg13g2_fill_2 FILLER_33_215 ();
 sg13g2_fill_1 FILLER_33_236 ();
 sg13g2_fill_2 FILLER_33_257 ();
 sg13g2_decap_8 FILLER_33_288 ();
 sg13g2_decap_8 FILLER_33_295 ();
 sg13g2_decap_4 FILLER_33_302 ();
 sg13g2_fill_2 FILLER_33_306 ();
 sg13g2_fill_2 FILLER_33_316 ();
 sg13g2_decap_8 FILLER_33_349 ();
 sg13g2_fill_2 FILLER_33_356 ();
 sg13g2_fill_2 FILLER_33_363 ();
 sg13g2_fill_1 FILLER_33_396 ();
 sg13g2_fill_1 FILLER_33_401 ();
 sg13g2_fill_2 FILLER_33_412 ();
 sg13g2_decap_4 FILLER_33_438 ();
 sg13g2_fill_1 FILLER_33_442 ();
 sg13g2_decap_4 FILLER_33_452 ();
 sg13g2_fill_1 FILLER_33_456 ();
 sg13g2_fill_2 FILLER_33_467 ();
 sg13g2_fill_1 FILLER_33_469 ();
 sg13g2_decap_8 FILLER_33_496 ();
 sg13g2_decap_8 FILLER_33_503 ();
 sg13g2_decap_8 FILLER_33_510 ();
 sg13g2_decap_8 FILLER_33_517 ();
 sg13g2_decap_8 FILLER_33_524 ();
 sg13g2_decap_8 FILLER_33_531 ();
 sg13g2_decap_8 FILLER_33_538 ();
 sg13g2_decap_8 FILLER_33_545 ();
 sg13g2_decap_8 FILLER_33_552 ();
 sg13g2_decap_8 FILLER_33_559 ();
 sg13g2_decap_8 FILLER_33_566 ();
 sg13g2_decap_8 FILLER_33_573 ();
 sg13g2_decap_8 FILLER_33_580 ();
 sg13g2_decap_8 FILLER_33_587 ();
 sg13g2_decap_8 FILLER_33_594 ();
 sg13g2_decap_8 FILLER_33_601 ();
 sg13g2_decap_8 FILLER_33_608 ();
 sg13g2_decap_8 FILLER_33_615 ();
 sg13g2_decap_8 FILLER_33_622 ();
 sg13g2_decap_8 FILLER_33_629 ();
 sg13g2_decap_8 FILLER_33_636 ();
 sg13g2_decap_8 FILLER_33_643 ();
 sg13g2_decap_8 FILLER_33_650 ();
 sg13g2_decap_8 FILLER_33_657 ();
 sg13g2_decap_8 FILLER_33_664 ();
 sg13g2_decap_8 FILLER_33_671 ();
 sg13g2_decap_8 FILLER_33_678 ();
 sg13g2_decap_8 FILLER_33_685 ();
 sg13g2_decap_8 FILLER_33_692 ();
 sg13g2_decap_8 FILLER_33_699 ();
 sg13g2_decap_8 FILLER_33_706 ();
 sg13g2_decap_8 FILLER_33_713 ();
 sg13g2_decap_8 FILLER_33_720 ();
 sg13g2_decap_8 FILLER_33_727 ();
 sg13g2_decap_8 FILLER_33_734 ();
 sg13g2_decap_8 FILLER_33_741 ();
 sg13g2_decap_8 FILLER_33_748 ();
 sg13g2_decap_8 FILLER_33_755 ();
 sg13g2_decap_8 FILLER_33_762 ();
 sg13g2_decap_8 FILLER_33_769 ();
 sg13g2_decap_8 FILLER_33_776 ();
 sg13g2_decap_8 FILLER_33_783 ();
 sg13g2_decap_8 FILLER_33_790 ();
 sg13g2_decap_8 FILLER_33_797 ();
 sg13g2_decap_8 FILLER_33_804 ();
 sg13g2_decap_8 FILLER_33_811 ();
 sg13g2_decap_8 FILLER_33_818 ();
 sg13g2_decap_8 FILLER_33_825 ();
 sg13g2_decap_8 FILLER_33_832 ();
 sg13g2_decap_8 FILLER_33_839 ();
 sg13g2_decap_8 FILLER_33_846 ();
 sg13g2_decap_8 FILLER_33_853 ();
 sg13g2_fill_2 FILLER_33_860 ();
 sg13g2_decap_4 FILLER_34_44 ();
 sg13g2_fill_2 FILLER_34_84 ();
 sg13g2_fill_1 FILLER_34_86 ();
 sg13g2_fill_1 FILLER_34_97 ();
 sg13g2_fill_2 FILLER_34_123 ();
 sg13g2_decap_4 FILLER_34_133 ();
 sg13g2_fill_2 FILLER_34_191 ();
 sg13g2_fill_2 FILLER_34_245 ();
 sg13g2_fill_1 FILLER_34_256 ();
 sg13g2_fill_1 FILLER_34_292 ();
 sg13g2_fill_1 FILLER_34_333 ();
 sg13g2_fill_2 FILLER_34_375 ();
 sg13g2_decap_4 FILLER_34_393 ();
 sg13g2_fill_1 FILLER_34_397 ();
 sg13g2_fill_1 FILLER_34_490 ();
 sg13g2_decap_8 FILLER_34_503 ();
 sg13g2_decap_8 FILLER_34_510 ();
 sg13g2_decap_8 FILLER_34_517 ();
 sg13g2_decap_8 FILLER_34_524 ();
 sg13g2_decap_8 FILLER_34_531 ();
 sg13g2_decap_8 FILLER_34_538 ();
 sg13g2_decap_8 FILLER_34_545 ();
 sg13g2_decap_8 FILLER_34_552 ();
 sg13g2_decap_8 FILLER_34_559 ();
 sg13g2_decap_8 FILLER_34_566 ();
 sg13g2_decap_8 FILLER_34_573 ();
 sg13g2_decap_8 FILLER_34_580 ();
 sg13g2_decap_8 FILLER_34_587 ();
 sg13g2_decap_8 FILLER_34_594 ();
 sg13g2_decap_8 FILLER_34_601 ();
 sg13g2_decap_8 FILLER_34_608 ();
 sg13g2_decap_8 FILLER_34_615 ();
 sg13g2_decap_8 FILLER_34_622 ();
 sg13g2_decap_8 FILLER_34_629 ();
 sg13g2_decap_8 FILLER_34_636 ();
 sg13g2_decap_8 FILLER_34_643 ();
 sg13g2_decap_8 FILLER_34_650 ();
 sg13g2_decap_8 FILLER_34_657 ();
 sg13g2_decap_8 FILLER_34_664 ();
 sg13g2_decap_8 FILLER_34_671 ();
 sg13g2_decap_8 FILLER_34_678 ();
 sg13g2_decap_8 FILLER_34_685 ();
 sg13g2_decap_8 FILLER_34_692 ();
 sg13g2_decap_8 FILLER_34_699 ();
 sg13g2_decap_8 FILLER_34_706 ();
 sg13g2_decap_8 FILLER_34_713 ();
 sg13g2_decap_8 FILLER_34_720 ();
 sg13g2_decap_8 FILLER_34_727 ();
 sg13g2_decap_8 FILLER_34_734 ();
 sg13g2_decap_8 FILLER_34_741 ();
 sg13g2_decap_8 FILLER_34_748 ();
 sg13g2_decap_8 FILLER_34_755 ();
 sg13g2_decap_8 FILLER_34_762 ();
 sg13g2_decap_8 FILLER_34_769 ();
 sg13g2_decap_8 FILLER_34_776 ();
 sg13g2_decap_8 FILLER_34_783 ();
 sg13g2_decap_8 FILLER_34_790 ();
 sg13g2_decap_8 FILLER_34_797 ();
 sg13g2_decap_8 FILLER_34_804 ();
 sg13g2_decap_8 FILLER_34_811 ();
 sg13g2_decap_8 FILLER_34_818 ();
 sg13g2_decap_8 FILLER_34_825 ();
 sg13g2_decap_8 FILLER_34_832 ();
 sg13g2_decap_8 FILLER_34_839 ();
 sg13g2_decap_8 FILLER_34_846 ();
 sg13g2_decap_8 FILLER_34_853 ();
 sg13g2_fill_2 FILLER_34_860 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_fill_2 FILLER_35_21 ();
 sg13g2_fill_1 FILLER_35_23 ();
 sg13g2_fill_1 FILLER_35_32 ();
 sg13g2_decap_8 FILLER_35_45 ();
 sg13g2_decap_4 FILLER_35_52 ();
 sg13g2_fill_1 FILLER_35_56 ();
 sg13g2_fill_2 FILLER_35_74 ();
 sg13g2_fill_1 FILLER_35_76 ();
 sg13g2_fill_2 FILLER_35_93 ();
 sg13g2_fill_2 FILLER_35_169 ();
 sg13g2_fill_1 FILLER_35_217 ();
 sg13g2_fill_1 FILLER_35_230 ();
 sg13g2_fill_1 FILLER_35_252 ();
 sg13g2_fill_2 FILLER_35_266 ();
 sg13g2_fill_2 FILLER_35_286 ();
 sg13g2_fill_1 FILLER_35_288 ();
 sg13g2_fill_2 FILLER_35_302 ();
 sg13g2_fill_2 FILLER_35_308 ();
 sg13g2_fill_1 FILLER_35_310 ();
 sg13g2_fill_2 FILLER_35_321 ();
 sg13g2_fill_1 FILLER_35_323 ();
 sg13g2_decap_4 FILLER_35_332 ();
 sg13g2_fill_1 FILLER_35_336 ();
 sg13g2_fill_2 FILLER_35_342 ();
 sg13g2_fill_2 FILLER_35_358 ();
 sg13g2_fill_1 FILLER_35_360 ();
 sg13g2_fill_2 FILLER_35_380 ();
 sg13g2_decap_4 FILLER_35_397 ();
 sg13g2_fill_2 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_406 ();
 sg13g2_fill_2 FILLER_35_417 ();
 sg13g2_fill_1 FILLER_35_419 ();
 sg13g2_fill_2 FILLER_35_460 ();
 sg13g2_fill_2 FILLER_35_472 ();
 sg13g2_fill_1 FILLER_35_474 ();
 sg13g2_decap_8 FILLER_35_505 ();
 sg13g2_decap_8 FILLER_35_512 ();
 sg13g2_decap_8 FILLER_35_519 ();
 sg13g2_decap_8 FILLER_35_526 ();
 sg13g2_decap_8 FILLER_35_533 ();
 sg13g2_decap_8 FILLER_35_540 ();
 sg13g2_decap_8 FILLER_35_547 ();
 sg13g2_decap_8 FILLER_35_554 ();
 sg13g2_decap_8 FILLER_35_561 ();
 sg13g2_decap_8 FILLER_35_568 ();
 sg13g2_decap_8 FILLER_35_575 ();
 sg13g2_decap_8 FILLER_35_582 ();
 sg13g2_decap_8 FILLER_35_589 ();
 sg13g2_decap_8 FILLER_35_596 ();
 sg13g2_decap_8 FILLER_35_603 ();
 sg13g2_decap_8 FILLER_35_610 ();
 sg13g2_decap_8 FILLER_35_617 ();
 sg13g2_decap_8 FILLER_35_624 ();
 sg13g2_decap_8 FILLER_35_631 ();
 sg13g2_decap_8 FILLER_35_638 ();
 sg13g2_decap_8 FILLER_35_645 ();
 sg13g2_decap_8 FILLER_35_652 ();
 sg13g2_decap_8 FILLER_35_659 ();
 sg13g2_decap_8 FILLER_35_666 ();
 sg13g2_decap_8 FILLER_35_673 ();
 sg13g2_decap_8 FILLER_35_680 ();
 sg13g2_decap_8 FILLER_35_687 ();
 sg13g2_decap_8 FILLER_35_694 ();
 sg13g2_decap_8 FILLER_35_701 ();
 sg13g2_decap_8 FILLER_35_708 ();
 sg13g2_decap_8 FILLER_35_715 ();
 sg13g2_decap_8 FILLER_35_722 ();
 sg13g2_decap_8 FILLER_35_729 ();
 sg13g2_decap_8 FILLER_35_736 ();
 sg13g2_decap_8 FILLER_35_743 ();
 sg13g2_decap_8 FILLER_35_750 ();
 sg13g2_decap_8 FILLER_35_757 ();
 sg13g2_decap_8 FILLER_35_764 ();
 sg13g2_decap_8 FILLER_35_771 ();
 sg13g2_decap_8 FILLER_35_778 ();
 sg13g2_decap_8 FILLER_35_785 ();
 sg13g2_decap_8 FILLER_35_792 ();
 sg13g2_decap_8 FILLER_35_799 ();
 sg13g2_decap_8 FILLER_35_806 ();
 sg13g2_decap_8 FILLER_35_813 ();
 sg13g2_decap_8 FILLER_35_820 ();
 sg13g2_decap_8 FILLER_35_827 ();
 sg13g2_decap_8 FILLER_35_834 ();
 sg13g2_decap_8 FILLER_35_841 ();
 sg13g2_decap_8 FILLER_35_848 ();
 sg13g2_decap_8 FILLER_35_855 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_fill_2 FILLER_36_21 ();
 sg13g2_fill_1 FILLER_36_23 ();
 sg13g2_fill_1 FILLER_36_32 ();
 sg13g2_fill_2 FILLER_36_38 ();
 sg13g2_fill_1 FILLER_36_40 ();
 sg13g2_fill_2 FILLER_36_85 ();
 sg13g2_fill_2 FILLER_36_99 ();
 sg13g2_fill_1 FILLER_36_101 ();
 sg13g2_fill_1 FILLER_36_111 ();
 sg13g2_decap_4 FILLER_36_182 ();
 sg13g2_fill_2 FILLER_36_259 ();
 sg13g2_decap_8 FILLER_36_283 ();
 sg13g2_fill_2 FILLER_36_290 ();
 sg13g2_fill_1 FILLER_36_292 ();
 sg13g2_fill_1 FILLER_36_298 ();
 sg13g2_fill_1 FILLER_36_344 ();
 sg13g2_fill_2 FILLER_36_364 ();
 sg13g2_fill_2 FILLER_36_432 ();
 sg13g2_fill_2 FILLER_36_452 ();
 sg13g2_fill_1 FILLER_36_454 ();
 sg13g2_fill_2 FILLER_36_460 ();
 sg13g2_fill_1 FILLER_36_462 ();
 sg13g2_fill_1 FILLER_36_487 ();
 sg13g2_decap_8 FILLER_36_505 ();
 sg13g2_decap_8 FILLER_36_512 ();
 sg13g2_decap_8 FILLER_36_519 ();
 sg13g2_decap_8 FILLER_36_526 ();
 sg13g2_decap_8 FILLER_36_533 ();
 sg13g2_decap_8 FILLER_36_540 ();
 sg13g2_decap_8 FILLER_36_547 ();
 sg13g2_decap_8 FILLER_36_554 ();
 sg13g2_decap_8 FILLER_36_561 ();
 sg13g2_decap_8 FILLER_36_568 ();
 sg13g2_decap_8 FILLER_36_575 ();
 sg13g2_decap_8 FILLER_36_582 ();
 sg13g2_decap_8 FILLER_36_589 ();
 sg13g2_decap_8 FILLER_36_596 ();
 sg13g2_decap_8 FILLER_36_603 ();
 sg13g2_decap_8 FILLER_36_610 ();
 sg13g2_decap_8 FILLER_36_617 ();
 sg13g2_decap_8 FILLER_36_624 ();
 sg13g2_decap_8 FILLER_36_631 ();
 sg13g2_decap_8 FILLER_36_638 ();
 sg13g2_decap_8 FILLER_36_645 ();
 sg13g2_decap_8 FILLER_36_652 ();
 sg13g2_decap_8 FILLER_36_659 ();
 sg13g2_decap_8 FILLER_36_666 ();
 sg13g2_decap_8 FILLER_36_673 ();
 sg13g2_decap_8 FILLER_36_680 ();
 sg13g2_decap_8 FILLER_36_687 ();
 sg13g2_decap_8 FILLER_36_694 ();
 sg13g2_decap_8 FILLER_36_701 ();
 sg13g2_decap_8 FILLER_36_708 ();
 sg13g2_decap_8 FILLER_36_715 ();
 sg13g2_decap_8 FILLER_36_722 ();
 sg13g2_decap_8 FILLER_36_729 ();
 sg13g2_decap_8 FILLER_36_736 ();
 sg13g2_decap_8 FILLER_36_743 ();
 sg13g2_decap_8 FILLER_36_750 ();
 sg13g2_decap_8 FILLER_36_757 ();
 sg13g2_decap_8 FILLER_36_764 ();
 sg13g2_decap_8 FILLER_36_771 ();
 sg13g2_decap_8 FILLER_36_778 ();
 sg13g2_decap_8 FILLER_36_785 ();
 sg13g2_decap_8 FILLER_36_792 ();
 sg13g2_decap_8 FILLER_36_799 ();
 sg13g2_decap_8 FILLER_36_806 ();
 sg13g2_decap_8 FILLER_36_813 ();
 sg13g2_decap_8 FILLER_36_820 ();
 sg13g2_decap_8 FILLER_36_827 ();
 sg13g2_decap_8 FILLER_36_834 ();
 sg13g2_decap_8 FILLER_36_841 ();
 sg13g2_decap_8 FILLER_36_848 ();
 sg13g2_decap_8 FILLER_36_855 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_4 FILLER_37_14 ();
 sg13g2_fill_1 FILLER_37_31 ();
 sg13g2_fill_2 FILLER_37_40 ();
 sg13g2_fill_1 FILLER_37_42 ();
 sg13g2_decap_4 FILLER_37_56 ();
 sg13g2_fill_2 FILLER_37_60 ();
 sg13g2_fill_2 FILLER_37_106 ();
 sg13g2_fill_1 FILLER_37_108 ();
 sg13g2_fill_2 FILLER_37_114 ();
 sg13g2_fill_1 FILLER_37_116 ();
 sg13g2_fill_2 FILLER_37_126 ();
 sg13g2_fill_1 FILLER_37_132 ();
 sg13g2_decap_4 FILLER_37_145 ();
 sg13g2_fill_1 FILLER_37_149 ();
 sg13g2_decap_8 FILLER_37_158 ();
 sg13g2_fill_1 FILLER_37_165 ();
 sg13g2_fill_2 FILLER_37_171 ();
 sg13g2_decap_8 FILLER_37_209 ();
 sg13g2_fill_1 FILLER_37_216 ();
 sg13g2_decap_4 FILLER_37_236 ();
 sg13g2_fill_1 FILLER_37_240 ();
 sg13g2_decap_8 FILLER_37_249 ();
 sg13g2_decap_4 FILLER_37_256 ();
 sg13g2_fill_2 FILLER_37_260 ();
 sg13g2_fill_2 FILLER_37_308 ();
 sg13g2_fill_1 FILLER_37_310 ();
 sg13g2_fill_1 FILLER_37_324 ();
 sg13g2_decap_4 FILLER_37_334 ();
 sg13g2_fill_2 FILLER_37_338 ();
 sg13g2_fill_2 FILLER_37_361 ();
 sg13g2_fill_2 FILLER_37_367 ();
 sg13g2_fill_1 FILLER_37_369 ();
 sg13g2_decap_8 FILLER_37_379 ();
 sg13g2_fill_2 FILLER_37_386 ();
 sg13g2_decap_4 FILLER_37_396 ();
 sg13g2_fill_2 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_413 ();
 sg13g2_fill_1 FILLER_37_415 ();
 sg13g2_decap_8 FILLER_37_421 ();
 sg13g2_decap_8 FILLER_37_510 ();
 sg13g2_decap_8 FILLER_37_517 ();
 sg13g2_decap_8 FILLER_37_524 ();
 sg13g2_decap_8 FILLER_37_531 ();
 sg13g2_decap_8 FILLER_37_538 ();
 sg13g2_decap_8 FILLER_37_545 ();
 sg13g2_decap_8 FILLER_37_552 ();
 sg13g2_decap_8 FILLER_37_559 ();
 sg13g2_decap_8 FILLER_37_566 ();
 sg13g2_decap_8 FILLER_37_573 ();
 sg13g2_decap_8 FILLER_37_580 ();
 sg13g2_decap_8 FILLER_37_587 ();
 sg13g2_decap_8 FILLER_37_594 ();
 sg13g2_decap_8 FILLER_37_601 ();
 sg13g2_decap_8 FILLER_37_608 ();
 sg13g2_decap_8 FILLER_37_615 ();
 sg13g2_decap_8 FILLER_37_622 ();
 sg13g2_decap_8 FILLER_37_629 ();
 sg13g2_decap_8 FILLER_37_636 ();
 sg13g2_decap_8 FILLER_37_643 ();
 sg13g2_decap_8 FILLER_37_650 ();
 sg13g2_decap_8 FILLER_37_657 ();
 sg13g2_decap_8 FILLER_37_664 ();
 sg13g2_decap_8 FILLER_37_671 ();
 sg13g2_decap_8 FILLER_37_678 ();
 sg13g2_decap_8 FILLER_37_685 ();
 sg13g2_decap_8 FILLER_37_692 ();
 sg13g2_decap_8 FILLER_37_699 ();
 sg13g2_decap_8 FILLER_37_706 ();
 sg13g2_decap_8 FILLER_37_713 ();
 sg13g2_decap_8 FILLER_37_720 ();
 sg13g2_decap_8 FILLER_37_727 ();
 sg13g2_decap_8 FILLER_37_734 ();
 sg13g2_decap_8 FILLER_37_741 ();
 sg13g2_decap_8 FILLER_37_748 ();
 sg13g2_decap_8 FILLER_37_755 ();
 sg13g2_decap_8 FILLER_37_762 ();
 sg13g2_decap_8 FILLER_37_769 ();
 sg13g2_decap_8 FILLER_37_776 ();
 sg13g2_decap_8 FILLER_37_783 ();
 sg13g2_decap_8 FILLER_37_790 ();
 sg13g2_decap_8 FILLER_37_797 ();
 sg13g2_decap_8 FILLER_37_804 ();
 sg13g2_decap_8 FILLER_37_811 ();
 sg13g2_decap_8 FILLER_37_818 ();
 sg13g2_decap_8 FILLER_37_825 ();
 sg13g2_decap_8 FILLER_37_832 ();
 sg13g2_decap_8 FILLER_37_839 ();
 sg13g2_decap_8 FILLER_37_846 ();
 sg13g2_decap_8 FILLER_37_853 ();
 sg13g2_fill_2 FILLER_37_860 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_58 ();
 sg13g2_decap_4 FILLER_38_65 ();
 sg13g2_fill_1 FILLER_38_69 ();
 sg13g2_fill_2 FILLER_38_84 ();
 sg13g2_fill_1 FILLER_38_86 ();
 sg13g2_fill_2 FILLER_38_105 ();
 sg13g2_fill_1 FILLER_38_107 ();
 sg13g2_fill_1 FILLER_38_116 ();
 sg13g2_fill_1 FILLER_38_127 ();
 sg13g2_decap_8 FILLER_38_164 ();
 sg13g2_fill_2 FILLER_38_171 ();
 sg13g2_decap_4 FILLER_38_178 ();
 sg13g2_fill_2 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_188 ();
 sg13g2_fill_2 FILLER_38_222 ();
 sg13g2_fill_1 FILLER_38_224 ();
 sg13g2_fill_2 FILLER_38_230 ();
 sg13g2_fill_1 FILLER_38_232 ();
 sg13g2_fill_2 FILLER_38_249 ();
 sg13g2_fill_1 FILLER_38_251 ();
 sg13g2_decap_8 FILLER_38_257 ();
 sg13g2_fill_1 FILLER_38_264 ();
 sg13g2_fill_1 FILLER_38_274 ();
 sg13g2_fill_2 FILLER_38_294 ();
 sg13g2_decap_4 FILLER_38_309 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_decap_4 FILLER_38_356 ();
 sg13g2_decap_8 FILLER_38_364 ();
 sg13g2_fill_1 FILLER_38_371 ();
 sg13g2_fill_2 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_decap_4 FILLER_38_407 ();
 sg13g2_decap_4 FILLER_38_419 ();
 sg13g2_fill_2 FILLER_38_433 ();
 sg13g2_decap_8 FILLER_38_444 ();
 sg13g2_decap_4 FILLER_38_451 ();
 sg13g2_fill_2 FILLER_38_455 ();
 sg13g2_fill_2 FILLER_38_466 ();
 sg13g2_decap_8 FILLER_38_472 ();
 sg13g2_decap_8 FILLER_38_479 ();
 sg13g2_decap_8 FILLER_38_486 ();
 sg13g2_decap_8 FILLER_38_493 ();
 sg13g2_decap_8 FILLER_38_500 ();
 sg13g2_decap_8 FILLER_38_507 ();
 sg13g2_decap_8 FILLER_38_514 ();
 sg13g2_decap_8 FILLER_38_521 ();
 sg13g2_decap_8 FILLER_38_528 ();
 sg13g2_decap_8 FILLER_38_535 ();
 sg13g2_decap_8 FILLER_38_542 ();
 sg13g2_decap_8 FILLER_38_549 ();
 sg13g2_decap_8 FILLER_38_556 ();
 sg13g2_decap_8 FILLER_38_563 ();
 sg13g2_decap_8 FILLER_38_570 ();
 sg13g2_decap_8 FILLER_38_577 ();
 sg13g2_decap_8 FILLER_38_584 ();
 sg13g2_decap_8 FILLER_38_591 ();
 sg13g2_decap_8 FILLER_38_598 ();
 sg13g2_decap_8 FILLER_38_605 ();
 sg13g2_decap_8 FILLER_38_612 ();
 sg13g2_decap_8 FILLER_38_619 ();
 sg13g2_decap_8 FILLER_38_626 ();
 sg13g2_decap_8 FILLER_38_633 ();
 sg13g2_decap_8 FILLER_38_640 ();
 sg13g2_decap_8 FILLER_38_647 ();
 sg13g2_decap_8 FILLER_38_654 ();
 sg13g2_decap_8 FILLER_38_661 ();
 sg13g2_decap_8 FILLER_38_668 ();
 sg13g2_decap_8 FILLER_38_675 ();
 sg13g2_decap_8 FILLER_38_682 ();
 sg13g2_decap_8 FILLER_38_689 ();
 sg13g2_decap_8 FILLER_38_696 ();
 sg13g2_decap_8 FILLER_38_703 ();
 sg13g2_decap_8 FILLER_38_710 ();
 sg13g2_decap_8 FILLER_38_717 ();
 sg13g2_decap_8 FILLER_38_724 ();
 sg13g2_decap_8 FILLER_38_731 ();
 sg13g2_decap_8 FILLER_38_738 ();
 sg13g2_decap_8 FILLER_38_745 ();
 sg13g2_decap_8 FILLER_38_752 ();
 sg13g2_decap_8 FILLER_38_759 ();
 sg13g2_decap_8 FILLER_38_766 ();
 sg13g2_decap_8 FILLER_38_773 ();
 sg13g2_decap_8 FILLER_38_780 ();
 sg13g2_decap_8 FILLER_38_787 ();
 sg13g2_decap_8 FILLER_38_794 ();
 sg13g2_decap_8 FILLER_38_801 ();
 sg13g2_decap_8 FILLER_38_808 ();
 sg13g2_decap_8 FILLER_38_815 ();
 sg13g2_decap_8 FILLER_38_822 ();
 sg13g2_decap_8 FILLER_38_829 ();
 sg13g2_decap_8 FILLER_38_836 ();
 sg13g2_decap_8 FILLER_38_843 ();
 sg13g2_decap_8 FILLER_38_850 ();
 sg13g2_decap_4 FILLER_38_857 ();
 sg13g2_fill_1 FILLER_38_861 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_4 FILLER_39_7 ();
 sg13g2_fill_2 FILLER_39_11 ();
 sg13g2_decap_8 FILLER_39_17 ();
 sg13g2_decap_4 FILLER_39_24 ();
 sg13g2_fill_2 FILLER_39_28 ();
 sg13g2_fill_2 FILLER_39_71 ();
 sg13g2_fill_1 FILLER_39_73 ();
 sg13g2_fill_1 FILLER_39_100 ();
 sg13g2_fill_1 FILLER_39_122 ();
 sg13g2_decap_4 FILLER_39_155 ();
 sg13g2_fill_2 FILLER_39_162 ();
 sg13g2_fill_2 FILLER_39_197 ();
 sg13g2_fill_2 FILLER_39_265 ();
 sg13g2_fill_1 FILLER_39_267 ();
 sg13g2_fill_2 FILLER_39_292 ();
 sg13g2_fill_1 FILLER_39_294 ();
 sg13g2_decap_8 FILLER_39_331 ();
 sg13g2_fill_2 FILLER_39_338 ();
 sg13g2_fill_1 FILLER_39_340 ();
 sg13g2_fill_1 FILLER_39_355 ();
 sg13g2_fill_1 FILLER_39_383 ();
 sg13g2_decap_4 FILLER_39_433 ();
 sg13g2_fill_1 FILLER_39_443 ();
 sg13g2_decap_8 FILLER_39_479 ();
 sg13g2_decap_8 FILLER_39_486 ();
 sg13g2_decap_8 FILLER_39_493 ();
 sg13g2_decap_8 FILLER_39_500 ();
 sg13g2_decap_8 FILLER_39_507 ();
 sg13g2_decap_8 FILLER_39_514 ();
 sg13g2_decap_8 FILLER_39_521 ();
 sg13g2_decap_8 FILLER_39_528 ();
 sg13g2_decap_8 FILLER_39_535 ();
 sg13g2_decap_8 FILLER_39_542 ();
 sg13g2_decap_8 FILLER_39_549 ();
 sg13g2_decap_8 FILLER_39_556 ();
 sg13g2_decap_8 FILLER_39_563 ();
 sg13g2_decap_8 FILLER_39_570 ();
 sg13g2_decap_8 FILLER_39_577 ();
 sg13g2_decap_8 FILLER_39_584 ();
 sg13g2_decap_8 FILLER_39_591 ();
 sg13g2_decap_8 FILLER_39_598 ();
 sg13g2_decap_8 FILLER_39_605 ();
 sg13g2_decap_8 FILLER_39_612 ();
 sg13g2_decap_8 FILLER_39_619 ();
 sg13g2_decap_8 FILLER_39_626 ();
 sg13g2_decap_8 FILLER_39_633 ();
 sg13g2_decap_8 FILLER_39_640 ();
 sg13g2_decap_8 FILLER_39_647 ();
 sg13g2_decap_8 FILLER_39_654 ();
 sg13g2_decap_8 FILLER_39_661 ();
 sg13g2_decap_8 FILLER_39_668 ();
 sg13g2_decap_8 FILLER_39_675 ();
 sg13g2_decap_8 FILLER_39_682 ();
 sg13g2_decap_8 FILLER_39_689 ();
 sg13g2_decap_8 FILLER_39_696 ();
 sg13g2_decap_8 FILLER_39_703 ();
 sg13g2_decap_8 FILLER_39_710 ();
 sg13g2_decap_8 FILLER_39_717 ();
 sg13g2_decap_8 FILLER_39_724 ();
 sg13g2_decap_8 FILLER_39_731 ();
 sg13g2_decap_8 FILLER_39_738 ();
 sg13g2_decap_8 FILLER_39_745 ();
 sg13g2_decap_8 FILLER_39_752 ();
 sg13g2_decap_8 FILLER_39_759 ();
 sg13g2_decap_8 FILLER_39_766 ();
 sg13g2_decap_8 FILLER_39_773 ();
 sg13g2_decap_8 FILLER_39_780 ();
 sg13g2_decap_8 FILLER_39_787 ();
 sg13g2_decap_8 FILLER_39_794 ();
 sg13g2_decap_8 FILLER_39_801 ();
 sg13g2_decap_8 FILLER_39_808 ();
 sg13g2_decap_8 FILLER_39_815 ();
 sg13g2_decap_8 FILLER_39_822 ();
 sg13g2_decap_8 FILLER_39_829 ();
 sg13g2_decap_8 FILLER_39_836 ();
 sg13g2_decap_8 FILLER_39_843 ();
 sg13g2_decap_8 FILLER_39_850 ();
 sg13g2_decap_4 FILLER_39_857 ();
 sg13g2_fill_1 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_4 FILLER_40_14 ();
 sg13g2_fill_1 FILLER_40_18 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_4 FILLER_40_35 ();
 sg13g2_decap_4 FILLER_40_61 ();
 sg13g2_fill_2 FILLER_40_65 ();
 sg13g2_decap_4 FILLER_40_77 ();
 sg13g2_fill_2 FILLER_40_81 ();
 sg13g2_decap_4 FILLER_40_97 ();
 sg13g2_decap_8 FILLER_40_123 ();
 sg13g2_decap_8 FILLER_40_157 ();
 sg13g2_decap_4 FILLER_40_164 ();
 sg13g2_decap_4 FILLER_40_177 ();
 sg13g2_fill_2 FILLER_40_185 ();
 sg13g2_fill_2 FILLER_40_217 ();
 sg13g2_fill_1 FILLER_40_225 ();
 sg13g2_fill_2 FILLER_40_258 ();
 sg13g2_fill_1 FILLER_40_281 ();
 sg13g2_decap_8 FILLER_40_290 ();
 sg13g2_decap_8 FILLER_40_297 ();
 sg13g2_fill_2 FILLER_40_304 ();
 sg13g2_decap_4 FILLER_40_310 ();
 sg13g2_fill_2 FILLER_40_314 ();
 sg13g2_decap_4 FILLER_40_357 ();
 sg13g2_fill_2 FILLER_40_371 ();
 sg13g2_fill_2 FILLER_40_383 ();
 sg13g2_fill_2 FILLER_40_403 ();
 sg13g2_decap_4 FILLER_40_416 ();
 sg13g2_fill_2 FILLER_40_420 ();
 sg13g2_decap_4 FILLER_40_431 ();
 sg13g2_fill_2 FILLER_40_435 ();
 sg13g2_decap_4 FILLER_40_441 ();
 sg13g2_fill_1 FILLER_40_463 ();
 sg13g2_decap_8 FILLER_40_468 ();
 sg13g2_decap_8 FILLER_40_475 ();
 sg13g2_decap_8 FILLER_40_482 ();
 sg13g2_decap_8 FILLER_40_489 ();
 sg13g2_decap_8 FILLER_40_496 ();
 sg13g2_decap_8 FILLER_40_503 ();
 sg13g2_decap_8 FILLER_40_510 ();
 sg13g2_decap_8 FILLER_40_517 ();
 sg13g2_decap_8 FILLER_40_524 ();
 sg13g2_decap_8 FILLER_40_531 ();
 sg13g2_decap_8 FILLER_40_538 ();
 sg13g2_decap_8 FILLER_40_545 ();
 sg13g2_decap_8 FILLER_40_552 ();
 sg13g2_decap_8 FILLER_40_559 ();
 sg13g2_decap_8 FILLER_40_566 ();
 sg13g2_decap_8 FILLER_40_573 ();
 sg13g2_decap_8 FILLER_40_580 ();
 sg13g2_decap_8 FILLER_40_587 ();
 sg13g2_decap_8 FILLER_40_594 ();
 sg13g2_decap_8 FILLER_40_601 ();
 sg13g2_decap_8 FILLER_40_608 ();
 sg13g2_decap_8 FILLER_40_615 ();
 sg13g2_decap_8 FILLER_40_622 ();
 sg13g2_decap_8 FILLER_40_629 ();
 sg13g2_decap_8 FILLER_40_636 ();
 sg13g2_decap_8 FILLER_40_643 ();
 sg13g2_decap_8 FILLER_40_650 ();
 sg13g2_decap_8 FILLER_40_657 ();
 sg13g2_decap_8 FILLER_40_664 ();
 sg13g2_decap_8 FILLER_40_671 ();
 sg13g2_decap_8 FILLER_40_678 ();
 sg13g2_decap_8 FILLER_40_685 ();
 sg13g2_decap_8 FILLER_40_692 ();
 sg13g2_decap_8 FILLER_40_699 ();
 sg13g2_decap_8 FILLER_40_706 ();
 sg13g2_decap_8 FILLER_40_713 ();
 sg13g2_decap_8 FILLER_40_720 ();
 sg13g2_decap_8 FILLER_40_727 ();
 sg13g2_decap_8 FILLER_40_734 ();
 sg13g2_decap_8 FILLER_40_741 ();
 sg13g2_decap_8 FILLER_40_748 ();
 sg13g2_decap_8 FILLER_40_755 ();
 sg13g2_decap_8 FILLER_40_762 ();
 sg13g2_decap_8 FILLER_40_769 ();
 sg13g2_decap_8 FILLER_40_776 ();
 sg13g2_decap_8 FILLER_40_783 ();
 sg13g2_decap_8 FILLER_40_790 ();
 sg13g2_decap_8 FILLER_40_797 ();
 sg13g2_decap_8 FILLER_40_804 ();
 sg13g2_decap_8 FILLER_40_811 ();
 sg13g2_decap_8 FILLER_40_818 ();
 sg13g2_decap_8 FILLER_40_825 ();
 sg13g2_decap_8 FILLER_40_832 ();
 sg13g2_decap_8 FILLER_40_839 ();
 sg13g2_decap_8 FILLER_40_846 ();
 sg13g2_decap_8 FILLER_40_853 ();
 sg13g2_fill_2 FILLER_40_860 ();
 sg13g2_decap_4 FILLER_41_34 ();
 sg13g2_fill_2 FILLER_41_43 ();
 sg13g2_fill_1 FILLER_41_45 ();
 sg13g2_decap_4 FILLER_41_59 ();
 sg13g2_decap_8 FILLER_41_115 ();
 sg13g2_fill_2 FILLER_41_122 ();
 sg13g2_fill_1 FILLER_41_124 ();
 sg13g2_fill_2 FILLER_41_183 ();
 sg13g2_fill_2 FILLER_41_215 ();
 sg13g2_decap_8 FILLER_41_243 ();
 sg13g2_fill_1 FILLER_41_250 ();
 sg13g2_fill_1 FILLER_41_287 ();
 sg13g2_fill_2 FILLER_41_300 ();
 sg13g2_decap_4 FILLER_41_312 ();
 sg13g2_fill_2 FILLER_41_321 ();
 sg13g2_fill_2 FILLER_41_337 ();
 sg13g2_decap_8 FILLER_41_348 ();
 sg13g2_fill_2 FILLER_41_355 ();
 sg13g2_fill_1 FILLER_41_357 ();
 sg13g2_fill_2 FILLER_41_380 ();
 sg13g2_decap_4 FILLER_41_403 ();
 sg13g2_fill_2 FILLER_41_407 ();
 sg13g2_fill_1 FILLER_41_418 ();
 sg13g2_decap_4 FILLER_41_434 ();
 sg13g2_fill_1 FILLER_41_443 ();
 sg13g2_decap_8 FILLER_41_459 ();
 sg13g2_decap_4 FILLER_41_466 ();
 sg13g2_fill_1 FILLER_41_470 ();
 sg13g2_decap_8 FILLER_41_475 ();
 sg13g2_decap_8 FILLER_41_482 ();
 sg13g2_decap_8 FILLER_41_489 ();
 sg13g2_decap_8 FILLER_41_496 ();
 sg13g2_decap_8 FILLER_41_503 ();
 sg13g2_decap_8 FILLER_41_510 ();
 sg13g2_decap_8 FILLER_41_517 ();
 sg13g2_decap_8 FILLER_41_524 ();
 sg13g2_decap_8 FILLER_41_531 ();
 sg13g2_decap_8 FILLER_41_538 ();
 sg13g2_decap_8 FILLER_41_545 ();
 sg13g2_decap_8 FILLER_41_552 ();
 sg13g2_decap_8 FILLER_41_559 ();
 sg13g2_decap_8 FILLER_41_566 ();
 sg13g2_decap_8 FILLER_41_573 ();
 sg13g2_decap_8 FILLER_41_580 ();
 sg13g2_decap_8 FILLER_41_587 ();
 sg13g2_decap_8 FILLER_41_594 ();
 sg13g2_decap_8 FILLER_41_601 ();
 sg13g2_decap_8 FILLER_41_608 ();
 sg13g2_decap_8 FILLER_41_615 ();
 sg13g2_decap_8 FILLER_41_622 ();
 sg13g2_decap_8 FILLER_41_629 ();
 sg13g2_decap_8 FILLER_41_636 ();
 sg13g2_decap_8 FILLER_41_643 ();
 sg13g2_decap_8 FILLER_41_650 ();
 sg13g2_decap_8 FILLER_41_657 ();
 sg13g2_decap_8 FILLER_41_664 ();
 sg13g2_decap_8 FILLER_41_671 ();
 sg13g2_decap_8 FILLER_41_678 ();
 sg13g2_decap_8 FILLER_41_685 ();
 sg13g2_decap_8 FILLER_41_692 ();
 sg13g2_decap_8 FILLER_41_699 ();
 sg13g2_decap_8 FILLER_41_706 ();
 sg13g2_decap_8 FILLER_41_713 ();
 sg13g2_decap_8 FILLER_41_720 ();
 sg13g2_decap_8 FILLER_41_727 ();
 sg13g2_decap_8 FILLER_41_734 ();
 sg13g2_decap_8 FILLER_41_741 ();
 sg13g2_decap_8 FILLER_41_748 ();
 sg13g2_decap_8 FILLER_41_755 ();
 sg13g2_decap_8 FILLER_41_762 ();
 sg13g2_decap_8 FILLER_41_769 ();
 sg13g2_decap_8 FILLER_41_776 ();
 sg13g2_decap_8 FILLER_41_783 ();
 sg13g2_decap_8 FILLER_41_790 ();
 sg13g2_decap_8 FILLER_41_797 ();
 sg13g2_decap_8 FILLER_41_804 ();
 sg13g2_decap_8 FILLER_41_811 ();
 sg13g2_decap_8 FILLER_41_818 ();
 sg13g2_decap_8 FILLER_41_825 ();
 sg13g2_decap_8 FILLER_41_832 ();
 sg13g2_decap_8 FILLER_41_839 ();
 sg13g2_decap_8 FILLER_41_846 ();
 sg13g2_decap_8 FILLER_41_853 ();
 sg13g2_fill_2 FILLER_41_860 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_7 ();
 sg13g2_fill_1 FILLER_42_9 ();
 sg13g2_fill_2 FILLER_42_74 ();
 sg13g2_decap_8 FILLER_42_89 ();
 sg13g2_fill_1 FILLER_42_96 ();
 sg13g2_fill_2 FILLER_42_137 ();
 sg13g2_fill_1 FILLER_42_139 ();
 sg13g2_fill_1 FILLER_42_166 ();
 sg13g2_decap_4 FILLER_42_180 ();
 sg13g2_fill_2 FILLER_42_198 ();
 sg13g2_fill_2 FILLER_42_220 ();
 sg13g2_fill_2 FILLER_42_226 ();
 sg13g2_fill_2 FILLER_42_235 ();
 sg13g2_fill_1 FILLER_42_237 ();
 sg13g2_decap_4 FILLER_42_248 ();
 sg13g2_fill_1 FILLER_42_252 ();
 sg13g2_fill_2 FILLER_42_257 ();
 sg13g2_decap_4 FILLER_42_277 ();
 sg13g2_fill_2 FILLER_42_281 ();
 sg13g2_fill_2 FILLER_42_287 ();
 sg13g2_decap_4 FILLER_42_298 ();
 sg13g2_fill_2 FILLER_42_302 ();
 sg13g2_decap_8 FILLER_42_350 ();
 sg13g2_decap_8 FILLER_42_357 ();
 sg13g2_fill_1 FILLER_42_364 ();
 sg13g2_decap_8 FILLER_42_375 ();
 sg13g2_decap_8 FILLER_42_387 ();
 sg13g2_decap_4 FILLER_42_394 ();
 sg13g2_fill_1 FILLER_42_398 ();
 sg13g2_decap_4 FILLER_42_414 ();
 sg13g2_fill_2 FILLER_42_418 ();
 sg13g2_decap_4 FILLER_42_430 ();
 sg13g2_fill_1 FILLER_42_444 ();
 sg13g2_fill_1 FILLER_42_455 ();
 sg13g2_decap_8 FILLER_42_489 ();
 sg13g2_decap_4 FILLER_42_496 ();
 sg13g2_decap_4 FILLER_42_504 ();
 sg13g2_fill_2 FILLER_42_508 ();
 sg13g2_decap_4 FILLER_42_523 ();
 sg13g2_fill_1 FILLER_42_527 ();
 sg13g2_decap_4 FILLER_42_533 ();
 sg13g2_fill_1 FILLER_42_537 ();
 sg13g2_decap_8 FILLER_42_542 ();
 sg13g2_decap_8 FILLER_42_549 ();
 sg13g2_decap_8 FILLER_42_556 ();
 sg13g2_decap_8 FILLER_42_563 ();
 sg13g2_decap_4 FILLER_42_570 ();
 sg13g2_fill_2 FILLER_42_574 ();
 sg13g2_decap_8 FILLER_42_581 ();
 sg13g2_decap_8 FILLER_42_588 ();
 sg13g2_decap_8 FILLER_42_595 ();
 sg13g2_decap_8 FILLER_42_602 ();
 sg13g2_decap_8 FILLER_42_609 ();
 sg13g2_decap_8 FILLER_42_616 ();
 sg13g2_decap_8 FILLER_42_623 ();
 sg13g2_decap_8 FILLER_42_630 ();
 sg13g2_decap_8 FILLER_42_637 ();
 sg13g2_decap_8 FILLER_42_644 ();
 sg13g2_decap_8 FILLER_42_651 ();
 sg13g2_decap_8 FILLER_42_658 ();
 sg13g2_decap_8 FILLER_42_665 ();
 sg13g2_decap_8 FILLER_42_672 ();
 sg13g2_decap_8 FILLER_42_679 ();
 sg13g2_decap_8 FILLER_42_686 ();
 sg13g2_decap_8 FILLER_42_693 ();
 sg13g2_decap_8 FILLER_42_700 ();
 sg13g2_decap_8 FILLER_42_707 ();
 sg13g2_decap_8 FILLER_42_714 ();
 sg13g2_decap_8 FILLER_42_721 ();
 sg13g2_decap_8 FILLER_42_728 ();
 sg13g2_decap_8 FILLER_42_735 ();
 sg13g2_decap_8 FILLER_42_742 ();
 sg13g2_decap_8 FILLER_42_749 ();
 sg13g2_decap_8 FILLER_42_756 ();
 sg13g2_decap_8 FILLER_42_763 ();
 sg13g2_decap_8 FILLER_42_770 ();
 sg13g2_decap_8 FILLER_42_777 ();
 sg13g2_decap_8 FILLER_42_784 ();
 sg13g2_decap_8 FILLER_42_791 ();
 sg13g2_decap_8 FILLER_42_798 ();
 sg13g2_decap_8 FILLER_42_805 ();
 sg13g2_decap_8 FILLER_42_812 ();
 sg13g2_decap_8 FILLER_42_819 ();
 sg13g2_decap_8 FILLER_42_826 ();
 sg13g2_decap_8 FILLER_42_833 ();
 sg13g2_decap_8 FILLER_42_840 ();
 sg13g2_decap_8 FILLER_42_847 ();
 sg13g2_decap_8 FILLER_42_854 ();
 sg13g2_fill_1 FILLER_42_861 ();
 sg13g2_decap_8 FILLER_43_37 ();
 sg13g2_fill_2 FILLER_43_49 ();
 sg13g2_decap_4 FILLER_43_97 ();
 sg13g2_fill_2 FILLER_43_101 ();
 sg13g2_decap_4 FILLER_43_107 ();
 sg13g2_fill_2 FILLER_43_148 ();
 sg13g2_fill_1 FILLER_43_150 ();
 sg13g2_decap_4 FILLER_43_155 ();
 sg13g2_fill_1 FILLER_43_195 ();
 sg13g2_fill_1 FILLER_43_215 ();
 sg13g2_fill_1 FILLER_43_275 ();
 sg13g2_fill_1 FILLER_43_289 ();
 sg13g2_fill_2 FILLER_43_294 ();
 sg13g2_fill_2 FILLER_43_306 ();
 sg13g2_fill_1 FILLER_43_308 ();
 sg13g2_fill_1 FILLER_43_318 ();
 sg13g2_fill_2 FILLER_43_323 ();
 sg13g2_decap_4 FILLER_43_332 ();
 sg13g2_fill_2 FILLER_43_336 ();
 sg13g2_fill_2 FILLER_43_353 ();
 sg13g2_fill_2 FILLER_43_398 ();
 sg13g2_decap_4 FILLER_43_421 ();
 sg13g2_fill_1 FILLER_43_425 ();
 sg13g2_decap_8 FILLER_43_435 ();
 sg13g2_decap_4 FILLER_43_442 ();
 sg13g2_fill_2 FILLER_43_446 ();
 sg13g2_decap_4 FILLER_43_452 ();
 sg13g2_fill_1 FILLER_43_456 ();
 sg13g2_decap_4 FILLER_43_476 ();
 sg13g2_fill_1 FILLER_43_480 ();
 sg13g2_fill_2 FILLER_43_491 ();
 sg13g2_decap_4 FILLER_43_558 ();
 sg13g2_decap_8 FILLER_43_588 ();
 sg13g2_decap_8 FILLER_43_595 ();
 sg13g2_decap_8 FILLER_43_602 ();
 sg13g2_decap_8 FILLER_43_609 ();
 sg13g2_decap_8 FILLER_43_616 ();
 sg13g2_decap_8 FILLER_43_623 ();
 sg13g2_decap_8 FILLER_43_630 ();
 sg13g2_decap_8 FILLER_43_637 ();
 sg13g2_decap_8 FILLER_43_644 ();
 sg13g2_decap_8 FILLER_43_651 ();
 sg13g2_decap_8 FILLER_43_658 ();
 sg13g2_decap_8 FILLER_43_665 ();
 sg13g2_decap_8 FILLER_43_672 ();
 sg13g2_decap_8 FILLER_43_679 ();
 sg13g2_decap_8 FILLER_43_686 ();
 sg13g2_decap_8 FILLER_43_693 ();
 sg13g2_decap_8 FILLER_43_700 ();
 sg13g2_decap_8 FILLER_43_707 ();
 sg13g2_decap_8 FILLER_43_714 ();
 sg13g2_decap_8 FILLER_43_721 ();
 sg13g2_decap_8 FILLER_43_728 ();
 sg13g2_decap_8 FILLER_43_735 ();
 sg13g2_decap_8 FILLER_43_742 ();
 sg13g2_decap_8 FILLER_43_749 ();
 sg13g2_decap_8 FILLER_43_756 ();
 sg13g2_decap_8 FILLER_43_763 ();
 sg13g2_decap_8 FILLER_43_770 ();
 sg13g2_decap_8 FILLER_43_777 ();
 sg13g2_decap_8 FILLER_43_784 ();
 sg13g2_decap_8 FILLER_43_791 ();
 sg13g2_decap_8 FILLER_43_798 ();
 sg13g2_decap_8 FILLER_43_805 ();
 sg13g2_decap_8 FILLER_43_812 ();
 sg13g2_decap_8 FILLER_43_819 ();
 sg13g2_decap_8 FILLER_43_826 ();
 sg13g2_decap_8 FILLER_43_833 ();
 sg13g2_decap_8 FILLER_43_840 ();
 sg13g2_decap_8 FILLER_43_847 ();
 sg13g2_decap_8 FILLER_43_854 ();
 sg13g2_fill_1 FILLER_43_861 ();
 sg13g2_decap_4 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_4 ();
 sg13g2_fill_1 FILLER_44_24 ();
 sg13g2_decap_4 FILLER_44_51 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_fill_1 FILLER_44_91 ();
 sg13g2_fill_1 FILLER_44_148 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_fill_2 FILLER_44_161 ();
 sg13g2_fill_1 FILLER_44_163 ();
 sg13g2_fill_2 FILLER_44_225 ();
 sg13g2_fill_1 FILLER_44_227 ();
 sg13g2_fill_2 FILLER_44_241 ();
 sg13g2_decap_8 FILLER_44_270 ();
 sg13g2_decap_4 FILLER_44_277 ();
 sg13g2_fill_1 FILLER_44_285 ();
 sg13g2_decap_4 FILLER_44_306 ();
 sg13g2_fill_2 FILLER_44_361 ();
 sg13g2_fill_2 FILLER_44_381 ();
 sg13g2_fill_1 FILLER_44_383 ();
 sg13g2_decap_8 FILLER_44_393 ();
 sg13g2_fill_2 FILLER_44_400 ();
 sg13g2_fill_1 FILLER_44_402 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_4 FILLER_44_419 ();
 sg13g2_fill_2 FILLER_44_423 ();
 sg13g2_decap_4 FILLER_44_455 ();
 sg13g2_fill_1 FILLER_44_459 ();
 sg13g2_decap_4 FILLER_44_474 ();
 sg13g2_fill_1 FILLER_44_478 ();
 sg13g2_decap_4 FILLER_44_495 ();
 sg13g2_fill_1 FILLER_44_514 ();
 sg13g2_decap_4 FILLER_44_523 ();
 sg13g2_fill_2 FILLER_44_542 ();
 sg13g2_fill_2 FILLER_44_590 ();
 sg13g2_decap_4 FILLER_44_618 ();
 sg13g2_fill_2 FILLER_44_622 ();
 sg13g2_decap_8 FILLER_44_630 ();
 sg13g2_decap_8 FILLER_44_637 ();
 sg13g2_decap_8 FILLER_44_644 ();
 sg13g2_decap_8 FILLER_44_651 ();
 sg13g2_decap_8 FILLER_44_658 ();
 sg13g2_decap_8 FILLER_44_665 ();
 sg13g2_decap_8 FILLER_44_672 ();
 sg13g2_decap_8 FILLER_44_679 ();
 sg13g2_decap_8 FILLER_44_686 ();
 sg13g2_decap_8 FILLER_44_693 ();
 sg13g2_decap_8 FILLER_44_700 ();
 sg13g2_decap_8 FILLER_44_707 ();
 sg13g2_decap_8 FILLER_44_714 ();
 sg13g2_decap_8 FILLER_44_721 ();
 sg13g2_decap_8 FILLER_44_728 ();
 sg13g2_decap_8 FILLER_44_735 ();
 sg13g2_decap_8 FILLER_44_742 ();
 sg13g2_decap_8 FILLER_44_749 ();
 sg13g2_decap_8 FILLER_44_756 ();
 sg13g2_decap_8 FILLER_44_763 ();
 sg13g2_decap_8 FILLER_44_770 ();
 sg13g2_decap_8 FILLER_44_777 ();
 sg13g2_decap_8 FILLER_44_784 ();
 sg13g2_decap_8 FILLER_44_791 ();
 sg13g2_decap_8 FILLER_44_798 ();
 sg13g2_decap_8 FILLER_44_805 ();
 sg13g2_decap_8 FILLER_44_812 ();
 sg13g2_decap_8 FILLER_44_819 ();
 sg13g2_decap_8 FILLER_44_826 ();
 sg13g2_decap_8 FILLER_44_833 ();
 sg13g2_decap_8 FILLER_44_840 ();
 sg13g2_decap_8 FILLER_44_847 ();
 sg13g2_decap_8 FILLER_44_854 ();
 sg13g2_fill_1 FILLER_44_861 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_fill_1 FILLER_45_14 ();
 sg13g2_decap_4 FILLER_45_23 ();
 sg13g2_fill_2 FILLER_45_27 ();
 sg13g2_fill_1 FILLER_45_71 ();
 sg13g2_fill_2 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_113 ();
 sg13g2_decap_4 FILLER_45_120 ();
 sg13g2_fill_1 FILLER_45_124 ();
 sg13g2_fill_2 FILLER_45_138 ();
 sg13g2_fill_1 FILLER_45_140 ();
 sg13g2_fill_2 FILLER_45_167 ();
 sg13g2_fill_1 FILLER_45_169 ();
 sg13g2_fill_2 FILLER_45_205 ();
 sg13g2_fill_2 FILLER_45_268 ();
 sg13g2_fill_1 FILLER_45_319 ();
 sg13g2_fill_2 FILLER_45_330 ();
 sg13g2_fill_1 FILLER_45_332 ();
 sg13g2_decap_4 FILLER_45_347 ();
 sg13g2_fill_1 FILLER_45_351 ();
 sg13g2_fill_1 FILLER_45_376 ();
 sg13g2_fill_1 FILLER_45_382 ();
 sg13g2_fill_1 FILLER_45_416 ();
 sg13g2_decap_8 FILLER_45_462 ();
 sg13g2_fill_2 FILLER_45_495 ();
 sg13g2_decap_8 FILLER_45_506 ();
 sg13g2_fill_1 FILLER_45_513 ();
 sg13g2_fill_1 FILLER_45_518 ();
 sg13g2_decap_4 FILLER_45_528 ();
 sg13g2_fill_2 FILLER_45_532 ();
 sg13g2_fill_1 FILLER_45_553 ();
 sg13g2_fill_2 FILLER_45_571 ();
 sg13g2_fill_2 FILLER_45_607 ();
 sg13g2_decap_8 FILLER_45_631 ();
 sg13g2_decap_8 FILLER_45_638 ();
 sg13g2_decap_8 FILLER_45_645 ();
 sg13g2_decap_8 FILLER_45_652 ();
 sg13g2_decap_8 FILLER_45_659 ();
 sg13g2_decap_8 FILLER_45_666 ();
 sg13g2_decap_8 FILLER_45_673 ();
 sg13g2_decap_8 FILLER_45_680 ();
 sg13g2_decap_8 FILLER_45_687 ();
 sg13g2_decap_8 FILLER_45_694 ();
 sg13g2_decap_8 FILLER_45_701 ();
 sg13g2_decap_8 FILLER_45_708 ();
 sg13g2_decap_8 FILLER_45_715 ();
 sg13g2_decap_8 FILLER_45_722 ();
 sg13g2_decap_8 FILLER_45_729 ();
 sg13g2_decap_8 FILLER_45_736 ();
 sg13g2_decap_8 FILLER_45_743 ();
 sg13g2_decap_8 FILLER_45_750 ();
 sg13g2_decap_8 FILLER_45_757 ();
 sg13g2_decap_8 FILLER_45_764 ();
 sg13g2_decap_8 FILLER_45_771 ();
 sg13g2_decap_8 FILLER_45_778 ();
 sg13g2_decap_8 FILLER_45_785 ();
 sg13g2_decap_8 FILLER_45_792 ();
 sg13g2_decap_8 FILLER_45_799 ();
 sg13g2_decap_8 FILLER_45_806 ();
 sg13g2_decap_8 FILLER_45_813 ();
 sg13g2_decap_8 FILLER_45_820 ();
 sg13g2_decap_8 FILLER_45_827 ();
 sg13g2_decap_8 FILLER_45_834 ();
 sg13g2_decap_8 FILLER_45_841 ();
 sg13g2_decap_8 FILLER_45_848 ();
 sg13g2_decap_8 FILLER_45_855 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_2 ();
 sg13g2_fill_2 FILLER_46_82 ();
 sg13g2_fill_1 FILLER_46_96 ();
 sg13g2_fill_1 FILLER_46_101 ();
 sg13g2_decap_8 FILLER_46_165 ();
 sg13g2_fill_1 FILLER_46_172 ();
 sg13g2_fill_1 FILLER_46_231 ();
 sg13g2_fill_1 FILLER_46_265 ();
 sg13g2_fill_1 FILLER_46_284 ();
 sg13g2_fill_2 FILLER_46_294 ();
 sg13g2_fill_1 FILLER_46_296 ();
 sg13g2_fill_2 FILLER_46_322 ();
 sg13g2_fill_2 FILLER_46_333 ();
 sg13g2_fill_1 FILLER_46_349 ();
 sg13g2_fill_2 FILLER_46_362 ();
 sg13g2_fill_1 FILLER_46_364 ();
 sg13g2_fill_1 FILLER_46_398 ();
 sg13g2_fill_1 FILLER_46_411 ();
 sg13g2_decap_4 FILLER_46_416 ();
 sg13g2_fill_2 FILLER_46_420 ();
 sg13g2_fill_1 FILLER_46_432 ();
 sg13g2_decap_8 FILLER_46_443 ();
 sg13g2_fill_2 FILLER_46_450 ();
 sg13g2_fill_1 FILLER_46_452 ();
 sg13g2_fill_2 FILLER_46_483 ();
 sg13g2_fill_1 FILLER_46_485 ();
 sg13g2_fill_2 FILLER_46_517 ();
 sg13g2_decap_4 FILLER_46_524 ();
 sg13g2_fill_2 FILLER_46_540 ();
 sg13g2_fill_1 FILLER_46_542 ();
 sg13g2_fill_1 FILLER_46_564 ();
 sg13g2_fill_1 FILLER_46_584 ();
 sg13g2_fill_2 FILLER_46_612 ();
 sg13g2_decap_8 FILLER_46_640 ();
 sg13g2_decap_8 FILLER_46_647 ();
 sg13g2_decap_8 FILLER_46_654 ();
 sg13g2_decap_8 FILLER_46_661 ();
 sg13g2_decap_8 FILLER_46_668 ();
 sg13g2_decap_8 FILLER_46_675 ();
 sg13g2_decap_8 FILLER_46_682 ();
 sg13g2_decap_8 FILLER_46_689 ();
 sg13g2_decap_8 FILLER_46_696 ();
 sg13g2_decap_8 FILLER_46_703 ();
 sg13g2_decap_8 FILLER_46_710 ();
 sg13g2_decap_8 FILLER_46_717 ();
 sg13g2_decap_8 FILLER_46_724 ();
 sg13g2_decap_8 FILLER_46_731 ();
 sg13g2_decap_8 FILLER_46_738 ();
 sg13g2_decap_8 FILLER_46_745 ();
 sg13g2_decap_8 FILLER_46_752 ();
 sg13g2_decap_8 FILLER_46_759 ();
 sg13g2_decap_8 FILLER_46_766 ();
 sg13g2_decap_8 FILLER_46_773 ();
 sg13g2_decap_8 FILLER_46_780 ();
 sg13g2_decap_8 FILLER_46_787 ();
 sg13g2_decap_8 FILLER_46_794 ();
 sg13g2_decap_8 FILLER_46_801 ();
 sg13g2_decap_8 FILLER_46_808 ();
 sg13g2_decap_8 FILLER_46_815 ();
 sg13g2_decap_8 FILLER_46_822 ();
 sg13g2_decap_8 FILLER_46_829 ();
 sg13g2_decap_8 FILLER_46_836 ();
 sg13g2_decap_8 FILLER_46_843 ();
 sg13g2_decap_8 FILLER_46_850 ();
 sg13g2_decap_4 FILLER_46_857 ();
 sg13g2_fill_1 FILLER_46_861 ();
 sg13g2_fill_2 FILLER_47_40 ();
 sg13g2_fill_1 FILLER_47_58 ();
 sg13g2_decap_4 FILLER_47_74 ();
 sg13g2_decap_8 FILLER_47_108 ();
 sg13g2_fill_2 FILLER_47_115 ();
 sg13g2_fill_1 FILLER_47_117 ();
 sg13g2_decap_4 FILLER_47_122 ();
 sg13g2_fill_2 FILLER_47_152 ();
 sg13g2_fill_1 FILLER_47_154 ();
 sg13g2_fill_2 FILLER_47_198 ();
 sg13g2_fill_2 FILLER_47_236 ();
 sg13g2_fill_1 FILLER_47_251 ();
 sg13g2_fill_1 FILLER_47_297 ();
 sg13g2_decap_4 FILLER_47_353 ();
 sg13g2_fill_2 FILLER_47_357 ();
 sg13g2_decap_8 FILLER_47_363 ();
 sg13g2_decap_4 FILLER_47_370 ();
 sg13g2_fill_1 FILLER_47_379 ();
 sg13g2_decap_8 FILLER_47_387 ();
 sg13g2_fill_2 FILLER_47_394 ();
 sg13g2_fill_1 FILLER_47_396 ();
 sg13g2_decap_4 FILLER_47_420 ();
 sg13g2_decap_4 FILLER_47_430 ();
 sg13g2_fill_1 FILLER_47_434 ();
 sg13g2_fill_2 FILLER_47_454 ();
 sg13g2_fill_1 FILLER_47_456 ();
 sg13g2_decap_4 FILLER_47_467 ();
 sg13g2_fill_2 FILLER_47_499 ();
 sg13g2_fill_1 FILLER_47_515 ();
 sg13g2_fill_1 FILLER_47_525 ();
 sg13g2_decap_4 FILLER_47_538 ();
 sg13g2_fill_2 FILLER_47_542 ();
 sg13g2_decap_4 FILLER_47_549 ();
 sg13g2_fill_2 FILLER_47_553 ();
 sg13g2_fill_2 FILLER_47_563 ();
 sg13g2_fill_1 FILLER_47_565 ();
 sg13g2_decap_4 FILLER_47_587 ();
 sg13g2_fill_1 FILLER_47_591 ();
 sg13g2_fill_1 FILLER_47_597 ();
 sg13g2_decap_4 FILLER_47_613 ();
 sg13g2_fill_2 FILLER_47_617 ();
 sg13g2_decap_8 FILLER_47_637 ();
 sg13g2_decap_8 FILLER_47_644 ();
 sg13g2_decap_8 FILLER_47_651 ();
 sg13g2_decap_8 FILLER_47_658 ();
 sg13g2_decap_8 FILLER_47_665 ();
 sg13g2_decap_8 FILLER_47_672 ();
 sg13g2_decap_8 FILLER_47_679 ();
 sg13g2_decap_8 FILLER_47_686 ();
 sg13g2_decap_8 FILLER_47_693 ();
 sg13g2_decap_8 FILLER_47_700 ();
 sg13g2_decap_8 FILLER_47_707 ();
 sg13g2_decap_8 FILLER_47_714 ();
 sg13g2_fill_2 FILLER_47_721 ();
 sg13g2_fill_1 FILLER_47_723 ();
 sg13g2_decap_8 FILLER_47_727 ();
 sg13g2_decap_8 FILLER_47_734 ();
 sg13g2_decap_8 FILLER_47_741 ();
 sg13g2_decap_8 FILLER_47_748 ();
 sg13g2_decap_8 FILLER_47_755 ();
 sg13g2_decap_8 FILLER_47_762 ();
 sg13g2_decap_8 FILLER_47_769 ();
 sg13g2_decap_8 FILLER_47_776 ();
 sg13g2_decap_8 FILLER_47_783 ();
 sg13g2_decap_8 FILLER_47_790 ();
 sg13g2_decap_8 FILLER_47_797 ();
 sg13g2_decap_8 FILLER_47_804 ();
 sg13g2_decap_8 FILLER_47_811 ();
 sg13g2_decap_8 FILLER_47_818 ();
 sg13g2_decap_8 FILLER_47_825 ();
 sg13g2_decap_8 FILLER_47_832 ();
 sg13g2_decap_8 FILLER_47_839 ();
 sg13g2_decap_8 FILLER_47_846 ();
 sg13g2_decap_8 FILLER_47_853 ();
 sg13g2_fill_2 FILLER_47_860 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_4 FILLER_48_7 ();
 sg13g2_fill_1 FILLER_48_29 ();
 sg13g2_fill_2 FILLER_48_40 ();
 sg13g2_fill_1 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_48 ();
 sg13g2_decap_8 FILLER_48_55 ();
 sg13g2_decap_4 FILLER_48_62 ();
 sg13g2_fill_1 FILLER_48_66 ();
 sg13g2_fill_2 FILLER_48_72 ();
 sg13g2_fill_1 FILLER_48_74 ();
 sg13g2_fill_2 FILLER_48_95 ();
 sg13g2_fill_1 FILLER_48_97 ();
 sg13g2_fill_2 FILLER_48_116 ();
 sg13g2_fill_2 FILLER_48_160 ();
 sg13g2_fill_1 FILLER_48_162 ();
 sg13g2_fill_2 FILLER_48_207 ();
 sg13g2_fill_2 FILLER_48_222 ();
 sg13g2_fill_2 FILLER_48_243 ();
 sg13g2_fill_1 FILLER_48_245 ();
 sg13g2_fill_1 FILLER_48_260 ();
 sg13g2_fill_1 FILLER_48_266 ();
 sg13g2_fill_2 FILLER_48_336 ();
 sg13g2_decap_8 FILLER_48_342 ();
 sg13g2_fill_2 FILLER_48_359 ();
 sg13g2_decap_4 FILLER_48_393 ();
 sg13g2_fill_2 FILLER_48_397 ();
 sg13g2_decap_8 FILLER_48_414 ();
 sg13g2_fill_2 FILLER_48_421 ();
 sg13g2_fill_1 FILLER_48_423 ();
 sg13g2_fill_2 FILLER_48_432 ();
 sg13g2_decap_8 FILLER_48_438 ();
 sg13g2_decap_8 FILLER_48_445 ();
 sg13g2_decap_8 FILLER_48_452 ();
 sg13g2_decap_4 FILLER_48_459 ();
 sg13g2_decap_8 FILLER_48_515 ();
 sg13g2_decap_4 FILLER_48_539 ();
 sg13g2_fill_2 FILLER_48_549 ();
 sg13g2_decap_8 FILLER_48_559 ();
 sg13g2_fill_1 FILLER_48_566 ();
 sg13g2_fill_2 FILLER_48_589 ();
 sg13g2_fill_1 FILLER_48_627 ();
 sg13g2_decap_8 FILLER_48_637 ();
 sg13g2_decap_8 FILLER_48_644 ();
 sg13g2_decap_8 FILLER_48_651 ();
 sg13g2_decap_8 FILLER_48_658 ();
 sg13g2_decap_8 FILLER_48_665 ();
 sg13g2_decap_8 FILLER_48_672 ();
 sg13g2_decap_4 FILLER_48_679 ();
 sg13g2_fill_2 FILLER_48_683 ();
 sg13g2_decap_8 FILLER_48_695 ();
 sg13g2_fill_1 FILLER_48_702 ();
 sg13g2_decap_8 FILLER_48_706 ();
 sg13g2_decap_4 FILLER_48_713 ();
 sg13g2_fill_1 FILLER_48_717 ();
 sg13g2_fill_2 FILLER_48_723 ();
 sg13g2_decap_8 FILLER_48_738 ();
 sg13g2_decap_8 FILLER_48_745 ();
 sg13g2_decap_8 FILLER_48_752 ();
 sg13g2_decap_8 FILLER_48_759 ();
 sg13g2_decap_8 FILLER_48_766 ();
 sg13g2_decap_8 FILLER_48_773 ();
 sg13g2_decap_8 FILLER_48_780 ();
 sg13g2_decap_8 FILLER_48_787 ();
 sg13g2_decap_8 FILLER_48_794 ();
 sg13g2_decap_8 FILLER_48_801 ();
 sg13g2_decap_8 FILLER_48_808 ();
 sg13g2_decap_8 FILLER_48_815 ();
 sg13g2_decap_8 FILLER_48_822 ();
 sg13g2_decap_8 FILLER_48_829 ();
 sg13g2_decap_8 FILLER_48_836 ();
 sg13g2_decap_8 FILLER_48_843 ();
 sg13g2_decap_8 FILLER_48_850 ();
 sg13g2_decap_4 FILLER_48_857 ();
 sg13g2_fill_1 FILLER_48_861 ();
 sg13g2_decap_4 FILLER_49_26 ();
 sg13g2_fill_2 FILLER_49_46 ();
 sg13g2_fill_1 FILLER_49_48 ();
 sg13g2_fill_2 FILLER_49_92 ();
 sg13g2_fill_1 FILLER_49_94 ();
 sg13g2_fill_1 FILLER_49_100 ();
 sg13g2_fill_1 FILLER_49_115 ();
 sg13g2_fill_2 FILLER_49_121 ();
 sg13g2_fill_1 FILLER_49_123 ();
 sg13g2_fill_2 FILLER_49_129 ();
 sg13g2_fill_2 FILLER_49_161 ();
 sg13g2_fill_1 FILLER_49_163 ();
 sg13g2_fill_2 FILLER_49_225 ();
 sg13g2_fill_1 FILLER_49_227 ();
 sg13g2_fill_1 FILLER_49_252 ();
 sg13g2_fill_1 FILLER_49_266 ();
 sg13g2_fill_2 FILLER_49_279 ();
 sg13g2_decap_8 FILLER_49_338 ();
 sg13g2_decap_4 FILLER_49_345 ();
 sg13g2_fill_1 FILLER_49_349 ();
 sg13g2_fill_1 FILLER_49_355 ();
 sg13g2_fill_1 FILLER_49_360 ();
 sg13g2_decap_4 FILLER_49_369 ();
 sg13g2_fill_2 FILLER_49_381 ();
 sg13g2_fill_1 FILLER_49_383 ();
 sg13g2_fill_1 FILLER_49_389 ();
 sg13g2_fill_1 FILLER_49_395 ();
 sg13g2_decap_4 FILLER_49_400 ();
 sg13g2_fill_1 FILLER_49_404 ();
 sg13g2_fill_2 FILLER_49_434 ();
 sg13g2_decap_8 FILLER_49_482 ();
 sg13g2_fill_2 FILLER_49_489 ();
 sg13g2_fill_1 FILLER_49_491 ();
 sg13g2_decap_8 FILLER_49_496 ();
 sg13g2_decap_4 FILLER_49_503 ();
 sg13g2_decap_4 FILLER_49_513 ();
 sg13g2_fill_2 FILLER_49_517 ();
 sg13g2_fill_1 FILLER_49_529 ();
 sg13g2_decap_8 FILLER_49_586 ();
 sg13g2_decap_4 FILLER_49_593 ();
 sg13g2_fill_1 FILLER_49_597 ();
 sg13g2_fill_2 FILLER_49_602 ();
 sg13g2_fill_2 FILLER_49_622 ();
 sg13g2_decap_8 FILLER_49_647 ();
 sg13g2_decap_8 FILLER_49_654 ();
 sg13g2_decap_8 FILLER_49_661 ();
 sg13g2_decap_8 FILLER_49_668 ();
 sg13g2_fill_1 FILLER_49_675 ();
 sg13g2_fill_1 FILLER_49_702 ();
 sg13g2_fill_2 FILLER_49_721 ();
 sg13g2_decap_8 FILLER_49_752 ();
 sg13g2_decap_8 FILLER_49_759 ();
 sg13g2_fill_2 FILLER_49_766 ();
 sg13g2_fill_1 FILLER_49_768 ();
 sg13g2_decap_8 FILLER_49_772 ();
 sg13g2_decap_8 FILLER_49_779 ();
 sg13g2_decap_8 FILLER_49_786 ();
 sg13g2_decap_8 FILLER_49_793 ();
 sg13g2_decap_8 FILLER_49_800 ();
 sg13g2_decap_8 FILLER_49_807 ();
 sg13g2_decap_8 FILLER_49_814 ();
 sg13g2_decap_8 FILLER_49_821 ();
 sg13g2_decap_8 FILLER_49_828 ();
 sg13g2_decap_8 FILLER_49_835 ();
 sg13g2_decap_8 FILLER_49_842 ();
 sg13g2_decap_8 FILLER_49_849 ();
 sg13g2_decap_4 FILLER_49_856 ();
 sg13g2_fill_2 FILLER_49_860 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_4 FILLER_50_7 ();
 sg13g2_fill_2 FILLER_50_15 ();
 sg13g2_fill_2 FILLER_50_26 ();
 sg13g2_fill_1 FILLER_50_33 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_4 FILLER_50_56 ();
 sg13g2_fill_2 FILLER_50_64 ();
 sg13g2_decap_8 FILLER_50_76 ();
 sg13g2_fill_1 FILLER_50_83 ();
 sg13g2_fill_2 FILLER_50_95 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_decap_4 FILLER_50_119 ();
 sg13g2_fill_1 FILLER_50_123 ();
 sg13g2_fill_2 FILLER_50_128 ();
 sg13g2_fill_1 FILLER_50_173 ();
 sg13g2_fill_2 FILLER_50_184 ();
 sg13g2_fill_2 FILLER_50_196 ();
 sg13g2_fill_2 FILLER_50_225 ();
 sg13g2_fill_1 FILLER_50_227 ();
 sg13g2_decap_4 FILLER_50_238 ();
 sg13g2_fill_2 FILLER_50_282 ();
 sg13g2_fill_1 FILLER_50_302 ();
 sg13g2_fill_2 FILLER_50_321 ();
 sg13g2_decap_4 FILLER_50_348 ();
 sg13g2_decap_8 FILLER_50_360 ();
 sg13g2_fill_1 FILLER_50_380 ();
 sg13g2_fill_1 FILLER_50_395 ();
 sg13g2_decap_8 FILLER_50_409 ();
 sg13g2_decap_8 FILLER_50_416 ();
 sg13g2_fill_2 FILLER_50_423 ();
 sg13g2_fill_1 FILLER_50_425 ();
 sg13g2_fill_1 FILLER_50_432 ();
 sg13g2_decap_8 FILLER_50_444 ();
 sg13g2_fill_1 FILLER_50_451 ();
 sg13g2_fill_2 FILLER_50_465 ();
 sg13g2_fill_1 FILLER_50_472 ();
 sg13g2_fill_1 FILLER_50_482 ();
 sg13g2_fill_2 FILLER_50_499 ();
 sg13g2_fill_2 FILLER_50_533 ();
 sg13g2_fill_2 FILLER_50_540 ();
 sg13g2_fill_2 FILLER_50_547 ();
 sg13g2_fill_1 FILLER_50_549 ();
 sg13g2_fill_2 FILLER_50_555 ();
 sg13g2_fill_1 FILLER_50_557 ();
 sg13g2_fill_1 FILLER_50_589 ();
 sg13g2_fill_2 FILLER_50_598 ();
 sg13g2_fill_1 FILLER_50_600 ();
 sg13g2_decap_8 FILLER_50_612 ();
 sg13g2_fill_2 FILLER_50_623 ();
 sg13g2_decap_4 FILLER_50_646 ();
 sg13g2_fill_2 FILLER_50_650 ();
 sg13g2_decap_4 FILLER_50_675 ();
 sg13g2_fill_2 FILLER_50_679 ();
 sg13g2_decap_4 FILLER_50_759 ();
 sg13g2_fill_1 FILLER_50_763 ();
 sg13g2_fill_1 FILLER_50_769 ();
 sg13g2_decap_4 FILLER_50_783 ();
 sg13g2_decap_8 FILLER_50_813 ();
 sg13g2_decap_8 FILLER_50_820 ();
 sg13g2_decap_8 FILLER_50_827 ();
 sg13g2_decap_8 FILLER_50_834 ();
 sg13g2_decap_8 FILLER_50_841 ();
 sg13g2_decap_8 FILLER_50_848 ();
 sg13g2_decap_8 FILLER_50_855 ();
 sg13g2_fill_2 FILLER_51_26 ();
 sg13g2_fill_2 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_61 ();
 sg13g2_fill_1 FILLER_51_68 ();
 sg13g2_fill_2 FILLER_51_74 ();
 sg13g2_fill_1 FILLER_51_112 ();
 sg13g2_fill_2 FILLER_51_148 ();
 sg13g2_decap_8 FILLER_51_240 ();
 sg13g2_fill_2 FILLER_51_247 ();
 sg13g2_fill_1 FILLER_51_249 ();
 sg13g2_fill_1 FILLER_51_277 ();
 sg13g2_fill_1 FILLER_51_291 ();
 sg13g2_fill_2 FILLER_51_342 ();
 sg13g2_fill_1 FILLER_51_344 ();
 sg13g2_fill_1 FILLER_51_388 ();
 sg13g2_fill_2 FILLER_51_400 ();
 sg13g2_fill_1 FILLER_51_413 ();
 sg13g2_fill_2 FILLER_51_429 ();
 sg13g2_fill_1 FILLER_51_431 ();
 sg13g2_decap_4 FILLER_51_438 ();
 sg13g2_decap_4 FILLER_51_447 ();
 sg13g2_fill_1 FILLER_51_451 ();
 sg13g2_decap_4 FILLER_51_465 ();
 sg13g2_fill_1 FILLER_51_478 ();
 sg13g2_fill_2 FILLER_51_510 ();
 sg13g2_decap_4 FILLER_51_532 ();
 sg13g2_decap_8 FILLER_51_555 ();
 sg13g2_fill_1 FILLER_51_562 ();
 sg13g2_decap_8 FILLER_51_577 ();
 sg13g2_fill_1 FILLER_51_584 ();
 sg13g2_fill_1 FILLER_51_617 ();
 sg13g2_decap_8 FILLER_51_644 ();
 sg13g2_fill_2 FILLER_51_651 ();
 sg13g2_fill_1 FILLER_51_653 ();
 sg13g2_fill_2 FILLER_51_664 ();
 sg13g2_fill_1 FILLER_51_686 ();
 sg13g2_decap_4 FILLER_51_706 ();
 sg13g2_fill_1 FILLER_51_710 ();
 sg13g2_fill_1 FILLER_51_809 ();
 sg13g2_decap_8 FILLER_51_819 ();
 sg13g2_decap_8 FILLER_51_826 ();
 sg13g2_decap_8 FILLER_51_833 ();
 sg13g2_decap_8 FILLER_51_840 ();
 sg13g2_decap_8 FILLER_51_847 ();
 sg13g2_decap_8 FILLER_51_854 ();
 sg13g2_fill_1 FILLER_51_861 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_4 FILLER_52_7 ();
 sg13g2_decap_4 FILLER_52_24 ();
 sg13g2_decap_4 FILLER_52_43 ();
 sg13g2_fill_2 FILLER_52_77 ();
 sg13g2_fill_2 FILLER_52_93 ();
 sg13g2_fill_1 FILLER_52_95 ();
 sg13g2_fill_2 FILLER_52_131 ();
 sg13g2_fill_2 FILLER_52_171 ();
 sg13g2_fill_1 FILLER_52_202 ();
 sg13g2_fill_2 FILLER_52_211 ();
 sg13g2_fill_2 FILLER_52_241 ();
 sg13g2_fill_1 FILLER_52_243 ();
 sg13g2_decap_8 FILLER_52_255 ();
 sg13g2_decap_8 FILLER_52_291 ();
 sg13g2_fill_2 FILLER_52_298 ();
 sg13g2_fill_1 FILLER_52_300 ();
 sg13g2_fill_1 FILLER_52_327 ();
 sg13g2_decap_4 FILLER_52_364 ();
 sg13g2_fill_1 FILLER_52_368 ();
 sg13g2_fill_1 FILLER_52_373 ();
 sg13g2_decap_8 FILLER_52_378 ();
 sg13g2_fill_1 FILLER_52_395 ();
 sg13g2_fill_1 FILLER_52_406 ();
 sg13g2_fill_2 FILLER_52_414 ();
 sg13g2_fill_1 FILLER_52_425 ();
 sg13g2_fill_1 FILLER_52_432 ();
 sg13g2_fill_2 FILLER_52_538 ();
 sg13g2_fill_1 FILLER_52_540 ();
 sg13g2_decap_8 FILLER_52_558 ();
 sg13g2_fill_2 FILLER_52_571 ();
 sg13g2_fill_2 FILLER_52_576 ();
 sg13g2_fill_1 FILLER_52_578 ();
 sg13g2_decap_4 FILLER_52_583 ();
 sg13g2_fill_1 FILLER_52_587 ();
 sg13g2_decap_4 FILLER_52_591 ();
 sg13g2_fill_2 FILLER_52_611 ();
 sg13g2_fill_2 FILLER_52_626 ();
 sg13g2_fill_1 FILLER_52_628 ();
 sg13g2_decap_8 FILLER_52_638 ();
 sg13g2_decap_4 FILLER_52_645 ();
 sg13g2_decap_4 FILLER_52_654 ();
 sg13g2_decap_4 FILLER_52_682 ();
 sg13g2_decap_4 FILLER_52_700 ();
 sg13g2_fill_1 FILLER_52_704 ();
 sg13g2_fill_1 FILLER_52_744 ();
 sg13g2_fill_1 FILLER_52_798 ();
 sg13g2_decap_8 FILLER_52_820 ();
 sg13g2_decap_8 FILLER_52_827 ();
 sg13g2_decap_8 FILLER_52_834 ();
 sg13g2_decap_8 FILLER_52_841 ();
 sg13g2_decap_8 FILLER_52_848 ();
 sg13g2_decap_8 FILLER_52_855 ();
 sg13g2_fill_2 FILLER_53_31 ();
 sg13g2_fill_1 FILLER_53_54 ();
 sg13g2_fill_2 FILLER_53_69 ();
 sg13g2_fill_1 FILLER_53_100 ();
 sg13g2_fill_1 FILLER_53_131 ();
 sg13g2_decap_8 FILLER_53_172 ();
 sg13g2_decap_4 FILLER_53_179 ();
 sg13g2_decap_4 FILLER_53_193 ();
 sg13g2_fill_2 FILLER_53_197 ();
 sg13g2_decap_8 FILLER_53_213 ();
 sg13g2_fill_2 FILLER_53_220 ();
 sg13g2_decap_8 FILLER_53_242 ();
 sg13g2_fill_2 FILLER_53_249 ();
 sg13g2_fill_2 FILLER_53_269 ();
 sg13g2_fill_2 FILLER_53_294 ();
 sg13g2_fill_2 FILLER_53_306 ();
 sg13g2_fill_2 FILLER_53_338 ();
 sg13g2_fill_1 FILLER_53_358 ();
 sg13g2_decap_8 FILLER_53_398 ();
 sg13g2_fill_2 FILLER_53_405 ();
 sg13g2_decap_4 FILLER_53_429 ();
 sg13g2_decap_4 FILLER_53_437 ();
 sg13g2_fill_2 FILLER_53_441 ();
 sg13g2_fill_1 FILLER_53_453 ();
 sg13g2_fill_1 FILLER_53_485 ();
 sg13g2_decap_8 FILLER_53_495 ();
 sg13g2_decap_4 FILLER_53_502 ();
 sg13g2_fill_2 FILLER_53_506 ();
 sg13g2_fill_2 FILLER_53_512 ();
 sg13g2_fill_1 FILLER_53_514 ();
 sg13g2_fill_2 FILLER_53_556 ();
 sg13g2_fill_1 FILLER_53_558 ();
 sg13g2_fill_2 FILLER_53_586 ();
 sg13g2_fill_1 FILLER_53_588 ();
 sg13g2_fill_2 FILLER_53_610 ();
 sg13g2_fill_1 FILLER_53_612 ();
 sg13g2_decap_8 FILLER_53_654 ();
 sg13g2_fill_2 FILLER_53_661 ();
 sg13g2_decap_8 FILLER_53_668 ();
 sg13g2_fill_1 FILLER_53_675 ();
 sg13g2_fill_1 FILLER_53_680 ();
 sg13g2_fill_2 FILLER_53_706 ();
 sg13g2_fill_1 FILLER_53_708 ();
 sg13g2_fill_1 FILLER_53_726 ();
 sg13g2_fill_1 FILLER_53_764 ();
 sg13g2_decap_8 FILLER_53_833 ();
 sg13g2_decap_8 FILLER_53_840 ();
 sg13g2_decap_8 FILLER_53_847 ();
 sg13g2_decap_8 FILLER_53_854 ();
 sg13g2_fill_1 FILLER_53_861 ();
 sg13g2_decap_4 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_4 ();
 sg13g2_fill_1 FILLER_54_57 ();
 sg13g2_fill_2 FILLER_54_85 ();
 sg13g2_fill_1 FILLER_54_113 ();
 sg13g2_fill_2 FILLER_54_123 ();
 sg13g2_fill_1 FILLER_54_145 ();
 sg13g2_fill_2 FILLER_54_152 ();
 sg13g2_fill_1 FILLER_54_158 ();
 sg13g2_fill_2 FILLER_54_176 ();
 sg13g2_fill_1 FILLER_54_178 ();
 sg13g2_decap_8 FILLER_54_189 ();
 sg13g2_fill_2 FILLER_54_196 ();
 sg13g2_fill_2 FILLER_54_209 ();
 sg13g2_fill_1 FILLER_54_211 ();
 sg13g2_fill_2 FILLER_54_222 ();
 sg13g2_decap_4 FILLER_54_239 ();
 sg13g2_fill_2 FILLER_54_243 ();
 sg13g2_fill_2 FILLER_54_271 ();
 sg13g2_fill_1 FILLER_54_292 ();
 sg13g2_fill_1 FILLER_54_328 ();
 sg13g2_fill_2 FILLER_54_344 ();
 sg13g2_decap_8 FILLER_54_370 ();
 sg13g2_decap_4 FILLER_54_377 ();
 sg13g2_fill_1 FILLER_54_381 ();
 sg13g2_decap_4 FILLER_54_394 ();
 sg13g2_fill_2 FILLER_54_398 ();
 sg13g2_fill_2 FILLER_54_422 ();
 sg13g2_fill_1 FILLER_54_440 ();
 sg13g2_decap_8 FILLER_54_515 ();
 sg13g2_decap_4 FILLER_54_522 ();
 sg13g2_fill_2 FILLER_54_530 ();
 sg13g2_fill_1 FILLER_54_532 ();
 sg13g2_fill_2 FILLER_54_539 ();
 sg13g2_decap_4 FILLER_54_559 ();
 sg13g2_fill_2 FILLER_54_563 ();
 sg13g2_decap_8 FILLER_54_574 ();
 sg13g2_decap_8 FILLER_54_581 ();
 sg13g2_decap_4 FILLER_54_588 ();
 sg13g2_fill_2 FILLER_54_592 ();
 sg13g2_fill_2 FILLER_54_604 ();
 sg13g2_fill_1 FILLER_54_606 ();
 sg13g2_fill_2 FILLER_54_611 ();
 sg13g2_fill_2 FILLER_54_617 ();
 sg13g2_fill_2 FILLER_54_632 ();
 sg13g2_fill_1 FILLER_54_634 ();
 sg13g2_fill_2 FILLER_54_688 ();
 sg13g2_fill_1 FILLER_54_690 ();
 sg13g2_fill_2 FILLER_54_718 ();
 sg13g2_fill_2 FILLER_54_730 ();
 sg13g2_fill_1 FILLER_54_732 ();
 sg13g2_fill_2 FILLER_54_802 ();
 sg13g2_decap_8 FILLER_54_822 ();
 sg13g2_decap_8 FILLER_54_829 ();
 sg13g2_decap_8 FILLER_54_836 ();
 sg13g2_decap_8 FILLER_54_843 ();
 sg13g2_decap_8 FILLER_54_850 ();
 sg13g2_decap_4 FILLER_54_857 ();
 sg13g2_fill_1 FILLER_54_861 ();
 sg13g2_fill_2 FILLER_55_40 ();
 sg13g2_decap_8 FILLER_55_90 ();
 sg13g2_fill_2 FILLER_55_159 ();
 sg13g2_fill_1 FILLER_55_161 ();
 sg13g2_fill_2 FILLER_55_188 ();
 sg13g2_fill_1 FILLER_55_190 ();
 sg13g2_decap_4 FILLER_55_196 ();
 sg13g2_fill_2 FILLER_55_204 ();
 sg13g2_decap_4 FILLER_55_223 ();
 sg13g2_fill_1 FILLER_55_227 ();
 sg13g2_fill_2 FILLER_55_313 ();
 sg13g2_decap_8 FILLER_55_352 ();
 sg13g2_fill_1 FILLER_55_359 ();
 sg13g2_decap_8 FILLER_55_365 ();
 sg13g2_fill_1 FILLER_55_372 ();
 sg13g2_fill_2 FILLER_55_403 ();
 sg13g2_fill_1 FILLER_55_405 ();
 sg13g2_fill_2 FILLER_55_414 ();
 sg13g2_fill_1 FILLER_55_416 ();
 sg13g2_decap_8 FILLER_55_427 ();
 sg13g2_decap_8 FILLER_55_434 ();
 sg13g2_decap_4 FILLER_55_441 ();
 sg13g2_fill_2 FILLER_55_445 ();
 sg13g2_fill_1 FILLER_55_456 ();
 sg13g2_fill_2 FILLER_55_461 ();
 sg13g2_fill_1 FILLER_55_463 ();
 sg13g2_fill_2 FILLER_55_492 ();
 sg13g2_decap_4 FILLER_55_525 ();
 sg13g2_fill_1 FILLER_55_529 ();
 sg13g2_decap_8 FILLER_55_579 ();
 sg13g2_fill_2 FILLER_55_586 ();
 sg13g2_fill_2 FILLER_55_615 ();
 sg13g2_fill_1 FILLER_55_617 ();
 sg13g2_decap_8 FILLER_55_626 ();
 sg13g2_fill_2 FILLER_55_633 ();
 sg13g2_fill_1 FILLER_55_635 ();
 sg13g2_fill_1 FILLER_55_645 ();
 sg13g2_decap_8 FILLER_55_656 ();
 sg13g2_decap_8 FILLER_55_663 ();
 sg13g2_decap_8 FILLER_55_670 ();
 sg13g2_fill_1 FILLER_55_677 ();
 sg13g2_fill_2 FILLER_55_715 ();
 sg13g2_fill_1 FILLER_55_717 ();
 sg13g2_fill_1 FILLER_55_738 ();
 sg13g2_fill_2 FILLER_55_748 ();
 sg13g2_fill_1 FILLER_55_803 ();
 sg13g2_decap_8 FILLER_55_833 ();
 sg13g2_decap_8 FILLER_55_840 ();
 sg13g2_decap_8 FILLER_55_847 ();
 sg13g2_decap_8 FILLER_55_854 ();
 sg13g2_fill_1 FILLER_55_861 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_7 ();
 sg13g2_fill_2 FILLER_56_66 ();
 sg13g2_fill_2 FILLER_56_81 ();
 sg13g2_decap_4 FILLER_56_98 ();
 sg13g2_fill_1 FILLER_56_102 ();
 sg13g2_fill_2 FILLER_56_177 ();
 sg13g2_decap_4 FILLER_56_188 ();
 sg13g2_fill_2 FILLER_56_205 ();
 sg13g2_fill_1 FILLER_56_207 ();
 sg13g2_fill_2 FILLER_56_218 ();
 sg13g2_fill_1 FILLER_56_237 ();
 sg13g2_fill_2 FILLER_56_252 ();
 sg13g2_fill_1 FILLER_56_254 ();
 sg13g2_fill_2 FILLER_56_278 ();
 sg13g2_fill_1 FILLER_56_280 ();
 sg13g2_decap_4 FILLER_56_290 ();
 sg13g2_fill_1 FILLER_56_309 ();
 sg13g2_fill_2 FILLER_56_339 ();
 sg13g2_fill_2 FILLER_56_378 ();
 sg13g2_decap_8 FILLER_56_405 ();
 sg13g2_fill_1 FILLER_56_412 ();
 sg13g2_fill_1 FILLER_56_450 ();
 sg13g2_decap_8 FILLER_56_468 ();
 sg13g2_decap_4 FILLER_56_475 ();
 sg13g2_fill_2 FILLER_56_479 ();
 sg13g2_decap_8 FILLER_56_503 ();
 sg13g2_fill_2 FILLER_56_510 ();
 sg13g2_fill_1 FILLER_56_512 ();
 sg13g2_fill_1 FILLER_56_526 ();
 sg13g2_fill_2 FILLER_56_545 ();
 sg13g2_decap_4 FILLER_56_566 ();
 sg13g2_fill_2 FILLER_56_592 ();
 sg13g2_fill_2 FILLER_56_613 ();
 sg13g2_fill_1 FILLER_56_615 ();
 sg13g2_fill_1 FILLER_56_633 ();
 sg13g2_decap_8 FILLER_56_675 ();
 sg13g2_fill_2 FILLER_56_682 ();
 sg13g2_fill_1 FILLER_56_684 ();
 sg13g2_fill_2 FILLER_56_712 ();
 sg13g2_fill_1 FILLER_56_714 ();
 sg13g2_fill_1 FILLER_56_723 ();
 sg13g2_fill_1 FILLER_56_766 ();
 sg13g2_decap_4 FILLER_56_789 ();
 sg13g2_decap_8 FILLER_56_833 ();
 sg13g2_decap_8 FILLER_56_840 ();
 sg13g2_decap_8 FILLER_56_847 ();
 sg13g2_decap_8 FILLER_56_854 ();
 sg13g2_fill_1 FILLER_56_861 ();
 sg13g2_fill_2 FILLER_57_54 ();
 sg13g2_decap_4 FILLER_57_84 ();
 sg13g2_fill_1 FILLER_57_88 ();
 sg13g2_fill_2 FILLER_57_125 ();
 sg13g2_fill_1 FILLER_57_127 ();
 sg13g2_fill_2 FILLER_57_137 ();
 sg13g2_fill_1 FILLER_57_139 ();
 sg13g2_decap_8 FILLER_57_153 ();
 sg13g2_fill_2 FILLER_57_160 ();
 sg13g2_decap_8 FILLER_57_166 ();
 sg13g2_fill_2 FILLER_57_200 ();
 sg13g2_fill_1 FILLER_57_202 ();
 sg13g2_decap_4 FILLER_57_219 ();
 sg13g2_fill_2 FILLER_57_223 ();
 sg13g2_fill_2 FILLER_57_322 ();
 sg13g2_decap_4 FILLER_57_334 ();
 sg13g2_decap_8 FILLER_57_346 ();
 sg13g2_decap_8 FILLER_57_353 ();
 sg13g2_fill_2 FILLER_57_360 ();
 sg13g2_decap_8 FILLER_57_369 ();
 sg13g2_decap_8 FILLER_57_376 ();
 sg13g2_decap_8 FILLER_57_410 ();
 sg13g2_decap_4 FILLER_57_417 ();
 sg13g2_fill_1 FILLER_57_421 ();
 sg13g2_fill_2 FILLER_57_425 ();
 sg13g2_fill_2 FILLER_57_433 ();
 sg13g2_fill_1 FILLER_57_435 ();
 sg13g2_fill_1 FILLER_57_455 ();
 sg13g2_decap_8 FILLER_57_492 ();
 sg13g2_decap_8 FILLER_57_499 ();
 sg13g2_decap_4 FILLER_57_506 ();
 sg13g2_fill_1 FILLER_57_510 ();
 sg13g2_decap_8 FILLER_57_523 ();
 sg13g2_fill_2 FILLER_57_530 ();
 sg13g2_fill_1 FILLER_57_532 ();
 sg13g2_fill_2 FILLER_57_549 ();
 sg13g2_decap_8 FILLER_57_574 ();
 sg13g2_decap_4 FILLER_57_581 ();
 sg13g2_fill_2 FILLER_57_585 ();
 sg13g2_fill_2 FILLER_57_596 ();
 sg13g2_fill_1 FILLER_57_602 ();
 sg13g2_decap_8 FILLER_57_608 ();
 sg13g2_decap_8 FILLER_57_615 ();
 sg13g2_fill_2 FILLER_57_639 ();
 sg13g2_decap_8 FILLER_57_655 ();
 sg13g2_decap_4 FILLER_57_662 ();
 sg13g2_fill_2 FILLER_57_666 ();
 sg13g2_decap_8 FILLER_57_689 ();
 sg13g2_decap_4 FILLER_57_696 ();
 sg13g2_fill_1 FILLER_57_700 ();
 sg13g2_decap_8 FILLER_57_720 ();
 sg13g2_fill_2 FILLER_57_727 ();
 sg13g2_fill_1 FILLER_57_729 ();
 sg13g2_fill_1 FILLER_57_735 ();
 sg13g2_fill_1 FILLER_57_776 ();
 sg13g2_fill_1 FILLER_57_813 ();
 sg13g2_decap_8 FILLER_57_840 ();
 sg13g2_decap_8 FILLER_57_847 ();
 sg13g2_decap_8 FILLER_57_854 ();
 sg13g2_fill_1 FILLER_57_861 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_7 ();
 sg13g2_fill_1 FILLER_58_9 ();
 sg13g2_fill_1 FILLER_58_55 ();
 sg13g2_fill_1 FILLER_58_64 ();
 sg13g2_decap_4 FILLER_58_94 ();
 sg13g2_fill_1 FILLER_58_118 ();
 sg13g2_fill_1 FILLER_58_123 ();
 sg13g2_fill_2 FILLER_58_137 ();
 sg13g2_decap_8 FILLER_58_151 ();
 sg13g2_fill_2 FILLER_58_158 ();
 sg13g2_fill_1 FILLER_58_160 ();
 sg13g2_fill_2 FILLER_58_187 ();
 sg13g2_fill_2 FILLER_58_203 ();
 sg13g2_fill_2 FILLER_58_215 ();
 sg13g2_fill_1 FILLER_58_217 ();
 sg13g2_decap_4 FILLER_58_221 ();
 sg13g2_fill_2 FILLER_58_225 ();
 sg13g2_fill_2 FILLER_58_232 ();
 sg13g2_fill_1 FILLER_58_262 ();
 sg13g2_fill_1 FILLER_58_273 ();
 sg13g2_decap_4 FILLER_58_292 ();
 sg13g2_fill_2 FILLER_58_296 ();
 sg13g2_decap_8 FILLER_58_302 ();
 sg13g2_decap_4 FILLER_58_313 ();
 sg13g2_fill_1 FILLER_58_328 ();
 sg13g2_decap_8 FILLER_58_341 ();
 sg13g2_fill_2 FILLER_58_348 ();
 sg13g2_decap_4 FILLER_58_376 ();
 sg13g2_fill_2 FILLER_58_380 ();
 sg13g2_fill_2 FILLER_58_392 ();
 sg13g2_fill_2 FILLER_58_430 ();
 sg13g2_fill_1 FILLER_58_432 ();
 sg13g2_decap_4 FILLER_58_457 ();
 sg13g2_fill_2 FILLER_58_461 ();
 sg13g2_fill_2 FILLER_58_470 ();
 sg13g2_fill_2 FILLER_58_476 ();
 sg13g2_fill_1 FILLER_58_478 ();
 sg13g2_decap_4 FILLER_58_488 ();
 sg13g2_fill_2 FILLER_58_514 ();
 sg13g2_decap_4 FILLER_58_520 ();
 sg13g2_fill_2 FILLER_58_524 ();
 sg13g2_fill_1 FILLER_58_531 ();
 sg13g2_decap_8 FILLER_58_537 ();
 sg13g2_decap_4 FILLER_58_544 ();
 sg13g2_fill_2 FILLER_58_548 ();
 sg13g2_fill_1 FILLER_58_559 ();
 sg13g2_fill_2 FILLER_58_565 ();
 sg13g2_fill_2 FILLER_58_580 ();
 sg13g2_fill_1 FILLER_58_582 ();
 sg13g2_fill_2 FILLER_58_587 ();
 sg13g2_fill_2 FILLER_58_615 ();
 sg13g2_fill_2 FILLER_58_651 ();
 sg13g2_fill_2 FILLER_58_697 ();
 sg13g2_fill_1 FILLER_58_699 ();
 sg13g2_decap_8 FILLER_58_710 ();
 sg13g2_fill_2 FILLER_58_717 ();
 sg13g2_fill_2 FILLER_58_739 ();
 sg13g2_decap_8 FILLER_58_835 ();
 sg13g2_decap_8 FILLER_58_842 ();
 sg13g2_decap_8 FILLER_58_849 ();
 sg13g2_decap_4 FILLER_58_856 ();
 sg13g2_fill_2 FILLER_58_860 ();
 sg13g2_fill_1 FILLER_59_44 ();
 sg13g2_decap_4 FILLER_59_61 ();
 sg13g2_fill_1 FILLER_59_65 ();
 sg13g2_fill_1 FILLER_59_85 ();
 sg13g2_fill_2 FILLER_59_96 ();
 sg13g2_fill_2 FILLER_59_116 ();
 sg13g2_decap_8 FILLER_59_124 ();
 sg13g2_fill_1 FILLER_59_131 ();
 sg13g2_decap_4 FILLER_59_151 ();
 sg13g2_fill_2 FILLER_59_161 ();
 sg13g2_decap_4 FILLER_59_202 ();
 sg13g2_fill_1 FILLER_59_241 ();
 sg13g2_decap_4 FILLER_59_324 ();
 sg13g2_decap_4 FILLER_59_375 ();
 sg13g2_fill_2 FILLER_59_379 ();
 sg13g2_fill_1 FILLER_59_389 ();
 sg13g2_fill_1 FILLER_59_395 ();
 sg13g2_decap_8 FILLER_59_400 ();
 sg13g2_fill_1 FILLER_59_407 ();
 sg13g2_fill_1 FILLER_59_413 ();
 sg13g2_fill_1 FILLER_59_480 ();
 sg13g2_fill_1 FILLER_59_495 ();
 sg13g2_fill_2 FILLER_59_525 ();
 sg13g2_fill_2 FILLER_59_566 ();
 sg13g2_decap_8 FILLER_59_573 ();
 sg13g2_decap_8 FILLER_59_580 ();
 sg13g2_fill_2 FILLER_59_597 ();
 sg13g2_decap_8 FILLER_59_608 ();
 sg13g2_fill_2 FILLER_59_615 ();
 sg13g2_fill_2 FILLER_59_637 ();
 sg13g2_fill_1 FILLER_59_639 ();
 sg13g2_fill_1 FILLER_59_645 ();
 sg13g2_fill_2 FILLER_59_655 ();
 sg13g2_fill_1 FILLER_59_657 ();
 sg13g2_decap_4 FILLER_59_662 ();
 sg13g2_fill_1 FILLER_59_666 ();
 sg13g2_decap_8 FILLER_59_686 ();
 sg13g2_fill_2 FILLER_59_693 ();
 sg13g2_fill_1 FILLER_59_721 ();
 sg13g2_fill_2 FILLER_59_749 ();
 sg13g2_fill_1 FILLER_59_756 ();
 sg13g2_fill_2 FILLER_59_766 ();
 sg13g2_fill_1 FILLER_59_801 ();
 sg13g2_decap_8 FILLER_59_840 ();
 sg13g2_decap_8 FILLER_59_847 ();
 sg13g2_decap_8 FILLER_59_854 ();
 sg13g2_fill_1 FILLER_59_861 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_7 ();
 sg13g2_fill_1 FILLER_60_9 ();
 sg13g2_fill_1 FILLER_60_41 ();
 sg13g2_decap_8 FILLER_60_61 ();
 sg13g2_fill_1 FILLER_60_68 ();
 sg13g2_fill_2 FILLER_60_78 ();
 sg13g2_fill_2 FILLER_60_84 ();
 sg13g2_fill_1 FILLER_60_86 ();
 sg13g2_decap_4 FILLER_60_92 ();
 sg13g2_decap_4 FILLER_60_118 ();
 sg13g2_decap_8 FILLER_60_127 ();
 sg13g2_fill_1 FILLER_60_134 ();
 sg13g2_decap_8 FILLER_60_150 ();
 sg13g2_decap_4 FILLER_60_157 ();
 sg13g2_fill_2 FILLER_60_175 ();
 sg13g2_fill_1 FILLER_60_177 ();
 sg13g2_decap_4 FILLER_60_225 ();
 sg13g2_fill_1 FILLER_60_247 ();
 sg13g2_decap_4 FILLER_60_280 ();
 sg13g2_fill_2 FILLER_60_284 ();
 sg13g2_fill_2 FILLER_60_357 ();
 sg13g2_fill_1 FILLER_60_359 ();
 sg13g2_fill_2 FILLER_60_393 ();
 sg13g2_decap_4 FILLER_60_417 ();
 sg13g2_decap_4 FILLER_60_425 ();
 sg13g2_fill_2 FILLER_60_429 ();
 sg13g2_decap_4 FILLER_60_437 ();
 sg13g2_fill_1 FILLER_60_441 ();
 sg13g2_decap_8 FILLER_60_447 ();
 sg13g2_decap_4 FILLER_60_458 ();
 sg13g2_fill_1 FILLER_60_462 ();
 sg13g2_fill_2 FILLER_60_469 ();
 sg13g2_fill_1 FILLER_60_471 ();
 sg13g2_fill_1 FILLER_60_484 ();
 sg13g2_fill_1 FILLER_60_493 ();
 sg13g2_decap_4 FILLER_60_503 ();
 sg13g2_fill_1 FILLER_60_512 ();
 sg13g2_decap_8 FILLER_60_517 ();
 sg13g2_decap_4 FILLER_60_530 ();
 sg13g2_fill_2 FILLER_60_534 ();
 sg13g2_decap_4 FILLER_60_540 ();
 sg13g2_fill_1 FILLER_60_544 ();
 sg13g2_fill_1 FILLER_60_552 ();
 sg13g2_decap_8 FILLER_60_568 ();
 sg13g2_fill_2 FILLER_60_575 ();
 sg13g2_decap_4 FILLER_60_582 ();
 sg13g2_decap_8 FILLER_60_614 ();
 sg13g2_fill_1 FILLER_60_621 ();
 sg13g2_fill_1 FILLER_60_648 ();
 sg13g2_fill_2 FILLER_60_662 ();
 sg13g2_fill_2 FILLER_60_683 ();
 sg13g2_fill_1 FILLER_60_695 ();
 sg13g2_decap_4 FILLER_60_704 ();
 sg13g2_fill_1 FILLER_60_708 ();
 sg13g2_decap_4 FILLER_60_717 ();
 sg13g2_fill_2 FILLER_60_721 ();
 sg13g2_fill_2 FILLER_60_737 ();
 sg13g2_fill_2 FILLER_60_752 ();
 sg13g2_fill_1 FILLER_60_754 ();
 sg13g2_fill_2 FILLER_60_768 ();
 sg13g2_fill_1 FILLER_60_770 ();
 sg13g2_decap_4 FILLER_60_778 ();
 sg13g2_fill_2 FILLER_60_782 ();
 sg13g2_decap_8 FILLER_60_846 ();
 sg13g2_decap_8 FILLER_60_853 ();
 sg13g2_fill_2 FILLER_60_860 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_7 ();
 sg13g2_fill_2 FILLER_61_63 ();
 sg13g2_fill_1 FILLER_61_65 ();
 sg13g2_fill_2 FILLER_61_81 ();
 sg13g2_fill_1 FILLER_61_88 ();
 sg13g2_decap_8 FILLER_61_93 ();
 sg13g2_fill_2 FILLER_61_100 ();
 sg13g2_fill_2 FILLER_61_116 ();
 sg13g2_fill_1 FILLER_61_118 ();
 sg13g2_decap_8 FILLER_61_124 ();
 sg13g2_decap_4 FILLER_61_131 ();
 sg13g2_decap_8 FILLER_61_161 ();
 sg13g2_fill_1 FILLER_61_168 ();
 sg13g2_fill_2 FILLER_61_179 ();
 sg13g2_fill_1 FILLER_61_181 ();
 sg13g2_fill_1 FILLER_61_213 ();
 sg13g2_decap_4 FILLER_61_224 ();
 sg13g2_fill_2 FILLER_61_251 ();
 sg13g2_decap_4 FILLER_61_278 ();
 sg13g2_fill_1 FILLER_61_282 ();
 sg13g2_decap_4 FILLER_61_343 ();
 sg13g2_decap_4 FILLER_61_353 ();
 sg13g2_fill_2 FILLER_61_378 ();
 sg13g2_decap_4 FILLER_61_405 ();
 sg13g2_fill_1 FILLER_61_433 ();
 sg13g2_fill_2 FILLER_61_456 ();
 sg13g2_fill_1 FILLER_61_458 ();
 sg13g2_fill_1 FILLER_61_464 ();
 sg13g2_decap_8 FILLER_61_478 ();
 sg13g2_fill_1 FILLER_61_485 ();
 sg13g2_decap_4 FILLER_61_492 ();
 sg13g2_fill_2 FILLER_61_496 ();
 sg13g2_fill_1 FILLER_61_541 ();
 sg13g2_fill_2 FILLER_61_560 ();
 sg13g2_fill_1 FILLER_61_562 ();
 sg13g2_decap_4 FILLER_61_585 ();
 sg13g2_decap_8 FILLER_61_604 ();
 sg13g2_decap_4 FILLER_61_611 ();
 sg13g2_fill_1 FILLER_61_639 ();
 sg13g2_fill_2 FILLER_61_645 ();
 sg13g2_decap_4 FILLER_61_660 ();
 sg13g2_fill_2 FILLER_61_664 ();
 sg13g2_fill_1 FILLER_61_671 ();
 sg13g2_decap_8 FILLER_61_689 ();
 sg13g2_decap_4 FILLER_61_696 ();
 sg13g2_decap_8 FILLER_61_704 ();
 sg13g2_decap_4 FILLER_61_711 ();
 sg13g2_decap_4 FILLER_61_739 ();
 sg13g2_fill_2 FILLER_61_743 ();
 sg13g2_fill_2 FILLER_61_765 ();
 sg13g2_fill_1 FILLER_61_767 ();
 sg13g2_fill_2 FILLER_61_772 ();
 sg13g2_fill_1 FILLER_61_774 ();
 sg13g2_decap_4 FILLER_61_787 ();
 sg13g2_fill_2 FILLER_61_791 ();
 sg13g2_fill_1 FILLER_61_798 ();
 sg13g2_fill_2 FILLER_61_809 ();
 sg13g2_fill_1 FILLER_61_811 ();
 sg13g2_decap_8 FILLER_61_842 ();
 sg13g2_decap_8 FILLER_61_849 ();
 sg13g2_decap_4 FILLER_61_856 ();
 sg13g2_fill_2 FILLER_61_860 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_4 FILLER_62_14 ();
 sg13g2_fill_1 FILLER_62_18 ();
 sg13g2_decap_4 FILLER_62_23 ();
 sg13g2_fill_1 FILLER_62_31 ();
 sg13g2_decap_4 FILLER_62_36 ();
 sg13g2_fill_2 FILLER_62_40 ();
 sg13g2_fill_2 FILLER_62_46 ();
 sg13g2_fill_1 FILLER_62_48 ();
 sg13g2_fill_2 FILLER_62_61 ();
 sg13g2_fill_1 FILLER_62_63 ();
 sg13g2_fill_1 FILLER_62_74 ();
 sg13g2_fill_2 FILLER_62_94 ();
 sg13g2_fill_1 FILLER_62_96 ();
 sg13g2_fill_1 FILLER_62_107 ();
 sg13g2_fill_2 FILLER_62_117 ();
 sg13g2_decap_8 FILLER_62_129 ();
 sg13g2_decap_4 FILLER_62_136 ();
 sg13g2_decap_4 FILLER_62_159 ();
 sg13g2_fill_2 FILLER_62_163 ();
 sg13g2_fill_2 FILLER_62_191 ();
 sg13g2_fill_1 FILLER_62_193 ();
 sg13g2_fill_1 FILLER_62_200 ();
 sg13g2_fill_2 FILLER_62_224 ();
 sg13g2_fill_1 FILLER_62_226 ();
 sg13g2_fill_2 FILLER_62_248 ();
 sg13g2_fill_1 FILLER_62_250 ();
 sg13g2_fill_2 FILLER_62_259 ();
 sg13g2_fill_1 FILLER_62_266 ();
 sg13g2_fill_2 FILLER_62_280 ();
 sg13g2_fill_1 FILLER_62_282 ();
 sg13g2_fill_2 FILLER_62_320 ();
 sg13g2_decap_8 FILLER_62_348 ();
 sg13g2_decap_8 FILLER_62_355 ();
 sg13g2_decap_8 FILLER_62_374 ();
 sg13g2_decap_4 FILLER_62_381 ();
 sg13g2_fill_1 FILLER_62_385 ();
 sg13g2_decap_4 FILLER_62_398 ();
 sg13g2_fill_1 FILLER_62_402 ();
 sg13g2_fill_2 FILLER_62_429 ();
 sg13g2_fill_1 FILLER_62_431 ();
 sg13g2_decap_8 FILLER_62_464 ();
 sg13g2_decap_4 FILLER_62_498 ();
 sg13g2_fill_2 FILLER_62_502 ();
 sg13g2_decap_8 FILLER_62_510 ();
 sg13g2_fill_2 FILLER_62_517 ();
 sg13g2_fill_1 FILLER_62_519 ();
 sg13g2_fill_2 FILLER_62_525 ();
 sg13g2_decap_4 FILLER_62_536 ();
 sg13g2_decap_4 FILLER_62_564 ();
 sg13g2_fill_1 FILLER_62_568 ();
 sg13g2_decap_8 FILLER_62_574 ();
 sg13g2_decap_4 FILLER_62_581 ();
 sg13g2_decap_8 FILLER_62_608 ();
 sg13g2_decap_8 FILLER_62_615 ();
 sg13g2_fill_2 FILLER_62_622 ();
 sg13g2_fill_2 FILLER_62_632 ();
 sg13g2_fill_1 FILLER_62_634 ();
 sg13g2_decap_8 FILLER_62_646 ();
 sg13g2_decap_4 FILLER_62_662 ();
 sg13g2_decap_4 FILLER_62_670 ();
 sg13g2_fill_1 FILLER_62_674 ();
 sg13g2_decap_4 FILLER_62_721 ();
 sg13g2_fill_2 FILLER_62_733 ();
 sg13g2_fill_1 FILLER_62_735 ();
 sg13g2_decap_4 FILLER_62_758 ();
 sg13g2_fill_1 FILLER_62_762 ();
 sg13g2_decap_8 FILLER_62_833 ();
 sg13g2_decap_8 FILLER_62_840 ();
 sg13g2_decap_8 FILLER_62_847 ();
 sg13g2_decap_8 FILLER_62_854 ();
 sg13g2_fill_1 FILLER_62_861 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_4 FILLER_63_7 ();
 sg13g2_fill_1 FILLER_63_11 ();
 sg13g2_fill_1 FILLER_63_69 ();
 sg13g2_fill_2 FILLER_63_75 ();
 sg13g2_fill_2 FILLER_63_88 ();
 sg13g2_decap_8 FILLER_63_94 ();
 sg13g2_fill_1 FILLER_63_101 ();
 sg13g2_fill_2 FILLER_63_132 ();
 sg13g2_fill_1 FILLER_63_134 ();
 sg13g2_fill_1 FILLER_63_150 ();
 sg13g2_fill_2 FILLER_63_180 ();
 sg13g2_fill_1 FILLER_63_200 ();
 sg13g2_decap_8 FILLER_63_221 ();
 sg13g2_decap_4 FILLER_63_228 ();
 sg13g2_decap_4 FILLER_63_240 ();
 sg13g2_decap_8 FILLER_63_253 ();
 sg13g2_fill_2 FILLER_63_260 ();
 sg13g2_fill_1 FILLER_63_262 ();
 sg13g2_decap_8 FILLER_63_284 ();
 sg13g2_fill_2 FILLER_63_291 ();
 sg13g2_fill_2 FILLER_63_336 ();
 sg13g2_fill_2 FILLER_63_349 ();
 sg13g2_fill_1 FILLER_63_351 ();
 sg13g2_fill_2 FILLER_63_367 ();
 sg13g2_fill_1 FILLER_63_369 ();
 sg13g2_decap_8 FILLER_63_383 ();
 sg13g2_decap_4 FILLER_63_402 ();
 sg13g2_fill_2 FILLER_63_424 ();
 sg13g2_decap_8 FILLER_63_435 ();
 sg13g2_decap_8 FILLER_63_442 ();
 sg13g2_fill_1 FILLER_63_449 ();
 sg13g2_fill_2 FILLER_63_480 ();
 sg13g2_fill_2 FILLER_63_487 ();
 sg13g2_decap_4 FILLER_63_503 ();
 sg13g2_fill_2 FILLER_63_507 ();
 sg13g2_decap_4 FILLER_63_524 ();
 sg13g2_fill_1 FILLER_63_539 ();
 sg13g2_fill_1 FILLER_63_570 ();
 sg13g2_decap_4 FILLER_63_575 ();
 sg13g2_decap_4 FILLER_63_591 ();
 sg13g2_fill_2 FILLER_63_595 ();
 sg13g2_fill_1 FILLER_63_608 ();
 sg13g2_fill_2 FILLER_63_628 ();
 sg13g2_fill_2 FILLER_63_647 ();
 sg13g2_decap_4 FILLER_63_668 ();
 sg13g2_fill_1 FILLER_63_672 ();
 sg13g2_decap_8 FILLER_63_682 ();
 sg13g2_fill_2 FILLER_63_689 ();
 sg13g2_fill_1 FILLER_63_691 ();
 sg13g2_fill_2 FILLER_63_716 ();
 sg13g2_fill_2 FILLER_63_737 ();
 sg13g2_decap_4 FILLER_63_769 ();
 sg13g2_fill_2 FILLER_63_773 ();
 sg13g2_fill_1 FILLER_63_780 ();
 sg13g2_decap_8 FILLER_63_791 ();
 sg13g2_fill_2 FILLER_63_817 ();
 sg13g2_decap_8 FILLER_63_836 ();
 sg13g2_decap_8 FILLER_63_843 ();
 sg13g2_decap_8 FILLER_63_850 ();
 sg13g2_decap_4 FILLER_63_857 ();
 sg13g2_fill_1 FILLER_63_861 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_28 ();
 sg13g2_fill_2 FILLER_64_74 ();
 sg13g2_fill_2 FILLER_64_85 ();
 sg13g2_fill_1 FILLER_64_96 ();
 sg13g2_fill_1 FILLER_64_135 ();
 sg13g2_fill_2 FILLER_64_147 ();
 sg13g2_fill_2 FILLER_64_154 ();
 sg13g2_decap_8 FILLER_64_160 ();
 sg13g2_fill_2 FILLER_64_167 ();
 sg13g2_fill_2 FILLER_64_173 ();
 sg13g2_fill_1 FILLER_64_175 ();
 sg13g2_decap_4 FILLER_64_180 ();
 sg13g2_fill_2 FILLER_64_184 ();
 sg13g2_fill_1 FILLER_64_212 ();
 sg13g2_decap_4 FILLER_64_223 ();
 sg13g2_fill_2 FILLER_64_227 ();
 sg13g2_decap_8 FILLER_64_258 ();
 sg13g2_fill_2 FILLER_64_265 ();
 sg13g2_fill_1 FILLER_64_267 ();
 sg13g2_fill_2 FILLER_64_274 ();
 sg13g2_fill_2 FILLER_64_320 ();
 sg13g2_fill_2 FILLER_64_362 ();
 sg13g2_fill_1 FILLER_64_364 ();
 sg13g2_fill_1 FILLER_64_370 ();
 sg13g2_decap_4 FILLER_64_383 ();
 sg13g2_decap_8 FILLER_64_392 ();
 sg13g2_decap_8 FILLER_64_399 ();
 sg13g2_fill_1 FILLER_64_406 ();
 sg13g2_fill_2 FILLER_64_412 ();
 sg13g2_decap_4 FILLER_64_419 ();
 sg13g2_fill_1 FILLER_64_423 ();
 sg13g2_decap_8 FILLER_64_445 ();
 sg13g2_fill_2 FILLER_64_452 ();
 sg13g2_fill_1 FILLER_64_461 ();
 sg13g2_fill_2 FILLER_64_466 ();
 sg13g2_fill_2 FILLER_64_491 ();
 sg13g2_fill_2 FILLER_64_503 ();
 sg13g2_fill_2 FILLER_64_527 ();
 sg13g2_fill_1 FILLER_64_529 ();
 sg13g2_decap_4 FILLER_64_535 ();
 sg13g2_fill_1 FILLER_64_539 ();
 sg13g2_decap_8 FILLER_64_560 ();
 sg13g2_fill_2 FILLER_64_567 ();
 sg13g2_fill_1 FILLER_64_569 ();
 sg13g2_fill_2 FILLER_64_579 ();
 sg13g2_fill_2 FILLER_64_587 ();
 sg13g2_fill_1 FILLER_64_589 ();
 sg13g2_decap_4 FILLER_64_605 ();
 sg13g2_fill_2 FILLER_64_609 ();
 sg13g2_decap_8 FILLER_64_632 ();
 sg13g2_decap_8 FILLER_64_644 ();
 sg13g2_fill_1 FILLER_64_655 ();
 sg13g2_fill_2 FILLER_64_661 ();
 sg13g2_fill_2 FILLER_64_678 ();
 sg13g2_fill_1 FILLER_64_680 ();
 sg13g2_fill_1 FILLER_64_701 ();
 sg13g2_decap_8 FILLER_64_710 ();
 sg13g2_decap_4 FILLER_64_717 ();
 sg13g2_fill_1 FILLER_64_721 ();
 sg13g2_fill_2 FILLER_64_732 ();
 sg13g2_fill_1 FILLER_64_734 ();
 sg13g2_fill_1 FILLER_64_743 ();
 sg13g2_decap_8 FILLER_64_760 ();
 sg13g2_decap_4 FILLER_64_767 ();
 sg13g2_fill_2 FILLER_64_771 ();
 sg13g2_fill_2 FILLER_64_781 ();
 sg13g2_fill_1 FILLER_64_783 ();
 sg13g2_decap_8 FILLER_64_838 ();
 sg13g2_decap_8 FILLER_64_845 ();
 sg13g2_decap_8 FILLER_64_852 ();
 sg13g2_fill_2 FILLER_64_859 ();
 sg13g2_fill_1 FILLER_64_861 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_fill_2 FILLER_65_7 ();
 sg13g2_fill_1 FILLER_65_9 ();
 sg13g2_fill_1 FILLER_65_22 ();
 sg13g2_fill_1 FILLER_65_36 ();
 sg13g2_fill_1 FILLER_65_42 ();
 sg13g2_fill_2 FILLER_65_56 ();
 sg13g2_fill_1 FILLER_65_76 ();
 sg13g2_fill_1 FILLER_65_109 ();
 sg13g2_fill_2 FILLER_65_123 ();
 sg13g2_fill_2 FILLER_65_156 ();
 sg13g2_fill_2 FILLER_65_193 ();
 sg13g2_fill_2 FILLER_65_218 ();
 sg13g2_fill_1 FILLER_65_220 ();
 sg13g2_decap_8 FILLER_65_231 ();
 sg13g2_fill_2 FILLER_65_238 ();
 sg13g2_fill_1 FILLER_65_240 ();
 sg13g2_fill_2 FILLER_65_246 ();
 sg13g2_fill_1 FILLER_65_248 ();
 sg13g2_fill_2 FILLER_65_264 ();
 sg13g2_decap_4 FILLER_65_286 ();
 sg13g2_fill_2 FILLER_65_311 ();
 sg13g2_fill_1 FILLER_65_313 ();
 sg13g2_fill_2 FILLER_65_331 ();
 sg13g2_decap_4 FILLER_65_350 ();
 sg13g2_fill_2 FILLER_65_411 ();
 sg13g2_fill_1 FILLER_65_413 ();
 sg13g2_fill_1 FILLER_65_432 ();
 sg13g2_decap_4 FILLER_65_459 ();
 sg13g2_fill_2 FILLER_65_477 ();
 sg13g2_fill_2 FILLER_65_484 ();
 sg13g2_fill_1 FILLER_65_495 ();
 sg13g2_fill_2 FILLER_65_511 ();
 sg13g2_fill_1 FILLER_65_513 ();
 sg13g2_fill_2 FILLER_65_530 ();
 sg13g2_fill_1 FILLER_65_532 ();
 sg13g2_fill_1 FILLER_65_549 ();
 sg13g2_fill_2 FILLER_65_555 ();
 sg13g2_decap_8 FILLER_65_567 ();
 sg13g2_fill_2 FILLER_65_574 ();
 sg13g2_decap_4 FILLER_65_582 ();
 sg13g2_fill_1 FILLER_65_586 ();
 sg13g2_fill_2 FILLER_65_599 ();
 sg13g2_fill_1 FILLER_65_601 ();
 sg13g2_fill_2 FILLER_65_612 ();
 sg13g2_fill_1 FILLER_65_614 ();
 sg13g2_fill_2 FILLER_65_626 ();
 sg13g2_fill_1 FILLER_65_628 ();
 sg13g2_fill_2 FILLER_65_637 ();
 sg13g2_fill_1 FILLER_65_639 ();
 sg13g2_fill_2 FILLER_65_650 ();
 sg13g2_decap_4 FILLER_65_661 ();
 sg13g2_fill_1 FILLER_65_665 ();
 sg13g2_decap_8 FILLER_65_687 ();
 sg13g2_fill_1 FILLER_65_694 ();
 sg13g2_fill_1 FILLER_65_746 ();
 sg13g2_fill_2 FILLER_65_751 ();
 sg13g2_fill_1 FILLER_65_753 ();
 sg13g2_fill_2 FILLER_65_762 ();
 sg13g2_fill_1 FILLER_65_768 ();
 sg13g2_decap_4 FILLER_65_778 ();
 sg13g2_fill_1 FILLER_65_782 ();
 sg13g2_fill_1 FILLER_65_793 ();
 sg13g2_decap_8 FILLER_65_830 ();
 sg13g2_decap_8 FILLER_65_837 ();
 sg13g2_decap_8 FILLER_65_844 ();
 sg13g2_decap_8 FILLER_65_851 ();
 sg13g2_decap_4 FILLER_65_858 ();
 sg13g2_decap_4 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_4 ();
 sg13g2_fill_1 FILLER_66_51 ();
 sg13g2_fill_2 FILLER_66_72 ();
 sg13g2_fill_1 FILLER_66_102 ();
 sg13g2_fill_1 FILLER_66_138 ();
 sg13g2_fill_2 FILLER_66_148 ();
 sg13g2_fill_1 FILLER_66_150 ();
 sg13g2_fill_1 FILLER_66_182 ();
 sg13g2_fill_1 FILLER_66_223 ();
 sg13g2_fill_2 FILLER_66_253 ();
 sg13g2_fill_1 FILLER_66_255 ();
 sg13g2_fill_1 FILLER_66_264 ();
 sg13g2_decap_4 FILLER_66_285 ();
 sg13g2_fill_1 FILLER_66_289 ();
 sg13g2_fill_1 FILLER_66_310 ();
 sg13g2_fill_2 FILLER_66_347 ();
 sg13g2_fill_2 FILLER_66_354 ();
 sg13g2_decap_8 FILLER_66_361 ();
 sg13g2_decap_4 FILLER_66_368 ();
 sg13g2_decap_8 FILLER_66_381 ();
 sg13g2_decap_4 FILLER_66_388 ();
 sg13g2_fill_1 FILLER_66_392 ();
 sg13g2_fill_2 FILLER_66_405 ();
 sg13g2_fill_2 FILLER_66_414 ();
 sg13g2_fill_1 FILLER_66_430 ();
 sg13g2_fill_1 FILLER_66_435 ();
 sg13g2_fill_1 FILLER_66_452 ();
 sg13g2_fill_1 FILLER_66_468 ();
 sg13g2_decap_4 FILLER_66_486 ();
 sg13g2_fill_2 FILLER_66_490 ();
 sg13g2_fill_1 FILLER_66_512 ();
 sg13g2_fill_2 FILLER_66_539 ();
 sg13g2_decap_4 FILLER_66_553 ();
 sg13g2_decap_4 FILLER_66_564 ();
 sg13g2_decap_4 FILLER_66_580 ();
 sg13g2_fill_2 FILLER_66_598 ();
 sg13g2_fill_1 FILLER_66_606 ();
 sg13g2_fill_2 FILLER_66_623 ();
 sg13g2_fill_1 FILLER_66_625 ();
 sg13g2_decap_8 FILLER_66_631 ();
 sg13g2_decap_4 FILLER_66_645 ();
 sg13g2_fill_1 FILLER_66_653 ();
 sg13g2_fill_2 FILLER_66_659 ();
 sg13g2_fill_2 FILLER_66_664 ();
 sg13g2_fill_2 FILLER_66_674 ();
 sg13g2_fill_1 FILLER_66_710 ();
 sg13g2_decap_8 FILLER_66_737 ();
 sg13g2_fill_2 FILLER_66_787 ();
 sg13g2_decap_8 FILLER_66_828 ();
 sg13g2_decap_8 FILLER_66_835 ();
 sg13g2_decap_8 FILLER_66_842 ();
 sg13g2_decap_8 FILLER_66_849 ();
 sg13g2_decap_4 FILLER_66_856 ();
 sg13g2_fill_2 FILLER_66_860 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_7 ();
 sg13g2_fill_1 FILLER_67_34 ();
 sg13g2_fill_1 FILLER_67_96 ();
 sg13g2_fill_1 FILLER_67_133 ();
 sg13g2_fill_2 FILLER_67_165 ();
 sg13g2_fill_2 FILLER_67_171 ();
 sg13g2_fill_1 FILLER_67_181 ();
 sg13g2_fill_1 FILLER_67_191 ();
 sg13g2_fill_1 FILLER_67_212 ();
 sg13g2_fill_2 FILLER_67_227 ();
 sg13g2_decap_8 FILLER_67_233 ();
 sg13g2_decap_4 FILLER_67_240 ();
 sg13g2_fill_2 FILLER_67_244 ();
 sg13g2_decap_4 FILLER_67_253 ();
 sg13g2_fill_2 FILLER_67_257 ();
 sg13g2_decap_8 FILLER_67_271 ();
 sg13g2_decap_8 FILLER_67_278 ();
 sg13g2_fill_2 FILLER_67_285 ();
 sg13g2_fill_1 FILLER_67_311 ();
 sg13g2_decap_8 FILLER_67_316 ();
 sg13g2_decap_4 FILLER_67_323 ();
 sg13g2_decap_4 FILLER_67_331 ();
 sg13g2_fill_2 FILLER_67_335 ();
 sg13g2_fill_2 FILLER_67_364 ();
 sg13g2_fill_2 FILLER_67_388 ();
 sg13g2_fill_2 FILLER_67_402 ();
 sg13g2_fill_1 FILLER_67_404 ();
 sg13g2_fill_2 FILLER_67_413 ();
 sg13g2_fill_1 FILLER_67_415 ();
 sg13g2_fill_1 FILLER_67_426 ();
 sg13g2_decap_4 FILLER_67_449 ();
 sg13g2_fill_1 FILLER_67_453 ();
 sg13g2_fill_2 FILLER_67_509 ();
 sg13g2_fill_1 FILLER_67_511 ();
 sg13g2_fill_2 FILLER_67_520 ();
 sg13g2_fill_1 FILLER_67_522 ();
 sg13g2_decap_4 FILLER_67_531 ();
 sg13g2_fill_2 FILLER_67_539 ();
 sg13g2_fill_1 FILLER_67_541 ();
 sg13g2_decap_4 FILLER_67_552 ();
 sg13g2_fill_1 FILLER_67_556 ();
 sg13g2_fill_1 FILLER_67_567 ();
 sg13g2_fill_1 FILLER_67_585 ();
 sg13g2_decap_8 FILLER_67_590 ();
 sg13g2_decap_8 FILLER_67_597 ();
 sg13g2_fill_2 FILLER_67_604 ();
 sg13g2_fill_1 FILLER_67_606 ();
 sg13g2_fill_2 FILLER_67_622 ();
 sg13g2_decap_8 FILLER_67_661 ();
 sg13g2_decap_4 FILLER_67_678 ();
 sg13g2_fill_1 FILLER_67_682 ();
 sg13g2_decap_8 FILLER_67_693 ();
 sg13g2_decap_4 FILLER_67_700 ();
 sg13g2_fill_1 FILLER_67_704 ();
 sg13g2_decap_8 FILLER_67_710 ();
 sg13g2_decap_8 FILLER_67_717 ();
 sg13g2_fill_2 FILLER_67_729 ();
 sg13g2_fill_1 FILLER_67_731 ();
 sg13g2_decap_8 FILLER_67_751 ();
 sg13g2_fill_2 FILLER_67_775 ();
 sg13g2_fill_1 FILLER_67_777 ();
 sg13g2_decap_8 FILLER_67_808 ();
 sg13g2_decap_8 FILLER_67_815 ();
 sg13g2_decap_8 FILLER_67_822 ();
 sg13g2_decap_8 FILLER_67_829 ();
 sg13g2_decap_8 FILLER_67_836 ();
 sg13g2_decap_8 FILLER_67_843 ();
 sg13g2_decap_8 FILLER_67_850 ();
 sg13g2_decap_4 FILLER_67_857 ();
 sg13g2_fill_1 FILLER_67_861 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_2 ();
 sg13g2_fill_1 FILLER_68_29 ();
 sg13g2_fill_2 FILLER_68_91 ();
 sg13g2_fill_1 FILLER_68_102 ();
 sg13g2_fill_2 FILLER_68_127 ();
 sg13g2_decap_8 FILLER_68_151 ();
 sg13g2_fill_2 FILLER_68_158 ();
 sg13g2_fill_1 FILLER_68_160 ();
 sg13g2_fill_2 FILLER_68_219 ();
 sg13g2_fill_1 FILLER_68_221 ();
 sg13g2_fill_2 FILLER_68_238 ();
 sg13g2_decap_8 FILLER_68_264 ();
 sg13g2_decap_8 FILLER_68_271 ();
 sg13g2_fill_1 FILLER_68_278 ();
 sg13g2_decap_4 FILLER_68_286 ();
 sg13g2_fill_1 FILLER_68_290 ();
 sg13g2_fill_1 FILLER_68_312 ();
 sg13g2_decap_8 FILLER_68_330 ();
 sg13g2_fill_2 FILLER_68_337 ();
 sg13g2_fill_1 FILLER_68_339 ();
 sg13g2_decap_4 FILLER_68_364 ();
 sg13g2_fill_2 FILLER_68_380 ();
 sg13g2_decap_4 FILLER_68_398 ();
 sg13g2_fill_2 FILLER_68_402 ();
 sg13g2_decap_8 FILLER_68_420 ();
 sg13g2_fill_1 FILLER_68_427 ();
 sg13g2_fill_2 FILLER_68_443 ();
 sg13g2_decap_4 FILLER_68_453 ();
 sg13g2_fill_2 FILLER_68_457 ();
 sg13g2_fill_1 FILLER_68_465 ();
 sg13g2_fill_2 FILLER_68_475 ();
 sg13g2_fill_2 FILLER_68_486 ();
 sg13g2_fill_1 FILLER_68_488 ();
 sg13g2_decap_4 FILLER_68_515 ();
 sg13g2_fill_2 FILLER_68_523 ();
 sg13g2_fill_1 FILLER_68_565 ();
 sg13g2_fill_1 FILLER_68_570 ();
 sg13g2_decap_4 FILLER_68_576 ();
 sg13g2_fill_2 FILLER_68_595 ();
 sg13g2_fill_1 FILLER_68_597 ();
 sg13g2_fill_2 FILLER_68_632 ();
 sg13g2_fill_2 FILLER_68_652 ();
 sg13g2_decap_4 FILLER_68_668 ();
 sg13g2_fill_1 FILLER_68_672 ();
 sg13g2_fill_2 FILLER_68_678 ();
 sg13g2_fill_2 FILLER_68_689 ();
 sg13g2_fill_1 FILLER_68_691 ();
 sg13g2_fill_1 FILLER_68_735 ();
 sg13g2_fill_2 FILLER_68_771 ();
 sg13g2_fill_1 FILLER_68_773 ();
 sg13g2_fill_2 FILLER_68_793 ();
 sg13g2_fill_1 FILLER_68_795 ();
 sg13g2_decap_8 FILLER_68_805 ();
 sg13g2_decap_8 FILLER_68_812 ();
 sg13g2_decap_8 FILLER_68_819 ();
 sg13g2_decap_8 FILLER_68_826 ();
 sg13g2_decap_8 FILLER_68_833 ();
 sg13g2_decap_8 FILLER_68_840 ();
 sg13g2_decap_8 FILLER_68_847 ();
 sg13g2_decap_8 FILLER_68_854 ();
 sg13g2_fill_1 FILLER_68_861 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_4 FILLER_69_7 ();
 sg13g2_fill_1 FILLER_69_11 ();
 sg13g2_fill_2 FILLER_69_38 ();
 sg13g2_fill_1 FILLER_69_62 ();
 sg13g2_fill_2 FILLER_69_72 ();
 sg13g2_fill_1 FILLER_69_128 ();
 sg13g2_fill_2 FILLER_69_135 ();
 sg13g2_fill_1 FILLER_69_142 ();
 sg13g2_decap_4 FILLER_69_149 ();
 sg13g2_fill_1 FILLER_69_153 ();
 sg13g2_decap_4 FILLER_69_158 ();
 sg13g2_fill_2 FILLER_69_183 ();
 sg13g2_fill_1 FILLER_69_185 ();
 sg13g2_fill_2 FILLER_69_192 ();
 sg13g2_decap_8 FILLER_69_200 ();
 sg13g2_decap_4 FILLER_69_207 ();
 sg13g2_fill_2 FILLER_69_211 ();
 sg13g2_fill_1 FILLER_69_225 ();
 sg13g2_fill_2 FILLER_69_244 ();
 sg13g2_decap_4 FILLER_69_261 ();
 sg13g2_fill_1 FILLER_69_265 ();
 sg13g2_fill_2 FILLER_69_311 ();
 sg13g2_fill_2 FILLER_69_332 ();
 sg13g2_fill_1 FILLER_69_334 ();
 sg13g2_decap_8 FILLER_69_351 ();
 sg13g2_fill_1 FILLER_69_358 ();
 sg13g2_decap_4 FILLER_69_367 ();
 sg13g2_fill_1 FILLER_69_371 ();
 sg13g2_decap_4 FILLER_69_380 ();
 sg13g2_decap_4 FILLER_69_392 ();
 sg13g2_decap_8 FILLER_69_403 ();
 sg13g2_decap_4 FILLER_69_416 ();
 sg13g2_fill_2 FILLER_69_452 ();
 sg13g2_fill_2 FILLER_69_472 ();
 sg13g2_fill_1 FILLER_69_474 ();
 sg13g2_fill_2 FILLER_69_492 ();
 sg13g2_fill_2 FILLER_69_498 ();
 sg13g2_decap_4 FILLER_69_511 ();
 sg13g2_fill_2 FILLER_69_515 ();
 sg13g2_decap_8 FILLER_69_530 ();
 sg13g2_fill_2 FILLER_69_537 ();
 sg13g2_fill_2 FILLER_69_549 ();
 sg13g2_fill_1 FILLER_69_551 ();
 sg13g2_fill_2 FILLER_69_563 ();
 sg13g2_fill_1 FILLER_69_572 ();
 sg13g2_decap_4 FILLER_69_578 ();
 sg13g2_fill_2 FILLER_69_582 ();
 sg13g2_decap_4 FILLER_69_588 ();
 sg13g2_fill_1 FILLER_69_592 ();
 sg13g2_fill_2 FILLER_69_598 ();
 sg13g2_decap_8 FILLER_69_606 ();
 sg13g2_fill_2 FILLER_69_613 ();
 sg13g2_fill_1 FILLER_69_644 ();
 sg13g2_fill_2 FILLER_69_688 ();
 sg13g2_fill_1 FILLER_69_721 ();
 sg13g2_decap_4 FILLER_69_747 ();
 sg13g2_fill_2 FILLER_69_768 ();
 sg13g2_fill_1 FILLER_69_770 ();
 sg13g2_fill_2 FILLER_69_797 ();
 sg13g2_decap_8 FILLER_69_825 ();
 sg13g2_decap_8 FILLER_69_832 ();
 sg13g2_decap_8 FILLER_69_839 ();
 sg13g2_decap_8 FILLER_69_846 ();
 sg13g2_decap_8 FILLER_69_853 ();
 sg13g2_fill_2 FILLER_69_860 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_fill_2 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_20 ();
 sg13g2_decap_4 FILLER_70_27 ();
 sg13g2_fill_2 FILLER_70_40 ();
 sg13g2_fill_1 FILLER_70_42 ();
 sg13g2_fill_2 FILLER_70_47 ();
 sg13g2_decap_8 FILLER_70_57 ();
 sg13g2_decap_8 FILLER_70_64 ();
 sg13g2_decap_8 FILLER_70_71 ();
 sg13g2_fill_2 FILLER_70_78 ();
 sg13g2_fill_1 FILLER_70_80 ();
 sg13g2_fill_1 FILLER_70_105 ();
 sg13g2_fill_2 FILLER_70_126 ();
 sg13g2_fill_2 FILLER_70_137 ();
 sg13g2_fill_1 FILLER_70_139 ();
 sg13g2_fill_2 FILLER_70_151 ();
 sg13g2_fill_2 FILLER_70_168 ();
 sg13g2_fill_1 FILLER_70_170 ();
 sg13g2_fill_1 FILLER_70_202 ();
 sg13g2_fill_2 FILLER_70_209 ();
 sg13g2_fill_1 FILLER_70_237 ();
 sg13g2_fill_2 FILLER_70_244 ();
 sg13g2_fill_1 FILLER_70_246 ();
 sg13g2_fill_2 FILLER_70_264 ();
 sg13g2_fill_1 FILLER_70_295 ();
 sg13g2_fill_1 FILLER_70_319 ();
 sg13g2_fill_2 FILLER_70_379 ();
 sg13g2_fill_1 FILLER_70_381 ();
 sg13g2_fill_2 FILLER_70_386 ();
 sg13g2_decap_8 FILLER_70_422 ();
 sg13g2_decap_8 FILLER_70_429 ();
 sg13g2_fill_2 FILLER_70_436 ();
 sg13g2_fill_1 FILLER_70_438 ();
 sg13g2_fill_2 FILLER_70_460 ();
 sg13g2_fill_1 FILLER_70_462 ();
 sg13g2_decap_8 FILLER_70_479 ();
 sg13g2_decap_4 FILLER_70_486 ();
 sg13g2_fill_1 FILLER_70_494 ();
 sg13g2_fill_2 FILLER_70_517 ();
 sg13g2_fill_1 FILLER_70_519 ();
 sg13g2_fill_1 FILLER_70_530 ();
 sg13g2_decap_4 FILLER_70_537 ();
 sg13g2_fill_2 FILLER_70_541 ();
 sg13g2_fill_2 FILLER_70_562 ();
 sg13g2_fill_1 FILLER_70_564 ();
 sg13g2_fill_1 FILLER_70_600 ();
 sg13g2_fill_2 FILLER_70_613 ();
 sg13g2_fill_1 FILLER_70_615 ();
 sg13g2_decap_4 FILLER_70_691 ();
 sg13g2_fill_2 FILLER_70_695 ();
 sg13g2_decap_4 FILLER_70_702 ();
 sg13g2_decap_4 FILLER_70_802 ();
 sg13g2_fill_1 FILLER_70_806 ();
 sg13g2_decap_8 FILLER_70_820 ();
 sg13g2_decap_8 FILLER_70_827 ();
 sg13g2_decap_8 FILLER_70_834 ();
 sg13g2_decap_8 FILLER_70_841 ();
 sg13g2_decap_8 FILLER_70_848 ();
 sg13g2_decap_8 FILLER_70_855 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_4 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_43 ();
 sg13g2_decap_8 FILLER_71_50 ();
 sg13g2_decap_8 FILLER_71_57 ();
 sg13g2_decap_8 FILLER_71_64 ();
 sg13g2_decap_8 FILLER_71_71 ();
 sg13g2_fill_1 FILLER_71_127 ();
 sg13g2_decap_8 FILLER_71_145 ();
 sg13g2_fill_1 FILLER_71_152 ();
 sg13g2_fill_2 FILLER_71_163 ();
 sg13g2_fill_1 FILLER_71_165 ();
 sg13g2_fill_1 FILLER_71_208 ();
 sg13g2_decap_8 FILLER_71_217 ();
 sg13g2_fill_2 FILLER_71_224 ();
 sg13g2_fill_1 FILLER_71_226 ();
 sg13g2_decap_4 FILLER_71_255 ();
 sg13g2_fill_2 FILLER_71_269 ();
 sg13g2_fill_1 FILLER_71_271 ();
 sg13g2_fill_2 FILLER_71_298 ();
 sg13g2_fill_1 FILLER_71_340 ();
 sg13g2_decap_4 FILLER_71_366 ();
 sg13g2_fill_1 FILLER_71_370 ();
 sg13g2_fill_2 FILLER_71_397 ();
 sg13g2_fill_1 FILLER_71_436 ();
 sg13g2_decap_8 FILLER_71_448 ();
 sg13g2_decap_8 FILLER_71_455 ();
 sg13g2_decap_8 FILLER_71_462 ();
 sg13g2_decap_4 FILLER_71_469 ();
 sg13g2_fill_1 FILLER_71_473 ();
 sg13g2_fill_2 FILLER_71_479 ();
 sg13g2_fill_1 FILLER_71_481 ();
 sg13g2_fill_2 FILLER_71_485 ();
 sg13g2_fill_1 FILLER_71_487 ();
 sg13g2_fill_1 FILLER_71_504 ();
 sg13g2_fill_2 FILLER_71_512 ();
 sg13g2_fill_2 FILLER_71_522 ();
 sg13g2_fill_1 FILLER_71_532 ();
 sg13g2_decap_8 FILLER_71_546 ();
 sg13g2_fill_1 FILLER_71_553 ();
 sg13g2_decap_4 FILLER_71_579 ();
 sg13g2_fill_2 FILLER_71_583 ();
 sg13g2_fill_2 FILLER_71_597 ();
 sg13g2_fill_2 FILLER_71_687 ();
 sg13g2_fill_2 FILLER_71_704 ();
 sg13g2_fill_2 FILLER_71_712 ();
 sg13g2_fill_1 FILLER_71_714 ();
 sg13g2_fill_1 FILLER_71_745 ();
 sg13g2_fill_1 FILLER_71_752 ();
 sg13g2_fill_2 FILLER_71_766 ();
 sg13g2_fill_2 FILLER_71_773 ();
 sg13g2_decap_8 FILLER_71_806 ();
 sg13g2_decap_8 FILLER_71_813 ();
 sg13g2_decap_8 FILLER_71_820 ();
 sg13g2_decap_8 FILLER_71_827 ();
 sg13g2_decap_8 FILLER_71_834 ();
 sg13g2_decap_8 FILLER_71_841 ();
 sg13g2_decap_8 FILLER_71_848 ();
 sg13g2_decap_8 FILLER_71_855 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_fill_2 FILLER_72_84 ();
 sg13g2_fill_1 FILLER_72_86 ();
 sg13g2_fill_2 FILLER_72_97 ();
 sg13g2_fill_1 FILLER_72_99 ();
 sg13g2_fill_2 FILLER_72_105 ();
 sg13g2_fill_1 FILLER_72_107 ();
 sg13g2_fill_2 FILLER_72_133 ();
 sg13g2_fill_1 FILLER_72_135 ();
 sg13g2_fill_2 FILLER_72_146 ();
 sg13g2_fill_2 FILLER_72_161 ();
 sg13g2_fill_1 FILLER_72_163 ();
 sg13g2_decap_4 FILLER_72_179 ();
 sg13g2_fill_2 FILLER_72_199 ();
 sg13g2_fill_2 FILLER_72_227 ();
 sg13g2_fill_1 FILLER_72_229 ();
 sg13g2_fill_2 FILLER_72_259 ();
 sg13g2_fill_1 FILLER_72_261 ();
 sg13g2_fill_2 FILLER_72_316 ();
 sg13g2_fill_1 FILLER_72_318 ();
 sg13g2_fill_1 FILLER_72_338 ();
 sg13g2_decap_4 FILLER_72_365 ();
 sg13g2_fill_2 FILLER_72_369 ();
 sg13g2_decap_8 FILLER_72_375 ();
 sg13g2_fill_1 FILLER_72_382 ();
 sg13g2_fill_1 FILLER_72_422 ();
 sg13g2_fill_2 FILLER_72_506 ();
 sg13g2_decap_4 FILLER_72_533 ();
 sg13g2_fill_1 FILLER_72_537 ();
 sg13g2_fill_1 FILLER_72_547 ();
 sg13g2_fill_1 FILLER_72_551 ();
 sg13g2_decap_4 FILLER_72_581 ();
 sg13g2_fill_2 FILLER_72_740 ();
 sg13g2_fill_1 FILLER_72_742 ();
 sg13g2_decap_8 FILLER_72_807 ();
 sg13g2_decap_8 FILLER_72_814 ();
 sg13g2_decap_8 FILLER_72_821 ();
 sg13g2_decap_8 FILLER_72_828 ();
 sg13g2_decap_8 FILLER_72_835 ();
 sg13g2_decap_8 FILLER_72_842 ();
 sg13g2_decap_8 FILLER_72_849 ();
 sg13g2_decap_4 FILLER_72_856 ();
 sg13g2_fill_2 FILLER_72_860 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_4 FILLER_73_70 ();
 sg13g2_fill_2 FILLER_73_106 ();
 sg13g2_fill_1 FILLER_73_124 ();
 sg13g2_fill_2 FILLER_73_130 ();
 sg13g2_fill_1 FILLER_73_132 ();
 sg13g2_fill_2 FILLER_73_138 ();
 sg13g2_fill_1 FILLER_73_149 ();
 sg13g2_fill_2 FILLER_73_165 ();
 sg13g2_fill_1 FILLER_73_167 ();
 sg13g2_fill_2 FILLER_73_178 ();
 sg13g2_fill_1 FILLER_73_195 ();
 sg13g2_fill_2 FILLER_73_205 ();
 sg13g2_fill_1 FILLER_73_212 ();
 sg13g2_decap_4 FILLER_73_218 ();
 sg13g2_decap_4 FILLER_73_228 ();
 sg13g2_fill_1 FILLER_73_232 ();
 sg13g2_fill_2 FILLER_73_249 ();
 sg13g2_fill_1 FILLER_73_251 ();
 sg13g2_fill_2 FILLER_73_271 ();
 sg13g2_fill_1 FILLER_73_273 ();
 sg13g2_fill_2 FILLER_73_328 ();
 sg13g2_fill_2 FILLER_73_387 ();
 sg13g2_fill_2 FILLER_73_403 ();
 sg13g2_fill_1 FILLER_73_409 ();
 sg13g2_fill_1 FILLER_73_455 ();
 sg13g2_decap_8 FILLER_73_468 ();
 sg13g2_decap_4 FILLER_73_475 ();
 sg13g2_fill_1 FILLER_73_479 ();
 sg13g2_fill_1 FILLER_73_497 ();
 sg13g2_fill_1 FILLER_73_571 ();
 sg13g2_fill_2 FILLER_73_594 ();
 sg13g2_fill_2 FILLER_73_609 ();
 sg13g2_fill_1 FILLER_73_620 ();
 sg13g2_fill_1 FILLER_73_629 ();
 sg13g2_fill_1 FILLER_73_657 ();
 sg13g2_fill_2 FILLER_73_667 ();
 sg13g2_fill_1 FILLER_73_678 ();
 sg13g2_fill_1 FILLER_73_731 ();
 sg13g2_decap_8 FILLER_73_807 ();
 sg13g2_decap_8 FILLER_73_814 ();
 sg13g2_decap_8 FILLER_73_821 ();
 sg13g2_decap_8 FILLER_73_828 ();
 sg13g2_decap_8 FILLER_73_835 ();
 sg13g2_decap_8 FILLER_73_842 ();
 sg13g2_decap_8 FILLER_73_849 ();
 sg13g2_decap_4 FILLER_73_856 ();
 sg13g2_fill_2 FILLER_73_860 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_4 FILLER_74_63 ();
 sg13g2_fill_2 FILLER_74_82 ();
 sg13g2_fill_2 FILLER_74_89 ();
 sg13g2_fill_2 FILLER_74_100 ();
 sg13g2_fill_2 FILLER_74_108 ();
 sg13g2_fill_1 FILLER_74_110 ();
 sg13g2_fill_2 FILLER_74_124 ();
 sg13g2_fill_1 FILLER_74_146 ();
 sg13g2_fill_2 FILLER_74_157 ();
 sg13g2_fill_1 FILLER_74_159 ();
 sg13g2_decap_4 FILLER_74_173 ();
 sg13g2_fill_2 FILLER_74_177 ();
 sg13g2_fill_2 FILLER_74_189 ();
 sg13g2_fill_2 FILLER_74_207 ();
 sg13g2_fill_1 FILLER_74_209 ();
 sg13g2_fill_1 FILLER_74_220 ();
 sg13g2_fill_1 FILLER_74_235 ();
 sg13g2_fill_1 FILLER_74_241 ();
 sg13g2_decap_8 FILLER_74_247 ();
 sg13g2_decap_4 FILLER_74_259 ();
 sg13g2_fill_2 FILLER_74_263 ();
 sg13g2_decap_8 FILLER_74_279 ();
 sg13g2_fill_2 FILLER_74_286 ();
 sg13g2_fill_2 FILLER_74_293 ();
 sg13g2_fill_1 FILLER_74_295 ();
 sg13g2_fill_1 FILLER_74_354 ();
 sg13g2_fill_2 FILLER_74_369 ();
 sg13g2_fill_1 FILLER_74_371 ();
 sg13g2_decap_8 FILLER_74_420 ();
 sg13g2_decap_4 FILLER_74_427 ();
 sg13g2_decap_4 FILLER_74_435 ();
 sg13g2_fill_1 FILLER_74_439 ();
 sg13g2_fill_2 FILLER_74_471 ();
 sg13g2_fill_2 FILLER_74_534 ();
 sg13g2_fill_1 FILLER_74_536 ();
 sg13g2_fill_1 FILLER_74_548 ();
 sg13g2_fill_2 FILLER_74_692 ();
 sg13g2_fill_2 FILLER_74_789 ();
 sg13g2_decap_8 FILLER_74_803 ();
 sg13g2_decap_8 FILLER_74_810 ();
 sg13g2_decap_8 FILLER_74_817 ();
 sg13g2_decap_8 FILLER_74_824 ();
 sg13g2_decap_8 FILLER_74_831 ();
 sg13g2_decap_8 FILLER_74_838 ();
 sg13g2_decap_8 FILLER_74_845 ();
 sg13g2_decap_8 FILLER_74_852 ();
 sg13g2_fill_2 FILLER_74_859 ();
 sg13g2_fill_1 FILLER_74_861 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_4 FILLER_75_70 ();
 sg13g2_fill_2 FILLER_75_74 ();
 sg13g2_fill_2 FILLER_75_81 ();
 sg13g2_fill_2 FILLER_75_89 ();
 sg13g2_fill_1 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_fill_1 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_164 ();
 sg13g2_fill_1 FILLER_75_171 ();
 sg13g2_decap_4 FILLER_75_191 ();
 sg13g2_fill_2 FILLER_75_195 ();
 sg13g2_fill_2 FILLER_75_217 ();
 sg13g2_fill_1 FILLER_75_223 ();
 sg13g2_fill_1 FILLER_75_230 ();
 sg13g2_fill_2 FILLER_75_250 ();
 sg13g2_fill_1 FILLER_75_252 ();
 sg13g2_decap_4 FILLER_75_275 ();
 sg13g2_decap_4 FILLER_75_285 ();
 sg13g2_fill_2 FILLER_75_289 ();
 sg13g2_fill_2 FILLER_75_386 ();
 sg13g2_fill_1 FILLER_75_397 ();
 sg13g2_decap_4 FILLER_75_402 ();
 sg13g2_decap_4 FILLER_75_415 ();
 sg13g2_fill_1 FILLER_75_419 ();
 sg13g2_fill_1 FILLER_75_435 ();
 sg13g2_decap_4 FILLER_75_464 ();
 sg13g2_fill_1 FILLER_75_468 ();
 sg13g2_decap_4 FILLER_75_473 ();
 sg13g2_fill_1 FILLER_75_477 ();
 sg13g2_fill_1 FILLER_75_496 ();
 sg13g2_fill_2 FILLER_75_501 ();
 sg13g2_fill_1 FILLER_75_566 ();
 sg13g2_fill_1 FILLER_75_603 ();
 sg13g2_fill_2 FILLER_75_610 ();
 sg13g2_fill_2 FILLER_75_621 ();
 sg13g2_fill_1 FILLER_75_636 ();
 sg13g2_fill_2 FILLER_75_653 ();
 sg13g2_fill_2 FILLER_75_664 ();
 sg13g2_fill_1 FILLER_75_671 ();
 sg13g2_fill_2 FILLER_75_742 ();
 sg13g2_decap_8 FILLER_75_752 ();
 sg13g2_decap_8 FILLER_75_759 ();
 sg13g2_decap_8 FILLER_75_780 ();
 sg13g2_decap_8 FILLER_75_787 ();
 sg13g2_decap_8 FILLER_75_794 ();
 sg13g2_decap_8 FILLER_75_801 ();
 sg13g2_decap_8 FILLER_75_808 ();
 sg13g2_decap_8 FILLER_75_815 ();
 sg13g2_decap_8 FILLER_75_822 ();
 sg13g2_decap_8 FILLER_75_829 ();
 sg13g2_decap_8 FILLER_75_836 ();
 sg13g2_decap_8 FILLER_75_843 ();
 sg13g2_decap_8 FILLER_75_850 ();
 sg13g2_decap_4 FILLER_75_857 ();
 sg13g2_fill_1 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_fill_2 FILLER_76_63 ();
 sg13g2_fill_1 FILLER_76_85 ();
 sg13g2_decap_8 FILLER_76_100 ();
 sg13g2_fill_1 FILLER_76_107 ();
 sg13g2_fill_2 FILLER_76_126 ();
 sg13g2_fill_1 FILLER_76_128 ();
 sg13g2_decap_8 FILLER_76_134 ();
 sg13g2_decap_8 FILLER_76_141 ();
 sg13g2_decap_4 FILLER_76_172 ();
 sg13g2_fill_2 FILLER_76_176 ();
 sg13g2_fill_2 FILLER_76_196 ();
 sg13g2_fill_1 FILLER_76_212 ();
 sg13g2_fill_2 FILLER_76_217 ();
 sg13g2_fill_2 FILLER_76_232 ();
 sg13g2_decap_4 FILLER_76_238 ();
 sg13g2_fill_1 FILLER_76_246 ();
 sg13g2_fill_1 FILLER_76_265 ();
 sg13g2_decap_8 FILLER_76_292 ();
 sg13g2_fill_2 FILLER_76_299 ();
 sg13g2_fill_1 FILLER_76_301 ();
 sg13g2_fill_1 FILLER_76_311 ();
 sg13g2_fill_1 FILLER_76_326 ();
 sg13g2_fill_2 FILLER_76_351 ();
 sg13g2_fill_1 FILLER_76_353 ();
 sg13g2_fill_1 FILLER_76_359 ();
 sg13g2_fill_1 FILLER_76_380 ();
 sg13g2_fill_2 FILLER_76_386 ();
 sg13g2_fill_1 FILLER_76_388 ();
 sg13g2_fill_1 FILLER_76_415 ();
 sg13g2_fill_1 FILLER_76_450 ();
 sg13g2_fill_2 FILLER_76_477 ();
 sg13g2_fill_1 FILLER_76_479 ();
 sg13g2_fill_2 FILLER_76_489 ();
 sg13g2_fill_1 FILLER_76_491 ();
 sg13g2_fill_1 FILLER_76_505 ();
 sg13g2_fill_2 FILLER_76_528 ();
 sg13g2_fill_2 FILLER_76_538 ();
 sg13g2_fill_1 FILLER_76_594 ();
 sg13g2_decap_4 FILLER_76_631 ();
 sg13g2_fill_1 FILLER_76_635 ();
 sg13g2_fill_2 FILLER_76_688 ();
 sg13g2_fill_2 FILLER_76_695 ();
 sg13g2_fill_1 FILLER_76_708 ();
 sg13g2_decap_8 FILLER_76_744 ();
 sg13g2_decap_8 FILLER_76_751 ();
 sg13g2_decap_8 FILLER_76_758 ();
 sg13g2_decap_8 FILLER_76_765 ();
 sg13g2_decap_8 FILLER_76_772 ();
 sg13g2_decap_8 FILLER_76_779 ();
 sg13g2_decap_8 FILLER_76_786 ();
 sg13g2_decap_8 FILLER_76_793 ();
 sg13g2_decap_8 FILLER_76_800 ();
 sg13g2_decap_8 FILLER_76_807 ();
 sg13g2_decap_8 FILLER_76_814 ();
 sg13g2_decap_8 FILLER_76_821 ();
 sg13g2_decap_8 FILLER_76_828 ();
 sg13g2_decap_8 FILLER_76_835 ();
 sg13g2_decap_8 FILLER_76_842 ();
 sg13g2_decap_8 FILLER_76_849 ();
 sg13g2_decap_4 FILLER_76_856 ();
 sg13g2_fill_2 FILLER_76_860 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_4 FILLER_77_63 ();
 sg13g2_fill_1 FILLER_77_67 ();
 sg13g2_fill_2 FILLER_77_90 ();
 sg13g2_fill_1 FILLER_77_92 ();
 sg13g2_fill_2 FILLER_77_103 ();
 sg13g2_fill_1 FILLER_77_122 ();
 sg13g2_decap_8 FILLER_77_148 ();
 sg13g2_fill_1 FILLER_77_161 ();
 sg13g2_fill_1 FILLER_77_168 ();
 sg13g2_decap_4 FILLER_77_180 ();
 sg13g2_fill_1 FILLER_77_221 ();
 sg13g2_fill_1 FILLER_77_227 ();
 sg13g2_decap_4 FILLER_77_233 ();
 sg13g2_fill_1 FILLER_77_247 ();
 sg13g2_fill_2 FILLER_77_253 ();
 sg13g2_fill_1 FILLER_77_255 ();
 sg13g2_fill_2 FILLER_77_264 ();
 sg13g2_fill_1 FILLER_77_271 ();
 sg13g2_fill_1 FILLER_77_281 ();
 sg13g2_fill_2 FILLER_77_287 ();
 sg13g2_fill_2 FILLER_77_299 ();
 sg13g2_fill_1 FILLER_77_305 ();
 sg13g2_fill_2 FILLER_77_310 ();
 sg13g2_fill_1 FILLER_77_312 ();
 sg13g2_fill_2 FILLER_77_374 ();
 sg13g2_fill_1 FILLER_77_376 ();
 sg13g2_fill_2 FILLER_77_410 ();
 sg13g2_fill_2 FILLER_77_416 ();
 sg13g2_fill_1 FILLER_77_418 ();
 sg13g2_fill_2 FILLER_77_433 ();
 sg13g2_fill_1 FILLER_77_435 ();
 sg13g2_decap_8 FILLER_77_470 ();
 sg13g2_fill_1 FILLER_77_539 ();
 sg13g2_fill_2 FILLER_77_569 ();
 sg13g2_fill_1 FILLER_77_612 ();
 sg13g2_fill_2 FILLER_77_674 ();
 sg13g2_fill_1 FILLER_77_676 ();
 sg13g2_fill_2 FILLER_77_686 ();
 sg13g2_fill_2 FILLER_77_723 ();
 sg13g2_fill_1 FILLER_77_725 ();
 sg13g2_decap_8 FILLER_77_735 ();
 sg13g2_decap_8 FILLER_77_742 ();
 sg13g2_decap_8 FILLER_77_749 ();
 sg13g2_decap_8 FILLER_77_756 ();
 sg13g2_decap_8 FILLER_77_763 ();
 sg13g2_decap_8 FILLER_77_770 ();
 sg13g2_decap_8 FILLER_77_777 ();
 sg13g2_decap_8 FILLER_77_784 ();
 sg13g2_decap_8 FILLER_77_791 ();
 sg13g2_decap_8 FILLER_77_798 ();
 sg13g2_decap_8 FILLER_77_805 ();
 sg13g2_decap_8 FILLER_77_812 ();
 sg13g2_decap_8 FILLER_77_819 ();
 sg13g2_decap_8 FILLER_77_826 ();
 sg13g2_decap_8 FILLER_77_833 ();
 sg13g2_decap_8 FILLER_77_840 ();
 sg13g2_decap_8 FILLER_77_847 ();
 sg13g2_decap_8 FILLER_77_854 ();
 sg13g2_fill_1 FILLER_77_861 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_4 FILLER_78_56 ();
 sg13g2_fill_2 FILLER_78_60 ();
 sg13g2_decap_8 FILLER_78_66 ();
 sg13g2_decap_4 FILLER_78_73 ();
 sg13g2_fill_2 FILLER_78_91 ();
 sg13g2_fill_1 FILLER_78_93 ();
 sg13g2_fill_2 FILLER_78_109 ();
 sg13g2_fill_2 FILLER_78_144 ();
 sg13g2_decap_8 FILLER_78_151 ();
 sg13g2_decap_4 FILLER_78_158 ();
 sg13g2_fill_2 FILLER_78_172 ();
 sg13g2_fill_1 FILLER_78_174 ();
 sg13g2_decap_4 FILLER_78_193 ();
 sg13g2_fill_2 FILLER_78_197 ();
 sg13g2_decap_4 FILLER_78_213 ();
 sg13g2_fill_2 FILLER_78_222 ();
 sg13g2_fill_2 FILLER_78_238 ();
 sg13g2_fill_1 FILLER_78_260 ();
 sg13g2_fill_1 FILLER_78_266 ();
 sg13g2_decap_4 FILLER_78_286 ();
 sg13g2_fill_2 FILLER_78_377 ();
 sg13g2_fill_2 FILLER_78_406 ();
 sg13g2_fill_2 FILLER_78_450 ();
 sg13g2_fill_1 FILLER_78_478 ();
 sg13g2_decap_4 FILLER_78_483 ();
 sg13g2_fill_1 FILLER_78_487 ();
 sg13g2_fill_1 FILLER_78_497 ();
 sg13g2_fill_1 FILLER_78_514 ();
 sg13g2_fill_1 FILLER_78_565 ();
 sg13g2_fill_1 FILLER_78_613 ();
 sg13g2_fill_1 FILLER_78_633 ();
 sg13g2_fill_1 FILLER_78_660 ();
 sg13g2_fill_2 FILLER_78_696 ();
 sg13g2_fill_1 FILLER_78_698 ();
 sg13g2_fill_2 FILLER_78_706 ();
 sg13g2_fill_1 FILLER_78_708 ();
 sg13g2_decap_4 FILLER_78_720 ();
 sg13g2_fill_1 FILLER_78_724 ();
 sg13g2_decap_8 FILLER_78_729 ();
 sg13g2_decap_8 FILLER_78_736 ();
 sg13g2_decap_8 FILLER_78_743 ();
 sg13g2_decap_8 FILLER_78_750 ();
 sg13g2_decap_8 FILLER_78_757 ();
 sg13g2_decap_8 FILLER_78_764 ();
 sg13g2_decap_8 FILLER_78_771 ();
 sg13g2_decap_8 FILLER_78_778 ();
 sg13g2_decap_8 FILLER_78_785 ();
 sg13g2_decap_8 FILLER_78_792 ();
 sg13g2_decap_8 FILLER_78_799 ();
 sg13g2_decap_8 FILLER_78_806 ();
 sg13g2_decap_8 FILLER_78_813 ();
 sg13g2_decap_8 FILLER_78_820 ();
 sg13g2_decap_8 FILLER_78_827 ();
 sg13g2_decap_8 FILLER_78_834 ();
 sg13g2_decap_8 FILLER_78_841 ();
 sg13g2_decap_8 FILLER_78_848 ();
 sg13g2_decap_8 FILLER_78_855 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_fill_2 FILLER_79_49 ();
 sg13g2_fill_1 FILLER_79_87 ();
 sg13g2_decap_4 FILLER_79_108 ();
 sg13g2_fill_1 FILLER_79_142 ();
 sg13g2_decap_4 FILLER_79_149 ();
 sg13g2_fill_2 FILLER_79_168 ();
 sg13g2_fill_2 FILLER_79_206 ();
 sg13g2_fill_1 FILLER_79_208 ();
 sg13g2_fill_2 FILLER_79_225 ();
 sg13g2_fill_2 FILLER_79_233 ();
 sg13g2_decap_8 FILLER_79_241 ();
 sg13g2_fill_2 FILLER_79_248 ();
 sg13g2_fill_1 FILLER_79_250 ();
 sg13g2_fill_1 FILLER_79_269 ();
 sg13g2_fill_1 FILLER_79_305 ();
 sg13g2_fill_2 FILLER_79_384 ();
 sg13g2_fill_1 FILLER_79_386 ();
 sg13g2_fill_2 FILLER_79_397 ();
 sg13g2_fill_1 FILLER_79_399 ();
 sg13g2_fill_2 FILLER_79_422 ();
 sg13g2_fill_2 FILLER_79_450 ();
 sg13g2_decap_8 FILLER_79_456 ();
 sg13g2_decap_8 FILLER_79_467 ();
 sg13g2_decap_4 FILLER_79_500 ();
 sg13g2_fill_2 FILLER_79_504 ();
 sg13g2_fill_2 FILLER_79_518 ();
 sg13g2_fill_1 FILLER_79_543 ();
 sg13g2_fill_2 FILLER_79_584 ();
 sg13g2_decap_4 FILLER_79_641 ();
 sg13g2_fill_2 FILLER_79_649 ();
 sg13g2_fill_1 FILLER_79_680 ();
 sg13g2_decap_8 FILLER_79_685 ();
 sg13g2_decap_8 FILLER_79_692 ();
 sg13g2_decap_8 FILLER_79_699 ();
 sg13g2_decap_8 FILLER_79_706 ();
 sg13g2_decap_8 FILLER_79_713 ();
 sg13g2_decap_8 FILLER_79_720 ();
 sg13g2_decap_8 FILLER_79_727 ();
 sg13g2_decap_8 FILLER_79_734 ();
 sg13g2_decap_8 FILLER_79_741 ();
 sg13g2_decap_8 FILLER_79_748 ();
 sg13g2_decap_8 FILLER_79_755 ();
 sg13g2_decap_8 FILLER_79_762 ();
 sg13g2_decap_8 FILLER_79_769 ();
 sg13g2_decap_8 FILLER_79_776 ();
 sg13g2_decap_8 FILLER_79_783 ();
 sg13g2_decap_8 FILLER_79_790 ();
 sg13g2_decap_8 FILLER_79_797 ();
 sg13g2_decap_8 FILLER_79_804 ();
 sg13g2_decap_8 FILLER_79_811 ();
 sg13g2_decap_8 FILLER_79_818 ();
 sg13g2_decap_8 FILLER_79_825 ();
 sg13g2_decap_8 FILLER_79_832 ();
 sg13g2_decap_8 FILLER_79_839 ();
 sg13g2_decap_8 FILLER_79_846 ();
 sg13g2_decap_8 FILLER_79_853 ();
 sg13g2_fill_2 FILLER_79_860 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_fill_1 FILLER_80_68 ();
 sg13g2_decap_8 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_112 ();
 sg13g2_fill_1 FILLER_80_121 ();
 sg13g2_decap_4 FILLER_80_133 ();
 sg13g2_fill_2 FILLER_80_142 ();
 sg13g2_decap_8 FILLER_80_154 ();
 sg13g2_decap_8 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_171 ();
 sg13g2_fill_2 FILLER_80_175 ();
 sg13g2_fill_1 FILLER_80_184 ();
 sg13g2_decap_8 FILLER_80_195 ();
 sg13g2_fill_2 FILLER_80_202 ();
 sg13g2_fill_1 FILLER_80_204 ();
 sg13g2_decap_4 FILLER_80_210 ();
 sg13g2_decap_4 FILLER_80_224 ();
 sg13g2_decap_4 FILLER_80_238 ();
 sg13g2_fill_2 FILLER_80_242 ();
 sg13g2_fill_2 FILLER_80_280 ();
 sg13g2_fill_2 FILLER_80_358 ();
 sg13g2_fill_2 FILLER_80_372 ();
 sg13g2_fill_1 FILLER_80_408 ();
 sg13g2_fill_2 FILLER_80_439 ();
 sg13g2_fill_1 FILLER_80_467 ();
 sg13g2_fill_1 FILLER_80_494 ();
 sg13g2_fill_1 FILLER_80_521 ();
 sg13g2_fill_1 FILLER_80_557 ();
 sg13g2_decap_8 FILLER_80_634 ();
 sg13g2_decap_8 FILLER_80_641 ();
 sg13g2_decap_8 FILLER_80_648 ();
 sg13g2_decap_8 FILLER_80_655 ();
 sg13g2_decap_8 FILLER_80_662 ();
 sg13g2_decap_8 FILLER_80_669 ();
 sg13g2_decap_8 FILLER_80_676 ();
 sg13g2_decap_8 FILLER_80_683 ();
 sg13g2_decap_8 FILLER_80_690 ();
 sg13g2_decap_8 FILLER_80_697 ();
 sg13g2_decap_8 FILLER_80_704 ();
 sg13g2_decap_8 FILLER_80_711 ();
 sg13g2_decap_8 FILLER_80_718 ();
 sg13g2_decap_8 FILLER_80_725 ();
 sg13g2_decap_8 FILLER_80_732 ();
 sg13g2_decap_8 FILLER_80_739 ();
 sg13g2_decap_8 FILLER_80_746 ();
 sg13g2_decap_8 FILLER_80_753 ();
 sg13g2_decap_8 FILLER_80_760 ();
 sg13g2_decap_8 FILLER_80_767 ();
 sg13g2_decap_8 FILLER_80_774 ();
 sg13g2_decap_8 FILLER_80_781 ();
 sg13g2_decap_8 FILLER_80_788 ();
 sg13g2_decap_8 FILLER_80_795 ();
 sg13g2_decap_8 FILLER_80_802 ();
 sg13g2_decap_8 FILLER_80_809 ();
 sg13g2_decap_8 FILLER_80_816 ();
 sg13g2_decap_8 FILLER_80_823 ();
 sg13g2_decap_8 FILLER_80_830 ();
 sg13g2_decap_8 FILLER_80_837 ();
 sg13g2_decap_8 FILLER_80_844 ();
 sg13g2_decap_8 FILLER_80_851 ();
 sg13g2_decap_4 FILLER_80_858 ();
 assign uio_oe[6] = net316;
 assign uio_oe[7] = net317;
endmodule

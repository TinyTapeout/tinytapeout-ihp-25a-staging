module tt_um_gfg_development_tinymandelbrot (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire clk_regs;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire _2568_;
 wire combined_rst_n;
 wire \configuration[0] ;
 wire \configuration[10] ;
 wire \configuration[11] ;
 wire \configuration[12] ;
 wire \configuration[13] ;
 wire \configuration[14] ;
 wire \configuration[15] ;
 wire \configuration[16] ;
 wire \configuration[17] ;
 wire \configuration[18] ;
 wire \configuration[19] ;
 wire \configuration[1] ;
 wire \configuration[20] ;
 wire \configuration[21] ;
 wire \configuration[22] ;
 wire \configuration[23] ;
 wire \configuration[24] ;
 wire \configuration[25] ;
 wire \configuration[26] ;
 wire \configuration[27] ;
 wire \configuration[28] ;
 wire \configuration[29] ;
 wire \configuration[2] ;
 wire \configuration[30] ;
 wire \configuration[31] ;
 wire \configuration[32] ;
 wire \configuration[33] ;
 wire \configuration[34] ;
 wire \configuration[35] ;
 wire \configuration[36] ;
 wire \configuration[37] ;
 wire \configuration[38] ;
 wire \configuration[39] ;
 wire \configuration[3] ;
 wire \configuration[40] ;
 wire \configuration[41] ;
 wire \configuration[42] ;
 wire \configuration[43] ;
 wire \configuration[44] ;
 wire \configuration[45] ;
 wire \configuration[46] ;
 wire \configuration[47] ;
 wire \configuration[48] ;
 wire \configuration[49] ;
 wire \configuration[4] ;
 wire \configuration[50] ;
 wire \configuration[51] ;
 wire \configuration[52] ;
 wire \configuration[5] ;
 wire \configuration[6] ;
 wire \configuration[7] ;
 wire \configuration[8] ;
 wire \configuration[9] ;
 wire finished;
 wire l_running;
 wire \l_sclk[0] ;
 wire \l_sclk[1] ;
 wire \l_sclk[2] ;
 wire \l_sdata[0] ;
 wire \l_sdata[1] ;
 wire \l_sdata[2] ;
 wire \l_sen[0] ;
 wire \l_sen[1] ;
 wire \l_sen[2] ;
 wire latched_rst_n;
 wire \mandelbrot.alu.finished ;
 wire \mandelbrot.alu.first_iteration ;
 wire \mandelbrot.alu.in_ci[0] ;
 wire \mandelbrot.alu.in_ci[10] ;
 wire \mandelbrot.alu.in_ci[11] ;
 wire \mandelbrot.alu.in_ci[12] ;
 wire \mandelbrot.alu.in_ci[13] ;
 wire \mandelbrot.alu.in_ci[14] ;
 wire \mandelbrot.alu.in_ci[15] ;
 wire \mandelbrot.alu.in_ci[1] ;
 wire \mandelbrot.alu.in_ci[2] ;
 wire \mandelbrot.alu.in_ci[3] ;
 wire \mandelbrot.alu.in_ci[4] ;
 wire \mandelbrot.alu.in_ci[5] ;
 wire \mandelbrot.alu.in_ci[6] ;
 wire \mandelbrot.alu.in_ci[7] ;
 wire \mandelbrot.alu.in_ci[8] ;
 wire \mandelbrot.alu.in_ci[9] ;
 wire \mandelbrot.alu.in_cr[0] ;
 wire \mandelbrot.alu.in_cr[10] ;
 wire \mandelbrot.alu.in_cr[11] ;
 wire \mandelbrot.alu.in_cr[12] ;
 wire \mandelbrot.alu.in_cr[13] ;
 wire \mandelbrot.alu.in_cr[14] ;
 wire \mandelbrot.alu.in_cr[15] ;
 wire \mandelbrot.alu.in_cr[1] ;
 wire \mandelbrot.alu.in_cr[2] ;
 wire \mandelbrot.alu.in_cr[3] ;
 wire \mandelbrot.alu.in_cr[4] ;
 wire \mandelbrot.alu.in_cr[5] ;
 wire \mandelbrot.alu.in_cr[6] ;
 wire \mandelbrot.alu.in_cr[7] ;
 wire \mandelbrot.alu.in_cr[8] ;
 wire \mandelbrot.alu.in_cr[9] ;
 wire \mandelbrot.alu.in_zi[0] ;
 wire \mandelbrot.alu.in_zi[10] ;
 wire \mandelbrot.alu.in_zi[11] ;
 wire \mandelbrot.alu.in_zi[12] ;
 wire \mandelbrot.alu.in_zi[13] ;
 wire \mandelbrot.alu.in_zi[14] ;
 wire \mandelbrot.alu.in_zi[15] ;
 wire \mandelbrot.alu.in_zi[1] ;
 wire \mandelbrot.alu.in_zi[2] ;
 wire \mandelbrot.alu.in_zi[3] ;
 wire \mandelbrot.alu.in_zi[4] ;
 wire \mandelbrot.alu.in_zi[5] ;
 wire \mandelbrot.alu.in_zi[6] ;
 wire \mandelbrot.alu.in_zi[7] ;
 wire \mandelbrot.alu.in_zi[8] ;
 wire \mandelbrot.alu.in_zi[9] ;
 wire \mandelbrot.alu.in_zr[0] ;
 wire \mandelbrot.alu.in_zr[10] ;
 wire \mandelbrot.alu.in_zr[11] ;
 wire \mandelbrot.alu.in_zr[12] ;
 wire \mandelbrot.alu.in_zr[13] ;
 wire \mandelbrot.alu.in_zr[14] ;
 wire \mandelbrot.alu.in_zr[15] ;
 wire \mandelbrot.alu.in_zr[1] ;
 wire \mandelbrot.alu.in_zr[2] ;
 wire \mandelbrot.alu.in_zr[3] ;
 wire \mandelbrot.alu.in_zr[4] ;
 wire \mandelbrot.alu.in_zr[5] ;
 wire \mandelbrot.alu.in_zr[6] ;
 wire \mandelbrot.alu.in_zr[7] ;
 wire \mandelbrot.alu.in_zr[8] ;
 wire \mandelbrot.alu.in_zr[9] ;
 wire \mandelbrot.alu.m1[0] ;
 wire \mandelbrot.alu.m1[10] ;
 wire \mandelbrot.alu.m1[11] ;
 wire \mandelbrot.alu.m1[12] ;
 wire \mandelbrot.alu.m1[13] ;
 wire \mandelbrot.alu.m1[14] ;
 wire \mandelbrot.alu.m1[15] ;
 wire \mandelbrot.alu.m1[16] ;
 wire \mandelbrot.alu.m1[17] ;
 wire \mandelbrot.alu.m1[18] ;
 wire \mandelbrot.alu.m1[19] ;
 wire \mandelbrot.alu.m1[1] ;
 wire \mandelbrot.alu.m1[20] ;
 wire \mandelbrot.alu.m1[21] ;
 wire \mandelbrot.alu.m1[22] ;
 wire \mandelbrot.alu.m1[23] ;
 wire \mandelbrot.alu.m1[24] ;
 wire \mandelbrot.alu.m1[25] ;
 wire \mandelbrot.alu.m1[26] ;
 wire \mandelbrot.alu.m1[27] ;
 wire \mandelbrot.alu.m1[28] ;
 wire \mandelbrot.alu.m1[29] ;
 wire \mandelbrot.alu.m1[2] ;
 wire \mandelbrot.alu.m1[30] ;
 wire \mandelbrot.alu.m1[31] ;
 wire \mandelbrot.alu.m1[3] ;
 wire \mandelbrot.alu.m1[4] ;
 wire \mandelbrot.alu.m1[5] ;
 wire \mandelbrot.alu.m1[6] ;
 wire \mandelbrot.alu.m1[7] ;
 wire \mandelbrot.alu.m1[8] ;
 wire \mandelbrot.alu.m1[9] ;
 wire \mandelbrot.alu.m2[0] ;
 wire \mandelbrot.alu.m2[10] ;
 wire \mandelbrot.alu.m2[11] ;
 wire \mandelbrot.alu.m2[12] ;
 wire \mandelbrot.alu.m2[13] ;
 wire \mandelbrot.alu.m2[14] ;
 wire \mandelbrot.alu.m2[15] ;
 wire \mandelbrot.alu.m2[16] ;
 wire \mandelbrot.alu.m2[17] ;
 wire \mandelbrot.alu.m2[18] ;
 wire \mandelbrot.alu.m2[19] ;
 wire \mandelbrot.alu.m2[1] ;
 wire \mandelbrot.alu.m2[20] ;
 wire \mandelbrot.alu.m2[21] ;
 wire \mandelbrot.alu.m2[22] ;
 wire \mandelbrot.alu.m2[23] ;
 wire \mandelbrot.alu.m2[24] ;
 wire \mandelbrot.alu.m2[25] ;
 wire \mandelbrot.alu.m2[26] ;
 wire \mandelbrot.alu.m2[27] ;
 wire \mandelbrot.alu.m2[28] ;
 wire \mandelbrot.alu.m2[29] ;
 wire \mandelbrot.alu.m2[2] ;
 wire \mandelbrot.alu.m2[30] ;
 wire \mandelbrot.alu.m2[31] ;
 wire \mandelbrot.alu.m2[3] ;
 wire \mandelbrot.alu.m2[4] ;
 wire \mandelbrot.alu.m2[5] ;
 wire \mandelbrot.alu.m2[6] ;
 wire \mandelbrot.alu.m2[7] ;
 wire \mandelbrot.alu.m2[8] ;
 wire \mandelbrot.alu.m2[9] ;
 wire \mandelbrot.alu.m3[0] ;
 wire \mandelbrot.alu.m3[10] ;
 wire \mandelbrot.alu.m3[11] ;
 wire \mandelbrot.alu.m3[12] ;
 wire \mandelbrot.alu.m3[13] ;
 wire \mandelbrot.alu.m3[14] ;
 wire \mandelbrot.alu.m3[15] ;
 wire \mandelbrot.alu.m3[16] ;
 wire \mandelbrot.alu.m3[17] ;
 wire \mandelbrot.alu.m3[18] ;
 wire \mandelbrot.alu.m3[19] ;
 wire \mandelbrot.alu.m3[1] ;
 wire \mandelbrot.alu.m3[20] ;
 wire \mandelbrot.alu.m3[21] ;
 wire \mandelbrot.alu.m3[22] ;
 wire \mandelbrot.alu.m3[23] ;
 wire \mandelbrot.alu.m3[24] ;
 wire \mandelbrot.alu.m3[25] ;
 wire \mandelbrot.alu.m3[26] ;
 wire \mandelbrot.alu.m3[27] ;
 wire \mandelbrot.alu.m3[28] ;
 wire \mandelbrot.alu.m3[29] ;
 wire \mandelbrot.alu.m3[2] ;
 wire \mandelbrot.alu.m3[30] ;
 wire \mandelbrot.alu.m3[31] ;
 wire \mandelbrot.alu.m3[3] ;
 wire \mandelbrot.alu.m3[4] ;
 wire \mandelbrot.alu.m3[5] ;
 wire \mandelbrot.alu.m3[6] ;
 wire \mandelbrot.alu.m3[7] ;
 wire \mandelbrot.alu.m3[8] ;
 wire \mandelbrot.alu.m3[9] ;
 wire \mandelbrot.alu.mult_zi_zi.ctr[0] ;
 wire \mandelbrot.alu.mult_zi_zi.ctr[1] ;
 wire \mandelbrot.alu.mult_zi_zi.ctr[2] ;
 wire \mandelbrot.alu.mult_zi_zi.running ;
 wire \mandelbrot.alu.mult_zi_zi.shift_reg[0] ;
 wire \mandelbrot.alu.mult_zr_zi.ctr[0] ;
 wire \mandelbrot.alu.mult_zr_zi.ctr[1] ;
 wire \mandelbrot.alu.mult_zr_zi.ctr[2] ;
 wire \mandelbrot.alu.mult_zr_zi.running ;
 wire \mandelbrot.alu.mult_zr_zi.shift_reg[0] ;
 wire \mandelbrot.alu.mult_zr_zr.ctr[0] ;
 wire \mandelbrot.alu.mult_zr_zr.ctr[1] ;
 wire \mandelbrot.alu.mult_zr_zr.ctr[2] ;
 wire \mandelbrot.alu.mult_zr_zr.running ;
 wire \mandelbrot.alu.mult_zr_zr.shift_reg[0] ;
 wire \mandelbrot.ctr[0] ;
 wire \mandelbrot.ctr[1] ;
 wire \mandelbrot.ctr[2] ;
 wire \mandelbrot.ctr[3] ;
 wire \mandelbrot.ctr[4] ;
 wire \mandelbrot.ctr[5] ;
 wire \mandelbrot.ctr[6] ;
 wire \mandelbrot.ctr[7] ;
 wire \mandelbrot.ctr[8] ;
 wire \mandelbrot.ctr[9] ;
 wire \mandelbrot.l_alu_finished ;
 wire \mandelbrot.overflowed ;
 wire \mandelbrot.run ;
 wire \mandelbrot.running ;
 wire \mandelbrot.x[0] ;
 wire \mandelbrot.x[1] ;
 wire \mandelbrot.x[2] ;
 wire \mandelbrot.x[3] ;
 wire \mandelbrot.x[4] ;
 wire \mandelbrot.x[5] ;
 wire \mandelbrot.x[6] ;
 wire \mandelbrot.x[7] ;
 wire \mandelbrot.x[8] ;
 wire \mandelbrot.y[0] ;
 wire \mandelbrot.y[1] ;
 wire \mandelbrot.y[2] ;
 wire \mandelbrot.y[3] ;
 wire \mandelbrot.y[4] ;
 wire \mandelbrot.y[5] ;
 wire \mandelbrot.y[6] ;
 wire \mandelbrot.y[7] ;
 wire \mandelbrot.y[8] ;
 wire reset_write_ptr;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire valid_data;
 wire \vga.l_read ;
 wire \vga.pixel_buffer[0] ;
 wire \vga.pixel_buffer[1] ;
 wire \vga.pixel_buffer[2] ;
 wire \vga.pixel_buffer[3] ;
 wire \vga.pixel_ctr[0] ;
 wire \vga.pixel_ctr[10] ;
 wire \vga.pixel_ctr[1] ;
 wire \vga.pixel_ctr[2] ;
 wire \vga.pixel_ctr[3] ;
 wire \vga.pixel_ctr[4] ;
 wire \vga.pixel_ctr[5] ;
 wire \vga.pixel_ctr[6] ;
 wire \vga.pixel_ctr[7] ;
 wire \vga.pixel_ctr[8] ;
 wire \vga.pixel_ctr[9] ;
 wire \vga.read ;
 wire \vga.reset_read_ptr ;
 wire \vga.timing_v.pixel[0] ;
 wire \vga.timing_v.pixel[1] ;
 wire \vga.timing_v.pixel[2] ;
 wire \vga.timing_v.pixel[3] ;
 wire \vga.timing_v.pixel[4] ;
 wire \vga.timing_v.pixel[5] ;
 wire \vga.timing_v.pixel[6] ;
 wire \vga.timing_v.pixel[7] ;
 wire \vga.timing_v.pixel[8] ;
 wire \vga.timing_v.pixel[9] ;
 wire \vga.wrote_data ;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_leaf_0_clk_regs;
 wire clknet_leaf_1_clk_regs;
 wire clknet_leaf_2_clk_regs;
 wire clknet_leaf_3_clk_regs;
 wire clknet_leaf_4_clk_regs;
 wire clknet_leaf_5_clk_regs;
 wire clknet_leaf_6_clk_regs;
 wire clknet_leaf_7_clk_regs;
 wire clknet_leaf_8_clk_regs;
 wire clknet_leaf_9_clk_regs;
 wire clknet_leaf_10_clk_regs;
 wire clknet_leaf_11_clk_regs;
 wire clknet_leaf_12_clk_regs;
 wire clknet_leaf_13_clk_regs;
 wire clknet_leaf_14_clk_regs;
 wire clknet_leaf_15_clk_regs;
 wire clknet_leaf_16_clk_regs;
 wire clknet_leaf_17_clk_regs;
 wire clknet_leaf_18_clk_regs;
 wire clknet_leaf_19_clk_regs;
 wire clknet_leaf_20_clk_regs;
 wire clknet_leaf_21_clk_regs;
 wire clknet_leaf_22_clk_regs;
 wire clknet_leaf_23_clk_regs;
 wire clknet_leaf_24_clk_regs;
 wire clknet_leaf_25_clk_regs;
 wire clknet_leaf_26_clk_regs;
 wire clknet_leaf_27_clk_regs;
 wire clknet_leaf_28_clk_regs;
 wire clknet_leaf_29_clk_regs;
 wire clknet_leaf_30_clk_regs;
 wire clknet_leaf_31_clk_regs;
 wire clknet_leaf_32_clk_regs;
 wire clknet_leaf_33_clk_regs;
 wire clknet_leaf_34_clk_regs;
 wire clknet_leaf_35_clk_regs;
 wire clknet_leaf_36_clk_regs;
 wire clknet_leaf_37_clk_regs;
 wire clknet_leaf_38_clk_regs;
 wire clknet_leaf_39_clk_regs;
 wire clknet_leaf_40_clk_regs;
 wire clknet_leaf_41_clk_regs;
 wire clknet_leaf_42_clk_regs;
 wire clknet_0_clk_regs;
 wire clknet_3_0__leaf_clk_regs;
 wire clknet_3_1__leaf_clk_regs;
 wire clknet_3_2__leaf_clk_regs;
 wire clknet_3_3__leaf_clk_regs;
 wire clknet_3_4__leaf_clk_regs;
 wire clknet_3_5__leaf_clk_regs;
 wire clknet_3_6__leaf_clk_regs;
 wire clknet_3_7__leaf_clk_regs;
 wire delaynet_0_clk;
 wire delaynet_1_clk;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;

 sg13g2_inv_1 _2569_ (.Y(\mandelbrot.running ),
    .A(net677));
 sg13g2_inv_1 _2570_ (.Y(_1908_),
    .A(net219));
 sg13g2_inv_1 _2571_ (.Y(_1909_),
    .A(net217));
 sg13g2_inv_2 _2572_ (.Y(_1910_),
    .A(net685));
 sg13g2_inv_1 _2573_ (.Y(_1911_),
    .A(net692));
 sg13g2_inv_1 _2574_ (.Y(_1912_),
    .A(net680));
 sg13g2_inv_1 _2575_ (.Y(_1913_),
    .A(\mandelbrot.alu.mult_zr_zr.ctr[0] ));
 sg13g2_inv_1 _2576_ (.Y(_1914_),
    .A(\mandelbrot.alu.mult_zi_zi.ctr[0] ));
 sg13g2_inv_1 _2577_ (.Y(_1915_),
    .A(\mandelbrot.alu.mult_zr_zi.ctr[0] ));
 sg13g2_inv_1 _2578_ (.Y(_1916_),
    .A(\mandelbrot.ctr[0] ));
 sg13g2_inv_1 _2579_ (.Y(_1917_),
    .A(net204));
 sg13g2_inv_1 _2580_ (.Y(_1918_),
    .A(net208));
 sg13g2_inv_4 _2581_ (.A(\mandelbrot.alu.m2[27] ),
    .Y(_1919_));
 sg13g2_inv_1 _2582_ (.Y(_1920_),
    .A(\mandelbrot.alu.m1[27] ));
 sg13g2_inv_1 _2583_ (.Y(_1921_),
    .A(\mandelbrot.alu.m1[17] ));
 sg13g2_inv_1 _2584_ (.Y(_1922_),
    .A(\mandelbrot.alu.m2[16] ));
 sg13g2_inv_1 _2585_ (.Y(_1923_),
    .A(net816));
 sg13g2_inv_1 _2586_ (.Y(_1924_),
    .A(net724));
 sg13g2_inv_1 _2587_ (.Y(_1925_),
    .A(net523));
 sg13g2_inv_1 _2588_ (.Y(_1926_),
    .A(\mandelbrot.alu.m2[13] ));
 sg13g2_inv_1 _2589_ (.Y(_1927_),
    .A(net533));
 sg13g2_inv_1 _2590_ (.Y(_1928_),
    .A(\mandelbrot.alu.m2[12] ));
 sg13g2_inv_1 _2591_ (.Y(_1929_),
    .A(net470));
 sg13g2_inv_1 _2592_ (.Y(_1930_),
    .A(net750));
 sg13g2_inv_1 _2593_ (.Y(_1931_),
    .A(net513));
 sg13g2_inv_1 _2594_ (.Y(_1932_),
    .A(net738));
 sg13g2_inv_1 _2595_ (.Y(_1933_),
    .A(net499));
 sg13g2_inv_2 _2596_ (.Y(_1934_),
    .A(net703));
 sg13g2_inv_2 _2597_ (.Y(_1935_),
    .A(net669));
 sg13g2_inv_1 _2598_ (.Y(_1936_),
    .A(\configuration[42] ));
 sg13g2_inv_1 _2599_ (.Y(_1937_),
    .A(net420));
 sg13g2_inv_1 _2600_ (.Y(_1938_),
    .A(\mandelbrot.ctr[1] ));
 sg13g2_inv_1 _2601_ (.Y(_1939_),
    .A(\mandelbrot.ctr[3] ));
 sg13g2_inv_1 _2602_ (.Y(_1940_),
    .A(\mandelbrot.ctr[4] ));
 sg13g2_inv_2 _2603_ (.Y(_1941_),
    .A(\mandelbrot.ctr[6] ));
 sg13g2_inv_1 _2604_ (.Y(_1942_),
    .A(\mandelbrot.ctr[7] ));
 sg13g2_inv_2 _2605_ (.Y(_1943_),
    .A(net271));
 sg13g2_inv_1 _2606_ (.Y(_1944_),
    .A(net286));
 sg13g2_inv_1 _2607_ (.Y(_1945_),
    .A(net256));
 sg13g2_inv_1 _2608_ (.Y(_1946_),
    .A(\mandelbrot.x[0] ));
 sg13g2_inv_1 _2609_ (.Y(_1947_),
    .A(net458));
 sg13g2_inv_1 _2610_ (.Y(_1948_),
    .A(\vga.pixel_ctr[5] ));
 sg13g2_inv_1 _2611_ (.Y(_1949_),
    .A(net713));
 sg13g2_inv_1 _2612_ (.Y(_1950_),
    .A(_0053_));
 sg13g2_inv_1 _2613_ (.Y(_1951_),
    .A(\mandelbrot.alu.in_ci[12] ));
 sg13g2_inv_1 _2614_ (.Y(_1952_),
    .A(\mandelbrot.alu.m3[25] ));
 sg13g2_inv_1 _2615_ (.Y(_1953_),
    .A(\mandelbrot.alu.in_ci[9] ));
 sg13g2_inv_1 _2616_ (.Y(_1954_),
    .A(net380));
 sg13g2_inv_1 _2617_ (.Y(_1955_),
    .A(net729));
 sg13g2_inv_1 _2618_ (.Y(_1956_),
    .A(net371));
 sg13g2_inv_2 _2619_ (.Y(_1957_),
    .A(net697));
 sg13g2_inv_1 _2620_ (.Y(_1958_),
    .A(\vga.timing_v.pixel[7] ));
 sg13g2_inv_1 _2621_ (.Y(_1959_),
    .A(\vga.timing_v.pixel[5] ));
 sg13g2_inv_1 _2622_ (.Y(_1960_),
    .A(net406));
 sg13g2_inv_1 _2623_ (.Y(_1961_),
    .A(net269));
 sg13g2_inv_1 _2624_ (.Y(_1962_),
    .A(uio_out[1]));
 sg13g2_inv_1 _2625_ (.Y(_1963_),
    .A(net253));
 sg13g2_inv_1 _2626_ (.Y(_1964_),
    .A(_0027_));
 sg13g2_inv_1 _2627_ (.Y(_1965_),
    .A(_0069_));
 sg13g2_inv_1 _2628_ (.Y(_1966_),
    .A(_0059_));
 sg13g2_inv_1 _2629_ (.Y(_1967_),
    .A(_0017_));
 sg13g2_inv_1 _2630_ (.Y(_1968_),
    .A(net277));
 sg13g2_inv_1 _2631_ (.Y(_1969_),
    .A(_0047_));
 sg13g2_inv_1 _2632_ (.Y(_1970_),
    .A(net812));
 sg13g2_inv_1 _2633_ (.Y(_1971_),
    .A(net261));
 sg13g2_inv_1 _2634_ (.Y(_1972_),
    .A(net233));
 sg13g2_inv_1 _2635_ (.Y(_1973_),
    .A(net255));
 sg13g2_inv_1 _2636_ (.Y(_1974_),
    .A(net243));
 sg13g2_inv_1 _2637_ (.Y(_1975_),
    .A(\mandelbrot.alu.m3[10] ));
 sg13g2_inv_1 _2638_ (.Y(_1976_),
    .A(net300));
 sg13g2_inv_1 _2639_ (.Y(_1977_),
    .A(_0085_));
 sg13g2_inv_1 _2640_ (.Y(_1978_),
    .A(net315));
 sg13g2_inv_1 _2641_ (.Y(_1979_),
    .A(\configuration[13] ));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_xor2_1 _2643_ (.B(\mandelbrot.alu.m1[30] ),
    .A(\mandelbrot.alu.m2[30] ),
    .X(_1980_));
 sg13g2_xnor2_1 _2644_ (.Y(_1981_),
    .A(\mandelbrot.alu.m2[30] ),
    .B(\mandelbrot.alu.m1[30] ));
 sg13g2_nand2_1 _2645_ (.Y(_1982_),
    .A(\mandelbrot.alu.m2[26] ),
    .B(\mandelbrot.alu.m1[26] ));
 sg13g2_a21oi_1 _2646_ (.A1(_1919_),
    .A2(_1920_),
    .Y(_1983_),
    .B1(_1982_));
 sg13g2_xor2_1 _2647_ (.B(\mandelbrot.alu.m1[27] ),
    .A(\mandelbrot.alu.m2[27] ),
    .X(_1984_));
 sg13g2_nor2_1 _2648_ (.A(\mandelbrot.alu.m2[26] ),
    .B(\mandelbrot.alu.m1[26] ),
    .Y(_1985_));
 sg13g2_xor2_1 _2649_ (.B(\mandelbrot.alu.m1[26] ),
    .A(\mandelbrot.alu.m2[26] ),
    .X(_1986_));
 sg13g2_and2_1 _2650_ (.A(_1984_),
    .B(_1986_),
    .X(_1987_));
 sg13g2_or2_1 _2651_ (.X(_1988_),
    .B(\mandelbrot.alu.m1[23] ),
    .A(\mandelbrot.alu.m2[23] ));
 sg13g2_and3_1 _2652_ (.X(_1989_),
    .A(\mandelbrot.alu.m2[22] ),
    .B(\mandelbrot.alu.m1[22] ),
    .C(_1988_));
 sg13g2_xnor2_1 _2653_ (.Y(_1990_),
    .A(\mandelbrot.alu.m2[23] ),
    .B(\mandelbrot.alu.m1[23] ));
 sg13g2_nor2_1 _2654_ (.A(\mandelbrot.alu.m2[22] ),
    .B(\mandelbrot.alu.m1[22] ),
    .Y(_1991_));
 sg13g2_xnor2_1 _2655_ (.Y(_1992_),
    .A(\mandelbrot.alu.m2[22] ),
    .B(\mandelbrot.alu.m1[22] ));
 sg13g2_nor2_1 _2656_ (.A(_1990_),
    .B(_1992_),
    .Y(_1993_));
 sg13g2_nor2_1 _2657_ (.A(\mandelbrot.alu.m2[21] ),
    .B(\mandelbrot.alu.m1[21] ),
    .Y(_1994_));
 sg13g2_a22oi_1 _2658_ (.Y(_1995_),
    .B1(\mandelbrot.alu.m2[20] ),
    .B2(\mandelbrot.alu.m1[20] ),
    .A2(\mandelbrot.alu.m1[21] ),
    .A1(\mandelbrot.alu.m2[21] ));
 sg13g2_nor2_1 _2659_ (.A(_1994_),
    .B(_1995_),
    .Y(_1996_));
 sg13g2_nor2_1 _2660_ (.A(\mandelbrot.alu.m2[2] ),
    .B(\mandelbrot.alu.m1[2] ),
    .Y(_1997_));
 sg13g2_nor2_1 _2661_ (.A(net705),
    .B(net665),
    .Y(_1998_));
 sg13g2_a22oi_1 _2662_ (.Y(_1999_),
    .B1(\mandelbrot.alu.m2[0] ),
    .B2(\mandelbrot.alu.m1[0] ),
    .A2(net665),
    .A1(net704));
 sg13g2_or3_1 _2663_ (.A(_1997_),
    .B(_1998_),
    .C(_1999_),
    .X(_2000_));
 sg13g2_a22oi_1 _2664_ (.Y(_2001_),
    .B1(\mandelbrot.alu.m2[2] ),
    .B2(\mandelbrot.alu.m1[2] ),
    .A2(\mandelbrot.alu.m1[3] ),
    .A1(\mandelbrot.alu.m2[3] ));
 sg13g2_or2_1 _2665_ (.X(_2002_),
    .B(\mandelbrot.alu.m1[4] ),
    .A(\mandelbrot.alu.m2[4] ));
 sg13g2_o21ai_1 _2666_ (.B1(_2002_),
    .Y(_2003_),
    .A1(\mandelbrot.alu.m2[3] ),
    .A2(\mandelbrot.alu.m1[3] ));
 sg13g2_a21o_1 _2667_ (.A2(_2001_),
    .A1(_2000_),
    .B1(_2003_),
    .X(_2004_));
 sg13g2_a22oi_1 _2668_ (.Y(_2005_),
    .B1(\mandelbrot.alu.m2[4] ),
    .B2(\mandelbrot.alu.m1[4] ),
    .A2(\mandelbrot.alu.m1[5] ),
    .A1(\mandelbrot.alu.m2[5] ));
 sg13g2_nand2_1 _2669_ (.Y(_2006_),
    .A(\mandelbrot.alu.m2[7] ),
    .B(\mandelbrot.alu.m1[7] ));
 sg13g2_nor2_1 _2670_ (.A(\mandelbrot.alu.m2[7] ),
    .B(\mandelbrot.alu.m1[7] ),
    .Y(_2007_));
 sg13g2_xor2_1 _2671_ (.B(\mandelbrot.alu.m1[7] ),
    .A(\mandelbrot.alu.m2[7] ),
    .X(_2008_));
 sg13g2_nand2_1 _2672_ (.Y(_2009_),
    .A(\mandelbrot.alu.m2[6] ),
    .B(\mandelbrot.alu.m1[6] ));
 sg13g2_xor2_1 _2673_ (.B(\mandelbrot.alu.m1[6] ),
    .A(\mandelbrot.alu.m2[6] ),
    .X(_2010_));
 sg13g2_or2_1 _2674_ (.X(_2011_),
    .B(\mandelbrot.alu.m1[5] ),
    .A(\mandelbrot.alu.m2[5] ));
 sg13g2_nand3_1 _2675_ (.B(_2010_),
    .C(_2011_),
    .A(_2008_),
    .Y(_2012_));
 sg13g2_a21oi_1 _2676_ (.A1(_2004_),
    .A2(_2005_),
    .Y(_2013_),
    .B1(_2012_));
 sg13g2_o21ai_1 _2677_ (.B1(_2006_),
    .Y(_2014_),
    .A1(_2007_),
    .A2(_2009_));
 sg13g2_nand2b_1 _2678_ (.Y(_2015_),
    .B(\mandelbrot.alu.m2[11] ),
    .A_N(\mandelbrot.alu.m1[11] ));
 sg13g2_nand2b_1 _2679_ (.Y(_2016_),
    .B(\mandelbrot.alu.m1[11] ),
    .A_N(\mandelbrot.alu.m2[11] ));
 sg13g2_nand2_1 _2680_ (.Y(_2017_),
    .A(_2015_),
    .B(_2016_));
 sg13g2_xor2_1 _2681_ (.B(\mandelbrot.alu.m1[10] ),
    .A(\mandelbrot.alu.m2[10] ),
    .X(_2018_));
 sg13g2_nand2_1 _2682_ (.Y(_2019_),
    .A(_2017_),
    .B(_2018_));
 sg13g2_nor2b_1 _2683_ (.A(\mandelbrot.alu.m1[9] ),
    .B_N(\mandelbrot.alu.m2[9] ),
    .Y(_2020_));
 sg13g2_nand2b_1 _2684_ (.Y(_2021_),
    .B(\mandelbrot.alu.m1[9] ),
    .A_N(\mandelbrot.alu.m2[9] ));
 sg13g2_nor2b_1 _2685_ (.A(_2020_),
    .B_N(_2021_),
    .Y(_2022_));
 sg13g2_nand2b_1 _2686_ (.Y(_2023_),
    .B(\mandelbrot.alu.m1[8] ),
    .A_N(\mandelbrot.alu.m2[8] ));
 sg13g2_xnor2_1 _2687_ (.Y(_2024_),
    .A(\mandelbrot.alu.m2[8] ),
    .B(\mandelbrot.alu.m1[8] ));
 sg13g2_nor3_1 _2688_ (.A(_2019_),
    .B(_2022_),
    .C(_2024_),
    .Y(_2025_));
 sg13g2_o21ai_1 _2689_ (.B1(_2025_),
    .Y(_2026_),
    .A1(_2013_),
    .A2(_2014_));
 sg13g2_nand3b_1 _2690_ (.B(\mandelbrot.alu.m1[8] ),
    .C(\mandelbrot.alu.m2[8] ),
    .Y(_2027_),
    .A_N(_2022_));
 sg13g2_a22oi_1 _2691_ (.Y(_2028_),
    .B1(\mandelbrot.alu.m2[9] ),
    .B2(\mandelbrot.alu.m1[9] ),
    .A2(\mandelbrot.alu.m1[10] ),
    .A1(\mandelbrot.alu.m2[10] ));
 sg13g2_o21ai_1 _2692_ (.B1(_2017_),
    .Y(_2029_),
    .A1(\mandelbrot.alu.m2[10] ),
    .A2(\mandelbrot.alu.m1[10] ));
 sg13g2_a21oi_1 _2693_ (.A1(_2027_),
    .A2(_2028_),
    .Y(_2030_),
    .B1(_2029_));
 sg13g2_a21oi_1 _2694_ (.A1(\mandelbrot.alu.m2[11] ),
    .A2(\mandelbrot.alu.m1[11] ),
    .Y(_2031_),
    .B1(_2030_));
 sg13g2_xor2_1 _2695_ (.B(\mandelbrot.alu.m1[13] ),
    .A(\mandelbrot.alu.m2[13] ),
    .X(_2032_));
 sg13g2_xor2_1 _2696_ (.B(\mandelbrot.alu.m1[12] ),
    .A(\mandelbrot.alu.m2[12] ),
    .X(_2033_));
 sg13g2_nand2_1 _2697_ (.Y(_2034_),
    .A(_2032_),
    .B(_2033_));
 sg13g2_a21oi_1 _2698_ (.A1(_2026_),
    .A2(_2031_),
    .Y(_2035_),
    .B1(_2034_));
 sg13g2_nand3_1 _2699_ (.B(\mandelbrot.alu.m1[12] ),
    .C(_2032_),
    .A(\mandelbrot.alu.m2[12] ),
    .Y(_2036_));
 sg13g2_o21ai_1 _2700_ (.B1(_2036_),
    .Y(_2037_),
    .A1(_1926_),
    .A2(_1927_));
 sg13g2_nor2_1 _2701_ (.A(_2035_),
    .B(_2037_),
    .Y(_2038_));
 sg13g2_nor2_1 _2702_ (.A(\mandelbrot.alu.m2[14] ),
    .B(\mandelbrot.alu.m1[14] ),
    .Y(_2039_));
 sg13g2_xor2_1 _2703_ (.B(\mandelbrot.alu.m1[14] ),
    .A(\mandelbrot.alu.m2[14] ),
    .X(_2040_));
 sg13g2_o21ai_1 _2704_ (.B1(_2040_),
    .Y(_2041_),
    .A1(_2035_),
    .A2(_2037_));
 sg13g2_a22oi_1 _2705_ (.Y(_2042_),
    .B1(\mandelbrot.alu.m2[14] ),
    .B2(\mandelbrot.alu.m1[14] ),
    .A2(\mandelbrot.alu.m1[15] ),
    .A1(\mandelbrot.alu.m2[15] ));
 sg13g2_a22oi_1 _2706_ (.Y(_2043_),
    .B1(_2041_),
    .B2(_2042_),
    .A2(_1924_),
    .A1(_1923_));
 sg13g2_nor2_1 _2707_ (.A(\mandelbrot.alu.m2[17] ),
    .B(\mandelbrot.alu.m1[17] ),
    .Y(_2044_));
 sg13g2_nand2_1 _2708_ (.Y(_2045_),
    .A(\mandelbrot.alu.m2[17] ),
    .B(\mandelbrot.alu.m1[17] ));
 sg13g2_nand2b_2 _2709_ (.Y(_2046_),
    .B(_2045_),
    .A_N(_2044_));
 sg13g2_nand2_1 _2710_ (.Y(_2047_),
    .A(\mandelbrot.alu.m2[16] ),
    .B(\mandelbrot.alu.m1[16] ));
 sg13g2_nor2_1 _2711_ (.A(\mandelbrot.alu.m2[16] ),
    .B(\mandelbrot.alu.m1[16] ),
    .Y(_2048_));
 sg13g2_xor2_1 _2712_ (.B(\mandelbrot.alu.m1[16] ),
    .A(\mandelbrot.alu.m2[16] ),
    .X(_2049_));
 sg13g2_xnor2_1 _2713_ (.Y(_2050_),
    .A(\mandelbrot.alu.m2[16] ),
    .B(\mandelbrot.alu.m1[16] ));
 sg13g2_nand2b_1 _2714_ (.Y(_2051_),
    .B(_2049_),
    .A_N(_2046_));
 sg13g2_a221oi_1 _2715_ (.B2(_2042_),
    .C1(_2051_),
    .B1(_2041_),
    .A1(_1923_),
    .Y(_2052_),
    .A2(_1924_));
 sg13g2_o21ai_1 _2716_ (.B1(_2045_),
    .Y(_2053_),
    .A1(_2044_),
    .A2(_2047_));
 sg13g2_nor2_1 _2717_ (.A(_2052_),
    .B(_2053_),
    .Y(_2054_));
 sg13g2_nand2_1 _2718_ (.Y(_2055_),
    .A(\mandelbrot.alu.m2[19] ),
    .B(\mandelbrot.alu.m1[19] ));
 sg13g2_nor2_1 _2719_ (.A(\mandelbrot.alu.m2[19] ),
    .B(\mandelbrot.alu.m1[19] ),
    .Y(_2056_));
 sg13g2_nand2_1 _2720_ (.Y(_2057_),
    .A(\mandelbrot.alu.m2[18] ),
    .B(\mandelbrot.alu.m1[18] ));
 sg13g2_o21ai_1 _2721_ (.B1(_2055_),
    .Y(_2058_),
    .A1(_2056_),
    .A2(_2057_));
 sg13g2_nor3_2 _2722_ (.A(_2052_),
    .B(_2053_),
    .C(_2058_),
    .Y(_2059_));
 sg13g2_nor2_1 _2723_ (.A(\mandelbrot.alu.m2[18] ),
    .B(\mandelbrot.alu.m1[18] ),
    .Y(_2060_));
 sg13g2_a21o_2 _2724_ (.A2(_2060_),
    .A1(_2055_),
    .B1(_2056_),
    .X(_2061_));
 sg13g2_xnor2_1 _2725_ (.Y(_2062_),
    .A(\mandelbrot.alu.m2[21] ),
    .B(\mandelbrot.alu.m1[21] ));
 sg13g2_nor2_1 _2726_ (.A(\mandelbrot.alu.m2[20] ),
    .B(\mandelbrot.alu.m1[20] ),
    .Y(_2063_));
 sg13g2_xnor2_1 _2727_ (.Y(_2064_),
    .A(\mandelbrot.alu.m2[20] ),
    .B(\mandelbrot.alu.m1[20] ));
 sg13g2_inv_1 _2728_ (.Y(_2065_),
    .A(_2064_));
 sg13g2_nor4_2 _2729_ (.A(_2059_),
    .B(_2061_),
    .C(_2062_),
    .Y(_2066_),
    .D(_2064_));
 sg13g2_or4_1 _2730_ (.A(_1990_),
    .B(_1992_),
    .C(_2062_),
    .D(_2064_),
    .X(_2067_));
 sg13g2_or3_2 _2731_ (.A(_2059_),
    .B(_2061_),
    .C(_2067_),
    .X(_2068_));
 sg13g2_a221oi_1 _2732_ (.B2(_1996_),
    .C1(_1989_),
    .B1(_1993_),
    .A1(\mandelbrot.alu.m2[23] ),
    .Y(_2069_),
    .A2(\mandelbrot.alu.m1[23] ));
 sg13g2_xor2_1 _2733_ (.B(\mandelbrot.alu.m1[25] ),
    .A(\mandelbrot.alu.m2[25] ),
    .X(_2070_));
 sg13g2_xnor2_1 _2734_ (.Y(_2071_),
    .A(net700),
    .B(\mandelbrot.alu.m1[25] ));
 sg13g2_nor2_1 _2735_ (.A(\mandelbrot.alu.m2[24] ),
    .B(\mandelbrot.alu.m1[24] ),
    .Y(_2072_));
 sg13g2_xor2_1 _2736_ (.B(\mandelbrot.alu.m1[24] ),
    .A(\mandelbrot.alu.m2[24] ),
    .X(_2073_));
 sg13g2_nand2_1 _2737_ (.Y(_2074_),
    .A(_2070_),
    .B(_2073_));
 sg13g2_a21o_1 _2738_ (.A2(_2069_),
    .A1(_2068_),
    .B1(_2074_),
    .X(_2075_));
 sg13g2_a22oi_1 _2739_ (.Y(_2076_),
    .B1(\mandelbrot.alu.m2[24] ),
    .B2(\mandelbrot.alu.m1[24] ),
    .A2(\mandelbrot.alu.m1[25] ),
    .A1(net700));
 sg13g2_inv_1 _2740_ (.Y(_2077_),
    .A(_2076_));
 sg13g2_o21ai_1 _2741_ (.B1(_2077_),
    .Y(_2078_),
    .A1(net700),
    .A2(\mandelbrot.alu.m1[25] ));
 sg13g2_inv_1 _2742_ (.Y(_2079_),
    .A(_2078_));
 sg13g2_nand3_1 _2743_ (.B(_2070_),
    .C(_2073_),
    .A(_1987_),
    .Y(_2080_));
 sg13g2_a21o_1 _2744_ (.A2(_2069_),
    .A1(_2068_),
    .B1(_2080_),
    .X(_2081_));
 sg13g2_a221oi_1 _2745_ (.B2(_2079_),
    .C1(_1983_),
    .B1(_1987_),
    .A1(\mandelbrot.alu.m2[27] ),
    .Y(_2082_),
    .A2(\mandelbrot.alu.m1[27] ));
 sg13g2_nand2_1 _2746_ (.Y(_2083_),
    .A(_2081_),
    .B(_2082_));
 sg13g2_xor2_1 _2747_ (.B(\mandelbrot.alu.m1[29] ),
    .A(\mandelbrot.alu.m2[29] ),
    .X(_2084_));
 sg13g2_nor2_1 _2748_ (.A(\mandelbrot.alu.m2[28] ),
    .B(\mandelbrot.alu.m1[28] ),
    .Y(_2085_));
 sg13g2_xor2_1 _2749_ (.B(\mandelbrot.alu.m1[28] ),
    .A(\mandelbrot.alu.m2[28] ),
    .X(_2086_));
 sg13g2_nand2_1 _2750_ (.Y(_2087_),
    .A(_2084_),
    .B(_2086_));
 sg13g2_a21oi_2 _2751_ (.B1(_2087_),
    .Y(_2088_),
    .A2(_2082_),
    .A1(_2081_));
 sg13g2_a22oi_1 _2752_ (.Y(_2089_),
    .B1(\mandelbrot.alu.m2[28] ),
    .B2(\mandelbrot.alu.m1[28] ),
    .A2(\mandelbrot.alu.m1[29] ),
    .A1(\mandelbrot.alu.m2[29] ));
 sg13g2_inv_1 _2753_ (.Y(_2090_),
    .A(_2089_));
 sg13g2_o21ai_1 _2754_ (.B1(_2090_),
    .Y(_2091_),
    .A1(\mandelbrot.alu.m2[29] ),
    .A2(\mandelbrot.alu.m1[29] ));
 sg13g2_inv_1 _2755_ (.Y(_2092_),
    .A(_2091_));
 sg13g2_nor2_1 _2756_ (.A(_2088_),
    .B(_2092_),
    .Y(_2093_));
 sg13g2_xnor2_1 _2757_ (.Y(_2094_),
    .A(_2083_),
    .B(_2086_));
 sg13g2_a21oi_1 _2758_ (.A1(_2075_),
    .A2(_2078_),
    .Y(_2095_),
    .B1(_1986_));
 sg13g2_and3_1 _2759_ (.X(_2096_),
    .A(_1986_),
    .B(_2075_),
    .C(_2078_));
 sg13g2_a21oi_1 _2760_ (.A1(_2068_),
    .A2(_2069_),
    .Y(_2097_),
    .B1(_2073_));
 sg13g2_nand3_1 _2761_ (.B(_2069_),
    .C(_2073_),
    .A(_2068_),
    .Y(_2098_));
 sg13g2_o21ai_1 _2762_ (.B1(_1992_),
    .Y(_2099_),
    .A1(_1996_),
    .A2(_2066_));
 sg13g2_o21ai_1 _2763_ (.B1(_2065_),
    .Y(_2100_),
    .A1(_2059_),
    .A2(_2061_));
 sg13g2_xor2_1 _2764_ (.B(\mandelbrot.alu.m1[18] ),
    .A(\mandelbrot.alu.m2[18] ),
    .X(_2101_));
 sg13g2_xnor2_1 _2765_ (.Y(_2102_),
    .A(\mandelbrot.alu.m2[18] ),
    .B(\mandelbrot.alu.m1[18] ));
 sg13g2_xnor2_1 _2766_ (.Y(_2103_),
    .A(_2038_),
    .B(_2040_));
 sg13g2_xnor2_1 _2767_ (.Y(_2104_),
    .A(_2071_),
    .B(_2072_));
 sg13g2_xor2_1 _2768_ (.B(_1985_),
    .A(_1984_),
    .X(_2105_));
 sg13g2_xnor2_1 _2769_ (.Y(_2106_),
    .A(_2046_),
    .B(_2048_));
 sg13g2_xnor2_1 _2770_ (.Y(_2107_),
    .A(\mandelbrot.alu.m2[19] ),
    .B(\mandelbrot.alu.m1[19] ));
 sg13g2_xnor2_1 _2771_ (.Y(_2108_),
    .A(_2060_),
    .B(_2107_));
 sg13g2_xor2_1 _2772_ (.B(\mandelbrot.alu.m1[15] ),
    .A(\mandelbrot.alu.m2[15] ),
    .X(_2109_));
 sg13g2_xor2_1 _2773_ (.B(_2109_),
    .A(_2039_),
    .X(_2110_));
 sg13g2_xnor2_1 _2774_ (.Y(_2111_),
    .A(_2062_),
    .B(_2063_));
 sg13g2_xor2_1 _2775_ (.B(_2085_),
    .A(_2084_),
    .X(_2112_));
 sg13g2_xnor2_1 _2776_ (.Y(_2113_),
    .A(_1990_),
    .B(_1991_));
 sg13g2_nand4_1 _2777_ (.B(_2105_),
    .C(_2106_),
    .A(_2104_),
    .Y(_2114_),
    .D(_2112_));
 sg13g2_nand4_1 _2778_ (.B(_2110_),
    .C(_2111_),
    .A(_2108_),
    .Y(_2115_),
    .D(_2113_));
 sg13g2_xnor2_1 _2779_ (.Y(_2116_),
    .A(_2043_),
    .B(_2050_));
 sg13g2_nor4_1 _2780_ (.A(_2103_),
    .B(_2114_),
    .C(_2115_),
    .D(_2116_),
    .Y(_2117_));
 sg13g2_xnor2_1 _2781_ (.Y(_2118_),
    .A(_2054_),
    .B(_2102_));
 sg13g2_or3_1 _2782_ (.A(_2059_),
    .B(_2061_),
    .C(_2065_),
    .X(_2119_));
 sg13g2_and4_1 _2783_ (.A(_2100_),
    .B(_2117_),
    .C(_2118_),
    .D(_2119_),
    .X(_2120_));
 sg13g2_or3_1 _2784_ (.A(_1992_),
    .B(_1996_),
    .C(_2066_),
    .X(_2121_));
 sg13g2_nand4_1 _2785_ (.B(_2099_),
    .C(_2120_),
    .A(_2098_),
    .Y(_2122_),
    .D(_2121_));
 sg13g2_nor4_2 _2786_ (.A(_2095_),
    .B(_2096_),
    .C(_2097_),
    .Y(_2123_),
    .D(_2122_));
 sg13g2_a22oi_1 _2787_ (.Y(_2124_),
    .B1(_2094_),
    .B2(_2123_),
    .A2(_2093_),
    .A1(_1981_));
 sg13g2_xor2_1 _2788_ (.B(\mandelbrot.alu.m1[31] ),
    .A(\mandelbrot.alu.m2[31] ),
    .X(_2125_));
 sg13g2_xnor2_1 _2789_ (.Y(_2126_),
    .A(\mandelbrot.alu.m2[31] ),
    .B(\mandelbrot.alu.m1[31] ));
 sg13g2_and3_1 _2790_ (.X(_2127_),
    .A(\mandelbrot.alu.m2[30] ),
    .B(\mandelbrot.alu.m1[30] ),
    .C(_2125_));
 sg13g2_o21ai_1 _2791_ (.B1(_1980_),
    .Y(_2128_),
    .A1(_2088_),
    .A2(_2092_));
 sg13g2_a21oi_1 _2792_ (.A1(\mandelbrot.alu.m2[30] ),
    .A2(\mandelbrot.alu.m1[30] ),
    .Y(_2129_),
    .B1(_2125_));
 sg13g2_a21oi_1 _2793_ (.A1(_2128_),
    .A2(_2129_),
    .Y(_2130_),
    .B1(_2127_));
 sg13g2_or2_1 _2794_ (.X(_2131_),
    .B(_2128_),
    .A(_2126_));
 sg13g2_o21ai_1 _2795_ (.B1(_2131_),
    .Y(_2132_),
    .A1(_2124_),
    .A2(_2130_));
 sg13g2_nor2_1 _2796_ (.A(_1981_),
    .B(_2126_),
    .Y(_2133_));
 sg13g2_a21oi_1 _2797_ (.A1(\mandelbrot.alu.m2[31] ),
    .A2(\mandelbrot.alu.m1[31] ),
    .Y(_2134_),
    .B1(\mandelbrot.overflowed ));
 sg13g2_a21oi_1 _2798_ (.A1(_2092_),
    .A2(_2133_),
    .Y(_2135_),
    .B1(_2127_));
 sg13g2_nor2_1 _2799_ (.A(_1944_),
    .B(\mandelbrot.ctr[9] ),
    .Y(_2136_));
 sg13g2_a22oi_1 _2800_ (.Y(_2137_),
    .B1(_1944_),
    .B2(\mandelbrot.ctr[9] ),
    .A2(\mandelbrot.ctr[1] ),
    .A1(_1937_));
 sg13g2_nor2_1 _2801_ (.A(_1943_),
    .B(\mandelbrot.ctr[8] ),
    .Y(_2138_));
 sg13g2_nand2b_1 _2802_ (.Y(_2139_),
    .B(\mandelbrot.ctr[7] ),
    .A_N(\configuration[49] ));
 sg13g2_a22oi_1 _2803_ (.Y(_2140_),
    .B1(\configuration[48] ),
    .B2(_1941_),
    .A2(\configuration[42] ),
    .A1(_1916_));
 sg13g2_o21ai_1 _2804_ (.B1(_2139_),
    .Y(_2141_),
    .A1(\configuration[48] ),
    .A2(_1941_));
 sg13g2_nand2_1 _2805_ (.Y(_2142_),
    .A(\configuration[47] ),
    .B(net672));
 sg13g2_or2_1 _2806_ (.X(_2143_),
    .B(net672),
    .A(\configuration[47] ));
 sg13g2_a221oi_1 _2807_ (.B2(_2143_),
    .C1(_2141_),
    .B1(_2142_),
    .A1(\configuration[49] ),
    .Y(_2144_),
    .A2(_1942_));
 sg13g2_a22oi_1 _2808_ (.Y(_2145_),
    .B1(\configuration[43] ),
    .B2(_1938_),
    .A2(_1936_),
    .A1(\mandelbrot.ctr[0] ));
 sg13g2_xnor2_1 _2809_ (.Y(_2146_),
    .A(\configuration[44] ),
    .B(\mandelbrot.ctr[2] ));
 sg13g2_a22oi_1 _2810_ (.Y(_2147_),
    .B1(_1943_),
    .B2(\mandelbrot.ctr[8] ),
    .A2(_1940_),
    .A1(\configuration[46] ));
 sg13g2_xnor2_1 _2811_ (.Y(_2148_),
    .A(\configuration[45] ),
    .B(\mandelbrot.ctr[3] ));
 sg13g2_nand4_1 _2812_ (.B(_2146_),
    .C(_2147_),
    .A(_2145_),
    .Y(_2149_),
    .D(_2148_));
 sg13g2_nor2_1 _2813_ (.A(\configuration[46] ),
    .B(_1940_),
    .Y(_2150_));
 sg13g2_nor4_1 _2814_ (.A(_2136_),
    .B(_2138_),
    .C(_2149_),
    .D(_2150_),
    .Y(_2151_));
 sg13g2_nand4_1 _2815_ (.B(_2140_),
    .C(_2144_),
    .A(_2137_),
    .Y(_2152_),
    .D(_2151_));
 sg13g2_nand3_1 _2816_ (.B(_2135_),
    .C(_2152_),
    .A(_2134_),
    .Y(_2153_));
 sg13g2_a21oi_1 _2817_ (.A1(_2088_),
    .A2(_2133_),
    .Y(_2154_),
    .B1(_2153_));
 sg13g2_nor2_2 _2818_ (.A(net691),
    .B(\mandelbrot.l_alu_finished ),
    .Y(_2155_));
 sg13g2_nand2_1 _2819_ (.Y(_2156_),
    .A(net662),
    .B(_2155_));
 sg13g2_a21oi_2 _2820_ (.B1(_2156_),
    .Y(_2157_),
    .A2(_2154_),
    .A1(_2132_));
 sg13g2_a21oi_1 _2821_ (.A1(net677),
    .A2(net199),
    .Y(_0116_),
    .B1(_2157_));
 sg13g2_nand2b_1 _2822_ (.Y(_2158_),
    .B(\l_sen[2] ),
    .A_N(net202));
 sg13g2_nand2_1 _2823_ (.Y(_2159_),
    .A(net677),
    .B(net275));
 sg13g2_inv_1 _2824_ (.Y(valid_data),
    .A(_2159_));
 sg13g2_and2_1 _2825_ (.A(net282),
    .B(valid_data),
    .X(_2160_));
 sg13g2_a22oi_1 _2826_ (.Y(_0115_),
    .B1(_2160_),
    .B2(net208),
    .A2(_2158_),
    .A1(net204));
 sg13g2_nand2_2 _2827_ (.Y(_2161_),
    .A(net1),
    .B(latched_rst_n));
 sg13g2_inv_1 _2828_ (.Y(combined_rst_n),
    .A(_2161_));
 sg13g2_nor2b_1 _2829_ (.A(net292),
    .B_N(net313),
    .Y(_2162_));
 sg13g2_a21o_1 _2830_ (.A2(_2160_),
    .A1(_1918_),
    .B1(_2162_),
    .X(_0001_));
 sg13g2_a21o_1 _2831_ (.A2(net292),
    .A1(\state[1] ),
    .B1(net201),
    .X(_2568_));
 sg13g2_a21o_1 _2832_ (.A2(_2159_),
    .A1(net282),
    .B1(_2568_),
    .X(_0002_));
 sg13g2_nor3_1 _2833_ (.A(\vga.timing_v.pixel[9] ),
    .B(\vga.timing_v.pixel[8] ),
    .C(\vga.timing_v.pixel[6] ),
    .Y(_2163_));
 sg13g2_nand3_1 _2834_ (.B(_1959_),
    .C(_2163_),
    .A(_1958_),
    .Y(_2164_));
 sg13g2_nor2_1 _2835_ (.A(\vga.timing_v.pixel[1] ),
    .B(\vga.timing_v.pixel[0] ),
    .Y(_2165_));
 sg13g2_nand2b_1 _2836_ (.Y(_2166_),
    .B(_0103_),
    .A_N(\vga.timing_v.pixel[2] ));
 sg13g2_nor2_1 _2837_ (.A(\vga.timing_v.pixel[2] ),
    .B(_2165_),
    .Y(_2167_));
 sg13g2_a21oi_1 _2838_ (.A1(_2165_),
    .A2(_2166_),
    .Y(_2168_),
    .B1(_2167_));
 sg13g2_nor4_2 _2839_ (.A(\vga.timing_v.pixel[4] ),
    .B(\vga.timing_v.pixel[3] ),
    .C(_2164_),
    .Y(\vga.reset_read_ptr ),
    .D(_2168_));
 sg13g2_nor2_2 _2840_ (.A(net782),
    .B(net512),
    .Y(_2169_));
 sg13g2_nor3_2 _2841_ (.A(\vga.pixel_ctr[2] ),
    .B(\vga.pixel_ctr[1] ),
    .C(\vga.pixel_ctr[0] ),
    .Y(_2170_));
 sg13g2_nor2_1 _2842_ (.A(\vga.pixel_ctr[6] ),
    .B(\vga.pixel_ctr[7] ),
    .Y(_2171_));
 sg13g2_nor2_1 _2843_ (.A(\vga.pixel_ctr[4] ),
    .B(\vga.pixel_ctr[5] ),
    .Y(_2172_));
 sg13g2_nor4_1 _2844_ (.A(\vga.pixel_ctr[3] ),
    .B(\vga.pixel_ctr[9] ),
    .C(\vga.pixel_ctr[10] ),
    .D(_0110_),
    .Y(_2173_));
 sg13g2_and4_1 _2845_ (.A(_2170_),
    .B(_2171_),
    .C(_2172_),
    .D(_2173_),
    .X(_2174_));
 sg13g2_and2_1 _2846_ (.A(\vga.timing_v.pixel[4] ),
    .B(\vga.timing_v.pixel[3] ),
    .X(_2175_));
 sg13g2_a21oi_2 _2847_ (.B1(_2164_),
    .Y(_2176_),
    .A2(_2175_),
    .A1(\vga.timing_v.pixel[2] ));
 sg13g2_nor2_1 _2848_ (.A(\vga.pixel_ctr[9] ),
    .B(\vga.pixel_ctr[8] ),
    .Y(_2177_));
 sg13g2_nor3_1 _2849_ (.A(\vga.pixel_ctr[9] ),
    .B(\vga.pixel_ctr[8] ),
    .C(\vga.pixel_ctr[10] ),
    .Y(_2178_));
 sg13g2_nor3_2 _2850_ (.A(_2174_),
    .B(_2176_),
    .C(_2178_),
    .Y(_2179_));
 sg13g2_nand2_1 _2851_ (.Y(_2180_),
    .A(\vga.pixel_buffer[2] ),
    .B(_2179_));
 sg13g2_nand2_1 _2852_ (.Y(_2181_),
    .A(\vga.pixel_buffer[3] ),
    .B(_2179_));
 sg13g2_nand2_1 _2853_ (.Y(_0390_),
    .A(\vga.pixel_buffer[0] ),
    .B(_2179_));
 sg13g2_nand2_2 _2854_ (.Y(_0391_),
    .A(\vga.pixel_buffer[1] ),
    .B(_2179_));
 sg13g2_inv_1 _2855_ (.Y(_0392_),
    .A(_0391_));
 sg13g2_nand2_1 _2856_ (.Y(_0393_),
    .A(\vga.pixel_buffer[0] ),
    .B(_0392_));
 sg13g2_and2_1 _2857_ (.A(net583),
    .B(_0393_),
    .X(_0394_));
 sg13g2_nor2_1 _2858_ (.A(net664),
    .B(net583),
    .Y(_0395_));
 sg13g2_mux2_1 _2859_ (.A0(_0395_),
    .A1(net583),
    .S(_0393_),
    .X(_0396_));
 sg13g2_nor4_1 _2860_ (.A(\vga.pixel_buffer[1] ),
    .B(net664),
    .C(net584),
    .D(_2181_),
    .Y(_0397_));
 sg13g2_a221oi_1 _2861_ (.B2(net584),
    .C1(_0397_),
    .B1(_0396_),
    .A1(net664),
    .Y(_0398_),
    .A2(net583));
 sg13g2_mux2_2 _2862_ (.A0(_0398_),
    .A1(uio_out[0]),
    .S(net5),
    .X(uo_out[0]));
 sg13g2_nand2_1 _2863_ (.Y(_0399_),
    .A(_0390_),
    .B(_0391_));
 sg13g2_a21oi_1 _2864_ (.A1(_1961_),
    .A2(_0399_),
    .Y(_0400_),
    .B1(_2180_));
 sg13g2_nor3_1 _2865_ (.A(net5),
    .B(_0395_),
    .C(_0400_),
    .Y(_0401_));
 sg13g2_a21oi_2 _2866_ (.B1(_0401_),
    .Y(uo_out[1]),
    .A2(_1962_),
    .A1(net707));
 sg13g2_nand3_1 _2867_ (.B(net583),
    .C(_0399_),
    .A(net584),
    .Y(_0402_));
 sg13g2_a21oi_1 _2868_ (.A1(_1960_),
    .A2(_0392_),
    .Y(_0403_),
    .B1(net584));
 sg13g2_nor2_1 _2869_ (.A(net664),
    .B(_0403_),
    .Y(_0404_));
 sg13g2_a221oi_1 _2870_ (.B2(_0404_),
    .C1(net707),
    .B1(_0402_),
    .A1(net664),
    .Y(_0405_),
    .A2(_0391_));
 sg13g2_a21o_2 _2871_ (.A2(uio_out[2]),
    .A1(net707),
    .B1(_0405_),
    .X(uo_out[2]));
 sg13g2_mux2_2 _2872_ (.A0(\vga.reset_read_ptr ),
    .A1(uio_out[3]),
    .S(net707),
    .X(uo_out[3]));
 sg13g2_nor3_1 _2873_ (.A(\vga.pixel_buffer[3] ),
    .B(\vga.pixel_buffer[0] ),
    .C(_0391_),
    .Y(_0406_));
 sg13g2_nand2_1 _2874_ (.Y(_0407_),
    .A(\vga.pixel_buffer[1] ),
    .B(net584));
 sg13g2_o21ai_1 _2875_ (.B1(net584),
    .Y(_0408_),
    .A1(\vga.pixel_buffer[1] ),
    .A2(net583));
 sg13g2_nor3_1 _2876_ (.A(net664),
    .B(_0406_),
    .C(_0408_),
    .Y(_0409_));
 sg13g2_a21oi_1 _2877_ (.A1(net664),
    .A2(_0390_),
    .Y(_0410_),
    .B1(_0409_));
 sg13g2_mux2_2 _2878_ (.A0(_0410_),
    .A1(net663),
    .S(net707),
    .X(uo_out[4]));
 sg13g2_nand2b_1 _2879_ (.Y(_0411_),
    .B(_0399_),
    .A_N(net583));
 sg13g2_a21oi_1 _2880_ (.A1(net584),
    .A2(_0411_),
    .Y(_0412_),
    .B1(_0394_));
 sg13g2_mux2_1 _2881_ (.A0(_0412_),
    .A1(finished),
    .S(net707),
    .X(uo_out[5]));
 sg13g2_xnor2_1 _2882_ (.Y(_0413_),
    .A(\vga.pixel_buffer[0] ),
    .B(_0407_));
 sg13g2_nor2_1 _2883_ (.A(net583),
    .B(_0413_),
    .Y(_0414_));
 sg13g2_nor3_1 _2884_ (.A(\vga.pixel_buffer[0] ),
    .B(\vga.pixel_buffer[1] ),
    .C(net584),
    .Y(_0415_));
 sg13g2_o21ai_1 _2885_ (.B1(_0394_),
    .Y(_0416_),
    .A1(\vga.pixel_buffer[2] ),
    .A2(_0391_));
 sg13g2_nor2_1 _2886_ (.A(_0415_),
    .B(_0416_),
    .Y(_0417_));
 sg13g2_nor3_2 _2887_ (.A(net707),
    .B(_0414_),
    .C(_0417_),
    .Y(uo_out[6]));
 sg13g2_nor2_1 _2888_ (.A(\vga.pixel_ctr[4] ),
    .B(_1948_),
    .Y(_0418_));
 sg13g2_nand2b_1 _2889_ (.Y(_0419_),
    .B(\vga.pixel_ctr[3] ),
    .A_N(_2170_));
 sg13g2_a21o_1 _2890_ (.A2(_0419_),
    .A1(_0418_),
    .B1(_0107_),
    .X(_0420_));
 sg13g2_nand3_1 _2891_ (.B(_2170_),
    .C(_0418_),
    .A(\vga.pixel_ctr[3] ),
    .Y(_0421_));
 sg13g2_nand3b_1 _2892_ (.B(_0420_),
    .C(_0421_),
    .Y(_0422_),
    .A_N(\vga.pixel_ctr[6] ));
 sg13g2_nand4_1 _2893_ (.B(_2171_),
    .C(_0420_),
    .A(_0110_),
    .Y(_0423_),
    .D(_0421_));
 sg13g2_nand3b_1 _2894_ (.B(_2178_),
    .C(_0423_),
    .Y(_0424_),
    .A_N(net707));
 sg13g2_a21oi_2 _2895_ (.B1(_0424_),
    .Y(uo_out[7]),
    .A2(_0422_),
    .A1(\vga.pixel_ctr[7] ));
 sg13g2_and3_2 _2896_ (.X(_0425_),
    .A(net662),
    .B(_2132_),
    .C(_2154_));
 sg13g2_mux2_1 _2897_ (.A0(net805),
    .A1(_2155_),
    .S(_0425_),
    .X(_0426_));
 sg13g2_and2_1 _2898_ (.A(net657),
    .B(net580),
    .X(_0427_));
 sg13g2_nand2_1 _2899_ (.Y(_0428_),
    .A(net658),
    .B(_0426_));
 sg13g2_nand2_1 _2900_ (.Y(_0429_),
    .A(\mandelbrot.alu.mult_zr_zr.ctr[0] ),
    .B(net240));
 sg13g2_nand2_1 _2901_ (.Y(_0430_),
    .A(net691),
    .B(_0429_));
 sg13g2_o21ai_1 _2902_ (.B1(net691),
    .Y(_0431_),
    .A1(_1963_),
    .A2(_0429_));
 sg13g2_nand2_1 _2903_ (.Y(_0005_),
    .A(_0428_),
    .B(_0431_));
 sg13g2_nand2_1 _2904_ (.Y(_0432_),
    .A(_1910_),
    .B(net580));
 sg13g2_nand2_1 _2905_ (.Y(_0433_),
    .A(\mandelbrot.alu.mult_zi_zi.ctr[0] ),
    .B(net235));
 sg13g2_nand2_1 _2906_ (.Y(_0434_),
    .A(net688),
    .B(_0433_));
 sg13g2_o21ai_1 _2907_ (.B1(net688),
    .Y(_0435_),
    .A1(_1968_),
    .A2(_0433_));
 sg13g2_nand2_1 _2908_ (.Y(_0003_),
    .A(_0432_),
    .B(_0435_));
 sg13g2_and2_1 _2909_ (.A(net655),
    .B(net580),
    .X(_0436_));
 sg13g2_nand2_1 _2910_ (.Y(_0437_),
    .A(net656),
    .B(net580));
 sg13g2_nand2_1 _2911_ (.Y(_0438_),
    .A(net784),
    .B(net227));
 sg13g2_nand2_1 _2912_ (.Y(_0439_),
    .A(net682),
    .B(_0438_));
 sg13g2_o21ai_1 _2913_ (.B1(net682),
    .Y(_0440_),
    .A1(_1971_),
    .A2(_0438_));
 sg13g2_nand2_1 _2914_ (.Y(_0004_),
    .A(net564),
    .B(_0440_));
 sg13g2_and2_1 _2915_ (.A(net782),
    .B(\vga.pixel_ctr[0] ),
    .X(_0441_));
 sg13g2_nand3_1 _2916_ (.B(\vga.pixel_ctr[2] ),
    .C(\vga.pixel_ctr[3] ),
    .A(\vga.pixel_ctr[4] ),
    .Y(_0442_));
 sg13g2_and3_1 _2917_ (.X(_0443_),
    .A(\vga.pixel_ctr[2] ),
    .B(net447),
    .C(_0441_));
 sg13g2_and2_2 _2918_ (.A(net506),
    .B(_0443_),
    .X(_0444_));
 sg13g2_nand3_1 _2919_ (.B(_2171_),
    .C(_2177_),
    .A(_0107_),
    .Y(_0445_));
 sg13g2_a21oi_1 _2920_ (.A1(_1948_),
    .A2(_0444_),
    .Y(_0446_),
    .B1(_0445_));
 sg13g2_nor2b_1 _2921_ (.A(_0446_),
    .B_N(net828),
    .Y(_0447_));
 sg13g2_nand2b_2 _2922_ (.Y(_0448_),
    .B(net822),
    .A_N(_0446_));
 sg13g2_nor2_1 _2923_ (.A(net512),
    .B(net581),
    .Y(_0006_));
 sg13g2_nor3_1 _2924_ (.A(_2169_),
    .B(_0441_),
    .C(net581),
    .Y(_0008_));
 sg13g2_xor2_1 _2925_ (.B(_0441_),
    .A(net238),
    .X(_0449_));
 sg13g2_nor2_1 _2926_ (.A(net581),
    .B(net239),
    .Y(_0009_));
 sg13g2_a21oi_1 _2927_ (.A1(\vga.pixel_ctr[2] ),
    .A2(_0441_),
    .Y(_0450_),
    .B1(net447));
 sg13g2_nor3_1 _2928_ (.A(_0443_),
    .B(net581),
    .C(net448),
    .Y(_0010_));
 sg13g2_nor2_1 _2929_ (.A(net506),
    .B(_0443_),
    .Y(_0451_));
 sg13g2_nor3_1 _2930_ (.A(_0444_),
    .B(net581),
    .C(net507),
    .Y(_0011_));
 sg13g2_xor2_1 _2931_ (.B(_0444_),
    .A(net725),
    .X(_0452_));
 sg13g2_nor2_1 _2932_ (.A(net582),
    .B(_0452_),
    .Y(_0012_));
 sg13g2_and3_1 _2933_ (.X(_0453_),
    .A(net494),
    .B(\vga.pixel_ctr[5] ),
    .C(_0444_));
 sg13g2_a21oi_1 _2934_ (.A1(\vga.pixel_ctr[5] ),
    .A2(_0444_),
    .Y(_0454_),
    .B1(net494));
 sg13g2_nor3_1 _2935_ (.A(net582),
    .B(_0453_),
    .C(net495),
    .Y(_0013_));
 sg13g2_xor2_1 _2936_ (.B(_0453_),
    .A(net444),
    .X(_0455_));
 sg13g2_nor2_1 _2937_ (.A(net582),
    .B(net445),
    .Y(_0014_));
 sg13g2_and2_1 _2938_ (.A(\vga.pixel_ctr[7] ),
    .B(_0453_),
    .X(_0456_));
 sg13g2_xor2_1 _2939_ (.B(_0456_),
    .A(net319),
    .X(_0457_));
 sg13g2_nor2_1 _2940_ (.A(net582),
    .B(net320),
    .Y(_0015_));
 sg13g2_a21oi_1 _2941_ (.A1(\vga.pixel_ctr[8] ),
    .A2(_0456_),
    .Y(_0458_),
    .B1(net531));
 sg13g2_nand3_1 _2942_ (.B(\vga.pixel_ctr[8] ),
    .C(_0456_),
    .A(net531),
    .Y(_0459_));
 sg13g2_inv_1 _2943_ (.Y(_0460_),
    .A(_0459_));
 sg13g2_nor3_1 _2944_ (.A(net581),
    .B(net532),
    .C(_0460_),
    .Y(_0016_));
 sg13g2_o21ai_1 _2945_ (.B1(_0448_),
    .Y(_0461_),
    .A1(net221),
    .A2(_0459_));
 sg13g2_a21oi_1 _2946_ (.A1(net221),
    .A2(_0459_),
    .Y(_0007_),
    .B1(_0461_));
 sg13g2_nor2_1 _2947_ (.A(_2169_),
    .B(_0442_),
    .Y(_0462_));
 sg13g2_nor3_2 _2948_ (.A(_1948_),
    .B(_2169_),
    .C(_0442_),
    .Y(_0463_));
 sg13g2_o21ai_1 _2949_ (.B1(net444),
    .Y(_0464_),
    .A1(\vga.pixel_ctr[6] ),
    .A2(_0463_));
 sg13g2_xor2_1 _2950_ (.B(_0462_),
    .A(_0107_),
    .X(_0465_));
 sg13g2_and2_1 _2951_ (.A(\vga.pixel_ctr[6] ),
    .B(_0463_),
    .X(_0466_));
 sg13g2_o21ai_1 _2952_ (.B1(_0465_),
    .Y(_0467_),
    .A1(_0108_),
    .A2(_0466_));
 sg13g2_inv_1 _2953_ (.Y(_0468_),
    .A(_0467_));
 sg13g2_nand2_1 _2954_ (.Y(_0469_),
    .A(\vga.pixel_ctr[7] ),
    .B(_0466_));
 sg13g2_nand2b_1 _2955_ (.Y(_0470_),
    .B(_0109_),
    .A_N(\vga.pixel_ctr[8] ));
 sg13g2_xnor2_1 _2956_ (.Y(_0471_),
    .A(\vga.pixel_ctr[9] ),
    .B(_0470_));
 sg13g2_o21ai_1 _2957_ (.B1(_0471_),
    .Y(_0472_),
    .A1(\vga.pixel_ctr[8] ),
    .A2(_0469_));
 sg13g2_a221oi_1 _2958_ (.B2(\vga.pixel_ctr[8] ),
    .C1(_0472_),
    .B1(_0469_),
    .A1(_0464_),
    .Y(_0473_),
    .A2(_0468_));
 sg13g2_nand2_1 _2959_ (.Y(_0474_),
    .A(_2177_),
    .B(_0469_));
 sg13g2_xnor2_1 _2960_ (.Y(_0475_),
    .A(net785),
    .B(_0474_));
 sg13g2_nor4_2 _2961_ (.A(net512),
    .B(_2176_),
    .C(_0473_),
    .Y(\vga.read ),
    .D(_0475_));
 sg13g2_nor2_1 _2962_ (.A(_1917_),
    .B(_2158_),
    .Y(_0000_));
 sg13g2_and2_2 _2963_ (.A(net361),
    .B(net287),
    .X(_0476_));
 sg13g2_nor3_1 _2964_ (.A(\vga.timing_v.pixel[3] ),
    .B(\vga.timing_v.pixel[2] ),
    .C(_0476_),
    .Y(_0477_));
 sg13g2_nand4_1 _2965_ (.B(\vga.timing_v.pixel[6] ),
    .C(\vga.timing_v.pixel[5] ),
    .A(_1958_),
    .Y(_0478_),
    .D(\vga.timing_v.pixel[4] ));
 sg13g2_nor2b_1 _2966_ (.A(\vga.timing_v.pixel[8] ),
    .B_N(_0101_),
    .Y(_0479_));
 sg13g2_o21ai_1 _2967_ (.B1(_0479_),
    .Y(_0480_),
    .A1(_0477_),
    .A2(_0478_));
 sg13g2_nand2_1 _2968_ (.Y(_0481_),
    .A(net311),
    .B(_0480_));
 sg13g2_nand2_2 _2969_ (.Y(_0482_),
    .A(net581),
    .B(_0481_));
 sg13g2_nand2_1 _2970_ (.Y(_0483_),
    .A(net287),
    .B(_0448_));
 sg13g2_o21ai_1 _2971_ (.B1(_0483_),
    .Y(_0217_),
    .A1(net287),
    .A2(_0482_));
 sg13g2_nor3_1 _2972_ (.A(_2165_),
    .B(_0476_),
    .C(_0482_),
    .Y(_0484_));
 sg13g2_a21o_1 _2973_ (.A2(_0448_),
    .A1(net361),
    .B1(_0484_),
    .X(_0218_));
 sg13g2_nand2_1 _2974_ (.Y(_0485_),
    .A(net752),
    .B(_0448_));
 sg13g2_xnor2_1 _2975_ (.Y(_0486_),
    .A(net752),
    .B(_0476_));
 sg13g2_o21ai_1 _2976_ (.B1(_0485_),
    .Y(_0219_),
    .A1(_0482_),
    .A2(_0486_));
 sg13g2_and3_1 _2977_ (.X(_0487_),
    .A(\vga.timing_v.pixel[2] ),
    .B(net582),
    .C(_0476_));
 sg13g2_nor2_2 _2978_ (.A(_0448_),
    .B(_0481_),
    .Y(_0488_));
 sg13g2_xnor2_1 _2979_ (.Y(_0489_),
    .A(net731),
    .B(_0487_));
 sg13g2_nor2_1 _2980_ (.A(_0488_),
    .B(_0489_),
    .Y(_0220_));
 sg13g2_a21oi_1 _2981_ (.A1(\vga.timing_v.pixel[3] ),
    .A2(_0487_),
    .Y(_0490_),
    .B1(net351));
 sg13g2_and3_1 _2982_ (.X(_0491_),
    .A(\vga.timing_v.pixel[2] ),
    .B(_2175_),
    .C(_0476_));
 sg13g2_a21oi_1 _2983_ (.A1(net582),
    .A2(_0491_),
    .Y(_0492_),
    .B1(_0488_));
 sg13g2_nor2b_1 _2984_ (.A(net352),
    .B_N(_0492_),
    .Y(_0221_));
 sg13g2_a21oi_1 _2985_ (.A1(net581),
    .A2(_0491_),
    .Y(_0493_),
    .B1(net396));
 sg13g2_and3_1 _2986_ (.X(_0494_),
    .A(net396),
    .B(_2175_),
    .C(_0487_));
 sg13g2_nor3_1 _2987_ (.A(_0488_),
    .B(_0493_),
    .C(_0494_),
    .Y(_0222_));
 sg13g2_xnor2_1 _2988_ (.Y(_0495_),
    .A(net481),
    .B(_0494_));
 sg13g2_and3_1 _2989_ (.X(_0496_),
    .A(\vga.timing_v.pixel[6] ),
    .B(\vga.timing_v.pixel[5] ),
    .C(_0491_));
 sg13g2_nor2_1 _2990_ (.A(_0488_),
    .B(_0495_),
    .Y(_0223_));
 sg13g2_nand2_1 _2991_ (.Y(_0497_),
    .A(net356),
    .B(_0448_));
 sg13g2_xor2_1 _2992_ (.B(_0496_),
    .A(_0101_),
    .X(_0498_));
 sg13g2_o21ai_1 _2993_ (.B1(_0497_),
    .Y(_0224_),
    .A1(_0482_),
    .A2(_0498_));
 sg13g2_nand3_1 _2994_ (.B(net356),
    .C(_0496_),
    .A(net408),
    .Y(_0499_));
 sg13g2_nand2_1 _2995_ (.Y(_0500_),
    .A(net408),
    .B(_0448_));
 sg13g2_a21o_1 _2996_ (.A2(_0496_),
    .A1(net356),
    .B1(net408),
    .X(_0501_));
 sg13g2_nand2_1 _2997_ (.Y(_0502_),
    .A(_0499_),
    .B(_0501_));
 sg13g2_o21ai_1 _2998_ (.B1(_0500_),
    .Y(_0225_),
    .A1(_0482_),
    .A2(_0502_));
 sg13g2_nand2_1 _2999_ (.Y(_0503_),
    .A(net311),
    .B(_0448_));
 sg13g2_xnor2_1 _3000_ (.Y(_0504_),
    .A(_0103_),
    .B(_0499_));
 sg13g2_o21ai_1 _3001_ (.B1(_0503_),
    .Y(_0226_),
    .A1(_0482_),
    .A2(_0504_));
 sg13g2_nor2_1 _3002_ (.A(net685),
    .B(net580),
    .Y(_0505_));
 sg13g2_a22oi_1 _3003_ (.Y(_0506_),
    .B1(net412),
    .B2(net562),
    .A2(net704),
    .A1(net687));
 sg13g2_inv_1 _3004_ (.Y(_0227_),
    .A(_0506_));
 sg13g2_nand2_1 _3005_ (.Y(_0507_),
    .A(net661),
    .B(_1910_));
 sg13g2_nand2b_1 _3006_ (.Y(_0508_),
    .B(net580),
    .A_N(_0507_));
 sg13g2_nand2_1 _3007_ (.Y(_0509_),
    .A(\mandelbrot.alu.in_ci[0] ),
    .B(\mandelbrot.alu.m3[13] ));
 sg13g2_xnor2_1 _3008_ (.Y(_0510_),
    .A(net768),
    .B(net371));
 sg13g2_nand2_1 _3009_ (.Y(_0511_),
    .A(net686),
    .B(net733));
 sg13g2_o21ai_1 _3010_ (.B1(_0511_),
    .Y(_0512_),
    .A1(net556),
    .A2(_0510_));
 sg13g2_a21o_1 _3011_ (.A2(net561),
    .A1(net762),
    .B1(_0512_),
    .X(_0228_));
 sg13g2_nand2_1 _3012_ (.Y(_0513_),
    .A(\mandelbrot.alu.in_ci[1] ),
    .B(\mandelbrot.alu.m3[14] ));
 sg13g2_xnor2_1 _3013_ (.Y(_0514_),
    .A(\mandelbrot.alu.in_ci[1] ),
    .B(\mandelbrot.alu.m3[14] ));
 sg13g2_xnor2_1 _3014_ (.Y(_0515_),
    .A(_0509_),
    .B(_0514_));
 sg13g2_a22oi_1 _3015_ (.Y(_0516_),
    .B1(net705),
    .B2(net561),
    .A2(net727),
    .A1(net686));
 sg13g2_o21ai_1 _3016_ (.B1(_0516_),
    .Y(_0229_),
    .A1(net556),
    .A2(_0515_));
 sg13g2_o21ai_1 _3017_ (.B1(_0513_),
    .Y(_0517_),
    .A1(_0509_),
    .A2(_0514_));
 sg13g2_and2_1 _3018_ (.A(\mandelbrot.alu.in_ci[2] ),
    .B(\mandelbrot.alu.m3[15] ),
    .X(_0518_));
 sg13g2_xor2_1 _3019_ (.B(\mandelbrot.alu.m3[15] ),
    .A(\mandelbrot.alu.in_ci[2] ),
    .X(_0519_));
 sg13g2_xnor2_1 _3020_ (.Y(_0520_),
    .A(_0517_),
    .B(_0519_));
 sg13g2_a22oi_1 _3021_ (.Y(_0521_),
    .B1(net733),
    .B2(net563),
    .A2(\mandelbrot.alu.m2[4] ),
    .A1(net686));
 sg13g2_o21ai_1 _3022_ (.B1(net734),
    .Y(_0230_),
    .A1(net556),
    .A2(_0520_));
 sg13g2_nand2_1 _3023_ (.Y(_0522_),
    .A(\mandelbrot.alu.in_ci[3] ),
    .B(\mandelbrot.alu.m3[16] ));
 sg13g2_xnor2_1 _3024_ (.Y(_0523_),
    .A(\mandelbrot.alu.in_ci[3] ),
    .B(\mandelbrot.alu.m3[16] ));
 sg13g2_a21oi_1 _3025_ (.A1(_0517_),
    .A2(_0519_),
    .Y(_0524_),
    .B1(_0518_));
 sg13g2_xnor2_1 _3026_ (.Y(_0525_),
    .A(_0523_),
    .B(_0524_));
 sg13g2_nand2_1 _3027_ (.Y(_0526_),
    .A(net686),
    .B(net710));
 sg13g2_o21ai_1 _3028_ (.B1(_0526_),
    .Y(_0527_),
    .A1(net556),
    .A2(_0525_));
 sg13g2_a21o_1 _3029_ (.A2(net561),
    .A1(net727),
    .B1(_0527_),
    .X(_0231_));
 sg13g2_o21ai_1 _3030_ (.B1(_0522_),
    .Y(_0528_),
    .A1(_0523_),
    .A2(_0524_));
 sg13g2_and2_1 _3031_ (.A(\mandelbrot.alu.in_ci[4] ),
    .B(\mandelbrot.alu.m3[17] ),
    .X(_0529_));
 sg13g2_xor2_1 _3032_ (.B(\mandelbrot.alu.m3[17] ),
    .A(\mandelbrot.alu.in_ci[4] ),
    .X(_0530_));
 sg13g2_xnor2_1 _3033_ (.Y(_0531_),
    .A(_0528_),
    .B(_0530_));
 sg13g2_nand2_1 _3034_ (.Y(_0532_),
    .A(net686),
    .B(\mandelbrot.alu.m2[6] ));
 sg13g2_o21ai_1 _3035_ (.B1(_0532_),
    .Y(_0533_),
    .A1(net556),
    .A2(_0531_));
 sg13g2_a21o_1 _3036_ (.A2(net561),
    .A1(net736),
    .B1(_0533_),
    .X(_0232_));
 sg13g2_a21oi_1 _3037_ (.A1(_0528_),
    .A2(_0530_),
    .Y(_0534_),
    .B1(_0529_));
 sg13g2_nor2_1 _3038_ (.A(\mandelbrot.alu.in_ci[5] ),
    .B(\mandelbrot.alu.m3[18] ),
    .Y(_0535_));
 sg13g2_xnor2_1 _3039_ (.Y(_0536_),
    .A(\mandelbrot.alu.in_ci[5] ),
    .B(\mandelbrot.alu.m3[18] ));
 sg13g2_xnor2_1 _3040_ (.Y(_0537_),
    .A(_0534_),
    .B(_0536_));
 sg13g2_nand2_1 _3041_ (.Y(_0538_),
    .A(net686),
    .B(\mandelbrot.alu.m2[7] ));
 sg13g2_o21ai_1 _3042_ (.B1(_0538_),
    .Y(_0539_),
    .A1(net556),
    .A2(_0537_));
 sg13g2_a21o_1 _3043_ (.A2(net563),
    .A1(net710),
    .B1(_0539_),
    .X(_0233_));
 sg13g2_nand2_1 _3044_ (.Y(_0540_),
    .A(net516),
    .B(\mandelbrot.alu.m3[19] ));
 sg13g2_xnor2_1 _3045_ (.Y(_0541_),
    .A(\mandelbrot.alu.in_ci[6] ),
    .B(\mandelbrot.alu.m3[19] ));
 sg13g2_a221oi_1 _3046_ (.B2(_0530_),
    .C1(_0529_),
    .B1(_0528_),
    .A1(\mandelbrot.alu.in_ci[5] ),
    .Y(_0542_),
    .A2(\mandelbrot.alu.m3[18] ));
 sg13g2_or3_1 _3047_ (.A(_0535_),
    .B(_0541_),
    .C(_0542_),
    .X(_0543_));
 sg13g2_o21ai_1 _3048_ (.B1(_0541_),
    .Y(_0544_),
    .A1(_0535_),
    .A2(_0542_));
 sg13g2_nand2_2 _3049_ (.Y(_0545_),
    .A(_0543_),
    .B(_0544_));
 sg13g2_nand2_1 _3050_ (.Y(_0546_),
    .A(net686),
    .B(\mandelbrot.alu.m2[8] ));
 sg13g2_o21ai_1 _3051_ (.B1(_0546_),
    .Y(_0547_),
    .A1(net556),
    .A2(_0545_));
 sg13g2_a21o_1 _3052_ (.A2(net563),
    .A1(net760),
    .B1(_0547_),
    .X(_0234_));
 sg13g2_and2_1 _3053_ (.A(\mandelbrot.alu.in_ci[7] ),
    .B(\mandelbrot.alu.m3[20] ),
    .X(_0548_));
 sg13g2_xnor2_1 _3054_ (.Y(_0549_),
    .A(\mandelbrot.alu.in_ci[7] ),
    .B(\mandelbrot.alu.m3[20] ));
 sg13g2_a21oi_1 _3055_ (.A1(_0540_),
    .A2(_0543_),
    .Y(_0550_),
    .B1(_0549_));
 sg13g2_nand3_1 _3056_ (.B(_0543_),
    .C(_0549_),
    .A(_0540_),
    .Y(_0551_));
 sg13g2_nand2b_2 _3057_ (.Y(_0552_),
    .B(_0551_),
    .A_N(_0550_));
 sg13g2_a22oi_1 _3058_ (.Y(_0553_),
    .B1(net795),
    .B2(net561),
    .A2(net527),
    .A1(net686));
 sg13g2_o21ai_1 _3059_ (.B1(_0553_),
    .Y(_0235_),
    .A1(net556),
    .A2(_0552_));
 sg13g2_nand2_1 _3060_ (.Y(_0554_),
    .A(\mandelbrot.alu.in_ci[8] ),
    .B(\mandelbrot.alu.m3[21] ));
 sg13g2_xor2_1 _3061_ (.B(\mandelbrot.alu.m3[21] ),
    .A(\mandelbrot.alu.in_ci[8] ),
    .X(_0555_));
 sg13g2_o21ai_1 _3062_ (.B1(_0555_),
    .Y(_0556_),
    .A1(_0548_),
    .A2(_0550_));
 sg13g2_or3_1 _3063_ (.A(_0548_),
    .B(_0550_),
    .C(_0555_),
    .X(_0557_));
 sg13g2_nand2_2 _3064_ (.Y(_0558_),
    .A(_0556_),
    .B(_0557_));
 sg13g2_nand2_1 _3065_ (.Y(_0559_),
    .A(net685),
    .B(net825));
 sg13g2_o21ai_1 _3066_ (.B1(_0559_),
    .Y(_0560_),
    .A1(net557),
    .A2(_0558_));
 sg13g2_a21o_1 _3067_ (.A2(net560),
    .A1(net771),
    .B1(_0560_),
    .X(_0236_));
 sg13g2_and2_1 _3068_ (.A(_0554_),
    .B(_0556_),
    .X(_0561_));
 sg13g2_and2_1 _3069_ (.A(\mandelbrot.alu.in_ci[9] ),
    .B(\mandelbrot.alu.m3[22] ),
    .X(_0562_));
 sg13g2_nor2_1 _3070_ (.A(\mandelbrot.alu.in_ci[9] ),
    .B(\mandelbrot.alu.m3[22] ),
    .Y(_0563_));
 sg13g2_nor2_1 _3071_ (.A(_0562_),
    .B(_0563_),
    .Y(_0564_));
 sg13g2_xor2_1 _3072_ (.B(_0564_),
    .A(_0561_),
    .X(_0565_));
 sg13g2_nand2_1 _3073_ (.Y(_0566_),
    .A(net687),
    .B(\mandelbrot.alu.m2[11] ));
 sg13g2_o21ai_1 _3074_ (.B1(_0566_),
    .Y(_0567_),
    .A1(net557),
    .A2(_0565_));
 sg13g2_a21o_1 _3075_ (.A2(net561),
    .A1(net527),
    .B1(_0567_),
    .X(_0237_));
 sg13g2_nand2_1 _3076_ (.Y(_0568_),
    .A(\mandelbrot.alu.in_ci[10] ),
    .B(\mandelbrot.alu.m3[23] ));
 sg13g2_xnor2_1 _3077_ (.Y(_0569_),
    .A(\mandelbrot.alu.in_ci[10] ),
    .B(\mandelbrot.alu.m3[23] ));
 sg13g2_inv_1 _3078_ (.Y(_0570_),
    .A(_0569_));
 sg13g2_a21oi_1 _3079_ (.A1(_0554_),
    .A2(_0556_),
    .Y(_0571_),
    .B1(_0563_));
 sg13g2_nor2_1 _3080_ (.A(_0562_),
    .B(_0571_),
    .Y(_0572_));
 sg13g2_o21ai_1 _3081_ (.B1(_0570_),
    .Y(_0573_),
    .A1(_0562_),
    .A2(_0571_));
 sg13g2_xnor2_1 _3082_ (.Y(_0574_),
    .A(_0569_),
    .B(_0572_));
 sg13g2_nand2_1 _3083_ (.Y(_0575_),
    .A(net685),
    .B(net792));
 sg13g2_o21ai_1 _3084_ (.B1(_0575_),
    .Y(_0576_),
    .A1(net557),
    .A2(_0574_));
 sg13g2_a21o_1 _3085_ (.A2(net560),
    .A1(net800),
    .B1(_0576_),
    .X(_0238_));
 sg13g2_nand2_1 _3086_ (.Y(_0577_),
    .A(_0568_),
    .B(_0573_));
 sg13g2_and2_1 _3087_ (.A(\mandelbrot.alu.in_ci[11] ),
    .B(\mandelbrot.alu.m3[24] ),
    .X(_0578_));
 sg13g2_nor2_1 _3088_ (.A(\mandelbrot.alu.in_ci[11] ),
    .B(\mandelbrot.alu.m3[24] ),
    .Y(_0579_));
 sg13g2_nor2_1 _3089_ (.A(_0578_),
    .B(_0579_),
    .Y(_0580_));
 sg13g2_xnor2_1 _3090_ (.Y(_0581_),
    .A(_0577_),
    .B(_0580_));
 sg13g2_nand2_1 _3091_ (.Y(_0582_),
    .A(net687),
    .B(\mandelbrot.alu.m2[13] ));
 sg13g2_o21ai_1 _3092_ (.B1(_0582_),
    .Y(_0583_),
    .A1(net557),
    .A2(_0581_));
 sg13g2_a21o_1 _3093_ (.A2(net561),
    .A1(net740),
    .B1(_0583_),
    .X(_0239_));
 sg13g2_xnor2_1 _3094_ (.Y(_0584_),
    .A(\mandelbrot.alu.in_ci[12] ),
    .B(\mandelbrot.alu.m3[25] ));
 sg13g2_inv_1 _3095_ (.Y(_0585_),
    .A(_0584_));
 sg13g2_a21oi_1 _3096_ (.A1(_0568_),
    .A2(_0573_),
    .Y(_0586_),
    .B1(_0579_));
 sg13g2_nor2_1 _3097_ (.A(_0578_),
    .B(_0586_),
    .Y(_0587_));
 sg13g2_o21ai_1 _3098_ (.B1(_0585_),
    .Y(_0588_),
    .A1(_0578_),
    .A2(_0586_));
 sg13g2_xnor2_1 _3099_ (.Y(_0589_),
    .A(_0584_),
    .B(_0587_));
 sg13g2_nand2_1 _3100_ (.Y(_0590_),
    .A(net685),
    .B(net827));
 sg13g2_o21ai_1 _3101_ (.B1(_0590_),
    .Y(_0591_),
    .A1(net557),
    .A2(_0589_));
 sg13g2_a21o_1 _3102_ (.A2(net560),
    .A1(net792),
    .B1(_0591_),
    .X(_0240_));
 sg13g2_nor2_1 _3103_ (.A(\mandelbrot.alu.in_ci[13] ),
    .B(\mandelbrot.alu.m3[26] ),
    .Y(_0592_));
 sg13g2_xor2_1 _3104_ (.B(\mandelbrot.alu.m3[26] ),
    .A(\mandelbrot.alu.in_ci[13] ),
    .X(_0593_));
 sg13g2_o21ai_1 _3105_ (.B1(_0588_),
    .Y(_0594_),
    .A1(_1951_),
    .A2(_1952_));
 sg13g2_xnor2_1 _3106_ (.Y(_0595_),
    .A(_0593_),
    .B(_0594_));
 sg13g2_nand2_1 _3107_ (.Y(_0596_),
    .A(net687),
    .B(\mandelbrot.alu.m2[15] ));
 sg13g2_o21ai_1 _3108_ (.B1(_0596_),
    .Y(_0597_),
    .A1(net557),
    .A2(_0595_));
 sg13g2_a21o_1 _3109_ (.A2(net561),
    .A1(net744),
    .B1(_0597_),
    .X(_0241_));
 sg13g2_and2_1 _3110_ (.A(\mandelbrot.alu.in_ci[14] ),
    .B(\mandelbrot.alu.m3[27] ),
    .X(_0598_));
 sg13g2_xor2_1 _3111_ (.B(\mandelbrot.alu.m3[27] ),
    .A(\mandelbrot.alu.in_ci[14] ),
    .X(_0599_));
 sg13g2_a22oi_1 _3112_ (.Y(_0600_),
    .B1(\mandelbrot.alu.in_ci[12] ),
    .B2(\mandelbrot.alu.m3[25] ),
    .A2(\mandelbrot.alu.m3[26] ),
    .A1(\mandelbrot.alu.in_ci[13] ));
 sg13g2_a21o_1 _3113_ (.A2(_0600_),
    .A1(_0588_),
    .B1(_0592_),
    .X(_0601_));
 sg13g2_nor2b_1 _3114_ (.A(_0601_),
    .B_N(_0599_),
    .Y(_0602_));
 sg13g2_xor2_1 _3115_ (.B(_0601_),
    .A(_0599_),
    .X(_0603_));
 sg13g2_nand2_1 _3116_ (.Y(_0604_),
    .A(\mandelbrot.alu.m2[0] ),
    .B(\mandelbrot.alu.mult_zi_zi.shift_reg[0] ));
 sg13g2_a21o_1 _3117_ (.A2(\mandelbrot.alu.mult_zi_zi.shift_reg[0] ),
    .A1(\mandelbrot.alu.m2[0] ),
    .B1(net704),
    .X(_0605_));
 sg13g2_nor2_1 _3118_ (.A(\mandelbrot.alu.m2[0] ),
    .B(\mandelbrot.alu.mult_zi_zi.shift_reg[0] ),
    .Y(_0606_));
 sg13g2_o21ai_1 _3119_ (.B1(net704),
    .Y(_0607_),
    .A1(\mandelbrot.alu.m2[0] ),
    .A2(\mandelbrot.alu.mult_zi_zi.shift_reg[0] ));
 sg13g2_nand2_2 _3120_ (.Y(_0608_),
    .A(_0605_),
    .B(_0607_));
 sg13g2_nor2_1 _3121_ (.A(net704),
    .B(_0606_),
    .Y(_0609_));
 sg13g2_a21oi_1 _3122_ (.A1(net706),
    .A2(_0604_),
    .Y(_0610_),
    .B1(_0609_));
 sg13g2_a21o_1 _3123_ (.A2(_0604_),
    .A1(net706),
    .B1(_0609_),
    .X(_0611_));
 sg13g2_nand3_1 _3124_ (.B(net644),
    .C(net605),
    .A(\mandelbrot.alu.in_zi[0] ),
    .Y(_0612_));
 sg13g2_a21oi_1 _3125_ (.A1(_1922_),
    .A2(_0612_),
    .Y(_0613_),
    .B1(_1910_));
 sg13g2_o21ai_1 _3126_ (.B1(_0613_),
    .Y(_0614_),
    .A1(_1922_),
    .A2(_0612_));
 sg13g2_o21ai_1 _3127_ (.B1(_0614_),
    .Y(_0615_),
    .A1(_0507_),
    .A2(_0603_));
 sg13g2_mux2_1 _3128_ (.A0(_0615_),
    .A1(net815),
    .S(net560),
    .X(_0242_));
 sg13g2_nand2_1 _3129_ (.Y(_0616_),
    .A(\mandelbrot.alu.in_ci[15] ),
    .B(\mandelbrot.alu.m3[28] ));
 sg13g2_xor2_1 _3130_ (.B(\mandelbrot.alu.m3[28] ),
    .A(\mandelbrot.alu.in_ci[15] ),
    .X(_0617_));
 sg13g2_nor2_1 _3131_ (.A(_0598_),
    .B(_0602_),
    .Y(_0618_));
 sg13g2_nand2_1 _3132_ (.Y(_0619_),
    .A(_0599_),
    .B(_0617_));
 sg13g2_xor2_1 _3133_ (.B(_0618_),
    .A(_0617_),
    .X(_0620_));
 sg13g2_nor2_1 _3134_ (.A(_0507_),
    .B(_0620_),
    .Y(_0621_));
 sg13g2_nand3_1 _3135_ (.B(net671),
    .C(net644),
    .A(\mandelbrot.alu.m2[16] ),
    .Y(_0622_));
 sg13g2_xnor2_1 _3136_ (.Y(_0623_),
    .A(net671),
    .B(\mandelbrot.alu.in_zi[1] ));
 sg13g2_nor2b_1 _3137_ (.A(net705),
    .B_N(_0046_),
    .Y(_0624_));
 sg13g2_a221oi_1 _3138_ (.B2(net704),
    .C1(_0624_),
    .B1(_0623_),
    .A1(_0605_),
    .Y(_0625_),
    .A2(_0607_));
 sg13g2_and3_1 _3139_ (.X(_0626_),
    .A(_1969_),
    .B(_0605_),
    .C(_0607_));
 sg13g2_nor2_1 _3140_ (.A(_0625_),
    .B(_0626_),
    .Y(_0627_));
 sg13g2_o21ai_1 _3141_ (.B1(\mandelbrot.alu.m2[17] ),
    .Y(_0628_),
    .A1(_0625_),
    .A2(_0626_));
 sg13g2_nor3_1 _3142_ (.A(\mandelbrot.alu.m2[17] ),
    .B(_0625_),
    .C(_0626_),
    .Y(_0629_));
 sg13g2_xor2_1 _3143_ (.B(_0627_),
    .A(\mandelbrot.alu.m2[17] ),
    .X(_0630_));
 sg13g2_xnor2_1 _3144_ (.Y(_0631_),
    .A(_0622_),
    .B(_0630_));
 sg13g2_o21ai_1 _3145_ (.B1(net688),
    .Y(_0632_),
    .A1(\mandelbrot.alu.m2[17] ),
    .A2(net604));
 sg13g2_a21oi_1 _3146_ (.A1(net604),
    .A2(_0631_),
    .Y(_0633_),
    .B1(_0632_));
 sg13g2_nor3_1 _3147_ (.A(net562),
    .B(_0621_),
    .C(_0633_),
    .Y(_0634_));
 sg13g2_a21oi_1 _3148_ (.A1(_1923_),
    .A2(net562),
    .Y(_0243_),
    .B1(_0634_));
 sg13g2_o21ai_1 _3149_ (.B1(_0628_),
    .Y(_0635_),
    .A1(_0622_),
    .A2(_0629_));
 sg13g2_nor3_1 _3150_ (.A(net671),
    .B(\mandelbrot.alu.in_zi[1] ),
    .C(\mandelbrot.alu.in_zi[2] ),
    .Y(_0636_));
 sg13g2_o21ai_1 _3151_ (.B1(\mandelbrot.alu.in_zi[2] ),
    .Y(_0637_),
    .A1(net671),
    .A2(\mandelbrot.alu.in_zi[1] ));
 sg13g2_nand2b_2 _3152_ (.Y(_0638_),
    .B(_0637_),
    .A_N(_0636_));
 sg13g2_mux2_1 _3153_ (.A0(_0045_),
    .A1(_0638_),
    .S(net706),
    .X(_0639_));
 sg13g2_mux4_1 _3154_ (.S0(net644),
    .A0(_0046_),
    .A1(_0045_),
    .A2(_0623_),
    .A3(_0638_),
    .S1(net704),
    .X(_0640_));
 sg13g2_xnor2_1 _3155_ (.Y(_0641_),
    .A(\mandelbrot.alu.m2[18] ),
    .B(_0640_));
 sg13g2_xor2_1 _3156_ (.B(_0641_),
    .A(_0635_),
    .X(_0642_));
 sg13g2_nor2_1 _3157_ (.A(net608),
    .B(_0642_),
    .Y(_0643_));
 sg13g2_a21oi_1 _3158_ (.A1(net378),
    .A2(net608),
    .Y(_0644_),
    .B1(_0643_));
 sg13g2_a22oi_1 _3159_ (.Y(_0645_),
    .B1(_0644_),
    .B2(net688),
    .A2(net562),
    .A1(\mandelbrot.alu.m2[16] ));
 sg13g2_inv_1 _3160_ (.Y(_0244_),
    .A(net379));
 sg13g2_nor2_1 _3161_ (.A(net706),
    .B(_0044_),
    .Y(_0646_));
 sg13g2_or4_2 _3162_ (.A(net671),
    .B(\mandelbrot.alu.in_zi[1] ),
    .C(\mandelbrot.alu.in_zi[2] ),
    .D(\mandelbrot.alu.in_zi[3] ),
    .X(_0647_));
 sg13g2_xnor2_1 _3163_ (.Y(_0648_),
    .A(\mandelbrot.alu.in_zi[3] ),
    .B(_0636_));
 sg13g2_a21oi_1 _3164_ (.A1(net706),
    .A2(_0648_),
    .Y(_0649_),
    .B1(_0646_));
 sg13g2_mux2_1 _3165_ (.A0(_0639_),
    .A1(_0649_),
    .S(net644),
    .X(_0650_));
 sg13g2_nand2b_1 _3166_ (.Y(_0651_),
    .B(\mandelbrot.alu.m2[19] ),
    .A_N(_0650_));
 sg13g2_nor2b_1 _3167_ (.A(\mandelbrot.alu.m2[19] ),
    .B_N(_0650_),
    .Y(_0652_));
 sg13g2_xnor2_1 _3168_ (.Y(_0653_),
    .A(\mandelbrot.alu.m2[19] ),
    .B(_0650_));
 sg13g2_nor2_1 _3169_ (.A(_0100_),
    .B(_0640_),
    .Y(_0654_));
 sg13g2_a21oi_1 _3170_ (.A1(_0635_),
    .A2(_0641_),
    .Y(_0655_),
    .B1(_0654_));
 sg13g2_xnor2_1 _3171_ (.Y(_0656_),
    .A(_0653_),
    .B(_0655_));
 sg13g2_nor2_1 _3172_ (.A(net608),
    .B(_0656_),
    .Y(_0657_));
 sg13g2_a21oi_1 _3173_ (.A1(net280),
    .A2(net608),
    .Y(_0658_),
    .B1(_0657_));
 sg13g2_a22oi_1 _3174_ (.Y(_0659_),
    .B1(_0658_),
    .B2(net688),
    .A2(net563),
    .A1(\mandelbrot.alu.m2[17] ));
 sg13g2_inv_1 _3175_ (.Y(_0245_),
    .A(net281));
 sg13g2_o21ai_1 _3176_ (.B1(_0651_),
    .Y(_0660_),
    .A1(_0652_),
    .A2(_0655_));
 sg13g2_nor2_1 _3177_ (.A(net706),
    .B(_0043_),
    .Y(_0661_));
 sg13g2_xor2_1 _3178_ (.B(_0647_),
    .A(\mandelbrot.alu.in_zi[4] ),
    .X(_0662_));
 sg13g2_a21oi_2 _3179_ (.B1(_0661_),
    .Y(_0663_),
    .A2(_0662_),
    .A1(net706));
 sg13g2_mux2_1 _3180_ (.A0(_0649_),
    .A1(_0663_),
    .S(_0608_),
    .X(_0664_));
 sg13g2_inv_1 _3181_ (.Y(_0665_),
    .A(_0664_));
 sg13g2_xnor2_1 _3182_ (.Y(_0666_),
    .A(\mandelbrot.alu.m2[20] ),
    .B(_0664_));
 sg13g2_xnor2_1 _3183_ (.Y(_0667_),
    .A(_0660_),
    .B(_0666_));
 sg13g2_o21ai_1 _3184_ (.B1(net688),
    .Y(_0668_),
    .A1(_1970_),
    .A2(net605));
 sg13g2_a21oi_1 _3185_ (.A1(net605),
    .A2(_0667_),
    .Y(_0669_),
    .B1(_0668_));
 sg13g2_a21o_1 _3186_ (.A2(net562),
    .A1(\mandelbrot.alu.m2[18] ),
    .B1(_0669_),
    .X(_0246_));
 sg13g2_a22oi_1 _3187_ (.Y(_0670_),
    .B1(_0666_),
    .B2(_0660_),
    .A2(_0665_),
    .A1(_1970_));
 sg13g2_or2_1 _3188_ (.X(_0671_),
    .B(_0042_),
    .A(net706));
 sg13g2_nor3_1 _3189_ (.A(\mandelbrot.alu.in_zi[4] ),
    .B(\mandelbrot.alu.in_zi[5] ),
    .C(_0647_),
    .Y(_0672_));
 sg13g2_o21ai_1 _3190_ (.B1(\mandelbrot.alu.in_zi[5] ),
    .Y(_0673_),
    .A1(\mandelbrot.alu.in_zi[4] ),
    .A2(_0647_));
 sg13g2_nand2b_1 _3191_ (.Y(_0674_),
    .B(_0673_),
    .A_N(_0672_));
 sg13g2_o21ai_1 _3192_ (.B1(_0671_),
    .Y(_0675_),
    .A1(_1934_),
    .A2(_0674_));
 sg13g2_nor2_1 _3193_ (.A(net644),
    .B(_0663_),
    .Y(_0676_));
 sg13g2_a21oi_1 _3194_ (.A1(net644),
    .A2(_0675_),
    .Y(_0677_),
    .B1(_0676_));
 sg13g2_nor2b_1 _3195_ (.A(_0677_),
    .B_N(\mandelbrot.alu.m2[21] ),
    .Y(_0678_));
 sg13g2_nor2b_1 _3196_ (.A(\mandelbrot.alu.m2[21] ),
    .B_N(_0677_),
    .Y(_0679_));
 sg13g2_nor2_1 _3197_ (.A(_0678_),
    .B(_0679_),
    .Y(_0680_));
 sg13g2_xor2_1 _3198_ (.B(_0680_),
    .A(_0670_),
    .X(_0681_));
 sg13g2_nand2_2 _3199_ (.Y(_0682_),
    .A(net684),
    .B(net604));
 sg13g2_nand2b_1 _3200_ (.Y(_0683_),
    .B(net684),
    .A_N(_0097_));
 sg13g2_a22oi_1 _3201_ (.Y(_0684_),
    .B1(_0682_),
    .B2(_0683_),
    .A2(_0681_),
    .A1(net605));
 sg13g2_a21o_1 _3202_ (.A2(net562),
    .A1(net807),
    .B1(_0684_),
    .X(_0247_));
 sg13g2_a221oi_1 _3203_ (.B2(_0660_),
    .C1(_0678_),
    .B1(_0666_),
    .A1(_1970_),
    .Y(_0685_),
    .A2(_0665_));
 sg13g2_nor2_1 _3204_ (.A(net703),
    .B(_0041_),
    .Y(_0686_));
 sg13g2_nor4_2 _3205_ (.A(\mandelbrot.alu.in_zi[4] ),
    .B(\mandelbrot.alu.in_zi[5] ),
    .C(\mandelbrot.alu.in_zi[6] ),
    .Y(_0687_),
    .D(_0647_));
 sg13g2_xnor2_1 _3206_ (.Y(_0688_),
    .A(\mandelbrot.alu.in_zi[6] ),
    .B(_0672_));
 sg13g2_a21oi_2 _3207_ (.B1(_0686_),
    .Y(_0689_),
    .A2(_0688_),
    .A1(net703));
 sg13g2_nand2_1 _3208_ (.Y(_0690_),
    .A(net644),
    .B(_0689_));
 sg13g2_o21ai_1 _3209_ (.B1(_0690_),
    .Y(_0691_),
    .A1(net644),
    .A2(_0675_));
 sg13g2_xor2_1 _3210_ (.B(_0691_),
    .A(\mandelbrot.alu.m2[22] ),
    .X(_0692_));
 sg13g2_nor3_2 _3211_ (.A(_0679_),
    .B(_0685_),
    .C(_0692_),
    .Y(_0693_));
 sg13g2_o21ai_1 _3212_ (.B1(_0692_),
    .Y(_0694_),
    .A1(_0679_),
    .A2(_0685_));
 sg13g2_nor2b_1 _3213_ (.A(_0693_),
    .B_N(_0694_),
    .Y(_0695_));
 sg13g2_o21ai_1 _3214_ (.B1(net685),
    .Y(_0696_),
    .A1(net608),
    .A2(_0695_));
 sg13g2_a21oi_1 _3215_ (.A1(net717),
    .A2(net608),
    .Y(_0697_),
    .B1(_0696_));
 sg13g2_a21o_1 _3216_ (.A2(net562),
    .A1(\mandelbrot.alu.m2[20] ),
    .B1(_0697_),
    .X(_0248_));
 sg13g2_nand2_1 _3217_ (.Y(_0698_),
    .A(\mandelbrot.alu.m2[21] ),
    .B(net559));
 sg13g2_nor2_1 _3218_ (.A(net703),
    .B(_0040_),
    .Y(_0699_));
 sg13g2_nand2b_2 _3219_ (.Y(_0700_),
    .B(_0687_),
    .A_N(\mandelbrot.alu.in_zi[7] ));
 sg13g2_xnor2_1 _3220_ (.Y(_0701_),
    .A(\mandelbrot.alu.in_zi[7] ),
    .B(_0687_));
 sg13g2_a21oi_2 _3221_ (.B1(_0699_),
    .Y(_0702_),
    .A2(_0701_),
    .A1(net703));
 sg13g2_mux2_1 _3222_ (.A0(_0689_),
    .A1(_0702_),
    .S(net643),
    .X(_0703_));
 sg13g2_nand2b_1 _3223_ (.Y(_0704_),
    .B(\mandelbrot.alu.m2[23] ),
    .A_N(_0703_));
 sg13g2_xnor2_1 _3224_ (.Y(_0705_),
    .A(\mandelbrot.alu.m2[23] ),
    .B(_0703_));
 sg13g2_nor2_1 _3225_ (.A(_0096_),
    .B(_0691_),
    .Y(_0706_));
 sg13g2_nor3_1 _3226_ (.A(_0693_),
    .B(_0705_),
    .C(_0706_),
    .Y(_0707_));
 sg13g2_o21ai_1 _3227_ (.B1(_0705_),
    .Y(_0708_),
    .A1(_0693_),
    .A2(_0706_));
 sg13g2_nand2b_1 _3228_ (.Y(_0709_),
    .B(_0708_),
    .A_N(_0707_));
 sg13g2_a21oi_1 _3229_ (.A1(net604),
    .A2(_0709_),
    .Y(_0710_),
    .B1(net267));
 sg13g2_o21ai_1 _3230_ (.B1(_0710_),
    .Y(_0711_),
    .A1(\mandelbrot.alu.m2[23] ),
    .A2(net604));
 sg13g2_o21ai_1 _3231_ (.B1(_0698_),
    .Y(_0249_),
    .A1(net559),
    .A2(_0711_));
 sg13g2_or2_1 _3232_ (.X(_0712_),
    .B(_0039_),
    .A(net703));
 sg13g2_xnor2_1 _3233_ (.Y(_0713_),
    .A(\mandelbrot.alu.in_zi[8] ),
    .B(_0700_));
 sg13g2_o21ai_1 _3234_ (.B1(_0712_),
    .Y(_0714_),
    .A1(_1934_),
    .A2(_0713_));
 sg13g2_nor2_1 _3235_ (.A(net643),
    .B(_0702_),
    .Y(_0715_));
 sg13g2_a21oi_1 _3236_ (.A1(net643),
    .A2(_0714_),
    .Y(_0716_),
    .B1(_0715_));
 sg13g2_xor2_1 _3237_ (.B(_0716_),
    .A(\mandelbrot.alu.m2[24] ),
    .X(_0717_));
 sg13g2_a21oi_1 _3238_ (.A1(_0704_),
    .A2(_0708_),
    .Y(_0718_),
    .B1(_0717_));
 sg13g2_nand3_1 _3239_ (.B(_0708_),
    .C(_0717_),
    .A(_0704_),
    .Y(_0719_));
 sg13g2_nor2b_1 _3240_ (.A(_0718_),
    .B_N(_0719_),
    .Y(_0720_));
 sg13g2_nor2_1 _3241_ (.A(net606),
    .B(_0720_),
    .Y(_0721_));
 sg13g2_a21oi_1 _3242_ (.A1(net440),
    .A2(net607),
    .Y(_0722_),
    .B1(_0721_));
 sg13g2_a22oi_1 _3243_ (.Y(_0723_),
    .B1(_0722_),
    .B2(net684),
    .A2(net559),
    .A1(\mandelbrot.alu.m2[22] ));
 sg13g2_inv_1 _3244_ (.Y(_0250_),
    .A(net441));
 sg13g2_nor2_1 _3245_ (.A(net701),
    .B(_0038_),
    .Y(_0724_));
 sg13g2_nor3_1 _3246_ (.A(\mandelbrot.alu.in_zi[8] ),
    .B(\mandelbrot.alu.in_zi[9] ),
    .C(_0700_),
    .Y(_0725_));
 sg13g2_o21ai_1 _3247_ (.B1(\mandelbrot.alu.in_zi[9] ),
    .Y(_0726_),
    .A1(\mandelbrot.alu.in_zi[8] ),
    .A2(_0700_));
 sg13g2_nor2b_1 _3248_ (.A(_0725_),
    .B_N(_0726_),
    .Y(_0727_));
 sg13g2_a21oi_1 _3249_ (.A1(net701),
    .A2(_0727_),
    .Y(_0728_),
    .B1(_0724_));
 sg13g2_nand2_1 _3250_ (.Y(_0729_),
    .A(net643),
    .B(_0728_));
 sg13g2_o21ai_1 _3251_ (.B1(_0729_),
    .Y(_0730_),
    .A1(net643),
    .A2(_0714_));
 sg13g2_nand2b_1 _3252_ (.Y(_0731_),
    .B(_0730_),
    .A_N(net700));
 sg13g2_nor2b_1 _3253_ (.A(_0730_),
    .B_N(net700),
    .Y(_0732_));
 sg13g2_xor2_1 _3254_ (.B(_0730_),
    .A(net700),
    .X(_0733_));
 sg13g2_nor2_1 _3255_ (.A(_0095_),
    .B(_0716_),
    .Y(_0734_));
 sg13g2_nor2_1 _3256_ (.A(_0718_),
    .B(_0734_),
    .Y(_0735_));
 sg13g2_or2_1 _3257_ (.X(_0736_),
    .B(_0734_),
    .A(_0732_));
 sg13g2_xnor2_1 _3258_ (.Y(_0737_),
    .A(_0733_),
    .B(_0735_));
 sg13g2_nand2b_1 _3259_ (.Y(_0738_),
    .B(net684),
    .A_N(net746));
 sg13g2_a22oi_1 _3260_ (.Y(_0739_),
    .B1(_0738_),
    .B2(_0682_),
    .A2(_0737_),
    .A1(net604));
 sg13g2_a21o_1 _3261_ (.A2(net558),
    .A1(\mandelbrot.alu.m2[23] ),
    .B1(_0739_),
    .X(_0251_));
 sg13g2_o21ai_1 _3262_ (.B1(_0731_),
    .Y(_0740_),
    .A1(_0718_),
    .A2(_0736_));
 sg13g2_or4_2 _3263_ (.A(\mandelbrot.alu.in_zi[8] ),
    .B(\mandelbrot.alu.in_zi[9] ),
    .C(\mandelbrot.alu.in_zi[10] ),
    .D(_0700_),
    .X(_0741_));
 sg13g2_xnor2_1 _3264_ (.Y(_0742_),
    .A(\mandelbrot.alu.in_zi[10] ),
    .B(_0725_));
 sg13g2_nand2_1 _3265_ (.Y(_0743_),
    .A(net701),
    .B(_0742_));
 sg13g2_o21ai_1 _3266_ (.B1(_0743_),
    .Y(_0744_),
    .A1(net701),
    .A2(_0037_));
 sg13g2_nor2_1 _3267_ (.A(net642),
    .B(_0728_),
    .Y(_0745_));
 sg13g2_a21oi_1 _3268_ (.A1(net642),
    .A2(_0744_),
    .Y(_0746_),
    .B1(_0745_));
 sg13g2_xnor2_1 _3269_ (.Y(_0747_),
    .A(\mandelbrot.alu.m2[26] ),
    .B(_0746_));
 sg13g2_nand2b_1 _3270_ (.Y(_0748_),
    .B(_0747_),
    .A_N(_0740_));
 sg13g2_xnor2_1 _3271_ (.Y(_0749_),
    .A(_0740_),
    .B(_0747_));
 sg13g2_o21ai_1 _3272_ (.B1(net684),
    .Y(_0750_),
    .A1(net606),
    .A2(_0749_));
 sg13g2_a21oi_1 _3273_ (.A1(net463),
    .A2(net607),
    .Y(_0751_),
    .B1(_0750_));
 sg13g2_a21o_1 _3274_ (.A2(net558),
    .A1(\mandelbrot.alu.m2[24] ),
    .B1(_0751_),
    .X(_0252_));
 sg13g2_nand2_1 _3275_ (.Y(_0752_),
    .A(net700),
    .B(net558));
 sg13g2_or2_1 _3276_ (.X(_0753_),
    .B(_0036_),
    .A(net701));
 sg13g2_xnor2_1 _3277_ (.Y(_0754_),
    .A(\mandelbrot.alu.in_zi[11] ),
    .B(_0741_));
 sg13g2_o21ai_1 _3278_ (.B1(_0753_),
    .Y(_0755_),
    .A1(_1934_),
    .A2(_0754_));
 sg13g2_nand2b_1 _3279_ (.Y(_0756_),
    .B(net642),
    .A_N(_0755_));
 sg13g2_o21ai_1 _3280_ (.B1(_0756_),
    .Y(_0757_),
    .A1(net642),
    .A2(_0744_));
 sg13g2_nand2b_1 _3281_ (.Y(_0758_),
    .B(\mandelbrot.alu.m2[27] ),
    .A_N(_0757_));
 sg13g2_and2_1 _3282_ (.A(_1919_),
    .B(_0757_),
    .X(_0759_));
 sg13g2_xnor2_1 _3283_ (.Y(_0760_),
    .A(\mandelbrot.alu.m2[27] ),
    .B(_0757_));
 sg13g2_or2_1 _3284_ (.X(_0761_),
    .B(_0746_),
    .A(_0093_));
 sg13g2_and2_1 _3285_ (.A(_0748_),
    .B(_0761_),
    .X(_0762_));
 sg13g2_xnor2_1 _3286_ (.Y(_0763_),
    .A(_0760_),
    .B(_0762_));
 sg13g2_a21oi_1 _3287_ (.A1(_1919_),
    .A2(net607),
    .Y(_0764_),
    .B1(net267));
 sg13g2_o21ai_1 _3288_ (.B1(_0764_),
    .Y(_0765_),
    .A1(net606),
    .A2(_0763_));
 sg13g2_o21ai_1 _3289_ (.B1(_0752_),
    .Y(_0253_),
    .A1(net559),
    .A2(_0765_));
 sg13g2_o21ai_1 _3290_ (.B1(_0758_),
    .Y(_0766_),
    .A1(_0759_),
    .A2(_0761_));
 sg13g2_nand3b_1 _3291_ (.B(_0747_),
    .C(_0760_),
    .Y(_0767_),
    .A_N(_0740_));
 sg13g2_nand2b_1 _3292_ (.Y(_0768_),
    .B(_0767_),
    .A_N(_0766_));
 sg13g2_nor2_1 _3293_ (.A(net702),
    .B(_0035_),
    .Y(_0769_));
 sg13g2_nor3_2 _3294_ (.A(\mandelbrot.alu.in_zi[11] ),
    .B(\mandelbrot.alu.in_zi[12] ),
    .C(_0741_),
    .Y(_0770_));
 sg13g2_o21ai_1 _3295_ (.B1(\mandelbrot.alu.in_zi[12] ),
    .Y(_0771_),
    .A1(\mandelbrot.alu.in_zi[11] ),
    .A2(_0741_));
 sg13g2_nor2b_1 _3296_ (.A(_0770_),
    .B_N(_0771_),
    .Y(_0772_));
 sg13g2_a21oi_1 _3297_ (.A1(net702),
    .A2(_0772_),
    .Y(_0773_),
    .B1(_0769_));
 sg13g2_nand2_1 _3298_ (.Y(_0774_),
    .A(net641),
    .B(_0773_));
 sg13g2_o21ai_1 _3299_ (.B1(_0774_),
    .Y(_0775_),
    .A1(net642),
    .A2(_0755_));
 sg13g2_xnor2_1 _3300_ (.Y(_0776_),
    .A(\mandelbrot.alu.m2[28] ),
    .B(_0775_));
 sg13g2_xor2_1 _3301_ (.B(_0776_),
    .A(_0768_),
    .X(_0777_));
 sg13g2_o21ai_1 _3302_ (.B1(net684),
    .Y(_0778_),
    .A1(net606),
    .A2(_0777_));
 sg13g2_a21oi_1 _3303_ (.A1(net364),
    .A2(net606),
    .Y(_0779_),
    .B1(_0778_));
 sg13g2_a21o_1 _3304_ (.A2(net558),
    .A1(\mandelbrot.alu.m2[26] ),
    .B1(_0779_),
    .X(_0254_));
 sg13g2_nor2_1 _3305_ (.A(net702),
    .B(_0034_),
    .Y(_0780_));
 sg13g2_nand2b_1 _3306_ (.Y(_0781_),
    .B(_0770_),
    .A_N(\mandelbrot.alu.in_zi[13] ));
 sg13g2_xnor2_1 _3307_ (.Y(_0782_),
    .A(\mandelbrot.alu.in_zi[13] ),
    .B(_0770_));
 sg13g2_a21oi_1 _3308_ (.A1(net702),
    .A2(_0782_),
    .Y(_0783_),
    .B1(_0780_));
 sg13g2_nand2b_1 _3309_ (.Y(_0784_),
    .B(_0773_),
    .A_N(net642));
 sg13g2_nand2_1 _3310_ (.Y(_0785_),
    .A(net641),
    .B(_0783_));
 sg13g2_and3_1 _3311_ (.X(_0786_),
    .A(\mandelbrot.alu.m2[29] ),
    .B(_0784_),
    .C(_0785_));
 sg13g2_a21oi_1 _3312_ (.A1(_0784_),
    .A2(_0785_),
    .Y(_0787_),
    .B1(\mandelbrot.alu.m2[29] ));
 sg13g2_nor2_1 _3313_ (.A(_0786_),
    .B(_0787_),
    .Y(_0788_));
 sg13g2_nor2_1 _3314_ (.A(_0092_),
    .B(_0775_),
    .Y(_0789_));
 sg13g2_a21oi_1 _3315_ (.A1(_0768_),
    .A2(_0776_),
    .Y(_0790_),
    .B1(_0789_));
 sg13g2_or2_1 _3316_ (.X(_0791_),
    .B(_0790_),
    .A(_0788_));
 sg13g2_a21oi_1 _3317_ (.A1(_0788_),
    .A2(_0790_),
    .Y(_0792_),
    .B1(net606));
 sg13g2_a221oi_1 _3318_ (.B2(_0792_),
    .C1(_1910_),
    .B1(_0791_),
    .A1(net409),
    .Y(_0793_),
    .A2(net607));
 sg13g2_a21o_1 _3319_ (.A2(net558),
    .A1(\mandelbrot.alu.m2[27] ),
    .B1(_0793_),
    .X(_0255_));
 sg13g2_and2_1 _3320_ (.A(_0776_),
    .B(_0788_),
    .X(_0794_));
 sg13g2_a21o_1 _3321_ (.A2(_0789_),
    .A1(_0788_),
    .B1(_0786_),
    .X(_0795_));
 sg13g2_a21o_1 _3322_ (.A2(_0794_),
    .A1(_0768_),
    .B1(_0795_),
    .X(_0796_));
 sg13g2_nor2_1 _3323_ (.A(\mandelbrot.alu.in_zi[14] ),
    .B(_0781_),
    .Y(_0797_));
 sg13g2_xor2_1 _3324_ (.B(_0781_),
    .A(\mandelbrot.alu.in_zi[14] ),
    .X(_0798_));
 sg13g2_nand2_1 _3325_ (.Y(_0799_),
    .A(net701),
    .B(_0798_));
 sg13g2_o21ai_1 _3326_ (.B1(_0799_),
    .Y(_0800_),
    .A1(net701),
    .A2(_0033_));
 sg13g2_nor2_1 _3327_ (.A(net641),
    .B(_0783_),
    .Y(_0801_));
 sg13g2_a21oi_1 _3328_ (.A1(net641),
    .A2(_0800_),
    .Y(_0802_),
    .B1(_0801_));
 sg13g2_xnor2_1 _3329_ (.Y(_0803_),
    .A(\mandelbrot.alu.m2[30] ),
    .B(_0802_));
 sg13g2_xor2_1 _3330_ (.B(_0803_),
    .A(_0796_),
    .X(_0804_));
 sg13g2_nor2_1 _3331_ (.A(net606),
    .B(_0804_),
    .Y(_0805_));
 sg13g2_a21oi_1 _3332_ (.A1(net446),
    .A2(net606),
    .Y(_0806_),
    .B1(_0805_));
 sg13g2_a22oi_1 _3333_ (.Y(_0807_),
    .B1(_0806_),
    .B2(net684),
    .A2(net558),
    .A1(\mandelbrot.alu.m2[28] ));
 sg13g2_inv_1 _3334_ (.Y(_0256_),
    .A(_0807_));
 sg13g2_nor2_1 _3335_ (.A(_0090_),
    .B(_0802_),
    .Y(_0808_));
 sg13g2_a21oi_2 _3336_ (.B1(_0808_),
    .Y(_0809_),
    .A2(_0803_),
    .A1(_0796_));
 sg13g2_inv_1 _3337_ (.Y(_0810_),
    .A(_0809_));
 sg13g2_nor2b_1 _3338_ (.A(net701),
    .B_N(_0032_),
    .Y(_0811_));
 sg13g2_or2_1 _3339_ (.X(_0812_),
    .B(_0797_),
    .A(\mandelbrot.alu.in_zi[15] ));
 sg13g2_xnor2_1 _3340_ (.Y(_0813_),
    .A(\mandelbrot.alu.in_zi[15] ),
    .B(_0797_));
 sg13g2_nor2_1 _3341_ (.A(_1934_),
    .B(_0813_),
    .Y(_0814_));
 sg13g2_or2_1 _3342_ (.X(_0815_),
    .B(_0814_),
    .A(_0811_));
 sg13g2_nand2_1 _3343_ (.Y(_0816_),
    .A(net641),
    .B(_0815_));
 sg13g2_o21ai_1 _3344_ (.B1(_0816_),
    .Y(_0817_),
    .A1(net641),
    .A2(_0800_));
 sg13g2_xnor2_1 _3345_ (.Y(_0818_),
    .A(\mandelbrot.alu.m2[31] ),
    .B(_0817_));
 sg13g2_xor2_1 _3346_ (.B(_0818_),
    .A(_0809_),
    .X(_0819_));
 sg13g2_nand2b_1 _3347_ (.Y(_0820_),
    .B(net684),
    .A_N(net823));
 sg13g2_a22oi_1 _3348_ (.Y(_0821_),
    .B1(_0820_),
    .B2(_0682_),
    .A2(_0819_),
    .A1(net604));
 sg13g2_a21o_1 _3349_ (.A2(net558),
    .A1(\mandelbrot.alu.m2[29] ),
    .B1(_0821_),
    .X(_0257_));
 sg13g2_nor2_1 _3350_ (.A(_0105_),
    .B(_0817_),
    .Y(_0822_));
 sg13g2_a21oi_1 _3351_ (.A1(_0810_),
    .A2(_0818_),
    .Y(_0823_),
    .B1(_0822_));
 sg13g2_a21oi_2 _3352_ (.B1(_0811_),
    .Y(_0824_),
    .A2(_0812_),
    .A1(net702));
 sg13g2_nor2_1 _3353_ (.A(net641),
    .B(_0815_),
    .Y(_0825_));
 sg13g2_a21oi_1 _3354_ (.A1(net641),
    .A2(_0824_),
    .Y(_0826_),
    .B1(_0825_));
 sg13g2_nor2_1 _3355_ (.A(_0105_),
    .B(_0826_),
    .Y(_0827_));
 sg13g2_xnor2_1 _3356_ (.Y(_0828_),
    .A(_0105_),
    .B(_0826_));
 sg13g2_nor2_1 _3357_ (.A(_0823_),
    .B(_0828_),
    .Y(_0829_));
 sg13g2_xnor2_1 _3358_ (.Y(_0830_),
    .A(_0823_),
    .B(_0828_));
 sg13g2_a22oi_1 _3359_ (.Y(_0831_),
    .B1(_0830_),
    .B2(net604),
    .A2(_0820_),
    .A1(_0682_));
 sg13g2_a21o_1 _3360_ (.A2(net558),
    .A1(\mandelbrot.alu.m2[30] ),
    .B1(_0831_),
    .X(_0258_));
 sg13g2_nor2_1 _3361_ (.A(net681),
    .B(net580),
    .Y(_0832_));
 sg13g2_nor2_2 _3362_ (.A(_2161_),
    .B(net555),
    .Y(_0833_));
 sg13g2_nand3_1 _3363_ (.B(net206),
    .C(net611),
    .A(net682),
    .Y(_0834_));
 sg13g2_o21ai_1 _3364_ (.B1(_0834_),
    .Y(_0259_),
    .A1(_1915_),
    .A2(_0833_));
 sg13g2_a21oi_1 _3365_ (.A1(\mandelbrot.alu.mult_zr_zi.ctr[0] ),
    .A2(_0833_),
    .Y(_0835_),
    .B1(net227));
 sg13g2_nand2b_1 _3366_ (.Y(_0836_),
    .B(_0833_),
    .A_N(_0438_));
 sg13g2_a21oi_1 _3367_ (.A1(_0439_),
    .A2(_0833_),
    .Y(_0260_),
    .B1(net228));
 sg13g2_a22oi_1 _3368_ (.Y(_0261_),
    .B1(_0836_),
    .B2(_1971_),
    .A2(_0833_),
    .A1(_0440_));
 sg13g2_nor2_1 _3369_ (.A(net691),
    .B(net580),
    .Y(_0837_));
 sg13g2_nor2_2 _3370_ (.A(_2161_),
    .B(net548),
    .Y(_0838_));
 sg13g2_nand3_1 _3371_ (.B(net210),
    .C(net629),
    .A(net691),
    .Y(_0839_));
 sg13g2_o21ai_1 _3372_ (.B1(_0839_),
    .Y(_0262_),
    .A1(_1913_),
    .A2(_0838_));
 sg13g2_a21oi_1 _3373_ (.A1(\mandelbrot.alu.mult_zr_zr.ctr[0] ),
    .A2(_0838_),
    .Y(_0840_),
    .B1(net240));
 sg13g2_nand2b_1 _3374_ (.Y(_0841_),
    .B(_0838_),
    .A_N(_0429_));
 sg13g2_a21oi_1 _3375_ (.A1(_0430_),
    .A2(_0838_),
    .Y(_0263_),
    .B1(net241));
 sg13g2_a22oi_1 _3376_ (.Y(_0264_),
    .B1(_0841_),
    .B2(_1963_),
    .A2(_0838_),
    .A1(_0431_));
 sg13g2_a22oi_1 _3377_ (.Y(_0842_),
    .B1(net552),
    .B2(net400),
    .A2(net698),
    .A1(net681));
 sg13g2_inv_1 _3378_ (.Y(_0265_),
    .A(net401));
 sg13g2_xnor2_1 _3379_ (.Y(_0843_),
    .A(\mandelbrot.alu.m2[3] ),
    .B(\mandelbrot.alu.m1[3] ));
 sg13g2_nor2b_1 _3380_ (.A(net704),
    .B_N(net665),
    .Y(_0844_));
 sg13g2_nand2b_1 _3381_ (.Y(_0845_),
    .B(\mandelbrot.alu.m2[0] ),
    .A_N(\mandelbrot.alu.m1[0] ));
 sg13g2_xnor2_1 _3382_ (.Y(_0846_),
    .A(\mandelbrot.alu.m2[2] ),
    .B(\mandelbrot.alu.m1[2] ));
 sg13g2_o21ai_1 _3383_ (.B1(_0846_),
    .Y(_0847_),
    .A1(_1934_),
    .A2(net665));
 sg13g2_o21ai_1 _3384_ (.B1(_0843_),
    .Y(_0848_),
    .A1(_0844_),
    .A2(_0845_));
 sg13g2_nor2b_1 _3385_ (.A(\mandelbrot.alu.m2[2] ),
    .B_N(\mandelbrot.alu.m1[2] ),
    .Y(_0849_));
 sg13g2_nor2b_1 _3386_ (.A(\mandelbrot.alu.m2[3] ),
    .B_N(\mandelbrot.alu.m1[3] ),
    .Y(_0850_));
 sg13g2_a21oi_1 _3387_ (.A1(_0843_),
    .A2(_0849_),
    .Y(_0851_),
    .B1(_0850_));
 sg13g2_o21ai_1 _3388_ (.B1(_0851_),
    .Y(_0852_),
    .A1(_0847_),
    .A2(_0848_));
 sg13g2_nor2_1 _3389_ (.A(_2008_),
    .B(_2010_),
    .Y(_0853_));
 sg13g2_xor2_1 _3390_ (.B(\mandelbrot.alu.m1[4] ),
    .A(\mandelbrot.alu.m2[4] ),
    .X(_0854_));
 sg13g2_xor2_1 _3391_ (.B(\mandelbrot.alu.m1[5] ),
    .A(\mandelbrot.alu.m2[5] ),
    .X(_0855_));
 sg13g2_nor4_1 _3392_ (.A(_2008_),
    .B(_2010_),
    .C(_0854_),
    .D(_0855_),
    .Y(_0856_));
 sg13g2_nand2b_1 _3393_ (.Y(_0857_),
    .B(\mandelbrot.alu.m1[5] ),
    .A_N(\mandelbrot.alu.m2[5] ));
 sg13g2_nand2b_1 _3394_ (.Y(_0858_),
    .B(\mandelbrot.alu.m1[4] ),
    .A_N(\mandelbrot.alu.m2[4] ));
 sg13g2_o21ai_1 _3395_ (.B1(_0857_),
    .Y(_0859_),
    .A1(_0855_),
    .A2(_0858_));
 sg13g2_nand2b_1 _3396_ (.Y(_0860_),
    .B(\mandelbrot.alu.m1[6] ),
    .A_N(\mandelbrot.alu.m2[6] ));
 sg13g2_nand2b_1 _3397_ (.Y(_0861_),
    .B(\mandelbrot.alu.m1[7] ),
    .A_N(\mandelbrot.alu.m2[7] ));
 sg13g2_o21ai_1 _3398_ (.B1(_0861_),
    .Y(_0862_),
    .A1(_2008_),
    .A2(_0860_));
 sg13g2_a221oi_1 _3399_ (.B2(_0853_),
    .C1(_0862_),
    .B1(_0859_),
    .A1(_0852_),
    .Y(_0863_),
    .A2(_0856_));
 sg13g2_nor2_1 _3400_ (.A(_2017_),
    .B(_2018_),
    .Y(_0864_));
 sg13g2_nand3_1 _3401_ (.B(_2024_),
    .C(_0864_),
    .A(_2022_),
    .Y(_0865_));
 sg13g2_a21oi_1 _3402_ (.A1(_2021_),
    .A2(_2023_),
    .Y(_0866_),
    .B1(_2020_));
 sg13g2_o21ai_1 _3403_ (.B1(_2016_),
    .Y(_0867_),
    .A1(\mandelbrot.alu.m2[10] ),
    .A2(_1930_));
 sg13g2_a22oi_1 _3404_ (.Y(_0868_),
    .B1(_0867_),
    .B2(_2015_),
    .A2(_0866_),
    .A1(_0864_));
 sg13g2_o21ai_1 _3405_ (.B1(_0868_),
    .Y(_0869_),
    .A1(_0863_),
    .A2(_0865_));
 sg13g2_nor2_1 _3406_ (.A(_2032_),
    .B(_2033_),
    .Y(_0870_));
 sg13g2_a22oi_1 _3407_ (.Y(_0871_),
    .B1(_1928_),
    .B2(\mandelbrot.alu.m1[12] ),
    .A2(\mandelbrot.alu.m1[13] ),
    .A1(_1926_));
 sg13g2_a21oi_1 _3408_ (.A1(\mandelbrot.alu.m2[13] ),
    .A2(_1927_),
    .Y(_0872_),
    .B1(_0871_));
 sg13g2_a21oi_1 _3409_ (.A1(_0869_),
    .A2(_0870_),
    .Y(_0873_),
    .B1(_0872_));
 sg13g2_xor2_1 _3410_ (.B(_0873_),
    .A(_2040_),
    .X(_0874_));
 sg13g2_nand2_1 _3411_ (.Y(_0875_),
    .A(\mandelbrot.alu.in_cr[0] ),
    .B(_0874_));
 sg13g2_xnor2_1 _3412_ (.Y(_0876_),
    .A(\mandelbrot.alu.in_cr[0] ),
    .B(_0874_));
 sg13g2_nor2_2 _3413_ (.A(net675),
    .B(_0876_),
    .Y(_0877_));
 sg13g2_a22oi_1 _3414_ (.Y(_0878_),
    .B1(_0877_),
    .B2(net565),
    .A2(net555),
    .A1(\mandelbrot.alu.m3[0] ));
 sg13g2_o21ai_1 _3415_ (.B1(_0878_),
    .Y(_0266_),
    .A1(net655),
    .A2(_1972_));
 sg13g2_nand2b_1 _3416_ (.Y(_0879_),
    .B(\mandelbrot.alu.m1[14] ),
    .A_N(\mandelbrot.alu.m2[14] ));
 sg13g2_o21ai_1 _3417_ (.B1(_0879_),
    .Y(_0880_),
    .A1(_2040_),
    .A2(_0873_));
 sg13g2_xnor2_1 _3418_ (.Y(_0881_),
    .A(_2109_),
    .B(_0880_));
 sg13g2_nand2b_1 _3419_ (.Y(_0882_),
    .B(_0881_),
    .A_N(_0056_));
 sg13g2_xor2_1 _3420_ (.B(_0881_),
    .A(_0056_),
    .X(_0883_));
 sg13g2_xnor2_1 _3421_ (.Y(_0884_),
    .A(_0875_),
    .B(_0883_));
 sg13g2_nand2b_2 _3422_ (.Y(_0885_),
    .B(net661),
    .A_N(_0884_));
 sg13g2_nor2_1 _3423_ (.A(_0437_),
    .B(_0885_),
    .Y(_0886_));
 sg13g2_a221oi_1 _3424_ (.B2(net699),
    .C1(_0886_),
    .B1(net554),
    .A1(net682),
    .Y(_0887_),
    .A2(net708));
 sg13g2_inv_1 _3425_ (.Y(_0267_),
    .A(net709));
 sg13g2_o21ai_1 _3426_ (.B1(_0882_),
    .Y(_0888_),
    .A1(_0875_),
    .A2(_0883_));
 sg13g2_nand2_1 _3427_ (.Y(_0889_),
    .A(_1923_),
    .B(\mandelbrot.alu.m1[15] ));
 sg13g2_o21ai_1 _3428_ (.B1(_0889_),
    .Y(_0890_),
    .A1(_2109_),
    .A2(_0879_));
 sg13g2_nor2_1 _3429_ (.A(_2040_),
    .B(_2109_),
    .Y(_0891_));
 sg13g2_and2_1 _3430_ (.A(_0870_),
    .B(_0891_),
    .X(_0892_));
 sg13g2_a221oi_1 _3431_ (.B2(_0869_),
    .C1(_0890_),
    .B1(_0892_),
    .A1(_0872_),
    .Y(_0893_),
    .A2(_0891_));
 sg13g2_nor2_1 _3432_ (.A(_2049_),
    .B(_0893_),
    .Y(_0894_));
 sg13g2_xnor2_1 _3433_ (.Y(_0895_),
    .A(_2050_),
    .B(_0893_));
 sg13g2_and2_1 _3434_ (.A(\mandelbrot.alu.in_cr[2] ),
    .B(_0895_),
    .X(_0896_));
 sg13g2_xnor2_1 _3435_ (.Y(_0897_),
    .A(\mandelbrot.alu.in_cr[2] ),
    .B(_0895_));
 sg13g2_nor2b_1 _3436_ (.A(_0897_),
    .B_N(_0888_),
    .Y(_0898_));
 sg13g2_xor2_1 _3437_ (.B(_0897_),
    .A(_0888_),
    .X(_0899_));
 sg13g2_nor2_1 _3438_ (.A(net675),
    .B(_0899_),
    .Y(_0900_));
 sg13g2_a22oi_1 _3439_ (.Y(_0901_),
    .B1(_0900_),
    .B2(net565),
    .A2(net554),
    .A1(net233));
 sg13g2_o21ai_1 _3440_ (.B1(_0901_),
    .Y(_0268_),
    .A1(net655),
    .A2(_1973_));
 sg13g2_nor2_1 _3441_ (.A(_0896_),
    .B(_0898_),
    .Y(_0902_));
 sg13g2_nor2b_1 _3442_ (.A(\mandelbrot.alu.m2[16] ),
    .B_N(\mandelbrot.alu.m1[16] ),
    .Y(_0903_));
 sg13g2_nor2_1 _3443_ (.A(_0894_),
    .B(_0903_),
    .Y(_0904_));
 sg13g2_nand2_1 _3444_ (.Y(_0905_),
    .A(_2046_),
    .B(_2050_));
 sg13g2_xor2_1 _3445_ (.B(_0904_),
    .A(_2046_),
    .X(_0906_));
 sg13g2_nand2_1 _3446_ (.Y(_0907_),
    .A(_0055_),
    .B(_0906_));
 sg13g2_nor2_1 _3447_ (.A(_0055_),
    .B(_0906_),
    .Y(_0908_));
 sg13g2_xor2_1 _3448_ (.B(_0906_),
    .A(_0055_),
    .X(_0909_));
 sg13g2_xor2_1 _3449_ (.B(_0909_),
    .A(_0902_),
    .X(_0910_));
 sg13g2_nor2_2 _3450_ (.A(net678),
    .B(_0910_),
    .Y(_0911_));
 sg13g2_a22oi_1 _3451_ (.Y(_0912_),
    .B1(_0911_),
    .B2(_0436_),
    .A2(net553),
    .A1(\mandelbrot.alu.m3[3] ));
 sg13g2_o21ai_1 _3452_ (.B1(_0912_),
    .Y(_0269_),
    .A1(net656),
    .A2(_1974_));
 sg13g2_nand3b_1 _3453_ (.B(_0909_),
    .C(_0888_),
    .Y(_0913_),
    .A_N(_0897_));
 sg13g2_o21ai_1 _3454_ (.B1(_0907_),
    .Y(_0914_),
    .A1(_0896_),
    .A2(_0908_));
 sg13g2_and2_1 _3455_ (.A(_0913_),
    .B(_0914_),
    .X(_0915_));
 sg13g2_nor2_1 _3456_ (.A(\mandelbrot.alu.m2[17] ),
    .B(_1921_),
    .Y(_0916_));
 sg13g2_a21oi_1 _3457_ (.A1(_2046_),
    .A2(_0903_),
    .Y(_0917_),
    .B1(_0916_));
 sg13g2_o21ai_1 _3458_ (.B1(_0917_),
    .Y(_0918_),
    .A1(_0893_),
    .A2(_0905_));
 sg13g2_xnor2_1 _3459_ (.Y(_0919_),
    .A(_2101_),
    .B(_0918_));
 sg13g2_nand2_1 _3460_ (.Y(_0920_),
    .A(\mandelbrot.alu.in_cr[4] ),
    .B(_0919_));
 sg13g2_xnor2_1 _3461_ (.Y(_0921_),
    .A(\mandelbrot.alu.in_cr[4] ),
    .B(_0919_));
 sg13g2_inv_1 _3462_ (.Y(_0922_),
    .A(_0921_));
 sg13g2_nand2b_1 _3463_ (.Y(_0923_),
    .B(_0922_),
    .A_N(_0915_));
 sg13g2_xnor2_1 _3464_ (.Y(_0924_),
    .A(_0915_),
    .B(_0922_));
 sg13g2_nand2_1 _3465_ (.Y(_0925_),
    .A(net662),
    .B(_0924_));
 sg13g2_nor2_1 _3466_ (.A(net564),
    .B(_0925_),
    .Y(_0926_));
 sg13g2_a221oi_1 _3467_ (.B2(net255),
    .C1(_0926_),
    .B1(net553),
    .A1(net683),
    .Y(_0927_),
    .A2(net492));
 sg13g2_inv_1 _3468_ (.Y(_0270_),
    .A(net493));
 sg13g2_nor2b_1 _3469_ (.A(\mandelbrot.alu.m2[18] ),
    .B_N(\mandelbrot.alu.m1[18] ),
    .Y(_0928_));
 sg13g2_a21oi_1 _3470_ (.A1(_2102_),
    .A2(_0918_),
    .Y(_0929_),
    .B1(_0928_));
 sg13g2_xor2_1 _3471_ (.B(_0929_),
    .A(_2107_),
    .X(_0930_));
 sg13g2_nand2_1 _3472_ (.Y(_0931_),
    .A(_0054_),
    .B(_0930_));
 sg13g2_xor2_1 _3473_ (.B(_0930_),
    .A(_0054_),
    .X(_0932_));
 sg13g2_nand2_1 _3474_ (.Y(_0933_),
    .A(_0920_),
    .B(_0923_));
 sg13g2_xor2_1 _3475_ (.B(_0933_),
    .A(_0932_),
    .X(_0934_));
 sg13g2_nand2_1 _3476_ (.Y(_0935_),
    .A(net662),
    .B(_0934_));
 sg13g2_nor2_1 _3477_ (.A(net564),
    .B(_0935_),
    .Y(_0936_));
 sg13g2_a221oi_1 _3478_ (.B2(net243),
    .C1(_0936_),
    .B1(net553),
    .A1(net683),
    .Y(_0937_),
    .A2(net345));
 sg13g2_inv_1 _3479_ (.Y(_0271_),
    .A(_0937_));
 sg13g2_nand4_1 _3480_ (.B(_2050_),
    .C(_2102_),
    .A(_2046_),
    .Y(_0938_),
    .D(_2107_));
 sg13g2_nand2b_1 _3481_ (.Y(_0939_),
    .B(\mandelbrot.alu.m1[19] ),
    .A_N(\mandelbrot.alu.m2[19] ));
 sg13g2_nor2_1 _3482_ (.A(_2101_),
    .B(_0917_),
    .Y(_0940_));
 sg13g2_o21ai_1 _3483_ (.B1(_2107_),
    .Y(_0941_),
    .A1(_0928_),
    .A2(_0940_));
 sg13g2_and2_1 _3484_ (.A(_0939_),
    .B(_0941_),
    .X(_0942_));
 sg13g2_o21ai_1 _3485_ (.B1(_0942_),
    .Y(_0943_),
    .A1(_0893_),
    .A2(_0938_));
 sg13g2_xnor2_1 _3486_ (.Y(_0944_),
    .A(_2065_),
    .B(_0943_));
 sg13g2_and2_1 _3487_ (.A(\mandelbrot.alu.in_cr[6] ),
    .B(_0944_),
    .X(_0945_));
 sg13g2_xor2_1 _3488_ (.B(_0944_),
    .A(\mandelbrot.alu.in_cr[6] ),
    .X(_0946_));
 sg13g2_nor2b_1 _3489_ (.A(_0923_),
    .B_N(_0932_),
    .Y(_0947_));
 sg13g2_o21ai_1 _3490_ (.B1(_0920_),
    .Y(_0948_),
    .A1(_0054_),
    .A2(_0930_));
 sg13g2_a21o_1 _3491_ (.A2(_0948_),
    .A1(_0931_),
    .B1(_0947_),
    .X(_0949_));
 sg13g2_xnor2_1 _3492_ (.Y(_0950_),
    .A(_0946_),
    .B(_0949_));
 sg13g2_nand2b_1 _3493_ (.Y(_0951_),
    .B(net662),
    .A_N(_0950_));
 sg13g2_nor2_1 _3494_ (.A(net564),
    .B(_0951_),
    .Y(_0952_));
 sg13g2_a221oi_1 _3495_ (.B2(net492),
    .C1(_0952_),
    .B1(net553),
    .A1(net683),
    .Y(_0953_),
    .A2(net338));
 sg13g2_inv_1 _3496_ (.Y(_0272_),
    .A(_0953_));
 sg13g2_a21oi_1 _3497_ (.A1(_0946_),
    .A2(_0949_),
    .Y(_0954_),
    .B1(_0945_));
 sg13g2_nor2b_1 _3498_ (.A(\mandelbrot.alu.m2[20] ),
    .B_N(\mandelbrot.alu.m1[20] ),
    .Y(_0955_));
 sg13g2_a21oi_1 _3499_ (.A1(_2064_),
    .A2(_0943_),
    .Y(_0956_),
    .B1(_0955_));
 sg13g2_xnor2_1 _3500_ (.Y(_0957_),
    .A(_2062_),
    .B(_0956_));
 sg13g2_nand2_1 _3501_ (.Y(_0958_),
    .A(_1950_),
    .B(_0957_));
 sg13g2_xnor2_1 _3502_ (.Y(_0959_),
    .A(_0053_),
    .B(_0957_));
 sg13g2_xor2_1 _3503_ (.B(_0959_),
    .A(_0954_),
    .X(_0960_));
 sg13g2_nand2b_1 _3504_ (.Y(_0961_),
    .B(net662),
    .A_N(_0960_));
 sg13g2_a22oi_1 _3505_ (.Y(_0962_),
    .B1(net554),
    .B2(net345),
    .A2(\mandelbrot.alu.m3[9] ),
    .A1(net682));
 sg13g2_o21ai_1 _3506_ (.B1(net346),
    .Y(_0273_),
    .A1(net564),
    .A2(_0961_));
 sg13g2_o21ai_1 _3507_ (.B1(_0945_),
    .Y(_0963_),
    .A1(_1950_),
    .A2(_0957_));
 sg13g2_nand4_1 _3508_ (.B(_0946_),
    .C(_0948_),
    .A(_0931_),
    .Y(_0964_),
    .D(_0959_));
 sg13g2_nand3_1 _3509_ (.B(_0963_),
    .C(_0964_),
    .A(_0958_),
    .Y(_0965_));
 sg13g2_nand4_1 _3510_ (.B(_0932_),
    .C(_0946_),
    .A(_0922_),
    .Y(_0966_),
    .D(_0959_));
 sg13g2_a21oi_1 _3511_ (.A1(_0913_),
    .A2(_0914_),
    .Y(_0967_),
    .B1(_0966_));
 sg13g2_or2_1 _3512_ (.X(_0968_),
    .B(_0967_),
    .A(_0965_));
 sg13g2_inv_1 _3513_ (.Y(_0969_),
    .A(_0968_));
 sg13g2_and2_1 _3514_ (.A(_2062_),
    .B(_2064_),
    .X(_0970_));
 sg13g2_nor2b_1 _3515_ (.A(\mandelbrot.alu.m2[21] ),
    .B_N(\mandelbrot.alu.m1[21] ),
    .Y(_0971_));
 sg13g2_a21o_1 _3516_ (.A2(_0955_),
    .A1(_2062_),
    .B1(_0971_),
    .X(_0972_));
 sg13g2_a21o_1 _3517_ (.A2(_0970_),
    .A1(_0943_),
    .B1(_0972_),
    .X(_0973_));
 sg13g2_xor2_1 _3518_ (.B(_0973_),
    .A(_1992_),
    .X(_0974_));
 sg13g2_xnor2_1 _3519_ (.Y(_0975_),
    .A(\mandelbrot.alu.in_cr[8] ),
    .B(_0974_));
 sg13g2_xor2_1 _3520_ (.B(_0975_),
    .A(_0968_),
    .X(_0976_));
 sg13g2_nor2_2 _3521_ (.A(net678),
    .B(_0976_),
    .Y(_0977_));
 sg13g2_a22oi_1 _3522_ (.Y(_0978_),
    .B1(_0977_),
    .B2(net565),
    .A2(net553),
    .A1(net338));
 sg13g2_o21ai_1 _3523_ (.B1(_0978_),
    .Y(_0274_),
    .A1(net655),
    .A2(_1975_));
 sg13g2_nor2b_1 _3524_ (.A(\mandelbrot.alu.m2[22] ),
    .B_N(\mandelbrot.alu.m1[22] ),
    .Y(_0979_));
 sg13g2_a21oi_1 _3525_ (.A1(_1992_),
    .A2(_0973_),
    .Y(_0980_),
    .B1(_0979_));
 sg13g2_xor2_1 _3526_ (.B(_0980_),
    .A(_1990_),
    .X(_0981_));
 sg13g2_xnor2_1 _3527_ (.Y(_0982_),
    .A(_0051_),
    .B(_0981_));
 sg13g2_nand2b_1 _3528_ (.Y(_0983_),
    .B(_0974_),
    .A_N(_0052_));
 sg13g2_o21ai_1 _3529_ (.B1(_0983_),
    .Y(_0984_),
    .A1(_0969_),
    .A2(_0975_));
 sg13g2_xor2_1 _3530_ (.B(_0984_),
    .A(_0982_),
    .X(_0985_));
 sg13g2_nor2_2 _3531_ (.A(net678),
    .B(_0985_),
    .Y(_0986_));
 sg13g2_a22oi_1 _3532_ (.Y(_0987_),
    .B1(_0986_),
    .B2(net565),
    .A2(net553),
    .A1(\mandelbrot.alu.m3[9] ));
 sg13g2_o21ai_1 _3533_ (.B1(_0987_),
    .Y(_0275_),
    .A1(net655),
    .A2(_1976_));
 sg13g2_nor2b_1 _3534_ (.A(\mandelbrot.alu.m2[23] ),
    .B_N(\mandelbrot.alu.m1[23] ),
    .Y(_0988_));
 sg13g2_a21oi_1 _3535_ (.A1(_1990_),
    .A2(_0979_),
    .Y(_0989_),
    .B1(_0988_));
 sg13g2_inv_1 _3536_ (.Y(_0990_),
    .A(_0989_));
 sg13g2_a21oi_1 _3537_ (.A1(_1990_),
    .A2(_1992_),
    .Y(_0991_),
    .B1(_0990_));
 sg13g2_nand2b_1 _3538_ (.Y(_0992_),
    .B(_0989_),
    .A_N(_0972_));
 sg13g2_a21oi_1 _3539_ (.A1(_0943_),
    .A2(_0970_),
    .Y(_0993_),
    .B1(_0992_));
 sg13g2_nor2_1 _3540_ (.A(_0991_),
    .B(_0993_),
    .Y(_0994_));
 sg13g2_nor3_2 _3541_ (.A(_2073_),
    .B(_0991_),
    .C(_0993_),
    .Y(_0995_));
 sg13g2_xnor2_1 _3542_ (.Y(_0996_),
    .A(_2073_),
    .B(_0994_));
 sg13g2_nand2_1 _3543_ (.Y(_0997_),
    .A(\mandelbrot.alu.in_cr[10] ),
    .B(_0996_));
 sg13g2_nor2_1 _3544_ (.A(\mandelbrot.alu.in_cr[10] ),
    .B(_0996_),
    .Y(_0998_));
 sg13g2_xor2_1 _3545_ (.B(_0996_),
    .A(\mandelbrot.alu.in_cr[10] ),
    .X(_0999_));
 sg13g2_nor2_1 _3546_ (.A(_0975_),
    .B(_0982_),
    .Y(_1000_));
 sg13g2_o21ai_1 _3547_ (.B1(_1000_),
    .Y(_1001_),
    .A1(_0965_),
    .A2(_0967_));
 sg13g2_a21o_1 _3548_ (.A2(_0981_),
    .A1(_0051_),
    .B1(_0983_),
    .X(_1002_));
 sg13g2_o21ai_1 _3549_ (.B1(_1002_),
    .Y(_1003_),
    .A1(_0051_),
    .A2(_0981_));
 sg13g2_nor2b_1 _3550_ (.A(_1003_),
    .B_N(_1001_),
    .Y(_1004_));
 sg13g2_xnor2_1 _3551_ (.Y(_1005_),
    .A(_0999_),
    .B(_1004_));
 sg13g2_inv_1 _3552_ (.Y(_1006_),
    .A(_1005_));
 sg13g2_nand2_2 _3553_ (.Y(_1007_),
    .A(net662),
    .B(_1005_));
 sg13g2_nor2_1 _3554_ (.A(net564),
    .B(_1007_),
    .Y(_1008_));
 sg13g2_a221oi_1 _3555_ (.B2(net417),
    .C1(_1008_),
    .B1(net553),
    .A1(net682),
    .Y(_1009_),
    .A2(net369));
 sg13g2_inv_1 _3556_ (.Y(_0276_),
    .A(_1009_));
 sg13g2_o21ai_1 _3557_ (.B1(_0997_),
    .Y(_1010_),
    .A1(_0998_),
    .A2(_1004_));
 sg13g2_nor2b_1 _3558_ (.A(\mandelbrot.alu.m2[24] ),
    .B_N(\mandelbrot.alu.m1[24] ),
    .Y(_1011_));
 sg13g2_nor2_1 _3559_ (.A(_0995_),
    .B(_1011_),
    .Y(_1012_));
 sg13g2_o21ai_1 _3560_ (.B1(_2071_),
    .Y(_1013_),
    .A1(_0995_),
    .A2(_1011_));
 sg13g2_xnor2_1 _3561_ (.Y(_1014_),
    .A(_2070_),
    .B(_1012_));
 sg13g2_nor2_1 _3562_ (.A(_1949_),
    .B(_1014_),
    .Y(_1015_));
 sg13g2_xnor2_1 _3563_ (.Y(_1016_),
    .A(\mandelbrot.alu.in_cr[11] ),
    .B(_1014_));
 sg13g2_xnor2_1 _3564_ (.Y(_1017_),
    .A(_1010_),
    .B(_1016_));
 sg13g2_nor2_2 _3565_ (.A(net678),
    .B(_1017_),
    .Y(_1018_));
 sg13g2_a22oi_1 _3566_ (.Y(_1019_),
    .B1(_1018_),
    .B2(net565),
    .A2(net554),
    .A1(net300));
 sg13g2_o21ai_1 _3567_ (.B1(_1019_),
    .Y(_0277_),
    .A1(net655),
    .A2(_1956_));
 sg13g2_nand2b_1 _3568_ (.Y(_1020_),
    .B(\mandelbrot.alu.m1[25] ),
    .A_N(net700));
 sg13g2_a21o_1 _3569_ (.A2(_1020_),
    .A1(_1013_),
    .B1(_1986_),
    .X(_1021_));
 sg13g2_nand3_1 _3570_ (.B(_1013_),
    .C(_1020_),
    .A(_1986_),
    .Y(_1022_));
 sg13g2_and2_1 _3571_ (.A(_1021_),
    .B(_1022_),
    .X(_1023_));
 sg13g2_nand2_1 _3572_ (.Y(_1024_),
    .A(\mandelbrot.alu.in_cr[12] ),
    .B(_1023_));
 sg13g2_xnor2_1 _3573_ (.Y(_1025_),
    .A(\mandelbrot.alu.in_cr[12] ),
    .B(_1023_));
 sg13g2_a21oi_1 _3574_ (.A1(_1949_),
    .A2(_1014_),
    .Y(_1026_),
    .B1(_0997_));
 sg13g2_nor2_1 _3575_ (.A(_1015_),
    .B(_1026_),
    .Y(_1027_));
 sg13g2_nor3_1 _3576_ (.A(_1003_),
    .B(_1015_),
    .C(_1026_),
    .Y(_1028_));
 sg13g2_nand2_1 _3577_ (.Y(_1029_),
    .A(_0999_),
    .B(_1016_));
 sg13g2_nor2b_1 _3578_ (.A(_1029_),
    .B_N(_1003_),
    .Y(_1030_));
 sg13g2_nor4_1 _3579_ (.A(_0969_),
    .B(_0975_),
    .C(_0982_),
    .D(_1029_),
    .Y(_1031_));
 sg13g2_nor4_1 _3580_ (.A(_1015_),
    .B(_1026_),
    .C(_1030_),
    .D(_1031_),
    .Y(_1032_));
 sg13g2_a221oi_1 _3581_ (.B2(_1027_),
    .C1(_1025_),
    .B1(_1029_),
    .A1(_1001_),
    .Y(_1033_),
    .A2(_1028_));
 sg13g2_xor2_1 _3582_ (.B(_1032_),
    .A(_1025_),
    .X(_1034_));
 sg13g2_inv_1 _3583_ (.Y(_1035_),
    .A(_1034_));
 sg13g2_nor2_2 _3584_ (.A(net678),
    .B(_1035_),
    .Y(_1036_));
 sg13g2_a22oi_1 _3585_ (.Y(_1037_),
    .B1(_1036_),
    .B2(net565),
    .A2(net553),
    .A1(net369));
 sg13g2_o21ai_1 _3586_ (.B1(_1037_),
    .Y(_0278_),
    .A1(net655),
    .A2(_1955_));
 sg13g2_a21oi_1 _3587_ (.A1(\mandelbrot.alu.in_cr[12] ),
    .A2(_1023_),
    .Y(_1038_),
    .B1(_1033_));
 sg13g2_nor2b_1 _3588_ (.A(\mandelbrot.alu.m2[26] ),
    .B_N(\mandelbrot.alu.m1[26] ),
    .Y(_1039_));
 sg13g2_inv_1 _3589_ (.Y(_1040_),
    .A(_1039_));
 sg13g2_nand3_1 _3590_ (.B(_1021_),
    .C(_1040_),
    .A(_1984_),
    .Y(_1041_));
 sg13g2_a21o_1 _3591_ (.A2(_1040_),
    .A1(_1021_),
    .B1(_1984_),
    .X(_1042_));
 sg13g2_a21oi_1 _3592_ (.A1(_1041_),
    .A2(_1042_),
    .Y(_1043_),
    .B1(\mandelbrot.alu.in_cr[13] ));
 sg13g2_nand3_1 _3593_ (.B(_1041_),
    .C(_1042_),
    .A(\mandelbrot.alu.in_cr[13] ),
    .Y(_1044_));
 sg13g2_nor2b_1 _3594_ (.A(_1043_),
    .B_N(_1044_),
    .Y(_1045_));
 sg13g2_xnor2_1 _3595_ (.Y(_1046_),
    .A(_1038_),
    .B(_1045_));
 sg13g2_inv_1 _3596_ (.Y(_1047_),
    .A(_1046_));
 sg13g2_nor2_2 _3597_ (.A(net677),
    .B(_1047_),
    .Y(_1048_));
 sg13g2_a22oi_1 _3598_ (.Y(_1049_),
    .B1(_1048_),
    .B2(net565),
    .A2(net554),
    .A1(net371));
 sg13g2_o21ai_1 _3599_ (.B1(_1049_),
    .Y(_0279_),
    .A1(net655),
    .A2(_1954_));
 sg13g2_a21oi_1 _3600_ (.A1(_1024_),
    .A2(_1044_),
    .Y(_1050_),
    .B1(_1043_));
 sg13g2_a21oi_1 _3601_ (.A1(_1033_),
    .A2(_1045_),
    .Y(_1051_),
    .B1(_1050_));
 sg13g2_nor3_1 _3602_ (.A(_1984_),
    .B(_1986_),
    .C(_2070_),
    .Y(_1052_));
 sg13g2_nand2_1 _3603_ (.Y(_1053_),
    .A(_2071_),
    .B(_1011_));
 sg13g2_a21o_1 _3604_ (.A2(_1053_),
    .A1(_1020_),
    .B1(_1986_),
    .X(_1054_));
 sg13g2_a21oi_1 _3605_ (.A1(_1040_),
    .A2(_1054_),
    .Y(_1055_),
    .B1(_1984_));
 sg13g2_a221oi_1 _3606_ (.B2(_1052_),
    .C1(_1055_),
    .B1(_0995_),
    .A1(_1919_),
    .Y(_1056_),
    .A2(\mandelbrot.alu.m1[27] ));
 sg13g2_xor2_1 _3607_ (.B(_1056_),
    .A(_2086_),
    .X(_1057_));
 sg13g2_xnor2_1 _3608_ (.Y(_1058_),
    .A(\mandelbrot.alu.in_cr[14] ),
    .B(_1057_));
 sg13g2_xnor2_1 _3609_ (.Y(_1059_),
    .A(_1051_),
    .B(_1058_));
 sg13g2_nor2_2 _3610_ (.A(net679),
    .B(_1059_),
    .Y(_1060_));
 sg13g2_nor2_1 _3611_ (.A(net564),
    .B(_1060_),
    .Y(_1061_));
 sg13g2_a21o_1 _3612_ (.A2(\mandelbrot.alu.m3[0] ),
    .A1(\mandelbrot.alu.mult_zr_zi.shift_reg[0] ),
    .B1(net699),
    .X(_1062_));
 sg13g2_nor2_1 _3613_ (.A(\mandelbrot.alu.mult_zr_zi.shift_reg[0] ),
    .B(\mandelbrot.alu.m3[0] ),
    .Y(_1063_));
 sg13g2_o21ai_1 _3614_ (.B1(net699),
    .Y(_1064_),
    .A1(\mandelbrot.alu.mult_zr_zi.shift_reg[0] ),
    .A2(\mandelbrot.alu.m3[0] ));
 sg13g2_nand2_1 _3615_ (.Y(_1065_),
    .A(_1062_),
    .B(_1064_));
 sg13g2_nor2_1 _3616_ (.A(net698),
    .B(_1063_),
    .Y(_1066_));
 sg13g2_a21o_1 _3617_ (.A2(\mandelbrot.alu.m3[0] ),
    .A1(\mandelbrot.alu.mult_zr_zi.shift_reg[0] ),
    .B1(_1957_),
    .X(_1067_));
 sg13g2_nor2b_1 _3618_ (.A(_1066_),
    .B_N(_1067_),
    .Y(_1068_));
 sg13g2_nand2b_2 _3619_ (.Y(_1069_),
    .B(_1067_),
    .A_N(_1066_));
 sg13g2_nand3_1 _3620_ (.B(net640),
    .C(_1069_),
    .A(net671),
    .Y(_1070_));
 sg13g2_xor2_1 _3621_ (.B(_1070_),
    .A(\mandelbrot.alu.m3[16] ),
    .X(_1071_));
 sg13g2_a221oi_1 _3622_ (.B2(net682),
    .C1(_1061_),
    .B1(_1071_),
    .A1(_1955_),
    .Y(_0280_),
    .A2(net555));
 sg13g2_nand2b_1 _3623_ (.Y(_1072_),
    .B(\mandelbrot.alu.m1[28] ),
    .A_N(\mandelbrot.alu.m2[28] ));
 sg13g2_o21ai_1 _3624_ (.B1(_1072_),
    .Y(_1073_),
    .A1(_2086_),
    .A2(_1056_));
 sg13g2_xnor2_1 _3625_ (.Y(_1074_),
    .A(_2084_),
    .B(_1073_));
 sg13g2_nor2_1 _3626_ (.A(\mandelbrot.alu.in_cr[15] ),
    .B(_1074_),
    .Y(_1075_));
 sg13g2_inv_1 _3627_ (.Y(_1076_),
    .A(_1075_));
 sg13g2_nand2_1 _3628_ (.Y(_1077_),
    .A(\mandelbrot.alu.in_cr[15] ),
    .B(_1074_));
 sg13g2_nor2b_1 _3629_ (.A(_1075_),
    .B_N(_1077_),
    .Y(_1078_));
 sg13g2_nand2b_1 _3630_ (.Y(_1079_),
    .B(_1057_),
    .A_N(_0050_));
 sg13g2_o21ai_1 _3631_ (.B1(_1079_),
    .Y(_1080_),
    .A1(_1051_),
    .A2(_1058_));
 sg13g2_xnor2_1 _3632_ (.Y(_1081_),
    .A(_1078_),
    .B(_1080_));
 sg13g2_nor2_2 _3633_ (.A(net679),
    .B(_1081_),
    .Y(_1082_));
 sg13g2_nand3_1 _3634_ (.B(net671),
    .C(net640),
    .A(\mandelbrot.alu.m3[16] ),
    .Y(_1083_));
 sg13g2_nor2b_1 _3635_ (.A(\mandelbrot.alu.m3[1] ),
    .B_N(_0046_),
    .Y(_1084_));
 sg13g2_a221oi_1 _3636_ (.B2(_1064_),
    .C1(_1084_),
    .B1(_1062_),
    .A1(net699),
    .Y(_1085_),
    .A2(_0623_));
 sg13g2_and3_1 _3637_ (.X(_1086_),
    .A(_1969_),
    .B(_1062_),
    .C(_1064_));
 sg13g2_nor2_1 _3638_ (.A(_1085_),
    .B(_1086_),
    .Y(_1087_));
 sg13g2_o21ai_1 _3639_ (.B1(\mandelbrot.alu.m3[17] ),
    .Y(_1088_),
    .A1(_1085_),
    .A2(_1086_));
 sg13g2_nor3_1 _3640_ (.A(\mandelbrot.alu.m3[17] ),
    .B(_1085_),
    .C(_1086_),
    .Y(_1089_));
 sg13g2_xnor2_1 _3641_ (.Y(_1090_),
    .A(\mandelbrot.alu.m3[17] ),
    .B(_1087_));
 sg13g2_xor2_1 _3642_ (.B(_1090_),
    .A(_1083_),
    .X(_1091_));
 sg13g2_nand2_1 _3643_ (.Y(_1092_),
    .A(net600),
    .B(_1091_));
 sg13g2_o21ai_1 _3644_ (.B1(_1092_),
    .Y(_1093_),
    .A1(\mandelbrot.alu.m3[17] ),
    .A2(_1069_));
 sg13g2_a22oi_1 _3645_ (.Y(_1094_),
    .B1(_1082_),
    .B2(net565),
    .A2(net554),
    .A1(net380));
 sg13g2_o21ai_1 _3646_ (.B1(_1094_),
    .Y(_0281_),
    .A1(net656),
    .A2(_1093_));
 sg13g2_o21ai_1 _3647_ (.B1(_1088_),
    .Y(_1095_),
    .A1(_1083_),
    .A2(_1089_));
 sg13g2_mux2_1 _3648_ (.A0(_0045_),
    .A1(_0638_),
    .S(\mandelbrot.alu.m3[1] ),
    .X(_1096_));
 sg13g2_mux4_1 _3649_ (.S0(net640),
    .A0(_0046_),
    .A1(_0045_),
    .A2(_0623_),
    .A3(_0638_),
    .S1(net699),
    .X(_1097_));
 sg13g2_xnor2_1 _3650_ (.Y(_1098_),
    .A(\mandelbrot.alu.m3[18] ),
    .B(_1097_));
 sg13g2_xor2_1 _3651_ (.B(_1098_),
    .A(_1095_),
    .X(_1099_));
 sg13g2_o21ai_1 _3652_ (.B1(net682),
    .Y(_1100_),
    .A1(net603),
    .A2(_1099_));
 sg13g2_a21oi_1 _3653_ (.A1(net404),
    .A2(net603),
    .Y(_1101_),
    .B1(_1100_));
 sg13g2_a21o_1 _3654_ (.A2(net555),
    .A1(\mandelbrot.alu.m3[16] ),
    .B1(_1101_),
    .X(_0282_));
 sg13g2_nor2_1 _3655_ (.A(net698),
    .B(_0044_),
    .Y(_1102_));
 sg13g2_a21oi_1 _3656_ (.A1(net698),
    .A2(_0648_),
    .Y(_1103_),
    .B1(_1102_));
 sg13g2_mux2_1 _3657_ (.A0(_1096_),
    .A1(_1103_),
    .S(net640),
    .X(_1104_));
 sg13g2_nand2b_1 _3658_ (.Y(_1105_),
    .B(\mandelbrot.alu.m3[19] ),
    .A_N(_1104_));
 sg13g2_xor2_1 _3659_ (.B(_1104_),
    .A(\mandelbrot.alu.m3[19] ),
    .X(_1106_));
 sg13g2_nor2_1 _3660_ (.A(_0087_),
    .B(_1097_),
    .Y(_1107_));
 sg13g2_a21oi_1 _3661_ (.A1(_1095_),
    .A2(_1098_),
    .Y(_1108_),
    .B1(_1107_));
 sg13g2_xnor2_1 _3662_ (.Y(_1109_),
    .A(_1106_),
    .B(_1108_));
 sg13g2_nand2_1 _3663_ (.Y(_1110_),
    .A(_1069_),
    .B(_1109_));
 sg13g2_a21oi_1 _3664_ (.A1(net245),
    .A2(net603),
    .Y(_1111_),
    .B1(net656));
 sg13g2_a22oi_1 _3665_ (.Y(_1112_),
    .B1(_1110_),
    .B2(_1111_),
    .A2(net555),
    .A1(\mandelbrot.alu.m3[17] ));
 sg13g2_inv_1 _3666_ (.Y(_0283_),
    .A(net246));
 sg13g2_o21ai_1 _3667_ (.B1(_1105_),
    .Y(_1113_),
    .A1(_1106_),
    .A2(_1108_));
 sg13g2_nor2_1 _3668_ (.A(net699),
    .B(_0043_),
    .Y(_1114_));
 sg13g2_a21oi_1 _3669_ (.A1(net698),
    .A2(_0662_),
    .Y(_1115_),
    .B1(_1114_));
 sg13g2_mux2_1 _3670_ (.A0(_1103_),
    .A1(_1115_),
    .S(net640),
    .X(_1116_));
 sg13g2_inv_1 _3671_ (.Y(_1117_),
    .A(_1116_));
 sg13g2_xnor2_1 _3672_ (.Y(_1118_),
    .A(\mandelbrot.alu.m3[20] ),
    .B(_1116_));
 sg13g2_xor2_1 _3673_ (.B(_1118_),
    .A(_1113_),
    .X(_1119_));
 sg13g2_nor2_1 _3674_ (.A(net603),
    .B(_1119_),
    .Y(_1120_));
 sg13g2_a21oi_1 _3675_ (.A1(net290),
    .A2(net603),
    .Y(_1121_),
    .B1(_1120_));
 sg13g2_a22oi_1 _3676_ (.Y(_1122_),
    .B1(_1121_),
    .B2(net681),
    .A2(net552),
    .A1(\mandelbrot.alu.m3[18] ));
 sg13g2_inv_1 _3677_ (.Y(_0284_),
    .A(net291));
 sg13g2_a22oi_1 _3678_ (.Y(_1123_),
    .B1(_1118_),
    .B2(_1113_),
    .A2(_1117_),
    .A1(_1977_));
 sg13g2_or2_1 _3679_ (.X(_1124_),
    .B(_0042_),
    .A(net698));
 sg13g2_o21ai_1 _3680_ (.B1(_1124_),
    .Y(_1125_),
    .A1(_1957_),
    .A2(_0674_));
 sg13g2_nor2_1 _3681_ (.A(net640),
    .B(_1115_),
    .Y(_1126_));
 sg13g2_a21oi_1 _3682_ (.A1(net640),
    .A2(_1125_),
    .Y(_1127_),
    .B1(_1126_));
 sg13g2_nor2b_1 _3683_ (.A(_1127_),
    .B_N(\mandelbrot.alu.m3[21] ),
    .Y(_1128_));
 sg13g2_nor2b_1 _3684_ (.A(\mandelbrot.alu.m3[21] ),
    .B_N(_1127_),
    .Y(_1129_));
 sg13g2_nor2_1 _3685_ (.A(_1128_),
    .B(_1129_),
    .Y(_1130_));
 sg13g2_xor2_1 _3686_ (.B(_1130_),
    .A(_1123_),
    .X(_1131_));
 sg13g2_nand2_2 _3687_ (.Y(_1132_),
    .A(net680),
    .B(net600));
 sg13g2_nand2b_1 _3688_ (.Y(_1133_),
    .B(net681),
    .A_N(_0084_));
 sg13g2_a22oi_1 _3689_ (.Y(_1134_),
    .B1(_1132_),
    .B2(_1133_),
    .A2(_1131_),
    .A1(net600));
 sg13g2_a21o_1 _3690_ (.A2(net552),
    .A1(net529),
    .B1(_1134_),
    .X(_0285_));
 sg13g2_a221oi_1 _3691_ (.B2(_1113_),
    .C1(_1128_),
    .B1(_1118_),
    .A1(_1977_),
    .Y(_1135_),
    .A2(_1117_));
 sg13g2_nor2_1 _3692_ (.A(net698),
    .B(_0041_),
    .Y(_1136_));
 sg13g2_a21oi_1 _3693_ (.A1(net698),
    .A2(_0688_),
    .Y(_1137_),
    .B1(_1136_));
 sg13g2_nand2_1 _3694_ (.Y(_1138_),
    .A(net639),
    .B(_1137_));
 sg13g2_o21ai_1 _3695_ (.B1(_1138_),
    .Y(_1139_),
    .A1(net639),
    .A2(_1125_));
 sg13g2_xor2_1 _3696_ (.B(_1139_),
    .A(\mandelbrot.alu.m3[22] ),
    .X(_1140_));
 sg13g2_or3_1 _3697_ (.A(_1129_),
    .B(_1135_),
    .C(_1140_),
    .X(_1141_));
 sg13g2_o21ai_1 _3698_ (.B1(_1140_),
    .Y(_1142_),
    .A1(_1129_),
    .A2(_1135_));
 sg13g2_a21oi_1 _3699_ (.A1(_1141_),
    .A2(_1142_),
    .Y(_1143_),
    .B1(net603));
 sg13g2_a21oi_1 _3700_ (.A1(_0083_),
    .A2(net603),
    .Y(_1144_),
    .B1(_1143_));
 sg13g2_a22oi_1 _3701_ (.Y(_1145_),
    .B1(_1144_),
    .B2(net681),
    .A2(net552),
    .A1(net435));
 sg13g2_inv_1 _3702_ (.Y(_0286_),
    .A(net436));
 sg13g2_nor2_1 _3703_ (.A(net697),
    .B(_0040_),
    .Y(_1146_));
 sg13g2_a21oi_1 _3704_ (.A1(net697),
    .A2(_0701_),
    .Y(_1147_),
    .B1(_1146_));
 sg13g2_mux2_1 _3705_ (.A0(_1137_),
    .A1(_1147_),
    .S(net639),
    .X(_1148_));
 sg13g2_nand2b_1 _3706_ (.Y(_1149_),
    .B(\mandelbrot.alu.m3[23] ),
    .A_N(_1148_));
 sg13g2_xnor2_1 _3707_ (.Y(_1150_),
    .A(\mandelbrot.alu.m3[23] ),
    .B(_1148_));
 sg13g2_inv_1 _3708_ (.Y(_1151_),
    .A(_1150_));
 sg13g2_nor2_1 _3709_ (.A(_0083_),
    .B(_1139_),
    .Y(_1152_));
 sg13g2_inv_1 _3710_ (.Y(_1153_),
    .A(_1152_));
 sg13g2_nand3_1 _3711_ (.B(_1151_),
    .C(_1153_),
    .A(_1141_),
    .Y(_1154_));
 sg13g2_a21o_1 _3712_ (.A2(_1153_),
    .A1(_1141_),
    .B1(_1151_),
    .X(_1155_));
 sg13g2_a21o_1 _3713_ (.A2(_1155_),
    .A1(_1154_),
    .B1(net602),
    .X(_1156_));
 sg13g2_o21ai_1 _3714_ (.B1(_1156_),
    .Y(_1157_),
    .A1(\mandelbrot.alu.m3[23] ),
    .A2(net600));
 sg13g2_nor3_1 _3715_ (.A(_0075_),
    .B(net550),
    .C(_1157_),
    .Y(_1158_));
 sg13g2_a21o_1 _3716_ (.A2(net552),
    .A1(net501),
    .B1(_1158_),
    .X(_0287_));
 sg13g2_nand2_1 _3717_ (.Y(_1159_),
    .A(_1149_),
    .B(_1155_));
 sg13g2_or2_1 _3718_ (.X(_1160_),
    .B(_0039_),
    .A(net696));
 sg13g2_o21ai_1 _3719_ (.B1(_1160_),
    .Y(_1161_),
    .A1(_1957_),
    .A2(_0713_));
 sg13g2_nor2_1 _3720_ (.A(net639),
    .B(_1147_),
    .Y(_1162_));
 sg13g2_a21oi_1 _3721_ (.A1(net639),
    .A2(_1161_),
    .Y(_1163_),
    .B1(_1162_));
 sg13g2_xnor2_1 _3722_ (.Y(_1164_),
    .A(\mandelbrot.alu.m3[24] ),
    .B(_1163_));
 sg13g2_inv_1 _3723_ (.Y(_1165_),
    .A(_1164_));
 sg13g2_a21o_1 _3724_ (.A2(_1155_),
    .A1(_1149_),
    .B1(_1165_),
    .X(_1166_));
 sg13g2_xnor2_1 _3725_ (.Y(_1167_),
    .A(_1159_),
    .B(_1165_));
 sg13g2_o21ai_1 _3726_ (.B1(net680),
    .Y(_1168_),
    .A1(net602),
    .A2(_1167_));
 sg13g2_a21oi_1 _3727_ (.A1(net415),
    .A2(net602),
    .Y(_1169_),
    .B1(_1168_));
 sg13g2_a21o_1 _3728_ (.A2(net551),
    .A1(\mandelbrot.alu.m3[22] ),
    .B1(_1169_),
    .X(_0288_));
 sg13g2_nor2_1 _3729_ (.A(net696),
    .B(_0038_),
    .Y(_1170_));
 sg13g2_a21oi_1 _3730_ (.A1(net696),
    .A2(_0727_),
    .Y(_1171_),
    .B1(_1170_));
 sg13g2_nand2_1 _3731_ (.Y(_1172_),
    .A(net638),
    .B(_1171_));
 sg13g2_o21ai_1 _3732_ (.B1(_1172_),
    .Y(_1173_),
    .A1(net638),
    .A2(_1161_));
 sg13g2_and2_1 _3733_ (.A(_1952_),
    .B(_1173_),
    .X(_1174_));
 sg13g2_nor2_1 _3734_ (.A(_1952_),
    .B(_1173_),
    .Y(_1175_));
 sg13g2_nor2_1 _3735_ (.A(_1174_),
    .B(_1175_),
    .Y(_1176_));
 sg13g2_nor2_1 _3736_ (.A(_0082_),
    .B(_1163_),
    .Y(_1177_));
 sg13g2_a21oi_1 _3737_ (.A1(_1159_),
    .A2(_1164_),
    .Y(_1178_),
    .B1(_1177_));
 sg13g2_nor2_1 _3738_ (.A(_1175_),
    .B(_1177_),
    .Y(_1179_));
 sg13g2_xor2_1 _3739_ (.B(_1178_),
    .A(_1176_),
    .X(_1180_));
 sg13g2_nand2b_1 _3740_ (.Y(_1181_),
    .B(net680),
    .A_N(_0081_));
 sg13g2_a22oi_1 _3741_ (.Y(_1182_),
    .B1(_1181_),
    .B2(_1132_),
    .A2(_1180_),
    .A1(net600));
 sg13g2_a21o_1 _3742_ (.A2(net550),
    .A1(net753),
    .B1(_1182_),
    .X(_0289_));
 sg13g2_a21o_1 _3743_ (.A2(_1179_),
    .A1(_1166_),
    .B1(_1174_),
    .X(_1183_));
 sg13g2_nand2_1 _3744_ (.Y(_1184_),
    .A(net695),
    .B(_0742_));
 sg13g2_o21ai_1 _3745_ (.B1(_1184_),
    .Y(_1185_),
    .A1(net695),
    .A2(_0037_));
 sg13g2_nor2_1 _3746_ (.A(net638),
    .B(_1171_),
    .Y(_1186_));
 sg13g2_a21oi_2 _3747_ (.B1(_1186_),
    .Y(_1187_),
    .A2(_1185_),
    .A1(net638));
 sg13g2_xnor2_1 _3748_ (.Y(_1188_),
    .A(\mandelbrot.alu.m3[26] ),
    .B(_1187_));
 sg13g2_nand2b_1 _3749_ (.Y(_1189_),
    .B(_1188_),
    .A_N(_1183_));
 sg13g2_xnor2_1 _3750_ (.Y(_1190_),
    .A(_1183_),
    .B(_1188_));
 sg13g2_o21ai_1 _3751_ (.B1(net680),
    .Y(_1191_),
    .A1(net601),
    .A2(_1190_));
 sg13g2_a21oi_1 _3752_ (.A1(net413),
    .A2(net601),
    .Y(_1192_),
    .B1(_1191_));
 sg13g2_a21o_1 _3753_ (.A2(net550),
    .A1(\mandelbrot.alu.m3[24] ),
    .B1(_1192_),
    .X(_0290_));
 sg13g2_or2_1 _3754_ (.X(_1193_),
    .B(_0036_),
    .A(net695));
 sg13g2_o21ai_1 _3755_ (.B1(_1193_),
    .Y(_1194_),
    .A1(_1957_),
    .A2(_0754_));
 sg13g2_nand2b_1 _3756_ (.Y(_1195_),
    .B(net636),
    .A_N(_1194_));
 sg13g2_o21ai_1 _3757_ (.B1(_1195_),
    .Y(_1196_),
    .A1(net638),
    .A2(_1185_));
 sg13g2_nand2b_1 _3758_ (.Y(_1197_),
    .B(\mandelbrot.alu.m3[27] ),
    .A_N(_1196_));
 sg13g2_nor2b_1 _3759_ (.A(\mandelbrot.alu.m3[27] ),
    .B_N(_1196_),
    .Y(_1198_));
 sg13g2_xnor2_1 _3760_ (.Y(_1199_),
    .A(\mandelbrot.alu.m3[27] ),
    .B(_1196_));
 sg13g2_or2_1 _3761_ (.X(_1200_),
    .B(_1187_),
    .A(_0080_));
 sg13g2_and2_1 _3762_ (.A(_1189_),
    .B(_1200_),
    .X(_1201_));
 sg13g2_a21oi_1 _3763_ (.A1(_1199_),
    .A2(_1201_),
    .Y(_1202_),
    .B1(net601));
 sg13g2_o21ai_1 _3764_ (.B1(_1202_),
    .Y(_1203_),
    .A1(_1199_),
    .A2(_1201_));
 sg13g2_o21ai_1 _3765_ (.B1(_1203_),
    .Y(_1204_),
    .A1(\mandelbrot.alu.m3[27] ),
    .A2(net600));
 sg13g2_nor3_1 _3766_ (.A(_0075_),
    .B(net550),
    .C(_1204_),
    .Y(_1205_));
 sg13g2_a21o_1 _3767_ (.A2(net550),
    .A1(net474),
    .B1(_1205_),
    .X(_0291_));
 sg13g2_o21ai_1 _3768_ (.B1(_1197_),
    .Y(_1206_),
    .A1(_1198_),
    .A2(_1200_));
 sg13g2_nand2_1 _3769_ (.Y(_1207_),
    .A(_1188_),
    .B(_1199_));
 sg13g2_a221oi_1 _3770_ (.B2(_1166_),
    .C1(_1207_),
    .B1(_1179_),
    .A1(_1952_),
    .Y(_1208_),
    .A2(_1173_));
 sg13g2_nor2_1 _3771_ (.A(_1206_),
    .B(_1208_),
    .Y(_1209_));
 sg13g2_nor2_1 _3772_ (.A(net694),
    .B(_0035_),
    .Y(_1210_));
 sg13g2_a21oi_1 _3773_ (.A1(net694),
    .A2(_0772_),
    .Y(_1211_),
    .B1(_1210_));
 sg13g2_nand2_1 _3774_ (.Y(_1212_),
    .A(net637),
    .B(_1211_));
 sg13g2_o21ai_1 _3775_ (.B1(_1212_),
    .Y(_1213_),
    .A1(net636),
    .A2(_1194_));
 sg13g2_xnor2_1 _3776_ (.Y(_1214_),
    .A(\mandelbrot.alu.m3[28] ),
    .B(_1213_));
 sg13g2_o21ai_1 _3777_ (.B1(_1214_),
    .Y(_1215_),
    .A1(_1206_),
    .A2(_1208_));
 sg13g2_xnor2_1 _3778_ (.Y(_1216_),
    .A(_1209_),
    .B(_1214_));
 sg13g2_o21ai_1 _3779_ (.B1(net680),
    .Y(_1217_),
    .A1(net601),
    .A2(_1216_));
 sg13g2_a21oi_1 _3780_ (.A1(net386),
    .A2(net601),
    .Y(_1218_),
    .B1(_1217_));
 sg13g2_a21o_1 _3781_ (.A2(net550),
    .A1(\mandelbrot.alu.m3[26] ),
    .B1(_1218_),
    .X(_0292_));
 sg13g2_nand2_1 _3782_ (.Y(_1219_),
    .A(\mandelbrot.alu.m3[27] ),
    .B(net550));
 sg13g2_or2_1 _3783_ (.X(_1220_),
    .B(_1213_),
    .A(_0079_));
 sg13g2_nor2_1 _3784_ (.A(net694),
    .B(_0034_),
    .Y(_1221_));
 sg13g2_a21oi_1 _3785_ (.A1(net694),
    .A2(_0782_),
    .Y(_1222_),
    .B1(_1221_));
 sg13g2_nand2b_1 _3786_ (.Y(_1223_),
    .B(_1211_),
    .A_N(net636));
 sg13g2_nand2_1 _3787_ (.Y(_1224_),
    .A(net636),
    .B(_1222_));
 sg13g2_a21oi_2 _3788_ (.B1(\mandelbrot.alu.m3[29] ),
    .Y(_1225_),
    .A2(_1224_),
    .A1(_1223_));
 sg13g2_nand3_1 _3789_ (.B(_1223_),
    .C(_1224_),
    .A(\mandelbrot.alu.m3[29] ),
    .Y(_1226_));
 sg13g2_nor2b_1 _3790_ (.A(_1225_),
    .B_N(_1226_),
    .Y(_1227_));
 sg13g2_a21oi_1 _3791_ (.A1(_1215_),
    .A2(_1220_),
    .Y(_1228_),
    .B1(_1227_));
 sg13g2_and3_1 _3792_ (.X(_1229_),
    .A(_1215_),
    .B(_1220_),
    .C(_1226_));
 sg13g2_nor2b_1 _3793_ (.A(_1225_),
    .B_N(_1229_),
    .Y(_1230_));
 sg13g2_nor3_1 _3794_ (.A(net601),
    .B(_1228_),
    .C(_1230_),
    .Y(_1231_));
 sg13g2_a21o_1 _3795_ (.A2(net601),
    .A1(net329),
    .B1(net656),
    .X(_1232_));
 sg13g2_o21ai_1 _3796_ (.B1(_1219_),
    .Y(_0293_),
    .A1(_1231_),
    .A2(_1232_));
 sg13g2_nand2_1 _3797_ (.Y(_1233_),
    .A(net694),
    .B(_0798_));
 sg13g2_o21ai_1 _3798_ (.B1(_1233_),
    .Y(_1234_),
    .A1(net694),
    .A2(_0033_));
 sg13g2_nor2_1 _3799_ (.A(net636),
    .B(_1222_),
    .Y(_1235_));
 sg13g2_a21oi_1 _3800_ (.A1(net636),
    .A2(_1234_),
    .Y(_1236_),
    .B1(_1235_));
 sg13g2_xor2_1 _3801_ (.B(_1236_),
    .A(\mandelbrot.alu.m3[30] ),
    .X(_1237_));
 sg13g2_nor3_1 _3802_ (.A(_1225_),
    .B(_1229_),
    .C(_1237_),
    .Y(_1238_));
 sg13g2_o21ai_1 _3803_ (.B1(_1237_),
    .Y(_1239_),
    .A1(_1225_),
    .A2(_1229_));
 sg13g2_nor2b_1 _3804_ (.A(_1238_),
    .B_N(_1239_),
    .Y(_1240_));
 sg13g2_nor2_1 _3805_ (.A(net601),
    .B(_1240_),
    .Y(_1241_));
 sg13g2_a21oi_1 _3806_ (.A1(net425),
    .A2(net602),
    .Y(_1242_),
    .B1(_1241_));
 sg13g2_a22oi_1 _3807_ (.Y(_1243_),
    .B1(_1242_),
    .B2(net680),
    .A2(net550),
    .A1(\mandelbrot.alu.m3[28] ));
 sg13g2_inv_1 _3808_ (.Y(_0294_),
    .A(net426));
 sg13g2_nor2_1 _3809_ (.A(_0104_),
    .B(_1236_),
    .Y(_1244_));
 sg13g2_nor2_1 _3810_ (.A(_1238_),
    .B(_1244_),
    .Y(_1245_));
 sg13g2_nor2b_1 _3811_ (.A(net694),
    .B_N(_0032_),
    .Y(_1246_));
 sg13g2_nor2_1 _3812_ (.A(_1957_),
    .B(_0813_),
    .Y(_1247_));
 sg13g2_or2_1 _3813_ (.X(_1248_),
    .B(_1247_),
    .A(_1246_));
 sg13g2_nand2_1 _3814_ (.Y(_1249_),
    .A(net637),
    .B(_1248_));
 sg13g2_o21ai_1 _3815_ (.B1(_1249_),
    .Y(_1250_),
    .A1(net636),
    .A2(_1234_));
 sg13g2_xnor2_1 _3816_ (.Y(_1251_),
    .A(\mandelbrot.alu.m3[31] ),
    .B(_1250_));
 sg13g2_nor2b_1 _3817_ (.A(_1245_),
    .B_N(_1251_),
    .Y(_1252_));
 sg13g2_xor2_1 _3818_ (.B(_1251_),
    .A(_1245_),
    .X(_1253_));
 sg13g2_nand2b_1 _3819_ (.Y(_1254_),
    .B(net680),
    .A_N(_0030_));
 sg13g2_a22oi_1 _3820_ (.Y(_1255_),
    .B1(_1254_),
    .B2(_1132_),
    .A2(_1253_),
    .A1(net600));
 sg13g2_a21o_1 _3821_ (.A2(net551),
    .A1(net739),
    .B1(_1255_),
    .X(_0295_));
 sg13g2_nor2_1 _3822_ (.A(_0030_),
    .B(_1250_),
    .Y(_1256_));
 sg13g2_nor2_1 _3823_ (.A(_1252_),
    .B(_1256_),
    .Y(_1257_));
 sg13g2_a21oi_2 _3824_ (.B1(_1246_),
    .Y(_1258_),
    .A2(_0812_),
    .A1(net694));
 sg13g2_nor2_1 _3825_ (.A(net637),
    .B(_1248_),
    .Y(_1259_));
 sg13g2_a21oi_2 _3826_ (.B1(_1259_),
    .Y(_1260_),
    .A2(_1258_),
    .A1(net636));
 sg13g2_or2_1 _3827_ (.X(_1261_),
    .B(_1260_),
    .A(_0030_));
 sg13g2_xnor2_1 _3828_ (.Y(_1262_),
    .A(_0030_),
    .B(_1260_));
 sg13g2_xnor2_1 _3829_ (.Y(_1263_),
    .A(_1257_),
    .B(_1262_));
 sg13g2_a22oi_1 _3830_ (.Y(_1264_),
    .B1(_1263_),
    .B2(net600),
    .A2(_1254_),
    .A1(_1132_));
 sg13g2_a21o_1 _3831_ (.A2(net551),
    .A1(net515),
    .B1(_1264_),
    .X(_0296_));
 sg13g2_nor2_2 _3832_ (.A(_2161_),
    .B(net562),
    .Y(_1265_));
 sg13g2_nand3_1 _3833_ (.B(net214),
    .C(net620),
    .A(net688),
    .Y(_1266_));
 sg13g2_o21ai_1 _3834_ (.B1(net215),
    .Y(_0297_),
    .A1(_1914_),
    .A2(_1265_));
 sg13g2_a21oi_1 _3835_ (.A1(\mandelbrot.alu.mult_zi_zi.ctr[0] ),
    .A2(_1265_),
    .Y(_1267_),
    .B1(net235));
 sg13g2_nand2b_1 _3836_ (.Y(_1268_),
    .B(_1265_),
    .A_N(_0433_));
 sg13g2_a21oi_1 _3837_ (.A1(_0434_),
    .A2(_1265_),
    .Y(_0298_),
    .B1(net236));
 sg13g2_a22oi_1 _3838_ (.Y(_0299_),
    .B1(_1268_),
    .B2(_1968_),
    .A2(_1265_),
    .A1(_0435_));
 sg13g2_xor2_1 _3839_ (.B(_0824_),
    .A(net817),
    .X(_1269_));
 sg13g2_o21ai_1 _3840_ (.B1(_1269_),
    .Y(_1270_),
    .A1(_0827_),
    .A2(_0829_));
 sg13g2_nor3_1 _3841_ (.A(_0827_),
    .B(_0829_),
    .C(_1269_),
    .Y(_1271_));
 sg13g2_nor2_1 _3842_ (.A(_0682_),
    .B(_1271_),
    .Y(_1272_));
 sg13g2_nand2_1 _3843_ (.Y(_1273_),
    .A(\mandelbrot.alu.m2[31] ),
    .B(_0432_));
 sg13g2_a22oi_1 _3844_ (.Y(_0300_),
    .B1(_1273_),
    .B2(_0682_),
    .A2(_1272_),
    .A1(net818));
 sg13g2_a21oi_2 _3845_ (.B1(_2161_),
    .Y(_1274_),
    .A2(_1918_),
    .A1(net677));
 sg13g2_o21ai_1 _3846_ (.B1(_1274_),
    .Y(_1275_),
    .A1(net677),
    .A2(_2155_));
 sg13g2_nand2_1 _3847_ (.Y(_1276_),
    .A(net772),
    .B(net587));
 sg13g2_and3_1 _3848_ (.X(_1277_),
    .A(_2155_),
    .B(_0425_),
    .C(_1274_));
 sg13g2_nand3_1 _3849_ (.B(_0425_),
    .C(_1274_),
    .A(_2155_),
    .Y(_1278_));
 sg13g2_o21ai_1 _3850_ (.B1(_1276_),
    .Y(_0301_),
    .A1(_0876_),
    .A2(net576));
 sg13g2_nand2_1 _3851_ (.Y(_1279_),
    .A(net491),
    .B(net587));
 sg13g2_o21ai_1 _3852_ (.B1(_1279_),
    .Y(_0302_),
    .A1(_0884_),
    .A2(net576));
 sg13g2_nand2_1 _3853_ (.Y(_1280_),
    .A(net374),
    .B(net591));
 sg13g2_o21ai_1 _3854_ (.B1(_1280_),
    .Y(_0303_),
    .A1(_0899_),
    .A2(net579));
 sg13g2_nand2_1 _3855_ (.Y(_1281_),
    .A(net331),
    .B(net591));
 sg13g2_o21ai_1 _3856_ (.B1(_1281_),
    .Y(_0304_),
    .A1(_0910_),
    .A2(net579));
 sg13g2_a22oi_1 _3857_ (.Y(_1282_),
    .B1(_1277_),
    .B2(_0924_),
    .A2(net591),
    .A1(net497));
 sg13g2_inv_1 _3858_ (.Y(_0305_),
    .A(net498));
 sg13g2_and2_1 _3859_ (.A(net773),
    .B(net591),
    .X(_1283_));
 sg13g2_a21o_1 _3860_ (.A2(_1277_),
    .A1(_0934_),
    .B1(_1283_),
    .X(_0306_));
 sg13g2_nand2_1 _3861_ (.Y(_1284_),
    .A(net279),
    .B(net591));
 sg13g2_o21ai_1 _3862_ (.B1(_1284_),
    .Y(_0307_),
    .A1(_0950_),
    .A2(net579));
 sg13g2_nand2_1 _3863_ (.Y(_1285_),
    .A(net296),
    .B(net591));
 sg13g2_o21ai_1 _3864_ (.B1(_1285_),
    .Y(_0308_),
    .A1(_0960_),
    .A2(net579));
 sg13g2_nand2_1 _3865_ (.Y(_1286_),
    .A(net427),
    .B(net591));
 sg13g2_o21ai_1 _3866_ (.B1(_1286_),
    .Y(_0309_),
    .A1(_0976_),
    .A2(net579));
 sg13g2_nand2_1 _3867_ (.Y(_1287_),
    .A(net297),
    .B(net591));
 sg13g2_o21ai_1 _3868_ (.B1(_1287_),
    .Y(_0310_),
    .A1(_0985_),
    .A2(net579));
 sg13g2_nand2_1 _3869_ (.Y(_1288_),
    .A(net258),
    .B(net590));
 sg13g2_o21ai_1 _3870_ (.B1(_1288_),
    .Y(_0311_),
    .A1(_1006_),
    .A2(net578));
 sg13g2_nand2_1 _3871_ (.Y(_1289_),
    .A(net388),
    .B(net590));
 sg13g2_o21ai_1 _3872_ (.B1(_1289_),
    .Y(_0312_),
    .A1(_1017_),
    .A2(net578));
 sg13g2_nand2_1 _3873_ (.Y(_1290_),
    .A(net381),
    .B(net590));
 sg13g2_o21ai_1 _3874_ (.B1(_1290_),
    .Y(_0313_),
    .A1(_1035_),
    .A2(_1278_));
 sg13g2_nand2_1 _3875_ (.Y(_1291_),
    .A(net294),
    .B(net590));
 sg13g2_o21ai_1 _3876_ (.B1(_1291_),
    .Y(_0314_),
    .A1(_1047_),
    .A2(net579));
 sg13g2_nand2_1 _3877_ (.Y(_1292_),
    .A(net260),
    .B(net590));
 sg13g2_o21ai_1 _3878_ (.B1(_1292_),
    .Y(_0315_),
    .A1(_1059_),
    .A2(net578));
 sg13g2_nand2_1 _3879_ (.Y(_1293_),
    .A(net259),
    .B(net590));
 sg13g2_o21ai_1 _3880_ (.B1(_1293_),
    .Y(_0316_),
    .A1(_1081_),
    .A2(net578));
 sg13g2_or2_1 _3881_ (.X(_1294_),
    .B(net589),
    .A(_0425_));
 sg13g2_inv_1 _3882_ (.Y(_1295_),
    .A(net573));
 sg13g2_nand4_1 _3883_ (.B(\mandelbrot.x[1] ),
    .C(\mandelbrot.x[3] ),
    .A(\mandelbrot.x[0] ),
    .Y(_1296_),
    .D(\mandelbrot.x[2] ));
 sg13g2_nand3b_1 _3884_ (.B(\mandelbrot.x[7] ),
    .C(\mandelbrot.x[8] ),
    .Y(_1297_),
    .A_N(\mandelbrot.x[6] ));
 sg13g2_nor4_2 _3885_ (.A(\mandelbrot.x[5] ),
    .B(\mandelbrot.x[4] ),
    .C(_1296_),
    .Y(_1298_),
    .D(_1297_));
 sg13g2_nor2_1 _3886_ (.A(net678),
    .B(_1298_),
    .Y(_1299_));
 sg13g2_or2_2 _3887_ (.X(_1300_),
    .B(_1298_),
    .A(net678));
 sg13g2_nor2_1 _3888_ (.A(net573),
    .B(net599),
    .Y(_1301_));
 sg13g2_nand2_2 _3889_ (.Y(_1302_),
    .A(_1295_),
    .B(_1300_));
 sg13g2_xor2_1 _3890_ (.B(\configuration[32] ),
    .A(\mandelbrot.alu.in_ci[0] ),
    .X(_1303_));
 sg13g2_nor2_1 _3891_ (.A(net674),
    .B(_1303_),
    .Y(_1304_));
 sg13g2_a21oi_1 _3892_ (.A1(net674),
    .A2(net383),
    .Y(_1305_),
    .B1(_1304_));
 sg13g2_nor2_1 _3893_ (.A(net768),
    .B(net541),
    .Y(_1306_));
 sg13g2_a21oi_1 _3894_ (.A1(net541),
    .A2(_1305_),
    .Y(_0317_),
    .B1(_1306_));
 sg13g2_nor2_1 _3895_ (.A(net510),
    .B(net541),
    .Y(_1307_));
 sg13g2_nand2_1 _3896_ (.Y(_1308_),
    .A(\mandelbrot.alu.in_ci[1] ),
    .B(\configuration[33] ));
 sg13g2_xor2_1 _3897_ (.B(\configuration[33] ),
    .A(\mandelbrot.alu.in_ci[1] ),
    .X(_1309_));
 sg13g2_o21ai_1 _3898_ (.B1(_1309_),
    .Y(_1310_),
    .A1(\mandelbrot.alu.in_ci[0] ),
    .A2(\configuration[32] ));
 sg13g2_nor3_1 _3899_ (.A(\mandelbrot.alu.in_ci[0] ),
    .B(\configuration[32] ),
    .C(_1309_),
    .Y(_1311_));
 sg13g2_nor2_1 _3900_ (.A(net675),
    .B(_1311_),
    .Y(_1312_));
 sg13g2_a22oi_1 _3901_ (.Y(_1313_),
    .B1(_1310_),
    .B2(_1312_),
    .A2(net424),
    .A1(net674));
 sg13g2_a21oi_1 _3902_ (.A1(net541),
    .A2(_1313_),
    .Y(_0318_),
    .B1(_1307_));
 sg13g2_nor2_1 _3903_ (.A(net763),
    .B(net541),
    .Y(_1314_));
 sg13g2_nand2_1 _3904_ (.Y(_1315_),
    .A(\mandelbrot.alu.in_ci[2] ),
    .B(\configuration[34] ));
 sg13g2_xnor2_1 _3905_ (.Y(_1316_),
    .A(\mandelbrot.alu.in_ci[2] ),
    .B(\configuration[34] ));
 sg13g2_nand3_1 _3906_ (.B(_1310_),
    .C(_1316_),
    .A(_1308_),
    .Y(_1317_));
 sg13g2_a21o_1 _3907_ (.A2(_1310_),
    .A1(_1308_),
    .B1(_1316_),
    .X(_1318_));
 sg13g2_a21o_1 _3908_ (.A2(_1318_),
    .A1(_1317_),
    .B1(net675),
    .X(_1319_));
 sg13g2_o21ai_1 _3909_ (.B1(_1319_),
    .Y(_1320_),
    .A1(net661),
    .A2(net398));
 sg13g2_a21oi_1 _3910_ (.A1(net541),
    .A2(_1320_),
    .Y(_0319_),
    .B1(_1314_));
 sg13g2_nand2_1 _3911_ (.Y(_1321_),
    .A(\mandelbrot.alu.in_ci[3] ),
    .B(\configuration[35] ));
 sg13g2_xnor2_1 _3912_ (.Y(_1322_),
    .A(\mandelbrot.alu.in_ci[3] ),
    .B(\configuration[35] ));
 sg13g2_a21o_1 _3913_ (.A2(_1318_),
    .A1(_1315_),
    .B1(_1322_),
    .X(_1323_));
 sg13g2_nand3_1 _3914_ (.B(_1318_),
    .C(_1322_),
    .A(_1315_),
    .Y(_1324_));
 sg13g2_and2_1 _3915_ (.A(net661),
    .B(_1324_),
    .X(_1325_));
 sg13g2_a22oi_1 _3916_ (.Y(_1326_),
    .B1(_1323_),
    .B2(_1325_),
    .A2(net298),
    .A1(net674));
 sg13g2_nor2_1 _3917_ (.A(net456),
    .B(net540),
    .Y(_1327_));
 sg13g2_a21oi_1 _3918_ (.A1(net543),
    .A2(_1326_),
    .Y(_0320_),
    .B1(_1327_));
 sg13g2_xnor2_1 _3919_ (.Y(_1328_),
    .A(\mandelbrot.alu.in_ci[4] ),
    .B(\configuration[36] ));
 sg13g2_a21oi_1 _3920_ (.A1(_1321_),
    .A2(_1323_),
    .Y(_1329_),
    .B1(_1328_));
 sg13g2_and3_1 _3921_ (.X(_1330_),
    .A(_1321_),
    .B(_1323_),
    .C(_1328_));
 sg13g2_nor3_1 _3922_ (.A(net674),
    .B(_1329_),
    .C(_1330_),
    .Y(_1331_));
 sg13g2_a21o_1 _3923_ (.A2(net365),
    .A1(net674),
    .B1(_1331_),
    .X(_1332_));
 sg13g2_mux2_1 _3924_ (.A0(net525),
    .A1(_1332_),
    .S(net540),
    .X(_0321_));
 sg13g2_a21oi_1 _3925_ (.A1(\mandelbrot.alu.in_ci[4] ),
    .A2(\configuration[36] ),
    .Y(_1333_),
    .B1(_1329_));
 sg13g2_nor2_1 _3926_ (.A(\mandelbrot.alu.in_ci[5] ),
    .B(\configuration[37] ),
    .Y(_1334_));
 sg13g2_nand2_1 _3927_ (.Y(_1335_),
    .A(\mandelbrot.alu.in_ci[5] ),
    .B(\configuration[37] ));
 sg13g2_nand2b_1 _3928_ (.Y(_1336_),
    .B(_1335_),
    .A_N(_1334_));
 sg13g2_xnor2_1 _3929_ (.Y(_1337_),
    .A(_1333_),
    .B(_1336_));
 sg13g2_nor2_1 _3930_ (.A(net674),
    .B(_1337_),
    .Y(_1338_));
 sg13g2_a21oi_1 _3931_ (.A1(net674),
    .A2(net389),
    .Y(_1339_),
    .B1(_1338_));
 sg13g2_nor2_1 _3932_ (.A(net519),
    .B(net540),
    .Y(_1340_));
 sg13g2_a21oi_1 _3933_ (.A1(net540),
    .A2(_1339_),
    .Y(_0322_),
    .B1(_1340_));
 sg13g2_nor2_1 _3934_ (.A(net516),
    .B(net540),
    .Y(_1341_));
 sg13g2_and2_1 _3935_ (.A(\mandelbrot.alu.in_ci[6] ),
    .B(\configuration[38] ),
    .X(_1342_));
 sg13g2_or2_1 _3936_ (.X(_1343_),
    .B(\configuration[38] ),
    .A(\mandelbrot.alu.in_ci[6] ));
 sg13g2_nor2b_1 _3937_ (.A(_1342_),
    .B_N(_1343_),
    .Y(_1344_));
 sg13g2_o21ai_1 _3938_ (.B1(_1335_),
    .Y(_1345_),
    .A1(_1333_),
    .A2(_1334_));
 sg13g2_xnor2_1 _3939_ (.Y(_1346_),
    .A(_1344_),
    .B(_1345_));
 sg13g2_nand2_1 _3940_ (.Y(_1347_),
    .A(net660),
    .B(_1346_));
 sg13g2_o21ai_1 _3941_ (.B1(_1347_),
    .Y(_1348_),
    .A1(net660),
    .A2(net384));
 sg13g2_a21oi_1 _3942_ (.A1(net540),
    .A2(_1348_),
    .Y(_0323_),
    .B1(_1341_));
 sg13g2_a21oi_1 _3943_ (.A1(_1343_),
    .A2(_1345_),
    .Y(_1349_),
    .B1(_1342_));
 sg13g2_nor2_1 _3944_ (.A(_0058_),
    .B(_1349_),
    .Y(_1350_));
 sg13g2_and2_1 _3945_ (.A(_0058_),
    .B(_1349_),
    .X(_1351_));
 sg13g2_o21ai_1 _3946_ (.B1(net660),
    .Y(_1352_),
    .A1(_1350_),
    .A2(_1351_));
 sg13g2_o21ai_1 _3947_ (.B1(_1352_),
    .Y(_1353_),
    .A1(net660),
    .A2(net347));
 sg13g2_nor2_1 _3948_ (.A(net372),
    .B(net540),
    .Y(_1354_));
 sg13g2_a21oi_1 _3949_ (.A1(net540),
    .A2(_1353_),
    .Y(_0324_),
    .B1(_1354_));
 sg13g2_nor2_1 _3950_ (.A(net508),
    .B(net539),
    .Y(_1355_));
 sg13g2_nand2_1 _3951_ (.Y(_1356_),
    .A(\mandelbrot.alu.in_ci[8] ),
    .B(_1350_));
 sg13g2_or2_1 _3952_ (.X(_1357_),
    .B(_1350_),
    .A(\mandelbrot.alu.in_ci[8] ));
 sg13g2_a21o_1 _3953_ (.A2(_1357_),
    .A1(_1356_),
    .B1(net676),
    .X(_1358_));
 sg13g2_o21ai_1 _3954_ (.B1(_1358_),
    .Y(_1359_),
    .A1(net660),
    .A2(net375));
 sg13g2_a21oi_1 _3955_ (.A1(net539),
    .A2(_1359_),
    .Y(_0325_),
    .B1(_1355_));
 sg13g2_nor2_1 _3956_ (.A(net377),
    .B(net539),
    .Y(_1360_));
 sg13g2_nor2_2 _3957_ (.A(_1953_),
    .B(_1356_),
    .Y(_1361_));
 sg13g2_a21oi_1 _3958_ (.A1(_1953_),
    .A2(_1356_),
    .Y(_1362_),
    .B1(net676));
 sg13g2_nor2b_1 _3959_ (.A(_1361_),
    .B_N(_1362_),
    .Y(_1363_));
 sg13g2_a21oi_1 _3960_ (.A1(net676),
    .A2(net342),
    .Y(_1364_),
    .B1(_1363_));
 sg13g2_a21oi_1 _3961_ (.A1(net539),
    .A2(_1364_),
    .Y(_0326_),
    .B1(_1360_));
 sg13g2_nor2_1 _3962_ (.A(net518),
    .B(net538),
    .Y(_1365_));
 sg13g2_xnor2_1 _3963_ (.Y(_1366_),
    .A(\mandelbrot.alu.in_ci[10] ),
    .B(_1361_));
 sg13g2_nand2_1 _3964_ (.Y(_1367_),
    .A(net659),
    .B(_1366_));
 sg13g2_o21ai_1 _3965_ (.B1(_1367_),
    .Y(_1368_),
    .A1(net659),
    .A2(net368));
 sg13g2_a21oi_1 _3966_ (.A1(net539),
    .A2(_1368_),
    .Y(_0327_),
    .B1(_1365_));
 sg13g2_nor2_1 _3967_ (.A(net453),
    .B(net537),
    .Y(_1369_));
 sg13g2_and3_2 _3968_ (.X(_1370_),
    .A(\mandelbrot.alu.in_ci[11] ),
    .B(\mandelbrot.alu.in_ci[10] ),
    .C(_1361_));
 sg13g2_a21oi_1 _3969_ (.A1(\mandelbrot.alu.in_ci[10] ),
    .A2(_1361_),
    .Y(_1371_),
    .B1(net453));
 sg13g2_o21ai_1 _3970_ (.B1(net659),
    .Y(_1372_),
    .A1(_1370_),
    .A2(_1371_));
 sg13g2_o21ai_1 _3971_ (.B1(_1372_),
    .Y(_1373_),
    .A1(net659),
    .A2(net395));
 sg13g2_a21oi_1 _3972_ (.A1(net537),
    .A2(_1373_),
    .Y(_0328_),
    .B1(_1369_));
 sg13g2_nor2_1 _3973_ (.A(net712),
    .B(net537),
    .Y(_1374_));
 sg13g2_xnor2_1 _3974_ (.Y(_1375_),
    .A(\mandelbrot.alu.in_ci[12] ),
    .B(_1370_));
 sg13g2_nand2_1 _3975_ (.Y(_1376_),
    .A(net659),
    .B(_1375_));
 sg13g2_o21ai_1 _3976_ (.B1(_1376_),
    .Y(_1377_),
    .A1(net659),
    .A2(net353));
 sg13g2_a21oi_1 _3977_ (.A1(net537),
    .A2(_1377_),
    .Y(_0329_),
    .B1(_1374_));
 sg13g2_nor2_1 _3978_ (.A(net767),
    .B(net538),
    .Y(_1378_));
 sg13g2_nor2_1 _3979_ (.A(net659),
    .B(net355),
    .Y(_1379_));
 sg13g2_nand3_1 _3980_ (.B(\mandelbrot.alu.in_ci[12] ),
    .C(_1370_),
    .A(\mandelbrot.alu.in_ci[13] ),
    .Y(_1380_));
 sg13g2_a21o_1 _3981_ (.A2(_1370_),
    .A1(\mandelbrot.alu.in_ci[12] ),
    .B1(\mandelbrot.alu.in_ci[13] ),
    .X(_1381_));
 sg13g2_a21oi_1 _3982_ (.A1(_1380_),
    .A2(_1381_),
    .Y(_1382_),
    .B1(net676));
 sg13g2_or2_1 _3983_ (.X(_1383_),
    .B(_1382_),
    .A(_1379_));
 sg13g2_a21oi_1 _3984_ (.A1(net538),
    .A2(_1383_),
    .Y(_0330_),
    .B1(_1378_));
 sg13g2_nor2_1 _3985_ (.A(net732),
    .B(net537),
    .Y(_1384_));
 sg13g2_nand2b_1 _3986_ (.Y(_1385_),
    .B(net676),
    .A_N(net340));
 sg13g2_nand4_1 _3987_ (.B(\mandelbrot.alu.in_ci[13] ),
    .C(\mandelbrot.alu.in_ci[12] ),
    .A(net826),
    .Y(_1386_),
    .D(_1370_));
 sg13g2_xnor2_1 _3988_ (.Y(_1387_),
    .A(\mandelbrot.alu.in_ci[14] ),
    .B(_1380_));
 sg13g2_o21ai_1 _3989_ (.B1(_1385_),
    .Y(_1388_),
    .A1(net676),
    .A2(_1387_));
 sg13g2_a21oi_1 _3990_ (.A1(net537),
    .A2(_1388_),
    .Y(_0331_),
    .B1(_1384_));
 sg13g2_a21oi_1 _3991_ (.A1(net673),
    .A2(_1386_),
    .Y(_1389_),
    .B1(net676));
 sg13g2_o21ai_1 _3992_ (.B1(_1389_),
    .Y(_1390_),
    .A1(net673),
    .A2(_1386_));
 sg13g2_o21ai_1 _3993_ (.B1(_1390_),
    .Y(_1391_),
    .A1(net659),
    .A2(net393));
 sg13g2_nor2_1 _3994_ (.A(net673),
    .B(net537),
    .Y(_1392_));
 sg13g2_a21oi_1 _3995_ (.A1(net537),
    .A2(_1391_),
    .Y(_0332_),
    .B1(_1392_));
 sg13g2_nand2_1 _3996_ (.Y(_1393_),
    .A(\mandelbrot.ctr[0] ),
    .B(net588));
 sg13g2_o21ai_1 _3997_ (.B1(_1393_),
    .Y(_0333_),
    .A1(_1909_),
    .A2(net577));
 sg13g2_nand2_1 _3998_ (.Y(_1394_),
    .A(net722),
    .B(net589));
 sg13g2_xnor2_1 _3999_ (.Y(_1395_),
    .A(\mandelbrot.ctr[0] ),
    .B(net722));
 sg13g2_o21ai_1 _4000_ (.B1(_1394_),
    .Y(_0334_),
    .A1(net578),
    .A2(_1395_));
 sg13g2_nand2_1 _4001_ (.Y(_1396_),
    .A(net517),
    .B(net588));
 sg13g2_nand3_1 _4002_ (.B(\mandelbrot.ctr[1] ),
    .C(\mandelbrot.ctr[2] ),
    .A(\mandelbrot.ctr[0] ),
    .Y(_1397_));
 sg13g2_a21o_1 _4003_ (.A2(\mandelbrot.ctr[1] ),
    .A1(\mandelbrot.ctr[0] ),
    .B1(net517),
    .X(_1398_));
 sg13g2_nand2_1 _4004_ (.Y(_1399_),
    .A(_1397_),
    .B(_1398_));
 sg13g2_o21ai_1 _4005_ (.B1(_1396_),
    .Y(_0335_),
    .A1(net577),
    .A2(_1399_));
 sg13g2_nand2_1 _4006_ (.Y(_1400_),
    .A(net509),
    .B(net588));
 sg13g2_nor2_2 _4007_ (.A(_1939_),
    .B(_1397_),
    .Y(_1401_));
 sg13g2_xnor2_1 _4008_ (.Y(_1402_),
    .A(_1939_),
    .B(_1397_));
 sg13g2_o21ai_1 _4009_ (.B1(_1400_),
    .Y(_0336_),
    .A1(net577),
    .A2(_1402_));
 sg13g2_nand2_1 _4010_ (.Y(_1403_),
    .A(net774),
    .B(net588));
 sg13g2_xnor2_1 _4011_ (.Y(_1404_),
    .A(net774),
    .B(_1401_));
 sg13g2_o21ai_1 _4012_ (.B1(_1403_),
    .Y(_0337_),
    .A1(net577),
    .A2(_1404_));
 sg13g2_nand2_1 _4013_ (.Y(_1405_),
    .A(net230),
    .B(net588));
 sg13g2_nand3_1 _4014_ (.B(net672),
    .C(_1401_),
    .A(\mandelbrot.ctr[4] ),
    .Y(_1406_));
 sg13g2_a21o_1 _4015_ (.A2(_1401_),
    .A1(net821),
    .B1(net672),
    .X(_1407_));
 sg13g2_nand2_1 _4016_ (.Y(_1408_),
    .A(_1406_),
    .B(_1407_));
 sg13g2_o21ai_1 _4017_ (.B1(_1405_),
    .Y(_0338_),
    .A1(net577),
    .A2(_1408_));
 sg13g2_nand2_1 _4018_ (.Y(_1409_),
    .A(net505),
    .B(net588));
 sg13g2_or2_1 _4019_ (.X(_1410_),
    .B(_1406_),
    .A(_1941_));
 sg13g2_xnor2_1 _4020_ (.Y(_1411_),
    .A(_1941_),
    .B(_1406_));
 sg13g2_o21ai_1 _4021_ (.B1(_1409_),
    .Y(_0339_),
    .A1(net577),
    .A2(_1411_));
 sg13g2_nand2_1 _4022_ (.Y(_1412_),
    .A(net485),
    .B(net588));
 sg13g2_nor2_1 _4023_ (.A(_1942_),
    .B(_1410_),
    .Y(_1413_));
 sg13g2_xnor2_1 _4024_ (.Y(_1414_),
    .A(_1942_),
    .B(_1410_));
 sg13g2_o21ai_1 _4025_ (.B1(_1412_),
    .Y(_0340_),
    .A1(net577),
    .A2(_1414_));
 sg13g2_nand2_1 _4026_ (.Y(_1415_),
    .A(net735),
    .B(net589));
 sg13g2_nand2_1 _4027_ (.Y(_1416_),
    .A(net824),
    .B(_1413_));
 sg13g2_xnor2_1 _4028_ (.Y(_1417_),
    .A(net735),
    .B(_1413_));
 sg13g2_o21ai_1 _4029_ (.B1(_1415_),
    .Y(_0341_),
    .A1(net578),
    .A2(_1417_));
 sg13g2_nand2_1 _4030_ (.Y(_1418_),
    .A(net715),
    .B(net588));
 sg13g2_xor2_1 _4031_ (.B(_1416_),
    .A(net715),
    .X(_1419_));
 sg13g2_o21ai_1 _4032_ (.B1(_1418_),
    .Y(_0342_),
    .A1(net577),
    .A2(_1419_));
 sg13g2_xor2_1 _4033_ (.B(\configuration[32] ),
    .A(\mandelbrot.alu.in_cr[0] ),
    .X(_1420_));
 sg13g2_nand2_1 _4034_ (.Y(_1421_),
    .A(net596),
    .B(_1420_));
 sg13g2_o21ai_1 _4035_ (.B1(_1421_),
    .Y(_1422_),
    .A1(net376),
    .A2(net596));
 sg13g2_nand2_1 _4036_ (.Y(_1423_),
    .A(net716),
    .B(net568));
 sg13g2_o21ai_1 _4037_ (.B1(_1423_),
    .Y(_0343_),
    .A1(net568),
    .A2(_1422_));
 sg13g2_nand2_1 _4038_ (.Y(_1424_),
    .A(\mandelbrot.alu.in_cr[1] ),
    .B(\configuration[33] ));
 sg13g2_xor2_1 _4039_ (.B(\configuration[33] ),
    .A(\mandelbrot.alu.in_cr[1] ),
    .X(_1425_));
 sg13g2_o21ai_1 _4040_ (.B1(_1425_),
    .Y(_1426_),
    .A1(\mandelbrot.alu.in_cr[0] ),
    .A2(\configuration[32] ));
 sg13g2_or3_1 _4041_ (.A(\mandelbrot.alu.in_cr[0] ),
    .B(\configuration[32] ),
    .C(_1425_),
    .X(_1427_));
 sg13g2_nand3_1 _4042_ (.B(_1426_),
    .C(_1427_),
    .A(net596),
    .Y(_1428_));
 sg13g2_nand2_1 _4043_ (.Y(_1429_),
    .A(\mandelbrot.alu.in_cr[1] ),
    .B(net568));
 sg13g2_o21ai_1 _4044_ (.B1(_1429_),
    .Y(_1430_),
    .A1(net568),
    .A2(_1428_));
 sg13g2_a21o_1 _4045_ (.A2(net541),
    .A1(net308),
    .B1(_1430_),
    .X(_0344_));
 sg13g2_and2_1 _4046_ (.A(\mandelbrot.alu.in_cr[2] ),
    .B(\configuration[34] ),
    .X(_1431_));
 sg13g2_xnor2_1 _4047_ (.Y(_1432_),
    .A(\mandelbrot.alu.in_cr[2] ),
    .B(\configuration[34] ));
 sg13g2_a21oi_1 _4048_ (.A1(_1424_),
    .A2(_1426_),
    .Y(_1433_),
    .B1(_1432_));
 sg13g2_nand3_1 _4049_ (.B(_1426_),
    .C(_1432_),
    .A(_1424_),
    .Y(_1434_));
 sg13g2_nand2_1 _4050_ (.Y(_1435_),
    .A(net596),
    .B(_1434_));
 sg13g2_nand2_1 _4051_ (.Y(_1436_),
    .A(net247),
    .B(_1300_));
 sg13g2_o21ai_1 _4052_ (.B1(_1436_),
    .Y(_1437_),
    .A1(_1433_),
    .A2(_1435_));
 sg13g2_mux2_1 _4053_ (.A0(_1437_),
    .A1(net794),
    .S(net568),
    .X(_0345_));
 sg13g2_nand2_1 _4054_ (.Y(_1438_),
    .A(\mandelbrot.alu.in_cr[3] ),
    .B(\configuration[35] ));
 sg13g2_xor2_1 _4055_ (.B(\configuration[35] ),
    .A(\mandelbrot.alu.in_cr[3] ),
    .X(_1439_));
 sg13g2_o21ai_1 _4056_ (.B1(_1439_),
    .Y(_1440_),
    .A1(_1431_),
    .A2(_1433_));
 sg13g2_or3_1 _4057_ (.A(_1431_),
    .B(_1433_),
    .C(_1439_),
    .X(_1441_));
 sg13g2_nand3_1 _4058_ (.B(_1440_),
    .C(_1441_),
    .A(net596),
    .Y(_1442_));
 sg13g2_o21ai_1 _4059_ (.B1(_1442_),
    .Y(_1443_),
    .A1(_1978_),
    .A2(net596));
 sg13g2_mux2_1 _4060_ (.A0(_1443_),
    .A1(net460),
    .S(net568),
    .X(_0346_));
 sg13g2_xnor2_1 _4061_ (.Y(_1444_),
    .A(\mandelbrot.alu.in_cr[4] ),
    .B(\configuration[36] ));
 sg13g2_a21oi_1 _4062_ (.A1(_1438_),
    .A2(_1440_),
    .Y(_1445_),
    .B1(_1444_));
 sg13g2_and3_1 _4063_ (.X(_1446_),
    .A(_1438_),
    .B(_1440_),
    .C(_1444_));
 sg13g2_nor3_1 _4064_ (.A(_1300_),
    .B(_1445_),
    .C(_1446_),
    .Y(_1447_));
 sg13g2_a21o_1 _4065_ (.A2(_1300_),
    .A1(\configuration[4] ),
    .B1(_1447_),
    .X(_1448_));
 sg13g2_mux2_1 _4066_ (.A0(_1448_),
    .A1(net765),
    .S(net569),
    .X(_0347_));
 sg13g2_a21o_1 _4067_ (.A2(\configuration[36] ),
    .A1(\mandelbrot.alu.in_cr[4] ),
    .B1(_1445_),
    .X(_1449_));
 sg13g2_nor2_1 _4068_ (.A(\mandelbrot.alu.in_cr[5] ),
    .B(\configuration[37] ),
    .Y(_1450_));
 sg13g2_xor2_1 _4069_ (.B(\configuration[37] ),
    .A(\mandelbrot.alu.in_cr[5] ),
    .X(_1451_));
 sg13g2_xnor2_1 _4070_ (.Y(_1452_),
    .A(_1449_),
    .B(_1451_));
 sg13g2_nand2_1 _4071_ (.Y(_1453_),
    .A(net596),
    .B(_1452_));
 sg13g2_o21ai_1 _4072_ (.B1(_1453_),
    .Y(_1454_),
    .A1(net349),
    .A2(net596));
 sg13g2_nand2_1 _4073_ (.Y(_1455_),
    .A(net363),
    .B(net568));
 sg13g2_o21ai_1 _4074_ (.B1(_1455_),
    .Y(_0348_),
    .A1(net568),
    .A2(_1454_));
 sg13g2_and2_1 _4075_ (.A(\mandelbrot.alu.in_cr[6] ),
    .B(\configuration[38] ),
    .X(_1456_));
 sg13g2_xor2_1 _4076_ (.B(\configuration[38] ),
    .A(\mandelbrot.alu.in_cr[6] ),
    .X(_1457_));
 sg13g2_a21oi_1 _4077_ (.A1(\mandelbrot.alu.in_cr[5] ),
    .A2(\configuration[37] ),
    .Y(_1458_),
    .B1(_1449_));
 sg13g2_nor2_1 _4078_ (.A(_1450_),
    .B(_1458_),
    .Y(_1459_));
 sg13g2_xnor2_1 _4079_ (.Y(_1460_),
    .A(_1457_),
    .B(_1459_));
 sg13g2_nand2_1 _4080_ (.Y(_1461_),
    .A(net597),
    .B(_1460_));
 sg13g2_o21ai_1 _4081_ (.B1(_1461_),
    .Y(_1462_),
    .A1(net390),
    .A2(net597));
 sg13g2_nand2_1 _4082_ (.Y(_1463_),
    .A(net482),
    .B(net569));
 sg13g2_o21ai_1 _4083_ (.B1(_1463_),
    .Y(_0349_),
    .A1(net569),
    .A2(_1462_));
 sg13g2_a21oi_1 _4084_ (.A1(_1457_),
    .A2(_1459_),
    .Y(_1464_),
    .B1(_1456_));
 sg13g2_nor2_2 _4085_ (.A(_0053_),
    .B(_1464_),
    .Y(_1465_));
 sg13g2_and2_1 _4086_ (.A(_0053_),
    .B(_1464_),
    .X(_1466_));
 sg13g2_o21ai_1 _4087_ (.B1(net597),
    .Y(_1467_),
    .A1(_1465_),
    .A2(_1466_));
 sg13g2_o21ai_1 _4088_ (.B1(_1467_),
    .Y(_1468_),
    .A1(\configuration[7] ),
    .A2(net597));
 sg13g2_nand2_1 _4089_ (.Y(_1469_),
    .A(net225),
    .B(net570));
 sg13g2_o21ai_1 _4090_ (.B1(_1469_),
    .Y(_0350_),
    .A1(net570),
    .A2(_1468_));
 sg13g2_nand2_1 _4091_ (.Y(_1470_),
    .A(net442),
    .B(net570));
 sg13g2_xor2_1 _4092_ (.B(_1465_),
    .A(_0052_),
    .X(_1471_));
 sg13g2_nand2_1 _4093_ (.Y(_1472_),
    .A(net597),
    .B(_1471_));
 sg13g2_o21ai_1 _4094_ (.B1(_1472_),
    .Y(_1473_),
    .A1(net397),
    .A2(net597));
 sg13g2_o21ai_1 _4095_ (.B1(_1470_),
    .Y(_0351_),
    .A1(net570),
    .A2(_1473_));
 sg13g2_a21oi_1 _4096_ (.A1(net442),
    .A2(_1465_),
    .Y(_1474_),
    .B1(net450));
 sg13g2_nand3_1 _4097_ (.B(\mandelbrot.alu.in_cr[8] ),
    .C(_1465_),
    .A(net450),
    .Y(_1475_));
 sg13g2_nand2_1 _4098_ (.Y(_1476_),
    .A(net598),
    .B(_1475_));
 sg13g2_nand2_1 _4099_ (.Y(_1477_),
    .A(net335),
    .B(_1300_));
 sg13g2_o21ai_1 _4100_ (.B1(_1477_),
    .Y(_1478_),
    .A1(_1474_),
    .A2(_1476_));
 sg13g2_mux2_1 _4101_ (.A0(_1478_),
    .A1(net450),
    .S(net571),
    .X(_0352_));
 sg13g2_nand2b_1 _4102_ (.Y(_1479_),
    .B(_1475_),
    .A_N(net465));
 sg13g2_nand4_1 _4103_ (.B(\mandelbrot.alu.in_cr[9] ),
    .C(\mandelbrot.alu.in_cr[8] ),
    .A(\mandelbrot.alu.in_cr[10] ),
    .Y(_1480_),
    .D(_1465_));
 sg13g2_and2_1 _4104_ (.A(net598),
    .B(_1480_),
    .X(_1481_));
 sg13g2_a22oi_1 _4105_ (.Y(_1482_),
    .B1(_1479_),
    .B2(_1481_),
    .A2(_1300_),
    .A1(net326));
 sg13g2_nand2_1 _4106_ (.Y(_1483_),
    .A(net465),
    .B(net571));
 sg13g2_o21ai_1 _4107_ (.B1(_1483_),
    .Y(_0353_),
    .A1(net571),
    .A2(_1482_));
 sg13g2_nand2_1 _4108_ (.Y(_1484_),
    .A(_1949_),
    .B(_1480_));
 sg13g2_nor2_2 _4109_ (.A(_1949_),
    .B(_1480_),
    .Y(_1485_));
 sg13g2_nor2_1 _4110_ (.A(_1300_),
    .B(_1485_),
    .Y(_1486_));
 sg13g2_a221oi_1 _4111_ (.B2(_1486_),
    .C1(net571),
    .B1(_1484_),
    .A1(net310),
    .Y(_1487_),
    .A2(_1300_));
 sg13g2_a21oi_1 _4112_ (.A1(_1949_),
    .A2(net571),
    .Y(_0354_),
    .B1(_1487_));
 sg13g2_xnor2_1 _4113_ (.Y(_1488_),
    .A(\mandelbrot.alu.in_cr[12] ),
    .B(_1485_));
 sg13g2_nand2_1 _4114_ (.Y(_1489_),
    .A(net598),
    .B(_1488_));
 sg13g2_o21ai_1 _4115_ (.B1(_1489_),
    .Y(_1490_),
    .A1(net231),
    .A2(net598));
 sg13g2_nand2_1 _4116_ (.Y(_1491_),
    .A(net726),
    .B(net572));
 sg13g2_o21ai_1 _4117_ (.B1(_1491_),
    .Y(_0355_),
    .A1(net572),
    .A2(_1490_));
 sg13g2_nand3_1 _4118_ (.B(\mandelbrot.alu.in_cr[12] ),
    .C(_1485_),
    .A(\mandelbrot.alu.in_cr[13] ),
    .Y(_1492_));
 sg13g2_a21o_1 _4119_ (.A2(_1485_),
    .A1(\mandelbrot.alu.in_cr[12] ),
    .B1(\mandelbrot.alu.in_cr[13] ),
    .X(_1493_));
 sg13g2_nand3_1 _4120_ (.B(_1492_),
    .C(_1493_),
    .A(net598),
    .Y(_1494_));
 sg13g2_o21ai_1 _4121_ (.B1(_1494_),
    .Y(_1495_),
    .A1(_1979_),
    .A2(net598));
 sg13g2_mux2_1 _4122_ (.A0(_1495_),
    .A1(net520),
    .S(net572),
    .X(_0356_));
 sg13g2_xor2_1 _4123_ (.B(_1492_),
    .A(\mandelbrot.alu.in_cr[14] ),
    .X(_1496_));
 sg13g2_nand2_1 _4124_ (.Y(_1497_),
    .A(net598),
    .B(_1496_));
 sg13g2_o21ai_1 _4125_ (.B1(_1497_),
    .Y(_1498_),
    .A1(net324),
    .A2(net598));
 sg13g2_nand2_1 _4126_ (.Y(_1499_),
    .A(net394),
    .B(net571));
 sg13g2_o21ai_1 _4127_ (.B1(_1499_),
    .Y(_0357_),
    .A1(net572),
    .A2(_1498_));
 sg13g2_nor2_1 _4128_ (.A(_0050_),
    .B(_1492_),
    .Y(_1500_));
 sg13g2_xnor2_1 _4129_ (.Y(_1501_),
    .A(\mandelbrot.alu.in_cr[15] ),
    .B(_1500_));
 sg13g2_nand2_1 _4130_ (.Y(_1502_),
    .A(net599),
    .B(_1501_));
 sg13g2_o21ai_1 _4131_ (.B1(_1502_),
    .Y(_1503_),
    .A1(net344),
    .A2(net599));
 sg13g2_nand2_1 _4132_ (.Y(_1504_),
    .A(net720),
    .B(net571));
 sg13g2_o21ai_1 _4133_ (.B1(_1504_),
    .Y(_0358_),
    .A1(net571),
    .A2(_1503_));
 sg13g2_nand3b_1 _4134_ (.B(\mandelbrot.y[1] ),
    .C(\mandelbrot.y[0] ),
    .Y(_1505_),
    .A_N(net410));
 sg13g2_nand4_1 _4135_ (.B(_1945_),
    .C(\mandelbrot.y[5] ),
    .A(\mandelbrot.y[3] ),
    .Y(_1506_),
    .D(\mandelbrot.y[8] ));
 sg13g2_nor4_2 _4136_ (.A(\mandelbrot.y[7] ),
    .B(\mandelbrot.y[6] ),
    .C(_1505_),
    .Y(_1507_),
    .D(_1506_));
 sg13g2_nand3_1 _4137_ (.B(_1298_),
    .C(_1507_),
    .A(_2157_),
    .Y(_1508_));
 sg13g2_a22oi_1 _4138_ (.Y(_1509_),
    .B1(_1508_),
    .B2(net223),
    .A2(\mandelbrot.run ),
    .A1(net677));
 sg13g2_inv_1 _4139_ (.Y(_0359_),
    .A(net224));
 sg13g2_nand2_2 _4140_ (.Y(_1510_),
    .A(_2157_),
    .B(net626));
 sg13g2_nor2_1 _4141_ (.A(\configuration[40] ),
    .B(\configuration[39] ),
    .Y(_1511_));
 sg13g2_o21ai_1 _4142_ (.B1(_0018_),
    .Y(_1512_),
    .A1(\configuration[41] ),
    .A2(_1511_));
 sg13g2_inv_1 _4143_ (.Y(_1513_),
    .A(_1512_));
 sg13g2_nand2_1 _4144_ (.Y(_1514_),
    .A(\configuration[40] ),
    .B(\configuration[39] ));
 sg13g2_nor2_1 _4145_ (.A(_0018_),
    .B(_1514_),
    .Y(_1515_));
 sg13g2_o21ai_1 _4146_ (.B1(\mandelbrot.ctr[0] ),
    .Y(_1516_),
    .A1(_1513_),
    .A2(_1515_));
 sg13g2_nand2b_1 _4147_ (.Y(_1517_),
    .B(\configuration[39] ),
    .A_N(\configuration[40] ));
 sg13g2_nor2_1 _4148_ (.A(\configuration[41] ),
    .B(_1517_),
    .Y(_1518_));
 sg13g2_nand2b_1 _4149_ (.Y(_1519_),
    .B(\configuration[40] ),
    .A_N(\configuration[39] ));
 sg13g2_nor2_1 _4150_ (.A(\configuration[41] ),
    .B(_1519_),
    .Y(_1520_));
 sg13g2_nor2_1 _4151_ (.A(_0018_),
    .B(_1519_),
    .Y(_1521_));
 sg13g2_nor2_2 _4152_ (.A(_0018_),
    .B(_1517_),
    .Y(_1522_));
 sg13g2_nor3_2 _4153_ (.A(\configuration[40] ),
    .B(\configuration[39] ),
    .C(_0018_),
    .Y(_1523_));
 sg13g2_nor2_1 _4154_ (.A(\configuration[41] ),
    .B(_1514_),
    .Y(_1524_));
 sg13g2_a22oi_1 _4155_ (.Y(_1525_),
    .B1(_1523_),
    .B2(\mandelbrot.ctr[4] ),
    .A2(_1520_),
    .A1(\mandelbrot.ctr[2] ));
 sg13g2_a22oi_1 _4156_ (.Y(_1526_),
    .B1(_1524_),
    .B2(\mandelbrot.ctr[3] ),
    .A2(_1522_),
    .A1(net672));
 sg13g2_a22oi_1 _4157_ (.Y(_1527_),
    .B1(_1521_),
    .B2(\mandelbrot.ctr[6] ),
    .A2(_1518_),
    .A1(\mandelbrot.ctr[1] ));
 sg13g2_nand4_1 _4158_ (.B(_1525_),
    .C(_1526_),
    .A(_1516_),
    .Y(_1528_),
    .D(_1527_));
 sg13g2_mux2_1 _4159_ (.A0(_1528_),
    .A1(net781),
    .S(_1510_),
    .X(_0360_));
 sg13g2_nand2_1 _4160_ (.Y(_1529_),
    .A(net486),
    .B(_1510_));
 sg13g2_a22oi_1 _4161_ (.Y(_1530_),
    .B1(_1524_),
    .B2(\mandelbrot.ctr[4] ),
    .A2(_1522_),
    .A1(\mandelbrot.ctr[6] ));
 sg13g2_a22oi_1 _4162_ (.Y(_1531_),
    .B1(_1521_),
    .B2(\mandelbrot.ctr[7] ),
    .A2(_1518_),
    .A1(\mandelbrot.ctr[2] ));
 sg13g2_and2_1 _4163_ (.A(_1530_),
    .B(_1531_),
    .X(_1532_));
 sg13g2_o21ai_1 _4164_ (.B1(\mandelbrot.ctr[3] ),
    .Y(_1533_),
    .A1(_1515_),
    .A2(_1520_));
 sg13g2_a21oi_1 _4165_ (.A1(net672),
    .A2(_1511_),
    .Y(_1534_),
    .B1(_1513_));
 sg13g2_nand3_1 _4166_ (.B(_1533_),
    .C(_1534_),
    .A(_1532_),
    .Y(_1535_));
 sg13g2_o21ai_1 _4167_ (.B1(_1535_),
    .Y(_1536_),
    .A1(net820),
    .A2(_1512_));
 sg13g2_o21ai_1 _4168_ (.B1(_1529_),
    .Y(_0361_),
    .A1(_1510_),
    .A2(_1536_));
 sg13g2_nor3_1 _4169_ (.A(_1940_),
    .B(\configuration[41] ),
    .C(_1519_),
    .Y(_1537_));
 sg13g2_o21ai_1 _4170_ (.B1(\mandelbrot.ctr[6] ),
    .Y(_1538_),
    .A1(_1515_),
    .A2(_1523_));
 sg13g2_a22oi_1 _4171_ (.Y(_1539_),
    .B1(_1522_),
    .B2(\mandelbrot.ctr[7] ),
    .A2(_1521_),
    .A1(\mandelbrot.ctr[8] ));
 sg13g2_a221oi_1 _4172_ (.B2(net672),
    .C1(_1537_),
    .B1(_1524_),
    .A1(\mandelbrot.ctr[3] ),
    .Y(_1540_),
    .A2(_1518_));
 sg13g2_nand4_1 _4173_ (.B(_1538_),
    .C(_1539_),
    .A(_1512_),
    .Y(_1541_),
    .D(_1540_));
 sg13g2_o21ai_1 _4174_ (.B1(_1541_),
    .Y(_1542_),
    .A1(\mandelbrot.ctr[2] ),
    .A2(_1512_));
 sg13g2_nand2_1 _4175_ (.Y(_1543_),
    .A(net503),
    .B(_1510_));
 sg13g2_o21ai_1 _4176_ (.B1(_1543_),
    .Y(_0362_),
    .A1(_1510_),
    .A2(_1542_));
 sg13g2_nor3_1 _4177_ (.A(_1941_),
    .B(\configuration[41] ),
    .C(_1514_),
    .Y(_1544_));
 sg13g2_nand2_1 _4178_ (.Y(_1545_),
    .A(\mandelbrot.ctr[9] ),
    .B(\configuration[40] ));
 sg13g2_o21ai_1 _4179_ (.B1(_1512_),
    .Y(_1546_),
    .A1(_0018_),
    .A2(_1545_));
 sg13g2_a221oi_1 _4180_ (.B2(\mandelbrot.ctr[7] ),
    .C1(_1544_),
    .B1(_1523_),
    .A1(\mandelbrot.ctr[8] ),
    .Y(_1547_),
    .A2(_1522_));
 sg13g2_a221oi_1 _4181_ (.B2(net672),
    .C1(_1546_),
    .B1(_1520_),
    .A1(\mandelbrot.ctr[4] ),
    .Y(_1548_),
    .A2(_1518_));
 sg13g2_a22oi_1 _4182_ (.Y(_1549_),
    .B1(_1547_),
    .B2(_1548_),
    .A2(_1513_),
    .A1(_1939_));
 sg13g2_mux2_1 _4183_ (.A0(_1549_),
    .A1(net793),
    .S(_1510_),
    .X(_0363_));
 sg13g2_nand2_1 _4184_ (.Y(_1550_),
    .A(net252),
    .B(net590));
 sg13g2_nand2_1 _4185_ (.Y(_1551_),
    .A(\mandelbrot.alu.in_ci[15] ),
    .B(\mandelbrot.alu.m3[29] ));
 sg13g2_nor2_1 _4186_ (.A(net673),
    .B(\mandelbrot.alu.m3[29] ),
    .Y(_1552_));
 sg13g2_xor2_1 _4187_ (.B(\mandelbrot.alu.m3[29] ),
    .A(net673),
    .X(_1553_));
 sg13g2_o21ai_1 _4188_ (.B1(_0616_),
    .Y(_1554_),
    .A1(_0601_),
    .A2(_0619_));
 sg13g2_a21oi_2 _4189_ (.B1(_1554_),
    .Y(_1555_),
    .A2(_0617_),
    .A1(_0598_));
 sg13g2_nand2_1 _4190_ (.Y(_1556_),
    .A(net673),
    .B(\mandelbrot.alu.m3[30] ));
 sg13g2_xor2_1 _4191_ (.B(\mandelbrot.alu.m3[30] ),
    .A(net673),
    .X(_1557_));
 sg13g2_nand3b_1 _4192_ (.B(_1557_),
    .C(_1553_),
    .Y(_1558_),
    .A_N(_1555_));
 sg13g2_nand3_1 _4193_ (.B(_1556_),
    .C(_1558_),
    .A(_1551_),
    .Y(_1559_));
 sg13g2_xor2_1 _4194_ (.B(\mandelbrot.alu.m3[31] ),
    .A(net673),
    .X(_1560_));
 sg13g2_xnor2_1 _4195_ (.Y(_1561_),
    .A(_1559_),
    .B(_1560_));
 sg13g2_o21ai_1 _4196_ (.B1(_1551_),
    .Y(_1562_),
    .A1(_1552_),
    .A2(_1555_));
 sg13g2_xnor2_1 _4197_ (.Y(_1563_),
    .A(_1557_),
    .B(_1562_));
 sg13g2_xor2_1 _4198_ (.B(_1555_),
    .A(_1553_),
    .X(_1564_));
 sg13g2_nand3_1 _4199_ (.B(_1563_),
    .C(_1564_),
    .A(_0620_),
    .Y(_1565_));
 sg13g2_nor3_2 _4200_ (.A(_0620_),
    .B(_1563_),
    .C(_1564_),
    .Y(_1566_));
 sg13g2_nor2_2 _4201_ (.A(_1561_),
    .B(_1566_),
    .Y(_1567_));
 sg13g2_nand2b_1 _4202_ (.Y(_1568_),
    .B(\mandelbrot.alu.m2[29] ),
    .A_N(\mandelbrot.alu.m1[29] ));
 sg13g2_nor2b_1 _4203_ (.A(\mandelbrot.alu.m2[29] ),
    .B_N(\mandelbrot.alu.m1[29] ),
    .Y(_1569_));
 sg13g2_a21o_1 _4204_ (.A2(_1568_),
    .A1(_1073_),
    .B1(_1569_),
    .X(_1570_));
 sg13g2_xnor2_1 _4205_ (.Y(_1571_),
    .A(_1980_),
    .B(_1570_));
 sg13g2_xnor2_1 _4206_ (.Y(_1572_),
    .A(\mandelbrot.alu.in_cr[15] ),
    .B(_1571_));
 sg13g2_nand2_1 _4207_ (.Y(_1573_),
    .A(_1077_),
    .B(_1079_));
 sg13g2_a221oi_1 _4208_ (.B2(_1573_),
    .C1(_1050_),
    .B1(_1076_),
    .A1(_1033_),
    .Y(_1574_),
    .A2(_1045_));
 sg13g2_nand3_1 _4209_ (.B(_1077_),
    .C(_1079_),
    .A(_1058_),
    .Y(_1575_));
 sg13g2_nand2_1 _4210_ (.Y(_1576_),
    .A(_1076_),
    .B(_1575_));
 sg13g2_or2_1 _4211_ (.X(_1577_),
    .B(_1576_),
    .A(_1574_));
 sg13g2_nor3_1 _4212_ (.A(_1572_),
    .B(_1574_),
    .C(_1576_),
    .Y(_1578_));
 sg13g2_nor2b_1 _4213_ (.A(\mandelbrot.alu.m2[30] ),
    .B_N(\mandelbrot.alu.m1[30] ),
    .Y(_1579_));
 sg13g2_a21oi_1 _4214_ (.A1(_1981_),
    .A2(_1570_),
    .Y(_1580_),
    .B1(_1579_));
 sg13g2_xnor2_1 _4215_ (.Y(_1581_),
    .A(_2126_),
    .B(_1580_));
 sg13g2_xor2_1 _4216_ (.B(_1581_),
    .A(\mandelbrot.alu.in_cr[15] ),
    .X(_1582_));
 sg13g2_a21oi_1 _4217_ (.A1(\mandelbrot.alu.in_cr[15] ),
    .A2(_1571_),
    .Y(_1583_),
    .B1(_1581_));
 sg13g2_nor2_1 _4218_ (.A(_0049_),
    .B(_1583_),
    .Y(_1584_));
 sg13g2_a21oi_1 _4219_ (.A1(_1578_),
    .A2(_1582_),
    .Y(_1585_),
    .B1(_1584_));
 sg13g2_nor2b_1 _4220_ (.A(\mandelbrot.alu.m2[31] ),
    .B_N(\mandelbrot.alu.m1[31] ),
    .Y(_1586_));
 sg13g2_a21oi_1 _4221_ (.A1(_2126_),
    .A2(_1580_),
    .Y(_1587_),
    .B1(_1586_));
 sg13g2_xnor2_1 _4222_ (.Y(_1588_),
    .A(\mandelbrot.alu.in_cr[15] ),
    .B(_1587_));
 sg13g2_xor2_1 _4223_ (.B(_1588_),
    .A(_1585_),
    .X(_1589_));
 sg13g2_nand2b_1 _4224_ (.Y(_1590_),
    .B(_1571_),
    .A_N(_0049_));
 sg13g2_nand2b_1 _4225_ (.Y(_1591_),
    .B(_1590_),
    .A_N(_1578_));
 sg13g2_xnor2_1 _4226_ (.Y(_1592_),
    .A(_1582_),
    .B(_1591_));
 sg13g2_xnor2_1 _4227_ (.Y(_1593_),
    .A(_1572_),
    .B(_1577_));
 sg13g2_nand4_1 _4228_ (.B(_1589_),
    .C(_1592_),
    .A(_1081_),
    .Y(_1594_),
    .D(_1593_));
 sg13g2_or4_1 _4229_ (.A(_1081_),
    .B(_1589_),
    .C(_1592_),
    .D(_1593_),
    .X(_1595_));
 sg13g2_a221oi_1 _4230_ (.B2(_1595_),
    .C1(_1567_),
    .B1(_1594_),
    .A1(_1561_),
    .Y(_1596_),
    .A2(_1565_));
 sg13g2_o21ai_1 _4231_ (.B1(_1550_),
    .Y(_0364_),
    .A1(net578),
    .A2(_1596_));
 sg13g2_a21oi_1 _4232_ (.A1(net212),
    .A2(net599),
    .Y(_1597_),
    .B1(net573));
 sg13g2_a21oi_1 _4233_ (.A1(_1946_),
    .A2(net573),
    .Y(_0365_),
    .B1(_1597_));
 sg13g2_and3_1 _4234_ (.X(_1598_),
    .A(\mandelbrot.x[0] ),
    .B(net249),
    .C(_1295_));
 sg13g2_a21oi_1 _4235_ (.A1(\mandelbrot.x[0] ),
    .A2(_1295_),
    .Y(_1599_),
    .B1(net249));
 sg13g2_nor3_1 _4236_ (.A(net542),
    .B(_1598_),
    .C(net250),
    .Y(_0366_));
 sg13g2_xnor2_1 _4237_ (.Y(_1600_),
    .A(net432),
    .B(_1598_));
 sg13g2_a21oi_1 _4238_ (.A1(net678),
    .A2(_1295_),
    .Y(_0367_),
    .B1(net433));
 sg13g2_a21oi_1 _4239_ (.A1(\mandelbrot.x[2] ),
    .A2(_1598_),
    .Y(_1601_),
    .B1(net264));
 sg13g2_nor2_1 _4240_ (.A(net573),
    .B(_1296_),
    .Y(_1602_));
 sg13g2_a21oi_1 _4241_ (.A1(net662),
    .A2(_1296_),
    .Y(_1603_),
    .B1(net573));
 sg13g2_nor2_1 _4242_ (.A(net265),
    .B(_1603_),
    .Y(_0368_));
 sg13g2_nor2_1 _4243_ (.A(net458),
    .B(_1602_),
    .Y(_1604_));
 sg13g2_nor3_2 _4244_ (.A(_1947_),
    .B(net573),
    .C(_1296_),
    .Y(_1605_));
 sg13g2_nor3_1 _4245_ (.A(net542),
    .B(net459),
    .C(_1605_),
    .Y(_0369_));
 sg13g2_o21ai_1 _4246_ (.B1(net536),
    .Y(_1606_),
    .A1(net454),
    .A2(_1605_));
 sg13g2_a21oi_1 _4247_ (.A1(net454),
    .A2(_1605_),
    .Y(_0370_),
    .B1(_1606_));
 sg13g2_a21oi_1 _4248_ (.A1(\mandelbrot.x[5] ),
    .A2(_1605_),
    .Y(_1607_),
    .B1(net305));
 sg13g2_and3_1 _4249_ (.X(_1608_),
    .A(net454),
    .B(net305),
    .C(_1605_));
 sg13g2_nor3_1 _4250_ (.A(net542),
    .B(net306),
    .C(_1608_),
    .Y(_0371_));
 sg13g2_and4_1 _4251_ (.A(net454),
    .B(net305),
    .C(net477),
    .D(_1605_),
    .X(_1609_));
 sg13g2_o21ai_1 _4252_ (.B1(net536),
    .Y(_1610_),
    .A1(net477),
    .A2(_1608_));
 sg13g2_nor2_1 _4253_ (.A(_1609_),
    .B(_1610_),
    .Y(_0372_));
 sg13g2_xnor2_1 _4254_ (.Y(_1611_),
    .A(net391),
    .B(_1609_));
 sg13g2_nor2_1 _4255_ (.A(net542),
    .B(net392),
    .Y(_0373_));
 sg13g2_nand2_1 _4256_ (.Y(_1612_),
    .A(net671),
    .B(net587));
 sg13g2_o21ai_1 _4257_ (.B1(_1612_),
    .Y(_0374_),
    .A1(_0510_),
    .A2(net576));
 sg13g2_nand2_1 _4258_ (.Y(_1613_),
    .A(net422),
    .B(net587));
 sg13g2_o21ai_1 _4259_ (.B1(_1613_),
    .Y(_0375_),
    .A1(_0515_),
    .A2(net576));
 sg13g2_nand2_1 _4260_ (.Y(_1614_),
    .A(net323),
    .B(net587));
 sg13g2_o21ai_1 _4261_ (.B1(_1614_),
    .Y(_0376_),
    .A1(_0520_),
    .A2(net576));
 sg13g2_nand2_1 _4262_ (.Y(_1615_),
    .A(net276),
    .B(net587));
 sg13g2_o21ai_1 _4263_ (.B1(_1615_),
    .Y(_0377_),
    .A1(_0525_),
    .A2(net576));
 sg13g2_nand2_1 _4264_ (.Y(_1616_),
    .A(net469),
    .B(net585));
 sg13g2_o21ai_1 _4265_ (.B1(_1616_),
    .Y(_0378_),
    .A1(_0531_),
    .A2(net574));
 sg13g2_nand2_1 _4266_ (.Y(_1617_),
    .A(net358),
    .B(net585));
 sg13g2_o21ai_1 _4267_ (.B1(_1617_),
    .Y(_0379_),
    .A1(_0537_),
    .A2(net574));
 sg13g2_nand2_1 _4268_ (.Y(_1618_),
    .A(net332),
    .B(net585));
 sg13g2_o21ai_1 _4269_ (.B1(_1618_),
    .Y(_0380_),
    .A1(_0545_),
    .A2(net574));
 sg13g2_nand2_1 _4270_ (.Y(_1619_),
    .A(net263),
    .B(net585));
 sg13g2_o21ai_1 _4271_ (.B1(_1619_),
    .Y(_0381_),
    .A1(_0552_),
    .A2(net574));
 sg13g2_nand2_1 _4272_ (.Y(_1620_),
    .A(net487),
    .B(net586));
 sg13g2_o21ai_1 _4273_ (.B1(_1620_),
    .Y(_0382_),
    .A1(_0558_),
    .A2(net575));
 sg13g2_nand2_1 _4274_ (.Y(_1621_),
    .A(net337),
    .B(net585));
 sg13g2_o21ai_1 _4275_ (.B1(_1621_),
    .Y(_0383_),
    .A1(_0565_),
    .A2(net575));
 sg13g2_nand2_1 _4276_ (.Y(_1622_),
    .A(net295),
    .B(net586));
 sg13g2_o21ai_1 _4277_ (.B1(_1622_),
    .Y(_0384_),
    .A1(_0574_),
    .A2(net575));
 sg13g2_nand2_1 _4278_ (.Y(_1623_),
    .A(net431),
    .B(net586));
 sg13g2_o21ai_1 _4279_ (.B1(_1623_),
    .Y(_0385_),
    .A1(_0581_),
    .A2(net574));
 sg13g2_nand2_1 _4280_ (.Y(_1624_),
    .A(net304),
    .B(net586));
 sg13g2_o21ai_1 _4281_ (.B1(_1624_),
    .Y(_0386_),
    .A1(_0589_),
    .A2(net575));
 sg13g2_nand2_1 _4282_ (.Y(_1625_),
    .A(net328),
    .B(net585));
 sg13g2_o21ai_1 _4283_ (.B1(_1625_),
    .Y(_0387_),
    .A1(_0595_),
    .A2(net574));
 sg13g2_nand2_1 _4284_ (.Y(_1626_),
    .A(net314),
    .B(net585));
 sg13g2_o21ai_1 _4285_ (.B1(_1626_),
    .Y(_0388_),
    .A1(_0603_),
    .A2(net574));
 sg13g2_nand2_1 _4286_ (.Y(_1627_),
    .A(net289),
    .B(net585));
 sg13g2_o21ai_1 _4287_ (.B1(_1627_),
    .Y(_0389_),
    .A1(_0620_),
    .A2(net574));
 sg13g2_nand2_1 _4288_ (.Y(_1628_),
    .A(\mandelbrot.y[0] ),
    .B(_1302_));
 sg13g2_nand3_1 _4289_ (.B(_1274_),
    .C(_1298_),
    .A(_2157_),
    .Y(_1629_));
 sg13g2_o21ai_1 _4290_ (.B1(_1628_),
    .Y(_0117_),
    .A1(_1908_),
    .A2(_1629_));
 sg13g2_a21oi_1 _4291_ (.A1(\mandelbrot.y[0] ),
    .A2(net428),
    .Y(_1630_),
    .B1(net677));
 sg13g2_nor2_1 _4292_ (.A(net536),
    .B(_1630_),
    .Y(_1631_));
 sg13g2_a21oi_1 _4293_ (.A1(\mandelbrot.y[0] ),
    .A2(net541),
    .Y(_1632_),
    .B1(net428));
 sg13g2_nor2_1 _4294_ (.A(_1631_),
    .B(net429),
    .Y(_0118_));
 sg13g2_o21ai_1 _4295_ (.B1(net410),
    .Y(_1633_),
    .A1(_1302_),
    .A2(_1630_));
 sg13g2_o21ai_1 _4296_ (.B1(_1633_),
    .Y(_0119_),
    .A1(_1505_),
    .A2(_1629_));
 sg13g2_nand2_1 _4297_ (.Y(_1634_),
    .A(net439),
    .B(_1302_));
 sg13g2_nand3_1 _4298_ (.B(net428),
    .C(net410),
    .A(\mandelbrot.y[0] ),
    .Y(_1635_));
 sg13g2_nand4_1 _4299_ (.B(\mandelbrot.y[1] ),
    .C(\mandelbrot.y[3] ),
    .A(\mandelbrot.y[0] ),
    .Y(_1636_),
    .D(\mandelbrot.y[2] ));
 sg13g2_xor2_1 _4300_ (.B(_1635_),
    .A(net439),
    .X(_1637_));
 sg13g2_o21ai_1 _4301_ (.B1(_1634_),
    .Y(_0120_),
    .A1(_1629_),
    .A2(_1637_));
 sg13g2_nand2_1 _4302_ (.Y(_1638_),
    .A(net256),
    .B(net536));
 sg13g2_nor2_2 _4303_ (.A(_1945_),
    .B(_1636_),
    .Y(_1639_));
 sg13g2_xnor2_1 _4304_ (.Y(_1640_),
    .A(_1945_),
    .B(_1636_));
 sg13g2_o21ai_1 _4305_ (.B1(_1638_),
    .Y(_0121_),
    .A1(_1629_),
    .A2(_1640_));
 sg13g2_nand2_1 _4306_ (.Y(_1641_),
    .A(net483),
    .B(net536));
 sg13g2_xnor2_1 _4307_ (.Y(_1642_),
    .A(net483),
    .B(_1639_));
 sg13g2_o21ai_1 _4308_ (.B1(_1641_),
    .Y(_0122_),
    .A1(_1629_),
    .A2(_1642_));
 sg13g2_nand2_1 _4309_ (.Y(_1643_),
    .A(net418),
    .B(net536));
 sg13g2_nand3_1 _4310_ (.B(net418),
    .C(_1639_),
    .A(\mandelbrot.y[5] ),
    .Y(_1644_));
 sg13g2_a21o_1 _4311_ (.A2(_1639_),
    .A1(\mandelbrot.y[5] ),
    .B1(net418),
    .X(_1645_));
 sg13g2_nand2_1 _4312_ (.Y(_1646_),
    .A(_1644_),
    .B(_1645_));
 sg13g2_o21ai_1 _4313_ (.B1(_1643_),
    .Y(_0123_),
    .A1(_1629_),
    .A2(_1646_));
 sg13g2_nand2_1 _4314_ (.Y(_1647_),
    .A(net488),
    .B(net536));
 sg13g2_nand4_1 _4315_ (.B(\mandelbrot.y[7] ),
    .C(\mandelbrot.y[6] ),
    .A(\mandelbrot.y[5] ),
    .Y(_1648_),
    .D(_1639_));
 sg13g2_xor2_1 _4316_ (.B(_1644_),
    .A(net488),
    .X(_1649_));
 sg13g2_o21ai_1 _4317_ (.B1(_1647_),
    .Y(_0124_),
    .A1(_1629_),
    .A2(_1649_));
 sg13g2_nand2_1 _4318_ (.Y(_1650_),
    .A(net284),
    .B(net536));
 sg13g2_xor2_1 _4319_ (.B(_1648_),
    .A(net284),
    .X(_1651_));
 sg13g2_o21ai_1 _4320_ (.B1(_1650_),
    .Y(_0125_),
    .A1(_1629_),
    .A2(_1651_));
 sg13g2_o21ai_1 _4321_ (.B1(_1261_),
    .Y(_1652_),
    .A1(_1257_),
    .A2(_1262_));
 sg13g2_xor2_1 _4322_ (.B(_1258_),
    .A(_0030_),
    .X(_1653_));
 sg13g2_xnor2_1 _4323_ (.Y(_1654_),
    .A(_1652_),
    .B(_1653_));
 sg13g2_nor2_1 _4324_ (.A(_1132_),
    .B(_1654_),
    .Y(_1655_));
 sg13g2_nand2_1 _4325_ (.Y(_1656_),
    .A(net421),
    .B(net564));
 sg13g2_a21oi_1 _4326_ (.A1(_1132_),
    .A2(_1656_),
    .Y(_0126_),
    .B1(_1655_));
 sg13g2_a22oi_1 _4327_ (.Y(_1657_),
    .B1(net526),
    .B2(net546),
    .A2(net665),
    .A1(net689));
 sg13g2_inv_1 _4328_ (.Y(_0127_),
    .A(_1657_));
 sg13g2_a22oi_1 _4329_ (.Y(_1658_),
    .B1(_0877_),
    .B2(net567),
    .A2(net546),
    .A1(\mandelbrot.alu.m1[0] ));
 sg13g2_o21ai_1 _4330_ (.B1(_1658_),
    .Y(_0128_),
    .A1(net657),
    .A2(_1933_));
 sg13g2_a22oi_1 _4331_ (.Y(_1659_),
    .B1(net667),
    .B2(net545),
    .A2(net809),
    .A1(net689));
 sg13g2_o21ai_1 _4332_ (.B1(net810),
    .Y(_0129_),
    .A1(net566),
    .A2(_0885_));
 sg13g2_a22oi_1 _4333_ (.Y(_1660_),
    .B1(_0900_),
    .B2(net567),
    .A2(net544),
    .A1(net499));
 sg13g2_o21ai_1 _4334_ (.B1(_1660_),
    .Y(_0130_),
    .A1(net657),
    .A2(_1932_));
 sg13g2_a22oi_1 _4335_ (.Y(_1661_),
    .B1(_0911_),
    .B2(_0427_),
    .A2(net545),
    .A1(\mandelbrot.alu.m1[3] ));
 sg13g2_o21ai_1 _4336_ (.B1(_1661_),
    .Y(_0131_),
    .A1(net658),
    .A2(_1931_));
 sg13g2_nor2_1 _4337_ (.A(net566),
    .B(_0925_),
    .Y(_1662_));
 sg13g2_a221oi_1 _4338_ (.B2(net544),
    .C1(_1662_),
    .B1(net738),
    .A1(net689),
    .Y(_1663_),
    .A2(net534));
 sg13g2_inv_1 _4339_ (.Y(_0132_),
    .A(_1663_));
 sg13g2_a22oi_1 _4340_ (.Y(_1664_),
    .B1(net513),
    .B2(net545),
    .A2(net791),
    .A1(net689));
 sg13g2_o21ai_1 _4341_ (.B1(_1664_),
    .Y(_0133_),
    .A1(net566),
    .A2(_0935_));
 sg13g2_a22oi_1 _4342_ (.Y(_1665_),
    .B1(net534),
    .B2(net544),
    .A2(\mandelbrot.alu.m1[8] ),
    .A1(net689));
 sg13g2_o21ai_1 _4343_ (.B1(net535),
    .Y(_0134_),
    .A1(net566),
    .A2(_0951_));
 sg13g2_nor2_1 _4344_ (.A(net566),
    .B(_0961_),
    .Y(_1666_));
 sg13g2_a221oi_1 _4345_ (.B2(net544),
    .C1(_1666_),
    .B1(net791),
    .A1(net689),
    .Y(_1667_),
    .A2(net814));
 sg13g2_inv_1 _4346_ (.Y(_0135_),
    .A(_1667_));
 sg13g2_a22oi_1 _4347_ (.Y(_1668_),
    .B1(_0977_),
    .B2(net567),
    .A2(net544),
    .A1(net759));
 sg13g2_o21ai_1 _4348_ (.B1(_1668_),
    .Y(_0136_),
    .A1(net657),
    .A2(_1930_));
 sg13g2_a22oi_1 _4349_ (.Y(_1669_),
    .B1(_0986_),
    .B2(net567),
    .A2(net544),
    .A1(\mandelbrot.alu.m1[9] ));
 sg13g2_o21ai_1 _4350_ (.B1(_1669_),
    .Y(_0137_),
    .A1(net657),
    .A2(_1929_));
 sg13g2_a22oi_1 _4351_ (.Y(_1670_),
    .B1(net750),
    .B2(net544),
    .A2(\mandelbrot.alu.m1[12] ),
    .A1(net689));
 sg13g2_o21ai_1 _4352_ (.B1(net751),
    .Y(_0138_),
    .A1(net566),
    .A2(_1007_));
 sg13g2_a22oi_1 _4353_ (.Y(_1671_),
    .B1(_1018_),
    .B2(net567),
    .A2(net544),
    .A1(net470));
 sg13g2_o21ai_1 _4354_ (.B1(_1671_),
    .Y(_0139_),
    .A1(net657),
    .A2(_1927_));
 sg13g2_a22oi_1 _4355_ (.Y(_1672_),
    .B1(_1036_),
    .B2(net567),
    .A2(net545),
    .A1(\mandelbrot.alu.m1[12] ));
 sg13g2_o21ai_1 _4356_ (.B1(_1672_),
    .Y(_0140_),
    .A1(net657),
    .A2(_1925_));
 sg13g2_a22oi_1 _4357_ (.Y(_1673_),
    .B1(_1048_),
    .B2(net567),
    .A2(net545),
    .A1(net533));
 sg13g2_o21ai_1 _4358_ (.B1(_1673_),
    .Y(_0141_),
    .A1(net657),
    .A2(_1924_));
 sg13g2_nor2_1 _4359_ (.A(net566),
    .B(_1060_),
    .Y(_1674_));
 sg13g2_nand2_1 _4360_ (.Y(_1675_),
    .A(\mandelbrot.alu.m1[0] ),
    .B(\mandelbrot.alu.mult_zr_zr.shift_reg[0] ));
 sg13g2_a21o_2 _4361_ (.A2(\mandelbrot.alu.mult_zr_zr.shift_reg[0] ),
    .A1(\mandelbrot.alu.m1[0] ),
    .B1(net665),
    .X(_1676_));
 sg13g2_nor2_1 _4362_ (.A(\mandelbrot.alu.m1[0] ),
    .B(\mandelbrot.alu.mult_zr_zr.shift_reg[0] ),
    .Y(_1677_));
 sg13g2_o21ai_1 _4363_ (.B1(net665),
    .Y(_1678_),
    .A1(\mandelbrot.alu.m1[0] ),
    .A2(\mandelbrot.alu.mult_zr_zr.shift_reg[0] ));
 sg13g2_and2_1 _4364_ (.A(_1676_),
    .B(_1678_),
    .X(_1679_));
 sg13g2_nand2_2 _4365_ (.Y(_1680_),
    .A(_1676_),
    .B(_1678_));
 sg13g2_nor2_1 _4366_ (.A(net666),
    .B(_1677_),
    .Y(_1681_));
 sg13g2_a21oi_2 _4367_ (.B1(_1681_),
    .Y(_1682_),
    .A2(_1675_),
    .A1(net666));
 sg13g2_a21o_1 _4368_ (.A2(_1675_),
    .A1(net666),
    .B1(_1681_),
    .X(_1683_));
 sg13g2_nand3_1 _4369_ (.B(net634),
    .C(net592),
    .A(\mandelbrot.alu.in_zr[0] ),
    .Y(_1684_));
 sg13g2_xor2_1 _4370_ (.B(_1684_),
    .A(net764),
    .X(_1685_));
 sg13g2_a221oi_1 _4371_ (.B2(net689),
    .C1(_1674_),
    .B1(_1685_),
    .A1(_1925_),
    .Y(_0142_),
    .A2(net545));
 sg13g2_and3_1 _4372_ (.X(_1686_),
    .A(\mandelbrot.alu.m1[16] ),
    .B(\mandelbrot.alu.in_zr[0] ),
    .C(net634));
 sg13g2_nor2_1 _4373_ (.A(net666),
    .B(_0073_),
    .Y(_1687_));
 sg13g2_nor2_1 _4374_ (.A(\mandelbrot.alu.in_zr[0] ),
    .B(\mandelbrot.alu.in_zr[1] ),
    .Y(_1688_));
 sg13g2_xor2_1 _4375_ (.B(\mandelbrot.alu.in_zr[1] ),
    .A(\mandelbrot.alu.in_zr[0] ),
    .X(_1689_));
 sg13g2_xnor2_1 _4376_ (.Y(_1690_),
    .A(\mandelbrot.alu.in_zr[0] ),
    .B(\mandelbrot.alu.in_zr[1] ));
 sg13g2_a221oi_1 _4377_ (.B2(net666),
    .C1(_1687_),
    .B1(_1689_),
    .A1(_1676_),
    .Y(_1691_),
    .A2(_1678_));
 sg13g2_and3_1 _4378_ (.X(_1692_),
    .A(_0074_),
    .B(_1676_),
    .C(_1678_));
 sg13g2_nor3_1 _4379_ (.A(_1921_),
    .B(_1691_),
    .C(_1692_),
    .Y(_1693_));
 sg13g2_o21ai_1 _4380_ (.B1(_1921_),
    .Y(_1694_),
    .A1(_1691_),
    .A2(_1692_));
 sg13g2_nor2b_1 _4381_ (.A(_1693_),
    .B_N(_1694_),
    .Y(_1695_));
 sg13g2_xnor2_1 _4382_ (.Y(_1696_),
    .A(_1686_),
    .B(_1695_));
 sg13g2_o21ai_1 _4383_ (.B1(net690),
    .Y(_1697_),
    .A1(\mandelbrot.alu.m1[17] ),
    .A2(net592));
 sg13g2_a21oi_1 _4384_ (.A1(net592),
    .A2(_1696_),
    .Y(_1698_),
    .B1(_1697_));
 sg13g2_a221oi_1 _4385_ (.B2(net567),
    .C1(_1698_),
    .B1(_1082_),
    .A1(net724),
    .Y(_1699_),
    .A2(net545));
 sg13g2_inv_1 _4386_ (.Y(_0143_),
    .A(_1699_));
 sg13g2_a21o_1 _4387_ (.A2(_1694_),
    .A1(_1686_),
    .B1(_1693_),
    .X(_1700_));
 sg13g2_nor3_1 _4388_ (.A(\mandelbrot.alu.in_zr[0] ),
    .B(\mandelbrot.alu.in_zr[1] ),
    .C(\mandelbrot.alu.in_zr[2] ),
    .Y(_1701_));
 sg13g2_xor2_1 _4389_ (.B(_1688_),
    .A(\mandelbrot.alu.in_zr[2] ),
    .X(_1702_));
 sg13g2_mux2_1 _4390_ (.A0(_0072_),
    .A1(_1702_),
    .S(net667),
    .X(_1703_));
 sg13g2_mux4_1 _4391_ (.S0(net634),
    .A0(_0073_),
    .A1(_0072_),
    .A2(_1690_),
    .A3(_1702_),
    .S1(net665),
    .X(_1704_));
 sg13g2_xnor2_1 _4392_ (.Y(_1705_),
    .A(\mandelbrot.alu.m1[18] ),
    .B(_1704_));
 sg13g2_nand2_2 _4393_ (.Y(_1706_),
    .A(net691),
    .B(net593));
 sg13g2_xor2_1 _4394_ (.B(_1705_),
    .A(_1700_),
    .X(_1707_));
 sg13g2_nor2_1 _4395_ (.A(net594),
    .B(_1707_),
    .Y(_1708_));
 sg13g2_a21oi_1 _4396_ (.A1(net451),
    .A2(net594),
    .Y(_1709_),
    .B1(_1708_));
 sg13g2_a22oi_1 _4397_ (.Y(_1710_),
    .B1(_1709_),
    .B2(net690),
    .A2(net549),
    .A1(\mandelbrot.alu.m1[16] ));
 sg13g2_inv_1 _4398_ (.Y(_0144_),
    .A(net452));
 sg13g2_or2_1 _4399_ (.X(_1711_),
    .B(_0071_),
    .A(net667));
 sg13g2_or4_2 _4400_ (.A(\mandelbrot.alu.in_zr[0] ),
    .B(\mandelbrot.alu.in_zr[1] ),
    .C(\mandelbrot.alu.in_zr[2] ),
    .D(\mandelbrot.alu.in_zr[3] ),
    .X(_1712_));
 sg13g2_xor2_1 _4401_ (.B(_1701_),
    .A(\mandelbrot.alu.in_zr[3] ),
    .X(_1713_));
 sg13g2_o21ai_1 _4402_ (.B1(_1711_),
    .Y(_1714_),
    .A1(_1935_),
    .A2(_1713_));
 sg13g2_nand2_1 _4403_ (.Y(_1715_),
    .A(net635),
    .B(_1703_));
 sg13g2_nand2b_1 _4404_ (.Y(_1716_),
    .B(net634),
    .A_N(_1714_));
 sg13g2_nand3_1 _4405_ (.B(_1715_),
    .C(_1716_),
    .A(\mandelbrot.alu.m1[19] ),
    .Y(_1717_));
 sg13g2_a21oi_1 _4406_ (.A1(_1715_),
    .A2(_1716_),
    .Y(_1718_),
    .B1(\mandelbrot.alu.m1[19] ));
 sg13g2_a21o_1 _4407_ (.A2(_1716_),
    .A1(_1715_),
    .B1(\mandelbrot.alu.m1[19] ),
    .X(_1719_));
 sg13g2_nand2_1 _4408_ (.Y(_1720_),
    .A(_1717_),
    .B(_1719_));
 sg13g2_nor2_1 _4409_ (.A(_0029_),
    .B(_1704_),
    .Y(_1721_));
 sg13g2_a21oi_1 _4410_ (.A1(_1700_),
    .A2(_1705_),
    .Y(_1722_),
    .B1(_1721_));
 sg13g2_xnor2_1 _4411_ (.Y(_1723_),
    .A(_1720_),
    .B(_1722_));
 sg13g2_nand2_1 _4412_ (.Y(_1724_),
    .A(net592),
    .B(_1723_));
 sg13g2_a21oi_1 _4413_ (.A1(net273),
    .A2(net594),
    .Y(_1725_),
    .B1(net658));
 sg13g2_a22oi_1 _4414_ (.Y(_1726_),
    .B1(_1724_),
    .B2(_1725_),
    .A2(net549),
    .A1(\mandelbrot.alu.m1[17] ));
 sg13g2_inv_1 _4415_ (.Y(_0145_),
    .A(net274));
 sg13g2_o21ai_1 _4416_ (.B1(_1717_),
    .Y(_1727_),
    .A1(_1718_),
    .A2(_1722_));
 sg13g2_nor2_1 _4417_ (.A(net667),
    .B(_0070_),
    .Y(_1728_));
 sg13g2_xor2_1 _4418_ (.B(_1712_),
    .A(\mandelbrot.alu.in_zr[4] ),
    .X(_1729_));
 sg13g2_a21oi_1 _4419_ (.A1(net667),
    .A2(_1729_),
    .Y(_1730_),
    .B1(_1728_));
 sg13g2_nand2_1 _4420_ (.Y(_1731_),
    .A(net635),
    .B(_1714_));
 sg13g2_o21ai_1 _4421_ (.B1(_1731_),
    .Y(_1732_),
    .A1(net635),
    .A2(_1730_));
 sg13g2_xor2_1 _4422_ (.B(_1732_),
    .A(\mandelbrot.alu.m1[20] ),
    .X(_1733_));
 sg13g2_xor2_1 _4423_ (.B(_1733_),
    .A(_1727_),
    .X(_1734_));
 sg13g2_nor2_1 _4424_ (.A(net594),
    .B(_1734_),
    .Y(_1735_));
 sg13g2_a21oi_1 _4425_ (.A1(net478),
    .A2(net594),
    .Y(_1736_),
    .B1(_1735_));
 sg13g2_a22oi_1 _4426_ (.Y(_1737_),
    .B1(_1736_),
    .B2(net690),
    .A2(net546),
    .A1(\mandelbrot.alu.m1[18] ));
 sg13g2_inv_1 _4427_ (.Y(_0146_),
    .A(net479));
 sg13g2_a22oi_1 _4428_ (.Y(_1738_),
    .B1(_1733_),
    .B2(_1727_),
    .A2(_1732_),
    .A1(_1964_));
 sg13g2_o21ai_1 _4429_ (.B1(\mandelbrot.alu.in_zr[5] ),
    .Y(_1739_),
    .A1(\mandelbrot.alu.in_zr[4] ),
    .A2(_1712_));
 sg13g2_nor3_2 _4430_ (.A(\mandelbrot.alu.in_zr[4] ),
    .B(\mandelbrot.alu.in_zr[5] ),
    .C(_1712_),
    .Y(_1740_));
 sg13g2_nor2_1 _4431_ (.A(_1935_),
    .B(_1740_),
    .Y(_1741_));
 sg13g2_a22oi_1 _4432_ (.Y(_1742_),
    .B1(_1739_),
    .B2(_1741_),
    .A2(_1965_),
    .A1(_1935_));
 sg13g2_nand2_1 _4433_ (.Y(_1743_),
    .A(net635),
    .B(_1730_));
 sg13g2_nand2_1 _4434_ (.Y(_1744_),
    .A(net634),
    .B(_1742_));
 sg13g2_and3_1 _4435_ (.X(_1745_),
    .A(\mandelbrot.alu.m1[21] ),
    .B(_1743_),
    .C(_1744_));
 sg13g2_a21oi_2 _4436_ (.B1(\mandelbrot.alu.m1[21] ),
    .Y(_1746_),
    .A2(_1744_),
    .A1(_1743_));
 sg13g2_nor2_1 _4437_ (.A(_1745_),
    .B(_1746_),
    .Y(_1747_));
 sg13g2_o21ai_1 _4438_ (.B1(net592),
    .Y(_1748_),
    .A1(_1738_),
    .A2(_1747_));
 sg13g2_a21oi_1 _4439_ (.A1(_1738_),
    .A2(_1747_),
    .Y(_1749_),
    .B1(_1748_));
 sg13g2_a21oi_1 _4440_ (.A1(net472),
    .A2(net594),
    .Y(_1750_),
    .B1(_1749_));
 sg13g2_a22oi_1 _4441_ (.Y(_1751_),
    .B1(_1750_),
    .B2(net690),
    .A2(net546),
    .A1(\mandelbrot.alu.m1[19] ));
 sg13g2_inv_1 _4442_ (.Y(_0147_),
    .A(net473));
 sg13g2_a221oi_1 _4443_ (.B2(_1727_),
    .C1(_1745_),
    .B1(_1733_),
    .A1(_1964_),
    .Y(_1752_),
    .A2(_1732_));
 sg13g2_nor2_1 _4444_ (.A(net668),
    .B(_0068_),
    .Y(_1753_));
 sg13g2_nor2b_1 _4445_ (.A(\mandelbrot.alu.in_zr[6] ),
    .B_N(_1740_),
    .Y(_1754_));
 sg13g2_xnor2_1 _4446_ (.Y(_1755_),
    .A(\mandelbrot.alu.in_zr[6] ),
    .B(_1740_));
 sg13g2_a21oi_1 _4447_ (.A1(net668),
    .A2(_1755_),
    .Y(_1756_),
    .B1(_1753_));
 sg13g2_mux2_1 _4448_ (.A0(_1742_),
    .A1(_1756_),
    .S(net634),
    .X(_1757_));
 sg13g2_xor2_1 _4449_ (.B(_1757_),
    .A(\mandelbrot.alu.m1[22] ),
    .X(_1758_));
 sg13g2_nor3_1 _4450_ (.A(_1746_),
    .B(_1752_),
    .C(_1758_),
    .Y(_1759_));
 sg13g2_or3_1 _4451_ (.A(_1746_),
    .B(_1752_),
    .C(_1758_),
    .X(_1760_));
 sg13g2_o21ai_1 _4452_ (.B1(_1758_),
    .Y(_1761_),
    .A1(_1746_),
    .A2(_1752_));
 sg13g2_a21oi_1 _4453_ (.A1(_1760_),
    .A2(_1761_),
    .Y(_1762_),
    .B1(net594));
 sg13g2_a21oi_1 _4454_ (.A1(net467),
    .A2(net594),
    .Y(_1763_),
    .B1(_1762_));
 sg13g2_a22oi_1 _4455_ (.Y(_1764_),
    .B1(_1763_),
    .B2(net693),
    .A2(net546),
    .A1(\mandelbrot.alu.m1[20] ));
 sg13g2_inv_1 _4456_ (.Y(_0148_),
    .A(net468));
 sg13g2_nand2_1 _4457_ (.Y(_1765_),
    .A(net461),
    .B(net546));
 sg13g2_nor2_1 _4458_ (.A(net668),
    .B(_0067_),
    .Y(_1766_));
 sg13g2_nand2b_2 _4459_ (.Y(_1767_),
    .B(_1754_),
    .A_N(\mandelbrot.alu.in_zr[7] ));
 sg13g2_xnor2_1 _4460_ (.Y(_1768_),
    .A(\mandelbrot.alu.in_zr[7] ),
    .B(_1754_));
 sg13g2_a21oi_1 _4461_ (.A1(net668),
    .A2(_1768_),
    .Y(_1769_),
    .B1(_1766_));
 sg13g2_mux2_1 _4462_ (.A0(_1756_),
    .A1(_1769_),
    .S(net634),
    .X(_1770_));
 sg13g2_nand2b_1 _4463_ (.Y(_1771_),
    .B(\mandelbrot.alu.m1[23] ),
    .A_N(_1770_));
 sg13g2_xnor2_1 _4464_ (.Y(_1772_),
    .A(\mandelbrot.alu.m1[23] ),
    .B(_1770_));
 sg13g2_nor2_1 _4465_ (.A(_0025_),
    .B(_1757_),
    .Y(_1773_));
 sg13g2_nor3_1 _4466_ (.A(_1759_),
    .B(_1772_),
    .C(_1773_),
    .Y(_1774_));
 sg13g2_o21ai_1 _4467_ (.B1(_1772_),
    .Y(_1775_),
    .A1(_1759_),
    .A2(_1773_));
 sg13g2_nand2b_1 _4468_ (.Y(_1776_),
    .B(_1775_),
    .A_N(_1774_));
 sg13g2_a21oi_1 _4469_ (.A1(net593),
    .A2(_1776_),
    .Y(_1777_),
    .B1(net203));
 sg13g2_o21ai_1 _4470_ (.B1(_1777_),
    .Y(_1778_),
    .A1(\mandelbrot.alu.m1[23] ),
    .A2(net592));
 sg13g2_o21ai_1 _4471_ (.B1(_1765_),
    .Y(_0149_),
    .A1(net546),
    .A2(_1778_));
 sg13g2_a21oi_1 _4472_ (.A1(\mandelbrot.alu.in_zr[8] ),
    .A2(_1767_),
    .Y(_1779_),
    .B1(_1935_));
 sg13g2_o21ai_1 _4473_ (.B1(_1779_),
    .Y(_1780_),
    .A1(\mandelbrot.alu.in_zr[8] ),
    .A2(_1767_));
 sg13g2_o21ai_1 _4474_ (.B1(_1780_),
    .Y(_1781_),
    .A1(net668),
    .A2(_0066_));
 sg13g2_nor2_1 _4475_ (.A(net634),
    .B(_1769_),
    .Y(_1782_));
 sg13g2_a21oi_2 _4476_ (.B1(_1782_),
    .Y(_1783_),
    .A2(_1781_),
    .A1(net633));
 sg13g2_xor2_1 _4477_ (.B(_1783_),
    .A(\mandelbrot.alu.m1[24] ),
    .X(_1784_));
 sg13g2_a21oi_1 _4478_ (.A1(_1771_),
    .A2(_1775_),
    .Y(_1785_),
    .B1(_1784_));
 sg13g2_nand3_1 _4479_ (.B(_1775_),
    .C(_1784_),
    .A(_1771_),
    .Y(_1786_));
 sg13g2_nor2b_1 _4480_ (.A(_1785_),
    .B_N(_1786_),
    .Y(_1787_));
 sg13g2_nor2_1 _4481_ (.A(net595),
    .B(_1787_),
    .Y(_1788_));
 sg13g2_a21oi_1 _4482_ (.A1(net317),
    .A2(net595),
    .Y(_1789_),
    .B1(_1788_));
 sg13g2_a22oi_1 _4483_ (.Y(_1790_),
    .B1(_1789_),
    .B2(net692),
    .A2(net547),
    .A1(\mandelbrot.alu.m1[22] ));
 sg13g2_inv_1 _4484_ (.Y(_0150_),
    .A(net318));
 sg13g2_nor2_1 _4485_ (.A(_0024_),
    .B(_1783_),
    .Y(_1791_));
 sg13g2_nor2_1 _4486_ (.A(_1785_),
    .B(_1791_),
    .Y(_1792_));
 sg13g2_nor2_1 _4487_ (.A(net668),
    .B(_0065_),
    .Y(_1793_));
 sg13g2_nor3_2 _4488_ (.A(\mandelbrot.alu.in_zr[8] ),
    .B(\mandelbrot.alu.in_zr[9] ),
    .C(_1767_),
    .Y(_1794_));
 sg13g2_o21ai_1 _4489_ (.B1(\mandelbrot.alu.in_zr[9] ),
    .Y(_1795_),
    .A1(\mandelbrot.alu.in_zr[8] ),
    .A2(_1767_));
 sg13g2_nor2b_1 _4490_ (.A(_1794_),
    .B_N(_1795_),
    .Y(_1796_));
 sg13g2_a21oi_1 _4491_ (.A1(net670),
    .A2(_1796_),
    .Y(_1797_),
    .B1(_1793_));
 sg13g2_nor2_1 _4492_ (.A(_1679_),
    .B(_1797_),
    .Y(_1798_));
 sg13g2_a21oi_1 _4493_ (.A1(net635),
    .A2(_1781_),
    .Y(_1799_),
    .B1(_1798_));
 sg13g2_nor2b_1 _4494_ (.A(\mandelbrot.alu.m1[25] ),
    .B_N(_1799_),
    .Y(_1800_));
 sg13g2_nor2b_1 _4495_ (.A(_1799_),
    .B_N(\mandelbrot.alu.m1[25] ),
    .Y(_1801_));
 sg13g2_inv_1 _4496_ (.Y(_1802_),
    .A(_1801_));
 sg13g2_nor2_1 _4497_ (.A(_1800_),
    .B(_1801_),
    .Y(_1803_));
 sg13g2_xor2_1 _4498_ (.B(_1803_),
    .A(_1792_),
    .X(_1804_));
 sg13g2_nand2b_1 _4499_ (.Y(_1805_),
    .B(net692),
    .A_N(net755));
 sg13g2_a22oi_1 _4500_ (.Y(_1806_),
    .B1(_1805_),
    .B2(_1706_),
    .A2(_1804_),
    .A1(net593));
 sg13g2_a21o_1 _4501_ (.A2(net547),
    .A1(\mandelbrot.alu.m1[23] ),
    .B1(_1806_),
    .X(_0151_));
 sg13g2_a21oi_2 _4502_ (.B1(_1800_),
    .Y(_1807_),
    .A2(_1802_),
    .A1(_1792_));
 sg13g2_nand2b_2 _4503_ (.Y(_1808_),
    .B(_1794_),
    .A_N(\mandelbrot.alu.in_zr[10] ));
 sg13g2_nand2b_1 _4504_ (.Y(_1809_),
    .B(\mandelbrot.alu.in_zr[10] ),
    .A_N(_1794_));
 sg13g2_nand3_1 _4505_ (.B(_1808_),
    .C(_1809_),
    .A(net668),
    .Y(_1810_));
 sg13g2_o21ai_1 _4506_ (.B1(_1810_),
    .Y(_1811_),
    .A1(net668),
    .A2(_0064_));
 sg13g2_nor2_1 _4507_ (.A(net633),
    .B(_1797_),
    .Y(_1812_));
 sg13g2_a21oi_1 _4508_ (.A1(net633),
    .A2(_1811_),
    .Y(_1813_),
    .B1(_1812_));
 sg13g2_xnor2_1 _4509_ (.Y(_1814_),
    .A(\mandelbrot.alu.m1[26] ),
    .B(_1813_));
 sg13g2_xor2_1 _4510_ (.B(_1814_),
    .A(_1807_),
    .X(_1815_));
 sg13g2_o21ai_1 _4511_ (.B1(net692),
    .Y(_1816_),
    .A1(net595),
    .A2(_1815_));
 sg13g2_a21oi_1 _4512_ (.A1(net366),
    .A2(net595),
    .Y(_1817_),
    .B1(_1816_));
 sg13g2_a21o_1 _4513_ (.A2(net547),
    .A1(\mandelbrot.alu.m1[24] ),
    .B1(_1817_),
    .X(_0152_));
 sg13g2_a21oi_1 _4514_ (.A1(\mandelbrot.alu.in_zr[11] ),
    .A2(_1808_),
    .Y(_1818_),
    .B1(_1935_));
 sg13g2_o21ai_1 _4515_ (.B1(_1818_),
    .Y(_1819_),
    .A1(\mandelbrot.alu.in_zr[11] ),
    .A2(_1808_));
 sg13g2_o21ai_1 _4516_ (.B1(_1819_),
    .Y(_1820_),
    .A1(net669),
    .A2(_0063_));
 sg13g2_mux2_1 _4517_ (.A0(_1811_),
    .A1(_1820_),
    .S(net633),
    .X(_1821_));
 sg13g2_nand2_1 _4518_ (.Y(_1822_),
    .A(\mandelbrot.alu.m1[27] ),
    .B(_1821_));
 sg13g2_nor2_1 _4519_ (.A(\mandelbrot.alu.m1[27] ),
    .B(_1821_),
    .Y(_1823_));
 sg13g2_xnor2_1 _4520_ (.Y(_1824_),
    .A(_1920_),
    .B(_1821_));
 sg13g2_nor2_1 _4521_ (.A(_0022_),
    .B(_1813_),
    .Y(_1825_));
 sg13g2_a21oi_2 _4522_ (.B1(_1825_),
    .Y(_1826_),
    .A2(_1814_),
    .A1(_1807_));
 sg13g2_a21oi_1 _4523_ (.A1(_1824_),
    .A2(_1826_),
    .Y(_1827_),
    .B1(net595));
 sg13g2_o21ai_1 _4524_ (.B1(_1827_),
    .Y(_1828_),
    .A1(_1824_),
    .A2(_1826_));
 sg13g2_o21ai_1 _4525_ (.B1(_1828_),
    .Y(_1829_),
    .A1(\mandelbrot.alu.m1[27] ),
    .A2(net593));
 sg13g2_nor3_1 _4526_ (.A(net203),
    .B(net548),
    .C(_1829_),
    .Y(_1830_));
 sg13g2_a21o_1 _4527_ (.A2(net548),
    .A1(net476),
    .B1(_1830_),
    .X(_0153_));
 sg13g2_a21oi_2 _4528_ (.B1(_1823_),
    .Y(_1831_),
    .A2(_1826_),
    .A1(_1822_));
 sg13g2_nor2_1 _4529_ (.A(net669),
    .B(_0062_),
    .Y(_1832_));
 sg13g2_nor3_1 _4530_ (.A(\mandelbrot.alu.in_zr[11] ),
    .B(\mandelbrot.alu.in_zr[12] ),
    .C(_1808_),
    .Y(_1833_));
 sg13g2_o21ai_1 _4531_ (.B1(\mandelbrot.alu.in_zr[12] ),
    .Y(_1834_),
    .A1(\mandelbrot.alu.in_zr[11] ),
    .A2(_1808_));
 sg13g2_nand3b_1 _4532_ (.B(_1834_),
    .C(net669),
    .Y(_1835_),
    .A_N(_1833_));
 sg13g2_nor2b_1 _4533_ (.A(_1832_),
    .B_N(_1835_),
    .Y(_1836_));
 sg13g2_nor2_1 _4534_ (.A(net635),
    .B(_1836_),
    .Y(_1837_));
 sg13g2_a21oi_1 _4535_ (.A1(net635),
    .A2(_1820_),
    .Y(_1838_),
    .B1(_1837_));
 sg13g2_xnor2_1 _4536_ (.Y(_1839_),
    .A(\mandelbrot.alu.m1[28] ),
    .B(_1838_));
 sg13g2_xor2_1 _4537_ (.B(_1839_),
    .A(_1831_),
    .X(_1840_));
 sg13g2_nor2_1 _4538_ (.A(net595),
    .B(_1840_),
    .Y(_1841_));
 sg13g2_a21oi_1 _4539_ (.A1(net359),
    .A2(net595),
    .Y(_1842_),
    .B1(_1841_));
 sg13g2_a22oi_1 _4540_ (.Y(_1843_),
    .B1(_1842_),
    .B2(net692),
    .A2(net547),
    .A1(\mandelbrot.alu.m1[26] ));
 sg13g2_inv_1 _4541_ (.Y(_0154_),
    .A(net360));
 sg13g2_nor2_1 _4542_ (.A(net669),
    .B(_0061_),
    .Y(_1844_));
 sg13g2_nor2b_1 _4543_ (.A(\mandelbrot.alu.in_zr[13] ),
    .B_N(_1833_),
    .Y(_1845_));
 sg13g2_xnor2_1 _4544_ (.Y(_1846_),
    .A(\mandelbrot.alu.in_zr[13] ),
    .B(_1833_));
 sg13g2_a21oi_1 _4545_ (.A1(net670),
    .A2(_1846_),
    .Y(_1847_),
    .B1(_1844_));
 sg13g2_nand2_1 _4546_ (.Y(_1848_),
    .A(net635),
    .B(_1836_));
 sg13g2_nand2_1 _4547_ (.Y(_1849_),
    .A(net633),
    .B(_1847_));
 sg13g2_and3_1 _4548_ (.X(_1850_),
    .A(\mandelbrot.alu.m1[29] ),
    .B(_1848_),
    .C(_1849_));
 sg13g2_a21oi_1 _4549_ (.A1(_1848_),
    .A2(_1849_),
    .Y(_1851_),
    .B1(\mandelbrot.alu.m1[29] ));
 sg13g2_nor2_1 _4550_ (.A(_1850_),
    .B(_1851_),
    .Y(_1852_));
 sg13g2_nor2_1 _4551_ (.A(_0021_),
    .B(_1838_),
    .Y(_1853_));
 sg13g2_a21oi_1 _4552_ (.A1(_1831_),
    .A2(_1839_),
    .Y(_1854_),
    .B1(_1853_));
 sg13g2_xor2_1 _4553_ (.B(_1854_),
    .A(_1852_),
    .X(_1855_));
 sg13g2_nand2b_1 _4554_ (.Y(_1856_),
    .B(net691),
    .A_N(net769));
 sg13g2_a22oi_1 _4555_ (.Y(_1857_),
    .B1(_1856_),
    .B2(_1706_),
    .A2(_1855_),
    .A1(net593));
 sg13g2_a21o_1 _4556_ (.A2(net547),
    .A1(\mandelbrot.alu.m1[27] ),
    .B1(_1857_),
    .X(_0155_));
 sg13g2_and2_1 _4557_ (.A(_1839_),
    .B(_1852_),
    .X(_1858_));
 sg13g2_a21o_1 _4558_ (.A2(_1853_),
    .A1(_1852_),
    .B1(_1850_),
    .X(_1859_));
 sg13g2_a21o_1 _4559_ (.A2(_1858_),
    .A1(_1831_),
    .B1(_1859_),
    .X(_1860_));
 sg13g2_nand2b_1 _4560_ (.Y(_1861_),
    .B(\mandelbrot.alu.in_zr[14] ),
    .A_N(_1845_));
 sg13g2_nand2b_1 _4561_ (.Y(_1862_),
    .B(_1845_),
    .A_N(\mandelbrot.alu.in_zr[14] ));
 sg13g2_nand3_1 _4562_ (.B(_1861_),
    .C(_1862_),
    .A(net669),
    .Y(_1863_));
 sg13g2_o21ai_1 _4563_ (.B1(_1863_),
    .Y(_1864_),
    .A1(net669),
    .A2(_0060_));
 sg13g2_nor2_1 _4564_ (.A(net633),
    .B(_1847_),
    .Y(_1865_));
 sg13g2_a21oi_1 _4565_ (.A1(net633),
    .A2(_1864_),
    .Y(_1866_),
    .B1(_1865_));
 sg13g2_xnor2_1 _4566_ (.Y(_1867_),
    .A(\mandelbrot.alu.m1[30] ),
    .B(_1866_));
 sg13g2_xnor2_1 _4567_ (.Y(_1868_),
    .A(_1860_),
    .B(_1867_));
 sg13g2_a21o_1 _4568_ (.A2(net595),
    .A1(_0019_),
    .B1(net658),
    .X(_1869_));
 sg13g2_a21oi_1 _4569_ (.A1(net593),
    .A2(_1868_),
    .Y(_1870_),
    .B1(_1869_));
 sg13g2_a21o_1 _4570_ (.A2(net547),
    .A1(net757),
    .B1(_1870_),
    .X(_0156_));
 sg13g2_nor2_1 _4571_ (.A(_0019_),
    .B(_1866_),
    .Y(_1871_));
 sg13g2_a21oi_1 _4572_ (.A1(_1860_),
    .A2(_1867_),
    .Y(_1872_),
    .B1(_1871_));
 sg13g2_nand2_1 _4573_ (.Y(_1873_),
    .A(net669),
    .B(\mandelbrot.alu.in_zr[15] ));
 sg13g2_nor2_1 _4574_ (.A(_1935_),
    .B(\mandelbrot.alu.in_zr[15] ),
    .Y(_1874_));
 sg13g2_a22oi_1 _4575_ (.Y(_1875_),
    .B1(_1862_),
    .B2(_1874_),
    .A2(_1966_),
    .A1(_1935_));
 sg13g2_o21ai_1 _4576_ (.B1(_1875_),
    .Y(_1876_),
    .A1(_1862_),
    .A2(_1873_));
 sg13g2_mux2_1 _4577_ (.A0(_1864_),
    .A1(_1876_),
    .S(_1680_),
    .X(_1877_));
 sg13g2_xnor2_1 _4578_ (.Y(_1878_),
    .A(\mandelbrot.alu.m1[31] ),
    .B(_1877_));
 sg13g2_nor2_1 _4579_ (.A(_1872_),
    .B(_1878_),
    .Y(_1879_));
 sg13g2_xnor2_1 _4580_ (.Y(_1880_),
    .A(_1872_),
    .B(_1878_));
 sg13g2_nand2_1 _4581_ (.Y(_1881_),
    .A(net691),
    .B(_1967_));
 sg13g2_a22oi_1 _4582_ (.Y(_1882_),
    .B1(_1881_),
    .B2(_1706_),
    .A2(_1880_),
    .A1(net592));
 sg13g2_a21o_1 _4583_ (.A2(net547),
    .A1(net798),
    .B1(_1882_),
    .X(_0157_));
 sg13g2_and2_1 _4584_ (.A(_1967_),
    .B(_1877_),
    .X(_1883_));
 sg13g2_nor2_1 _4585_ (.A(_1879_),
    .B(_1883_),
    .Y(_1884_));
 sg13g2_nand2_1 _4586_ (.Y(_1885_),
    .A(net633),
    .B(_1875_));
 sg13g2_nand2_1 _4587_ (.Y(_1886_),
    .A(_1876_),
    .B(_1885_));
 sg13g2_xnor2_1 _4588_ (.Y(_1887_),
    .A(_1967_),
    .B(_1886_));
 sg13g2_o21ai_1 _4589_ (.B1(_1887_),
    .Y(_1888_),
    .A1(_1879_),
    .A2(_1883_));
 sg13g2_xor2_1 _4590_ (.B(_1887_),
    .A(_1884_),
    .X(_1889_));
 sg13g2_a22oi_1 _4591_ (.Y(_1890_),
    .B1(_1889_),
    .B2(net592),
    .A2(_1881_),
    .A1(_1706_));
 sg13g2_a21o_1 _4592_ (.A2(net547),
    .A1(net803),
    .B1(_1890_),
    .X(_0158_));
 sg13g2_nand3b_1 _4593_ (.B(\l_sclk[1] ),
    .C(\l_sen[2] ),
    .Y(_1891_),
    .A_N(\l_sclk[2] ));
 sg13g2_mux2_1 _4594_ (.A0(net308),
    .A1(net376),
    .S(net646),
    .X(_0159_));
 sg13g2_mux2_1 _4595_ (.A0(net247),
    .A1(net308),
    .S(net647),
    .X(_0160_));
 sg13g2_nand2_1 _4596_ (.Y(_1892_),
    .A(net247),
    .B(net649));
 sg13g2_o21ai_1 _4597_ (.B1(_1892_),
    .Y(_0161_),
    .A1(_1978_),
    .A2(net649));
 sg13g2_nor2_1 _4598_ (.A(\configuration[4] ),
    .B(net649),
    .Y(_1893_));
 sg13g2_a21oi_1 _4599_ (.A1(_1978_),
    .A2(net649),
    .Y(_0162_),
    .B1(_1893_));
 sg13g2_mux2_1 _4600_ (.A0(net349),
    .A1(\configuration[4] ),
    .S(net649),
    .X(_0163_));
 sg13g2_mux2_1 _4601_ (.A0(net390),
    .A1(net349),
    .S(net649),
    .X(_0164_));
 sg13g2_mux2_1 _4602_ (.A0(net321),
    .A1(\configuration[6] ),
    .S(net649),
    .X(_0165_));
 sg13g2_mux2_1 _4603_ (.A0(net397),
    .A1(net321),
    .S(net650),
    .X(_0166_));
 sg13g2_mux2_1 _4604_ (.A0(net335),
    .A1(\configuration[8] ),
    .S(net649),
    .X(_0167_));
 sg13g2_mux2_1 _4605_ (.A0(net326),
    .A1(\configuration[9] ),
    .S(net650),
    .X(_0168_));
 sg13g2_mux2_1 _4606_ (.A0(net310),
    .A1(net326),
    .S(net650),
    .X(_0169_));
 sg13g2_mux2_1 _4607_ (.A0(net231),
    .A1(net310),
    .S(net650),
    .X(_0170_));
 sg13g2_nand2_1 _4608_ (.Y(_1894_),
    .A(net231),
    .B(net651));
 sg13g2_o21ai_1 _4609_ (.B1(_1894_),
    .Y(_0171_),
    .A1(_1979_),
    .A2(net651));
 sg13g2_nor2_1 _4610_ (.A(net324),
    .B(net650),
    .Y(_1895_));
 sg13g2_a21oi_1 _4611_ (.A1(_1979_),
    .A2(net651),
    .Y(_0172_),
    .B1(_1895_));
 sg13g2_mux2_1 _4612_ (.A0(net344),
    .A1(net324),
    .S(net650),
    .X(_0173_));
 sg13g2_mux2_1 _4613_ (.A0(net383),
    .A1(net344),
    .S(net651),
    .X(_0174_));
 sg13g2_mux2_1 _4614_ (.A0(net424),
    .A1(net383),
    .S(net647),
    .X(_0175_));
 sg13g2_mux2_1 _4615_ (.A0(net398),
    .A1(\configuration[17] ),
    .S(net646),
    .X(_0176_));
 sg13g2_mux2_1 _4616_ (.A0(net298),
    .A1(\configuration[18] ),
    .S(net646),
    .X(_0177_));
 sg13g2_mux2_1 _4617_ (.A0(net365),
    .A1(net298),
    .S(net646),
    .X(_0178_));
 sg13g2_mux2_1 _4618_ (.A0(net389),
    .A1(net365),
    .S(net646),
    .X(_0179_));
 sg13g2_mux2_1 _4619_ (.A0(net384),
    .A1(\configuration[21] ),
    .S(net645),
    .X(_0180_));
 sg13g2_mux2_1 _4620_ (.A0(net347),
    .A1(\configuration[22] ),
    .S(net648),
    .X(_0181_));
 sg13g2_mux2_1 _4621_ (.A0(net375),
    .A1(net347),
    .S(net648),
    .X(_0182_));
 sg13g2_mux2_1 _4622_ (.A0(net342),
    .A1(\configuration[24] ),
    .S(net645),
    .X(_0183_));
 sg13g2_mux2_1 _4623_ (.A0(net368),
    .A1(net342),
    .S(net645),
    .X(_0184_));
 sg13g2_mux2_1 _4624_ (.A0(net395),
    .A1(net368),
    .S(net645),
    .X(_0185_));
 sg13g2_mux2_1 _4625_ (.A0(net353),
    .A1(\configuration[27] ),
    .S(net645),
    .X(_0186_));
 sg13g2_mux2_1 _4626_ (.A0(net355),
    .A1(net353),
    .S(net645),
    .X(_0187_));
 sg13g2_mux2_1 _4627_ (.A0(net340),
    .A1(\configuration[29] ),
    .S(net645),
    .X(_0188_));
 sg13g2_mux2_1 _4628_ (.A0(net393),
    .A1(net340),
    .S(net645),
    .X(_0189_));
 sg13g2_mux2_1 _4629_ (.A0(net719),
    .A1(net393),
    .S(net646),
    .X(_0190_));
 sg13g2_mux2_1 _4630_ (.A0(net789),
    .A1(net719),
    .S(net647),
    .X(_0191_));
 sg13g2_mux2_1 _4631_ (.A0(net790),
    .A1(net789),
    .S(net647),
    .X(_0192_));
 sg13g2_mux2_1 _4632_ (.A0(net777),
    .A1(\configuration[34] ),
    .S(net647),
    .X(_0193_));
 sg13g2_mux2_1 _4633_ (.A0(net804),
    .A1(net777),
    .S(net647),
    .X(_0194_));
 sg13g2_mux2_1 _4634_ (.A0(net801),
    .A1(\configuration[36] ),
    .S(net646),
    .X(_0195_));
 sg13g2_mux2_1 _4635_ (.A0(net799),
    .A1(net801),
    .S(net646),
    .X(_0196_));
 sg13g2_mux2_1 _4636_ (.A0(net796),
    .A1(net799),
    .S(net650),
    .X(_0197_));
 sg13g2_mux2_1 _4637_ (.A0(\configuration[40] ),
    .A1(net796),
    .S(net653),
    .X(_0198_));
 sg13g2_mux2_1 _4638_ (.A0(net775),
    .A1(\configuration[40] ),
    .S(net653),
    .X(_0199_));
 sg13g2_mux2_1 _4639_ (.A0(net333),
    .A1(\configuration[41] ),
    .S(net653),
    .X(_0200_));
 sg13g2_nand2_1 _4640_ (.Y(_1896_),
    .A(net333),
    .B(net652));
 sg13g2_o21ai_1 _4641_ (.B1(_1896_),
    .Y(_0201_),
    .A1(_1937_),
    .A2(net652));
 sg13g2_nor2_1 _4642_ (.A(net438),
    .B(net654),
    .Y(_1897_));
 sg13g2_a21oi_1 _4643_ (.A1(_1937_),
    .A2(net652),
    .Y(_0202_),
    .B1(_1897_));
 sg13g2_mux2_1 _4644_ (.A0(net480),
    .A1(net438),
    .S(net652),
    .X(_0203_));
 sg13g2_mux2_1 _4645_ (.A0(net490),
    .A1(net480),
    .S(net652),
    .X(_0204_));
 sg13g2_mux2_1 _4646_ (.A0(net302),
    .A1(\configuration[46] ),
    .S(net653),
    .X(_0205_));
 sg13g2_mux2_1 _4647_ (.A0(net437),
    .A1(net302),
    .S(net653),
    .X(_0206_));
 sg13g2_mux2_1 _4648_ (.A0(net457),
    .A1(net437),
    .S(net653),
    .X(_0207_));
 sg13g2_nand2_1 _4649_ (.Y(_1898_),
    .A(\configuration[49] ),
    .B(net653));
 sg13g2_o21ai_1 _4650_ (.B1(_1898_),
    .Y(_0208_),
    .A1(_1943_),
    .A2(net653));
 sg13g2_nor2_1 _4651_ (.A(net286),
    .B(net652),
    .Y(_1899_));
 sg13g2_a21oi_1 _4652_ (.A1(_1943_),
    .A2(net652),
    .Y(_0209_),
    .B1(_1899_));
 sg13g2_nor2_1 _4653_ (.A(net664),
    .B(net654),
    .Y(_1900_));
 sg13g2_a21oi_1 _4654_ (.A1(_1944_),
    .A2(net652),
    .Y(_0210_),
    .B1(_1900_));
 sg13g2_nor2_1 _4655_ (.A(\l_sdata[2] ),
    .B(net654),
    .Y(_1901_));
 sg13g2_a21oi_1 _4656_ (.A1(_1961_),
    .A2(net654),
    .Y(_0211_),
    .B1(_1901_));
 sg13g2_mux2_1 _4657_ (.A0(net742),
    .A1(net6),
    .S(\vga.l_read ),
    .X(_0212_));
 sg13g2_mux2_1 _4658_ (.A0(net748),
    .A1(net7),
    .S(\vga.l_read ),
    .X(_0213_));
 sg13g2_mux2_1 _4659_ (.A0(net402),
    .A1(net8),
    .S(\vga.l_read ),
    .X(_0214_));
 sg13g2_nand2_1 _4660_ (.Y(_1902_),
    .A(\vga.l_read ),
    .B(net9));
 sg13g2_o21ai_1 _4661_ (.B1(_1902_),
    .Y(_0215_),
    .A1(_1960_),
    .A2(\vga.l_read ));
 sg13g2_o21ai_1 _4662_ (.B1(_1888_),
    .Y(_1903_),
    .A1(_0017_),
    .A2(_1886_));
 sg13g2_and2_1 _4663_ (.A(_0017_),
    .B(_1875_),
    .X(_1904_));
 sg13g2_xnor2_1 _4664_ (.Y(_1905_),
    .A(_1967_),
    .B(_1875_));
 sg13g2_a221oi_1 _4665_ (.B2(_1903_),
    .C1(_1706_),
    .B1(_1905_),
    .A1(_1888_),
    .Y(_1906_),
    .A2(_1904_));
 sg13g2_nand3_1 _4666_ (.B(net566),
    .C(_1706_),
    .A(net779),
    .Y(_1907_));
 sg13g2_nand2b_1 _4667_ (.Y(_0216_),
    .B(_1907_),
    .A_N(_1906_));
 sg13g2_dfrbp_1 _4668_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net630),
    .D(net293),
    .Q_N(_0102_),
    .Q(\mandelbrot.run ));
 sg13g2_dfrbp_1 _4669_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net626),
    .D(net201),
    .Q_N(_2371_),
    .Q(reset_write_ptr));
 sg13g2_dfrbp_1 _4670_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net11),
    .D(net663),
    .Q_N(_2370_),
    .Q(l_running));
 sg13g2_dfrbp_1 _4671_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net626),
    .D(net288),
    .Q_N(_2369_),
    .Q(\vga.timing_v.pixel[0] ));
 sg13g2_dfrbp_1 _4672_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net626),
    .D(net362),
    .Q_N(_2368_),
    .Q(\vga.timing_v.pixel[1] ));
 sg13g2_dfrbp_1 _4673_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net623),
    .D(_0219_),
    .Q_N(_2367_),
    .Q(\vga.timing_v.pixel[2] ));
 sg13g2_dfrbp_1 _4674_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net624),
    .D(_0220_),
    .Q_N(_2366_),
    .Q(\vga.timing_v.pixel[3] ));
 sg13g2_dfrbp_1 _4675_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net624),
    .D(_0221_),
    .Q_N(_2365_),
    .Q(\vga.timing_v.pixel[4] ));
 sg13g2_dfrbp_1 _4676_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net624),
    .D(_0222_),
    .Q_N(_2364_),
    .Q(\vga.timing_v.pixel[5] ));
 sg13g2_dfrbp_1 _4677_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net624),
    .D(_0223_),
    .Q_N(_2363_),
    .Q(\vga.timing_v.pixel[6] ));
 sg13g2_dfrbp_1 _4678_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net623),
    .D(net357),
    .Q_N(_0101_),
    .Q(\vga.timing_v.pixel[7] ));
 sg13g2_dfrbp_1 _4679_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net623),
    .D(_0225_),
    .Q_N(_2362_),
    .Q(\vga.timing_v.pixel[8] ));
 sg13g2_dfrbp_1 _4680_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net623),
    .D(net312),
    .Q_N(_0103_),
    .Q(\vga.timing_v.pixel[9] ));
 sg13g2_dfrbp_1 _4681_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net22),
    .D(net3),
    .Q_N(_2372_),
    .Q(\l_sdata[0] ));
 sg13g2_dfrbp_1 _4682_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net23),
    .D(net200),
    .Q_N(_2373_),
    .Q(\l_sdata[1] ));
 sg13g2_dfrbp_1 _4683_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net24),
    .D(net196),
    .Q_N(_2374_),
    .Q(\l_sdata[2] ));
 sg13g2_dfrbp_1 _4684_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net25),
    .D(net4),
    .Q_N(_2375_),
    .Q(\l_sclk[0] ));
 sg13g2_dfrbp_1 _4685_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net26),
    .D(net197),
    .Q_N(_2376_),
    .Q(\l_sclk[1] ));
 sg13g2_dfrbp_1 _4686_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net27),
    .D(net195),
    .Q_N(_2377_),
    .Q(\l_sclk[2] ));
 sg13g2_dfrbp_1 _4687_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net28),
    .D(net2),
    .Q_N(_2378_),
    .Q(\l_sen[0] ));
 sg13g2_dfrbp_1 _4688_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net31),
    .D(net198),
    .Q_N(_2379_),
    .Q(\l_sen[1] ));
 sg13g2_dfrbp_1 _4689_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net152),
    .D(net202),
    .Q_N(_2361_),
    .Q(\l_sen[2] ));
 sg13g2_dfrbp_1 _4690_ (.CLK(net194),
    .RESET_B(net151),
    .D(net1),
    .Q_N(_2360_),
    .Q(latched_rst_n));
 sg13g2_dfrbp_1 _4691_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net630),
    .D(net209),
    .Q_N(\state[0] ),
    .Q(_0111_));
 sg13g2_dfrbp_1 _4692_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net630),
    .D(_0001_),
    .Q_N(_2380_),
    .Q(\state[1] ));
 sg13g2_dfrbp_1 _4693_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net630),
    .D(net205),
    .Q_N(_2381_),
    .Q(\state[2] ));
 sg13g2_dfrbp_1 _4694_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net626),
    .D(net283),
    .Q_N(_2359_),
    .Q(\state[3] ));
 sg13g2_dfrbp_1 _4695_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net620),
    .D(_0227_),
    .Q_N(_2358_),
    .Q(\mandelbrot.alu.mult_zi_zi.shift_reg[0] ));
 sg13g2_dfrbp_1 _4696_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net617),
    .D(_0228_),
    .Q_N(_2357_),
    .Q(\mandelbrot.alu.m2[0] ));
 sg13g2_dfrbp_1 _4697_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net619),
    .D(net788),
    .Q_N(_2356_),
    .Q(\mandelbrot.alu.m2[1] ));
 sg13g2_dfrbp_1 _4698_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net617),
    .D(_0230_),
    .Q_N(_2355_),
    .Q(\mandelbrot.alu.m2[2] ));
 sg13g2_dfrbp_1 _4699_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net617),
    .D(_0231_),
    .Q_N(_2354_),
    .Q(\mandelbrot.alu.m2[3] ));
 sg13g2_dfrbp_1 _4700_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net617),
    .D(net737),
    .Q_N(_2353_),
    .Q(\mandelbrot.alu.m2[4] ));
 sg13g2_dfrbp_1 _4701_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net617),
    .D(net711),
    .Q_N(_2352_),
    .Q(\mandelbrot.alu.m2[5] ));
 sg13g2_dfrbp_1 _4702_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net617),
    .D(net761),
    .Q_N(_2351_),
    .Q(\mandelbrot.alu.m2[6] ));
 sg13g2_dfrbp_1 _4703_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net617),
    .D(_0235_),
    .Q_N(_2350_),
    .Q(\mandelbrot.alu.m2[7] ));
 sg13g2_dfrbp_1 _4704_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net616),
    .D(_0236_),
    .Q_N(_2349_),
    .Q(\mandelbrot.alu.m2[8] ));
 sg13g2_dfrbp_1 _4705_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net616),
    .D(net528),
    .Q_N(_2348_),
    .Q(\mandelbrot.alu.m2[9] ));
 sg13g2_dfrbp_1 _4706_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net616),
    .D(_0238_),
    .Q_N(_2347_),
    .Q(\mandelbrot.alu.m2[10] ));
 sg13g2_dfrbp_1 _4707_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net616),
    .D(net741),
    .Q_N(_2346_),
    .Q(\mandelbrot.alu.m2[11] ));
 sg13g2_dfrbp_1 _4708_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net616),
    .D(_0240_),
    .Q_N(_2345_),
    .Q(\mandelbrot.alu.m2[12] ));
 sg13g2_dfrbp_1 _4709_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net616),
    .D(net745),
    .Q_N(_2344_),
    .Q(\mandelbrot.alu.m2[13] ));
 sg13g2_dfrbp_1 _4710_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net615),
    .D(_0242_),
    .Q_N(_2343_),
    .Q(\mandelbrot.alu.m2[14] ));
 sg13g2_dfrbp_1 _4711_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net620),
    .D(_0243_),
    .Q_N(_2342_),
    .Q(\mandelbrot.alu.m2[15] ));
 sg13g2_dfrbp_1 _4712_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net620),
    .D(_0244_),
    .Q_N(_2341_),
    .Q(\mandelbrot.alu.m2[16] ));
 sg13g2_dfrbp_1 _4713_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net620),
    .D(_0245_),
    .Q_N(_2340_),
    .Q(\mandelbrot.alu.m2[17] ));
 sg13g2_dfrbp_1 _4714_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net615),
    .D(net813),
    .Q_N(_0100_),
    .Q(\mandelbrot.alu.m2[18] ));
 sg13g2_dfrbp_1 _4715_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net621),
    .D(net808),
    .Q_N(_0099_),
    .Q(\mandelbrot.alu.m2[19] ));
 sg13g2_dfrbp_1 _4716_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net615),
    .D(net718),
    .Q_N(_0098_),
    .Q(\mandelbrot.alu.m2[20] ));
 sg13g2_dfrbp_1 _4717_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net615),
    .D(net268),
    .Q_N(_0097_),
    .Q(\mandelbrot.alu.m2[21] ));
 sg13g2_dfrbp_1 _4718_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net615),
    .D(_0250_),
    .Q_N(_0096_),
    .Q(\mandelbrot.alu.m2[22] ));
 sg13g2_dfrbp_1 _4719_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net614),
    .D(net747),
    .Q_N(_2339_),
    .Q(\mandelbrot.alu.m2[23] ));
 sg13g2_dfrbp_1 _4720_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net615),
    .D(net464),
    .Q_N(_0095_),
    .Q(\mandelbrot.alu.m2[24] ));
 sg13g2_dfrbp_1 _4721_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net614),
    .D(_0253_),
    .Q_N(_0094_),
    .Q(\mandelbrot.alu.m2[25] ));
 sg13g2_dfrbp_1 _4722_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net614),
    .D(_0254_),
    .Q_N(_0093_),
    .Q(\mandelbrot.alu.m2[26] ));
 sg13g2_dfrbp_1 _4723_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net614),
    .D(_0255_),
    .Q_N(_2338_),
    .Q(\mandelbrot.alu.m2[27] ));
 sg13g2_dfrbp_1 _4724_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net614),
    .D(_0256_),
    .Q_N(_0092_),
    .Q(\mandelbrot.alu.m2[28] ));
 sg13g2_dfrbp_1 _4725_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net614),
    .D(_0257_),
    .Q_N(_0091_),
    .Q(\mandelbrot.alu.m2[29] ));
 sg13g2_dfrbp_1 _4726_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net614),
    .D(_0258_),
    .Q_N(_0090_),
    .Q(\mandelbrot.alu.m2[30] ));
 sg13g2_dfrbp_1 _4727_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net150),
    .D(net207),
    .Q_N(_0089_),
    .Q(\mandelbrot.alu.mult_zr_zi.ctr[0] ));
 sg13g2_dfrbp_1 _4728_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net149),
    .D(net229),
    .Q_N(_2337_),
    .Q(\mandelbrot.alu.mult_zr_zi.ctr[1] ));
 sg13g2_dfrbp_1 _4729_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net148),
    .D(net262),
    .Q_N(_2336_),
    .Q(\mandelbrot.alu.mult_zr_zi.ctr[2] ));
 sg13g2_dfrbp_1 _4730_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net147),
    .D(net211),
    .Q_N(_0088_),
    .Q(\mandelbrot.alu.mult_zr_zr.ctr[0] ));
 sg13g2_dfrbp_1 _4731_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net146),
    .D(net242),
    .Q_N(_2335_),
    .Q(\mandelbrot.alu.mult_zr_zr.ctr[1] ));
 sg13g2_dfrbp_1 _4732_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net145),
    .D(net254),
    .Q_N(_2334_),
    .Q(\mandelbrot.alu.mult_zr_zr.ctr[2] ));
 sg13g2_dfrbp_1 _4733_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net610),
    .D(_0265_),
    .Q_N(_2333_),
    .Q(\mandelbrot.alu.mult_zr_zi.shift_reg[0] ));
 sg13g2_dfrbp_1 _4734_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net618),
    .D(net234),
    .Q_N(_2332_),
    .Q(\mandelbrot.alu.m3[0] ));
 sg13g2_dfrbp_1 _4735_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net618),
    .D(_0267_),
    .Q_N(_2331_),
    .Q(\mandelbrot.alu.m3[1] ));
 sg13g2_dfrbp_1 _4736_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net612),
    .D(_0268_),
    .Q_N(_2330_),
    .Q(\mandelbrot.alu.m3[2] ));
 sg13g2_dfrbp_1 _4737_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net618),
    .D(net244),
    .Q_N(_2329_),
    .Q(\mandelbrot.alu.m3[3] ));
 sg13g2_dfrbp_1 _4738_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net612),
    .D(_0270_),
    .Q_N(_2328_),
    .Q(\mandelbrot.alu.m3[4] ));
 sg13g2_dfrbp_1 _4739_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net627),
    .D(_0271_),
    .Q_N(_2327_),
    .Q(\mandelbrot.alu.m3[5] ));
 sg13g2_dfrbp_1 _4740_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net627),
    .D(_0272_),
    .Q_N(_2326_),
    .Q(\mandelbrot.alu.m3[6] ));
 sg13g2_dfrbp_1 _4741_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net628),
    .D(_0273_),
    .Q_N(_2325_),
    .Q(\mandelbrot.alu.m3[7] ));
 sg13g2_dfrbp_1 _4742_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net627),
    .D(net339),
    .Q_N(_2324_),
    .Q(\mandelbrot.alu.m3[8] ));
 sg13g2_dfrbp_1 _4743_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net628),
    .D(net301),
    .Q_N(_2323_),
    .Q(\mandelbrot.alu.m3[9] ));
 sg13g2_dfrbp_1 _4744_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net612),
    .D(_0276_),
    .Q_N(_2322_),
    .Q(\mandelbrot.alu.m3[10] ));
 sg13g2_dfrbp_1 _4745_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net611),
    .D(_0277_),
    .Q_N(_2321_),
    .Q(\mandelbrot.alu.m3[11] ));
 sg13g2_dfrbp_1 _4746_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net612),
    .D(net370),
    .Q_N(_2320_),
    .Q(\mandelbrot.alu.m3[12] ));
 sg13g2_dfrbp_1 _4747_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net611),
    .D(_0279_),
    .Q_N(_2319_),
    .Q(\mandelbrot.alu.m3[13] ));
 sg13g2_dfrbp_1 _4748_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net611),
    .D(net730),
    .Q_N(_2318_),
    .Q(\mandelbrot.alu.m3[14] ));
 sg13g2_dfrbp_1 _4749_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net611),
    .D(_0281_),
    .Q_N(_2317_),
    .Q(\mandelbrot.alu.m3[15] ));
 sg13g2_dfrbp_1 _4750_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net611),
    .D(net405),
    .Q_N(_2316_),
    .Q(\mandelbrot.alu.m3[16] ));
 sg13g2_dfrbp_1 _4751_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net611),
    .D(_0283_),
    .Q_N(_2315_),
    .Q(\mandelbrot.alu.m3[17] ));
 sg13g2_dfrbp_1 _4752_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net611),
    .D(_0284_),
    .Q_N(_0087_),
    .Q(\mandelbrot.alu.m3[18] ));
 sg13g2_dfrbp_1 _4753_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net610),
    .D(net530),
    .Q_N(_0086_),
    .Q(\mandelbrot.alu.m3[19] ));
 sg13g2_dfrbp_1 _4754_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net610),
    .D(_0286_),
    .Q_N(_0085_),
    .Q(\mandelbrot.alu.m3[20] ));
 sg13g2_dfrbp_1 _4755_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net610),
    .D(net502),
    .Q_N(_0084_),
    .Q(\mandelbrot.alu.m3[21] ));
 sg13g2_dfrbp_1 _4756_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net610),
    .D(net416),
    .Q_N(_0083_),
    .Q(\mandelbrot.alu.m3[22] ));
 sg13g2_dfrbp_1 _4757_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net609),
    .D(net754),
    .Q_N(_2314_),
    .Q(\mandelbrot.alu.m3[23] ));
 sg13g2_dfrbp_1 _4758_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net609),
    .D(net414),
    .Q_N(_0082_),
    .Q(\mandelbrot.alu.m3[24] ));
 sg13g2_dfrbp_1 _4759_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net609),
    .D(net475),
    .Q_N(_0081_),
    .Q(\mandelbrot.alu.m3[25] ));
 sg13g2_dfrbp_1 _4760_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net609),
    .D(net387),
    .Q_N(_0080_),
    .Q(\mandelbrot.alu.m3[26] ));
 sg13g2_dfrbp_1 _4761_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net609),
    .D(net330),
    .Q_N(_2313_),
    .Q(\mandelbrot.alu.m3[27] ));
 sg13g2_dfrbp_1 _4762_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net609),
    .D(_0294_),
    .Q_N(_0079_),
    .Q(\mandelbrot.alu.m3[28] ));
 sg13g2_dfrbp_1 _4763_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net609),
    .D(_0295_),
    .Q_N(_0078_),
    .Q(\mandelbrot.alu.m3[29] ));
 sg13g2_dfrbp_1 _4764_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net609),
    .D(_0296_),
    .Q_N(_0104_),
    .Q(\mandelbrot.alu.m3[30] ));
 sg13g2_dfrbp_1 _4765_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net629),
    .D(net806),
    .Q_N(\mandelbrot.alu.finished ),
    .Q(\mandelbrot.alu.mult_zr_zr.running ));
 sg13g2_dfrbp_1 _4766_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net144),
    .D(net216),
    .Q_N(_0077_),
    .Q(\mandelbrot.alu.mult_zi_zi.ctr[0] ));
 sg13g2_dfrbp_1 _4767_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net143),
    .D(net237),
    .Q_N(_2312_),
    .Q(\mandelbrot.alu.mult_zi_zi.ctr[1] ));
 sg13g2_dfrbp_1 _4768_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net105),
    .D(net278),
    .Q_N(_2382_),
    .Q(\mandelbrot.alu.mult_zi_zi.ctr[2] ));
 sg13g2_dfrbp_1 _4769_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net615),
    .D(_0003_),
    .Q_N(_0076_),
    .Q(\mandelbrot.alu.mult_zi_zi.running ));
 sg13g2_dfrbp_1 _4770_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net614),
    .D(net819),
    .Q_N(_0105_),
    .Q(\mandelbrot.alu.m2[31] ));
 sg13g2_dfrbp_1 _4771_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net610),
    .D(_0004_),
    .Q_N(_0075_),
    .Q(\mandelbrot.alu.mult_zr_zi.running ));
 sg13g2_dfrbp_1 _4772_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net630),
    .D(_0116_),
    .Q_N(\mandelbrot.alu.first_iteration ),
    .Q(_0112_));
 sg13g2_dfrbp_1 _4773_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net142),
    .D(_0301_),
    .Q_N(_0074_),
    .Q(\mandelbrot.alu.in_zr[0] ));
 sg13g2_dfrbp_1 _4774_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net141),
    .D(_0302_),
    .Q_N(_0073_),
    .Q(\mandelbrot.alu.in_zr[1] ));
 sg13g2_dfrbp_1 _4775_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net140),
    .D(_0303_),
    .Q_N(_0072_),
    .Q(\mandelbrot.alu.in_zr[2] ));
 sg13g2_dfrbp_1 _4776_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net139),
    .D(_0304_),
    .Q_N(_0071_),
    .Q(\mandelbrot.alu.in_zr[3] ));
 sg13g2_dfrbp_1 _4777_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net138),
    .D(_0305_),
    .Q_N(_0070_),
    .Q(\mandelbrot.alu.in_zr[4] ));
 sg13g2_dfrbp_1 _4778_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net136),
    .D(_0306_),
    .Q_N(_0069_),
    .Q(\mandelbrot.alu.in_zr[5] ));
 sg13g2_dfrbp_1 _4779_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net134),
    .D(_0307_),
    .Q_N(_0068_),
    .Q(\mandelbrot.alu.in_zr[6] ));
 sg13g2_dfrbp_1 _4780_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net132),
    .D(_0308_),
    .Q_N(_0067_),
    .Q(\mandelbrot.alu.in_zr[7] ));
 sg13g2_dfrbp_1 _4781_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net130),
    .D(_0309_),
    .Q_N(_0066_),
    .Q(\mandelbrot.alu.in_zr[8] ));
 sg13g2_dfrbp_1 _4782_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net128),
    .D(_0310_),
    .Q_N(_0065_),
    .Q(\mandelbrot.alu.in_zr[9] ));
 sg13g2_dfrbp_1 _4783_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net126),
    .D(_0311_),
    .Q_N(_0064_),
    .Q(\mandelbrot.alu.in_zr[10] ));
 sg13g2_dfrbp_1 _4784_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net124),
    .D(_0312_),
    .Q_N(_0063_),
    .Q(\mandelbrot.alu.in_zr[11] ));
 sg13g2_dfrbp_1 _4785_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net122),
    .D(net382),
    .Q_N(_0062_),
    .Q(\mandelbrot.alu.in_zr[12] ));
 sg13g2_dfrbp_1 _4786_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net120),
    .D(_0314_),
    .Q_N(_0061_),
    .Q(\mandelbrot.alu.in_zr[13] ));
 sg13g2_dfrbp_1 _4787_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net118),
    .D(_0315_),
    .Q_N(_0060_),
    .Q(\mandelbrot.alu.in_zr[14] ));
 sg13g2_dfrbp_1 _4788_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net116),
    .D(_0316_),
    .Q_N(_0059_),
    .Q(\mandelbrot.alu.in_zr[15] ));
 sg13g2_dfrbp_1 _4789_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net114),
    .D(_0317_),
    .Q_N(_2311_),
    .Q(\mandelbrot.alu.in_ci[0] ));
 sg13g2_dfrbp_1 _4790_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net113),
    .D(_0318_),
    .Q_N(_2310_),
    .Q(\mandelbrot.alu.in_ci[1] ));
 sg13g2_dfrbp_1 _4791_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net112),
    .D(_0319_),
    .Q_N(_2309_),
    .Q(\mandelbrot.alu.in_ci[2] ));
 sg13g2_dfrbp_1 _4792_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net111),
    .D(_0320_),
    .Q_N(_2308_),
    .Q(\mandelbrot.alu.in_ci[3] ));
 sg13g2_dfrbp_1 _4793_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net110),
    .D(_0321_),
    .Q_N(_2307_),
    .Q(\mandelbrot.alu.in_ci[4] ));
 sg13g2_dfrbp_1 _4794_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net109),
    .D(_0322_),
    .Q_N(_2306_),
    .Q(\mandelbrot.alu.in_ci[5] ));
 sg13g2_dfrbp_1 _4795_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net108),
    .D(_0323_),
    .Q_N(_2305_),
    .Q(\mandelbrot.alu.in_ci[6] ));
 sg13g2_dfrbp_1 _4796_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net107),
    .D(net373),
    .Q_N(_0058_),
    .Q(\mandelbrot.alu.in_ci[7] ));
 sg13g2_dfrbp_1 _4797_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net106),
    .D(_0325_),
    .Q_N(_2304_),
    .Q(\mandelbrot.alu.in_ci[8] ));
 sg13g2_dfrbp_1 _4798_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net104),
    .D(_0326_),
    .Q_N(_2303_),
    .Q(\mandelbrot.alu.in_ci[9] ));
 sg13g2_dfrbp_1 _4799_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net103),
    .D(_0327_),
    .Q_N(_2302_),
    .Q(\mandelbrot.alu.in_ci[10] ));
 sg13g2_dfrbp_1 _4800_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net102),
    .D(_0328_),
    .Q_N(_2301_),
    .Q(\mandelbrot.alu.in_ci[11] ));
 sg13g2_dfrbp_1 _4801_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net101),
    .D(_0329_),
    .Q_N(_2300_),
    .Q(\mandelbrot.alu.in_ci[12] ));
 sg13g2_dfrbp_1 _4802_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net100),
    .D(_0330_),
    .Q_N(_2299_),
    .Q(\mandelbrot.alu.in_ci[13] ));
 sg13g2_dfrbp_1 _4803_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net99),
    .D(_0331_),
    .Q_N(_2298_),
    .Q(\mandelbrot.alu.in_ci[14] ));
 sg13g2_dfrbp_1 _4804_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net98),
    .D(_0332_),
    .Q_N(_2297_),
    .Q(\mandelbrot.alu.in_ci[15] ));
 sg13g2_dfrbp_1 _4805_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net97),
    .D(net218),
    .Q_N(_0057_),
    .Q(\mandelbrot.ctr[0] ));
 sg13g2_dfrbp_1 _4806_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net95),
    .D(net723),
    .Q_N(_2296_),
    .Q(\mandelbrot.ctr[1] ));
 sg13g2_dfrbp_1 _4807_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net93),
    .D(_0335_),
    .Q_N(_2295_),
    .Q(\mandelbrot.ctr[2] ));
 sg13g2_dfrbp_1 _4808_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net91),
    .D(_0336_),
    .Q_N(_2294_),
    .Q(\mandelbrot.ctr[3] ));
 sg13g2_dfrbp_1 _4809_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net89),
    .D(_0337_),
    .Q_N(_2293_),
    .Q(\mandelbrot.ctr[4] ));
 sg13g2_dfrbp_1 _4810_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net87),
    .D(_0338_),
    .Q_N(_2292_),
    .Q(\mandelbrot.ctr[5] ));
 sg13g2_dfrbp_1 _4811_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net85),
    .D(_0339_),
    .Q_N(_2291_),
    .Q(\mandelbrot.ctr[6] ));
 sg13g2_dfrbp_1 _4812_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net83),
    .D(_0340_),
    .Q_N(_2290_),
    .Q(\mandelbrot.ctr[7] ));
 sg13g2_dfrbp_1 _4813_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net81),
    .D(_0341_),
    .Q_N(_2289_),
    .Q(\mandelbrot.ctr[8] ));
 sg13g2_dfrbp_1 _4814_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net79),
    .D(_0342_),
    .Q_N(_2288_),
    .Q(\mandelbrot.ctr[9] ));
 sg13g2_dfrbp_1 _4815_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net77),
    .D(_0343_),
    .Q_N(_2287_),
    .Q(\mandelbrot.alu.in_cr[0] ));
 sg13g2_dfrbp_1 _4816_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net76),
    .D(net309),
    .Q_N(_0056_),
    .Q(\mandelbrot.alu.in_cr[1] ));
 sg13g2_dfrbp_1 _4817_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net75),
    .D(_0345_),
    .Q_N(_2286_),
    .Q(\mandelbrot.alu.in_cr[2] ));
 sg13g2_dfrbp_1 _4818_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net74),
    .D(_0346_),
    .Q_N(_0055_),
    .Q(\mandelbrot.alu.in_cr[3] ));
 sg13g2_dfrbp_1 _4819_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net73),
    .D(net766),
    .Q_N(_2285_),
    .Q(\mandelbrot.alu.in_cr[4] ));
 sg13g2_dfrbp_1 _4820_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net72),
    .D(_0348_),
    .Q_N(_0054_),
    .Q(\mandelbrot.alu.in_cr[5] ));
 sg13g2_dfrbp_1 _4821_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net71),
    .D(_0349_),
    .Q_N(_2284_),
    .Q(\mandelbrot.alu.in_cr[6] ));
 sg13g2_dfrbp_1 _4822_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net70),
    .D(net226),
    .Q_N(_0053_),
    .Q(\mandelbrot.alu.in_cr[7] ));
 sg13g2_dfrbp_1 _4823_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net69),
    .D(net443),
    .Q_N(_0052_),
    .Q(\mandelbrot.alu.in_cr[8] ));
 sg13g2_dfrbp_1 _4824_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net68),
    .D(_0352_),
    .Q_N(_0051_),
    .Q(\mandelbrot.alu.in_cr[9] ));
 sg13g2_dfrbp_1 _4825_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net67),
    .D(net466),
    .Q_N(_2283_),
    .Q(\mandelbrot.alu.in_cr[10] ));
 sg13g2_dfrbp_1 _4826_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net66),
    .D(net714),
    .Q_N(_2282_),
    .Q(\mandelbrot.alu.in_cr[11] ));
 sg13g2_dfrbp_1 _4827_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net65),
    .D(_0355_),
    .Q_N(_2281_),
    .Q(\mandelbrot.alu.in_cr[12] ));
 sg13g2_dfrbp_1 _4828_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net64),
    .D(net521),
    .Q_N(_2280_),
    .Q(\mandelbrot.alu.in_cr[13] ));
 sg13g2_dfrbp_1 _4829_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net63),
    .D(_0357_),
    .Q_N(_0050_),
    .Q(\mandelbrot.alu.in_cr[14] ));
 sg13g2_dfrbp_1 _4830_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net62),
    .D(net721),
    .Q_N(_0049_),
    .Q(\mandelbrot.alu.in_cr[15] ));
 sg13g2_dfrbp_1 _4831_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net630),
    .D(_0359_),
    .Q_N(finished),
    .Q(_0113_));
 sg13g2_dfrbp_1 _4832_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net59),
    .D(_0360_),
    .Q_N(_2279_),
    .Q(uio_out[0]));
 sg13g2_dfrbp_1 _4833_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net58),
    .D(_0361_),
    .Q_N(_2278_),
    .Q(uio_out[1]));
 sg13g2_dfrbp_1 _4834_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net57),
    .D(net504),
    .Q_N(_2277_),
    .Q(uio_out[2]));
 sg13g2_dfrbp_1 _4835_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net56),
    .D(_0363_),
    .Q_N(_2276_),
    .Q(uio_out[3]));
 sg13g2_dfrbp_1 _4836_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net55),
    .D(_0364_),
    .Q_N(_2275_),
    .Q(\mandelbrot.overflowed ));
 sg13g2_dfrbp_1 _4837_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net53),
    .D(net213),
    .Q_N(_0048_),
    .Q(\mandelbrot.x[0] ));
 sg13g2_dfrbp_1 _4838_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net51),
    .D(net251),
    .Q_N(_2274_),
    .Q(\mandelbrot.x[1] ));
 sg13g2_dfrbp_1 _4839_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net49),
    .D(net434),
    .Q_N(_2273_),
    .Q(\mandelbrot.x[2] ));
 sg13g2_dfrbp_1 _4840_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net47),
    .D(net266),
    .Q_N(_2272_),
    .Q(\mandelbrot.x[3] ));
 sg13g2_dfrbp_1 _4841_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net45),
    .D(_0369_),
    .Q_N(_2271_),
    .Q(\mandelbrot.x[4] ));
 sg13g2_dfrbp_1 _4842_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net43),
    .D(net455),
    .Q_N(_2270_),
    .Q(\mandelbrot.x[5] ));
 sg13g2_dfrbp_1 _4843_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net41),
    .D(net307),
    .Q_N(_2269_),
    .Q(\mandelbrot.x[6] ));
 sg13g2_dfrbp_1 _4844_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net39),
    .D(_0372_),
    .Q_N(_2268_),
    .Q(\mandelbrot.x[7] ));
 sg13g2_dfrbp_1 _4845_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net37),
    .D(_0373_),
    .Q_N(_2267_),
    .Q(\mandelbrot.x[8] ));
 sg13g2_dfrbp_1 _4846_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net35),
    .D(_0374_),
    .Q_N(_0047_),
    .Q(\mandelbrot.alu.in_zi[0] ));
 sg13g2_dfrbp_1 _4847_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net33),
    .D(net423),
    .Q_N(_0046_),
    .Q(\mandelbrot.alu.in_zi[1] ));
 sg13g2_dfrbp_1 _4848_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net30),
    .D(_0376_),
    .Q_N(_0045_),
    .Q(\mandelbrot.alu.in_zi[2] ));
 sg13g2_dfrbp_1 _4849_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net21),
    .D(_0377_),
    .Q_N(_0044_),
    .Q(\mandelbrot.alu.in_zi[3] ));
 sg13g2_dfrbp_1 _4850_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net19),
    .D(_0378_),
    .Q_N(_0043_),
    .Q(\mandelbrot.alu.in_zi[4] ));
 sg13g2_dfrbp_1 _4851_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net17),
    .D(_0379_),
    .Q_N(_0042_),
    .Q(\mandelbrot.alu.in_zi[5] ));
 sg13g2_dfrbp_1 _4852_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net15),
    .D(_0380_),
    .Q_N(_0041_),
    .Q(\mandelbrot.alu.in_zi[6] ));
 sg13g2_dfrbp_1 _4853_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net13),
    .D(_0381_),
    .Q_N(_0040_),
    .Q(\mandelbrot.alu.in_zi[7] ));
 sg13g2_dfrbp_1 _4854_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net10),
    .D(_0382_),
    .Q_N(_0039_),
    .Q(\mandelbrot.alu.in_zi[8] ));
 sg13g2_dfrbp_1 _4855_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net182),
    .D(_0383_),
    .Q_N(_0038_),
    .Q(\mandelbrot.alu.in_zi[9] ));
 sg13g2_dfrbp_1 _4856_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net180),
    .D(_0384_),
    .Q_N(_0037_),
    .Q(\mandelbrot.alu.in_zi[10] ));
 sg13g2_dfrbp_1 _4857_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net178),
    .D(_0385_),
    .Q_N(_0036_),
    .Q(\mandelbrot.alu.in_zi[11] ));
 sg13g2_dfrbp_1 _4858_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net176),
    .D(_0386_),
    .Q_N(_0035_),
    .Q(\mandelbrot.alu.in_zi[12] ));
 sg13g2_dfrbp_1 _4859_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net174),
    .D(_0387_),
    .Q_N(_0034_),
    .Q(\mandelbrot.alu.in_zi[13] ));
 sg13g2_dfrbp_1 _4860_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net172),
    .D(_0388_),
    .Q_N(_0033_),
    .Q(\mandelbrot.alu.in_zi[14] ));
 sg13g2_dfrbp_1 _4861_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net170),
    .D(_0389_),
    .Q_N(_0032_),
    .Q(\mandelbrot.alu.in_zi[15] ));
 sg13g2_dfrbp_1 _4862_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net168),
    .D(net220),
    .Q_N(_0031_),
    .Q(\mandelbrot.y[0] ));
 sg13g2_dfrbp_1 _4863_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net166),
    .D(net430),
    .Q_N(_2266_),
    .Q(\mandelbrot.y[1] ));
 sg13g2_dfrbp_1 _4864_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net164),
    .D(net411),
    .Q_N(_2265_),
    .Q(\mandelbrot.y[2] ));
 sg13g2_dfrbp_1 _4865_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net162),
    .D(_0120_),
    .Q_N(_2264_),
    .Q(\mandelbrot.y[3] ));
 sg13g2_dfrbp_1 _4866_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net160),
    .D(net257),
    .Q_N(_2263_),
    .Q(\mandelbrot.y[4] ));
 sg13g2_dfrbp_1 _4867_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net158),
    .D(net484),
    .Q_N(_2262_),
    .Q(\mandelbrot.y[5] ));
 sg13g2_dfrbp_1 _4868_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net156),
    .D(net419),
    .Q_N(_2261_),
    .Q(\mandelbrot.y[6] ));
 sg13g2_dfrbp_1 _4869_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net154),
    .D(net489),
    .Q_N(_2260_),
    .Q(\mandelbrot.y[7] ));
 sg13g2_dfrbp_1 _4870_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net183),
    .D(net285),
    .Q_N(_2383_),
    .Q(\mandelbrot.y[8] ));
 sg13g2_dfrbp_1 _4871_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net629),
    .D(net203),
    .Q_N(_2259_),
    .Q(\mandelbrot.l_alu_finished ));
 sg13g2_dfrbp_1 _4872_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net616),
    .D(_0126_),
    .Q_N(_0030_),
    .Q(\mandelbrot.alu.m3[31] ));
 sg13g2_dfrbp_1 _4873_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net620),
    .D(_0127_),
    .Q_N(_2258_),
    .Q(\mandelbrot.alu.mult_zr_zr.shift_reg[0] ));
 sg13g2_dfrbp_1 _4874_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net620),
    .D(net500),
    .Q_N(_2257_),
    .Q(\mandelbrot.alu.m1[0] ));
 sg13g2_dfrbp_1 _4875_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net628),
    .D(_0129_),
    .Q_N(_2256_),
    .Q(\mandelbrot.alu.m1[1] ));
 sg13g2_dfrbp_1 _4876_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net617),
    .D(_0130_),
    .Q_N(_2255_),
    .Q(\mandelbrot.alu.m1[2] ));
 sg13g2_dfrbp_1 _4877_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net618),
    .D(net514),
    .Q_N(_2254_),
    .Q(\mandelbrot.alu.m1[3] ));
 sg13g2_dfrbp_1 _4878_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net618),
    .D(_0132_),
    .Q_N(_2253_),
    .Q(\mandelbrot.alu.m1[4] ));
 sg13g2_dfrbp_1 _4879_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net628),
    .D(_0133_),
    .Q_N(_2252_),
    .Q(\mandelbrot.alu.m1[5] ));
 sg13g2_dfrbp_1 _4880_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net618),
    .D(_0134_),
    .Q_N(_2251_),
    .Q(\mandelbrot.alu.m1[6] ));
 sg13g2_dfrbp_1 _4881_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net618),
    .D(_0135_),
    .Q_N(_2250_),
    .Q(\mandelbrot.alu.m1[7] ));
 sg13g2_dfrbp_1 _4882_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net619),
    .D(_0136_),
    .Q_N(_2249_),
    .Q(\mandelbrot.alu.m1[8] ));
 sg13g2_dfrbp_1 _4883_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net619),
    .D(net471),
    .Q_N(_2248_),
    .Q(\mandelbrot.alu.m1[9] ));
 sg13g2_dfrbp_1 _4884_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net628),
    .D(_0138_),
    .Q_N(_2247_),
    .Q(\mandelbrot.alu.m1[10] ));
 sg13g2_dfrbp_1 _4885_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net618),
    .D(_0139_),
    .Q_N(_2246_),
    .Q(\mandelbrot.alu.m1[11] ));
 sg13g2_dfrbp_1 _4886_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net621),
    .D(net524),
    .Q_N(_2245_),
    .Q(\mandelbrot.alu.m1[12] ));
 sg13g2_dfrbp_1 _4887_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net622),
    .D(_0141_),
    .Q_N(_2244_),
    .Q(\mandelbrot.alu.m1[13] ));
 sg13g2_dfrbp_1 _4888_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net621),
    .D(_0142_),
    .Q_N(_2243_),
    .Q(\mandelbrot.alu.m1[14] ));
 sg13g2_dfrbp_1 _4889_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net620),
    .D(_0143_),
    .Q_N(_2242_),
    .Q(\mandelbrot.alu.m1[15] ));
 sg13g2_dfrbp_1 _4890_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net621),
    .D(_0144_),
    .Q_N(_2241_),
    .Q(\mandelbrot.alu.m1[16] ));
 sg13g2_dfrbp_1 _4891_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net621),
    .D(_0145_),
    .Q_N(_2240_),
    .Q(\mandelbrot.alu.m1[17] ));
 sg13g2_dfrbp_1 _4892_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net621),
    .D(_0146_),
    .Q_N(_0029_),
    .Q(\mandelbrot.alu.m1[18] ));
 sg13g2_dfrbp_1 _4893_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net621),
    .D(_0147_),
    .Q_N(_0028_),
    .Q(\mandelbrot.alu.m1[19] ));
 sg13g2_dfrbp_1 _4894_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net631),
    .D(_0148_),
    .Q_N(_0027_),
    .Q(\mandelbrot.alu.m1[20] ));
 sg13g2_dfrbp_1 _4895_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net631),
    .D(net462),
    .Q_N(_0026_),
    .Q(\mandelbrot.alu.m1[21] ));
 sg13g2_dfrbp_1 _4896_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net628),
    .D(_0150_),
    .Q_N(_0025_),
    .Q(\mandelbrot.alu.m1[22] ));
 sg13g2_dfrbp_1 _4897_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net628),
    .D(net756),
    .Q_N(_2239_),
    .Q(\mandelbrot.alu.m1[23] ));
 sg13g2_dfrbp_1 _4898_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net628),
    .D(net367),
    .Q_N(_0024_),
    .Q(\mandelbrot.alu.m1[24] ));
 sg13g2_dfrbp_1 _4899_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net630),
    .D(_0153_),
    .Q_N(_0023_),
    .Q(\mandelbrot.alu.m1[25] ));
 sg13g2_dfrbp_1 _4900_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net629),
    .D(_0154_),
    .Q_N(_0022_),
    .Q(\mandelbrot.alu.m1[26] ));
 sg13g2_dfrbp_1 _4901_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net629),
    .D(net770),
    .Q_N(_2238_),
    .Q(\mandelbrot.alu.m1[27] ));
 sg13g2_dfrbp_1 _4902_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net629),
    .D(net758),
    .Q_N(_0021_),
    .Q(\mandelbrot.alu.m1[28] ));
 sg13g2_dfrbp_1 _4903_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net629),
    .D(_0157_),
    .Q_N(_0020_),
    .Q(\mandelbrot.alu.m1[29] ));
 sg13g2_dfrbp_1 _4904_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net629),
    .D(_0158_),
    .Q_N(_0019_),
    .Q(\mandelbrot.alu.m1[30] ));
 sg13g2_dfrbp_1 _4905_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net137),
    .D(_0159_),
    .Q_N(_2237_),
    .Q(\configuration[0] ));
 sg13g2_dfrbp_1 _4906_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net135),
    .D(_0160_),
    .Q_N(_2236_),
    .Q(\configuration[1] ));
 sg13g2_dfrbp_1 _4907_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net133),
    .D(net248),
    .Q_N(_2235_),
    .Q(\configuration[2] ));
 sg13g2_dfrbp_1 _4908_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net131),
    .D(net316),
    .Q_N(_2234_),
    .Q(\configuration[3] ));
 sg13g2_dfrbp_1 _4909_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net129),
    .D(net350),
    .Q_N(_2233_),
    .Q(\configuration[4] ));
 sg13g2_dfrbp_1 _4910_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net127),
    .D(_0164_),
    .Q_N(_2232_),
    .Q(\configuration[5] ));
 sg13g2_dfrbp_1 _4911_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net125),
    .D(net322),
    .Q_N(_2231_),
    .Q(\configuration[6] ));
 sg13g2_dfrbp_1 _4912_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net123),
    .D(_0166_),
    .Q_N(_2230_),
    .Q(\configuration[7] ));
 sg13g2_dfrbp_1 _4913_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net121),
    .D(net336),
    .Q_N(_2229_),
    .Q(\configuration[8] ));
 sg13g2_dfrbp_1 _4914_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net119),
    .D(net327),
    .Q_N(_2228_),
    .Q(\configuration[9] ));
 sg13g2_dfrbp_1 _4915_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net117),
    .D(_0169_),
    .Q_N(_2227_),
    .Q(\configuration[10] ));
 sg13g2_dfrbp_1 _4916_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net115),
    .D(_0170_),
    .Q_N(_2226_),
    .Q(\configuration[11] ));
 sg13g2_dfrbp_1 _4917_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net96),
    .D(net232),
    .Q_N(_2225_),
    .Q(\configuration[12] ));
 sg13g2_dfrbp_1 _4918_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net94),
    .D(net325),
    .Q_N(_2224_),
    .Q(\configuration[13] ));
 sg13g2_dfrbp_1 _4919_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net92),
    .D(_0173_),
    .Q_N(_2223_),
    .Q(\configuration[14] ));
 sg13g2_dfrbp_1 _4920_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net90),
    .D(_0174_),
    .Q_N(_2222_),
    .Q(\configuration[15] ));
 sg13g2_dfrbp_1 _4921_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net88),
    .D(_0175_),
    .Q_N(_2221_),
    .Q(\configuration[16] ));
 sg13g2_dfrbp_1 _4922_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net86),
    .D(net399),
    .Q_N(_2220_),
    .Q(\configuration[17] ));
 sg13g2_dfrbp_1 _4923_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net84),
    .D(net299),
    .Q_N(_2219_),
    .Q(\configuration[18] ));
 sg13g2_dfrbp_1 _4924_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net82),
    .D(_0178_),
    .Q_N(_2218_),
    .Q(\configuration[19] ));
 sg13g2_dfrbp_1 _4925_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net80),
    .D(_0179_),
    .Q_N(_2217_),
    .Q(\configuration[20] ));
 sg13g2_dfrbp_1 _4926_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net78),
    .D(net385),
    .Q_N(_2216_),
    .Q(\configuration[21] ));
 sg13g2_dfrbp_1 _4927_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net61),
    .D(net348),
    .Q_N(_2215_),
    .Q(\configuration[22] ));
 sg13g2_dfrbp_1 _4928_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net60),
    .D(_0182_),
    .Q_N(_2214_),
    .Q(\configuration[23] ));
 sg13g2_dfrbp_1 _4929_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net54),
    .D(net343),
    .Q_N(_2213_),
    .Q(\configuration[24] ));
 sg13g2_dfrbp_1 _4930_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net52),
    .D(_0184_),
    .Q_N(_2212_),
    .Q(\configuration[25] ));
 sg13g2_dfrbp_1 _4931_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net50),
    .D(_0185_),
    .Q_N(_2211_),
    .Q(\configuration[26] ));
 sg13g2_dfrbp_1 _4932_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net48),
    .D(net354),
    .Q_N(_2210_),
    .Q(\configuration[27] ));
 sg13g2_dfrbp_1 _4933_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net46),
    .D(_0187_),
    .Q_N(_2209_),
    .Q(\configuration[28] ));
 sg13g2_dfrbp_1 _4934_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net44),
    .D(net341),
    .Q_N(_2208_),
    .Q(\configuration[29] ));
 sg13g2_dfrbp_1 _4935_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net42),
    .D(_0189_),
    .Q_N(_2207_),
    .Q(\configuration[30] ));
 sg13g2_dfrbp_1 _4936_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net40),
    .D(_0190_),
    .Q_N(_2206_),
    .Q(\configuration[31] ));
 sg13g2_dfrbp_1 _4937_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net38),
    .D(_0191_),
    .Q_N(_2205_),
    .Q(\configuration[32] ));
 sg13g2_dfrbp_1 _4938_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net36),
    .D(_0192_),
    .Q_N(_2204_),
    .Q(\configuration[33] ));
 sg13g2_dfrbp_1 _4939_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net34),
    .D(net778),
    .Q_N(_2203_),
    .Q(\configuration[34] ));
 sg13g2_dfrbp_1 _4940_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net32),
    .D(_0194_),
    .Q_N(_2202_),
    .Q(\configuration[35] ));
 sg13g2_dfrbp_1 _4941_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net29),
    .D(net802),
    .Q_N(_2201_),
    .Q(\configuration[36] ));
 sg13g2_dfrbp_1 _4942_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net20),
    .D(_0196_),
    .Q_N(_2200_),
    .Q(\configuration[37] ));
 sg13g2_dfrbp_1 _4943_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net18),
    .D(_0197_),
    .Q_N(_2199_),
    .Q(\configuration[38] ));
 sg13g2_dfrbp_1 _4944_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net16),
    .D(net797),
    .Q_N(_2198_),
    .Q(\configuration[39] ));
 sg13g2_dfrbp_1 _4945_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net14),
    .D(net776),
    .Q_N(_2197_),
    .Q(\configuration[40] ));
 sg13g2_dfrbp_1 _4946_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net12),
    .D(net334),
    .Q_N(_0018_),
    .Q(\configuration[41] ));
 sg13g2_dfrbp_1 _4947_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net185),
    .D(_0201_),
    .Q_N(_2196_),
    .Q(\configuration[42] ));
 sg13g2_dfrbp_1 _4948_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net181),
    .D(_0202_),
    .Q_N(_2195_),
    .Q(\configuration[43] ));
 sg13g2_dfrbp_1 _4949_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net179),
    .D(_0203_),
    .Q_N(_2194_),
    .Q(\configuration[44] ));
 sg13g2_dfrbp_1 _4950_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net177),
    .D(_0204_),
    .Q_N(_2193_),
    .Q(\configuration[45] ));
 sg13g2_dfrbp_1 _4951_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net175),
    .D(net303),
    .Q_N(_2192_),
    .Q(\configuration[46] ));
 sg13g2_dfrbp_1 _4952_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net173),
    .D(_0206_),
    .Q_N(_2191_),
    .Q(\configuration[47] ));
 sg13g2_dfrbp_1 _4953_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net171),
    .D(_0207_),
    .Q_N(_2190_),
    .Q(\configuration[48] ));
 sg13g2_dfrbp_1 _4954_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net169),
    .D(net272),
    .Q_N(_2189_),
    .Q(\configuration[49] ));
 sg13g2_dfrbp_1 _4955_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net167),
    .D(_0209_),
    .Q_N(_2188_),
    .Q(\configuration[50] ));
 sg13g2_dfrbp_1 _4956_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net165),
    .D(_0210_),
    .Q_N(_2187_),
    .Q(\configuration[51] ));
 sg13g2_dfrbp_1 _4957_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net163),
    .D(net270),
    .Q_N(_2186_),
    .Q(\configuration[52] ));
 sg13g2_dfrbp_1 _4958_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net161),
    .D(net743),
    .Q_N(_2185_),
    .Q(\vga.pixel_buffer[0] ));
 sg13g2_dfrbp_1 _4959_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net159),
    .D(net749),
    .Q_N(_2184_),
    .Q(\vga.pixel_buffer[1] ));
 sg13g2_dfrbp_1 _4960_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net157),
    .D(net403),
    .Q_N(_2183_),
    .Q(\vga.pixel_buffer[2] ));
 sg13g2_dfrbp_1 _4961_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net184),
    .D(net407),
    .Q_N(_2384_),
    .Q(\vga.pixel_buffer[3] ));
 sg13g2_dfrbp_1 _4962_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net625),
    .D(_0006_),
    .Q_N(_2385_),
    .Q(\vga.pixel_ctr[0] ));
 sg13g2_dfrbp_1 _4963_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net625),
    .D(net783),
    .Q_N(_2386_),
    .Q(\vga.pixel_ctr[1] ));
 sg13g2_dfrbp_1 _4964_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net623),
    .D(_0009_),
    .Q_N(_0106_),
    .Q(\vga.pixel_ctr[2] ));
 sg13g2_dfrbp_1 _4965_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net625),
    .D(net449),
    .Q_N(_2387_),
    .Q(\vga.pixel_ctr[3] ));
 sg13g2_dfrbp_1 _4966_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net623),
    .D(_0011_),
    .Q_N(_2388_),
    .Q(\vga.pixel_ctr[4] ));
 sg13g2_dfrbp_1 _4967_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net625),
    .D(_0012_),
    .Q_N(_0107_),
    .Q(\vga.pixel_ctr[5] ));
 sg13g2_dfrbp_1 _4968_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net625),
    .D(net496),
    .Q_N(_2389_),
    .Q(\vga.pixel_ctr[6] ));
 sg13g2_dfrbp_1 _4969_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net625),
    .D(_0014_),
    .Q_N(_0108_),
    .Q(\vga.pixel_ctr[7] ));
 sg13g2_dfrbp_1 _4970_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net623),
    .D(_0015_),
    .Q_N(_0109_),
    .Q(\vga.pixel_ctr[8] ));
 sg13g2_dfrbp_1 _4971_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net624),
    .D(_0016_),
    .Q_N(_2390_),
    .Q(\vga.pixel_ctr[9] ));
 sg13g2_dfrbp_1 _4972_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net623),
    .D(net222),
    .Q_N(_0110_),
    .Q(\vga.pixel_ctr[10] ));
 sg13g2_dfrbp_1 _4973_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net153),
    .D(valid_data),
    .Q_N(_2391_),
    .Q(\vga.wrote_data ));
 sg13g2_dfrbp_1 _4974_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net155),
    .D(net786),
    .Q_N(_2182_),
    .Q(\vga.l_read ));
 sg13g2_dfrbp_1 _4975_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net630),
    .D(net780),
    .Q_N(_0017_),
    .Q(\mandelbrot.alu.m1[31] ));
 sg13g2_tiehi _4670__11 (.L_HI(net11));
 sg13g2_tiehi _4946__12 (.L_HI(net12));
 sg13g2_tiehi _4853__13 (.L_HI(net13));
 sg13g2_tiehi _4945__14 (.L_HI(net14));
 sg13g2_tiehi _4852__15 (.L_HI(net15));
 sg13g2_tiehi _4944__16 (.L_HI(net16));
 sg13g2_tiehi _4851__17 (.L_HI(net17));
 sg13g2_tiehi _4943__18 (.L_HI(net18));
 sg13g2_tiehi _4850__19 (.L_HI(net19));
 sg13g2_tiehi _4942__20 (.L_HI(net20));
 sg13g2_tiehi _4849__21 (.L_HI(net21));
 sg13g2_tiehi _4681__22 (.L_HI(net22));
 sg13g2_tiehi _4682__23 (.L_HI(net23));
 sg13g2_tiehi _4683__24 (.L_HI(net24));
 sg13g2_tiehi _4684__25 (.L_HI(net25));
 sg13g2_tiehi _4685__26 (.L_HI(net26));
 sg13g2_tiehi _4686__27 (.L_HI(net27));
 sg13g2_tiehi _4687__28 (.L_HI(net28));
 sg13g2_tiehi _4941__29 (.L_HI(net29));
 sg13g2_tiehi _4848__30 (.L_HI(net30));
 sg13g2_tiehi _4688__31 (.L_HI(net31));
 sg13g2_tiehi _4940__32 (.L_HI(net32));
 sg13g2_tiehi _4847__33 (.L_HI(net33));
 sg13g2_tiehi _4939__34 (.L_HI(net34));
 sg13g2_tiehi _4846__35 (.L_HI(net35));
 sg13g2_tiehi _4938__36 (.L_HI(net36));
 sg13g2_tiehi _4845__37 (.L_HI(net37));
 sg13g2_tiehi _4937__38 (.L_HI(net38));
 sg13g2_tiehi _4844__39 (.L_HI(net39));
 sg13g2_tiehi _4936__40 (.L_HI(net40));
 sg13g2_tiehi _4843__41 (.L_HI(net41));
 sg13g2_tiehi _4935__42 (.L_HI(net42));
 sg13g2_tiehi _4842__43 (.L_HI(net43));
 sg13g2_tiehi _4934__44 (.L_HI(net44));
 sg13g2_tiehi _4841__45 (.L_HI(net45));
 sg13g2_tiehi _4933__46 (.L_HI(net46));
 sg13g2_tiehi _4840__47 (.L_HI(net47));
 sg13g2_tiehi _4932__48 (.L_HI(net48));
 sg13g2_tiehi _4839__49 (.L_HI(net49));
 sg13g2_tiehi _4931__50 (.L_HI(net50));
 sg13g2_tiehi _4838__51 (.L_HI(net51));
 sg13g2_tiehi _4930__52 (.L_HI(net52));
 sg13g2_tiehi _4837__53 (.L_HI(net53));
 sg13g2_tiehi _4929__54 (.L_HI(net54));
 sg13g2_tiehi _4836__55 (.L_HI(net55));
 sg13g2_tiehi _4835__56 (.L_HI(net56));
 sg13g2_tiehi _4834__57 (.L_HI(net57));
 sg13g2_tiehi _4833__58 (.L_HI(net58));
 sg13g2_tiehi _4832__59 (.L_HI(net59));
 sg13g2_tiehi _4928__60 (.L_HI(net60));
 sg13g2_tiehi _4927__61 (.L_HI(net61));
 sg13g2_tiehi _4830__62 (.L_HI(net62));
 sg13g2_tiehi _4829__63 (.L_HI(net63));
 sg13g2_tiehi _4828__64 (.L_HI(net64));
 sg13g2_tiehi _4827__65 (.L_HI(net65));
 sg13g2_tiehi _4826__66 (.L_HI(net66));
 sg13g2_tiehi _4825__67 (.L_HI(net67));
 sg13g2_tiehi _4824__68 (.L_HI(net68));
 sg13g2_tiehi _4823__69 (.L_HI(net69));
 sg13g2_tiehi _4822__70 (.L_HI(net70));
 sg13g2_tiehi _4821__71 (.L_HI(net71));
 sg13g2_tiehi _4820__72 (.L_HI(net72));
 sg13g2_tiehi _4819__73 (.L_HI(net73));
 sg13g2_tiehi _4818__74 (.L_HI(net74));
 sg13g2_tiehi _4817__75 (.L_HI(net75));
 sg13g2_tiehi _4816__76 (.L_HI(net76));
 sg13g2_tiehi _4815__77 (.L_HI(net77));
 sg13g2_tiehi _4926__78 (.L_HI(net78));
 sg13g2_tiehi _4814__79 (.L_HI(net79));
 sg13g2_tiehi _4925__80 (.L_HI(net80));
 sg13g2_tiehi _4813__81 (.L_HI(net81));
 sg13g2_tiehi _4924__82 (.L_HI(net82));
 sg13g2_tiehi _4812__83 (.L_HI(net83));
 sg13g2_tiehi _4923__84 (.L_HI(net84));
 sg13g2_tiehi _4811__85 (.L_HI(net85));
 sg13g2_tiehi _4922__86 (.L_HI(net86));
 sg13g2_tiehi _4810__87 (.L_HI(net87));
 sg13g2_tiehi _4921__88 (.L_HI(net88));
 sg13g2_tiehi _4809__89 (.L_HI(net89));
 sg13g2_tiehi _4920__90 (.L_HI(net90));
 sg13g2_tiehi _4808__91 (.L_HI(net91));
 sg13g2_tiehi _4919__92 (.L_HI(net92));
 sg13g2_tiehi _4807__93 (.L_HI(net93));
 sg13g2_tiehi _4918__94 (.L_HI(net94));
 sg13g2_tiehi _4806__95 (.L_HI(net95));
 sg13g2_tiehi _4917__96 (.L_HI(net96));
 sg13g2_tiehi _4805__97 (.L_HI(net97));
 sg13g2_tiehi _4804__98 (.L_HI(net98));
 sg13g2_tiehi _4803__99 (.L_HI(net99));
 sg13g2_tiehi _4802__100 (.L_HI(net100));
 sg13g2_tiehi _4801__101 (.L_HI(net101));
 sg13g2_tiehi _4800__102 (.L_HI(net102));
 sg13g2_tiehi _4799__103 (.L_HI(net103));
 sg13g2_tiehi _4798__104 (.L_HI(net104));
 sg13g2_tiehi _4768__105 (.L_HI(net105));
 sg13g2_tiehi _4797__106 (.L_HI(net106));
 sg13g2_tiehi _4796__107 (.L_HI(net107));
 sg13g2_tiehi _4795__108 (.L_HI(net108));
 sg13g2_tiehi _4794__109 (.L_HI(net109));
 sg13g2_tiehi _4793__110 (.L_HI(net110));
 sg13g2_tiehi _4792__111 (.L_HI(net111));
 sg13g2_tiehi _4791__112 (.L_HI(net112));
 sg13g2_tiehi _4790__113 (.L_HI(net113));
 sg13g2_tiehi _4789__114 (.L_HI(net114));
 sg13g2_tiehi _4916__115 (.L_HI(net115));
 sg13g2_tiehi _4788__116 (.L_HI(net116));
 sg13g2_tiehi _4915__117 (.L_HI(net117));
 sg13g2_tiehi _4787__118 (.L_HI(net118));
 sg13g2_tiehi _4914__119 (.L_HI(net119));
 sg13g2_tiehi _4786__120 (.L_HI(net120));
 sg13g2_tiehi _4913__121 (.L_HI(net121));
 sg13g2_tiehi _4785__122 (.L_HI(net122));
 sg13g2_tiehi _4912__123 (.L_HI(net123));
 sg13g2_tiehi _4784__124 (.L_HI(net124));
 sg13g2_tiehi _4911__125 (.L_HI(net125));
 sg13g2_tiehi _4783__126 (.L_HI(net126));
 sg13g2_tiehi _4910__127 (.L_HI(net127));
 sg13g2_tiehi _4782__128 (.L_HI(net128));
 sg13g2_tiehi _4909__129 (.L_HI(net129));
 sg13g2_tiehi _4781__130 (.L_HI(net130));
 sg13g2_tiehi _4908__131 (.L_HI(net131));
 sg13g2_tiehi _4780__132 (.L_HI(net132));
 sg13g2_tiehi _4907__133 (.L_HI(net133));
 sg13g2_tiehi _4779__134 (.L_HI(net134));
 sg13g2_tiehi _4906__135 (.L_HI(net135));
 sg13g2_tiehi _4778__136 (.L_HI(net136));
 sg13g2_tiehi _4905__137 (.L_HI(net137));
 sg13g2_tiehi _4777__138 (.L_HI(net138));
 sg13g2_tiehi _4776__139 (.L_HI(net139));
 sg13g2_tiehi _4775__140 (.L_HI(net140));
 sg13g2_tiehi _4774__141 (.L_HI(net141));
 sg13g2_tiehi _4773__142 (.L_HI(net142));
 sg13g2_tiehi _4767__143 (.L_HI(net143));
 sg13g2_tiehi _4766__144 (.L_HI(net144));
 sg13g2_tiehi _4732__145 (.L_HI(net145));
 sg13g2_tiehi _4731__146 (.L_HI(net146));
 sg13g2_tiehi _4730__147 (.L_HI(net147));
 sg13g2_tiehi _4729__148 (.L_HI(net148));
 sg13g2_tiehi _4728__149 (.L_HI(net149));
 sg13g2_tiehi _4727__150 (.L_HI(net150));
 sg13g2_tiehi _4690__151 (.L_HI(net151));
 sg13g2_tiehi _4689__152 (.L_HI(net152));
 sg13g2_tiehi _4973__153 (.L_HI(net153));
 sg13g2_tiehi _4869__154 (.L_HI(net154));
 sg13g2_tiehi _4974__155 (.L_HI(net155));
 sg13g2_tiehi _4868__156 (.L_HI(net156));
 sg13g2_tiehi _4960__157 (.L_HI(net157));
 sg13g2_tiehi _4867__158 (.L_HI(net158));
 sg13g2_tiehi _4959__159 (.L_HI(net159));
 sg13g2_tiehi _4866__160 (.L_HI(net160));
 sg13g2_tiehi _4958__161 (.L_HI(net161));
 sg13g2_tiehi _4865__162 (.L_HI(net162));
 sg13g2_tiehi _4957__163 (.L_HI(net163));
 sg13g2_tiehi _4864__164 (.L_HI(net164));
 sg13g2_tiehi _4956__165 (.L_HI(net165));
 sg13g2_tiehi _4863__166 (.L_HI(net166));
 sg13g2_tiehi _4955__167 (.L_HI(net167));
 sg13g2_tiehi _4862__168 (.L_HI(net168));
 sg13g2_tiehi _4954__169 (.L_HI(net169));
 sg13g2_tiehi _4861__170 (.L_HI(net170));
 sg13g2_tiehi _4953__171 (.L_HI(net171));
 sg13g2_tiehi _4860__172 (.L_HI(net172));
 sg13g2_tiehi _4952__173 (.L_HI(net173));
 sg13g2_tiehi _4859__174 (.L_HI(net174));
 sg13g2_tiehi _4951__175 (.L_HI(net175));
 sg13g2_tiehi _4858__176 (.L_HI(net176));
 sg13g2_tiehi _4950__177 (.L_HI(net177));
 sg13g2_tiehi _4857__178 (.L_HI(net178));
 sg13g2_tiehi _4949__179 (.L_HI(net179));
 sg13g2_tiehi _4856__180 (.L_HI(net180));
 sg13g2_tiehi _4948__181 (.L_HI(net181));
 sg13g2_tiehi _4855__182 (.L_HI(net182));
 sg13g2_tiehi _4870__183 (.L_HI(net183));
 sg13g2_tiehi _4961__184 (.L_HI(net184));
 sg13g2_tiehi _4947__185 (.L_HI(net185));
 sg13g2_tiehi tt_um_gfg_development_tinymandelbrot_186 (.L_HI(net186));
 sg13g2_tiehi tt_um_gfg_development_tinymandelbrot_187 (.L_HI(net187));
 sg13g2_tiehi tt_um_gfg_development_tinymandelbrot_188 (.L_HI(net188));
 sg13g2_tiehi tt_um_gfg_development_tinymandelbrot_189 (.L_HI(net189));
 sg13g2_tiehi tt_um_gfg_development_tinymandelbrot_190 (.L_HI(net190));
 sg13g2_tiehi tt_um_gfg_development_tinymandelbrot_191 (.L_HI(net191));
 sg13g2_tiehi tt_um_gfg_development_tinymandelbrot_192 (.L_HI(net192));
 sg13g2_tiehi tt_um_gfg_development_tinymandelbrot_193 (.L_HI(net193));
 sg13g2_inv_1 _2642__1 (.Y(net194),
    .A(clknet_1_0__leaf_clk));
 sg13g2_buf_1 _5160_ (.A(reset_write_ptr),
    .X(uio_out[4]));
 sg13g2_buf_1 _5161_ (.A(valid_data),
    .X(uio_out[5]));
 sg13g2_buf_2 _5162_ (.A(\vga.reset_read_ptr ),
    .X(uio_out[6]));
 sg13g2_buf_1 _5163_ (.A(\vga.read ),
    .X(uio_out[7]));
 sg13g2_buf_2 fanout536 (.A(_1302_),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(net538),
    .X(net537));
 sg13g2_buf_1 fanout538 (.A(net539),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(net543),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(net543),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(net543),
    .X(net541));
 sg13g2_buf_1 fanout542 (.A(net543),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(_1301_),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(net545),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(net546),
    .X(net545));
 sg13g2_buf_4 fanout546 (.X(net546),
    .A(net549));
 sg13g2_buf_2 fanout547 (.A(net548),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(net549),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(_0837_),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(net551),
    .X(net550));
 sg13g2_buf_1 fanout551 (.A(net552),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(_0832_),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(net554),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(net555),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(_0832_),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(net557),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(_0508_),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(net559),
    .X(net558));
 sg13g2_buf_1 fanout559 (.A(net560),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(_0505_),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(net563),
    .X(net561));
 sg13g2_buf_4 fanout562 (.X(net562),
    .A(net563));
 sg13g2_buf_2 fanout563 (.A(_0505_),
    .X(net563));
 sg13g2_buf_4 fanout564 (.X(net564),
    .A(_0437_));
 sg13g2_buf_4 fanout565 (.X(net565),
    .A(_0436_));
 sg13g2_buf_4 fanout566 (.X(net566),
    .A(_0428_));
 sg13g2_buf_4 fanout567 (.X(net567),
    .A(_0427_));
 sg13g2_buf_2 fanout568 (.A(net569),
    .X(net568));
 sg13g2_buf_1 fanout569 (.A(net570),
    .X(net569));
 sg13g2_buf_1 fanout570 (.A(_1294_),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(_1294_),
    .X(net571));
 sg13g2_buf_1 fanout572 (.A(net573),
    .X(net572));
 sg13g2_buf_4 fanout573 (.X(net573),
    .A(_1294_));
 sg13g2_buf_4 fanout574 (.X(net574),
    .A(net576));
 sg13g2_buf_2 fanout575 (.A(net576),
    .X(net575));
 sg13g2_buf_4 fanout576 (.X(net576),
    .A(_1278_));
 sg13g2_buf_4 fanout577 (.X(net577),
    .A(net578));
 sg13g2_buf_4 fanout578 (.X(net578),
    .A(net579));
 sg13g2_buf_4 fanout579 (.X(net579),
    .A(_1278_));
 sg13g2_buf_4 fanout580 (.X(net580),
    .A(_0426_));
 sg13g2_buf_4 fanout581 (.X(net581),
    .A(_0447_));
 sg13g2_buf_2 fanout582 (.A(_0447_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_2181_),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(_2180_),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(net587),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(net587),
    .X(net586));
 sg13g2_buf_4 fanout587 (.X(net587),
    .A(_1275_));
 sg13g2_buf_4 fanout588 (.X(net588),
    .A(net589));
 sg13g2_buf_2 fanout589 (.A(net590),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(_1275_),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(_1275_),
    .X(net591));
 sg13g2_buf_4 fanout592 (.X(net592),
    .A(_1683_));
 sg13g2_buf_4 fanout593 (.X(net593),
    .A(_1683_));
 sg13g2_buf_2 fanout594 (.A(_1682_),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(_1682_),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(net597),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(_1299_),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(net599),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(_1299_),
    .X(net599));
 sg13g2_buf_4 fanout600 (.X(net600),
    .A(_1069_));
 sg13g2_buf_2 fanout601 (.A(net602),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(net603),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(_1068_),
    .X(net603));
 sg13g2_buf_4 fanout604 (.X(net604),
    .A(_0611_));
 sg13g2_buf_1 fanout605 (.A(_0611_),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(net607),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(net608),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(_0610_),
    .X(net608));
 sg13g2_buf_4 fanout609 (.X(net609),
    .A(net613));
 sg13g2_buf_4 fanout610 (.X(net610),
    .A(net613));
 sg13g2_buf_4 fanout611 (.X(net611),
    .A(net613));
 sg13g2_buf_2 fanout612 (.A(net613),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(net632),
    .X(net613));
 sg13g2_buf_4 fanout614 (.X(net614),
    .A(net615));
 sg13g2_buf_4 fanout615 (.X(net615),
    .A(net616));
 sg13g2_buf_4 fanout616 (.X(net616),
    .A(net622));
 sg13g2_buf_4 fanout617 (.X(net617),
    .A(net619));
 sg13g2_buf_4 fanout618 (.X(net618),
    .A(net619));
 sg13g2_buf_2 fanout619 (.A(net622),
    .X(net619));
 sg13g2_buf_4 fanout620 (.X(net620),
    .A(net621));
 sg13g2_buf_4 fanout621 (.X(net621),
    .A(net622));
 sg13g2_buf_2 fanout622 (.A(net632),
    .X(net622));
 sg13g2_buf_4 fanout623 (.X(net623),
    .A(net625));
 sg13g2_buf_4 fanout624 (.X(net624),
    .A(net625));
 sg13g2_buf_4 fanout625 (.X(net625),
    .A(net626));
 sg13g2_buf_4 fanout626 (.X(net626),
    .A(net627));
 sg13g2_buf_2 fanout627 (.A(net632),
    .X(net627));
 sg13g2_buf_4 fanout628 (.X(net628),
    .A(net631));
 sg13g2_buf_4 fanout629 (.X(net629),
    .A(net631));
 sg13g2_buf_4 fanout630 (.X(net630),
    .A(net631));
 sg13g2_buf_4 fanout631 (.X(net631),
    .A(net632));
 sg13g2_buf_2 fanout632 (.A(combined_rst_n),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(_1680_),
    .X(net633));
 sg13g2_buf_4 fanout634 (.X(net634),
    .A(_1680_));
 sg13g2_buf_2 fanout635 (.A(_1679_),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(net637),
    .X(net636));
 sg13g2_buf_1 fanout637 (.A(net638),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(net639),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(net640),
    .X(net639));
 sg13g2_buf_4 fanout640 (.X(net640),
    .A(_1065_));
 sg13g2_buf_2 fanout641 (.A(net643),
    .X(net641));
 sg13g2_buf_1 fanout642 (.A(net643),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(_0608_),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(_0608_),
    .X(net644));
 sg13g2_buf_4 fanout645 (.X(net645),
    .A(net648));
 sg13g2_buf_4 fanout646 (.X(net646),
    .A(net648));
 sg13g2_buf_2 fanout647 (.A(net648),
    .X(net647));
 sg13g2_buf_4 fanout648 (.X(net648),
    .A(_1891_));
 sg13g2_buf_2 fanout649 (.A(net650),
    .X(net649));
 sg13g2_buf_4 fanout650 (.X(net650),
    .A(net651));
 sg13g2_buf_2 fanout651 (.A(_1891_),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(net654),
    .X(net652));
 sg13g2_buf_4 fanout653 (.X(net653),
    .A(net654));
 sg13g2_buf_2 fanout654 (.A(_1891_),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(net656),
    .X(net655));
 sg13g2_buf_4 fanout656 (.X(net656),
    .A(_1912_));
 sg13g2_buf_2 fanout657 (.A(net658),
    .X(net657));
 sg13g2_buf_4 fanout658 (.X(net658),
    .A(_1911_));
 sg13g2_buf_2 fanout659 (.A(net661),
    .X(net659));
 sg13g2_buf_1 fanout660 (.A(net661),
    .X(net660));
 sg13g2_buf_4 fanout661 (.X(net661),
    .A(net663));
 sg13g2_buf_4 fanout662 (.X(net662),
    .A(net663));
 sg13g2_buf_2 fanout663 (.A(\mandelbrot.running ),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(net269),
    .X(net664));
 sg13g2_buf_4 fanout665 (.X(net665),
    .A(net667));
 sg13g2_buf_1 fanout666 (.A(net667),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(\mandelbrot.alu.m1[1] ),
    .X(net667));
 sg13g2_buf_2 fanout668 (.A(net670),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(net670),
    .X(net669));
 sg13g2_buf_2 fanout670 (.A(\mandelbrot.alu.m1[1] ),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(net811),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(\mandelbrot.ctr[5] ),
    .X(net672));
 sg13g2_buf_4 fanout673 (.X(net673),
    .A(net728));
 sg13g2_buf_2 fanout674 (.A(net675),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(net676),
    .X(net675));
 sg13g2_buf_4 fanout676 (.X(net676),
    .A(net679));
 sg13g2_buf_4 fanout677 (.X(net677),
    .A(net679));
 sg13g2_buf_4 fanout678 (.X(net678),
    .A(net679));
 sg13g2_buf_4 fanout679 (.X(net679),
    .A(net522));
 sg13g2_buf_2 fanout680 (.A(net683),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(net683),
    .X(net681));
 sg13g2_buf_4 fanout682 (.X(net682),
    .A(net683));
 sg13g2_buf_4 fanout683 (.X(net683),
    .A(net511));
 sg13g2_buf_4 fanout684 (.X(net684),
    .A(net685));
 sg13g2_buf_2 fanout685 (.A(\mandelbrot.alu.mult_zi_zi.running ),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(net687),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(net688),
    .X(net687));
 sg13g2_buf_4 fanout688 (.X(net688),
    .A(\mandelbrot.alu.mult_zi_zi.running ));
 sg13g2_buf_4 fanout689 (.X(net689),
    .A(net693));
 sg13g2_buf_2 fanout690 (.A(net693),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(net692),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(net693),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(\mandelbrot.alu.mult_zr_zr.running ),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(net695),
    .X(net694));
 sg13g2_buf_1 fanout695 (.A(net696),
    .X(net695));
 sg13g2_buf_1 fanout696 (.A(net697),
    .X(net696));
 sg13g2_buf_1 fanout697 (.A(net699),
    .X(net697));
 sg13g2_buf_2 fanout698 (.A(net699),
    .X(net698));
 sg13g2_buf_4 fanout699 (.X(net699),
    .A(\mandelbrot.alu.m3[1] ));
 sg13g2_buf_4 fanout700 (.X(net700),
    .A(\mandelbrot.alu.m2[25] ));
 sg13g2_buf_2 fanout701 (.A(net703),
    .X(net701));
 sg13g2_buf_2 fanout702 (.A(net703),
    .X(net702));
 sg13g2_buf_4 fanout703 (.X(net703),
    .A(\mandelbrot.alu.m2[1] ));
 sg13g2_buf_2 fanout704 (.A(net705),
    .X(net704));
 sg13g2_buf_1 fanout705 (.A(net787),
    .X(net705));
 sg13g2_buf_4 fanout706 (.X(net706),
    .A(\mandelbrot.alu.m2[1] ));
 sg13g2_buf_4 fanout707 (.X(net707),
    .A(net5));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_tiehi _4854__10 (.L_HI(net10));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(delaynet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_leaf_0_clk_regs (.A(clknet_3_1__leaf_clk_regs),
    .X(clknet_leaf_0_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_1_clk_regs (.A(clknet_3_1__leaf_clk_regs),
    .X(clknet_leaf_1_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_2_clk_regs (.A(clknet_3_1__leaf_clk_regs),
    .X(clknet_leaf_2_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_3_clk_regs (.A(clknet_3_1__leaf_clk_regs),
    .X(clknet_leaf_3_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_4_clk_regs (.A(clknet_3_1__leaf_clk_regs),
    .X(clknet_leaf_4_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_5_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_5_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_6_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_6_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_7_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_7_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_8_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_8_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_9_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_9_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_10_clk_regs (.A(clknet_3_5__leaf_clk_regs),
    .X(clknet_leaf_10_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_11_clk_regs (.A(clknet_3_5__leaf_clk_regs),
    .X(clknet_leaf_11_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_12_clk_regs (.A(clknet_3_5__leaf_clk_regs),
    .X(clknet_leaf_12_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_13_clk_regs (.A(clknet_3_5__leaf_clk_regs),
    .X(clknet_leaf_13_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_14_clk_regs (.A(clknet_3_5__leaf_clk_regs),
    .X(clknet_leaf_14_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_15_clk_regs (.A(clknet_3_7__leaf_clk_regs),
    .X(clknet_leaf_15_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_16_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_16_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_17_clk_regs (.A(clknet_3_6__leaf_clk_regs),
    .X(clknet_leaf_17_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_18_clk_regs (.A(clknet_3_6__leaf_clk_regs),
    .X(clknet_leaf_18_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_19_clk_regs (.A(clknet_3_6__leaf_clk_regs),
    .X(clknet_leaf_19_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_20_clk_regs (.A(clknet_3_7__leaf_clk_regs),
    .X(clknet_leaf_20_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_21_clk_regs (.A(clknet_3_7__leaf_clk_regs),
    .X(clknet_leaf_21_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_22_clk_regs (.A(clknet_3_7__leaf_clk_regs),
    .X(clknet_leaf_22_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_23_clk_regs (.A(clknet_3_7__leaf_clk_regs),
    .X(clknet_leaf_23_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_24_clk_regs (.A(clknet_3_6__leaf_clk_regs),
    .X(clknet_leaf_24_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_25_clk_regs (.A(clknet_3_6__leaf_clk_regs),
    .X(clknet_leaf_25_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_26_clk_regs (.A(clknet_3_3__leaf_clk_regs),
    .X(clknet_leaf_26_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_27_clk_regs (.A(clknet_3_3__leaf_clk_regs),
    .X(clknet_leaf_27_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_28_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_28_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_29_clk_regs (.A(clknet_3_3__leaf_clk_regs),
    .X(clknet_leaf_29_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_30_clk_regs (.A(clknet_3_3__leaf_clk_regs),
    .X(clknet_leaf_30_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_31_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_31_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_32_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_32_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_33_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_33_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_34_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_34_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_35_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_35_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_36_clk_regs (.A(clknet_3_3__leaf_clk_regs),
    .X(clknet_leaf_36_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_37_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_37_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_38_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_38_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_39_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_39_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_40_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_40_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_41_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_41_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_42_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_42_clk_regs));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_3_0__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_1__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_1__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_2__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_2__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_3__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_3__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_4__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_4__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_5__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_5__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_6__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_6__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_7__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_7__leaf_clk_regs));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk_regs));
 sg13g2_buf_2 clkload1 (.A(clknet_3_3__leaf_clk_regs));
 sg13g2_buf_2 clkload2 (.A(clknet_3_5__leaf_clk_regs));
 sg13g2_buf_2 clkload3 (.A(clknet_3_6__leaf_clk_regs));
 sg13g2_buf_2 clkload4 (.A(clknet_3_7__leaf_clk_regs));
 sg13g2_inv_4 clkload5 (.A(clknet_leaf_39_clk_regs));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_40_clk_regs));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_0_clk_regs));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_28_clk_regs));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_31_clk_regs));
 sg13g2_inv_2 clkload10 (.A(clknet_leaf_32_clk_regs));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_33_clk_regs));
 sg13g2_inv_4 clkload12 (.A(clknet_leaf_34_clk_regs));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_27_clk_regs));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_30_clk_regs));
 sg13g2_inv_1 clkload15 (.A(clknet_leaf_36_clk_regs));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_18_clk_regs));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_24_clk_regs));
 sg13g2_inv_2 clkload18 (.A(clknet_leaf_21_clk_regs));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_23_clk_regs));
 sg13g2_buf_2 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(delaynet_1_clk));
 sg13g2_buf_2 delaybuf_1_clk (.A(delaynet_1_clk),
    .X(clknet_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\l_sclk[1] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold2 (.A(\l_sdata[1] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold3 (.A(\l_sclk[0] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold4 (.A(\l_sen[0] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0102_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold6 (.A(\l_sdata[0] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold7 (.A(\state[2] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold8 (.A(\l_sen[1] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold9 (.A(\mandelbrot.alu.finished ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold10 (.A(\state[0] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0000_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0089_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0259_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold14 (.A(finished),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0115_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0088_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0262_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0048_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0365_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0077_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold21 (.A(_1266_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0297_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0057_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0333_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0031_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0117_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0110_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0007_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0113_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold30 (.A(_1509_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold31 (.A(\mandelbrot.alu.in_cr[7] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0350_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold33 (.A(\mandelbrot.alu.mult_zr_zi.ctr[1] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0835_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0260_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold36 (.A(\mandelbrot.ctr[5] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold37 (.A(\configuration[12] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0171_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold39 (.A(\mandelbrot.alu.m3[2] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0266_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold41 (.A(\mandelbrot.alu.mult_zi_zi.ctr[1] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold42 (.A(_1267_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0298_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0106_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0449_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold46 (.A(\mandelbrot.alu.mult_zr_zr.ctr[1] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0840_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0263_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold49 (.A(\mandelbrot.alu.m3[5] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0269_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0086_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold52 (.A(_1112_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold53 (.A(\configuration[2] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0161_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold55 (.A(\mandelbrot.x[1] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold56 (.A(_1599_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0366_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold58 (.A(\mandelbrot.overflowed ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold59 (.A(\mandelbrot.alu.mult_zr_zr.ctr[2] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0264_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold61 (.A(\mandelbrot.alu.m3[4] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold62 (.A(\mandelbrot.y[4] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0121_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold64 (.A(\mandelbrot.alu.in_zr[10] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold65 (.A(\mandelbrot.alu.in_zr[15] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold66 (.A(\mandelbrot.alu.in_zr[14] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold67 (.A(\mandelbrot.alu.mult_zr_zi.ctr[2] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0261_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold69 (.A(\mandelbrot.alu.in_zi[7] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold70 (.A(\mandelbrot.x[3] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold71 (.A(_1601_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0368_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0076_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0249_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold75 (.A(\configuration[52] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0211_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold77 (.A(\configuration[50] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0208_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0028_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold80 (.A(_1726_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold81 (.A(l_running),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold82 (.A(\mandelbrot.alu.in_zi[3] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold83 (.A(\mandelbrot.alu.mult_zi_zi.ctr[2] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0299_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold85 (.A(\mandelbrot.alu.in_zr[6] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0099_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0659_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold88 (.A(\state[3] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0002_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold90 (.A(\mandelbrot.y[8] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0125_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold92 (.A(\configuration[51] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold93 (.A(\vga.timing_v.pixel[0] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0217_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold95 (.A(\mandelbrot.alu.in_zi[15] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0085_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold97 (.A(_1122_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold98 (.A(\vga.wrote_data ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold99 (.A(_2568_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold100 (.A(\mandelbrot.alu.in_zr[13] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold101 (.A(\mandelbrot.alu.in_zi[10] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold102 (.A(\mandelbrot.alu.in_zr[7] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold103 (.A(\mandelbrot.alu.in_zr[9] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold104 (.A(\configuration[19] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0177_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold106 (.A(\mandelbrot.alu.m3[11] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0275_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold108 (.A(\configuration[47] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0205_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold110 (.A(\mandelbrot.alu.in_zi[12] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold111 (.A(\mandelbrot.x[6] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold112 (.A(_1607_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0371_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold114 (.A(\configuration[1] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0344_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold116 (.A(\configuration[11] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold117 (.A(\vga.timing_v.pixel[9] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0226_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold119 (.A(\state[1] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold120 (.A(\mandelbrot.alu.in_zi[14] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold121 (.A(\configuration[3] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0162_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0024_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold124 (.A(_1790_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0109_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0457_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold127 (.A(\configuration[7] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0165_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold129 (.A(\mandelbrot.alu.in_zi[2] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold130 (.A(\configuration[14] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0172_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold132 (.A(\configuration[10] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0168_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold134 (.A(\mandelbrot.alu.in_zi[13] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0078_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0293_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold137 (.A(\mandelbrot.alu.in_zr[3] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold138 (.A(\mandelbrot.alu.in_zi[6] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold139 (.A(\configuration[42] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0200_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold141 (.A(\configuration[9] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0167_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold143 (.A(\mandelbrot.alu.in_zi[9] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold144 (.A(\mandelbrot.alu.m3[8] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0274_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold146 (.A(\configuration[30] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0188_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold148 (.A(\configuration[25] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0183_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold150 (.A(\configuration[15] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold151 (.A(\mandelbrot.alu.m3[7] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0962_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold153 (.A(\configuration[23] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0181_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold155 (.A(\configuration[5] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0163_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold157 (.A(\vga.timing_v.pixel[4] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0490_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold159 (.A(\configuration[28] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0186_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold161 (.A(\configuration[29] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold162 (.A(\vga.timing_v.pixel[7] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0224_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold164 (.A(\mandelbrot.alu.in_zi[5] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0021_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold166 (.A(_1843_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold167 (.A(\vga.timing_v.pixel[1] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0218_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold169 (.A(\mandelbrot.alu.in_cr[5] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0092_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold171 (.A(\configuration[20] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0022_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0152_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold174 (.A(\configuration[26] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold175 (.A(\mandelbrot.alu.m3[12] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0278_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold177 (.A(\mandelbrot.alu.m3[13] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold178 (.A(\mandelbrot.alu.in_ci[7] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0324_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold180 (.A(\mandelbrot.alu.in_zr[2] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold181 (.A(\configuration[24] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold182 (.A(\configuration[0] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold183 (.A(\mandelbrot.alu.in_ci[9] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0100_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0645_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold186 (.A(\mandelbrot.alu.m3[15] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold187 (.A(\mandelbrot.alu.in_zr[12] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0313_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold189 (.A(\configuration[16] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold190 (.A(\configuration[22] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0180_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0079_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0292_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold194 (.A(\mandelbrot.alu.in_zr[11] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold195 (.A(\configuration[21] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold196 (.A(\configuration[6] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold197 (.A(\mandelbrot.x[8] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold198 (.A(_1611_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold199 (.A(\configuration[31] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold200 (.A(\mandelbrot.alu.in_cr[14] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold201 (.A(\configuration[27] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold202 (.A(\vga.timing_v.pixel[5] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold203 (.A(\configuration[8] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold204 (.A(\configuration[18] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0176_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold206 (.A(\mandelbrot.alu.mult_zr_zi.shift_reg[0] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0842_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold208 (.A(\vga.pixel_buffer[2] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0214_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0087_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0282_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold212 (.A(\vga.pixel_buffer[3] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0215_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold214 (.A(\vga.timing_v.pixel[8] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0091_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold216 (.A(\mandelbrot.y[2] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0119_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold218 (.A(\mandelbrot.alu.mult_zi_zi.shift_reg[0] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0080_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0290_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0082_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0288_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold223 (.A(\mandelbrot.alu.m3[10] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold224 (.A(\mandelbrot.y[6] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0123_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold226 (.A(\configuration[43] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold227 (.A(\mandelbrot.alu.m3[31] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold228 (.A(\mandelbrot.alu.in_zi[1] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0375_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold230 (.A(\configuration[17] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0104_),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold232 (.A(_1243_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold233 (.A(\mandelbrot.alu.in_zr[8] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold234 (.A(\mandelbrot.y[1] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold235 (.A(_1632_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0118_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold237 (.A(\mandelbrot.alu.in_zi[11] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold238 (.A(\mandelbrot.x[2] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold239 (.A(_1600_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0367_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold241 (.A(\mandelbrot.alu.m3[20] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold242 (.A(_1145_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold243 (.A(\configuration[48] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold244 (.A(\configuration[44] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold245 (.A(\mandelbrot.y[3] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0095_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0723_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold248 (.A(\mandelbrot.alu.in_cr[8] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0351_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0108_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0455_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0090_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold253 (.A(\vga.pixel_ctr[3] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0450_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0010_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold256 (.A(\mandelbrot.alu.in_cr[9] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0029_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold258 (.A(_1710_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold259 (.A(\mandelbrot.alu.in_ci[11] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold260 (.A(\mandelbrot.x[5] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold261 (.A(_0370_),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold262 (.A(\mandelbrot.alu.in_ci[3] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold263 (.A(\configuration[49] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold264 (.A(\mandelbrot.x[4] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold265 (.A(_1604_),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold266 (.A(\mandelbrot.alu.in_cr[3] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold267 (.A(\mandelbrot.alu.m1[21] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0149_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0093_),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0252_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold271 (.A(\mandelbrot.alu.in_cr[10] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold272 (.A(_0353_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0025_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold274 (.A(_1764_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold275 (.A(\mandelbrot.alu.in_zi[4] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold276 (.A(\mandelbrot.alu.m1[11] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0137_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0026_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold279 (.A(_1751_),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold280 (.A(\mandelbrot.alu.m3[25] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0291_),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold282 (.A(\mandelbrot.alu.m1[25] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold283 (.A(\mandelbrot.x[7] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold284 (.A(_0027_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold285 (.A(_1737_),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold286 (.A(\configuration[45] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold287 (.A(\vga.timing_v.pixel[6] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold288 (.A(\mandelbrot.alu.in_cr[6] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold289 (.A(\mandelbrot.y[5] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0122_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold291 (.A(\mandelbrot.ctr[7] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold292 (.A(uio_out[1]),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold293 (.A(\mandelbrot.alu.in_zi[8] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold294 (.A(\mandelbrot.y[7] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0124_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold296 (.A(\configuration[46] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold297 (.A(\mandelbrot.alu.in_zr[1] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold298 (.A(\mandelbrot.alu.m3[6] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold299 (.A(_0927_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold300 (.A(\vga.pixel_ctr[6] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0454_),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0013_),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold303 (.A(\mandelbrot.alu.in_zr[4] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold304 (.A(_1282_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold305 (.A(\mandelbrot.alu.m1[2] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold306 (.A(_0128_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold307 (.A(\mandelbrot.alu.m3[21] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0287_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold309 (.A(uio_out[2]),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold310 (.A(_0362_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold311 (.A(\mandelbrot.ctr[6] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold312 (.A(\vga.pixel_ctr[4] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold313 (.A(_0451_),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold314 (.A(\mandelbrot.alu.in_ci[8] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold315 (.A(\mandelbrot.ctr[3] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold316 (.A(\mandelbrot.alu.in_ci[1] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold317 (.A(\mandelbrot.alu.mult_zr_zi.running ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold318 (.A(\vga.pixel_ctr[0] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold319 (.A(\mandelbrot.alu.m1[5] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0131_),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold321 (.A(\mandelbrot.alu.m3[30] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold322 (.A(\mandelbrot.alu.in_ci[6] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold323 (.A(\mandelbrot.ctr[2] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold324 (.A(\mandelbrot.alu.in_ci[10] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold325 (.A(\mandelbrot.alu.in_ci[5] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold326 (.A(\mandelbrot.alu.in_cr[13] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold327 (.A(_0356_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold328 (.A(\mandelbrot.alu.first_iteration ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold329 (.A(\mandelbrot.alu.m1[14] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold330 (.A(_0140_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold331 (.A(\mandelbrot.alu.in_ci[4] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold332 (.A(\mandelbrot.alu.mult_zr_zr.shift_reg[0] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold333 (.A(\mandelbrot.alu.m2[9] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold334 (.A(_0237_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold335 (.A(\mandelbrot.alu.m3[19] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold336 (.A(_0285_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold337 (.A(\vga.pixel_ctr[9] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold338 (.A(_0458_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold339 (.A(\mandelbrot.alu.m1[13] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold340 (.A(\mandelbrot.alu.m1[6] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold341 (.A(_1665_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold342 (.A(\mandelbrot.alu.m3[3] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold343 (.A(_0887_),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold344 (.A(\mandelbrot.alu.m2[5] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0233_),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold346 (.A(\mandelbrot.alu.in_ci[12] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold347 (.A(\mandelbrot.alu.in_cr[11] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0354_),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold349 (.A(\mandelbrot.ctr[9] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold350 (.A(\mandelbrot.alu.in_cr[0] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0096_),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0248_),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold353 (.A(\configuration[32] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold354 (.A(\mandelbrot.alu.in_cr[15] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0358_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold356 (.A(\mandelbrot.ctr[1] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0334_),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold358 (.A(\mandelbrot.alu.m1[15] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0107_),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold360 (.A(\mandelbrot.alu.in_cr[12] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold361 (.A(\mandelbrot.alu.m2[3] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold362 (.A(\mandelbrot.alu.in_ci[15] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold363 (.A(\mandelbrot.alu.m3[14] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold364 (.A(_0280_),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold365 (.A(\vga.timing_v.pixel[3] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold366 (.A(\mandelbrot.alu.in_ci[14] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold367 (.A(\mandelbrot.alu.m2[2] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold368 (.A(_0521_),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold369 (.A(\mandelbrot.ctr[8] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold370 (.A(\mandelbrot.alu.m2[4] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold371 (.A(_0232_),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold372 (.A(\mandelbrot.alu.m1[4] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold373 (.A(\mandelbrot.alu.m3[29] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold374 (.A(\mandelbrot.alu.m2[11] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold375 (.A(_0239_),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold376 (.A(\vga.pixel_buffer[0] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold377 (.A(_0212_),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold378 (.A(\mandelbrot.alu.m2[13] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold379 (.A(_0241_),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0094_),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold381 (.A(_0251_),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold382 (.A(\vga.pixel_buffer[1] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold383 (.A(_0213_),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold384 (.A(\mandelbrot.alu.m1[10] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold385 (.A(_1670_),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold386 (.A(\vga.timing_v.pixel[2] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold387 (.A(\mandelbrot.alu.m3[23] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold388 (.A(_0289_),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold389 (.A(_0023_),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold390 (.A(_0151_),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold391 (.A(\mandelbrot.alu.m1[28] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold392 (.A(_0156_),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold393 (.A(\mandelbrot.alu.m1[8] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold394 (.A(\mandelbrot.alu.m2[6] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold395 (.A(_0234_),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold396 (.A(\mandelbrot.alu.m2[0] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold397 (.A(\mandelbrot.alu.in_ci[2] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold398 (.A(\mandelbrot.alu.m1[16] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold399 (.A(\mandelbrot.alu.in_cr[4] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold400 (.A(_0347_),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold401 (.A(\mandelbrot.alu.in_ci[13] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold402 (.A(\mandelbrot.alu.in_ci[0] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold403 (.A(_0020_),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold404 (.A(_0155_),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold405 (.A(\mandelbrot.alu.m2[8] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold406 (.A(\mandelbrot.alu.in_zr[0] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold407 (.A(\mandelbrot.alu.in_zr[5] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold408 (.A(\mandelbrot.ctr[4] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold409 (.A(\configuration[41] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold410 (.A(_0199_),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold411 (.A(\configuration[35] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold412 (.A(_0193_),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold413 (.A(\mandelbrot.alu.m1[31] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold414 (.A(_0216_),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold415 (.A(uio_out[0]),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold416 (.A(\vga.pixel_ctr[1] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold417 (.A(_0008_),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold418 (.A(\mandelbrot.alu.mult_zr_zi.ctr[0] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold419 (.A(\vga.pixel_ctr[10] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold420 (.A(\vga.read ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold421 (.A(\mandelbrot.alu.m2[1] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold422 (.A(_0229_),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold423 (.A(\configuration[33] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold424 (.A(\configuration[34] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold425 (.A(\mandelbrot.alu.m1[7] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold426 (.A(\mandelbrot.alu.m2[12] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold427 (.A(uio_out[3]),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold428 (.A(\mandelbrot.alu.in_cr[2] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold429 (.A(\mandelbrot.alu.m2[7] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold430 (.A(\configuration[39] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold431 (.A(_0198_),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold432 (.A(\mandelbrot.alu.m1[29] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold433 (.A(\configuration[38] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold434 (.A(\mandelbrot.alu.m2[10] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold435 (.A(\configuration[37] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold436 (.A(_0195_),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold437 (.A(\mandelbrot.alu.m1[30] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold438 (.A(\configuration[36] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold439 (.A(\mandelbrot.run ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold440 (.A(_0005_),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold441 (.A(\mandelbrot.alu.m2[19] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold442 (.A(_0247_),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold443 (.A(\mandelbrot.alu.m1[3] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold444 (.A(_1659_),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold445 (.A(\mandelbrot.alu.in_zi[0] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold446 (.A(_0098_),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold447 (.A(_0246_),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold448 (.A(\mandelbrot.alu.m1[9] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold449 (.A(\mandelbrot.alu.m2[14] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold450 (.A(\mandelbrot.alu.m2[15] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold451 (.A(_0105_),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold452 (.A(_1270_),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold453 (.A(_0300_),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold454 (.A(\mandelbrot.ctr[1] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold455 (.A(\mandelbrot.ctr[4] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold456 (.A(\vga.pixel_ctr[10] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold457 (.A(_0105_),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold458 (.A(\mandelbrot.ctr[8] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold459 (.A(\mandelbrot.alu.m2[10] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold460 (.A(\mandelbrot.alu.in_ci[14] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold461 (.A(\mandelbrot.alu.m2[14] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold462 (.A(\vga.pixel_ctr[10] ),
    .X(net828));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_fill_2 FILLER_0_105 ();
 sg13g2_fill_1 FILLER_0_107 ();
 sg13g2_fill_2 FILLER_0_122 ();
 sg13g2_fill_1 FILLER_0_124 ();
 sg13g2_decap_4 FILLER_0_138 ();
 sg13g2_fill_2 FILLER_0_142 ();
 sg13g2_fill_2 FILLER_0_177 ();
 sg13g2_fill_1 FILLER_0_188 ();
 sg13g2_decap_8 FILLER_0_199 ();
 sg13g2_decap_8 FILLER_0_206 ();
 sg13g2_decap_8 FILLER_0_213 ();
 sg13g2_fill_1 FILLER_0_220 ();
 sg13g2_decap_8 FILLER_0_225 ();
 sg13g2_decap_8 FILLER_0_232 ();
 sg13g2_decap_8 FILLER_0_239 ();
 sg13g2_decap_4 FILLER_0_246 ();
 sg13g2_fill_1 FILLER_0_250 ();
 sg13g2_decap_4 FILLER_0_255 ();
 sg13g2_fill_2 FILLER_0_263 ();
 sg13g2_decap_4 FILLER_0_270 ();
 sg13g2_fill_1 FILLER_0_274 ();
 sg13g2_fill_1 FILLER_0_279 ();
 sg13g2_fill_2 FILLER_0_284 ();
 sg13g2_decap_8 FILLER_0_290 ();
 sg13g2_decap_8 FILLER_0_297 ();
 sg13g2_decap_8 FILLER_0_304 ();
 sg13g2_fill_2 FILLER_0_311 ();
 sg13g2_fill_1 FILLER_0_313 ();
 sg13g2_decap_4 FILLER_0_318 ();
 sg13g2_fill_2 FILLER_0_322 ();
 sg13g2_decap_4 FILLER_0_327 ();
 sg13g2_fill_1 FILLER_0_331 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_4 FILLER_1_95 ();
 sg13g2_fill_1 FILLER_1_146 ();
 sg13g2_fill_2 FILLER_1_213 ();
 sg13g2_fill_1 FILLER_1_220 ();
 sg13g2_decap_4 FILLER_1_234 ();
 sg13g2_fill_1 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_302 ();
 sg13g2_fill_1 FILLER_1_317 ();
 sg13g2_fill_1 FILLER_1_340 ();
 sg13g2_decap_8 FILLER_1_367 ();
 sg13g2_decap_8 FILLER_1_374 ();
 sg13g2_decap_8 FILLER_1_381 ();
 sg13g2_decap_8 FILLER_1_388 ();
 sg13g2_decap_8 FILLER_1_395 ();
 sg13g2_decap_8 FILLER_1_402 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_4 FILLER_2_77 ();
 sg13g2_fill_1 FILLER_2_112 ();
 sg13g2_decap_4 FILLER_2_165 ();
 sg13g2_fill_1 FILLER_2_198 ();
 sg13g2_fill_2 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_381 ();
 sg13g2_decap_8 FILLER_2_388 ();
 sg13g2_decap_8 FILLER_2_395 ();
 sg13g2_decap_8 FILLER_2_402 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_4 FILLER_3_70 ();
 sg13g2_fill_1 FILLER_3_74 ();
 sg13g2_fill_2 FILLER_3_147 ();
 sg13g2_fill_1 FILLER_3_165 ();
 sg13g2_fill_1 FILLER_3_171 ();
 sg13g2_fill_1 FILLER_3_185 ();
 sg13g2_fill_1 FILLER_3_194 ();
 sg13g2_fill_2 FILLER_3_207 ();
 sg13g2_fill_1 FILLER_3_209 ();
 sg13g2_fill_1 FILLER_3_223 ();
 sg13g2_fill_2 FILLER_3_250 ();
 sg13g2_fill_1 FILLER_3_266 ();
 sg13g2_fill_2 FILLER_3_314 ();
 sg13g2_fill_1 FILLER_3_349 ();
 sg13g2_decap_8 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_4 FILLER_3_403 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_4 FILLER_4_63 ();
 sg13g2_fill_1 FILLER_4_67 ();
 sg13g2_fill_1 FILLER_4_101 ();
 sg13g2_fill_2 FILLER_4_117 ();
 sg13g2_fill_2 FILLER_4_152 ();
 sg13g2_fill_1 FILLER_4_181 ();
 sg13g2_fill_1 FILLER_4_191 ();
 sg13g2_fill_2 FILLER_4_212 ();
 sg13g2_decap_4 FILLER_4_222 ();
 sg13g2_fill_2 FILLER_4_226 ();
 sg13g2_fill_2 FILLER_4_243 ();
 sg13g2_fill_1 FILLER_4_258 ();
 sg13g2_fill_2 FILLER_4_276 ();
 sg13g2_decap_4 FILLER_4_282 ();
 sg13g2_decap_8 FILLER_4_290 ();
 sg13g2_decap_8 FILLER_4_297 ();
 sg13g2_fill_1 FILLER_4_304 ();
 sg13g2_fill_2 FILLER_4_322 ();
 sg13g2_fill_2 FILLER_4_328 ();
 sg13g2_fill_2 FILLER_4_346 ();
 sg13g2_fill_1 FILLER_4_348 ();
 sg13g2_decap_8 FILLER_4_376 ();
 sg13g2_decap_8 FILLER_4_383 ();
 sg13g2_decap_8 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_397 ();
 sg13g2_decap_4 FILLER_4_404 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_fill_2 FILLER_5_70 ();
 sg13g2_decap_4 FILLER_5_187 ();
 sg13g2_fill_2 FILLER_5_191 ();
 sg13g2_fill_2 FILLER_5_197 ();
 sg13g2_fill_1 FILLER_5_199 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_fill_2 FILLER_5_224 ();
 sg13g2_fill_1 FILLER_5_226 ();
 sg13g2_fill_1 FILLER_5_255 ();
 sg13g2_fill_2 FILLER_5_269 ();
 sg13g2_fill_1 FILLER_5_276 ();
 sg13g2_fill_2 FILLER_5_281 ();
 sg13g2_decap_4 FILLER_5_296 ();
 sg13g2_fill_2 FILLER_5_314 ();
 sg13g2_decap_4 FILLER_5_347 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_fill_2 FILLER_6_108 ();
 sg13g2_fill_2 FILLER_6_119 ();
 sg13g2_fill_1 FILLER_6_134 ();
 sg13g2_fill_2 FILLER_6_173 ();
 sg13g2_decap_4 FILLER_6_185 ();
 sg13g2_fill_1 FILLER_6_189 ();
 sg13g2_fill_2 FILLER_6_195 ();
 sg13g2_fill_1 FILLER_6_197 ();
 sg13g2_fill_1 FILLER_6_215 ();
 sg13g2_fill_2 FILLER_6_251 ();
 sg13g2_fill_1 FILLER_6_253 ();
 sg13g2_fill_2 FILLER_6_328 ();
 sg13g2_fill_1 FILLER_6_330 ();
 sg13g2_fill_2 FILLER_6_345 ();
 sg13g2_fill_1 FILLER_6_347 ();
 sg13g2_decap_8 FILLER_6_381 ();
 sg13g2_decap_8 FILLER_6_388 ();
 sg13g2_decap_8 FILLER_6_395 ();
 sg13g2_decap_8 FILLER_6_402 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_4 FILLER_7_70 ();
 sg13g2_fill_1 FILLER_7_74 ();
 sg13g2_fill_1 FILLER_7_102 ();
 sg13g2_fill_2 FILLER_7_134 ();
 sg13g2_fill_2 FILLER_7_179 ();
 sg13g2_fill_1 FILLER_7_181 ();
 sg13g2_decap_4 FILLER_7_187 ();
 sg13g2_fill_1 FILLER_7_198 ();
 sg13g2_fill_2 FILLER_7_208 ();
 sg13g2_fill_1 FILLER_7_210 ();
 sg13g2_decap_4 FILLER_7_226 ();
 sg13g2_fill_1 FILLER_7_230 ();
 sg13g2_fill_2 FILLER_7_271 ();
 sg13g2_fill_1 FILLER_7_277 ();
 sg13g2_decap_8 FILLER_7_328 ();
 sg13g2_fill_2 FILLER_7_335 ();
 sg13g2_fill_1 FILLER_7_337 ();
 sg13g2_fill_2 FILLER_7_346 ();
 sg13g2_fill_1 FILLER_7_348 ();
 sg13g2_decap_8 FILLER_7_373 ();
 sg13g2_decap_8 FILLER_7_380 ();
 sg13g2_decap_8 FILLER_7_387 ();
 sg13g2_decap_8 FILLER_7_394 ();
 sg13g2_decap_8 FILLER_7_401 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_4 FILLER_8_70 ();
 sg13g2_fill_1 FILLER_8_74 ();
 sg13g2_fill_2 FILLER_8_109 ();
 sg13g2_fill_1 FILLER_8_111 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_fill_1 FILLER_8_161 ();
 sg13g2_fill_2 FILLER_8_180 ();
 sg13g2_fill_1 FILLER_8_182 ();
 sg13g2_fill_2 FILLER_8_209 ();
 sg13g2_fill_1 FILLER_8_249 ();
 sg13g2_fill_2 FILLER_8_258 ();
 sg13g2_fill_1 FILLER_8_260 ();
 sg13g2_decap_8 FILLER_8_270 ();
 sg13g2_fill_1 FILLER_8_281 ();
 sg13g2_decap_8 FILLER_8_312 ();
 sg13g2_fill_2 FILLER_8_319 ();
 sg13g2_fill_1 FILLER_8_321 ();
 sg13g2_decap_8 FILLER_8_388 ();
 sg13g2_decap_8 FILLER_8_395 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_fill_1 FILLER_9_77 ();
 sg13g2_fill_1 FILLER_9_91 ();
 sg13g2_fill_2 FILLER_9_105 ();
 sg13g2_fill_1 FILLER_9_107 ();
 sg13g2_fill_2 FILLER_9_118 ();
 sg13g2_decap_4 FILLER_9_133 ();
 sg13g2_fill_2 FILLER_9_137 ();
 sg13g2_decap_8 FILLER_9_143 ();
 sg13g2_decap_8 FILLER_9_150 ();
 sg13g2_decap_8 FILLER_9_157 ();
 sg13g2_decap_8 FILLER_9_164 ();
 sg13g2_fill_2 FILLER_9_174 ();
 sg13g2_fill_2 FILLER_9_207 ();
 sg13g2_fill_1 FILLER_9_233 ();
 sg13g2_decap_8 FILLER_9_239 ();
 sg13g2_decap_8 FILLER_9_246 ();
 sg13g2_decap_8 FILLER_9_253 ();
 sg13g2_decap_4 FILLER_9_260 ();
 sg13g2_fill_2 FILLER_9_264 ();
 sg13g2_decap_4 FILLER_9_270 ();
 sg13g2_fill_1 FILLER_9_274 ();
 sg13g2_decap_4 FILLER_9_307 ();
 sg13g2_fill_1 FILLER_9_311 ();
 sg13g2_fill_1 FILLER_9_319 ();
 sg13g2_fill_1 FILLER_9_341 ();
 sg13g2_decap_8 FILLER_9_372 ();
 sg13g2_decap_8 FILLER_9_379 ();
 sg13g2_decap_8 FILLER_9_386 ();
 sg13g2_decap_8 FILLER_9_393 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_fill_2 FILLER_10_77 ();
 sg13g2_decap_4 FILLER_10_98 ();
 sg13g2_fill_2 FILLER_10_102 ();
 sg13g2_fill_1 FILLER_10_121 ();
 sg13g2_fill_2 FILLER_10_126 ();
 sg13g2_fill_1 FILLER_10_128 ();
 sg13g2_fill_2 FILLER_10_163 ();
 sg13g2_decap_4 FILLER_10_183 ();
 sg13g2_fill_1 FILLER_10_187 ();
 sg13g2_fill_2 FILLER_10_200 ();
 sg13g2_fill_2 FILLER_10_223 ();
 sg13g2_fill_2 FILLER_10_239 ();
 sg13g2_decap_4 FILLER_10_250 ();
 sg13g2_fill_2 FILLER_10_254 ();
 sg13g2_fill_1 FILLER_10_264 ();
 sg13g2_fill_1 FILLER_10_299 ();
 sg13g2_fill_2 FILLER_10_346 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_fill_2 FILLER_11_70 ();
 sg13g2_fill_1 FILLER_11_120 ();
 sg13g2_fill_1 FILLER_11_199 ();
 sg13g2_fill_1 FILLER_11_209 ();
 sg13g2_decap_4 FILLER_11_223 ();
 sg13g2_fill_2 FILLER_11_227 ();
 sg13g2_fill_2 FILLER_11_281 ();
 sg13g2_decap_4 FILLER_11_300 ();
 sg13g2_fill_2 FILLER_11_334 ();
 sg13g2_fill_2 FILLER_11_356 ();
 sg13g2_fill_2 FILLER_11_366 ();
 sg13g2_decap_8 FILLER_11_387 ();
 sg13g2_decap_8 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_fill_1 FILLER_12_102 ();
 sg13g2_fill_2 FILLER_12_137 ();
 sg13g2_fill_1 FILLER_12_139 ();
 sg13g2_fill_1 FILLER_12_184 ();
 sg13g2_fill_2 FILLER_12_204 ();
 sg13g2_fill_1 FILLER_12_214 ();
 sg13g2_decap_4 FILLER_12_228 ();
 sg13g2_fill_2 FILLER_12_242 ();
 sg13g2_fill_2 FILLER_12_307 ();
 sg13g2_fill_1 FILLER_12_309 ();
 sg13g2_fill_1 FILLER_12_319 ();
 sg13g2_fill_2 FILLER_12_360 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_fill_2 FILLER_13_126 ();
 sg13g2_fill_1 FILLER_13_128 ();
 sg13g2_fill_2 FILLER_13_167 ();
 sg13g2_fill_1 FILLER_13_169 ();
 sg13g2_fill_2 FILLER_13_198 ();
 sg13g2_fill_1 FILLER_13_200 ();
 sg13g2_fill_2 FILLER_13_207 ();
 sg13g2_fill_1 FILLER_13_209 ();
 sg13g2_decap_8 FILLER_13_234 ();
 sg13g2_fill_2 FILLER_13_241 ();
 sg13g2_fill_1 FILLER_13_243 ();
 sg13g2_decap_8 FILLER_13_248 ();
 sg13g2_decap_4 FILLER_13_255 ();
 sg13g2_decap_8 FILLER_13_267 ();
 sg13g2_fill_2 FILLER_13_274 ();
 sg13g2_fill_1 FILLER_13_287 ();
 sg13g2_fill_1 FILLER_13_301 ();
 sg13g2_fill_1 FILLER_13_307 ();
 sg13g2_decap_8 FILLER_13_374 ();
 sg13g2_decap_8 FILLER_13_381 ();
 sg13g2_decap_8 FILLER_13_388 ();
 sg13g2_decap_8 FILLER_13_395 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_fill_2 FILLER_14_77 ();
 sg13g2_fill_1 FILLER_14_89 ();
 sg13g2_fill_2 FILLER_14_104 ();
 sg13g2_fill_2 FILLER_14_138 ();
 sg13g2_decap_8 FILLER_14_149 ();
 sg13g2_fill_1 FILLER_14_194 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_4 FILLER_14_210 ();
 sg13g2_fill_2 FILLER_14_214 ();
 sg13g2_fill_2 FILLER_14_229 ();
 sg13g2_fill_1 FILLER_14_231 ();
 sg13g2_fill_1 FILLER_14_262 ();
 sg13g2_fill_2 FILLER_14_312 ();
 sg13g2_fill_1 FILLER_14_314 ();
 sg13g2_decap_8 FILLER_14_342 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_4 FILLER_15_103 ();
 sg13g2_fill_1 FILLER_15_107 ();
 sg13g2_decap_4 FILLER_15_117 ();
 sg13g2_fill_1 FILLER_15_121 ();
 sg13g2_decap_8 FILLER_15_156 ();
 sg13g2_fill_2 FILLER_15_163 ();
 sg13g2_decap_8 FILLER_15_198 ();
 sg13g2_decap_4 FILLER_15_205 ();
 sg13g2_decap_8 FILLER_15_222 ();
 sg13g2_fill_2 FILLER_15_229 ();
 sg13g2_fill_1 FILLER_15_240 ();
 sg13g2_decap_4 FILLER_15_267 ();
 sg13g2_fill_2 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_fill_1 FILLER_15_322 ();
 sg13g2_decap_4 FILLER_15_327 ();
 sg13g2_fill_2 FILLER_15_341 ();
 sg13g2_fill_1 FILLER_15_347 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_fill_2 FILLER_16_77 ();
 sg13g2_fill_1 FILLER_16_88 ();
 sg13g2_decap_4 FILLER_16_124 ();
 sg13g2_decap_4 FILLER_16_132 ();
 sg13g2_fill_1 FILLER_16_136 ();
 sg13g2_fill_2 FILLER_16_158 ();
 sg13g2_fill_1 FILLER_16_160 ();
 sg13g2_fill_2 FILLER_16_253 ();
 sg13g2_fill_2 FILLER_16_300 ();
 sg13g2_fill_2 FILLER_16_318 ();
 sg13g2_fill_1 FILLER_16_329 ();
 sg13g2_fill_1 FILLER_16_343 ();
 sg13g2_fill_2 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_fill_1 FILLER_17_103 ();
 sg13g2_fill_1 FILLER_17_116 ();
 sg13g2_fill_2 FILLER_17_189 ();
 sg13g2_fill_1 FILLER_17_191 ();
 sg13g2_decap_8 FILLER_17_212 ();
 sg13g2_fill_1 FILLER_17_219 ();
 sg13g2_fill_1 FILLER_17_251 ();
 sg13g2_fill_2 FILLER_17_257 ();
 sg13g2_decap_8 FILLER_17_278 ();
 sg13g2_decap_4 FILLER_17_285 ();
 sg13g2_fill_2 FILLER_17_301 ();
 sg13g2_fill_1 FILLER_17_303 ();
 sg13g2_decap_4 FILLER_17_330 ();
 sg13g2_fill_1 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_394 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_4 FILLER_18_63 ();
 sg13g2_fill_2 FILLER_18_91 ();
 sg13g2_fill_1 FILLER_18_93 ();
 sg13g2_fill_2 FILLER_18_103 ();
 sg13g2_fill_1 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_124 ();
 sg13g2_fill_1 FILLER_18_131 ();
 sg13g2_fill_2 FILLER_18_141 ();
 sg13g2_fill_2 FILLER_18_158 ();
 sg13g2_fill_1 FILLER_18_160 ();
 sg13g2_fill_1 FILLER_18_184 ();
 sg13g2_fill_2 FILLER_18_205 ();
 sg13g2_fill_2 FILLER_18_231 ();
 sg13g2_fill_1 FILLER_18_238 ();
 sg13g2_decap_4 FILLER_18_275 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_4 FILLER_19_70 ();
 sg13g2_fill_2 FILLER_19_108 ();
 sg13g2_fill_1 FILLER_19_110 ();
 sg13g2_decap_8 FILLER_19_130 ();
 sg13g2_decap_4 FILLER_19_137 ();
 sg13g2_fill_1 FILLER_19_173 ();
 sg13g2_fill_2 FILLER_19_183 ();
 sg13g2_fill_2 FILLER_19_266 ();
 sg13g2_fill_1 FILLER_19_268 ();
 sg13g2_fill_1 FILLER_19_328 ();
 sg13g2_fill_1 FILLER_19_338 ();
 sg13g2_fill_2 FILLER_19_352 ();
 sg13g2_fill_1 FILLER_19_377 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_4 FILLER_20_77 ();
 sg13g2_fill_1 FILLER_20_81 ();
 sg13g2_fill_1 FILLER_20_91 ();
 sg13g2_fill_2 FILLER_20_96 ();
 sg13g2_fill_1 FILLER_20_124 ();
 sg13g2_decap_4 FILLER_20_215 ();
 sg13g2_fill_2 FILLER_20_219 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_fill_2 FILLER_20_256 ();
 sg13g2_fill_1 FILLER_20_258 ();
 sg13g2_decap_8 FILLER_20_271 ();
 sg13g2_fill_2 FILLER_20_278 ();
 sg13g2_fill_2 FILLER_20_284 ();
 sg13g2_fill_2 FILLER_20_306 ();
 sg13g2_fill_1 FILLER_20_308 ();
 sg13g2_fill_2 FILLER_20_335 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_4 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_fill_2 FILLER_21_77 ();
 sg13g2_fill_1 FILLER_21_111 ();
 sg13g2_fill_1 FILLER_21_121 ();
 sg13g2_fill_1 FILLER_21_130 ();
 sg13g2_fill_1 FILLER_21_150 ();
 sg13g2_fill_1 FILLER_21_180 ();
 sg13g2_fill_2 FILLER_21_202 ();
 sg13g2_decap_8 FILLER_21_230 ();
 sg13g2_decap_8 FILLER_21_237 ();
 sg13g2_decap_4 FILLER_21_244 ();
 sg13g2_fill_1 FILLER_21_257 ();
 sg13g2_fill_1 FILLER_21_263 ();
 sg13g2_fill_1 FILLER_21_285 ();
 sg13g2_fill_1 FILLER_21_296 ();
 sg13g2_fill_1 FILLER_21_321 ();
 sg13g2_fill_2 FILLER_21_332 ();
 sg13g2_fill_1 FILLER_21_334 ();
 sg13g2_fill_1 FILLER_21_340 ();
 sg13g2_fill_2 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_389 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_fill_2 FILLER_22_70 ();
 sg13g2_fill_2 FILLER_22_122 ();
 sg13g2_fill_1 FILLER_22_124 ();
 sg13g2_fill_1 FILLER_22_139 ();
 sg13g2_fill_2 FILLER_22_144 ();
 sg13g2_fill_1 FILLER_22_146 ();
 sg13g2_fill_1 FILLER_22_167 ();
 sg13g2_decap_4 FILLER_22_210 ();
 sg13g2_fill_2 FILLER_22_222 ();
 sg13g2_fill_1 FILLER_22_224 ();
 sg13g2_decap_4 FILLER_22_235 ();
 sg13g2_fill_2 FILLER_22_252 ();
 sg13g2_fill_1 FILLER_22_254 ();
 sg13g2_fill_2 FILLER_22_325 ();
 sg13g2_fill_1 FILLER_22_327 ();
 sg13g2_fill_1 FILLER_22_336 ();
 sg13g2_fill_2 FILLER_22_347 ();
 sg13g2_fill_1 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_358 ();
 sg13g2_fill_1 FILLER_22_365 ();
 sg13g2_fill_1 FILLER_22_374 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_4 FILLER_23_63 ();
 sg13g2_fill_1 FILLER_23_67 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_4 FILLER_23_119 ();
 sg13g2_fill_2 FILLER_23_123 ();
 sg13g2_decap_4 FILLER_23_155 ();
 sg13g2_fill_2 FILLER_23_159 ();
 sg13g2_fill_1 FILLER_23_171 ();
 sg13g2_fill_2 FILLER_23_183 ();
 sg13g2_fill_1 FILLER_23_204 ();
 sg13g2_fill_1 FILLER_23_213 ();
 sg13g2_fill_1 FILLER_23_219 ();
 sg13g2_fill_1 FILLER_23_228 ();
 sg13g2_fill_2 FILLER_23_255 ();
 sg13g2_fill_1 FILLER_23_257 ();
 sg13g2_decap_4 FILLER_23_340 ();
 sg13g2_decap_4 FILLER_23_370 ();
 sg13g2_decap_8 FILLER_23_395 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_fill_2 FILLER_24_70 ();
 sg13g2_fill_1 FILLER_24_72 ();
 sg13g2_decap_4 FILLER_24_109 ();
 sg13g2_fill_1 FILLER_24_113 ();
 sg13g2_fill_2 FILLER_24_123 ();
 sg13g2_fill_2 FILLER_24_135 ();
 sg13g2_fill_2 FILLER_24_166 ();
 sg13g2_fill_1 FILLER_24_168 ();
 sg13g2_fill_1 FILLER_24_208 ();
 sg13g2_decap_4 FILLER_24_221 ();
 sg13g2_fill_2 FILLER_24_225 ();
 sg13g2_fill_1 FILLER_24_232 ();
 sg13g2_fill_1 FILLER_24_238 ();
 sg13g2_fill_1 FILLER_24_260 ();
 sg13g2_decap_4 FILLER_24_265 ();
 sg13g2_fill_2 FILLER_24_307 ();
 sg13g2_fill_1 FILLER_24_309 ();
 sg13g2_fill_1 FILLER_24_337 ();
 sg13g2_fill_2 FILLER_24_351 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_fill_2 FILLER_25_77 ();
 sg13g2_decap_4 FILLER_25_83 ();
 sg13g2_decap_4 FILLER_25_110 ();
 sg13g2_fill_1 FILLER_25_119 ();
 sg13g2_fill_1 FILLER_25_138 ();
 sg13g2_fill_1 FILLER_25_148 ();
 sg13g2_fill_2 FILLER_25_165 ();
 sg13g2_fill_1 FILLER_25_206 ();
 sg13g2_fill_2 FILLER_25_222 ();
 sg13g2_fill_1 FILLER_25_224 ();
 sg13g2_fill_2 FILLER_25_257 ();
 sg13g2_fill_2 FILLER_25_279 ();
 sg13g2_fill_1 FILLER_25_281 ();
 sg13g2_fill_2 FILLER_25_289 ();
 sg13g2_fill_1 FILLER_25_291 ();
 sg13g2_fill_2 FILLER_25_333 ();
 sg13g2_fill_1 FILLER_25_347 ();
 sg13g2_fill_2 FILLER_25_361 ();
 sg13g2_fill_1 FILLER_25_363 ();
 sg13g2_fill_2 FILLER_25_380 ();
 sg13g2_decap_8 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_fill_1 FILLER_26_77 ();
 sg13g2_fill_2 FILLER_26_96 ();
 sg13g2_fill_1 FILLER_26_103 ();
 sg13g2_fill_1 FILLER_26_129 ();
 sg13g2_decap_4 FILLER_26_156 ();
 sg13g2_fill_2 FILLER_26_194 ();
 sg13g2_fill_1 FILLER_26_204 ();
 sg13g2_fill_2 FILLER_26_234 ();
 sg13g2_fill_1 FILLER_26_236 ();
 sg13g2_fill_1 FILLER_26_247 ();
 sg13g2_fill_2 FILLER_26_256 ();
 sg13g2_fill_1 FILLER_26_258 ();
 sg13g2_fill_2 FILLER_26_304 ();
 sg13g2_fill_2 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_391 ();
 sg13g2_decap_8 FILLER_26_398 ();
 sg13g2_decap_4 FILLER_26_405 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_fill_2 FILLER_27_63 ();
 sg13g2_fill_1 FILLER_27_65 ();
 sg13g2_fill_1 FILLER_27_125 ();
 sg13g2_decap_4 FILLER_27_175 ();
 sg13g2_fill_2 FILLER_27_179 ();
 sg13g2_fill_2 FILLER_27_200 ();
 sg13g2_fill_2 FILLER_27_210 ();
 sg13g2_fill_2 FILLER_27_264 ();
 sg13g2_fill_1 FILLER_27_266 ();
 sg13g2_fill_1 FILLER_27_377 ();
 sg13g2_decap_8 FILLER_27_397 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_fill_1 FILLER_28_75 ();
 sg13g2_fill_2 FILLER_28_145 ();
 sg13g2_decap_8 FILLER_28_151 ();
 sg13g2_decap_8 FILLER_28_163 ();
 sg13g2_decap_4 FILLER_28_170 ();
 sg13g2_fill_1 FILLER_28_174 ();
 sg13g2_fill_2 FILLER_28_204 ();
 sg13g2_fill_1 FILLER_28_206 ();
 sg13g2_decap_8 FILLER_28_215 ();
 sg13g2_decap_4 FILLER_28_222 ();
 sg13g2_fill_1 FILLER_28_226 ();
 sg13g2_fill_2 FILLER_28_231 ();
 sg13g2_decap_4 FILLER_28_238 ();
 sg13g2_fill_2 FILLER_28_255 ();
 sg13g2_fill_1 FILLER_28_257 ();
 sg13g2_fill_1 FILLER_28_350 ();
 sg13g2_fill_1 FILLER_28_360 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_fill_2 FILLER_29_49 ();
 sg13g2_fill_2 FILLER_29_66 ();
 sg13g2_fill_1 FILLER_29_68 ();
 sg13g2_fill_2 FILLER_29_105 ();
 sg13g2_fill_2 FILLER_29_126 ();
 sg13g2_fill_1 FILLER_29_142 ();
 sg13g2_decap_8 FILLER_29_156 ();
 sg13g2_decap_8 FILLER_29_163 ();
 sg13g2_decap_4 FILLER_29_170 ();
 sg13g2_fill_2 FILLER_29_174 ();
 sg13g2_decap_8 FILLER_29_206 ();
 sg13g2_decap_4 FILLER_29_213 ();
 sg13g2_fill_1 FILLER_29_217 ();
 sg13g2_fill_2 FILLER_29_226 ();
 sg13g2_fill_1 FILLER_29_228 ();
 sg13g2_fill_2 FILLER_29_251 ();
 sg13g2_fill_1 FILLER_29_342 ();
 sg13g2_fill_2 FILLER_29_360 ();
 sg13g2_fill_1 FILLER_29_362 ();
 sg13g2_decap_8 FILLER_29_388 ();
 sg13g2_decap_8 FILLER_29_395 ();
 sg13g2_decap_8 FILLER_29_402 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_fill_1 FILLER_30_28 ();
 sg13g2_fill_2 FILLER_30_40 ();
 sg13g2_fill_1 FILLER_30_42 ();
 sg13g2_fill_2 FILLER_30_69 ();
 sg13g2_fill_1 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_99 ();
 sg13g2_fill_1 FILLER_30_101 ();
 sg13g2_decap_4 FILLER_30_192 ();
 sg13g2_fill_2 FILLER_30_196 ();
 sg13g2_fill_2 FILLER_30_202 ();
 sg13g2_fill_1 FILLER_30_204 ();
 sg13g2_fill_2 FILLER_30_215 ();
 sg13g2_fill_1 FILLER_30_217 ();
 sg13g2_fill_2 FILLER_30_310 ();
 sg13g2_fill_2 FILLER_30_331 ();
 sg13g2_fill_1 FILLER_30_333 ();
 sg13g2_fill_2 FILLER_30_357 ();
 sg13g2_fill_1 FILLER_30_359 ();
 sg13g2_decap_8 FILLER_30_397 ();
 sg13g2_decap_4 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_fill_2 FILLER_31_21 ();
 sg13g2_fill_1 FILLER_31_36 ();
 sg13g2_fill_1 FILLER_31_72 ();
 sg13g2_fill_2 FILLER_31_124 ();
 sg13g2_fill_1 FILLER_31_126 ();
 sg13g2_fill_2 FILLER_31_135 ();
 sg13g2_fill_1 FILLER_31_137 ();
 sg13g2_fill_1 FILLER_31_168 ();
 sg13g2_fill_1 FILLER_31_198 ();
 sg13g2_fill_1 FILLER_31_231 ();
 sg13g2_fill_2 FILLER_31_267 ();
 sg13g2_fill_2 FILLER_31_275 ();
 sg13g2_fill_1 FILLER_31_277 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_4 ();
 sg13g2_decap_8 FILLER_32_9 ();
 sg13g2_fill_1 FILLER_32_54 ();
 sg13g2_fill_1 FILLER_32_164 ();
 sg13g2_fill_2 FILLER_32_251 ();
 sg13g2_fill_2 FILLER_32_275 ();
 sg13g2_fill_1 FILLER_32_277 ();
 sg13g2_fill_2 FILLER_32_321 ();
 sg13g2_fill_1 FILLER_32_323 ();
 sg13g2_decap_8 FILLER_32_332 ();
 sg13g2_decap_4 FILLER_32_339 ();
 sg13g2_decap_8 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_2 ();
 sg13g2_fill_2 FILLER_33_34 ();
 sg13g2_fill_2 FILLER_33_62 ();
 sg13g2_fill_2 FILLER_33_91 ();
 sg13g2_fill_2 FILLER_33_114 ();
 sg13g2_fill_1 FILLER_33_141 ();
 sg13g2_fill_1 FILLER_33_160 ();
 sg13g2_fill_2 FILLER_33_192 ();
 sg13g2_decap_8 FILLER_33_202 ();
 sg13g2_decap_4 FILLER_33_209 ();
 sg13g2_fill_1 FILLER_33_221 ();
 sg13g2_fill_1 FILLER_33_227 ();
 sg13g2_decap_4 FILLER_33_231 ();
 sg13g2_fill_2 FILLER_33_235 ();
 sg13g2_decap_8 FILLER_33_240 ();
 sg13g2_decap_8 FILLER_33_247 ();
 sg13g2_decap_4 FILLER_33_254 ();
 sg13g2_fill_1 FILLER_33_263 ();
 sg13g2_decap_4 FILLER_33_319 ();
 sg13g2_decap_8 FILLER_33_379 ();
 sg13g2_decap_8 FILLER_33_386 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_fill_1 FILLER_34_74 ();
 sg13g2_fill_1 FILLER_34_80 ();
 sg13g2_fill_1 FILLER_34_94 ();
 sg13g2_fill_1 FILLER_34_116 ();
 sg13g2_fill_2 FILLER_34_122 ();
 sg13g2_fill_1 FILLER_34_124 ();
 sg13g2_fill_2 FILLER_34_135 ();
 sg13g2_fill_1 FILLER_34_137 ();
 sg13g2_fill_1 FILLER_34_155 ();
 sg13g2_fill_2 FILLER_34_175 ();
 sg13g2_fill_1 FILLER_34_227 ();
 sg13g2_decap_4 FILLER_34_253 ();
 sg13g2_fill_1 FILLER_34_257 ();
 sg13g2_fill_2 FILLER_34_297 ();
 sg13g2_fill_1 FILLER_34_304 ();
 sg13g2_fill_2 FILLER_34_309 ();
 sg13g2_decap_8 FILLER_34_347 ();
 sg13g2_decap_8 FILLER_34_354 ();
 sg13g2_fill_2 FILLER_34_361 ();
 sg13g2_fill_1 FILLER_34_363 ();
 sg13g2_fill_2 FILLER_34_367 ();
 sg13g2_fill_1 FILLER_34_369 ();
 sg13g2_decap_8 FILLER_34_386 ();
 sg13g2_decap_8 FILLER_34_393 ();
 sg13g2_decap_8 FILLER_34_400 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_fill_2 FILLER_35_39 ();
 sg13g2_fill_1 FILLER_35_68 ();
 sg13g2_fill_1 FILLER_35_125 ();
 sg13g2_fill_2 FILLER_35_196 ();
 sg13g2_fill_1 FILLER_35_207 ();
 sg13g2_decap_8 FILLER_35_256 ();
 sg13g2_fill_2 FILLER_35_263 ();
 sg13g2_fill_2 FILLER_35_290 ();
 sg13g2_decap_4 FILLER_35_306 ();
 sg13g2_fill_2 FILLER_35_310 ();
 sg13g2_fill_2 FILLER_35_317 ();
 sg13g2_fill_2 FILLER_35_335 ();
 sg13g2_fill_1 FILLER_35_337 ();
 sg13g2_decap_4 FILLER_35_405 ();
 sg13g2_fill_1 FILLER_36_37 ();
 sg13g2_fill_2 FILLER_36_94 ();
 sg13g2_fill_1 FILLER_36_96 ();
 sg13g2_fill_2 FILLER_36_159 ();
 sg13g2_fill_1 FILLER_36_189 ();
 sg13g2_fill_2 FILLER_36_216 ();
 sg13g2_fill_1 FILLER_36_286 ();
 sg13g2_fill_2 FILLER_36_337 ();
 sg13g2_fill_1 FILLER_36_339 ();
 sg13g2_fill_2 FILLER_36_346 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_49 ();
 sg13g2_fill_2 FILLER_37_145 ();
 sg13g2_fill_1 FILLER_37_147 ();
 sg13g2_fill_1 FILLER_37_202 ();
 sg13g2_fill_2 FILLER_37_208 ();
 sg13g2_fill_1 FILLER_37_243 ();
 sg13g2_decap_4 FILLER_37_259 ();
 sg13g2_fill_2 FILLER_37_263 ();
 sg13g2_fill_2 FILLER_37_282 ();
 sg13g2_fill_2 FILLER_37_315 ();
 sg13g2_decap_4 FILLER_37_351 ();
 sg13g2_fill_2 FILLER_37_355 ();
 sg13g2_fill_2 FILLER_38_70 ();
 sg13g2_fill_1 FILLER_38_72 ();
 sg13g2_fill_1 FILLER_38_97 ();
 sg13g2_fill_1 FILLER_38_108 ();
 sg13g2_fill_2 FILLER_38_127 ();
 sg13g2_fill_1 FILLER_38_129 ();
 sg13g2_fill_2 FILLER_38_135 ();
 sg13g2_fill_1 FILLER_38_137 ();
 sg13g2_fill_1 FILLER_38_157 ();
 sg13g2_fill_2 FILLER_38_177 ();
 sg13g2_fill_2 FILLER_38_218 ();
 sg13g2_fill_1 FILLER_38_243 ();
 sg13g2_fill_2 FILLER_38_253 ();
 sg13g2_decap_8 FILLER_38_268 ();
 sg13g2_decap_4 FILLER_38_275 ();
 sg13g2_fill_1 FILLER_38_279 ();
 sg13g2_fill_1 FILLER_38_336 ();
 sg13g2_decap_4 FILLER_38_363 ();
 sg13g2_fill_1 FILLER_38_399 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_2 ();
 sg13g2_fill_1 FILLER_39_108 ();
 sg13g2_fill_2 FILLER_39_182 ();
 sg13g2_fill_1 FILLER_39_293 ();
 sg13g2_fill_1 FILLER_39_309 ();
 sg13g2_fill_1 FILLER_39_313 ();
 sg13g2_decap_4 FILLER_39_364 ();
 sg13g2_fill_1 FILLER_39_395 ();
 sg13g2_decap_8 FILLER_39_399 ();
 sg13g2_fill_2 FILLER_39_406 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_2 ();
 sg13g2_fill_1 FILLER_40_59 ();
 sg13g2_fill_1 FILLER_40_74 ();
 sg13g2_fill_2 FILLER_40_101 ();
 sg13g2_fill_2 FILLER_40_138 ();
 sg13g2_fill_1 FILLER_40_149 ();
 sg13g2_decap_8 FILLER_40_159 ();
 sg13g2_decap_8 FILLER_40_170 ();
 sg13g2_fill_2 FILLER_40_177 ();
 sg13g2_fill_1 FILLER_40_179 ();
 sg13g2_fill_2 FILLER_40_193 ();
 sg13g2_fill_1 FILLER_40_195 ();
 sg13g2_fill_2 FILLER_40_255 ();
 sg13g2_decap_8 FILLER_40_299 ();
 sg13g2_decap_8 FILLER_40_306 ();
 sg13g2_fill_2 FILLER_40_313 ();
 sg13g2_fill_1 FILLER_40_337 ();
 sg13g2_decap_8 FILLER_40_360 ();
 sg13g2_decap_8 FILLER_40_367 ();
 sg13g2_decap_8 FILLER_40_374 ();
 sg13g2_decap_8 FILLER_40_381 ();
 sg13g2_decap_8 FILLER_40_388 ();
 sg13g2_decap_8 FILLER_40_395 ();
 sg13g2_decap_8 FILLER_40_402 ();
 sg13g2_fill_2 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_2 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_fill_2 FILLER_41_14 ();
 sg13g2_fill_1 FILLER_41_16 ();
 sg13g2_fill_2 FILLER_41_34 ();
 sg13g2_fill_2 FILLER_41_54 ();
 sg13g2_fill_2 FILLER_41_60 ();
 sg13g2_fill_1 FILLER_41_62 ();
 sg13g2_fill_2 FILLER_41_75 ();
 sg13g2_fill_2 FILLER_41_134 ();
 sg13g2_decap_4 FILLER_41_158 ();
 sg13g2_fill_1 FILLER_41_162 ();
 sg13g2_decap_4 FILLER_41_167 ();
 sg13g2_fill_1 FILLER_41_244 ();
 sg13g2_fill_1 FILLER_41_286 ();
 sg13g2_decap_8 FILLER_41_306 ();
 sg13g2_fill_1 FILLER_41_313 ();
 sg13g2_fill_2 FILLER_41_359 ();
 sg13g2_decap_4 FILLER_41_374 ();
 sg13g2_fill_1 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_41_383 ();
 sg13g2_decap_8 FILLER_41_390 ();
 sg13g2_decap_8 FILLER_41_397 ();
 sg13g2_decap_4 FILLER_41_404 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_fill_1 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_5 ();
 sg13g2_fill_1 FILLER_42_7 ();
 sg13g2_fill_2 FILLER_42_58 ();
 sg13g2_fill_1 FILLER_42_71 ();
 sg13g2_fill_1 FILLER_42_85 ();
 sg13g2_fill_2 FILLER_42_94 ();
 sg13g2_fill_1 FILLER_42_163 ();
 sg13g2_fill_1 FILLER_42_181 ();
 sg13g2_fill_2 FILLER_42_222 ();
 sg13g2_fill_2 FILLER_42_286 ();
 sg13g2_fill_2 FILLER_42_314 ();
 sg13g2_fill_1 FILLER_42_358 ();
 sg13g2_fill_1 FILLER_42_377 ();
 sg13g2_decap_8 FILLER_42_392 ();
 sg13g2_decap_8 FILLER_42_399 ();
 sg13g2_fill_2 FILLER_42_406 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_fill_2 FILLER_43_91 ();
 sg13g2_fill_1 FILLER_43_107 ();
 sg13g2_fill_1 FILLER_43_115 ();
 sg13g2_fill_2 FILLER_43_133 ();
 sg13g2_fill_1 FILLER_43_135 ();
 sg13g2_fill_1 FILLER_43_226 ();
 sg13g2_fill_1 FILLER_43_275 ();
 sg13g2_fill_2 FILLER_43_328 ();
 sg13g2_decap_8 FILLER_43_338 ();
 sg13g2_decap_4 FILLER_43_345 ();
 sg13g2_decap_8 FILLER_43_402 ();
 sg13g2_fill_2 FILLER_44_136 ();
 sg13g2_fill_1 FILLER_44_148 ();
 sg13g2_fill_2 FILLER_44_159 ();
 sg13g2_fill_1 FILLER_44_161 ();
 sg13g2_fill_1 FILLER_44_250 ();
 sg13g2_fill_2 FILLER_44_264 ();
 sg13g2_decap_8 FILLER_44_318 ();
 sg13g2_decap_8 FILLER_44_325 ();
 sg13g2_decap_8 FILLER_44_332 ();
 sg13g2_fill_1 FILLER_44_339 ();
 sg13g2_fill_2 FILLER_44_345 ();
 sg13g2_fill_1 FILLER_44_347 ();
 sg13g2_fill_1 FILLER_45_26 ();
 sg13g2_decap_4 FILLER_45_151 ();
 sg13g2_fill_2 FILLER_45_162 ();
 sg13g2_fill_1 FILLER_45_164 ();
 sg13g2_decap_8 FILLER_45_174 ();
 sg13g2_fill_1 FILLER_45_250 ();
 sg13g2_decap_8 FILLER_45_320 ();
 sg13g2_decap_4 FILLER_45_327 ();
 sg13g2_fill_1 FILLER_45_351 ();
 sg13g2_fill_1 FILLER_45_373 ();
 sg13g2_fill_1 FILLER_45_382 ();
 sg13g2_fill_1 FILLER_46_45 ();
 sg13g2_fill_1 FILLER_46_168 ();
 sg13g2_fill_1 FILLER_46_198 ();
 sg13g2_fill_2 FILLER_46_233 ();
 sg13g2_fill_2 FILLER_46_239 ();
 sg13g2_fill_1 FILLER_46_264 ();
 sg13g2_fill_2 FILLER_46_270 ();
 sg13g2_fill_2 FILLER_46_293 ();
 sg13g2_fill_1 FILLER_46_295 ();
 sg13g2_fill_2 FILLER_46_307 ();
 sg13g2_fill_1 FILLER_46_309 ();
 sg13g2_decap_4 FILLER_46_383 ();
 sg13g2_decap_8 FILLER_46_393 ();
 sg13g2_decap_8 FILLER_46_400 ();
 sg13g2_fill_2 FILLER_46_407 ();
 sg13g2_fill_1 FILLER_47_90 ();
 sg13g2_fill_2 FILLER_47_101 ();
 sg13g2_fill_2 FILLER_47_139 ();
 sg13g2_fill_1 FILLER_47_177 ();
 sg13g2_decap_4 FILLER_47_213 ();
 sg13g2_fill_2 FILLER_47_217 ();
 sg13g2_fill_2 FILLER_47_222 ();
 sg13g2_fill_1 FILLER_47_224 ();
 sg13g2_fill_2 FILLER_47_256 ();
 sg13g2_fill_2 FILLER_47_271 ();
 sg13g2_decap_4 FILLER_47_386 ();
 sg13g2_fill_1 FILLER_47_390 ();
 sg13g2_fill_1 FILLER_48_63 ();
 sg13g2_fill_2 FILLER_48_98 ();
 sg13g2_fill_1 FILLER_48_100 ();
 sg13g2_fill_2 FILLER_48_109 ();
 sg13g2_fill_1 FILLER_48_111 ();
 sg13g2_decap_4 FILLER_48_185 ();
 sg13g2_fill_1 FILLER_48_197 ();
 sg13g2_decap_8 FILLER_48_209 ();
 sg13g2_fill_2 FILLER_48_216 ();
 sg13g2_fill_2 FILLER_48_231 ();
 sg13g2_fill_1 FILLER_48_237 ();
 sg13g2_fill_2 FILLER_48_273 ();
 sg13g2_fill_2 FILLER_48_281 ();
 sg13g2_fill_1 FILLER_48_292 ();
 sg13g2_decap_4 FILLER_48_332 ();
 sg13g2_fill_1 FILLER_48_340 ();
 sg13g2_decap_4 FILLER_48_345 ();
 sg13g2_fill_1 FILLER_48_349 ();
 sg13g2_fill_2 FILLER_48_376 ();
 sg13g2_fill_1 FILLER_48_378 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_fill_1 FILLER_49_35 ();
 sg13g2_fill_1 FILLER_49_45 ();
 sg13g2_fill_2 FILLER_49_55 ();
 sg13g2_fill_2 FILLER_49_103 ();
 sg13g2_fill_2 FILLER_49_117 ();
 sg13g2_fill_1 FILLER_49_119 ();
 sg13g2_fill_2 FILLER_49_139 ();
 sg13g2_fill_1 FILLER_49_141 ();
 sg13g2_fill_1 FILLER_49_183 ();
 sg13g2_decap_4 FILLER_49_193 ();
 sg13g2_decap_8 FILLER_49_202 ();
 sg13g2_decap_4 FILLER_49_209 ();
 sg13g2_fill_1 FILLER_49_213 ();
 sg13g2_decap_4 FILLER_49_257 ();
 sg13g2_fill_2 FILLER_49_261 ();
 sg13g2_fill_2 FILLER_49_295 ();
 sg13g2_decap_8 FILLER_49_323 ();
 sg13g2_decap_8 FILLER_49_330 ();
 sg13g2_decap_8 FILLER_49_337 ();
 sg13g2_decap_8 FILLER_49_344 ();
 sg13g2_decap_8 FILLER_49_351 ();
 sg13g2_decap_4 FILLER_49_358 ();
 sg13g2_fill_1 FILLER_49_367 ();
 sg13g2_fill_2 FILLER_49_376 ();
 sg13g2_fill_1 FILLER_50_17 ();
 sg13g2_fill_2 FILLER_50_160 ();
 sg13g2_fill_1 FILLER_50_162 ();
 sg13g2_fill_2 FILLER_50_168 ();
 sg13g2_decap_8 FILLER_50_196 ();
 sg13g2_decap_4 FILLER_50_203 ();
 sg13g2_decap_4 FILLER_50_215 ();
 sg13g2_decap_8 FILLER_50_250 ();
 sg13g2_decap_4 FILLER_50_257 ();
 sg13g2_fill_2 FILLER_50_261 ();
 sg13g2_decap_4 FILLER_50_322 ();
 sg13g2_decap_4 FILLER_50_339 ();
 sg13g2_fill_1 FILLER_50_361 ();
 sg13g2_fill_2 FILLER_50_374 ();
 sg13g2_fill_1 FILLER_50_376 ();
 sg13g2_fill_2 FILLER_50_398 ();
 sg13g2_fill_2 FILLER_51_31 ();
 sg13g2_fill_1 FILLER_51_33 ();
 sg13g2_fill_2 FILLER_51_65 ();
 sg13g2_fill_1 FILLER_51_67 ();
 sg13g2_fill_1 FILLER_51_76 ();
 sg13g2_fill_2 FILLER_51_108 ();
 sg13g2_fill_1 FILLER_51_110 ();
 sg13g2_fill_2 FILLER_51_119 ();
 sg13g2_fill_2 FILLER_51_135 ();
 sg13g2_fill_1 FILLER_51_137 ();
 sg13g2_fill_2 FILLER_51_147 ();
 sg13g2_fill_1 FILLER_51_149 ();
 sg13g2_fill_2 FILLER_51_167 ();
 sg13g2_fill_1 FILLER_51_169 ();
 sg13g2_fill_1 FILLER_51_201 ();
 sg13g2_fill_2 FILLER_51_219 ();
 sg13g2_fill_1 FILLER_51_221 ();
 sg13g2_fill_2 FILLER_51_238 ();
 sg13g2_decap_8 FILLER_51_250 ();
 sg13g2_decap_8 FILLER_51_257 ();
 sg13g2_decap_8 FILLER_51_264 ();
 sg13g2_decap_8 FILLER_51_271 ();
 sg13g2_decap_8 FILLER_51_282 ();
 sg13g2_decap_4 FILLER_51_289 ();
 sg13g2_decap_4 FILLER_51_306 ();
 sg13g2_fill_1 FILLER_51_310 ();
 sg13g2_fill_2 FILLER_51_318 ();
 sg13g2_fill_1 FILLER_51_337 ();
 sg13g2_fill_1 FILLER_51_356 ();
 sg13g2_fill_2 FILLER_51_377 ();
 sg13g2_fill_1 FILLER_51_379 ();
 sg13g2_fill_1 FILLER_52_107 ();
 sg13g2_fill_1 FILLER_52_152 ();
 sg13g2_fill_1 FILLER_52_169 ();
 sg13g2_fill_2 FILLER_52_184 ();
 sg13g2_fill_2 FILLER_52_203 ();
 sg13g2_fill_1 FILLER_52_205 ();
 sg13g2_fill_2 FILLER_52_209 ();
 sg13g2_fill_1 FILLER_52_216 ();
 sg13g2_decap_8 FILLER_52_227 ();
 sg13g2_decap_4 FILLER_52_234 ();
 sg13g2_decap_4 FILLER_52_244 ();
 sg13g2_fill_2 FILLER_52_248 ();
 sg13g2_decap_8 FILLER_52_265 ();
 sg13g2_fill_2 FILLER_52_272 ();
 sg13g2_decap_8 FILLER_52_283 ();
 sg13g2_decap_4 FILLER_52_294 ();
 sg13g2_fill_1 FILLER_52_298 ();
 sg13g2_fill_1 FILLER_52_338 ();
 sg13g2_decap_4 FILLER_52_351 ();
 sg13g2_fill_1 FILLER_53_26 ();
 sg13g2_fill_2 FILLER_53_62 ();
 sg13g2_fill_2 FILLER_53_78 ();
 sg13g2_fill_1 FILLER_53_80 ();
 sg13g2_fill_1 FILLER_53_121 ();
 sg13g2_fill_2 FILLER_53_127 ();
 sg13g2_fill_1 FILLER_53_129 ();
 sg13g2_fill_2 FILLER_53_147 ();
 sg13g2_fill_1 FILLER_53_149 ();
 sg13g2_fill_1 FILLER_53_162 ();
 sg13g2_fill_1 FILLER_53_168 ();
 sg13g2_fill_2 FILLER_53_177 ();
 sg13g2_fill_1 FILLER_53_179 ();
 sg13g2_decap_8 FILLER_53_206 ();
 sg13g2_fill_1 FILLER_53_230 ();
 sg13g2_fill_1 FILLER_53_237 ();
 sg13g2_fill_2 FILLER_53_250 ();
 sg13g2_fill_1 FILLER_53_252 ();
 sg13g2_fill_1 FILLER_53_258 ();
 sg13g2_fill_2 FILLER_53_336 ();
 sg13g2_fill_1 FILLER_53_351 ();
 sg13g2_fill_2 FILLER_53_357 ();
 sg13g2_fill_1 FILLER_53_372 ();
 sg13g2_fill_2 FILLER_53_399 ();
 sg13g2_fill_2 FILLER_53_406 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_fill_2 FILLER_54_32 ();
 sg13g2_fill_2 FILLER_54_51 ();
 sg13g2_fill_2 FILLER_54_108 ();
 sg13g2_fill_2 FILLER_54_150 ();
 sg13g2_decap_4 FILLER_54_156 ();
 sg13g2_fill_1 FILLER_54_160 ();
 sg13g2_fill_1 FILLER_54_174 ();
 sg13g2_fill_2 FILLER_54_193 ();
 sg13g2_fill_1 FILLER_54_195 ();
 sg13g2_fill_2 FILLER_54_218 ();
 sg13g2_fill_2 FILLER_54_247 ();
 sg13g2_fill_1 FILLER_54_249 ();
 sg13g2_decap_4 FILLER_54_376 ();
 sg13g2_fill_2 FILLER_54_396 ();
 sg13g2_fill_1 FILLER_54_398 ();
 sg13g2_decap_4 FILLER_55_4 ();
 sg13g2_fill_2 FILLER_55_13 ();
 sg13g2_fill_1 FILLER_55_20 ();
 sg13g2_decap_4 FILLER_55_30 ();
 sg13g2_fill_1 FILLER_55_34 ();
 sg13g2_fill_1 FILLER_55_69 ();
 sg13g2_fill_2 FILLER_55_75 ();
 sg13g2_fill_2 FILLER_55_86 ();
 sg13g2_fill_2 FILLER_55_158 ();
 sg13g2_fill_1 FILLER_55_160 ();
 sg13g2_fill_2 FILLER_55_184 ();
 sg13g2_fill_2 FILLER_55_203 ();
 sg13g2_decap_8 FILLER_55_231 ();
 sg13g2_decap_8 FILLER_55_238 ();
 sg13g2_fill_2 FILLER_55_245 ();
 sg13g2_fill_1 FILLER_55_247 ();
 sg13g2_fill_2 FILLER_55_314 ();
 sg13g2_fill_1 FILLER_55_316 ();
 sg13g2_fill_2 FILLER_55_329 ();
 sg13g2_fill_1 FILLER_55_348 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_2 ();
 sg13g2_fill_2 FILLER_56_29 ();
 sg13g2_fill_1 FILLER_56_79 ();
 sg13g2_fill_1 FILLER_56_92 ();
 sg13g2_fill_2 FILLER_56_110 ();
 sg13g2_fill_1 FILLER_56_112 ();
 sg13g2_fill_2 FILLER_56_123 ();
 sg13g2_fill_1 FILLER_56_125 ();
 sg13g2_fill_2 FILLER_56_171 ();
 sg13g2_fill_1 FILLER_56_173 ();
 sg13g2_fill_2 FILLER_56_214 ();
 sg13g2_fill_1 FILLER_56_216 ();
 sg13g2_decap_8 FILLER_56_226 ();
 sg13g2_fill_2 FILLER_56_233 ();
 sg13g2_fill_1 FILLER_56_235 ();
 sg13g2_decap_8 FILLER_56_298 ();
 sg13g2_decap_4 FILLER_56_305 ();
 sg13g2_fill_1 FILLER_56_309 ();
 sg13g2_decap_4 FILLER_56_314 ();
 sg13g2_fill_1 FILLER_56_318 ();
 sg13g2_decap_4 FILLER_56_327 ();
 sg13g2_decap_8 FILLER_56_342 ();
 sg13g2_decap_8 FILLER_56_349 ();
 sg13g2_fill_2 FILLER_56_356 ();
 sg13g2_decap_8 FILLER_56_376 ();
 sg13g2_decap_4 FILLER_56_383 ();
 sg13g2_fill_1 FILLER_56_387 ();
 sg13g2_fill_2 FILLER_57_85 ();
 sg13g2_fill_1 FILLER_57_87 ();
 sg13g2_fill_2 FILLER_57_97 ();
 sg13g2_fill_2 FILLER_57_107 ();
 sg13g2_fill_1 FILLER_57_138 ();
 sg13g2_fill_2 FILLER_57_182 ();
 sg13g2_fill_2 FILLER_57_210 ();
 sg13g2_fill_1 FILLER_57_212 ();
 sg13g2_fill_2 FILLER_57_235 ();
 sg13g2_fill_1 FILLER_57_304 ();
 sg13g2_decap_8 FILLER_57_314 ();
 sg13g2_decap_8 FILLER_57_321 ();
 sg13g2_decap_8 FILLER_57_328 ();
 sg13g2_fill_2 FILLER_57_344 ();
 sg13g2_decap_8 FILLER_57_355 ();
 sg13g2_fill_2 FILLER_57_362 ();
 sg13g2_fill_1 FILLER_57_364 ();
 sg13g2_fill_2 FILLER_57_374 ();
 sg13g2_fill_2 FILLER_57_402 ();
 sg13g2_fill_2 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_2 ();
 sg13g2_fill_2 FILLER_58_20 ();
 sg13g2_fill_1 FILLER_58_37 ();
 sg13g2_fill_2 FILLER_58_43 ();
 sg13g2_fill_2 FILLER_58_100 ();
 sg13g2_fill_1 FILLER_58_102 ();
 sg13g2_fill_1 FILLER_58_117 ();
 sg13g2_fill_2 FILLER_58_177 ();
 sg13g2_fill_2 FILLER_58_193 ();
 sg13g2_fill_2 FILLER_58_209 ();
 sg13g2_fill_2 FILLER_58_238 ();
 sg13g2_fill_2 FILLER_58_258 ();
 sg13g2_fill_2 FILLER_58_277 ();
 sg13g2_fill_1 FILLER_58_279 ();
 sg13g2_decap_8 FILLER_58_294 ();
 sg13g2_decap_4 FILLER_58_301 ();
 sg13g2_fill_1 FILLER_58_305 ();
 sg13g2_decap_8 FILLER_58_310 ();
 sg13g2_fill_2 FILLER_58_317 ();
 sg13g2_fill_1 FILLER_58_319 ();
 sg13g2_fill_1 FILLER_58_359 ();
 sg13g2_fill_1 FILLER_58_368 ();
 sg13g2_fill_2 FILLER_58_382 ();
 sg13g2_fill_1 FILLER_58_384 ();
 sg13g2_fill_2 FILLER_58_407 ();
 sg13g2_fill_2 FILLER_59_26 ();
 sg13g2_fill_2 FILLER_59_37 ();
 sg13g2_fill_2 FILLER_59_58 ();
 sg13g2_fill_2 FILLER_59_78 ();
 sg13g2_fill_1 FILLER_59_210 ();
 sg13g2_fill_1 FILLER_59_235 ();
 sg13g2_fill_2 FILLER_59_246 ();
 sg13g2_decap_4 FILLER_59_274 ();
 sg13g2_decap_8 FILLER_59_282 ();
 sg13g2_decap_8 FILLER_59_289 ();
 sg13g2_fill_2 FILLER_59_316 ();
 sg13g2_fill_1 FILLER_59_326 ();
 sg13g2_fill_1 FILLER_59_372 ();
 sg13g2_fill_2 FILLER_59_407 ();
 sg13g2_fill_2 FILLER_60_51 ();
 sg13g2_fill_1 FILLER_60_95 ();
 sg13g2_decap_4 FILLER_60_132 ();
 sg13g2_fill_1 FILLER_60_146 ();
 sg13g2_fill_2 FILLER_60_164 ();
 sg13g2_fill_1 FILLER_60_166 ();
 sg13g2_fill_1 FILLER_60_175 ();
 sg13g2_fill_1 FILLER_60_182 ();
 sg13g2_fill_2 FILLER_60_192 ();
 sg13g2_fill_1 FILLER_60_194 ();
 sg13g2_fill_2 FILLER_60_208 ();
 sg13g2_decap_8 FILLER_60_227 ();
 sg13g2_fill_2 FILLER_60_234 ();
 sg13g2_decap_4 FILLER_60_239 ();
 sg13g2_fill_1 FILLER_60_279 ();
 sg13g2_fill_2 FILLER_60_293 ();
 sg13g2_fill_1 FILLER_60_295 ();
 sg13g2_decap_4 FILLER_60_314 ();
 sg13g2_fill_2 FILLER_60_340 ();
 sg13g2_fill_1 FILLER_60_342 ();
 sg13g2_decap_4 FILLER_60_376 ();
 sg13g2_fill_1 FILLER_60_380 ();
 sg13g2_decap_8 FILLER_60_398 ();
 sg13g2_fill_1 FILLER_60_405 ();
 sg13g2_fill_2 FILLER_61_35 ();
 sg13g2_fill_1 FILLER_61_45 ();
 sg13g2_fill_2 FILLER_61_56 ();
 sg13g2_fill_2 FILLER_61_67 ();
 sg13g2_fill_2 FILLER_61_141 ();
 sg13g2_fill_2 FILLER_61_147 ();
 sg13g2_fill_1 FILLER_61_149 ();
 sg13g2_fill_2 FILLER_61_163 ();
 sg13g2_fill_2 FILLER_61_169 ();
 sg13g2_fill_1 FILLER_61_171 ();
 sg13g2_fill_2 FILLER_61_177 ();
 sg13g2_decap_8 FILLER_61_184 ();
 sg13g2_decap_8 FILLER_61_191 ();
 sg13g2_decap_8 FILLER_61_198 ();
 sg13g2_decap_4 FILLER_61_205 ();
 sg13g2_decap_8 FILLER_61_212 ();
 sg13g2_fill_2 FILLER_61_227 ();
 sg13g2_fill_1 FILLER_61_229 ();
 sg13g2_decap_8 FILLER_61_235 ();
 sg13g2_decap_8 FILLER_61_242 ();
 sg13g2_fill_2 FILLER_61_266 ();
 sg13g2_fill_1 FILLER_61_268 ();
 sg13g2_fill_2 FILLER_61_295 ();
 sg13g2_fill_1 FILLER_61_340 ();
 sg13g2_fill_2 FILLER_61_364 ();
 sg13g2_fill_1 FILLER_61_366 ();
 sg13g2_decap_4 FILLER_61_403 ();
 sg13g2_fill_2 FILLER_61_407 ();
 sg13g2_fill_1 FILLER_62_61 ();
 sg13g2_fill_2 FILLER_62_67 ();
 sg13g2_fill_2 FILLER_62_74 ();
 sg13g2_fill_1 FILLER_62_107 ();
 sg13g2_fill_2 FILLER_62_208 ();
 sg13g2_fill_1 FILLER_62_210 ();
 sg13g2_decap_8 FILLER_62_216 ();
 sg13g2_fill_2 FILLER_62_243 ();
 sg13g2_fill_2 FILLER_62_258 ();
 sg13g2_fill_1 FILLER_62_260 ();
 sg13g2_decap_8 FILLER_62_300 ();
 sg13g2_decap_8 FILLER_62_307 ();
 sg13g2_decap_4 FILLER_62_314 ();
 sg13g2_fill_1 FILLER_62_318 ();
 sg13g2_fill_1 FILLER_62_324 ();
 sg13g2_fill_2 FILLER_62_337 ();
 sg13g2_decap_8 FILLER_62_351 ();
 sg13g2_decap_8 FILLER_62_358 ();
 sg13g2_fill_1 FILLER_62_365 ();
 sg13g2_decap_8 FILLER_62_397 ();
 sg13g2_decap_4 FILLER_62_404 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_83 ();
 sg13g2_fill_2 FILLER_63_90 ();
 sg13g2_fill_1 FILLER_63_92 ();
 sg13g2_fill_1 FILLER_63_98 ();
 sg13g2_fill_2 FILLER_63_108 ();
 sg13g2_fill_1 FILLER_63_110 ();
 sg13g2_fill_1 FILLER_63_129 ();
 sg13g2_fill_1 FILLER_63_216 ();
 sg13g2_fill_1 FILLER_63_239 ();
 sg13g2_fill_2 FILLER_63_295 ();
 sg13g2_fill_1 FILLER_63_301 ();
 sg13g2_decap_8 FILLER_63_306 ();
 sg13g2_decap_4 FILLER_63_313 ();
 sg13g2_fill_1 FILLER_63_317 ();
 sg13g2_decap_8 FILLER_63_326 ();
 sg13g2_decap_8 FILLER_63_333 ();
 sg13g2_decap_8 FILLER_63_340 ();
 sg13g2_decap_8 FILLER_63_347 ();
 sg13g2_fill_2 FILLER_63_354 ();
 sg13g2_fill_1 FILLER_63_356 ();
 sg13g2_fill_1 FILLER_63_370 ();
 sg13g2_decap_8 FILLER_63_389 ();
 sg13g2_decap_8 FILLER_63_396 ();
 sg13g2_decap_4 FILLER_63_403 ();
 sg13g2_fill_2 FILLER_63_407 ();
 sg13g2_fill_2 FILLER_64_9 ();
 sg13g2_fill_2 FILLER_64_43 ();
 sg13g2_fill_1 FILLER_64_45 ();
 sg13g2_fill_2 FILLER_64_88 ();
 sg13g2_fill_1 FILLER_64_96 ();
 sg13g2_fill_1 FILLER_64_103 ();
 sg13g2_fill_2 FILLER_64_161 ();
 sg13g2_fill_2 FILLER_64_179 ();
 sg13g2_fill_1 FILLER_64_181 ();
 sg13g2_fill_2 FILLER_64_191 ();
 sg13g2_decap_8 FILLER_64_233 ();
 sg13g2_decap_8 FILLER_64_240 ();
 sg13g2_fill_1 FILLER_64_296 ();
 sg13g2_fill_1 FILLER_64_310 ();
 sg13g2_fill_2 FILLER_64_319 ();
 sg13g2_decap_4 FILLER_64_342 ();
 sg13g2_fill_2 FILLER_64_354 ();
 sg13g2_decap_8 FILLER_64_390 ();
 sg13g2_decap_8 FILLER_64_397 ();
 sg13g2_decap_4 FILLER_64_404 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_2 ();
 sg13g2_fill_1 FILLER_65_56 ();
 sg13g2_fill_2 FILLER_65_66 ();
 sg13g2_fill_1 FILLER_65_68 ();
 sg13g2_decap_4 FILLER_65_90 ();
 sg13g2_fill_2 FILLER_65_172 ();
 sg13g2_fill_1 FILLER_65_233 ();
 sg13g2_fill_2 FILLER_65_253 ();
 sg13g2_fill_1 FILLER_65_255 ();
 sg13g2_fill_1 FILLER_65_264 ();
 sg13g2_decap_4 FILLER_65_284 ();
 sg13g2_fill_2 FILLER_65_297 ();
 sg13g2_fill_1 FILLER_65_299 ();
 sg13g2_fill_1 FILLER_65_358 ();
 sg13g2_decap_8 FILLER_65_378 ();
 sg13g2_decap_8 FILLER_65_394 ();
 sg13g2_decap_8 FILLER_65_401 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_fill_1 FILLER_66_34 ();
 sg13g2_fill_1 FILLER_66_83 ();
 sg13g2_fill_1 FILLER_66_115 ();
 sg13g2_fill_1 FILLER_66_169 ();
 sg13g2_fill_1 FILLER_66_175 ();
 sg13g2_decap_8 FILLER_66_225 ();
 sg13g2_decap_4 FILLER_66_232 ();
 sg13g2_fill_1 FILLER_66_236 ();
 sg13g2_decap_8 FILLER_66_256 ();
 sg13g2_decap_8 FILLER_66_263 ();
 sg13g2_fill_1 FILLER_66_285 ();
 sg13g2_decap_8 FILLER_66_386 ();
 sg13g2_decap_8 FILLER_66_393 ();
 sg13g2_decap_8 FILLER_66_400 ();
 sg13g2_fill_2 FILLER_66_407 ();
 sg13g2_fill_1 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_21 ();
 sg13g2_fill_2 FILLER_67_83 ();
 sg13g2_fill_2 FILLER_67_92 ();
 sg13g2_fill_1 FILLER_67_94 ();
 sg13g2_fill_2 FILLER_67_104 ();
 sg13g2_fill_1 FILLER_67_127 ();
 sg13g2_fill_1 FILLER_67_136 ();
 sg13g2_fill_2 FILLER_67_173 ();
 sg13g2_decap_4 FILLER_67_205 ();
 sg13g2_fill_1 FILLER_67_217 ();
 sg13g2_decap_8 FILLER_67_224 ();
 sg13g2_decap_4 FILLER_67_231 ();
 sg13g2_fill_2 FILLER_67_246 ();
 sg13g2_fill_1 FILLER_67_248 ();
 sg13g2_fill_2 FILLER_67_258 ();
 sg13g2_decap_4 FILLER_67_284 ();
 sg13g2_fill_1 FILLER_67_328 ();
 sg13g2_decap_8 FILLER_67_384 ();
 sg13g2_decap_8 FILLER_67_391 ();
 sg13g2_decap_8 FILLER_67_398 ();
 sg13g2_decap_4 FILLER_67_405 ();
 sg13g2_fill_2 FILLER_68_102 ();
 sg13g2_fill_1 FILLER_68_104 ();
 sg13g2_decap_8 FILLER_68_113 ();
 sg13g2_fill_1 FILLER_68_120 ();
 sg13g2_decap_4 FILLER_68_137 ();
 sg13g2_fill_2 FILLER_68_198 ();
 sg13g2_fill_1 FILLER_68_200 ();
 sg13g2_fill_2 FILLER_68_281 ();
 sg13g2_fill_2 FILLER_68_323 ();
 sg13g2_fill_2 FILLER_68_341 ();
 sg13g2_fill_2 FILLER_68_355 ();
 sg13g2_fill_1 FILLER_68_357 ();
 sg13g2_decap_8 FILLER_68_384 ();
 sg13g2_decap_8 FILLER_68_391 ();
 sg13g2_decap_8 FILLER_68_398 ();
 sg13g2_decap_4 FILLER_68_405 ();
 sg13g2_fill_1 FILLER_69_97 ();
 sg13g2_decap_4 FILLER_69_134 ();
 sg13g2_decap_8 FILLER_69_142 ();
 sg13g2_decap_4 FILLER_69_149 ();
 sg13g2_fill_1 FILLER_69_153 ();
 sg13g2_decap_8 FILLER_69_172 ();
 sg13g2_fill_2 FILLER_69_179 ();
 sg13g2_fill_2 FILLER_69_224 ();
 sg13g2_fill_1 FILLER_69_226 ();
 sg13g2_fill_2 FILLER_69_279 ();
 sg13g2_fill_2 FILLER_69_294 ();
 sg13g2_decap_8 FILLER_69_306 ();
 sg13g2_decap_8 FILLER_69_313 ();
 sg13g2_decap_8 FILLER_69_323 ();
 sg13g2_fill_1 FILLER_69_352 ();
 sg13g2_fill_2 FILLER_69_369 ();
 sg13g2_fill_1 FILLER_69_371 ();
 sg13g2_decap_8 FILLER_69_377 ();
 sg13g2_decap_8 FILLER_69_384 ();
 sg13g2_decap_8 FILLER_69_391 ();
 sg13g2_decap_8 FILLER_69_398 ();
 sg13g2_decap_4 FILLER_69_405 ();
 sg13g2_fill_1 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_20 ();
 sg13g2_fill_1 FILLER_70_22 ();
 sg13g2_fill_2 FILLER_70_55 ();
 sg13g2_fill_2 FILLER_70_65 ();
 sg13g2_fill_2 FILLER_70_125 ();
 sg13g2_fill_1 FILLER_70_127 ();
 sg13g2_decap_8 FILLER_70_182 ();
 sg13g2_fill_2 FILLER_70_243 ();
 sg13g2_fill_2 FILLER_70_262 ();
 sg13g2_fill_1 FILLER_70_264 ();
 sg13g2_fill_1 FILLER_70_282 ();
 sg13g2_decap_4 FILLER_70_288 ();
 sg13g2_fill_1 FILLER_70_292 ();
 sg13g2_decap_8 FILLER_70_302 ();
 sg13g2_decap_4 FILLER_70_309 ();
 sg13g2_fill_1 FILLER_70_313 ();
 sg13g2_fill_2 FILLER_70_368 ();
 sg13g2_fill_1 FILLER_70_370 ();
 sg13g2_fill_1 FILLER_70_379 ();
 sg13g2_decap_8 FILLER_70_385 ();
 sg13g2_decap_8 FILLER_70_392 ();
 sg13g2_decap_8 FILLER_70_399 ();
 sg13g2_fill_2 FILLER_70_406 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_23 ();
 sg13g2_fill_1 FILLER_71_25 ();
 sg13g2_fill_1 FILLER_71_31 ();
 sg13g2_fill_2 FILLER_71_45 ();
 sg13g2_fill_2 FILLER_71_73 ();
 sg13g2_decap_8 FILLER_71_129 ();
 sg13g2_decap_8 FILLER_71_194 ();
 sg13g2_fill_2 FILLER_71_201 ();
 sg13g2_fill_2 FILLER_71_221 ();
 sg13g2_fill_2 FILLER_71_227 ();
 sg13g2_fill_1 FILLER_71_229 ();
 sg13g2_decap_8 FILLER_71_250 ();
 sg13g2_decap_4 FILLER_71_257 ();
 sg13g2_fill_2 FILLER_71_261 ();
 sg13g2_fill_2 FILLER_71_273 ();
 sg13g2_fill_1 FILLER_71_275 ();
 sg13g2_fill_1 FILLER_71_295 ();
 sg13g2_fill_2 FILLER_71_349 ();
 sg13g2_decap_8 FILLER_71_396 ();
 sg13g2_decap_4 FILLER_71_403 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_fill_1 FILLER_72_35 ();
 sg13g2_fill_2 FILLER_72_48 ();
 sg13g2_fill_2 FILLER_72_85 ();
 sg13g2_fill_2 FILLER_72_124 ();
 sg13g2_fill_1 FILLER_72_126 ();
 sg13g2_fill_1 FILLER_72_214 ();
 sg13g2_fill_1 FILLER_72_234 ();
 sg13g2_fill_1 FILLER_72_290 ();
 sg13g2_decap_4 FILLER_72_301 ();
 sg13g2_decap_8 FILLER_72_395 ();
 sg13g2_decap_8 FILLER_72_402 ();
 sg13g2_fill_2 FILLER_73_0 ();
 sg13g2_fill_1 FILLER_73_2 ();
 sg13g2_fill_2 FILLER_73_17 ();
 sg13g2_fill_1 FILLER_73_19 ();
 sg13g2_fill_2 FILLER_73_44 ();
 sg13g2_fill_2 FILLER_73_64 ();
 sg13g2_fill_2 FILLER_73_117 ();
 sg13g2_fill_1 FILLER_73_163 ();
 sg13g2_fill_1 FILLER_73_235 ();
 sg13g2_fill_1 FILLER_73_271 ();
 sg13g2_fill_1 FILLER_73_294 ();
 sg13g2_decap_8 FILLER_73_384 ();
 sg13g2_decap_8 FILLER_73_391 ();
 sg13g2_decap_8 FILLER_73_398 ();
 sg13g2_decap_4 FILLER_73_405 ();
 sg13g2_fill_2 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_57 ();
 sg13g2_fill_1 FILLER_74_134 ();
 sg13g2_fill_2 FILLER_74_168 ();
 sg13g2_fill_1 FILLER_74_179 ();
 sg13g2_fill_1 FILLER_74_201 ();
 sg13g2_fill_2 FILLER_74_228 ();
 sg13g2_fill_1 FILLER_74_230 ();
 sg13g2_fill_1 FILLER_74_250 ();
 sg13g2_fill_1 FILLER_74_260 ();
 sg13g2_fill_1 FILLER_74_270 ();
 sg13g2_decap_4 FILLER_74_281 ();
 sg13g2_fill_1 FILLER_74_285 ();
 sg13g2_fill_2 FILLER_74_290 ();
 sg13g2_decap_8 FILLER_74_296 ();
 sg13g2_fill_1 FILLER_74_303 ();
 sg13g2_fill_2 FILLER_74_330 ();
 sg13g2_fill_1 FILLER_74_358 ();
 sg13g2_decap_8 FILLER_74_382 ();
 sg13g2_decap_8 FILLER_74_389 ();
 sg13g2_decap_8 FILLER_74_396 ();
 sg13g2_decap_4 FILLER_74_403 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_fill_1 FILLER_75_26 ();
 sg13g2_fill_1 FILLER_75_41 ();
 sg13g2_fill_1 FILLER_75_68 ();
 sg13g2_fill_1 FILLER_75_145 ();
 sg13g2_fill_2 FILLER_75_177 ();
 sg13g2_fill_1 FILLER_75_179 ();
 sg13g2_fill_2 FILLER_75_216 ();
 sg13g2_fill_1 FILLER_75_218 ();
 sg13g2_fill_2 FILLER_75_229 ();
 sg13g2_fill_1 FILLER_75_231 ();
 sg13g2_fill_1 FILLER_75_262 ();
 sg13g2_decap_4 FILLER_75_276 ();
 sg13g2_decap_4 FILLER_75_284 ();
 sg13g2_fill_2 FILLER_75_293 ();
 sg13g2_fill_1 FILLER_75_295 ();
 sg13g2_fill_1 FILLER_75_316 ();
 sg13g2_fill_2 FILLER_75_339 ();
 sg13g2_decap_4 FILLER_75_349 ();
 sg13g2_fill_1 FILLER_75_353 ();
 sg13g2_fill_2 FILLER_75_365 ();
 sg13g2_fill_1 FILLER_75_367 ();
 sg13g2_fill_2 FILLER_75_382 ();
 sg13g2_decap_8 FILLER_75_387 ();
 sg13g2_decap_8 FILLER_75_394 ();
 sg13g2_decap_8 FILLER_75_401 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_fill_1 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_122 ();
 sg13g2_decap_8 FILLER_76_197 ();
 sg13g2_decap_8 FILLER_76_204 ();
 sg13g2_decap_4 FILLER_76_211 ();
 sg13g2_fill_1 FILLER_76_215 ();
 sg13g2_decap_4 FILLER_76_225 ();
 sg13g2_fill_2 FILLER_76_255 ();
 sg13g2_fill_1 FILLER_76_257 ();
 sg13g2_fill_2 FILLER_76_279 ();
 sg13g2_fill_1 FILLER_76_281 ();
 sg13g2_fill_1 FILLER_76_301 ();
 sg13g2_decap_8 FILLER_76_320 ();
 sg13g2_decap_4 FILLER_76_327 ();
 sg13g2_fill_1 FILLER_76_331 ();
 sg13g2_decap_8 FILLER_76_336 ();
 sg13g2_decap_8 FILLER_76_343 ();
 sg13g2_decap_8 FILLER_76_350 ();
 sg13g2_fill_2 FILLER_76_357 ();
 sg13g2_decap_4 FILLER_76_404 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_fill_2 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_41 ();
 sg13g2_fill_2 FILLER_77_57 ();
 sg13g2_fill_1 FILLER_77_59 ();
 sg13g2_fill_1 FILLER_77_70 ();
 sg13g2_fill_2 FILLER_77_84 ();
 sg13g2_fill_1 FILLER_77_86 ();
 sg13g2_fill_2 FILLER_77_91 ();
 sg13g2_fill_2 FILLER_77_130 ();
 sg13g2_fill_2 FILLER_77_137 ();
 sg13g2_fill_1 FILLER_77_143 ();
 sg13g2_decap_8 FILLER_77_208 ();
 sg13g2_decap_8 FILLER_77_215 ();
 sg13g2_fill_2 FILLER_77_222 ();
 sg13g2_fill_2 FILLER_77_238 ();
 sg13g2_fill_2 FILLER_77_258 ();
 sg13g2_fill_2 FILLER_77_269 ();
 sg13g2_fill_2 FILLER_77_296 ();
 sg13g2_fill_2 FILLER_77_306 ();
 sg13g2_fill_1 FILLER_77_308 ();
 sg13g2_fill_2 FILLER_77_341 ();
 sg13g2_fill_1 FILLER_77_343 ();
 sg13g2_fill_2 FILLER_77_350 ();
 sg13g2_fill_1 FILLER_77_357 ();
 sg13g2_fill_2 FILLER_77_363 ();
 sg13g2_fill_1 FILLER_77_365 ();
 sg13g2_decap_4 FILLER_77_403 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_4 FILLER_78_7 ();
 sg13g2_decap_4 FILLER_78_15 ();
 sg13g2_fill_1 FILLER_78_19 ();
 sg13g2_fill_2 FILLER_78_33 ();
 sg13g2_fill_2 FILLER_78_183 ();
 sg13g2_fill_1 FILLER_78_237 ();
 sg13g2_decap_8 FILLER_78_250 ();
 sg13g2_fill_1 FILLER_78_260 ();
 sg13g2_decap_4 FILLER_78_296 ();
 sg13g2_fill_2 FILLER_78_326 ();
 sg13g2_fill_1 FILLER_78_328 ();
 sg13g2_decap_4 FILLER_78_355 ();
 sg13g2_decap_4 FILLER_78_403 ();
 sg13g2_fill_2 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_fill_1 FILLER_79_21 ();
 sg13g2_fill_1 FILLER_79_76 ();
 sg13g2_fill_1 FILLER_79_129 ();
 sg13g2_decap_8 FILLER_79_243 ();
 sg13g2_decap_8 FILLER_79_250 ();
 sg13g2_decap_8 FILLER_79_257 ();
 sg13g2_decap_4 FILLER_79_264 ();
 sg13g2_fill_1 FILLER_79_268 ();
 sg13g2_fill_1 FILLER_79_278 ();
 sg13g2_fill_2 FILLER_79_303 ();
 sg13g2_decap_4 FILLER_79_350 ();
 sg13g2_decap_8 FILLER_79_387 ();
 sg13g2_decap_8 FILLER_79_394 ();
 sg13g2_decap_8 FILLER_79_401 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_fill_2 FILLER_80_28 ();
 sg13g2_fill_2 FILLER_80_91 ();
 sg13g2_fill_1 FILLER_80_111 ();
 sg13g2_fill_2 FILLER_80_151 ();
 sg13g2_fill_2 FILLER_80_166 ();
 sg13g2_fill_1 FILLER_80_168 ();
 sg13g2_fill_2 FILLER_80_191 ();
 sg13g2_fill_1 FILLER_80_193 ();
 sg13g2_decap_8 FILLER_80_207 ();
 sg13g2_decap_4 FILLER_80_214 ();
 sg13g2_fill_1 FILLER_80_218 ();
 sg13g2_decap_8 FILLER_80_227 ();
 sg13g2_decap_8 FILLER_80_234 ();
 sg13g2_decap_8 FILLER_80_241 ();
 sg13g2_decap_8 FILLER_80_248 ();
 sg13g2_decap_8 FILLER_80_255 ();
 sg13g2_decap_8 FILLER_80_262 ();
 sg13g2_decap_4 FILLER_80_269 ();
 sg13g2_fill_1 FILLER_80_273 ();
 sg13g2_fill_2 FILLER_80_279 ();
 sg13g2_fill_1 FILLER_80_294 ();
 sg13g2_fill_2 FILLER_80_325 ();
 sg13g2_decap_8 FILLER_80_392 ();
 sg13g2_decap_8 FILLER_80_399 ();
 sg13g2_fill_2 FILLER_80_406 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net186;
 assign uio_oe[1] = net187;
 assign uio_oe[2] = net188;
 assign uio_oe[3] = net189;
 assign uio_oe[4] = net190;
 assign uio_oe[5] = net191;
 assign uio_oe[6] = net192;
 assign uio_oe[7] = net193;
endmodule

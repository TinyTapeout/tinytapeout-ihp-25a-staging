module tt_um_led_matrix_ayla_lin (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire clknet_0_clk;
 wire \top_inst.address[0] ;
 wire \top_inst.address[1] ;
 wire \top_inst.address[2] ;
 wire \top_inst.address[3] ;
 wire \top_inst.address[4] ;
 wire \top_inst.address[5] ;
 wire \top_inst.address[6] ;
 wire \top_inst.clk ;
 wire \top_inst.controller_inst.counter[0] ;
 wire \top_inst.controller_inst.counter[10] ;
 wire \top_inst.controller_inst.counter[11] ;
 wire \top_inst.controller_inst.counter[12] ;
 wire \top_inst.controller_inst.counter[13] ;
 wire \top_inst.controller_inst.counter[14] ;
 wire \top_inst.controller_inst.counter[15] ;
 wire \top_inst.controller_inst.counter[16] ;
 wire \top_inst.controller_inst.counter[17] ;
 wire \top_inst.controller_inst.counter[18] ;
 wire \top_inst.controller_inst.counter[19] ;
 wire \top_inst.controller_inst.counter[1] ;
 wire \top_inst.controller_inst.counter[20] ;
 wire \top_inst.controller_inst.counter[21] ;
 wire \top_inst.controller_inst.counter[2] ;
 wire \top_inst.controller_inst.counter[3] ;
 wire \top_inst.controller_inst.counter[4] ;
 wire \top_inst.controller_inst.counter[5] ;
 wire \top_inst.controller_inst.counter[6] ;
 wire \top_inst.controller_inst.counter[7] ;
 wire \top_inst.controller_inst.counter[8] ;
 wire \top_inst.controller_inst.counter[9] ;
 wire \top_inst.controller_inst.spi_load ;
 wire \top_inst.controller_inst.spi_load_next ;
 wire \top_inst.controller_inst.spi_load_pending ;
 wire \top_inst.controller_inst.spi_ready ;
 wire \top_inst.controller_inst.state[0] ;
 wire \top_inst.controller_inst.state[1] ;
 wire \top_inst.controller_inst.state[2] ;
 wire \top_inst.controller_inst.state[3] ;
 wire \top_inst.counter[0] ;
 wire \top_inst.counter[1] ;
 wire \top_inst.counter[2] ;
 wire \top_inst.counter[3] ;
 wire \top_inst.data[0] ;
 wire \top_inst.data[10] ;
 wire \top_inst.data[11] ;
 wire \top_inst.data[12] ;
 wire \top_inst.data[13] ;
 wire \top_inst.data[14] ;
 wire \top_inst.data[15] ;
 wire \top_inst.data[16] ;
 wire \top_inst.data[17] ;
 wire \top_inst.data[18] ;
 wire \top_inst.data[19] ;
 wire \top_inst.data[1] ;
 wire \top_inst.data[20] ;
 wire \top_inst.data[21] ;
 wire \top_inst.data[24] ;
 wire \top_inst.data[25] ;
 wire \top_inst.data[26] ;
 wire \top_inst.data[27] ;
 wire \top_inst.data[28] ;
 wire \top_inst.data[29] ;
 wire \top_inst.data[2] ;
 wire \top_inst.data[30] ;
 wire \top_inst.data[31] ;
 wire \top_inst.data[36] ;
 wire \top_inst.data[37] ;
 wire \top_inst.data[39] ;
 wire \top_inst.data[40] ;
 wire \top_inst.data[41] ;
 wire \top_inst.data[42] ;
 wire \top_inst.data[4] ;
 wire \top_inst.data[5] ;
 wire \top_inst.data[6] ;
 wire \top_inst.data[7] ;
 wire \top_inst.spi_cs_n ;
 wire \top_inst.spi_inst.buffer[0] ;
 wire \top_inst.spi_inst.buffer[10] ;
 wire \top_inst.spi_inst.buffer[11] ;
 wire \top_inst.spi_inst.buffer[12] ;
 wire \top_inst.spi_inst.buffer[13] ;
 wire \top_inst.spi_inst.buffer[14] ;
 wire \top_inst.spi_inst.buffer[15] ;
 wire \top_inst.spi_inst.buffer[16] ;
 wire \top_inst.spi_inst.buffer[17] ;
 wire \top_inst.spi_inst.buffer[18] ;
 wire \top_inst.spi_inst.buffer[19] ;
 wire \top_inst.spi_inst.buffer[1] ;
 wire \top_inst.spi_inst.buffer[20] ;
 wire \top_inst.spi_inst.buffer[21] ;
 wire \top_inst.spi_inst.buffer[22] ;
 wire \top_inst.spi_inst.buffer[23] ;
 wire \top_inst.spi_inst.buffer[24] ;
 wire \top_inst.spi_inst.buffer[25] ;
 wire \top_inst.spi_inst.buffer[26] ;
 wire \top_inst.spi_inst.buffer[27] ;
 wire \top_inst.spi_inst.buffer[28] ;
 wire \top_inst.spi_inst.buffer[29] ;
 wire \top_inst.spi_inst.buffer[2] ;
 wire \top_inst.spi_inst.buffer[30] ;
 wire \top_inst.spi_inst.buffer[31] ;
 wire \top_inst.spi_inst.buffer[32] ;
 wire \top_inst.spi_inst.buffer[33] ;
 wire \top_inst.spi_inst.buffer[34] ;
 wire \top_inst.spi_inst.buffer[35] ;
 wire \top_inst.spi_inst.buffer[36] ;
 wire \top_inst.spi_inst.buffer[37] ;
 wire \top_inst.spi_inst.buffer[38] ;
 wire \top_inst.spi_inst.buffer[39] ;
 wire \top_inst.spi_inst.buffer[3] ;
 wire \top_inst.spi_inst.buffer[40] ;
 wire \top_inst.spi_inst.buffer[41] ;
 wire \top_inst.spi_inst.buffer[42] ;
 wire \top_inst.spi_inst.buffer[43] ;
 wire \top_inst.spi_inst.buffer[44] ;
 wire \top_inst.spi_inst.buffer[45] ;
 wire \top_inst.spi_inst.buffer[46] ;
 wire \top_inst.spi_inst.buffer[47] ;
 wire \top_inst.spi_inst.buffer[48] ;
 wire \top_inst.spi_inst.buffer[49] ;
 wire \top_inst.spi_inst.buffer[4] ;
 wire \top_inst.spi_inst.buffer[50] ;
 wire \top_inst.spi_inst.buffer[51] ;
 wire \top_inst.spi_inst.buffer[52] ;
 wire \top_inst.spi_inst.buffer[53] ;
 wire \top_inst.spi_inst.buffer[54] ;
 wire \top_inst.spi_inst.buffer[55] ;
 wire \top_inst.spi_inst.buffer[56] ;
 wire \top_inst.spi_inst.buffer[57] ;
 wire \top_inst.spi_inst.buffer[58] ;
 wire \top_inst.spi_inst.buffer[59] ;
 wire \top_inst.spi_inst.buffer[5] ;
 wire \top_inst.spi_inst.buffer[60] ;
 wire \top_inst.spi_inst.buffer[61] ;
 wire \top_inst.spi_inst.buffer[62] ;
 wire \top_inst.spi_inst.buffer[63] ;
 wire \top_inst.spi_inst.buffer[6] ;
 wire \top_inst.spi_inst.buffer[7] ;
 wire \top_inst.spi_inst.buffer[8] ;
 wire \top_inst.spi_inst.buffer[9] ;
 wire \top_inst.spi_inst.counter[0] ;
 wire \top_inst.spi_inst.counter[1] ;
 wire \top_inst.spi_inst.counter[2] ;
 wire \top_inst.spi_inst.counter[3] ;
 wire \top_inst.spi_inst.counter[4] ;
 wire \top_inst.spi_inst.counter[5] ;
 wire \top_inst.spi_inst.counter[6] ;
 wire \top_inst.spi_inst.state[1] ;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net1;
 wire net2;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;

 sg13g2_inv_1 _0750_ (.Y(_0148_),
    .A(\top_inst.controller_inst.counter[15] ));
 sg13g2_inv_1 _0751_ (.Y(_0149_),
    .A(\top_inst.controller_inst.counter[6] ));
 sg13g2_inv_1 _0752_ (.Y(_0150_),
    .A(\top_inst.controller_inst.counter[5] ));
 sg13g2_inv_1 _0753_ (.Y(_0151_),
    .A(\top_inst.controller_inst.counter[4] ));
 sg13g2_inv_4 _0754_ (.A(\top_inst.address[0] ),
    .Y(_0152_));
 sg13g2_inv_1 _0755_ (.Y(_0153_),
    .A(\top_inst.address[2] ));
 sg13g2_inv_2 _0756_ (.Y(_0154_),
    .A(\top_inst.address[3] ));
 sg13g2_inv_1 _0757_ (.Y(_0155_),
    .A(\top_inst.address[4] ));
 sg13g2_inv_1 _0758_ (.Y(_0156_),
    .A(\top_inst.data[12] ));
 sg13g2_inv_1 _0759_ (.Y(_0157_),
    .A(\top_inst.data[13] ));
 sg13g2_inv_1 _0760_ (.Y(_0158_),
    .A(\top_inst.data[14] ));
 sg13g2_inv_1 _0761_ (.Y(_0159_),
    .A(\top_inst.data[15] ));
 sg13g2_inv_1 _0762_ (.Y(_0160_),
    .A(\top_inst.data[16] ));
 sg13g2_inv_1 _0763_ (.Y(_0161_),
    .A(\top_inst.data[17] ));
 sg13g2_inv_1 _0764_ (.Y(_0162_),
    .A(\top_inst.data[18] ));
 sg13g2_inv_1 _0765_ (.Y(_0163_),
    .A(\top_inst.data[19] ));
 sg13g2_inv_1 _0766_ (.Y(_0164_),
    .A(\top_inst.data[36] ));
 sg13g2_inv_1 _0767_ (.Y(_0165_),
    .A(\top_inst.data[39] ));
 sg13g2_inv_1 _0768_ (.Y(_0166_),
    .A(\top_inst.data[40] ));
 sg13g2_inv_1 _0769_ (.Y(_0167_),
    .A(\top_inst.data[41] ));
 sg13g2_inv_1 _0770_ (.Y(_0168_),
    .A(\top_inst.data[42] ));
 sg13g2_inv_1 _0771_ (.Y(_0169_),
    .A(\top_inst.data[24] ));
 sg13g2_inv_1 _0772_ (.Y(_0170_),
    .A(\top_inst.data[25] ));
 sg13g2_inv_1 _0773_ (.Y(_0171_),
    .A(\top_inst.data[26] ));
 sg13g2_inv_1 _0774_ (.Y(_0172_),
    .A(\top_inst.data[27] ));
 sg13g2_inv_1 _0775_ (.Y(_0173_),
    .A(\top_inst.data[28] ));
 sg13g2_inv_1 _0776_ (.Y(_0174_),
    .A(\top_inst.data[29] ));
 sg13g2_inv_1 _0777_ (.Y(_0175_),
    .A(\top_inst.data[30] ));
 sg13g2_inv_1 _0778_ (.Y(_0176_),
    .A(\top_inst.data[31] ));
 sg13g2_inv_1 _0779_ (.Y(_0177_),
    .A(\top_inst.data[1] ));
 sg13g2_inv_1 _0780_ (.Y(_0178_),
    .A(\top_inst.data[4] ));
 sg13g2_inv_1 _0781_ (.Y(_0179_),
    .A(\top_inst.data[5] ));
 sg13g2_inv_1 _0782_ (.Y(_0180_),
    .A(\top_inst.data[6] ));
 sg13g2_inv_1 _0783_ (.Y(_0181_),
    .A(\top_inst.data[7] ));
 sg13g2_inv_1 _0784_ (.Y(_0182_),
    .A(net244));
 sg13g2_nand4_1 _0785_ (.B(\top_inst.controller_inst.counter[2] ),
    .C(\top_inst.controller_inst.counter[1] ),
    .A(\top_inst.controller_inst.counter[3] ),
    .Y(_0183_),
    .D(\top_inst.controller_inst.counter[0] ));
 sg13g2_nor3_2 _0786_ (.A(_0150_),
    .B(_0151_),
    .C(_0183_),
    .Y(_0184_));
 sg13g2_or2_1 _0787_ (.X(_0185_),
    .B(_0184_),
    .A(\top_inst.controller_inst.counter[6] ));
 sg13g2_nor3_1 _0788_ (.A(\top_inst.controller_inst.counter[12] ),
    .B(\top_inst.controller_inst.counter[11] ),
    .C(\top_inst.controller_inst.counter[8] ),
    .Y(_0186_));
 sg13g2_nor4_1 _0789_ (.A(\top_inst.controller_inst.counter[13] ),
    .B(\top_inst.controller_inst.counter[10] ),
    .C(\top_inst.controller_inst.counter[9] ),
    .D(\top_inst.controller_inst.counter[7] ),
    .Y(_0187_));
 sg13g2_or4_1 _0790_ (.A(\top_inst.controller_inst.counter[17] ),
    .B(\top_inst.controller_inst.counter[16] ),
    .C(\top_inst.controller_inst.counter[15] ),
    .D(\top_inst.controller_inst.counter[14] ),
    .X(_0188_));
 sg13g2_nor4_1 _0791_ (.A(\top_inst.controller_inst.counter[21] ),
    .B(\top_inst.controller_inst.counter[20] ),
    .C(\top_inst.controller_inst.counter[19] ),
    .D(\top_inst.controller_inst.counter[18] ),
    .Y(_0189_));
 sg13g2_nand3_1 _0792_ (.B(_0187_),
    .C(_0189_),
    .A(_0186_),
    .Y(_0190_));
 sg13g2_nor4_2 _0793_ (.A(\top_inst.controller_inst.counter[6] ),
    .B(_0184_),
    .C(_0188_),
    .Y(_0191_),
    .D(_0190_));
 sg13g2_nand2b_1 _0794_ (.Y(_0192_),
    .B(net219),
    .A_N(\top_inst.controller_inst.spi_load_next ));
 sg13g2_or2_1 _0795_ (.X(_0193_),
    .B(_0192_),
    .A(_0191_));
 sg13g2_and2_2 _0796_ (.A(\top_inst.address[0] ),
    .B(net220),
    .X(_0194_));
 sg13g2_nand2_2 _0797_ (.Y(_0195_),
    .A(\top_inst.address[0] ),
    .B(net220));
 sg13g2_nor3_2 _0798_ (.A(\top_inst.address[4] ),
    .B(\top_inst.address[5] ),
    .C(\top_inst.address[6] ),
    .Y(_0196_));
 sg13g2_or3_1 _0799_ (.A(\top_inst.address[4] ),
    .B(\top_inst.address[5] ),
    .C(\top_inst.address[6] ),
    .X(_0197_));
 sg13g2_nand3_1 _0800_ (.B(\top_inst.address[3] ),
    .C(_0196_),
    .A(_0153_),
    .Y(_0198_));
 sg13g2_or2_1 _0801_ (.X(_0199_),
    .B(_0198_),
    .A(_0195_));
 sg13g2_nor2_1 _0802_ (.A(\top_inst.address[2] ),
    .B(\top_inst.address[3] ),
    .Y(_0200_));
 sg13g2_or2_1 _0803_ (.X(_0201_),
    .B(\top_inst.address[3] ),
    .A(\top_inst.address[2] ));
 sg13g2_nor4_2 _0804_ (.A(_0155_),
    .B(\top_inst.address[5] ),
    .C(\top_inst.address[6] ),
    .Y(_0202_),
    .D(_0201_));
 sg13g2_nand2_1 _0805_ (.Y(_0203_),
    .A(_0194_),
    .B(_0202_));
 sg13g2_a21oi_1 _0806_ (.A1(_0199_),
    .A2(_0203_),
    .Y(_0204_),
    .B1(_0193_));
 sg13g2_and2_1 _0807_ (.A(net1),
    .B(net247),
    .X(_0205_));
 sg13g2_nand2_2 _0808_ (.Y(_0206_),
    .A(net1),
    .B(net247));
 sg13g2_and2_1 _0809_ (.A(\top_inst.controller_inst.state[1] ),
    .B(net246),
    .X(_0207_));
 sg13g2_nand2_1 _0810_ (.Y(_0208_),
    .A(\top_inst.controller_inst.state[1] ),
    .B(net246));
 sg13g2_and2_2 _0811_ (.A(_0196_),
    .B(_0200_),
    .X(_0209_));
 sg13g2_nand2_1 _0812_ (.Y(_0210_),
    .A(_0196_),
    .B(_0200_));
 sg13g2_nor3_1 _0813_ (.A(_0193_),
    .B(_0195_),
    .C(_0210_),
    .Y(_0211_));
 sg13g2_nand2_1 _0814_ (.Y(_0212_),
    .A(\top_inst.controller_inst.state[2] ),
    .B(net246));
 sg13g2_nor4_1 _0815_ (.A(_0193_),
    .B(_0195_),
    .C(_0210_),
    .D(_0212_),
    .Y(_0213_));
 sg13g2_and2_1 _0816_ (.A(\top_inst.controller_inst.state[3] ),
    .B(_0205_),
    .X(_0214_));
 sg13g2_nor4_2 _0817_ (.A(_0149_),
    .B(_0150_),
    .C(_0151_),
    .Y(_0215_),
    .D(_0183_));
 sg13g2_nand2_1 _0818_ (.Y(_0216_),
    .A(\top_inst.controller_inst.counter[6] ),
    .B(_0184_));
 sg13g2_and2_1 _0819_ (.A(\top_inst.controller_inst.counter[10] ),
    .B(\top_inst.controller_inst.counter[9] ),
    .X(_0217_));
 sg13g2_and3_1 _0820_ (.X(_0218_),
    .A(\top_inst.controller_inst.counter[11] ),
    .B(\top_inst.controller_inst.counter[8] ),
    .C(_0217_));
 sg13g2_nand3_1 _0821_ (.B(_0215_),
    .C(_0218_),
    .A(\top_inst.controller_inst.counter[7] ),
    .Y(_0219_));
 sg13g2_nand3_1 _0822_ (.B(\top_inst.controller_inst.counter[13] ),
    .C(\top_inst.controller_inst.counter[12] ),
    .A(\top_inst.controller_inst.counter[14] ),
    .Y(_0220_));
 sg13g2_nor2_1 _0823_ (.A(_0148_),
    .B(_0220_),
    .Y(_0221_));
 sg13g2_nand4_1 _0824_ (.B(_0215_),
    .C(_0218_),
    .A(\top_inst.controller_inst.counter[7] ),
    .Y(_0222_),
    .D(_0221_));
 sg13g2_nand4_1 _0825_ (.B(\top_inst.controller_inst.counter[18] ),
    .C(\top_inst.controller_inst.counter[17] ),
    .A(\top_inst.controller_inst.counter[19] ),
    .Y(_0223_),
    .D(\top_inst.controller_inst.counter[16] ));
 sg13g2_nor2_2 _0826_ (.A(_0222_),
    .B(_0223_),
    .Y(_0224_));
 sg13g2_nand3_1 _0827_ (.B(\top_inst.controller_inst.counter[20] ),
    .C(_0224_),
    .A(\top_inst.controller_inst.counter[21] ),
    .Y(_0225_));
 sg13g2_nand4_1 _0828_ (.B(\top_inst.controller_inst.counter[20] ),
    .C(_0214_),
    .A(\top_inst.controller_inst.counter[21] ),
    .Y(_0226_),
    .D(_0224_));
 sg13g2_o21ai_1 _0829_ (.B1(_0226_),
    .Y(_0227_),
    .A1(_0204_),
    .A2(_0208_));
 sg13g2_or2_1 _0830_ (.X(_0001_),
    .B(_0227_),
    .A(_0213_));
 sg13g2_and2_1 _0831_ (.A(\top_inst.spi_inst.counter[0] ),
    .B(\top_inst.spi_inst.counter[1] ),
    .X(_0228_));
 sg13g2_and2_1 _0832_ (.A(\top_inst.spi_inst.counter[2] ),
    .B(_0228_),
    .X(_0229_));
 sg13g2_and3_1 _0833_ (.X(_0230_),
    .A(\top_inst.spi_inst.counter[3] ),
    .B(\top_inst.spi_inst.counter[2] ),
    .C(_0228_));
 sg13g2_and2_1 _0834_ (.A(\top_inst.spi_inst.counter[4] ),
    .B(_0230_),
    .X(_0231_));
 sg13g2_nand2_1 _0835_ (.Y(_0232_),
    .A(\top_inst.spi_inst.counter[5] ),
    .B(_0231_));
 sg13g2_nor2_1 _0836_ (.A(\top_inst.spi_inst.counter[6] ),
    .B(_0232_),
    .Y(_0233_));
 sg13g2_nand2_1 _0837_ (.Y(_0234_),
    .A(net213),
    .B(_0233_));
 sg13g2_nor2b_1 _0838_ (.A(\top_inst.controller_inst.spi_load ),
    .B_N(net217),
    .Y(_0235_));
 sg13g2_nand2b_1 _0839_ (.Y(_0236_),
    .B(net217),
    .A_N(\top_inst.controller_inst.spi_load ));
 sg13g2_nand3_1 _0840_ (.B(_0234_),
    .C(net211),
    .A(net248),
    .Y(_0004_));
 sg13g2_and3_1 _0841_ (.X(_0237_),
    .A(net217),
    .B(net247),
    .C(\top_inst.controller_inst.spi_load ));
 sg13g2_inv_1 _0842_ (.Y(_0238_),
    .A(_0237_));
 sg13g2_nand2_2 _0843_ (.Y(_0239_),
    .A(net248),
    .B(net216));
 sg13g2_o21ai_1 _0844_ (.B1(_0238_),
    .Y(_0005_),
    .A1(_0233_),
    .A2(_0239_));
 sg13g2_a22oi_1 _0845_ (.Y(_0240_),
    .B1(_0214_),
    .B2(_0225_),
    .A2(_0207_),
    .A1(_0204_));
 sg13g2_inv_1 _0846_ (.Y(_0003_),
    .A(_0240_));
 sg13g2_nor2b_2 _0847_ (.A(net219),
    .B_N(\top_inst.controller_inst.state[0] ),
    .Y(_0241_));
 sg13g2_nand2b_2 _0848_ (.Y(_0242_),
    .B(\top_inst.controller_inst.state[0] ),
    .A_N(net219));
 sg13g2_nand2_1 _0849_ (.Y(_0000_),
    .A(_0205_),
    .B(_0242_));
 sg13g2_nand2_1 _0850_ (.Y(_0243_),
    .A(net219),
    .B(net246));
 sg13g2_nand3_1 _0851_ (.B(\top_inst.controller_inst.state[0] ),
    .C(net246),
    .A(net219),
    .Y(_0244_));
 sg13g2_o21ai_1 _0852_ (.B1(_0244_),
    .Y(_0002_),
    .A1(_0211_),
    .A2(_0212_));
 sg13g2_nor2_2 _0853_ (.A(\top_inst.controller_inst.state[2] ),
    .B(\top_inst.controller_inst.state[1] ),
    .Y(_0245_));
 sg13g2_inv_1 _0854_ (.Y(_0246_),
    .A(_0245_));
 sg13g2_o21ai_1 _0855_ (.B1(_0246_),
    .Y(_0247_),
    .A1(_0191_),
    .A2(_0192_));
 sg13g2_nor2_1 _0856_ (.A(\top_inst.controller_inst.state[0] ),
    .B(_0246_),
    .Y(_0248_));
 sg13g2_nor2_1 _0857_ (.A(_0243_),
    .B(_0248_),
    .Y(_0249_));
 sg13g2_and2_2 _0858_ (.A(_0247_),
    .B(_0249_),
    .X(_0250_));
 sg13g2_nor3_2 _0859_ (.A(_0193_),
    .B(_0243_),
    .C(_0245_),
    .Y(_0009_));
 sg13g2_nor2_2 _0860_ (.A(\top_inst.address[0] ),
    .B(net220),
    .Y(_0251_));
 sg13g2_nor2_1 _0861_ (.A(_0194_),
    .B(_0251_),
    .Y(_0252_));
 sg13g2_or2_1 _0862_ (.X(_0253_),
    .B(_0251_),
    .A(_0194_));
 sg13g2_nand2_1 _0863_ (.Y(_0254_),
    .A(_0202_),
    .B(_0252_));
 sg13g2_nand4_1 _0864_ (.B(\top_inst.address[3] ),
    .C(_0196_),
    .A(\top_inst.address[2] ),
    .Y(_0255_),
    .D(_0252_));
 sg13g2_and2_1 _0865_ (.A(_0254_),
    .B(_0255_),
    .X(_0256_));
 sg13g2_nand2_1 _0866_ (.Y(_0048_),
    .A(_0198_),
    .B(_0256_));
 sg13g2_nor3_2 _0867_ (.A(_0153_),
    .B(\top_inst.address[3] ),
    .C(_0197_),
    .Y(_0257_));
 sg13g2_nand2_1 _0868_ (.Y(_0258_),
    .A(\top_inst.address[1] ),
    .B(_0257_));
 sg13g2_nand2_1 _0869_ (.Y(_0259_),
    .A(_0194_),
    .B(_0257_));
 sg13g2_nand3_1 _0870_ (.B(_0256_),
    .C(_0259_),
    .A(_0198_),
    .Y(_0010_));
 sg13g2_and2_1 _0871_ (.A(net250),
    .B(net170),
    .X(_0011_));
 sg13g2_o21ai_1 _0872_ (.B1(net250),
    .Y(_0260_),
    .A1(net174),
    .A2(\top_inst.counter[1] ));
 sg13g2_a21oi_1 _0873_ (.A1(net174),
    .A2(\top_inst.counter[1] ),
    .Y(_0012_),
    .B1(_0260_));
 sg13g2_a21oi_1 _0874_ (.A1(\top_inst.counter[0] ),
    .A2(\top_inst.counter[1] ),
    .Y(_0261_),
    .B1(net171));
 sg13g2_nand3_1 _0875_ (.B(net178),
    .C(net171),
    .A(net174),
    .Y(_0262_));
 sg13g2_nand2_1 _0876_ (.Y(_0263_),
    .A(net250),
    .B(_0262_));
 sg13g2_nor2_1 _0877_ (.A(net172),
    .B(_0263_),
    .Y(_0013_));
 sg13g2_nand2b_1 _0878_ (.Y(_0264_),
    .B(_0262_),
    .A_N(net176));
 sg13g2_nand4_1 _0879_ (.B(\top_inst.counter[1] ),
    .C(net171),
    .A(net174),
    .Y(_0265_),
    .D(net176));
 sg13g2_and3_1 _0880_ (.X(_0014_),
    .A(net250),
    .B(_0264_),
    .C(net177));
 sg13g2_o21ai_1 _0881_ (.B1(net250),
    .Y(_0266_),
    .A1(_0182_),
    .A2(net177));
 sg13g2_a21oi_1 _0882_ (.A1(_0182_),
    .A2(net177),
    .Y(_0015_),
    .B1(_0266_));
 sg13g2_nand2b_1 _0883_ (.Y(_0267_),
    .B(_0247_),
    .A_N(\top_inst.controller_inst.state[3] ));
 sg13g2_a21oi_1 _0884_ (.A1(_0006_),
    .A2(_0248_),
    .Y(_0268_),
    .B1(_0241_));
 sg13g2_a21oi_1 _0885_ (.A1(_0267_),
    .A2(_0268_),
    .Y(_0269_),
    .B1(\top_inst.controller_inst.counter[0] ));
 sg13g2_and2_1 _0886_ (.A(\top_inst.controller_inst.counter[0] ),
    .B(_0242_),
    .X(_0270_));
 sg13g2_nor3_1 _0887_ (.A(_0206_),
    .B(_0269_),
    .C(_0270_),
    .Y(_0016_));
 sg13g2_nand3_1 _0888_ (.B(_0242_),
    .C(_0247_),
    .A(_0006_),
    .Y(_0271_));
 sg13g2_nand2_1 _0889_ (.Y(_0272_),
    .A(net246),
    .B(_0271_));
 sg13g2_nor2_1 _0890_ (.A(\top_inst.controller_inst.counter[1] ),
    .B(_0270_),
    .Y(_0273_));
 sg13g2_and2_1 _0891_ (.A(\top_inst.controller_inst.counter[1] ),
    .B(_0270_),
    .X(_0274_));
 sg13g2_nor3_1 _0892_ (.A(net190),
    .B(_0273_),
    .C(_0274_),
    .Y(_0017_));
 sg13g2_xnor2_1 _0893_ (.Y(_0275_),
    .A(\top_inst.controller_inst.counter[2] ),
    .B(_0274_));
 sg13g2_nor2_1 _0894_ (.A(net190),
    .B(_0275_),
    .Y(_0018_));
 sg13g2_a21oi_1 _0895_ (.A1(\top_inst.controller_inst.counter[2] ),
    .A2(_0274_),
    .Y(_0276_),
    .B1(\top_inst.controller_inst.counter[3] ));
 sg13g2_nor2_1 _0896_ (.A(_0183_),
    .B(_0241_),
    .Y(_0277_));
 sg13g2_a21oi_1 _0897_ (.A1(_0006_),
    .A2(_0247_),
    .Y(_0278_),
    .B1(_0241_));
 sg13g2_nor3_1 _0898_ (.A(net190),
    .B(_0276_),
    .C(_0277_),
    .Y(_0019_));
 sg13g2_xnor2_1 _0899_ (.Y(_0279_),
    .A(\top_inst.controller_inst.counter[4] ),
    .B(_0277_));
 sg13g2_nor2_1 _0900_ (.A(_0272_),
    .B(_0279_),
    .Y(_0020_));
 sg13g2_a21oi_1 _0901_ (.A1(\top_inst.controller_inst.counter[4] ),
    .A2(_0277_),
    .Y(_0280_),
    .B1(\top_inst.controller_inst.counter[5] ));
 sg13g2_nor4_1 _0902_ (.A(_0150_),
    .B(_0151_),
    .C(_0183_),
    .D(_0241_),
    .Y(_0281_));
 sg13g2_nor3_1 _0903_ (.A(net190),
    .B(_0280_),
    .C(_0281_),
    .Y(_0021_));
 sg13g2_o21ai_1 _0904_ (.B1(\top_inst.controller_inst.state[0] ),
    .Y(_0282_),
    .A1(\top_inst.controller_inst.counter[6] ),
    .A2(net219));
 sg13g2_nand4_1 _0905_ (.B(_0216_),
    .C(_0267_),
    .A(_0185_),
    .Y(_0283_),
    .D(_0268_));
 sg13g2_a21oi_1 _0906_ (.A1(_0282_),
    .A2(_0283_),
    .Y(_0022_),
    .B1(_0206_));
 sg13g2_a21oi_1 _0907_ (.A1(_0215_),
    .A2(_0242_),
    .Y(_0284_),
    .B1(\top_inst.controller_inst.counter[7] ));
 sg13g2_and3_2 _0908_ (.X(_0285_),
    .A(\top_inst.controller_inst.counter[7] ),
    .B(_0215_),
    .C(_0242_));
 sg13g2_nor3_1 _0909_ (.A(net190),
    .B(_0284_),
    .C(_0285_),
    .Y(_0023_));
 sg13g2_xnor2_1 _0910_ (.Y(_0286_),
    .A(\top_inst.controller_inst.counter[8] ),
    .B(_0285_));
 sg13g2_nor2_1 _0911_ (.A(net190),
    .B(_0286_),
    .Y(_0024_));
 sg13g2_and3_1 _0912_ (.X(_0287_),
    .A(\top_inst.controller_inst.counter[9] ),
    .B(\top_inst.controller_inst.counter[8] ),
    .C(_0285_));
 sg13g2_a21oi_1 _0913_ (.A1(\top_inst.controller_inst.counter[8] ),
    .A2(_0285_),
    .Y(_0288_),
    .B1(\top_inst.controller_inst.counter[9] ));
 sg13g2_nor3_1 _0914_ (.A(net190),
    .B(_0287_),
    .C(_0288_),
    .Y(_0025_));
 sg13g2_nand3_1 _0915_ (.B(_0217_),
    .C(_0285_),
    .A(\top_inst.controller_inst.counter[8] ),
    .Y(_0289_));
 sg13g2_nand4_1 _0916_ (.B(\top_inst.controller_inst.counter[7] ),
    .C(_0215_),
    .A(\top_inst.controller_inst.counter[8] ),
    .Y(_0290_),
    .D(_0217_));
 sg13g2_o21ai_1 _0917_ (.B1(_0289_),
    .Y(_0291_),
    .A1(\top_inst.controller_inst.counter[10] ),
    .A2(_0287_));
 sg13g2_nor2_1 _0918_ (.A(net189),
    .B(_0291_),
    .Y(_0026_));
 sg13g2_nand2_1 _0919_ (.Y(_0292_),
    .A(\top_inst.controller_inst.counter[11] ),
    .B(_0241_));
 sg13g2_nand2b_1 _0920_ (.Y(_0293_),
    .B(_0290_),
    .A_N(\top_inst.controller_inst.counter[11] ));
 sg13g2_nand3_1 _0921_ (.B(_0278_),
    .C(_0293_),
    .A(_0219_),
    .Y(_0294_));
 sg13g2_a21oi_1 _0922_ (.A1(_0292_),
    .A2(_0294_),
    .Y(_0027_),
    .B1(_0206_));
 sg13g2_and2_1 _0923_ (.A(_0218_),
    .B(_0285_),
    .X(_0295_));
 sg13g2_nor2_1 _0924_ (.A(\top_inst.controller_inst.counter[12] ),
    .B(_0295_),
    .Y(_0296_));
 sg13g2_and2_1 _0925_ (.A(\top_inst.controller_inst.counter[12] ),
    .B(_0295_),
    .X(_0297_));
 sg13g2_nor3_1 _0926_ (.A(net189),
    .B(_0296_),
    .C(_0297_),
    .Y(_0028_));
 sg13g2_nor2_1 _0927_ (.A(\top_inst.controller_inst.counter[13] ),
    .B(_0297_),
    .Y(_0298_));
 sg13g2_and2_1 _0928_ (.A(\top_inst.controller_inst.counter[13] ),
    .B(_0297_),
    .X(_0299_));
 sg13g2_nor3_1 _0929_ (.A(net189),
    .B(_0298_),
    .C(_0299_),
    .Y(_0029_));
 sg13g2_a21oi_1 _0930_ (.A1(\top_inst.controller_inst.counter[13] ),
    .A2(_0297_),
    .Y(_0300_),
    .B1(\top_inst.controller_inst.counter[14] ));
 sg13g2_nor3_1 _0931_ (.A(_0219_),
    .B(_0220_),
    .C(_0241_),
    .Y(_0301_));
 sg13g2_nor3_1 _0932_ (.A(net189),
    .B(_0300_),
    .C(_0301_),
    .Y(_0030_));
 sg13g2_nand2_1 _0933_ (.Y(_0302_),
    .A(\top_inst.controller_inst.counter[15] ),
    .B(_0241_));
 sg13g2_o21ai_1 _0934_ (.B1(_0148_),
    .Y(_0303_),
    .A1(_0219_),
    .A2(_0220_));
 sg13g2_nand3_1 _0935_ (.B(_0278_),
    .C(_0303_),
    .A(_0222_),
    .Y(_0304_));
 sg13g2_a21oi_1 _0936_ (.A1(_0302_),
    .A2(_0304_),
    .Y(_0031_),
    .B1(_0206_));
 sg13g2_nor2_2 _0937_ (.A(_0222_),
    .B(_0241_),
    .Y(_0305_));
 sg13g2_xnor2_1 _0938_ (.Y(_0306_),
    .A(\top_inst.controller_inst.counter[16] ),
    .B(_0305_));
 sg13g2_nor2_1 _0939_ (.A(net189),
    .B(_0306_),
    .Y(_0032_));
 sg13g2_a21o_1 _0940_ (.A2(_0305_),
    .A1(\top_inst.controller_inst.counter[16] ),
    .B1(\top_inst.controller_inst.counter[17] ),
    .X(_0307_));
 sg13g2_nand3_1 _0941_ (.B(\top_inst.controller_inst.counter[16] ),
    .C(_0305_),
    .A(\top_inst.controller_inst.counter[17] ),
    .Y(_0308_));
 sg13g2_and4_1 _0942_ (.A(net246),
    .B(_0271_),
    .C(_0307_),
    .D(_0308_),
    .X(_0033_));
 sg13g2_nor2b_1 _0943_ (.A(\top_inst.controller_inst.counter[18] ),
    .B_N(_0308_),
    .Y(_0309_));
 sg13g2_and4_1 _0944_ (.A(\top_inst.controller_inst.counter[18] ),
    .B(\top_inst.controller_inst.counter[17] ),
    .C(\top_inst.controller_inst.counter[16] ),
    .D(_0305_),
    .X(_0310_));
 sg13g2_nor3_1 _0945_ (.A(net189),
    .B(_0309_),
    .C(_0310_),
    .Y(_0034_));
 sg13g2_nor2_1 _0946_ (.A(\top_inst.controller_inst.counter[19] ),
    .B(_0310_),
    .Y(_0311_));
 sg13g2_and2_1 _0947_ (.A(\top_inst.controller_inst.counter[19] ),
    .B(_0310_),
    .X(_0312_));
 sg13g2_nor3_1 _0948_ (.A(net189),
    .B(_0311_),
    .C(_0312_),
    .Y(_0035_));
 sg13g2_a21o_1 _0949_ (.A2(_0242_),
    .A1(_0224_),
    .B1(\top_inst.controller_inst.counter[20] ),
    .X(_0313_));
 sg13g2_nand3_1 _0950_ (.B(_0224_),
    .C(_0242_),
    .A(\top_inst.controller_inst.counter[20] ),
    .Y(_0314_));
 sg13g2_and4_1 _0951_ (.A(net246),
    .B(_0271_),
    .C(_0313_),
    .D(_0314_),
    .X(_0036_));
 sg13g2_xor2_1 _0952_ (.B(_0314_),
    .A(\top_inst.controller_inst.counter[21] ),
    .X(_0315_));
 sg13g2_nor2_1 _0953_ (.A(net189),
    .B(_0315_),
    .Y(_0037_));
 sg13g2_nand2_2 _0954_ (.Y(_0316_),
    .A(\top_inst.address[2] ),
    .B(_0194_));
 sg13g2_nor3_2 _0955_ (.A(_0154_),
    .B(_0155_),
    .C(_0316_),
    .Y(_0317_));
 sg13g2_inv_1 _0956_ (.Y(_0318_),
    .A(_0317_));
 sg13g2_and3_1 _0957_ (.X(_0319_),
    .A(\top_inst.address[5] ),
    .B(_0250_),
    .C(_0317_));
 sg13g2_nand4_1 _0958_ (.B(_0247_),
    .C(_0249_),
    .A(\top_inst.address[5] ),
    .Y(_0320_),
    .D(_0317_));
 sg13g2_nand2b_1 _0959_ (.Y(_0321_),
    .B(_0245_),
    .A_N(_0244_));
 sg13g2_o21ai_1 _0960_ (.B1(_0321_),
    .Y(_0322_),
    .A1(\top_inst.address[6] ),
    .A2(_0320_));
 sg13g2_a21o_1 _0961_ (.A2(_0320_),
    .A1(\top_inst.address[6] ),
    .B1(_0322_),
    .X(_0038_));
 sg13g2_a21oi_1 _0962_ (.A1(_0250_),
    .A2(_0317_),
    .Y(_0323_),
    .B1(\top_inst.address[5] ));
 sg13g2_o21ai_1 _0963_ (.B1(_0321_),
    .Y(_0039_),
    .A1(_0319_),
    .A2(_0323_));
 sg13g2_o21ai_1 _0964_ (.B1(_0246_),
    .Y(_0324_),
    .A1(_0154_),
    .A2(_0316_));
 sg13g2_a21oi_1 _0965_ (.A1(_0250_),
    .A2(_0324_),
    .Y(_0325_),
    .B1(\top_inst.address[4] ));
 sg13g2_o21ai_1 _0966_ (.B1(_0318_),
    .Y(_0326_),
    .A1(\top_inst.controller_inst.state[2] ),
    .A2(_0203_));
 sg13g2_a21oi_1 _0967_ (.A1(_0009_),
    .A2(_0326_),
    .Y(_0040_),
    .B1(_0325_));
 sg13g2_xnor2_1 _0968_ (.Y(_0327_),
    .A(_0154_),
    .B(_0316_));
 sg13g2_nor2_1 _0969_ (.A(\top_inst.address[3] ),
    .B(_0250_),
    .Y(_0328_));
 sg13g2_a21oi_1 _0970_ (.A1(_0009_),
    .A2(_0327_),
    .Y(_0041_),
    .B1(_0328_));
 sg13g2_o21ai_1 _0971_ (.B1(_0250_),
    .Y(_0329_),
    .A1(_0194_),
    .A2(_0245_));
 sg13g2_o21ai_1 _0972_ (.B1(_0316_),
    .Y(_0330_),
    .A1(\top_inst.controller_inst.state[2] ),
    .A2(_0203_));
 sg13g2_a22oi_1 _0973_ (.Y(_0042_),
    .B1(_0330_),
    .B2(_0009_),
    .A2(_0329_),
    .A1(_0153_));
 sg13g2_nand3_1 _0974_ (.B(_0194_),
    .C(_0202_),
    .A(\top_inst.controller_inst.state[1] ),
    .Y(_0331_));
 sg13g2_and2_1 _0975_ (.A(_0009_),
    .B(_0331_),
    .X(_0332_));
 sg13g2_nor2_1 _0976_ (.A(net220),
    .B(_0250_),
    .Y(_0333_));
 sg13g2_a21oi_1 _0977_ (.A1(_0253_),
    .A2(_0332_),
    .Y(_0043_),
    .B1(_0333_));
 sg13g2_nor2_1 _0978_ (.A(\top_inst.address[0] ),
    .B(_0250_),
    .Y(_0334_));
 sg13g2_a21oi_1 _0979_ (.A1(\top_inst.address[0] ),
    .A2(_0332_),
    .Y(_0044_),
    .B1(_0334_));
 sg13g2_nor4_1 _0980_ (.A(_0152_),
    .B(_0153_),
    .C(_0154_),
    .D(_0197_),
    .Y(_0335_));
 sg13g2_a21oi_2 _0981_ (.B1(_0335_),
    .Y(_0336_),
    .A2(_0202_),
    .A1(_0152_));
 sg13g2_or2_2 _0982_ (.X(_0337_),
    .B(_0336_),
    .A(_0252_));
 sg13g2_nor2_2 _0983_ (.A(_0152_),
    .B(\top_inst.address[1] ),
    .Y(_0338_));
 sg13g2_nand2_1 _0984_ (.Y(_0339_),
    .A(_0202_),
    .B(_0338_));
 sg13g2_and3_1 _0985_ (.X(_0340_),
    .A(_0152_),
    .B(net220),
    .C(_0196_));
 sg13g2_nand3_1 _0986_ (.B(\top_inst.address[3] ),
    .C(_0340_),
    .A(\top_inst.address[2] ),
    .Y(_0341_));
 sg13g2_nand3_1 _0987_ (.B(_0339_),
    .C(_0341_),
    .A(_0337_),
    .Y(_0045_));
 sg13g2_nor2_2 _0988_ (.A(net220),
    .B(_0198_),
    .Y(_0342_));
 sg13g2_nand2_2 _0989_ (.Y(_0343_),
    .A(_0152_),
    .B(_0342_));
 sg13g2_inv_1 _0990_ (.Y(_0047_),
    .A(_0343_));
 sg13g2_nand2_1 _0991_ (.Y(_0046_),
    .A(_0337_),
    .B(_0343_));
 sg13g2_and2_1 _0992_ (.A(_0254_),
    .B(_0337_),
    .X(_0344_));
 sg13g2_nor2_2 _0993_ (.A(\top_inst.address[0] ),
    .B(_0198_),
    .Y(_0345_));
 sg13g2_nor2_2 _0994_ (.A(_0342_),
    .B(_0345_),
    .Y(_0346_));
 sg13g2_nand2_1 _0995_ (.Y(_0049_),
    .A(_0344_),
    .B(_0346_));
 sg13g2_a22oi_1 _0996_ (.Y(_0347_),
    .B1(_0209_),
    .B2(_0194_),
    .A2(_0202_),
    .A1(_0152_));
 sg13g2_nor2_1 _0997_ (.A(_0340_),
    .B(_0345_),
    .Y(_0348_));
 sg13g2_nand3_1 _0998_ (.B(_0196_),
    .C(_0251_),
    .A(\top_inst.address[2] ),
    .Y(_0349_));
 sg13g2_nand3_1 _0999_ (.B(_0348_),
    .C(_0349_),
    .A(_0347_),
    .Y(_0050_));
 sg13g2_nand2_2 _1000_ (.Y(_0350_),
    .A(_0195_),
    .B(_0209_));
 sg13g2_nand2b_1 _1001_ (.Y(_0051_),
    .B(_0350_),
    .A_N(_0045_));
 sg13g2_nand2_1 _1002_ (.Y(_0351_),
    .A(_0209_),
    .B(_0338_));
 sg13g2_nand2_2 _1003_ (.Y(_0352_),
    .A(_0152_),
    .B(_0209_));
 sg13g2_nand3_1 _1004_ (.B(_0343_),
    .C(_0352_),
    .A(_0255_),
    .Y(_0076_));
 sg13g2_and2_2 _1005_ (.A(_0256_),
    .B(_0337_),
    .X(_0353_));
 sg13g2_nand2_1 _1006_ (.Y(_0077_),
    .A(_0352_),
    .B(_0353_));
 sg13g2_nand3_1 _1007_ (.B(_0352_),
    .C(_0353_),
    .A(_0343_),
    .Y(_0075_));
 sg13g2_nand2b_1 _1008_ (.Y(_0052_),
    .B(_0351_),
    .A_N(_0075_));
 sg13g2_nand2_1 _1009_ (.Y(_0354_),
    .A(_0251_),
    .B(_0257_));
 sg13g2_nand3_1 _1010_ (.B(_0353_),
    .C(_0354_),
    .A(_0350_),
    .Y(_0053_));
 sg13g2_a21oi_2 _1011_ (.B1(_0342_),
    .Y(_0355_),
    .A2(_0257_),
    .A1(net220));
 sg13g2_nand3_1 _1012_ (.B(_0350_),
    .C(_0355_),
    .A(_0344_),
    .Y(_0054_));
 sg13g2_and3_1 _1013_ (.X(_0055_),
    .A(net250),
    .B(net215),
    .C(_0007_));
 sg13g2_nor2_1 _1014_ (.A(\top_inst.spi_inst.counter[0] ),
    .B(\top_inst.spi_inst.counter[1] ),
    .Y(_0356_));
 sg13g2_nor3_1 _1015_ (.A(_0228_),
    .B(_0239_),
    .C(_0356_),
    .Y(_0056_));
 sg13g2_nor2_1 _1016_ (.A(\top_inst.spi_inst.counter[2] ),
    .B(_0228_),
    .Y(_0357_));
 sg13g2_nor3_1 _1017_ (.A(_0229_),
    .B(_0239_),
    .C(_0357_),
    .Y(_0057_));
 sg13g2_nor2_1 _1018_ (.A(\top_inst.spi_inst.counter[3] ),
    .B(_0229_),
    .Y(_0358_));
 sg13g2_nor3_1 _1019_ (.A(_0230_),
    .B(_0239_),
    .C(_0358_),
    .Y(_0058_));
 sg13g2_nor2_1 _1020_ (.A(\top_inst.spi_inst.counter[4] ),
    .B(_0230_),
    .Y(_0359_));
 sg13g2_nor3_1 _1021_ (.A(_0231_),
    .B(_0239_),
    .C(_0359_),
    .Y(_0059_));
 sg13g2_xnor2_1 _1022_ (.Y(_0360_),
    .A(\top_inst.spi_inst.counter[5] ),
    .B(_0231_));
 sg13g2_nor2_1 _1023_ (.A(_0239_),
    .B(_0360_),
    .Y(_0060_));
 sg13g2_xor2_1 _1024_ (.B(_0232_),
    .A(\top_inst.spi_inst.counter[6] ),
    .X(_0361_));
 sg13g2_nor2_1 _1025_ (.A(_0239_),
    .B(_0361_),
    .Y(_0061_));
 sg13g2_and2_1 _1026_ (.A(\top_inst.spi_cs_n ),
    .B(net211),
    .X(_0362_));
 sg13g2_nand2_1 _1027_ (.Y(_0363_),
    .A(net217),
    .B(\top_inst.data[0] ));
 sg13g2_o21ai_1 _1028_ (.B1(net248),
    .Y(_0364_),
    .A1(\top_inst.spi_inst.buffer[0] ),
    .A2(_0362_));
 sg13g2_a21oi_1 _1029_ (.A1(_0362_),
    .A2(_0363_),
    .Y(_0062_),
    .B1(_0364_));
 sg13g2_nand2b_1 _1030_ (.Y(_0365_),
    .B(_0252_),
    .A_N(_0198_));
 sg13g2_nand4_1 _1031_ (.B(_0337_),
    .C(_0343_),
    .A(_0258_),
    .Y(_0063_),
    .D(_0365_));
 sg13g2_nor2_1 _1032_ (.A(\top_inst.address[0] ),
    .B(_0258_),
    .Y(_0366_));
 sg13g2_a21o_1 _1033_ (.A2(_0345_),
    .A1(net220),
    .B1(_0366_),
    .X(_0367_));
 sg13g2_nand2b_1 _1034_ (.Y(_0064_),
    .B(_0254_),
    .A_N(_0367_));
 sg13g2_nand3b_1 _1035_ (.B(_0255_),
    .C(_0344_),
    .Y(_0065_),
    .A_N(_0367_));
 sg13g2_nand2b_1 _1036_ (.Y(_0066_),
    .B(_0343_),
    .A_N(_0065_));
 sg13g2_nand2_1 _1037_ (.Y(_0067_),
    .A(_0258_),
    .B(_0346_));
 sg13g2_nand2_1 _1038_ (.Y(_0068_),
    .A(_0336_),
    .B(_0355_));
 sg13g2_a21oi_2 _1039_ (.B1(_0067_),
    .Y(_0368_),
    .A2(_0338_),
    .A1(_0257_));
 sg13g2_inv_1 _1040_ (.Y(_0072_),
    .A(_0368_));
 sg13g2_nand4_1 _1041_ (.B(_0336_),
    .C(_0354_),
    .A(_0199_),
    .Y(_0069_),
    .D(_0368_));
 sg13g2_and3_1 _1042_ (.X(_0070_),
    .A(_0349_),
    .B(_0353_),
    .C(_0368_));
 sg13g2_nand2_1 _1043_ (.Y(_0071_),
    .A(_0336_),
    .B(_0368_));
 sg13g2_nand2_1 _1044_ (.Y(_0073_),
    .A(_0337_),
    .B(_0352_));
 sg13g2_nand3_1 _1045_ (.B(_0343_),
    .C(_0352_),
    .A(_0337_),
    .Y(_0074_));
 sg13g2_a22oi_1 _1046_ (.Y(_0369_),
    .B1(_0257_),
    .B2(_0338_),
    .A2(_0209_),
    .A1(_0152_));
 sg13g2_nand3_1 _1047_ (.B(_0354_),
    .C(_0369_),
    .A(_0353_),
    .Y(_0078_));
 sg13g2_nor2b_1 _1048_ (.A(_0366_),
    .B_N(_0369_),
    .Y(_0370_));
 sg13g2_nand3_1 _1049_ (.B(_0354_),
    .C(_0370_),
    .A(_0336_),
    .Y(_0079_));
 sg13g2_nand3_1 _1050_ (.B(_0336_),
    .C(_0352_),
    .A(_0259_),
    .Y(_0080_));
 sg13g2_nand4_1 _1051_ (.B(_0344_),
    .C(_0346_),
    .A(_0259_),
    .Y(_0081_),
    .D(_0351_));
 sg13g2_nand3_1 _1052_ (.B(_0352_),
    .C(_0355_),
    .A(_0256_),
    .Y(_0082_));
 sg13g2_nand4_1 _1053_ (.B(_0346_),
    .C(_0352_),
    .A(_0259_),
    .Y(_0083_),
    .D(_0353_));
 sg13g2_nand3_1 _1054_ (.B(_0365_),
    .C(_0370_),
    .A(_0256_),
    .Y(_0084_));
 sg13g2_nor2_2 _1055_ (.A(_0235_),
    .B(_0239_),
    .Y(_0371_));
 sg13g2_and2_1 _1056_ (.A(net247),
    .B(_0235_),
    .X(_0372_));
 sg13g2_a22oi_1 _1057_ (.Y(_0373_),
    .B1(net197),
    .B2(\top_inst.spi_inst.buffer[1] ),
    .A2(net204),
    .A1(\top_inst.spi_inst.buffer[0] ));
 sg13g2_o21ai_1 _1058_ (.B1(_0373_),
    .Y(_0085_),
    .A1(_0177_),
    .A2(net208));
 sg13g2_a221oi_1 _1059_ (.B2(net217),
    .C1(net212),
    .B1(\top_inst.data[2] ),
    .A1(\top_inst.spi_inst.buffer[1] ),
    .Y(_0374_),
    .A2(net213));
 sg13g2_o21ai_1 _1060_ (.B1(net247),
    .Y(_0375_),
    .A1(\top_inst.spi_inst.buffer[2] ),
    .A2(net211));
 sg13g2_nor2_1 _1061_ (.A(_0374_),
    .B(_0375_),
    .Y(_0086_));
 sg13g2_a221oi_1 _1062_ (.B2(net217),
    .C1(net212),
    .B1(\top_inst.data[2] ),
    .A1(\top_inst.spi_inst.buffer[2] ),
    .Y(_0376_),
    .A2(net213));
 sg13g2_o21ai_1 _1063_ (.B1(net247),
    .Y(_0377_),
    .A1(\top_inst.spi_inst.buffer[3] ),
    .A2(net211));
 sg13g2_nor2_1 _1064_ (.A(_0376_),
    .B(_0377_),
    .Y(_0087_));
 sg13g2_a22oi_1 _1065_ (.Y(_0378_),
    .B1(net197),
    .B2(\top_inst.spi_inst.buffer[4] ),
    .A2(net204),
    .A1(\top_inst.spi_inst.buffer[3] ));
 sg13g2_o21ai_1 _1066_ (.B1(_0378_),
    .Y(_0088_),
    .A1(_0178_),
    .A2(net208));
 sg13g2_a22oi_1 _1067_ (.Y(_0379_),
    .B1(net196),
    .B2(\top_inst.spi_inst.buffer[5] ),
    .A2(net203),
    .A1(\top_inst.spi_inst.buffer[4] ));
 sg13g2_o21ai_1 _1068_ (.B1(_0379_),
    .Y(_0089_),
    .A1(_0179_),
    .A2(net208));
 sg13g2_a22oi_1 _1069_ (.Y(_0380_),
    .B1(net196),
    .B2(\top_inst.spi_inst.buffer[6] ),
    .A2(net203),
    .A1(\top_inst.spi_inst.buffer[5] ));
 sg13g2_o21ai_1 _1070_ (.B1(_0380_),
    .Y(_0090_),
    .A1(_0180_),
    .A2(net208));
 sg13g2_a22oi_1 _1071_ (.Y(_0381_),
    .B1(net196),
    .B2(\top_inst.spi_inst.buffer[7] ),
    .A2(net203),
    .A1(\top_inst.spi_inst.buffer[6] ));
 sg13g2_o21ai_1 _1072_ (.B1(_0381_),
    .Y(_0091_),
    .A1(_0181_),
    .A2(net208));
 sg13g2_nand2_1 _1073_ (.Y(_0382_),
    .A(\top_inst.spi_inst.buffer[7] ),
    .B(net213));
 sg13g2_a21oi_2 _1074_ (.B1(net212),
    .Y(_0383_),
    .A2(\top_inst.data[20] ),
    .A1(net217));
 sg13g2_o21ai_1 _1075_ (.B1(net247),
    .Y(_0384_),
    .A1(\top_inst.spi_inst.buffer[8] ),
    .A2(net211));
 sg13g2_a21oi_1 _1076_ (.A1(_0382_),
    .A2(_0383_),
    .Y(_0092_),
    .B1(_0384_));
 sg13g2_nand2_1 _1077_ (.Y(_0385_),
    .A(\top_inst.spi_inst.buffer[8] ),
    .B(net213));
 sg13g2_a21oi_2 _1078_ (.B1(net212),
    .Y(_0386_),
    .A2(\top_inst.data[21] ),
    .A1(net218));
 sg13g2_o21ai_1 _1079_ (.B1(net249),
    .Y(_0387_),
    .A1(\top_inst.spi_inst.buffer[9] ),
    .A2(net210));
 sg13g2_a21oi_1 _1080_ (.A1(_0385_),
    .A2(_0386_),
    .Y(_0093_),
    .B1(_0387_));
 sg13g2_nand2_1 _1081_ (.Y(_0388_),
    .A(\top_inst.spi_inst.buffer[9] ),
    .B(net215));
 sg13g2_a21oi_2 _1082_ (.B1(net212),
    .Y(_0389_),
    .A2(\top_inst.data[10] ),
    .A1(net218));
 sg13g2_o21ai_1 _1083_ (.B1(net251),
    .Y(_0390_),
    .A1(\top_inst.spi_inst.buffer[10] ),
    .A2(net209));
 sg13g2_a21oi_1 _1084_ (.A1(_0388_),
    .A2(_0389_),
    .Y(_0094_),
    .B1(_0390_));
 sg13g2_nand2_1 _1085_ (.Y(_0391_),
    .A(\top_inst.spi_inst.buffer[10] ),
    .B(net214));
 sg13g2_a21oi_2 _1086_ (.B1(net212),
    .Y(_0392_),
    .A2(\top_inst.data[11] ),
    .A1(net218));
 sg13g2_o21ai_1 _1087_ (.B1(net249),
    .Y(_0393_),
    .A1(\top_inst.spi_inst.buffer[11] ),
    .A2(net209));
 sg13g2_a21oi_1 _1088_ (.A1(_0391_),
    .A2(_0392_),
    .Y(_0095_),
    .B1(_0393_));
 sg13g2_a22oi_1 _1089_ (.Y(_0394_),
    .B1(net194),
    .B2(\top_inst.spi_inst.buffer[12] ),
    .A2(net201),
    .A1(\top_inst.spi_inst.buffer[11] ));
 sg13g2_inv_1 _1090_ (.Y(_0096_),
    .A(_0394_));
 sg13g2_a22oi_1 _1091_ (.Y(_0395_),
    .B1(net192),
    .B2(\top_inst.spi_inst.buffer[13] ),
    .A2(net199),
    .A1(\top_inst.spi_inst.buffer[12] ));
 sg13g2_inv_1 _1092_ (.Y(_0097_),
    .A(_0395_));
 sg13g2_a22oi_1 _1093_ (.Y(_0396_),
    .B1(net192),
    .B2(\top_inst.spi_inst.buffer[14] ),
    .A2(net199),
    .A1(\top_inst.spi_inst.buffer[13] ));
 sg13g2_inv_1 _1094_ (.Y(_0098_),
    .A(_0396_));
 sg13g2_a22oi_1 _1095_ (.Y(_0397_),
    .B1(net192),
    .B2(\top_inst.spi_inst.buffer[15] ),
    .A2(net199),
    .A1(\top_inst.spi_inst.buffer[14] ));
 sg13g2_inv_1 _1096_ (.Y(_0099_),
    .A(_0397_));
 sg13g2_a22oi_1 _1097_ (.Y(_0398_),
    .B1(net191),
    .B2(\top_inst.spi_inst.buffer[16] ),
    .A2(net198),
    .A1(\top_inst.spi_inst.buffer[15] ));
 sg13g2_o21ai_1 _1098_ (.B1(_0398_),
    .Y(_0100_),
    .A1(_0156_),
    .A2(net205));
 sg13g2_a22oi_1 _1099_ (.Y(_0399_),
    .B1(net195),
    .B2(\top_inst.spi_inst.buffer[17] ),
    .A2(net202),
    .A1(\top_inst.spi_inst.buffer[16] ));
 sg13g2_o21ai_1 _1100_ (.B1(_0399_),
    .Y(_0101_),
    .A1(_0157_),
    .A2(net207));
 sg13g2_a22oi_1 _1101_ (.Y(_0400_),
    .B1(net195),
    .B2(\top_inst.spi_inst.buffer[18] ),
    .A2(net202),
    .A1(\top_inst.spi_inst.buffer[17] ));
 sg13g2_o21ai_1 _1102_ (.B1(_0400_),
    .Y(_0102_),
    .A1(_0158_),
    .A2(net207));
 sg13g2_a22oi_1 _1103_ (.Y(_0401_),
    .B1(net195),
    .B2(\top_inst.spi_inst.buffer[19] ),
    .A2(net202),
    .A1(\top_inst.spi_inst.buffer[18] ));
 sg13g2_o21ai_1 _1104_ (.B1(_0401_),
    .Y(_0103_),
    .A1(_0159_),
    .A2(net207));
 sg13g2_a22oi_1 _1105_ (.Y(_0402_),
    .B1(net195),
    .B2(\top_inst.spi_inst.buffer[20] ),
    .A2(net202),
    .A1(\top_inst.spi_inst.buffer[19] ));
 sg13g2_o21ai_1 _1106_ (.B1(_0402_),
    .Y(_0104_),
    .A1(_0160_),
    .A2(net207));
 sg13g2_a22oi_1 _1107_ (.Y(_0403_),
    .B1(net195),
    .B2(\top_inst.spi_inst.buffer[21] ),
    .A2(net202),
    .A1(\top_inst.spi_inst.buffer[20] ));
 sg13g2_o21ai_1 _1108_ (.B1(_0403_),
    .Y(_0105_),
    .A1(_0161_),
    .A2(net207));
 sg13g2_a22oi_1 _1109_ (.Y(_0404_),
    .B1(net195),
    .B2(\top_inst.spi_inst.buffer[22] ),
    .A2(net202),
    .A1(\top_inst.spi_inst.buffer[21] ));
 sg13g2_o21ai_1 _1110_ (.B1(_0404_),
    .Y(_0106_),
    .A1(_0162_),
    .A2(net207));
 sg13g2_a22oi_1 _1111_ (.Y(_0405_),
    .B1(net195),
    .B2(\top_inst.spi_inst.buffer[23] ),
    .A2(net202),
    .A1(\top_inst.spi_inst.buffer[22] ));
 sg13g2_o21ai_1 _1112_ (.B1(_0405_),
    .Y(_0107_),
    .A1(_0163_),
    .A2(net207));
 sg13g2_nand2_1 _1113_ (.Y(_0406_),
    .A(\top_inst.spi_inst.buffer[23] ),
    .B(net213));
 sg13g2_o21ai_1 _1114_ (.B1(net249),
    .Y(_0407_),
    .A1(\top_inst.spi_inst.buffer[24] ),
    .A2(net210));
 sg13g2_a21oi_1 _1115_ (.A1(_0383_),
    .A2(_0406_),
    .Y(_0108_),
    .B1(_0407_));
 sg13g2_nand2_1 _1116_ (.Y(_0408_),
    .A(\top_inst.spi_inst.buffer[24] ),
    .B(net214));
 sg13g2_o21ai_1 _1117_ (.B1(net249),
    .Y(_0409_),
    .A1(\top_inst.spi_inst.buffer[25] ),
    .A2(net209));
 sg13g2_a21oi_1 _1118_ (.A1(_0386_),
    .A2(_0408_),
    .Y(_0109_),
    .B1(_0409_));
 sg13g2_nand2_1 _1119_ (.Y(_0410_),
    .A(\top_inst.spi_inst.buffer[25] ),
    .B(net214));
 sg13g2_o21ai_1 _1120_ (.B1(net249),
    .Y(_0411_),
    .A1(\top_inst.spi_inst.buffer[26] ),
    .A2(net209));
 sg13g2_a21oi_1 _1121_ (.A1(_0389_),
    .A2(_0410_),
    .Y(_0110_),
    .B1(_0411_));
 sg13g2_nand2_1 _1122_ (.Y(_0412_),
    .A(\top_inst.spi_inst.buffer[26] ),
    .B(net214));
 sg13g2_o21ai_1 _1123_ (.B1(net249),
    .Y(_0413_),
    .A1(\top_inst.spi_inst.buffer[27] ),
    .A2(net209));
 sg13g2_a21oi_1 _1124_ (.A1(_0392_),
    .A2(_0412_),
    .Y(_0111_),
    .B1(_0413_));
 sg13g2_a22oi_1 _1125_ (.Y(_0414_),
    .B1(net193),
    .B2(\top_inst.spi_inst.buffer[28] ),
    .A2(net200),
    .A1(\top_inst.spi_inst.buffer[27] ));
 sg13g2_inv_1 _1126_ (.Y(_0112_),
    .A(_0414_));
 sg13g2_a22oi_1 _1127_ (.Y(_0415_),
    .B1(net193),
    .B2(\top_inst.spi_inst.buffer[29] ),
    .A2(net200),
    .A1(\top_inst.spi_inst.buffer[28] ));
 sg13g2_inv_1 _1128_ (.Y(_0113_),
    .A(_0415_));
 sg13g2_a22oi_1 _1129_ (.Y(_0416_),
    .B1(net192),
    .B2(\top_inst.spi_inst.buffer[30] ),
    .A2(net199),
    .A1(\top_inst.spi_inst.buffer[29] ));
 sg13g2_inv_1 _1130_ (.Y(_0114_),
    .A(_0416_));
 sg13g2_a22oi_1 _1131_ (.Y(_0417_),
    .B1(net191),
    .B2(\top_inst.spi_inst.buffer[31] ),
    .A2(net198),
    .A1(\top_inst.spi_inst.buffer[30] ));
 sg13g2_inv_1 _1132_ (.Y(_0115_),
    .A(_0417_));
 sg13g2_a22oi_1 _1133_ (.Y(_0418_),
    .B1(net191),
    .B2(\top_inst.spi_inst.buffer[32] ),
    .A2(net198),
    .A1(\top_inst.spi_inst.buffer[31] ));
 sg13g2_o21ai_1 _1134_ (.B1(_0418_),
    .Y(_0116_),
    .A1(_0169_),
    .A2(net205));
 sg13g2_a22oi_1 _1135_ (.Y(_0419_),
    .B1(net191),
    .B2(\top_inst.spi_inst.buffer[33] ),
    .A2(net198),
    .A1(\top_inst.spi_inst.buffer[32] ));
 sg13g2_o21ai_1 _1136_ (.B1(_0419_),
    .Y(_0117_),
    .A1(_0170_),
    .A2(net205));
 sg13g2_a22oi_1 _1137_ (.Y(_0420_),
    .B1(net191),
    .B2(\top_inst.spi_inst.buffer[34] ),
    .A2(net198),
    .A1(\top_inst.spi_inst.buffer[33] ));
 sg13g2_o21ai_1 _1138_ (.B1(_0420_),
    .Y(_0118_),
    .A1(_0171_),
    .A2(net205));
 sg13g2_a22oi_1 _1139_ (.Y(_0421_),
    .B1(net191),
    .B2(\top_inst.spi_inst.buffer[35] ),
    .A2(net198),
    .A1(\top_inst.spi_inst.buffer[34] ));
 sg13g2_o21ai_1 _1140_ (.B1(_0421_),
    .Y(_0119_),
    .A1(_0172_),
    .A2(net205));
 sg13g2_a22oi_1 _1141_ (.Y(_0422_),
    .B1(net191),
    .B2(\top_inst.spi_inst.buffer[36] ),
    .A2(net198),
    .A1(\top_inst.spi_inst.buffer[35] ));
 sg13g2_o21ai_1 _1142_ (.B1(_0422_),
    .Y(_0120_),
    .A1(_0173_),
    .A2(net205));
 sg13g2_a22oi_1 _1143_ (.Y(_0423_),
    .B1(net191),
    .B2(\top_inst.spi_inst.buffer[37] ),
    .A2(net198),
    .A1(\top_inst.spi_inst.buffer[36] ));
 sg13g2_o21ai_1 _1144_ (.B1(_0423_),
    .Y(_0121_),
    .A1(_0174_),
    .A2(net205));
 sg13g2_a22oi_1 _1145_ (.Y(_0424_),
    .B1(net193),
    .B2(\top_inst.spi_inst.buffer[38] ),
    .A2(net200),
    .A1(\top_inst.spi_inst.buffer[37] ));
 sg13g2_o21ai_1 _1146_ (.B1(_0424_),
    .Y(_0122_),
    .A1(_0175_),
    .A2(net205));
 sg13g2_a22oi_1 _1147_ (.Y(_0425_),
    .B1(net193),
    .B2(\top_inst.spi_inst.buffer[39] ),
    .A2(net200),
    .A1(\top_inst.spi_inst.buffer[38] ));
 sg13g2_o21ai_1 _1148_ (.B1(_0425_),
    .Y(_0123_),
    .A1(_0176_),
    .A2(net206));
 sg13g2_nand2_1 _1149_ (.Y(_0426_),
    .A(\top_inst.spi_inst.buffer[39] ),
    .B(net214));
 sg13g2_o21ai_1 _1150_ (.B1(net251),
    .Y(_0427_),
    .A1(\top_inst.spi_inst.buffer[40] ),
    .A2(net209));
 sg13g2_a21oi_1 _1151_ (.A1(_0383_),
    .A2(_0426_),
    .Y(_0124_),
    .B1(_0427_));
 sg13g2_nand2_1 _1152_ (.Y(_0428_),
    .A(\top_inst.spi_inst.buffer[40] ),
    .B(net214));
 sg13g2_o21ai_1 _1153_ (.B1(net249),
    .Y(_0429_),
    .A1(\top_inst.spi_inst.buffer[41] ),
    .A2(net210));
 sg13g2_a21oi_1 _1154_ (.A1(_0386_),
    .A2(_0428_),
    .Y(_0125_),
    .B1(_0429_));
 sg13g2_nand2_1 _1155_ (.Y(_0430_),
    .A(\top_inst.spi_inst.buffer[41] ),
    .B(net215));
 sg13g2_o21ai_1 _1156_ (.B1(net250),
    .Y(_0431_),
    .A1(\top_inst.spi_inst.buffer[42] ),
    .A2(net209));
 sg13g2_a21oi_1 _1157_ (.A1(_0389_),
    .A2(_0430_),
    .Y(_0126_),
    .B1(_0431_));
 sg13g2_nand2_1 _1158_ (.Y(_0432_),
    .A(\top_inst.spi_inst.buffer[42] ),
    .B(net215));
 sg13g2_o21ai_1 _1159_ (.B1(net251),
    .Y(_0433_),
    .A1(\top_inst.spi_inst.buffer[43] ),
    .A2(net210));
 sg13g2_a21oi_1 _1160_ (.A1(_0392_),
    .A2(_0432_),
    .Y(_0127_),
    .B1(_0433_));
 sg13g2_a22oi_1 _1161_ (.Y(_0434_),
    .B1(net197),
    .B2(\top_inst.spi_inst.buffer[44] ),
    .A2(net204),
    .A1(\top_inst.spi_inst.buffer[43] ));
 sg13g2_inv_1 _1162_ (.Y(_0128_),
    .A(_0434_));
 sg13g2_a22oi_1 _1163_ (.Y(_0435_),
    .B1(net197),
    .B2(\top_inst.spi_inst.buffer[45] ),
    .A2(net204),
    .A1(\top_inst.spi_inst.buffer[44] ));
 sg13g2_inv_1 _1164_ (.Y(_0129_),
    .A(_0435_));
 sg13g2_a22oi_1 _1165_ (.Y(_0436_),
    .B1(net197),
    .B2(\top_inst.spi_inst.buffer[46] ),
    .A2(net204),
    .A1(\top_inst.spi_inst.buffer[45] ));
 sg13g2_inv_1 _1166_ (.Y(_0130_),
    .A(_0436_));
 sg13g2_a22oi_1 _1167_ (.Y(_0437_),
    .B1(net197),
    .B2(\top_inst.spi_inst.buffer[47] ),
    .A2(net204),
    .A1(\top_inst.spi_inst.buffer[46] ));
 sg13g2_inv_1 _1168_ (.Y(_0131_),
    .A(_0437_));
 sg13g2_a22oi_1 _1169_ (.Y(_0438_),
    .B1(net196),
    .B2(\top_inst.spi_inst.buffer[48] ),
    .A2(net203),
    .A1(\top_inst.spi_inst.buffer[47] ));
 sg13g2_o21ai_1 _1170_ (.B1(_0438_),
    .Y(_0132_),
    .A1(_0164_),
    .A2(net208));
 sg13g2_a221oi_1 _1171_ (.B2(net218),
    .C1(net212),
    .B1(\top_inst.data[37] ),
    .A1(\top_inst.spi_inst.buffer[48] ),
    .Y(_0439_),
    .A2(net213));
 sg13g2_o21ai_1 _1172_ (.B1(net248),
    .Y(_0440_),
    .A1(\top_inst.spi_inst.buffer[49] ),
    .A2(net211));
 sg13g2_nor2_1 _1173_ (.A(_0439_),
    .B(_0440_),
    .Y(_0133_));
 sg13g2_a221oi_1 _1174_ (.B2(net217),
    .C1(net212),
    .B1(\top_inst.data[37] ),
    .A1(\top_inst.spi_inst.buffer[49] ),
    .Y(_0441_),
    .A2(net213));
 sg13g2_o21ai_1 _1175_ (.B1(net247),
    .Y(_0442_),
    .A1(\top_inst.spi_inst.buffer[50] ),
    .A2(net211));
 sg13g2_nor2_1 _1176_ (.A(_0441_),
    .B(_0442_),
    .Y(_0134_));
 sg13g2_a22oi_1 _1177_ (.Y(_0443_),
    .B1(net197),
    .B2(\top_inst.spi_inst.buffer[51] ),
    .A2(net204),
    .A1(\top_inst.spi_inst.buffer[50] ));
 sg13g2_o21ai_1 _1178_ (.B1(_0443_),
    .Y(_0135_),
    .A1(_0165_),
    .A2(_0238_));
 sg13g2_a22oi_1 _1179_ (.Y(_0444_),
    .B1(net193),
    .B2(\top_inst.spi_inst.buffer[52] ),
    .A2(net200),
    .A1(\top_inst.spi_inst.buffer[51] ));
 sg13g2_o21ai_1 _1180_ (.B1(_0444_),
    .Y(_0136_),
    .A1(_0166_),
    .A2(net206));
 sg13g2_a22oi_1 _1181_ (.Y(_0445_),
    .B1(net193),
    .B2(\top_inst.spi_inst.buffer[53] ),
    .A2(net200),
    .A1(\top_inst.spi_inst.buffer[52] ));
 sg13g2_o21ai_1 _1182_ (.B1(_0445_),
    .Y(_0137_),
    .A1(_0167_),
    .A2(net206));
 sg13g2_a22oi_1 _1183_ (.Y(_0446_),
    .B1(net193),
    .B2(\top_inst.spi_inst.buffer[54] ),
    .A2(net200),
    .A1(\top_inst.spi_inst.buffer[53] ));
 sg13g2_o21ai_1 _1184_ (.B1(_0446_),
    .Y(_0138_),
    .A1(_0168_),
    .A2(net206));
 sg13g2_a22oi_1 _1185_ (.Y(_0447_),
    .B1(net193),
    .B2(\top_inst.spi_inst.buffer[55] ),
    .A2(net200),
    .A1(\top_inst.spi_inst.buffer[54] ));
 sg13g2_inv_1 _1186_ (.Y(_0139_),
    .A(_0447_));
 sg13g2_nand2_1 _1187_ (.Y(_0448_),
    .A(\top_inst.spi_inst.buffer[55] ),
    .B(net214));
 sg13g2_o21ai_1 _1188_ (.B1(net251),
    .Y(_0449_),
    .A1(\top_inst.spi_inst.buffer[56] ),
    .A2(net209));
 sg13g2_a21oi_1 _1189_ (.A1(_0383_),
    .A2(_0448_),
    .Y(_0140_),
    .B1(_0449_));
 sg13g2_nand2_1 _1190_ (.Y(_0450_),
    .A(\top_inst.spi_inst.buffer[56] ),
    .B(net214));
 sg13g2_o21ai_1 _1191_ (.B1(net249),
    .Y(_0451_),
    .A1(\top_inst.spi_inst.buffer[57] ),
    .A2(net210));
 sg13g2_a21oi_1 _1192_ (.A1(_0386_),
    .A2(_0450_),
    .Y(_0141_),
    .B1(_0451_));
 sg13g2_nand2_1 _1193_ (.Y(_0452_),
    .A(\top_inst.spi_inst.buffer[57] ),
    .B(net215));
 sg13g2_o21ai_1 _1194_ (.B1(net250),
    .Y(_0453_),
    .A1(\top_inst.spi_inst.buffer[58] ),
    .A2(net210));
 sg13g2_a21oi_1 _1195_ (.A1(_0389_),
    .A2(_0452_),
    .Y(_0142_),
    .B1(_0453_));
 sg13g2_nand2_1 _1196_ (.Y(_0454_),
    .A(\top_inst.spi_inst.buffer[58] ),
    .B(net215));
 sg13g2_o21ai_1 _1197_ (.B1(net248),
    .Y(_0455_),
    .A1(\top_inst.spi_inst.buffer[59] ),
    .A2(net211));
 sg13g2_a21oi_1 _1198_ (.A1(_0392_),
    .A2(_0454_),
    .Y(_0143_),
    .B1(_0455_));
 sg13g2_a22oi_1 _1199_ (.Y(_0456_),
    .B1(net196),
    .B2(\top_inst.spi_inst.buffer[60] ),
    .A2(net203),
    .A1(\top_inst.spi_inst.buffer[59] ));
 sg13g2_inv_1 _1200_ (.Y(_0144_),
    .A(_0456_));
 sg13g2_a22oi_1 _1201_ (.Y(_0457_),
    .B1(net196),
    .B2(\top_inst.spi_inst.buffer[61] ),
    .A2(net203),
    .A1(\top_inst.spi_inst.buffer[60] ));
 sg13g2_inv_1 _1202_ (.Y(_0145_),
    .A(_0457_));
 sg13g2_a22oi_1 _1203_ (.Y(_0458_),
    .B1(net196),
    .B2(\top_inst.spi_inst.buffer[62] ),
    .A2(net203),
    .A1(\top_inst.spi_inst.buffer[61] ));
 sg13g2_inv_1 _1204_ (.Y(_0146_),
    .A(_0458_));
 sg13g2_a22oi_1 _1205_ (.Y(_0459_),
    .B1(net196),
    .B2(\top_inst.spi_inst.buffer[63] ),
    .A2(net203),
    .A1(\top_inst.spi_inst.buffer[62] ));
 sg13g2_inv_1 _1206_ (.Y(_0147_),
    .A(_0459_));
 sg13g2_dfrbp_1 _1207_ (.CLK(net228),
    .RESET_B(net30),
    .D(_0009_),
    .Q_N(_0594_),
    .Q(\top_inst.controller_inst.spi_load_next ));
 sg13g2_dfrbp_1 _1208_ (.CLK(net233),
    .RESET_B(net38),
    .D(_0010_),
    .Q_N(_0593_),
    .Q(\top_inst.data[40] ));
 sg13g2_dfrbp_1 _1209_ (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net37),
    .D(_0011_),
    .Q_N(_0008_),
    .Q(\top_inst.counter[0] ));
 sg13g2_dfrbp_1 _1210_ (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net36),
    .D(net175),
    .Q_N(_0592_),
    .Q(\top_inst.counter[1] ));
 sg13g2_dfrbp_1 _1211_ (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net35),
    .D(net173),
    .Q_N(_0591_),
    .Q(\top_inst.counter[2] ));
 sg13g2_dfrbp_1 _1212_ (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net34),
    .D(_0014_),
    .Q_N(_0590_),
    .Q(\top_inst.counter[3] ));
 sg13g2_dfrbp_1 _1213_ (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net53),
    .D(_0015_),
    .Q_N(_0595_),
    .Q(\top_inst.clk ));
 sg13g2_dfrbp_1 _1214_ (.CLK(net228),
    .RESET_B(net33),
    .D(\top_inst.controller_inst.spi_load_pending ),
    .Q_N(_0589_),
    .Q(\top_inst.controller_inst.spi_load ));
 sg13g2_dfrbp_1 _1215_ (.CLK(net229),
    .RESET_B(net32),
    .D(_0016_),
    .Q_N(_0588_),
    .Q(\top_inst.controller_inst.counter[0] ));
 sg13g2_dfrbp_1 _1216_ (.CLK(net229),
    .RESET_B(net29),
    .D(_0017_),
    .Q_N(_0587_),
    .Q(\top_inst.controller_inst.counter[1] ));
 sg13g2_dfrbp_1 _1217_ (.CLK(net230),
    .RESET_B(net27),
    .D(_0018_),
    .Q_N(_0586_),
    .Q(\top_inst.controller_inst.counter[2] ));
 sg13g2_dfrbp_1 _1218_ (.CLK(net229),
    .RESET_B(net25),
    .D(_0019_),
    .Q_N(_0585_),
    .Q(\top_inst.controller_inst.counter[3] ));
 sg13g2_dfrbp_1 _1219_ (.CLK(net225),
    .RESET_B(net23),
    .D(_0020_),
    .Q_N(_0584_),
    .Q(\top_inst.controller_inst.counter[4] ));
 sg13g2_dfrbp_1 _1220_ (.CLK(net226),
    .RESET_B(net168),
    .D(_0021_),
    .Q_N(_0583_),
    .Q(\top_inst.controller_inst.counter[5] ));
 sg13g2_dfrbp_1 _1221_ (.CLK(net226),
    .RESET_B(net166),
    .D(_0022_),
    .Q_N(_0582_),
    .Q(\top_inst.controller_inst.counter[6] ));
 sg13g2_dfrbp_1 _1222_ (.CLK(net225),
    .RESET_B(net164),
    .D(_0023_),
    .Q_N(_0581_),
    .Q(\top_inst.controller_inst.counter[7] ));
 sg13g2_dfrbp_1 _1223_ (.CLK(net225),
    .RESET_B(net162),
    .D(_0024_),
    .Q_N(_0580_),
    .Q(\top_inst.controller_inst.counter[8] ));
 sg13g2_dfrbp_1 _1224_ (.CLK(net225),
    .RESET_B(net160),
    .D(_0025_),
    .Q_N(_0579_),
    .Q(\top_inst.controller_inst.counter[9] ));
 sg13g2_dfrbp_1 _1225_ (.CLK(net225),
    .RESET_B(net158),
    .D(_0026_),
    .Q_N(_0578_),
    .Q(\top_inst.controller_inst.counter[10] ));
 sg13g2_dfrbp_1 _1226_ (.CLK(net225),
    .RESET_B(net156),
    .D(_0027_),
    .Q_N(_0577_),
    .Q(\top_inst.controller_inst.counter[11] ));
 sg13g2_dfrbp_1 _1227_ (.CLK(net225),
    .RESET_B(net154),
    .D(_0028_),
    .Q_N(_0576_),
    .Q(\top_inst.controller_inst.counter[12] ));
 sg13g2_dfrbp_1 _1228_ (.CLK(net225),
    .RESET_B(net152),
    .D(_0029_),
    .Q_N(_0575_),
    .Q(\top_inst.controller_inst.counter[13] ));
 sg13g2_dfrbp_1 _1229_ (.CLK(net224),
    .RESET_B(net150),
    .D(_0030_),
    .Q_N(_0574_),
    .Q(\top_inst.controller_inst.counter[14] ));
 sg13g2_dfrbp_1 _1230_ (.CLK(net224),
    .RESET_B(net148),
    .D(_0031_),
    .Q_N(_0573_),
    .Q(\top_inst.controller_inst.counter[15] ));
 sg13g2_dfrbp_1 _1231_ (.CLK(net224),
    .RESET_B(net146),
    .D(_0032_),
    .Q_N(_0572_),
    .Q(\top_inst.controller_inst.counter[16] ));
 sg13g2_dfrbp_1 _1232_ (.CLK(net224),
    .RESET_B(net144),
    .D(_0033_),
    .Q_N(_0571_),
    .Q(\top_inst.controller_inst.counter[17] ));
 sg13g2_dfrbp_1 _1233_ (.CLK(net224),
    .RESET_B(net142),
    .D(_0034_),
    .Q_N(_0570_),
    .Q(\top_inst.controller_inst.counter[18] ));
 sg13g2_dfrbp_1 _1234_ (.CLK(net224),
    .RESET_B(net140),
    .D(_0035_),
    .Q_N(_0569_),
    .Q(\top_inst.controller_inst.counter[19] ));
 sg13g2_dfrbp_1 _1235_ (.CLK(net224),
    .RESET_B(net138),
    .D(_0036_),
    .Q_N(_0568_),
    .Q(\top_inst.controller_inst.counter[20] ));
 sg13g2_dfrbp_1 _1236_ (.CLK(net224),
    .RESET_B(net71),
    .D(_0037_),
    .Q_N(_0596_),
    .Q(\top_inst.controller_inst.counter[21] ));
 sg13g2_dfrbp_1 _1237_ (.CLK(net228),
    .RESET_B(net136),
    .D(\top_inst.controller_inst.spi_load_next ),
    .Q_N(_0567_),
    .Q(\top_inst.controller_inst.spi_load_pending ));
 sg13g2_dfrbp_1 _1238_ (.CLK(net223),
    .RESET_B(net134),
    .D(_0038_),
    .Q_N(_0566_),
    .Q(\top_inst.address[6] ));
 sg13g2_dfrbp_1 _1239_ (.CLK(net223),
    .RESET_B(net132),
    .D(_0039_),
    .Q_N(_0565_),
    .Q(\top_inst.address[5] ));
 sg13g2_dfrbp_1 _1240_ (.CLK(net223),
    .RESET_B(net130),
    .D(_0040_),
    .Q_N(_0564_),
    .Q(\top_inst.address[4] ));
 sg13g2_dfrbp_1 _1241_ (.CLK(net223),
    .RESET_B(net128),
    .D(_0041_),
    .Q_N(_0563_),
    .Q(\top_inst.address[3] ));
 sg13g2_dfrbp_1 _1242_ (.CLK(net222),
    .RESET_B(net126),
    .D(_0042_),
    .Q_N(_0562_),
    .Q(\top_inst.address[2] ));
 sg13g2_dfrbp_1 _1243_ (.CLK(net221),
    .RESET_B(net124),
    .D(_0043_),
    .Q_N(_0561_),
    .Q(\top_inst.address[1] ));
 sg13g2_dfrbp_1 _1244_ (.CLK(net221),
    .RESET_B(net122),
    .D(_0044_),
    .Q_N(_0560_),
    .Q(\top_inst.address[0] ));
 sg13g2_dfrbp_1 _1245_ (.CLK(net227),
    .RESET_B(net120),
    .D(_0045_),
    .Q_N(_0559_),
    .Q(\top_inst.data[6] ));
 sg13g2_dfrbp_1 _1246_ (.CLK(net227),
    .RESET_B(net119),
    .D(_0046_),
    .Q_N(_0558_),
    .Q(\top_inst.data[4] ));
 sg13g2_dfrbp_1 _1247_ (.CLK(net227),
    .RESET_B(net118),
    .D(_0047_),
    .Q_N(_0557_),
    .Q(\top_inst.data[7] ));
 sg13g2_dfrbp_1 _1248_ (.CLK(net234),
    .RESET_B(net117),
    .D(_0048_),
    .Q_N(_0556_),
    .Q(\top_inst.data[41] ));
 sg13g2_dfrbp_1 _1249_ (.CLK(net236),
    .RESET_B(net116),
    .D(_0049_),
    .Q_N(_0555_),
    .Q(\top_inst.data[42] ));
 sg13g2_dfrbp_1 _1250_ (.CLK(net222),
    .RESET_B(net115),
    .D(_0050_),
    .Q_N(_0554_),
    .Q(\top_inst.data[20] ));
 sg13g2_dfrbp_1 _1251_ (.CLK(net227),
    .RESET_B(net114),
    .D(_0051_),
    .Q_N(_0553_),
    .Q(\top_inst.data[0] ));
 sg13g2_dfrbp_1 _1252_ (.CLK(net231),
    .RESET_B(net113),
    .D(_0052_),
    .Q_N(_0552_),
    .Q(\top_inst.data[12] ));
 sg13g2_dfrbp_1 _1253_ (.CLK(net232),
    .RESET_B(net112),
    .D(_0053_),
    .Q_N(_0551_),
    .Q(\top_inst.data[24] ));
 sg13g2_dfrbp_1 _1254_ (.CLK(net233),
    .RESET_B(net72),
    .D(_0054_),
    .Q_N(_0597_),
    .Q(\top_inst.data[36] ));
 sg13g2_dfrbp_1 _1255_ (.CLK(net226),
    .RESET_B(net73),
    .D(_0000_),
    .Q_N(_0598_),
    .Q(\top_inst.controller_inst.state[0] ));
 sg13g2_dfrbp_1 _1256_ (.CLK(net223),
    .RESET_B(net74),
    .D(_0001_),
    .Q_N(_0599_),
    .Q(\top_inst.controller_inst.state[1] ));
 sg13g2_dfrbp_1 _1257_ (.CLK(net223),
    .RESET_B(net82),
    .D(_0002_),
    .Q_N(_0600_),
    .Q(\top_inst.controller_inst.state[2] ));
 sg13g2_dfrbp_1 _1258_ (.CLK(net226),
    .RESET_B(net111),
    .D(_0003_),
    .Q_N(_0006_),
    .Q(\top_inst.controller_inst.state[3] ));
 sg13g2_dfrbp_1 _1259_ (.CLK(net244),
    .RESET_B(net110),
    .D(_0055_),
    .Q_N(_0007_),
    .Q(\top_inst.spi_inst.counter[0] ));
 sg13g2_dfrbp_1 _1260_ (.CLK(net244),
    .RESET_B(net109),
    .D(_0056_),
    .Q_N(_0550_),
    .Q(\top_inst.spi_inst.counter[1] ));
 sg13g2_dfrbp_1 _1261_ (.CLK(net240),
    .RESET_B(net108),
    .D(_0057_),
    .Q_N(_0549_),
    .Q(\top_inst.spi_inst.counter[2] ));
 sg13g2_dfrbp_1 _1262_ (.CLK(net240),
    .RESET_B(net107),
    .D(_0058_),
    .Q_N(_0548_),
    .Q(\top_inst.spi_inst.counter[3] ));
 sg13g2_dfrbp_1 _1263_ (.CLK(net241),
    .RESET_B(net106),
    .D(_0059_),
    .Q_N(_0547_),
    .Q(\top_inst.spi_inst.counter[4] ));
 sg13g2_dfrbp_1 _1264_ (.CLK(net240),
    .RESET_B(net105),
    .D(_0060_),
    .Q_N(_0546_),
    .Q(\top_inst.spi_inst.counter[5] ));
 sg13g2_dfrbp_1 _1265_ (.CLK(net240),
    .RESET_B(net83),
    .D(_0061_),
    .Q_N(_0601_),
    .Q(\top_inst.spi_inst.counter[6] ));
 sg13g2_dfrbp_1 _1266_ (.CLK(net240),
    .RESET_B(net102),
    .D(_0004_),
    .Q_N(_0602_),
    .Q(\top_inst.controller_inst.spi_ready ));
 sg13g2_dfrbp_1 _1267_ (.CLK(net240),
    .RESET_B(net104),
    .D(_0005_),
    .Q_N(\top_inst.spi_cs_n ),
    .Q(\top_inst.spi_inst.state[1] ));
 sg13g2_dfrbp_1 _1268_ (.CLK(net229),
    .RESET_B(net103),
    .D(_0062_),
    .Q_N(_0545_),
    .Q(\top_inst.spi_inst.buffer[0] ));
 sg13g2_dfrbp_1 _1269_ (.CLK(net222),
    .RESET_B(net101),
    .D(_0063_),
    .Q_N(_0544_),
    .Q(\top_inst.data[5] ));
 sg13g2_dfrbp_1 _1270_ (.CLK(net221),
    .RESET_B(net100),
    .D(_0064_),
    .Q_N(_0543_),
    .Q(\top_inst.data[16] ));
 sg13g2_dfrbp_1 _1271_ (.CLK(net222),
    .RESET_B(net99),
    .D(_0065_),
    .Q_N(_0542_),
    .Q(\top_inst.data[17] ));
 sg13g2_dfrbp_1 _1272_ (.CLK(net222),
    .RESET_B(net98),
    .D(_0066_),
    .Q_N(_0541_),
    .Q(\top_inst.data[18] ));
 sg13g2_dfrbp_1 _1273_ (.CLK(net231),
    .RESET_B(net97),
    .D(_0067_),
    .Q_N(_0540_),
    .Q(\top_inst.data[19] ));
 sg13g2_dfrbp_1 _1274_ (.CLK(net234),
    .RESET_B(net96),
    .D(_0068_),
    .Q_N(_0539_),
    .Q(\top_inst.data[29] ));
 sg13g2_dfrbp_1 _1275_ (.CLK(net233),
    .RESET_B(net95),
    .D(_0069_),
    .Q_N(_0538_),
    .Q(\top_inst.data[28] ));
 sg13g2_dfrbp_1 _1276_ (.CLK(net233),
    .RESET_B(net94),
    .D(_0070_),
    .Q_N(_0537_),
    .Q(\top_inst.data[11] ));
 sg13g2_dfrbp_1 _1277_ (.CLK(net234),
    .RESET_B(net93),
    .D(_0071_),
    .Q_N(_0536_),
    .Q(\top_inst.data[30] ));
 sg13g2_dfrbp_1 _1278_ (.CLK(net234),
    .RESET_B(net92),
    .D(_0072_),
    .Q_N(_0535_),
    .Q(\top_inst.data[31] ));
 sg13g2_dfrbp_1 _1279_ (.CLK(net227),
    .RESET_B(net91),
    .D(_0073_),
    .Q_N(_0534_),
    .Q(\top_inst.data[1] ));
 sg13g2_dfrbp_1 _1280_ (.CLK(net227),
    .RESET_B(net90),
    .D(_0074_),
    .Q_N(_0533_),
    .Q(\top_inst.data[2] ));
 sg13g2_dfrbp_1 _1281_ (.CLK(net231),
    .RESET_B(net89),
    .D(_0075_),
    .Q_N(_0532_),
    .Q(\top_inst.data[13] ));
 sg13g2_dfrbp_1 _1282_ (.CLK(net221),
    .RESET_B(net88),
    .D(_0076_),
    .Q_N(_0531_),
    .Q(\top_inst.data[14] ));
 sg13g2_dfrbp_1 _1283_ (.CLK(net221),
    .RESET_B(net87),
    .D(_0077_),
    .Q_N(_0530_),
    .Q(\top_inst.data[15] ));
 sg13g2_dfrbp_1 _1284_ (.CLK(net232),
    .RESET_B(net86),
    .D(_0078_),
    .Q_N(_0529_),
    .Q(\top_inst.data[25] ));
 sg13g2_dfrbp_1 _1285_ (.CLK(net231),
    .RESET_B(net85),
    .D(_0079_),
    .Q_N(_0528_),
    .Q(\top_inst.data[26] ));
 sg13g2_dfrbp_1 _1286_ (.CLK(net231),
    .RESET_B(net84),
    .D(_0080_),
    .Q_N(_0527_),
    .Q(\top_inst.data[27] ));
 sg13g2_dfrbp_1 _1287_ (.CLK(net239),
    .RESET_B(net81),
    .D(_0081_),
    .Q_N(_0526_),
    .Q(\top_inst.data[10] ));
 sg13g2_dfrbp_1 _1288_ (.CLK(net233),
    .RESET_B(net80),
    .D(_0082_),
    .Q_N(_0525_),
    .Q(\top_inst.data[37] ));
 sg13g2_dfrbp_1 _1289_ (.CLK(net233),
    .RESET_B(net79),
    .D(_0083_),
    .Q_N(_0524_),
    .Q(\top_inst.data[39] ));
 sg13g2_dfrbp_1 _1290_ (.CLK(net239),
    .RESET_B(net78),
    .D(_0084_),
    .Q_N(_0523_),
    .Q(\top_inst.data[21] ));
 sg13g2_dfrbp_1 _1291_ (.CLK(net240),
    .RESET_B(net77),
    .D(_0085_),
    .Q_N(_0522_),
    .Q(\top_inst.spi_inst.buffer[1] ));
 sg13g2_dfrbp_1 _1292_ (.CLK(net239),
    .RESET_B(net75),
    .D(_0086_),
    .Q_N(_0521_),
    .Q(\top_inst.spi_inst.buffer[2] ));
 sg13g2_dfrbp_1 _1293_ (.CLK(net239),
    .RESET_B(net69),
    .D(_0087_),
    .Q_N(_0520_),
    .Q(\top_inst.spi_inst.buffer[3] ));
 sg13g2_dfrbp_1 _1294_ (.CLK(net227),
    .RESET_B(net67),
    .D(_0088_),
    .Q_N(_0519_),
    .Q(\top_inst.spi_inst.buffer[4] ));
 sg13g2_dfrbp_1 _1295_ (.CLK(net227),
    .RESET_B(net65),
    .D(_0089_),
    .Q_N(_0518_),
    .Q(\top_inst.spi_inst.buffer[5] ));
 sg13g2_dfrbp_1 _1296_ (.CLK(net239),
    .RESET_B(net63),
    .D(_0090_),
    .Q_N(_0517_),
    .Q(\top_inst.spi_inst.buffer[6] ));
 sg13g2_dfrbp_1 _1297_ (.CLK(net239),
    .RESET_B(net61),
    .D(_0091_),
    .Q_N(_0516_),
    .Q(\top_inst.spi_inst.buffer[7] ));
 sg13g2_dfrbp_1 _1298_ (.CLK(net239),
    .RESET_B(net59),
    .D(_0092_),
    .Q_N(_0515_),
    .Q(\top_inst.spi_inst.buffer[8] ));
 sg13g2_dfrbp_1 _1299_ (.CLK(net242),
    .RESET_B(net57),
    .D(_0093_),
    .Q_N(_0514_),
    .Q(\top_inst.spi_inst.buffer[9] ));
 sg13g2_dfrbp_1 _1300_ (.CLK(net243),
    .RESET_B(net55),
    .D(_0094_),
    .Q_N(_0513_),
    .Q(\top_inst.spi_inst.buffer[10] ));
 sg13g2_dfrbp_1 _1301_ (.CLK(net243),
    .RESET_B(net52),
    .D(_0095_),
    .Q_N(_0512_),
    .Q(\top_inst.spi_inst.buffer[11] ));
 sg13g2_dfrbp_1 _1302_ (.CLK(net237),
    .RESET_B(net50),
    .D(_0096_),
    .Q_N(_0511_),
    .Q(\top_inst.spi_inst.buffer[12] ));
 sg13g2_dfrbp_1 _1303_ (.CLK(net237),
    .RESET_B(net48),
    .D(_0097_),
    .Q_N(_0510_),
    .Q(\top_inst.spi_inst.buffer[13] ));
 sg13g2_dfrbp_1 _1304_ (.CLK(net235),
    .RESET_B(net46),
    .D(_0098_),
    .Q_N(_0509_),
    .Q(\top_inst.spi_inst.buffer[14] ));
 sg13g2_dfrbp_1 _1305_ (.CLK(net235),
    .RESET_B(net44),
    .D(_0099_),
    .Q_N(_0508_),
    .Q(\top_inst.spi_inst.buffer[15] ));
 sg13g2_dfrbp_1 _1306_ (.CLK(net232),
    .RESET_B(net42),
    .D(_0100_),
    .Q_N(_0507_),
    .Q(\top_inst.spi_inst.buffer[16] ));
 sg13g2_dfrbp_1 _1307_ (.CLK(net231),
    .RESET_B(net40),
    .D(_0101_),
    .Q_N(_0506_),
    .Q(\top_inst.spi_inst.buffer[17] ));
 sg13g2_dfrbp_1 _1308_ (.CLK(net231),
    .RESET_B(net31),
    .D(_0102_),
    .Q_N(_0505_),
    .Q(\top_inst.spi_inst.buffer[18] ));
 sg13g2_dfrbp_1 _1309_ (.CLK(net221),
    .RESET_B(net26),
    .D(_0103_),
    .Q_N(_0504_),
    .Q(\top_inst.spi_inst.buffer[19] ));
 sg13g2_dfrbp_1 _1310_ (.CLK(net221),
    .RESET_B(net169),
    .D(_0104_),
    .Q_N(_0503_),
    .Q(\top_inst.spi_inst.buffer[20] ));
 sg13g2_dfrbp_1 _1311_ (.CLK(net221),
    .RESET_B(net165),
    .D(_0105_),
    .Q_N(_0502_),
    .Q(\top_inst.spi_inst.buffer[21] ));
 sg13g2_dfrbp_1 _1312_ (.CLK(net231),
    .RESET_B(net161),
    .D(_0106_),
    .Q_N(_0501_),
    .Q(\top_inst.spi_inst.buffer[22] ));
 sg13g2_dfrbp_1 _1313_ (.CLK(net232),
    .RESET_B(net157),
    .D(_0107_),
    .Q_N(_0500_),
    .Q(\top_inst.spi_inst.buffer[23] ));
 sg13g2_dfrbp_1 _1314_ (.CLK(net242),
    .RESET_B(net153),
    .D(_0108_),
    .Q_N(_0499_),
    .Q(\top_inst.spi_inst.buffer[24] ));
 sg13g2_dfrbp_1 _1315_ (.CLK(net242),
    .RESET_B(net149),
    .D(_0109_),
    .Q_N(_0498_),
    .Q(\top_inst.spi_inst.buffer[25] ));
 sg13g2_dfrbp_1 _1316_ (.CLK(net242),
    .RESET_B(net145),
    .D(_0110_),
    .Q_N(_0497_),
    .Q(\top_inst.spi_inst.buffer[26] ));
 sg13g2_dfrbp_1 _1317_ (.CLK(net243),
    .RESET_B(net141),
    .D(_0111_),
    .Q_N(_0496_),
    .Q(\top_inst.spi_inst.buffer[27] ));
 sg13g2_dfrbp_1 _1318_ (.CLK(net237),
    .RESET_B(net137),
    .D(_0112_),
    .Q_N(_0495_),
    .Q(\top_inst.spi_inst.buffer[28] ));
 sg13g2_dfrbp_1 _1319_ (.CLK(net237),
    .RESET_B(net133),
    .D(_0113_),
    .Q_N(_0494_),
    .Q(\top_inst.spi_inst.buffer[29] ));
 sg13g2_dfrbp_1 _1320_ (.CLK(net235),
    .RESET_B(net129),
    .D(_0114_),
    .Q_N(_0493_),
    .Q(\top_inst.spi_inst.buffer[30] ));
 sg13g2_dfrbp_1 _1321_ (.CLK(net235),
    .RESET_B(net125),
    .D(_0115_),
    .Q_N(_0492_),
    .Q(\top_inst.spi_inst.buffer[31] ));
 sg13g2_dfrbp_1 _1322_ (.CLK(net235),
    .RESET_B(net121),
    .D(_0116_),
    .Q_N(_0491_),
    .Q(\top_inst.spi_inst.buffer[32] ));
 sg13g2_dfrbp_1 _1323_ (.CLK(net235),
    .RESET_B(net76),
    .D(_0117_),
    .Q_N(_0490_),
    .Q(\top_inst.spi_inst.buffer[33] ));
 sg13g2_dfrbp_1 _1324_ (.CLK(net232),
    .RESET_B(net68),
    .D(_0118_),
    .Q_N(_0489_),
    .Q(\top_inst.spi_inst.buffer[34] ));
 sg13g2_dfrbp_1 _1325_ (.CLK(net232),
    .RESET_B(net64),
    .D(_0119_),
    .Q_N(_0488_),
    .Q(\top_inst.spi_inst.buffer[35] ));
 sg13g2_dfrbp_1 _1326_ (.CLK(net235),
    .RESET_B(net60),
    .D(_0120_),
    .Q_N(_0487_),
    .Q(\top_inst.spi_inst.buffer[36] ));
 sg13g2_dfrbp_1 _1327_ (.CLK(net235),
    .RESET_B(net56),
    .D(_0121_),
    .Q_N(_0486_),
    .Q(\top_inst.spi_inst.buffer[37] ));
 sg13g2_dfrbp_1 _1328_ (.CLK(net236),
    .RESET_B(net51),
    .D(_0122_),
    .Q_N(_0485_),
    .Q(\top_inst.spi_inst.buffer[38] ));
 sg13g2_dfrbp_1 _1329_ (.CLK(net236),
    .RESET_B(net47),
    .D(_0123_),
    .Q_N(_0484_),
    .Q(\top_inst.spi_inst.buffer[39] ));
 sg13g2_dfrbp_1 _1330_ (.CLK(net242),
    .RESET_B(net43),
    .D(_0124_),
    .Q_N(_0483_),
    .Q(\top_inst.spi_inst.buffer[40] ));
 sg13g2_dfrbp_1 _1331_ (.CLK(net242),
    .RESET_B(net39),
    .D(_0125_),
    .Q_N(_0482_),
    .Q(\top_inst.spi_inst.buffer[41] ));
 sg13g2_dfrbp_1 _1332_ (.CLK(net244),
    .RESET_B(net24),
    .D(_0126_),
    .Q_N(_0481_),
    .Q(\top_inst.spi_inst.buffer[42] ));
 sg13g2_dfrbp_1 _1333_ (.CLK(net244),
    .RESET_B(net163),
    .D(_0127_),
    .Q_N(_0480_),
    .Q(\top_inst.spi_inst.buffer[43] ));
 sg13g2_dfrbp_1 _1334_ (.CLK(net245),
    .RESET_B(net155),
    .D(_0128_),
    .Q_N(_0479_),
    .Q(\top_inst.spi_inst.buffer[44] ));
 sg13g2_dfrbp_1 _1335_ (.CLK(net243),
    .RESET_B(net147),
    .D(_0129_),
    .Q_N(_0478_),
    .Q(\top_inst.spi_inst.buffer[45] ));
 sg13g2_dfrbp_1 _1336_ (.CLK(net243),
    .RESET_B(net139),
    .D(_0130_),
    .Q_N(_0477_),
    .Q(\top_inst.spi_inst.buffer[46] ));
 sg13g2_dfrbp_1 _1337_ (.CLK(net236),
    .RESET_B(net131),
    .D(_0131_),
    .Q_N(_0476_),
    .Q(\top_inst.spi_inst.buffer[47] ));
 sg13g2_dfrbp_1 _1338_ (.CLK(net233),
    .RESET_B(net123),
    .D(_0132_),
    .Q_N(_0475_),
    .Q(\top_inst.spi_inst.buffer[48] ));
 sg13g2_dfrbp_1 _1339_ (.CLK(net239),
    .RESET_B(net70),
    .D(_0133_),
    .Q_N(_0474_),
    .Q(\top_inst.spi_inst.buffer[49] ));
 sg13g2_dfrbp_1 _1340_ (.CLK(net241),
    .RESET_B(net62),
    .D(_0134_),
    .Q_N(_0473_),
    .Q(\top_inst.spi_inst.buffer[50] ));
 sg13g2_dfrbp_1 _1341_ (.CLK(net233),
    .RESET_B(net54),
    .D(_0135_),
    .Q_N(_0472_),
    .Q(\top_inst.spi_inst.buffer[51] ));
 sg13g2_dfrbp_1 _1342_ (.CLK(net236),
    .RESET_B(net45),
    .D(_0136_),
    .Q_N(_0471_),
    .Q(\top_inst.spi_inst.buffer[52] ));
 sg13g2_dfrbp_1 _1343_ (.CLK(net236),
    .RESET_B(net28),
    .D(_0137_),
    .Q_N(_0470_),
    .Q(\top_inst.spi_inst.buffer[53] ));
 sg13g2_dfrbp_1 _1344_ (.CLK(net236),
    .RESET_B(net159),
    .D(_0138_),
    .Q_N(_0469_),
    .Q(\top_inst.spi_inst.buffer[54] ));
 sg13g2_dfrbp_1 _1345_ (.CLK(net236),
    .RESET_B(net143),
    .D(_0139_),
    .Q_N(_0468_),
    .Q(\top_inst.spi_inst.buffer[55] ));
 sg13g2_dfrbp_1 _1346_ (.CLK(net242),
    .RESET_B(net127),
    .D(_0140_),
    .Q_N(_0467_),
    .Q(\top_inst.spi_inst.buffer[56] ));
 sg13g2_dfrbp_1 _1347_ (.CLK(net242),
    .RESET_B(net66),
    .D(_0141_),
    .Q_N(_0466_),
    .Q(\top_inst.spi_inst.buffer[57] ));
 sg13g2_dfrbp_1 _1348_ (.CLK(net244),
    .RESET_B(net49),
    .D(_0142_),
    .Q_N(_0465_),
    .Q(\top_inst.spi_inst.buffer[58] ));
 sg13g2_dfrbp_1 _1349_ (.CLK(net241),
    .RESET_B(net167),
    .D(_0143_),
    .Q_N(_0464_),
    .Q(\top_inst.spi_inst.buffer[59] ));
 sg13g2_dfrbp_1 _1350_ (.CLK(net241),
    .RESET_B(net135),
    .D(_0144_),
    .Q_N(_0463_),
    .Q(\top_inst.spi_inst.buffer[60] ));
 sg13g2_dfrbp_1 _1351_ (.CLK(net229),
    .RESET_B(net58),
    .D(_0145_),
    .Q_N(_0462_),
    .Q(\top_inst.spi_inst.buffer[61] ));
 sg13g2_dfrbp_1 _1352_ (.CLK(net229),
    .RESET_B(net151),
    .D(_0146_),
    .Q_N(_0461_),
    .Q(\top_inst.spi_inst.buffer[62] ));
 sg13g2_dfrbp_1 _1353_ (.CLK(net229),
    .RESET_B(net41),
    .D(_0147_),
    .Q_N(_0460_),
    .Q(\top_inst.spi_inst.buffer[63] ));
 sg13g2_tiehi _1332__24 (.L_HI(net24));
 sg13g2_tiehi _1218__25 (.L_HI(net25));
 sg13g2_tiehi _1309__26 (.L_HI(net26));
 sg13g2_tiehi _1217__27 (.L_HI(net27));
 sg13g2_tiehi _1343__28 (.L_HI(net28));
 sg13g2_tiehi _1216__29 (.L_HI(net29));
 sg13g2_tiehi _1207__30 (.L_HI(net30));
 sg13g2_tiehi _1308__31 (.L_HI(net31));
 sg13g2_tiehi _1215__32 (.L_HI(net32));
 sg13g2_tiehi _1214__33 (.L_HI(net33));
 sg13g2_tiehi _1212__34 (.L_HI(net34));
 sg13g2_tiehi _1211__35 (.L_HI(net35));
 sg13g2_tiehi _1210__36 (.L_HI(net36));
 sg13g2_tiehi _1209__37 (.L_HI(net37));
 sg13g2_tiehi _1208__38 (.L_HI(net38));
 sg13g2_tiehi _1331__39 (.L_HI(net39));
 sg13g2_tiehi _1307__40 (.L_HI(net40));
 sg13g2_tiehi _1353__41 (.L_HI(net41));
 sg13g2_tiehi _1306__42 (.L_HI(net42));
 sg13g2_tiehi _1330__43 (.L_HI(net43));
 sg13g2_tiehi _1305__44 (.L_HI(net44));
 sg13g2_tiehi _1342__45 (.L_HI(net45));
 sg13g2_tiehi _1304__46 (.L_HI(net46));
 sg13g2_tiehi _1329__47 (.L_HI(net47));
 sg13g2_tiehi _1303__48 (.L_HI(net48));
 sg13g2_tiehi _1348__49 (.L_HI(net49));
 sg13g2_tiehi _1302__50 (.L_HI(net50));
 sg13g2_tiehi _1328__51 (.L_HI(net51));
 sg13g2_tiehi _1301__52 (.L_HI(net52));
 sg13g2_tiehi _1213__53 (.L_HI(net53));
 sg13g2_tiehi _1341__54 (.L_HI(net54));
 sg13g2_tiehi _1300__55 (.L_HI(net55));
 sg13g2_tiehi _1327__56 (.L_HI(net56));
 sg13g2_tiehi _1299__57 (.L_HI(net57));
 sg13g2_tiehi _1351__58 (.L_HI(net58));
 sg13g2_tiehi _1298__59 (.L_HI(net59));
 sg13g2_tiehi _1326__60 (.L_HI(net60));
 sg13g2_tiehi _1297__61 (.L_HI(net61));
 sg13g2_tiehi _1340__62 (.L_HI(net62));
 sg13g2_tiehi _1296__63 (.L_HI(net63));
 sg13g2_tiehi _1325__64 (.L_HI(net64));
 sg13g2_tiehi _1295__65 (.L_HI(net65));
 sg13g2_tiehi _1347__66 (.L_HI(net66));
 sg13g2_tiehi _1294__67 (.L_HI(net67));
 sg13g2_tiehi _1324__68 (.L_HI(net68));
 sg13g2_tiehi _1293__69 (.L_HI(net69));
 sg13g2_tiehi _1339__70 (.L_HI(net70));
 sg13g2_tiehi _1236__71 (.L_HI(net71));
 sg13g2_tiehi _1254__72 (.L_HI(net72));
 sg13g2_tiehi _1255__73 (.L_HI(net73));
 sg13g2_tiehi _1256__74 (.L_HI(net74));
 sg13g2_tiehi _1292__75 (.L_HI(net75));
 sg13g2_tiehi _1323__76 (.L_HI(net76));
 sg13g2_tiehi _1291__77 (.L_HI(net77));
 sg13g2_tiehi _1290__78 (.L_HI(net78));
 sg13g2_tiehi _1289__79 (.L_HI(net79));
 sg13g2_tiehi _1288__80 (.L_HI(net80));
 sg13g2_tiehi _1287__81 (.L_HI(net81));
 sg13g2_tiehi _1257__82 (.L_HI(net82));
 sg13g2_tiehi _1265__83 (.L_HI(net83));
 sg13g2_tiehi _1286__84 (.L_HI(net84));
 sg13g2_tiehi _1285__85 (.L_HI(net85));
 sg13g2_tiehi _1284__86 (.L_HI(net86));
 sg13g2_tiehi _1283__87 (.L_HI(net87));
 sg13g2_tiehi _1282__88 (.L_HI(net88));
 sg13g2_tiehi _1281__89 (.L_HI(net89));
 sg13g2_tiehi _1280__90 (.L_HI(net90));
 sg13g2_tiehi _1279__91 (.L_HI(net91));
 sg13g2_tiehi _1278__92 (.L_HI(net92));
 sg13g2_tiehi _1277__93 (.L_HI(net93));
 sg13g2_tiehi _1276__94 (.L_HI(net94));
 sg13g2_tiehi _1275__95 (.L_HI(net95));
 sg13g2_tiehi _1274__96 (.L_HI(net96));
 sg13g2_tiehi _1273__97 (.L_HI(net97));
 sg13g2_tiehi _1272__98 (.L_HI(net98));
 sg13g2_tiehi _1271__99 (.L_HI(net99));
 sg13g2_tiehi _1270__100 (.L_HI(net100));
 sg13g2_tiehi _1269__101 (.L_HI(net101));
 sg13g2_tiehi _1266__102 (.L_HI(net102));
 sg13g2_tiehi _1268__103 (.L_HI(net103));
 sg13g2_tiehi _1267__104 (.L_HI(net104));
 sg13g2_tiehi _1264__105 (.L_HI(net105));
 sg13g2_tiehi _1263__106 (.L_HI(net106));
 sg13g2_tiehi _1262__107 (.L_HI(net107));
 sg13g2_tiehi _1261__108 (.L_HI(net108));
 sg13g2_tiehi _1260__109 (.L_HI(net109));
 sg13g2_tiehi _1259__110 (.L_HI(net110));
 sg13g2_tiehi _1258__111 (.L_HI(net111));
 sg13g2_tiehi _1253__112 (.L_HI(net112));
 sg13g2_tiehi _1252__113 (.L_HI(net113));
 sg13g2_tiehi _1251__114 (.L_HI(net114));
 sg13g2_tiehi _1250__115 (.L_HI(net115));
 sg13g2_tiehi _1249__116 (.L_HI(net116));
 sg13g2_tiehi _1248__117 (.L_HI(net117));
 sg13g2_tiehi _1247__118 (.L_HI(net118));
 sg13g2_tiehi _1246__119 (.L_HI(net119));
 sg13g2_tiehi _1245__120 (.L_HI(net120));
 sg13g2_tiehi _1322__121 (.L_HI(net121));
 sg13g2_tiehi _1244__122 (.L_HI(net122));
 sg13g2_tiehi _1338__123 (.L_HI(net123));
 sg13g2_tiehi _1243__124 (.L_HI(net124));
 sg13g2_tiehi _1321__125 (.L_HI(net125));
 sg13g2_tiehi _1242__126 (.L_HI(net126));
 sg13g2_tiehi _1346__127 (.L_HI(net127));
 sg13g2_tiehi _1241__128 (.L_HI(net128));
 sg13g2_tiehi _1320__129 (.L_HI(net129));
 sg13g2_tiehi _1240__130 (.L_HI(net130));
 sg13g2_tiehi _1337__131 (.L_HI(net131));
 sg13g2_tiehi _1239__132 (.L_HI(net132));
 sg13g2_tiehi _1319__133 (.L_HI(net133));
 sg13g2_tiehi _1238__134 (.L_HI(net134));
 sg13g2_tiehi _1350__135 (.L_HI(net135));
 sg13g2_tiehi _1237__136 (.L_HI(net136));
 sg13g2_tiehi _1318__137 (.L_HI(net137));
 sg13g2_tiehi _1235__138 (.L_HI(net138));
 sg13g2_tiehi _1336__139 (.L_HI(net139));
 sg13g2_tiehi _1234__140 (.L_HI(net140));
 sg13g2_tiehi _1317__141 (.L_HI(net141));
 sg13g2_tiehi _1233__142 (.L_HI(net142));
 sg13g2_tiehi _1345__143 (.L_HI(net143));
 sg13g2_tiehi _1232__144 (.L_HI(net144));
 sg13g2_tiehi _1316__145 (.L_HI(net145));
 sg13g2_tiehi _1231__146 (.L_HI(net146));
 sg13g2_tiehi _1335__147 (.L_HI(net147));
 sg13g2_tiehi _1230__148 (.L_HI(net148));
 sg13g2_tiehi _1315__149 (.L_HI(net149));
 sg13g2_tiehi _1229__150 (.L_HI(net150));
 sg13g2_tiehi _1352__151 (.L_HI(net151));
 sg13g2_tiehi _1228__152 (.L_HI(net152));
 sg13g2_tiehi _1314__153 (.L_HI(net153));
 sg13g2_tiehi _1227__154 (.L_HI(net154));
 sg13g2_tiehi _1334__155 (.L_HI(net155));
 sg13g2_tiehi _1226__156 (.L_HI(net156));
 sg13g2_tiehi _1313__157 (.L_HI(net157));
 sg13g2_tiehi _1225__158 (.L_HI(net158));
 sg13g2_tiehi _1344__159 (.L_HI(net159));
 sg13g2_tiehi _1224__160 (.L_HI(net160));
 sg13g2_tiehi _1312__161 (.L_HI(net161));
 sg13g2_tiehi _1223__162 (.L_HI(net162));
 sg13g2_tiehi _1333__163 (.L_HI(net163));
 sg13g2_tiehi _1222__164 (.L_HI(net164));
 sg13g2_tiehi _1311__165 (.L_HI(net165));
 sg13g2_tiehi _1221__166 (.L_HI(net166));
 sg13g2_tiehi _1349__167 (.L_HI(net167));
 sg13g2_tiehi _1220__168 (.L_HI(net168));
 sg13g2_tiehi _1310__169 (.L_HI(net169));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_3 (.L_LO(net3));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_4 (.L_LO(net4));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_5 (.L_LO(net5));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_6 (.L_LO(net6));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_7 (.L_LO(net7));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_8 (.L_LO(net8));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_9 (.L_LO(net9));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_10 (.L_LO(net10));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_11 (.L_LO(net11));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_12 (.L_LO(net12));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_13 (.L_LO(net13));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_14 (.L_LO(net14));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_15 (.L_LO(net15));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_16 (.L_LO(net16));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_17 (.L_LO(net17));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_18 (.L_LO(net18));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_19 (.L_LO(net19));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_20 (.L_LO(net20));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_21 (.L_LO(net21));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_22 (.L_LO(net22));
 sg13g2_tiehi _1219__23 (.L_HI(net23));
 sg13g2_buf_1 _1522_ (.A(net240),
    .X(uo_out[0]));
 sg13g2_buf_1 _1523_ (.A(\top_inst.spi_cs_n ),
    .X(uo_out[1]));
 sg13g2_buf_1 _1524_ (.A(\top_inst.spi_inst.buffer[63] ),
    .X(uo_out[2]));
 sg13g2_buf_2 fanout189 (.A(net190),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_0272_),
    .X(net190));
 sg13g2_buf_4 fanout191 (.X(net191),
    .A(net194));
 sg13g2_buf_1 fanout192 (.A(net194),
    .X(net192));
 sg13g2_buf_4 fanout193 (.X(net193),
    .A(net194));
 sg13g2_buf_2 fanout194 (.A(net195),
    .X(net194));
 sg13g2_buf_4 fanout195 (.X(net195),
    .A(_0372_));
 sg13g2_buf_4 fanout196 (.X(net196),
    .A(net197));
 sg13g2_buf_4 fanout197 (.X(net197),
    .A(_0372_));
 sg13g2_buf_2 fanout198 (.A(net201),
    .X(net198));
 sg13g2_buf_1 fanout199 (.A(net201),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(net201),
    .X(net200));
 sg13g2_buf_1 fanout201 (.A(net202),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_0371_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(net204),
    .X(net203));
 sg13g2_buf_4 fanout204 (.X(net204),
    .A(_0371_));
 sg13g2_buf_2 fanout205 (.A(net208),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(net207),
    .X(net206));
 sg13g2_buf_4 fanout207 (.X(net207),
    .A(net208));
 sg13g2_buf_4 fanout208 (.X(net208),
    .A(_0238_));
 sg13g2_buf_2 fanout209 (.A(net210),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_0236_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_0236_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_0235_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(net216),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(net216),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(net216),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(\top_inst.spi_inst.state[1] ),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(net219),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(net219),
    .X(net218));
 sg13g2_buf_4 fanout219 (.X(net219),
    .A(\top_inst.controller_inst.spi_ready ));
 sg13g2_buf_4 fanout220 (.X(net220),
    .A(\top_inst.address[1] ));
 sg13g2_buf_2 fanout221 (.A(net222),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(net223),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(net230),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(net226),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(net226),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(net230),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(net228),
    .X(net227));
 sg13g2_buf_1 fanout228 (.A(net229),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(net230),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(\top_inst.clk ),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(net232),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(net238),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(net238),
    .X(net233));
 sg13g2_buf_1 fanout234 (.A(net238),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(net237),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(net237),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(net238),
    .X(net237));
 sg13g2_buf_1 fanout238 (.A(net245),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(net241),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(net241),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(net245),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(net244),
    .X(net242));
 sg13g2_buf_1 fanout243 (.A(net244),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(net245),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(\top_inst.clk ),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_0205_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(net248),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(rst_n),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(net251),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(net251),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(rst_n),
    .X(net251));
 sg13g2_buf_2 input1 (.A(ena),
    .X(net1));
 sg13g2_tielo tt_um_led_matrix_ayla_lin_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0008_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold2 (.A(\top_inst.counter[2] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0261_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0013_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold5 (.A(\top_inst.counter[0] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0012_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold7 (.A(\top_inst.counter[3] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0265_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold9 (.A(\top_inst.counter[1] ),
    .X(net178));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_fill_1 FILLER_10_164 ();
 sg13g2_decap_4 FILLER_10_170 ();
 sg13g2_fill_1 FILLER_10_174 ();
 sg13g2_decap_8 FILLER_10_179 ();
 sg13g2_decap_8 FILLER_10_186 ();
 sg13g2_decap_8 FILLER_10_193 ();
 sg13g2_decap_8 FILLER_10_200 ();
 sg13g2_decap_8 FILLER_10_207 ();
 sg13g2_decap_8 FILLER_10_214 ();
 sg13g2_decap_8 FILLER_10_221 ();
 sg13g2_decap_8 FILLER_10_228 ();
 sg13g2_fill_1 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_244 ();
 sg13g2_decap_8 FILLER_10_251 ();
 sg13g2_decap_8 FILLER_10_258 ();
 sg13g2_decap_8 FILLER_10_265 ();
 sg13g2_decap_8 FILLER_10_272 ();
 sg13g2_decap_8 FILLER_10_279 ();
 sg13g2_decap_8 FILLER_10_286 ();
 sg13g2_decap_8 FILLER_10_293 ();
 sg13g2_decap_8 FILLER_10_300 ();
 sg13g2_decap_8 FILLER_10_307 ();
 sg13g2_decap_8 FILLER_10_314 ();
 sg13g2_decap_8 FILLER_10_321 ();
 sg13g2_decap_8 FILLER_10_328 ();
 sg13g2_decap_8 FILLER_10_335 ();
 sg13g2_decap_8 FILLER_10_342 ();
 sg13g2_decap_8 FILLER_10_349 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_decap_8 FILLER_10_363 ();
 sg13g2_decap_8 FILLER_10_370 ();
 sg13g2_decap_8 FILLER_10_377 ();
 sg13g2_decap_8 FILLER_10_384 ();
 sg13g2_decap_8 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_398 ();
 sg13g2_decap_4 FILLER_10_405 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_4 FILLER_11_126 ();
 sg13g2_fill_2 FILLER_11_130 ();
 sg13g2_decap_8 FILLER_11_262 ();
 sg13g2_fill_2 FILLER_11_269 ();
 sg13g2_decap_8 FILLER_11_275 ();
 sg13g2_decap_8 FILLER_11_282 ();
 sg13g2_decap_8 FILLER_11_289 ();
 sg13g2_decap_8 FILLER_11_296 ();
 sg13g2_decap_8 FILLER_11_303 ();
 sg13g2_decap_8 FILLER_11_310 ();
 sg13g2_decap_8 FILLER_11_317 ();
 sg13g2_decap_8 FILLER_11_324 ();
 sg13g2_decap_8 FILLER_11_331 ();
 sg13g2_decap_8 FILLER_11_338 ();
 sg13g2_decap_8 FILLER_11_345 ();
 sg13g2_decap_8 FILLER_11_352 ();
 sg13g2_decap_8 FILLER_11_359 ();
 sg13g2_decap_8 FILLER_11_366 ();
 sg13g2_decap_8 FILLER_11_373 ();
 sg13g2_decap_8 FILLER_11_380 ();
 sg13g2_decap_8 FILLER_11_387 ();
 sg13g2_decap_8 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_4 FILLER_12_140 ();
 sg13g2_fill_2 FILLER_12_144 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_fill_2 FILLER_12_161 ();
 sg13g2_fill_1 FILLER_12_163 ();
 sg13g2_decap_4 FILLER_12_172 ();
 sg13g2_decap_8 FILLER_12_180 ();
 sg13g2_fill_2 FILLER_12_187 ();
 sg13g2_fill_1 FILLER_12_189 ();
 sg13g2_fill_2 FILLER_12_201 ();
 sg13g2_fill_1 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_214 ();
 sg13g2_fill_2 FILLER_12_225 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_4 FILLER_12_245 ();
 sg13g2_fill_1 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_286 ();
 sg13g2_decap_4 FILLER_12_293 ();
 sg13g2_fill_1 FILLER_12_297 ();
 sg13g2_decap_8 FILLER_12_324 ();
 sg13g2_decap_8 FILLER_12_331 ();
 sg13g2_decap_8 FILLER_12_338 ();
 sg13g2_decap_8 FILLER_12_345 ();
 sg13g2_decap_8 FILLER_12_352 ();
 sg13g2_decap_8 FILLER_12_359 ();
 sg13g2_decap_8 FILLER_12_366 ();
 sg13g2_decap_4 FILLER_12_373 ();
 sg13g2_fill_1 FILLER_12_377 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_4 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_fill_2 FILLER_13_133 ();
 sg13g2_decap_4 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_197 ();
 sg13g2_decap_4 FILLER_13_204 ();
 sg13g2_fill_1 FILLER_13_208 ();
 sg13g2_fill_2 FILLER_13_214 ();
 sg13g2_fill_1 FILLER_13_247 ();
 sg13g2_decap_8 FILLER_13_251 ();
 sg13g2_fill_1 FILLER_13_258 ();
 sg13g2_fill_2 FILLER_13_264 ();
 sg13g2_fill_1 FILLER_13_266 ();
 sg13g2_decap_4 FILLER_13_304 ();
 sg13g2_fill_1 FILLER_13_308 ();
 sg13g2_fill_2 FILLER_13_318 ();
 sg13g2_fill_1 FILLER_13_320 ();
 sg13g2_decap_4 FILLER_13_325 ();
 sg13g2_fill_2 FILLER_13_329 ();
 sg13g2_decap_4 FILLER_13_360 ();
 sg13g2_fill_1 FILLER_13_393 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_fill_2 FILLER_14_126 ();
 sg13g2_fill_1 FILLER_14_128 ();
 sg13g2_fill_1 FILLER_14_155 ();
 sg13g2_fill_1 FILLER_14_159 ();
 sg13g2_fill_1 FILLER_14_191 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_fill_1 FILLER_14_231 ();
 sg13g2_fill_1 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_270 ();
 sg13g2_fill_1 FILLER_14_277 ();
 sg13g2_decap_4 FILLER_14_286 ();
 sg13g2_fill_2 FILLER_14_290 ();
 sg13g2_fill_2 FILLER_14_301 ();
 sg13g2_fill_1 FILLER_14_303 ();
 sg13g2_fill_1 FILLER_14_348 ();
 sg13g2_fill_2 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_fill_2 FILLER_15_126 ();
 sg13g2_fill_1 FILLER_15_128 ();
 sg13g2_decap_4 FILLER_15_134 ();
 sg13g2_fill_1 FILLER_15_138 ();
 sg13g2_decap_4 FILLER_15_143 ();
 sg13g2_fill_1 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_152 ();
 sg13g2_decap_8 FILLER_15_167 ();
 sg13g2_fill_2 FILLER_15_174 ();
 sg13g2_decap_4 FILLER_15_180 ();
 sg13g2_fill_2 FILLER_15_184 ();
 sg13g2_decap_8 FILLER_15_200 ();
 sg13g2_fill_2 FILLER_15_207 ();
 sg13g2_decap_8 FILLER_15_213 ();
 sg13g2_fill_2 FILLER_15_220 ();
 sg13g2_fill_2 FILLER_15_225 ();
 sg13g2_fill_1 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_237 ();
 sg13g2_decap_4 FILLER_15_244 ();
 sg13g2_fill_2 FILLER_15_248 ();
 sg13g2_decap_4 FILLER_15_257 ();
 sg13g2_fill_1 FILLER_15_261 ();
 sg13g2_decap_4 FILLER_15_299 ();
 sg13g2_decap_8 FILLER_15_306 ();
 sg13g2_decap_4 FILLER_15_313 ();
 sg13g2_decap_8 FILLER_15_323 ();
 sg13g2_decap_8 FILLER_15_330 ();
 sg13g2_fill_2 FILLER_15_337 ();
 sg13g2_fill_2 FILLER_15_353 ();
 sg13g2_fill_2 FILLER_15_358 ();
 sg13g2_fill_1 FILLER_15_368 ();
 sg13g2_fill_1 FILLER_15_375 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_fill_2 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_4 FILLER_16_98 ();
 sg13g2_fill_2 FILLER_16_102 ();
 sg13g2_fill_1 FILLER_16_108 ();
 sg13g2_fill_2 FILLER_16_135 ();
 sg13g2_fill_1 FILLER_16_163 ();
 sg13g2_decap_8 FILLER_16_246 ();
 sg13g2_decap_4 FILLER_16_253 ();
 sg13g2_decap_8 FILLER_16_264 ();
 sg13g2_decap_8 FILLER_16_276 ();
 sg13g2_fill_1 FILLER_16_283 ();
 sg13g2_fill_2 FILLER_16_359 ();
 sg13g2_fill_2 FILLER_16_367 ();
 sg13g2_fill_1 FILLER_16_369 ();
 sg13g2_fill_2 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_fill_2 FILLER_17_91 ();
 sg13g2_fill_1 FILLER_17_119 ();
 sg13g2_decap_4 FILLER_17_124 ();
 sg13g2_fill_2 FILLER_17_128 ();
 sg13g2_decap_8 FILLER_17_136 ();
 sg13g2_fill_2 FILLER_17_152 ();
 sg13g2_fill_1 FILLER_17_154 ();
 sg13g2_fill_2 FILLER_17_162 ();
 sg13g2_fill_1 FILLER_17_164 ();
 sg13g2_decap_4 FILLER_17_169 ();
 sg13g2_fill_2 FILLER_17_173 ();
 sg13g2_decap_8 FILLER_17_179 ();
 sg13g2_decap_8 FILLER_17_186 ();
 sg13g2_fill_1 FILLER_17_193 ();
 sg13g2_fill_1 FILLER_17_198 ();
 sg13g2_decap_8 FILLER_17_213 ();
 sg13g2_decap_8 FILLER_17_220 ();
 sg13g2_fill_1 FILLER_17_305 ();
 sg13g2_decap_4 FILLER_17_310 ();
 sg13g2_decap_8 FILLER_17_319 ();
 sg13g2_fill_2 FILLER_17_326 ();
 sg13g2_decap_8 FILLER_17_332 ();
 sg13g2_fill_2 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_383 ();
 sg13g2_fill_2 FILLER_17_390 ();
 sg13g2_fill_1 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_4 FILLER_18_84 ();
 sg13g2_fill_1 FILLER_18_88 ();
 sg13g2_fill_1 FILLER_18_102 ();
 sg13g2_fill_1 FILLER_18_120 ();
 sg13g2_fill_1 FILLER_18_127 ();
 sg13g2_decap_4 FILLER_18_142 ();
 sg13g2_fill_1 FILLER_18_146 ();
 sg13g2_decap_4 FILLER_18_175 ();
 sg13g2_fill_2 FILLER_18_179 ();
 sg13g2_fill_2 FILLER_18_220 ();
 sg13g2_fill_2 FILLER_18_227 ();
 sg13g2_fill_1 FILLER_18_229 ();
 sg13g2_decap_4 FILLER_18_256 ();
 sg13g2_fill_2 FILLER_18_260 ();
 sg13g2_decap_4 FILLER_18_270 ();
 sg13g2_fill_2 FILLER_18_274 ();
 sg13g2_fill_2 FILLER_18_281 ();
 sg13g2_fill_2 FILLER_18_287 ();
 sg13g2_fill_1 FILLER_18_289 ();
 sg13g2_decap_8 FILLER_18_319 ();
 sg13g2_decap_4 FILLER_18_326 ();
 sg13g2_fill_2 FILLER_18_334 ();
 sg13g2_decap_8 FILLER_18_342 ();
 sg13g2_decap_4 FILLER_18_349 ();
 sg13g2_fill_1 FILLER_18_353 ();
 sg13g2_fill_2 FILLER_18_362 ();
 sg13g2_fill_1 FILLER_18_364 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_4 FILLER_19_56 ();
 sg13g2_fill_1 FILLER_19_60 ();
 sg13g2_fill_1 FILLER_19_87 ();
 sg13g2_fill_2 FILLER_19_97 ();
 sg13g2_fill_1 FILLER_19_99 ();
 sg13g2_fill_1 FILLER_19_105 ();
 sg13g2_fill_2 FILLER_19_111 ();
 sg13g2_decap_4 FILLER_19_117 ();
 sg13g2_fill_1 FILLER_19_121 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_fill_1 FILLER_19_140 ();
 sg13g2_fill_1 FILLER_19_150 ();
 sg13g2_fill_2 FILLER_19_157 ();
 sg13g2_decap_4 FILLER_19_173 ();
 sg13g2_fill_1 FILLER_19_177 ();
 sg13g2_fill_2 FILLER_19_206 ();
 sg13g2_fill_1 FILLER_19_208 ();
 sg13g2_decap_8 FILLER_19_230 ();
 sg13g2_fill_1 FILLER_19_237 ();
 sg13g2_fill_2 FILLER_19_250 ();
 sg13g2_fill_1 FILLER_19_252 ();
 sg13g2_fill_1 FILLER_19_313 ();
 sg13g2_fill_2 FILLER_19_345 ();
 sg13g2_fill_1 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_fill_2 FILLER_20_70 ();
 sg13g2_decap_4 FILLER_20_76 ();
 sg13g2_decap_4 FILLER_20_97 ();
 sg13g2_fill_2 FILLER_20_101 ();
 sg13g2_fill_2 FILLER_20_114 ();
 sg13g2_fill_1 FILLER_20_116 ();
 sg13g2_fill_1 FILLER_20_186 ();
 sg13g2_decap_8 FILLER_20_193 ();
 sg13g2_decap_8 FILLER_20_200 ();
 sg13g2_decap_4 FILLER_20_217 ();
 sg13g2_fill_2 FILLER_20_234 ();
 sg13g2_fill_1 FILLER_20_236 ();
 sg13g2_fill_1 FILLER_20_250 ();
 sg13g2_decap_4 FILLER_20_277 ();
 sg13g2_decap_8 FILLER_20_284 ();
 sg13g2_fill_1 FILLER_20_291 ();
 sg13g2_decap_8 FILLER_20_352 ();
 sg13g2_decap_8 FILLER_20_363 ();
 sg13g2_decap_4 FILLER_20_370 ();
 sg13g2_decap_8 FILLER_20_382 ();
 sg13g2_decap_4 FILLER_20_389 ();
 sg13g2_fill_1 FILLER_20_393 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_4 FILLER_21_42 ();
 sg13g2_fill_1 FILLER_21_46 ();
 sg13g2_fill_2 FILLER_21_73 ();
 sg13g2_fill_1 FILLER_21_84 ();
 sg13g2_fill_1 FILLER_21_105 ();
 sg13g2_fill_2 FILLER_21_110 ();
 sg13g2_fill_1 FILLER_21_123 ();
 sg13g2_fill_1 FILLER_21_129 ();
 sg13g2_decap_8 FILLER_21_135 ();
 sg13g2_decap_4 FILLER_21_142 ();
 sg13g2_fill_2 FILLER_21_151 ();
 sg13g2_fill_1 FILLER_21_153 ();
 sg13g2_fill_2 FILLER_21_164 ();
 sg13g2_decap_8 FILLER_21_170 ();
 sg13g2_decap_8 FILLER_21_177 ();
 sg13g2_fill_2 FILLER_21_184 ();
 sg13g2_decap_4 FILLER_21_190 ();
 sg13g2_decap_8 FILLER_21_201 ();
 sg13g2_fill_2 FILLER_21_208 ();
 sg13g2_fill_2 FILLER_21_262 ();
 sg13g2_decap_8 FILLER_21_268 ();
 sg13g2_fill_1 FILLER_21_278 ();
 sg13g2_decap_8 FILLER_21_313 ();
 sg13g2_decap_8 FILLER_21_320 ();
 sg13g2_decap_4 FILLER_21_327 ();
 sg13g2_decap_4 FILLER_21_350 ();
 sg13g2_fill_1 FILLER_21_354 ();
 sg13g2_decap_4 FILLER_21_366 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_fill_2 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_66 ();
 sg13g2_decap_8 FILLER_22_73 ();
 sg13g2_fill_2 FILLER_22_121 ();
 sg13g2_fill_2 FILLER_22_201 ();
 sg13g2_decap_8 FILLER_22_229 ();
 sg13g2_fill_2 FILLER_22_236 ();
 sg13g2_fill_1 FILLER_22_238 ();
 sg13g2_decap_4 FILLER_22_242 ();
 sg13g2_fill_1 FILLER_22_246 ();
 sg13g2_decap_8 FILLER_22_251 ();
 sg13g2_decap_4 FILLER_22_258 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_fill_2 FILLER_22_273 ();
 sg13g2_fill_1 FILLER_22_275 ();
 sg13g2_decap_8 FILLER_22_284 ();
 sg13g2_fill_2 FILLER_22_291 ();
 sg13g2_fill_1 FILLER_22_293 ();
 sg13g2_decap_8 FILLER_22_298 ();
 sg13g2_decap_8 FILLER_22_305 ();
 sg13g2_decap_8 FILLER_22_346 ();
 sg13g2_fill_1 FILLER_22_353 ();
 sg13g2_fill_2 FILLER_22_389 ();
 sg13g2_fill_1 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_4 FILLER_23_42 ();
 sg13g2_fill_2 FILLER_23_46 ();
 sg13g2_fill_2 FILLER_23_74 ();
 sg13g2_fill_1 FILLER_23_76 ();
 sg13g2_decap_4 FILLER_23_84 ();
 sg13g2_decap_4 FILLER_23_104 ();
 sg13g2_decap_8 FILLER_23_121 ();
 sg13g2_decap_8 FILLER_23_128 ();
 sg13g2_fill_1 FILLER_23_135 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_fill_2 FILLER_23_147 ();
 sg13g2_fill_1 FILLER_23_149 ();
 sg13g2_decap_8 FILLER_23_155 ();
 sg13g2_decap_4 FILLER_23_162 ();
 sg13g2_fill_1 FILLER_23_166 ();
 sg13g2_decap_8 FILLER_23_171 ();
 sg13g2_fill_1 FILLER_23_178 ();
 sg13g2_decap_8 FILLER_23_190 ();
 sg13g2_decap_8 FILLER_23_197 ();
 sg13g2_decap_4 FILLER_23_204 ();
 sg13g2_fill_2 FILLER_23_208 ();
 sg13g2_fill_2 FILLER_23_240 ();
 sg13g2_fill_1 FILLER_23_242 ();
 sg13g2_decap_8 FILLER_23_274 ();
 sg13g2_decap_8 FILLER_23_307 ();
 sg13g2_fill_2 FILLER_23_314 ();
 sg13g2_fill_1 FILLER_23_316 ();
 sg13g2_decap_8 FILLER_23_321 ();
 sg13g2_fill_2 FILLER_23_328 ();
 sg13g2_fill_1 FILLER_23_330 ();
 sg13g2_decap_4 FILLER_23_335 ();
 sg13g2_decap_4 FILLER_23_343 ();
 sg13g2_fill_1 FILLER_23_347 ();
 sg13g2_decap_4 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_369 ();
 sg13g2_decap_4 FILLER_23_376 ();
 sg13g2_fill_2 FILLER_23_380 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_4 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_72 ();
 sg13g2_fill_1 FILLER_24_102 ();
 sg13g2_fill_2 FILLER_24_120 ();
 sg13g2_fill_2 FILLER_24_148 ();
 sg13g2_fill_2 FILLER_24_176 ();
 sg13g2_decap_4 FILLER_24_204 ();
 sg13g2_decap_4 FILLER_24_220 ();
 sg13g2_fill_1 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_229 ();
 sg13g2_fill_2 FILLER_24_236 ();
 sg13g2_fill_1 FILLER_24_238 ();
 sg13g2_decap_4 FILLER_24_243 ();
 sg13g2_fill_2 FILLER_24_247 ();
 sg13g2_fill_2 FILLER_24_255 ();
 sg13g2_fill_1 FILLER_24_257 ();
 sg13g2_decap_4 FILLER_24_262 ();
 sg13g2_fill_1 FILLER_24_266 ();
 sg13g2_fill_2 FILLER_24_275 ();
 sg13g2_fill_1 FILLER_24_277 ();
 sg13g2_decap_8 FILLER_24_283 ();
 sg13g2_fill_1 FILLER_24_290 ();
 sg13g2_decap_8 FILLER_24_295 ();
 sg13g2_decap_4 FILLER_24_302 ();
 sg13g2_decap_4 FILLER_24_332 ();
 sg13g2_decap_4 FILLER_24_346 ();
 sg13g2_decap_8 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_fill_1 FILLER_25_56 ();
 sg13g2_fill_2 FILLER_25_61 ();
 sg13g2_fill_1 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_95 ();
 sg13g2_decap_4 FILLER_25_102 ();
 sg13g2_fill_2 FILLER_25_106 ();
 sg13g2_decap_4 FILLER_25_126 ();
 sg13g2_fill_2 FILLER_25_130 ();
 sg13g2_decap_8 FILLER_25_136 ();
 sg13g2_decap_8 FILLER_25_143 ();
 sg13g2_decap_8 FILLER_25_150 ();
 sg13g2_decap_4 FILLER_25_157 ();
 sg13g2_decap_8 FILLER_25_169 ();
 sg13g2_decap_8 FILLER_25_176 ();
 sg13g2_decap_4 FILLER_25_183 ();
 sg13g2_fill_2 FILLER_25_226 ();
 sg13g2_decap_4 FILLER_25_254 ();
 sg13g2_fill_1 FILLER_25_258 ();
 sg13g2_decap_8 FILLER_25_267 ();
 sg13g2_fill_1 FILLER_25_274 ();
 sg13g2_fill_2 FILLER_25_315 ();
 sg13g2_fill_1 FILLER_25_317 ();
 sg13g2_fill_2 FILLER_25_344 ();
 sg13g2_decap_8 FILLER_25_356 ();
 sg13g2_decap_8 FILLER_25_372 ();
 sg13g2_decap_4 FILLER_25_379 ();
 sg13g2_fill_1 FILLER_25_387 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_34 ();
 sg13g2_decap_8 FILLER_26_65 ();
 sg13g2_fill_2 FILLER_26_72 ();
 sg13g2_fill_1 FILLER_26_74 ();
 sg13g2_decap_4 FILLER_26_79 ();
 sg13g2_fill_1 FILLER_26_83 ();
 sg13g2_fill_2 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_122 ();
 sg13g2_decap_4 FILLER_26_129 ();
 sg13g2_decap_4 FILLER_26_184 ();
 sg13g2_fill_2 FILLER_26_225 ();
 sg13g2_decap_8 FILLER_26_239 ();
 sg13g2_decap_4 FILLER_26_246 ();
 sg13g2_decap_4 FILLER_26_295 ();
 sg13g2_fill_1 FILLER_26_299 ();
 sg13g2_decap_4 FILLER_26_304 ();
 sg13g2_fill_2 FILLER_26_308 ();
 sg13g2_fill_2 FILLER_26_333 ();
 sg13g2_fill_2 FILLER_26_344 ();
 sg13g2_decap_8 FILLER_26_398 ();
 sg13g2_decap_4 FILLER_26_405 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_66 ();
 sg13g2_fill_2 FILLER_27_73 ();
 sg13g2_fill_1 FILLER_27_75 ();
 sg13g2_decap_8 FILLER_27_93 ();
 sg13g2_decap_8 FILLER_27_100 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_fill_1 FILLER_27_119 ();
 sg13g2_decap_4 FILLER_27_146 ();
 sg13g2_fill_2 FILLER_27_150 ();
 sg13g2_fill_2 FILLER_27_186 ();
 sg13g2_fill_1 FILLER_27_188 ();
 sg13g2_decap_8 FILLER_27_193 ();
 sg13g2_fill_2 FILLER_27_200 ();
 sg13g2_fill_1 FILLER_27_202 ();
 sg13g2_decap_8 FILLER_27_207 ();
 sg13g2_decap_8 FILLER_27_214 ();
 sg13g2_decap_4 FILLER_27_252 ();
 sg13g2_fill_2 FILLER_27_256 ();
 sg13g2_decap_4 FILLER_27_263 ();
 sg13g2_fill_2 FILLER_27_267 ();
 sg13g2_decap_8 FILLER_27_274 ();
 sg13g2_fill_2 FILLER_27_281 ();
 sg13g2_decap_4 FILLER_27_296 ();
 sg13g2_fill_2 FILLER_27_300 ();
 sg13g2_decap_4 FILLER_27_306 ();
 sg13g2_fill_1 FILLER_27_310 ();
 sg13g2_decap_8 FILLER_27_316 ();
 sg13g2_fill_1 FILLER_27_323 ();
 sg13g2_decap_8 FILLER_27_347 ();
 sg13g2_fill_2 FILLER_27_354 ();
 sg13g2_fill_1 FILLER_27_365 ();
 sg13g2_decap_4 FILLER_27_375 ();
 sg13g2_fill_1 FILLER_27_379 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_11 ();
 sg13g2_fill_2 FILLER_28_17 ();
 sg13g2_fill_2 FILLER_28_27 ();
 sg13g2_fill_1 FILLER_28_29 ();
 sg13g2_fill_2 FILLER_28_40 ();
 sg13g2_fill_2 FILLER_28_96 ();
 sg13g2_fill_1 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_103 ();
 sg13g2_fill_1 FILLER_28_110 ();
 sg13g2_fill_1 FILLER_28_116 ();
 sg13g2_fill_1 FILLER_28_129 ();
 sg13g2_fill_1 FILLER_28_134 ();
 sg13g2_fill_2 FILLER_28_161 ();
 sg13g2_fill_1 FILLER_28_167 ();
 sg13g2_decap_4 FILLER_28_172 ();
 sg13g2_fill_2 FILLER_28_176 ();
 sg13g2_decap_4 FILLER_28_204 ();
 sg13g2_fill_1 FILLER_28_208 ();
 sg13g2_decap_4 FILLER_28_213 ();
 sg13g2_fill_1 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_fill_1 FILLER_28_236 ();
 sg13g2_decap_8 FILLER_28_241 ();
 sg13g2_fill_2 FILLER_28_252 ();
 sg13g2_fill_1 FILLER_28_254 ();
 sg13g2_fill_2 FILLER_28_267 ();
 sg13g2_fill_2 FILLER_28_321 ();
 sg13g2_fill_1 FILLER_28_323 ();
 sg13g2_decap_4 FILLER_28_355 ();
 sg13g2_fill_1 FILLER_28_390 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_1 FILLER_29_29 ();
 sg13g2_decap_8 FILLER_29_66 ();
 sg13g2_fill_2 FILLER_29_77 ();
 sg13g2_fill_1 FILLER_29_79 ();
 sg13g2_fill_2 FILLER_29_85 ();
 sg13g2_fill_1 FILLER_29_87 ();
 sg13g2_fill_2 FILLER_29_154 ();
 sg13g2_fill_2 FILLER_29_182 ();
 sg13g2_fill_1 FILLER_29_184 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_fill_2 FILLER_29_196 ();
 sg13g2_decap_4 FILLER_29_233 ();
 sg13g2_fill_2 FILLER_29_277 ();
 sg13g2_fill_1 FILLER_29_279 ();
 sg13g2_decap_8 FILLER_29_284 ();
 sg13g2_decap_8 FILLER_29_291 ();
 sg13g2_decap_4 FILLER_29_298 ();
 sg13g2_fill_1 FILLER_29_302 ();
 sg13g2_decap_8 FILLER_29_329 ();
 sg13g2_decap_4 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_348 ();
 sg13g2_decap_8 FILLER_29_355 ();
 sg13g2_fill_1 FILLER_29_362 ();
 sg13g2_fill_2 FILLER_29_372 ();
 sg13g2_fill_1 FILLER_29_374 ();
 sg13g2_decap_4 FILLER_29_379 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_4 ();
 sg13g2_decap_8 FILLER_30_44 ();
 sg13g2_fill_1 FILLER_30_51 ();
 sg13g2_decap_8 FILLER_30_58 ();
 sg13g2_decap_8 FILLER_30_100 ();
 sg13g2_decap_4 FILLER_30_107 ();
 sg13g2_fill_1 FILLER_30_121 ();
 sg13g2_decap_8 FILLER_30_128 ();
 sg13g2_decap_8 FILLER_30_139 ();
 sg13g2_decap_8 FILLER_30_146 ();
 sg13g2_decap_8 FILLER_30_158 ();
 sg13g2_fill_2 FILLER_30_165 ();
 sg13g2_fill_2 FILLER_30_239 ();
 sg13g2_decap_4 FILLER_30_251 ();
 sg13g2_fill_2 FILLER_30_255 ();
 sg13g2_fill_1 FILLER_30_272 ();
 sg13g2_fill_2 FILLER_30_315 ();
 sg13g2_fill_1 FILLER_30_317 ();
 sg13g2_decap_4 FILLER_30_332 ();
 sg13g2_fill_1 FILLER_30_336 ();
 sg13g2_fill_2 FILLER_30_346 ();
 sg13g2_fill_1 FILLER_30_358 ();
 sg13g2_fill_2 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_14 ();
 sg13g2_decap_4 FILLER_31_24 ();
 sg13g2_fill_1 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_33 ();
 sg13g2_decap_4 FILLER_31_40 ();
 sg13g2_fill_1 FILLER_31_59 ();
 sg13g2_fill_1 FILLER_31_74 ();
 sg13g2_decap_8 FILLER_31_79 ();
 sg13g2_decap_8 FILLER_31_86 ();
 sg13g2_decap_8 FILLER_31_93 ();
 sg13g2_fill_2 FILLER_31_100 ();
 sg13g2_fill_2 FILLER_31_121 ();
 sg13g2_fill_1 FILLER_31_123 ();
 sg13g2_fill_2 FILLER_31_150 ();
 sg13g2_fill_1 FILLER_31_152 ();
 sg13g2_fill_2 FILLER_31_179 ();
 sg13g2_decap_8 FILLER_31_185 ();
 sg13g2_fill_2 FILLER_31_192 ();
 sg13g2_fill_1 FILLER_31_194 ();
 sg13g2_decap_4 FILLER_31_203 ();
 sg13g2_fill_1 FILLER_31_207 ();
 sg13g2_decap_8 FILLER_31_212 ();
 sg13g2_decap_4 FILLER_31_219 ();
 sg13g2_fill_2 FILLER_31_223 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_fill_2 FILLER_31_268 ();
 sg13g2_decap_8 FILLER_31_275 ();
 sg13g2_decap_4 FILLER_31_282 ();
 sg13g2_fill_1 FILLER_31_286 ();
 sg13g2_decap_8 FILLER_31_296 ();
 sg13g2_decap_8 FILLER_31_303 ();
 sg13g2_decap_4 FILLER_31_310 ();
 sg13g2_decap_4 FILLER_31_338 ();
 sg13g2_fill_1 FILLER_31_342 ();
 sg13g2_decap_8 FILLER_31_362 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_38 ();
 sg13g2_fill_1 FILLER_32_47 ();
 sg13g2_fill_1 FILLER_32_68 ();
 sg13g2_fill_1 FILLER_32_74 ();
 sg13g2_decap_4 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_92 ();
 sg13g2_decap_4 FILLER_32_99 ();
 sg13g2_fill_1 FILLER_32_103 ();
 sg13g2_fill_1 FILLER_32_134 ();
 sg13g2_decap_8 FILLER_32_139 ();
 sg13g2_decap_4 FILLER_32_146 ();
 sg13g2_fill_2 FILLER_32_150 ();
 sg13g2_decap_8 FILLER_32_156 ();
 sg13g2_fill_1 FILLER_32_163 ();
 sg13g2_fill_2 FILLER_32_168 ();
 sg13g2_fill_1 FILLER_32_170 ();
 sg13g2_fill_2 FILLER_32_197 ();
 sg13g2_decap_8 FILLER_32_241 ();
 sg13g2_decap_4 FILLER_32_248 ();
 sg13g2_fill_1 FILLER_32_252 ();
 sg13g2_fill_2 FILLER_32_258 ();
 sg13g2_fill_1 FILLER_32_260 ();
 sg13g2_decap_8 FILLER_32_304 ();
 sg13g2_fill_2 FILLER_32_337 ();
 sg13g2_fill_1 FILLER_32_339 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_4 ();
 sg13g2_fill_2 FILLER_33_31 ();
 sg13g2_fill_2 FILLER_33_47 ();
 sg13g2_decap_4 FILLER_33_73 ();
 sg13g2_decap_4 FILLER_33_103 ();
 sg13g2_fill_2 FILLER_33_107 ();
 sg13g2_fill_1 FILLER_33_112 ();
 sg13g2_fill_2 FILLER_33_122 ();
 sg13g2_fill_2 FILLER_33_129 ();
 sg13g2_decap_8 FILLER_33_157 ();
 sg13g2_decap_8 FILLER_33_164 ();
 sg13g2_fill_1 FILLER_33_171 ();
 sg13g2_decap_8 FILLER_33_177 ();
 sg13g2_decap_4 FILLER_33_184 ();
 sg13g2_decap_8 FILLER_33_191 ();
 sg13g2_decap_8 FILLER_33_198 ();
 sg13g2_decap_4 FILLER_33_205 ();
 sg13g2_fill_1 FILLER_33_213 ();
 sg13g2_decap_8 FILLER_33_240 ();
 sg13g2_fill_2 FILLER_33_247 ();
 sg13g2_decap_8 FILLER_33_275 ();
 sg13g2_fill_2 FILLER_33_282 ();
 sg13g2_fill_2 FILLER_33_288 ();
 sg13g2_decap_4 FILLER_33_300 ();
 sg13g2_decap_8 FILLER_33_309 ();
 sg13g2_fill_2 FILLER_33_324 ();
 sg13g2_decap_4 FILLER_33_333 ();
 sg13g2_fill_1 FILLER_33_337 ();
 sg13g2_decap_8 FILLER_33_342 ();
 sg13g2_fill_2 FILLER_33_349 ();
 sg13g2_fill_1 FILLER_33_351 ();
 sg13g2_decap_4 FILLER_33_361 ();
 sg13g2_fill_2 FILLER_33_380 ();
 sg13g2_fill_2 FILLER_33_387 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_14 ();
 sg13g2_decap_4 FILLER_34_19 ();
 sg13g2_fill_2 FILLER_34_23 ();
 sg13g2_decap_8 FILLER_34_44 ();
 sg13g2_fill_1 FILLER_34_51 ();
 sg13g2_fill_1 FILLER_34_62 ();
 sg13g2_decap_8 FILLER_34_75 ();
 sg13g2_decap_4 FILLER_34_82 ();
 sg13g2_fill_2 FILLER_34_86 ();
 sg13g2_decap_4 FILLER_34_93 ();
 sg13g2_fill_1 FILLER_34_97 ();
 sg13g2_fill_2 FILLER_34_102 ();
 sg13g2_fill_2 FILLER_34_123 ();
 sg13g2_fill_2 FILLER_34_130 ();
 sg13g2_decap_4 FILLER_34_137 ();
 sg13g2_fill_1 FILLER_34_141 ();
 sg13g2_decap_4 FILLER_34_146 ();
 sg13g2_fill_1 FILLER_34_150 ();
 sg13g2_fill_1 FILLER_34_156 ();
 sg13g2_fill_1 FILLER_34_183 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_fill_2 FILLER_34_223 ();
 sg13g2_decap_4 FILLER_34_229 ();
 sg13g2_decap_8 FILLER_34_237 ();
 sg13g2_fill_2 FILLER_34_244 ();
 sg13g2_decap_4 FILLER_34_255 ();
 sg13g2_decap_4 FILLER_34_263 ();
 sg13g2_decap_8 FILLER_34_272 ();
 sg13g2_decap_4 FILLER_34_279 ();
 sg13g2_fill_2 FILLER_34_283 ();
 sg13g2_fill_2 FILLER_34_311 ();
 sg13g2_fill_1 FILLER_34_339 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_decap_8 FILLER_35_29 ();
 sg13g2_decap_8 FILLER_35_36 ();
 sg13g2_fill_1 FILLER_35_43 ();
 sg13g2_fill_2 FILLER_35_49 ();
 sg13g2_decap_4 FILLER_35_57 ();
 sg13g2_decap_8 FILLER_35_132 ();
 sg13g2_fill_1 FILLER_35_167 ();
 sg13g2_decap_8 FILLER_35_172 ();
 sg13g2_decap_8 FILLER_35_179 ();
 sg13g2_decap_4 FILLER_35_186 ();
 sg13g2_fill_2 FILLER_35_190 ();
 sg13g2_fill_2 FILLER_35_199 ();
 sg13g2_fill_2 FILLER_35_205 ();
 sg13g2_fill_1 FILLER_35_207 ();
 sg13g2_fill_2 FILLER_35_243 ();
 sg13g2_fill_1 FILLER_35_271 ();
 sg13g2_decap_8 FILLER_35_302 ();
 sg13g2_fill_2 FILLER_35_309 ();
 sg13g2_decap_8 FILLER_35_316 ();
 sg13g2_fill_1 FILLER_35_323 ();
 sg13g2_fill_2 FILLER_35_332 ();
 sg13g2_fill_1 FILLER_35_334 ();
 sg13g2_fill_2 FILLER_35_345 ();
 sg13g2_fill_1 FILLER_35_355 ();
 sg13g2_fill_1 FILLER_35_392 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_4 FILLER_36_18 ();
 sg13g2_fill_2 FILLER_36_48 ();
 sg13g2_fill_2 FILLER_36_69 ();
 sg13g2_fill_1 FILLER_36_75 ();
 sg13g2_decap_8 FILLER_36_80 ();
 sg13g2_decap_4 FILLER_36_87 ();
 sg13g2_fill_1 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_97 ();
 sg13g2_decap_8 FILLER_36_104 ();
 sg13g2_fill_1 FILLER_36_111 ();
 sg13g2_fill_1 FILLER_36_120 ();
 sg13g2_fill_1 FILLER_36_152 ();
 sg13g2_fill_1 FILLER_36_157 ();
 sg13g2_decap_4 FILLER_36_184 ();
 sg13g2_fill_2 FILLER_36_188 ();
 sg13g2_decap_8 FILLER_36_216 ();
 sg13g2_decap_4 FILLER_36_223 ();
 sg13g2_decap_8 FILLER_36_231 ();
 sg13g2_decap_8 FILLER_36_238 ();
 sg13g2_decap_4 FILLER_36_245 ();
 sg13g2_fill_2 FILLER_36_249 ();
 sg13g2_fill_1 FILLER_36_255 ();
 sg13g2_decap_4 FILLER_36_260 ();
 sg13g2_fill_1 FILLER_36_264 ();
 sg13g2_decap_4 FILLER_36_277 ();
 sg13g2_fill_1 FILLER_36_281 ();
 sg13g2_fill_2 FILLER_36_304 ();
 sg13g2_fill_1 FILLER_36_306 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_4 FILLER_37_21 ();
 sg13g2_fill_2 FILLER_37_25 ();
 sg13g2_fill_2 FILLER_37_31 ();
 sg13g2_fill_2 FILLER_37_37 ();
 sg13g2_fill_1 FILLER_37_39 ();
 sg13g2_fill_1 FILLER_37_66 ();
 sg13g2_fill_2 FILLER_37_75 ();
 sg13g2_fill_1 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_120 ();
 sg13g2_decap_8 FILLER_37_127 ();
 sg13g2_fill_2 FILLER_37_134 ();
 sg13g2_fill_1 FILLER_37_136 ();
 sg13g2_decap_8 FILLER_37_141 ();
 sg13g2_decap_8 FILLER_37_148 ();
 sg13g2_decap_8 FILLER_37_155 ();
 sg13g2_decap_8 FILLER_37_162 ();
 sg13g2_decap_8 FILLER_37_173 ();
 sg13g2_decap_8 FILLER_37_180 ();
 sg13g2_decap_8 FILLER_37_187 ();
 sg13g2_decap_8 FILLER_37_194 ();
 sg13g2_decap_8 FILLER_37_201 ();
 sg13g2_decap_8 FILLER_37_208 ();
 sg13g2_decap_8 FILLER_37_215 ();
 sg13g2_decap_8 FILLER_37_222 ();
 sg13g2_decap_4 FILLER_37_229 ();
 sg13g2_fill_2 FILLER_37_233 ();
 sg13g2_fill_2 FILLER_37_239 ();
 sg13g2_decap_8 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_fill_2 FILLER_37_315 ();
 sg13g2_decap_4 FILLER_37_325 ();
 sg13g2_fill_2 FILLER_37_329 ();
 sg13g2_fill_2 FILLER_37_341 ();
 sg13g2_fill_1 FILLER_37_343 ();
 sg13g2_fill_1 FILLER_37_363 ();
 sg13g2_fill_2 FILLER_37_378 ();
 sg13g2_fill_1 FILLER_37_380 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_fill_2 FILLER_38_65 ();
 sg13g2_fill_2 FILLER_38_101 ();
 sg13g2_fill_1 FILLER_38_103 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_4 FILLER_38_180 ();
 sg13g2_decap_4 FILLER_38_188 ();
 sg13g2_decap_4 FILLER_38_196 ();
 sg13g2_decap_4 FILLER_38_204 ();
 sg13g2_decap_4 FILLER_38_212 ();
 sg13g2_decap_8 FILLER_38_220 ();
 sg13g2_decap_8 FILLER_38_227 ();
 sg13g2_decap_8 FILLER_38_234 ();
 sg13g2_decap_8 FILLER_38_241 ();
 sg13g2_decap_8 FILLER_38_248 ();
 sg13g2_decap_8 FILLER_38_255 ();
 sg13g2_decap_8 FILLER_38_262 ();
 sg13g2_decap_4 FILLER_38_269 ();
 sg13g2_fill_1 FILLER_38_273 ();
 sg13g2_fill_2 FILLER_38_278 ();
 sg13g2_fill_1 FILLER_38_280 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_fill_1 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_292 ();
 sg13g2_decap_8 FILLER_38_299 ();
 sg13g2_fill_2 FILLER_38_306 ();
 sg13g2_decap_4 FILLER_38_334 ();
 sg13g2_fill_1 FILLER_38_338 ();
 sg13g2_fill_2 FILLER_38_374 ();
 sg13g2_fill_1 FILLER_38_376 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
 assign uo_out[3] = net18;
 assign uo_out[4] = net19;
 assign uo_out[5] = net20;
 assign uo_out[6] = net21;
 assign uo_out[7] = net22;
endmodule

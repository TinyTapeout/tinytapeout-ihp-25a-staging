module tt_um_ddc_arghunter (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire \u_ddc_top_level.cic_left_inst.comb_out0[0] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out0[10] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out0[11] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out0[12] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out0[13] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out0[14] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out0[15] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out0[16] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out0[1] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out0[2] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out0[3] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out0[4] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out0[5] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out0[6] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out0[7] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out0[8] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out0[9] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out1[0] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out1[10] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out1[11] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out1[12] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out1[13] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out1[14] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out1[15] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out1[16] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out1[17] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out1[1] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out1[2] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out1[3] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out1[4] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out1[5] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out1[6] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out1[7] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out1[8] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out1[9] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out2[0] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out2[10] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out2[11] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out2[12] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out2[13] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out2[14] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out2[15] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out2[16] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out2[17] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out2[18] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out2[1] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out2[2] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out2[3] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out2[4] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out2[5] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out2[6] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out2[7] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out2[8] ;
 wire \u_ddc_top_level.cic_left_inst.comb_out2[9] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg0[0] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg0[10] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg0[11] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg0[12] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg0[13] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg0[14] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg0[15] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg0[1] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg0[2] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg0[3] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg0[4] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg0[5] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg0[6] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg0[7] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg0[8] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg0[9] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg1[0] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg1[10] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg1[11] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg1[12] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg1[13] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg1[14] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg1[15] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg1[16] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg1[1] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg1[2] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg1[3] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg1[4] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg1[5] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg1[6] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg1[7] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg1[8] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg1[9] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg2[0] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg2[10] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg2[11] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg2[12] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg2[13] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg2[14] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg2[15] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg2[16] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg2[17] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg2[1] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg2[2] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg2[3] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg2[4] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg2[5] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg2[6] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg2[7] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg2[8] ;
 wire \u_ddc_top_level.cic_left_inst.comb_reg2[9] ;
 wire \u_ddc_top_level.cic_left_inst.in_data[0] ;
 wire \u_ddc_top_level.cic_left_inst.in_data[10] ;
 wire \u_ddc_top_level.cic_left_inst.in_data[11] ;
 wire \u_ddc_top_level.cic_left_inst.in_data[12] ;
 wire \u_ddc_top_level.cic_left_inst.in_data[13] ;
 wire \u_ddc_top_level.cic_left_inst.in_data[14] ;
 wire \u_ddc_top_level.cic_left_inst.in_data[15] ;
 wire \u_ddc_top_level.cic_left_inst.in_data[1] ;
 wire \u_ddc_top_level.cic_left_inst.in_data[2] ;
 wire \u_ddc_top_level.cic_left_inst.in_data[3] ;
 wire \u_ddc_top_level.cic_left_inst.in_data[4] ;
 wire \u_ddc_top_level.cic_left_inst.in_data[5] ;
 wire \u_ddc_top_level.cic_left_inst.in_data[6] ;
 wire \u_ddc_top_level.cic_left_inst.in_data[7] ;
 wire \u_ddc_top_level.cic_left_inst.in_data[8] ;
 wire \u_ddc_top_level.cic_left_inst.in_data[9] ;
 wire \u_ddc_top_level.cic_left_inst.in_valid ;
 wire \u_ddc_top_level.cic_left_inst.int_reg0[0] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg0[10] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg0[11] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg0[12] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg0[13] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg0[14] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg0[15] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg0[16] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg0[17] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg0[18] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg0[19] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg0[1] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg0[2] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg0[3] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg0[4] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg0[5] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg0[6] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg0[7] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg0[8] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg0[9] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[0] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[10] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[11] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[12] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[13] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[14] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[15] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[16] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[17] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[18] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[19] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[1] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[20] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[21] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[22] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[23] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[2] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[3] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[4] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[5] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[6] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[7] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[8] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg1[9] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[0] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[10] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[11] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[12] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[13] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[14] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[15] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[16] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[17] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[18] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[19] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[1] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[20] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[21] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[22] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[23] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[24] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[25] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[26] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[27] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[2] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[3] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[4] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[5] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[6] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[7] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[8] ;
 wire \u_ddc_top_level.cic_left_inst.int_reg2[9] ;
 wire \u_ddc_top_level.cic_out_right[0] ;
 wire \u_ddc_top_level.cic_out_right[10] ;
 wire \u_ddc_top_level.cic_out_right[11] ;
 wire \u_ddc_top_level.cic_out_right[12] ;
 wire \u_ddc_top_level.cic_out_right[13] ;
 wire \u_ddc_top_level.cic_out_right[14] ;
 wire \u_ddc_top_level.cic_out_right[15] ;
 wire \u_ddc_top_level.cic_out_right[1] ;
 wire \u_ddc_top_level.cic_out_right[2] ;
 wire \u_ddc_top_level.cic_out_right[3] ;
 wire \u_ddc_top_level.cic_out_right[4] ;
 wire \u_ddc_top_level.cic_out_right[5] ;
 wire \u_ddc_top_level.cic_out_right[6] ;
 wire \u_ddc_top_level.cic_out_right[7] ;
 wire \u_ddc_top_level.cic_out_right[8] ;
 wire \u_ddc_top_level.cic_out_right[9] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out0[0] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out0[10] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out0[11] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out0[12] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out0[13] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out0[14] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out0[15] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out0[16] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out0[1] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out0[2] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out0[3] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out0[4] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out0[5] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out0[6] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out0[7] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out0[8] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out0[9] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out1[0] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out1[10] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out1[11] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out1[12] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out1[13] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out1[14] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out1[15] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out1[16] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out1[17] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out1[1] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out1[2] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out1[3] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out1[4] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out1[5] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out1[6] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out1[7] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out1[8] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out1[9] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out2[0] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out2[10] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out2[11] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out2[12] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out2[13] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out2[14] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out2[15] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out2[16] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out2[17] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out2[18] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out2[1] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out2[2] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out2[3] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out2[4] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out2[5] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out2[6] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out2[7] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out2[8] ;
 wire \u_ddc_top_level.cic_right_inst.comb_out2[9] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg0[0] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg0[10] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg0[11] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg0[12] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg0[13] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg0[14] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg0[15] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg0[1] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg0[2] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg0[3] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg0[4] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg0[5] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg0[6] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg0[7] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg0[8] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg0[9] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg1[0] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg1[10] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg1[11] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg1[12] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg1[13] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg1[14] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg1[15] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg1[16] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg1[1] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg1[2] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg1[3] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg1[4] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg1[5] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg1[6] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg1[7] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg1[8] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg1[9] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg2[0] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg2[10] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg2[11] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg2[12] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg2[13] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg2[14] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg2[15] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg2[16] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg2[17] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg2[1] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg2[2] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg2[3] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg2[4] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg2[5] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg2[6] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg2[7] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg2[8] ;
 wire \u_ddc_top_level.cic_right_inst.comb_reg2[9] ;
 wire \u_ddc_top_level.cic_right_inst.in_data[0] ;
 wire \u_ddc_top_level.cic_right_inst.in_data[10] ;
 wire \u_ddc_top_level.cic_right_inst.in_data[11] ;
 wire \u_ddc_top_level.cic_right_inst.in_data[12] ;
 wire \u_ddc_top_level.cic_right_inst.in_data[13] ;
 wire \u_ddc_top_level.cic_right_inst.in_data[14] ;
 wire \u_ddc_top_level.cic_right_inst.in_data[15] ;
 wire \u_ddc_top_level.cic_right_inst.in_data[1] ;
 wire \u_ddc_top_level.cic_right_inst.in_data[2] ;
 wire \u_ddc_top_level.cic_right_inst.in_data[3] ;
 wire \u_ddc_top_level.cic_right_inst.in_data[4] ;
 wire \u_ddc_top_level.cic_right_inst.in_data[5] ;
 wire \u_ddc_top_level.cic_right_inst.in_data[6] ;
 wire \u_ddc_top_level.cic_right_inst.in_data[7] ;
 wire \u_ddc_top_level.cic_right_inst.in_data[8] ;
 wire \u_ddc_top_level.cic_right_inst.in_data[9] ;
 wire \u_ddc_top_level.cic_right_inst.in_valid ;
 wire \u_ddc_top_level.cic_right_inst.int_reg0[0] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg0[10] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg0[11] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg0[12] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg0[13] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg0[14] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg0[15] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg0[16] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg0[17] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg0[18] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg0[19] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg0[1] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg0[2] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg0[3] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg0[4] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg0[5] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg0[6] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg0[7] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg0[8] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg0[9] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[0] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[10] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[11] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[12] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[13] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[14] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[15] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[16] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[17] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[18] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[19] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[1] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[20] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[21] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[22] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[23] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[2] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[3] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[4] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[5] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[6] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[7] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[8] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg1[9] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg2[0] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg2[10] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg2[11] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg2[1] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg2[2] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg2[3] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg2[4] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg2[5] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg2[6] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg2[7] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg2[8] ;
 wire \u_ddc_top_level.cic_right_inst.int_reg2[9] ;
 wire \u_ddc_top_level.dsm_left_inst.feedback[17] ;
 wire \u_ddc_top_level.dsm_left_inst.in_dither ;
 wire \u_ddc_top_level.dsm_left_inst.integrator1[0] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator1[10] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator1[11] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator1[12] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator1[13] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator1[14] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator1[15] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator1[16] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator1[17] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator1[18] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator1[1] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator1[2] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator1[3] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator1[4] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator1[5] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator1[6] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator1[7] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator1[8] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator1[9] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator2[0] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator2[10] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator2[11] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator2[12] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator2[13] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator2[14] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator2[15] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator2[16] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator2[17] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator2[1] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator2[2] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator2[3] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator2[4] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator2[5] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator2[6] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator2[7] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator2[8] ;
 wire \u_ddc_top_level.dsm_left_inst.integrator2[9] ;
 wire \u_ddc_top_level.dsm_left_inst.out_bitstream ;
 wire \u_ddc_top_level.dsm_right_inst.feedback[17] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator1[0] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator1[10] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator1[11] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator1[12] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator1[13] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator1[14] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator1[15] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator1[16] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator1[17] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator1[18] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator1[1] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator1[2] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator1[3] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator1[4] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator1[5] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator1[6] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator1[7] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator1[8] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator1[9] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator2[0] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator2[10] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator2[11] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator2[12] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator2[13] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator2[14] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator2[15] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator2[16] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator2[17] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator2[1] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator2[2] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator2[3] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator2[4] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator2[5] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator2[6] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator2[7] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator2[8] ;
 wire \u_ddc_top_level.dsm_right_inst.integrator2[9] ;
 wire \u_ddc_top_level.dsm_right_inst.out_bitstream ;
 wire \u_ddc_top_level.i2s_rx_inst.bit_count[0] ;
 wire \u_ddc_top_level.i2s_rx_inst.bit_count[1] ;
 wire \u_ddc_top_level.i2s_rx_inst.bit_count[2] ;
 wire \u_ddc_top_level.i2s_rx_inst.bit_count[3] ;
 wire \u_ddc_top_level.i2s_rx_inst.bit_count[4] ;
 wire \u_ddc_top_level.i2s_rx_inst.bit_count[5] ;
 wire \u_ddc_top_level.i2s_rx_inst.lrclk_prev ;
 wire \u_ddc_top_level.i2s_rx_inst.shift_reg[0] ;
 wire \u_ddc_top_level.i2s_rx_inst.shift_reg[10] ;
 wire \u_ddc_top_level.i2s_rx_inst.shift_reg[11] ;
 wire \u_ddc_top_level.i2s_rx_inst.shift_reg[12] ;
 wire \u_ddc_top_level.i2s_rx_inst.shift_reg[13] ;
 wire \u_ddc_top_level.i2s_rx_inst.shift_reg[14] ;
 wire \u_ddc_top_level.i2s_rx_inst.shift_reg[15] ;
 wire \u_ddc_top_level.i2s_rx_inst.shift_reg[1] ;
 wire \u_ddc_top_level.i2s_rx_inst.shift_reg[2] ;
 wire \u_ddc_top_level.i2s_rx_inst.shift_reg[3] ;
 wire \u_ddc_top_level.i2s_rx_inst.shift_reg[4] ;
 wire \u_ddc_top_level.i2s_rx_inst.shift_reg[5] ;
 wire \u_ddc_top_level.i2s_rx_inst.shift_reg[6] ;
 wire \u_ddc_top_level.i2s_rx_inst.shift_reg[7] ;
 wire \u_ddc_top_level.i2s_rx_inst.shift_reg[8] ;
 wire \u_ddc_top_level.i2s_rx_inst.shift_reg[9] ;
 wire \u_ddc_top_level.lsfr_inst.lfsr_reg[0] ;
 wire \u_ddc_top_level.lsfr_inst.lfsr_reg[10] ;
 wire \u_ddc_top_level.lsfr_inst.lfsr_reg[11] ;
 wire \u_ddc_top_level.lsfr_inst.lfsr_reg[12] ;
 wire \u_ddc_top_level.lsfr_inst.lfsr_reg[13] ;
 wire \u_ddc_top_level.lsfr_inst.lfsr_reg[14] ;
 wire \u_ddc_top_level.lsfr_inst.lfsr_reg[15] ;
 wire \u_ddc_top_level.lsfr_inst.lfsr_reg[1] ;
 wire \u_ddc_top_level.lsfr_inst.lfsr_reg[2] ;
 wire \u_ddc_top_level.lsfr_inst.lfsr_reg[3] ;
 wire \u_ddc_top_level.lsfr_inst.lfsr_reg[4] ;
 wire \u_ddc_top_level.lsfr_inst.lfsr_reg[5] ;
 wire \u_ddc_top_level.lsfr_inst.lfsr_reg[6] ;
 wire \u_ddc_top_level.lsfr_inst.lfsr_reg[7] ;
 wire \u_ddc_top_level.lsfr_inst.lfsr_reg[8] ;
 wire \u_ddc_top_level.lsfr_inst.lfsr_reg[9] ;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1;
 wire net2;
 wire net3;
 wire net4;

 sg13g2_a22oi_1 _3069_ (.Y(_0449_),
    .B1(_1291_),
    .B2(_1292_),
    .A2(_0743_),
    .A1(net813));
 sg13g2_nand2_1 _3070_ (.Y(_1293_),
    .A(net816),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[17] ));
 sg13g2_nor2b_1 _3071_ (.A(\u_ddc_top_level.cic_right_inst.comb_reg1[16] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_out0[16] ),
    .Y(_1294_));
 sg13g2_xor2_1 _3072_ (.B(\u_ddc_top_level.cic_right_inst.comb_reg1[16] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_out0[16] ),
    .X(_1295_));
 sg13g2_nor2b_1 _3073_ (.A(\u_ddc_top_level.cic_right_inst.comb_reg1[7] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_out0[7] ),
    .Y(_1296_));
 sg13g2_nor2b_1 _3074_ (.A(\u_ddc_top_level.cic_right_inst.comb_reg1[5] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_out0[5] ),
    .Y(_1297_));
 sg13g2_nand2b_1 _3075_ (.Y(_1298_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg1[5] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_out0[5] ));
 sg13g2_nand2b_1 _3076_ (.Y(_1299_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg1[4] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_out0[4] ));
 sg13g2_nand2b_1 _3077_ (.Y(_1300_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg1[3] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_out0[3] ));
 sg13g2_xor2_1 _3078_ (.B(\u_ddc_top_level.cic_right_inst.comb_reg1[3] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_out0[3] ),
    .X(_1301_));
 sg13g2_nor2b_1 _3079_ (.A(\u_ddc_top_level.cic_right_inst.comb_out0[2] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg1[2] ),
    .Y(_1302_));
 sg13g2_nand2b_1 _3080_ (.Y(_1303_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg1[1] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_out0[1] ));
 sg13g2_nor2b_1 _3081_ (.A(\u_ddc_top_level.cic_right_inst.comb_reg1[0] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_out0[0] ),
    .Y(_1304_));
 sg13g2_nor2b_1 _3082_ (.A(\u_ddc_top_level.cic_right_inst.comb_reg1[1] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_out0[1] ),
    .Y(_1305_));
 sg13g2_xnor2_1 _3083_ (.Y(_1306_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out0[1] ),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg1[1] ));
 sg13g2_o21ai_1 _3084_ (.B1(_1303_),
    .Y(_1307_),
    .A1(_1304_),
    .A2(_1305_));
 sg13g2_xnor2_1 _3085_ (.Y(_1308_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out0[2] ),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg1[2] ));
 sg13g2_a21oi_1 _3086_ (.A1(_1307_),
    .A2(_1308_),
    .Y(_1309_),
    .B1(_1302_));
 sg13g2_o21ai_1 _3087_ (.B1(_1300_),
    .Y(_1310_),
    .A1(_1301_),
    .A2(_1309_));
 sg13g2_xnor2_1 _3088_ (.Y(_1311_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out0[4] ),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg1[4] ));
 sg13g2_nand2_1 _3089_ (.Y(_1312_),
    .A(_1310_),
    .B(_1311_));
 sg13g2_nand2_1 _3090_ (.Y(_1313_),
    .A(_1299_),
    .B(_1312_));
 sg13g2_o21ai_1 _3091_ (.B1(_1298_),
    .Y(_1314_),
    .A1(_1297_),
    .A2(_1299_));
 sg13g2_nor2b_1 _3092_ (.A(_1297_),
    .B_N(_1298_),
    .Y(_1315_));
 sg13g2_and2_1 _3093_ (.A(_1311_),
    .B(_1315_),
    .X(_1316_));
 sg13g2_a21o_1 _3094_ (.A2(_1316_),
    .A1(_1310_),
    .B1(_1314_),
    .X(_1317_));
 sg13g2_a21oi_1 _3095_ (.A1(_1310_),
    .A2(_1316_),
    .Y(_1318_),
    .B1(_1314_));
 sg13g2_nand2b_1 _3096_ (.Y(_1319_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg1[6] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_out0[6] ));
 sg13g2_xor2_1 _3097_ (.B(\u_ddc_top_level.cic_right_inst.comb_reg1[6] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_out0[6] ),
    .X(_1320_));
 sg13g2_nand2b_1 _3098_ (.Y(_1321_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg1[7] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_out0[7] ));
 sg13g2_o21ai_1 _3099_ (.B1(_1321_),
    .Y(_1322_),
    .A1(_1296_),
    .A2(_1319_));
 sg13g2_nor2b_1 _3100_ (.A(_1296_),
    .B_N(_1321_),
    .Y(_1323_));
 sg13g2_nor2b_1 _3101_ (.A(_1320_),
    .B_N(_1323_),
    .Y(_1324_));
 sg13g2_a21oi_2 _3102_ (.B1(_1322_),
    .Y(_1325_),
    .A2(_1324_),
    .A1(_1317_));
 sg13g2_nor2b_1 _3103_ (.A(\u_ddc_top_level.cic_right_inst.comb_reg1[9] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_out0[9] ),
    .Y(_1326_));
 sg13g2_nand2b_1 _3104_ (.Y(_1327_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg1[9] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_out0[9] ));
 sg13g2_nand2b_1 _3105_ (.Y(_1328_),
    .B(_1327_),
    .A_N(_1326_));
 sg13g2_nand2b_1 _3106_ (.Y(_1329_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg1[8] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_out0[8] ));
 sg13g2_xor2_1 _3107_ (.B(\u_ddc_top_level.cic_right_inst.comb_reg1[8] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_out0[8] ),
    .X(_1330_));
 sg13g2_nor3_1 _3108_ (.A(_1325_),
    .B(_1328_),
    .C(_1330_),
    .Y(_1331_));
 sg13g2_o21ai_1 _3109_ (.B1(_1327_),
    .Y(_1332_),
    .A1(_1326_),
    .A2(_1329_));
 sg13g2_nand2_1 _3110_ (.Y(_1333_),
    .A(_0717_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg1[10] ));
 sg13g2_nor2b_1 _3111_ (.A(\u_ddc_top_level.cic_right_inst.comb_reg1[11] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_out0[11] ),
    .Y(_1334_));
 sg13g2_nand2b_1 _3112_ (.Y(_1335_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg1[11] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_out0[11] ));
 sg13g2_o21ai_1 _3113_ (.B1(_1335_),
    .Y(_1336_),
    .A1(_1333_),
    .A2(_1334_));
 sg13g2_or2_1 _3114_ (.X(_1337_),
    .B(_1336_),
    .A(_1332_));
 sg13g2_nor2_1 _3115_ (.A(_0717_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg1[10] ),
    .Y(_1338_));
 sg13g2_o21ai_1 _3116_ (.B1(_1335_),
    .Y(_1339_),
    .A1(_1334_),
    .A2(_1338_));
 sg13g2_o21ai_1 _3117_ (.B1(_1339_),
    .Y(_1340_),
    .A1(_1331_),
    .A2(_1337_));
 sg13g2_xor2_1 _3118_ (.B(\u_ddc_top_level.cic_right_inst.comb_reg1[13] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_out0[13] ),
    .X(_1341_));
 sg13g2_nand2b_1 _3119_ (.Y(_1342_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg1[12] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_out0[12] ));
 sg13g2_xor2_1 _3120_ (.B(\u_ddc_top_level.cic_right_inst.comb_reg1[12] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_out0[12] ),
    .X(_1343_));
 sg13g2_or2_1 _3121_ (.X(_1344_),
    .B(_1343_),
    .A(_1341_));
 sg13g2_a21oi_1 _3122_ (.A1(\u_ddc_top_level.cic_right_inst.comb_out0[13] ),
    .A2(_0737_),
    .Y(_1345_),
    .B1(_1342_));
 sg13g2_a21oi_1 _3123_ (.A1(_0716_),
    .A2(\u_ddc_top_level.cic_right_inst.comb_reg1[13] ),
    .Y(_1346_),
    .B1(_1345_));
 sg13g2_o21ai_1 _3124_ (.B1(_1346_),
    .Y(_1347_),
    .A1(_1340_),
    .A2(_1344_));
 sg13g2_nor2b_1 _3125_ (.A(\u_ddc_top_level.cic_right_inst.comb_out0[15] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg1[15] ),
    .Y(_1348_));
 sg13g2_nand2b_1 _3126_ (.Y(_1349_),
    .B(\u_ddc_top_level.cic_right_inst.comb_out0[15] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_reg1[15] ));
 sg13g2_nand2b_1 _3127_ (.Y(_1350_),
    .B(_1349_),
    .A_N(_1348_));
 sg13g2_nor2b_1 _3128_ (.A(\u_ddc_top_level.cic_right_inst.comb_out0[14] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg1[14] ),
    .Y(_1351_));
 sg13g2_nand2b_1 _3129_ (.Y(_1352_),
    .B(\u_ddc_top_level.cic_right_inst.comb_out0[14] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_reg1[14] ));
 sg13g2_nand2b_1 _3130_ (.Y(_1353_),
    .B(_1352_),
    .A_N(_1351_));
 sg13g2_nor2_1 _3131_ (.A(_1350_),
    .B(_1353_),
    .Y(_1354_));
 sg13g2_a221oi_1 _3132_ (.B2(_1347_),
    .C1(_1348_),
    .B1(_1354_),
    .A1(_1349_),
    .Y(_1355_),
    .A2(_1351_));
 sg13g2_o21ai_1 _3133_ (.B1(net873),
    .Y(_1356_),
    .A1(_1295_),
    .A2(_1355_));
 sg13g2_o21ai_1 _3134_ (.B1(_1293_),
    .Y(_0448_),
    .A1(_1294_),
    .A2(_1356_));
 sg13g2_nand2_1 _3135_ (.Y(_1357_),
    .A(net816),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[16] ));
 sg13g2_and2_1 _3136_ (.A(_1295_),
    .B(_1355_),
    .X(_1358_));
 sg13g2_o21ai_1 _3137_ (.B1(_1357_),
    .Y(_0447_),
    .A1(_1356_),
    .A2(_1358_));
 sg13g2_a21oi_1 _3138_ (.A1(_1347_),
    .A2(_1352_),
    .Y(_1359_),
    .B1(_1351_));
 sg13g2_nand2_1 _3139_ (.Y(_1360_),
    .A(net815),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[15] ));
 sg13g2_xnor2_1 _3140_ (.Y(_1361_),
    .A(_1350_),
    .B(_1359_));
 sg13g2_o21ai_1 _3141_ (.B1(_1360_),
    .Y(_0446_),
    .A1(net815),
    .A2(_1361_));
 sg13g2_nor2_1 _3142_ (.A(net873),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[14] ),
    .Y(_1362_));
 sg13g2_xor2_1 _3143_ (.B(_1353_),
    .A(_1347_),
    .X(_1363_));
 sg13g2_a21oi_1 _3144_ (.A1(net873),
    .A2(_1363_),
    .Y(_0445_),
    .B1(_1362_));
 sg13g2_o21ai_1 _3145_ (.B1(_1342_),
    .Y(_1364_),
    .A1(_1340_),
    .A2(_1343_));
 sg13g2_o21ai_1 _3146_ (.B1(net874),
    .Y(_1365_),
    .A1(_1341_),
    .A2(_1364_));
 sg13g2_a21oi_1 _3147_ (.A1(_1341_),
    .A2(_1364_),
    .Y(_1366_),
    .B1(_1365_));
 sg13g2_a21oi_1 _3148_ (.A1(net816),
    .A2(_0733_),
    .Y(_0444_),
    .B1(_1366_));
 sg13g2_o21ai_1 _3149_ (.B1(net874),
    .Y(_1367_),
    .A1(_1340_),
    .A2(_1343_));
 sg13g2_a21oi_1 _3150_ (.A1(_1340_),
    .A2(_1343_),
    .Y(_1368_),
    .B1(_1367_));
 sg13g2_a21o_1 _3151_ (.A2(\u_ddc_top_level.cic_right_inst.comb_out1[12] ),
    .A1(net816),
    .B1(_1368_),
    .X(_0443_));
 sg13g2_nand2b_1 _3152_ (.Y(_1369_),
    .B(_1335_),
    .A_N(_1334_));
 sg13g2_xor2_1 _3153_ (.B(\u_ddc_top_level.cic_right_inst.comb_reg1[10] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_out0[10] ),
    .X(_1370_));
 sg13g2_nor2_1 _3154_ (.A(_1331_),
    .B(_1332_),
    .Y(_1371_));
 sg13g2_o21ai_1 _3155_ (.B1(_1333_),
    .Y(_1372_),
    .A1(_1338_),
    .A2(_1371_));
 sg13g2_xnor2_1 _3156_ (.Y(_1373_),
    .A(_1369_),
    .B(_1372_));
 sg13g2_mux2_1 _3157_ (.A0(\u_ddc_top_level.cic_right_inst.comb_out1[11] ),
    .A1(_1373_),
    .S(net872),
    .X(_0442_));
 sg13g2_o21ai_1 _3158_ (.B1(net874),
    .Y(_1374_),
    .A1(_1370_),
    .A2(_1371_));
 sg13g2_a21oi_1 _3159_ (.A1(_1370_),
    .A2(_1371_),
    .Y(_1375_),
    .B1(_1374_));
 sg13g2_a21o_1 _3160_ (.A2(\u_ddc_top_level.cic_right_inst.comb_out1[10] ),
    .A1(net816),
    .B1(_1375_),
    .X(_0441_));
 sg13g2_o21ai_1 _3161_ (.B1(_1329_),
    .Y(_1376_),
    .A1(_1325_),
    .A2(_1330_));
 sg13g2_o21ai_1 _3162_ (.B1(net866),
    .Y(_1377_),
    .A1(_1328_),
    .A2(_1376_));
 sg13g2_a21oi_1 _3163_ (.A1(_1328_),
    .A2(_1376_),
    .Y(_1378_),
    .B1(_1377_));
 sg13g2_a21oi_1 _3164_ (.A1(net814),
    .A2(_0734_),
    .Y(_0440_),
    .B1(_1378_));
 sg13g2_o21ai_1 _3165_ (.B1(net866),
    .Y(_1379_),
    .A1(_1325_),
    .A2(_1330_));
 sg13g2_a21oi_1 _3166_ (.A1(_1325_),
    .A2(_1330_),
    .Y(_1380_),
    .B1(_1379_));
 sg13g2_a21o_1 _3167_ (.A2(\u_ddc_top_level.cic_right_inst.comb_out1[8] ),
    .A1(net814),
    .B1(_1380_),
    .X(_0439_));
 sg13g2_o21ai_1 _3168_ (.B1(_1319_),
    .Y(_1381_),
    .A1(_1318_),
    .A2(_1320_));
 sg13g2_nand2_1 _3169_ (.Y(_1382_),
    .A(net814),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[7] ));
 sg13g2_and2_1 _3170_ (.A(_1323_),
    .B(_1381_),
    .X(_1383_));
 sg13g2_o21ai_1 _3171_ (.B1(net867),
    .Y(_1384_),
    .A1(_1323_),
    .A2(_1381_));
 sg13g2_o21ai_1 _3172_ (.B1(_1382_),
    .Y(_0438_),
    .A1(_1383_),
    .A2(_1384_));
 sg13g2_o21ai_1 _3173_ (.B1(net867),
    .Y(_1385_),
    .A1(_1318_),
    .A2(_1320_));
 sg13g2_a21oi_1 _3174_ (.A1(_1318_),
    .A2(_1320_),
    .Y(_1386_),
    .B1(_1385_));
 sg13g2_a21o_1 _3175_ (.A2(\u_ddc_top_level.cic_right_inst.comb_out1[6] ),
    .A1(net814),
    .B1(_1386_),
    .X(_0437_));
 sg13g2_o21ai_1 _3176_ (.B1(net865),
    .Y(_1387_),
    .A1(_1313_),
    .A2(_1315_));
 sg13g2_a21oi_1 _3177_ (.A1(_1313_),
    .A2(_1315_),
    .Y(_1388_),
    .B1(_1387_));
 sg13g2_a21o_1 _3178_ (.A2(\u_ddc_top_level.cic_right_inst.comb_out1[5] ),
    .A1(net814),
    .B1(_1388_),
    .X(_0436_));
 sg13g2_nor2_1 _3179_ (.A(net864),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[4] ),
    .Y(_1389_));
 sg13g2_xnor2_1 _3180_ (.Y(_1390_),
    .A(_1310_),
    .B(_1311_));
 sg13g2_a21oi_1 _3181_ (.A1(net864),
    .A2(_1390_),
    .Y(_0435_),
    .B1(_1389_));
 sg13g2_nor2_1 _3182_ (.A(net855),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[3] ),
    .Y(_1391_));
 sg13g2_xnor2_1 _3183_ (.Y(_1392_),
    .A(_1301_),
    .B(_1309_));
 sg13g2_a21oi_1 _3184_ (.A1(net855),
    .A2(_1392_),
    .Y(_0434_),
    .B1(_1391_));
 sg13g2_nor2_1 _3185_ (.A(net854),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[2] ),
    .Y(_1393_));
 sg13g2_xnor2_1 _3186_ (.Y(_1394_),
    .A(_1307_),
    .B(_1308_));
 sg13g2_a21oi_1 _3187_ (.A1(net855),
    .A2(_1394_),
    .Y(_0433_),
    .B1(_1393_));
 sg13g2_xnor2_1 _3188_ (.Y(_1395_),
    .A(_1304_),
    .B(_1306_));
 sg13g2_mux2_1 _3189_ (.A0(\u_ddc_top_level.cic_right_inst.comb_out1[1] ),
    .A1(_1395_),
    .S(net854),
    .X(_0432_));
 sg13g2_nor2b_1 _3190_ (.A(\u_ddc_top_level.cic_right_inst.comb_out0[0] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg1[0] ),
    .Y(_1396_));
 sg13g2_nor3_1 _3191_ (.A(net813),
    .B(_1304_),
    .C(_1396_),
    .Y(_1397_));
 sg13g2_a21oi_1 _3192_ (.A1(net813),
    .A2(_0736_),
    .Y(_0431_),
    .B1(_1397_));
 sg13g2_nor2b_1 _3193_ (.A(net1),
    .B_N(\u_ddc_top_level.i2s_rx_inst.lrclk_prev ),
    .Y(_1398_));
 sg13g2_nor2b_1 _3194_ (.A(\u_ddc_top_level.i2s_rx_inst.lrclk_prev ),
    .B_N(net1),
    .Y(_1399_));
 sg13g2_or2_2 _3195_ (.X(_1400_),
    .B(net819),
    .A(net822));
 sg13g2_nor2_1 _3196_ (.A(\u_ddc_top_level.i2s_rx_inst.bit_count[0] ),
    .B(_1400_),
    .Y(_0000_));
 sg13g2_and2_1 _3197_ (.A(\u_ddc_top_level.i2s_rx_inst.bit_count[0] ),
    .B(\u_ddc_top_level.i2s_rx_inst.bit_count[1] ),
    .X(_1401_));
 sg13g2_nor2_1 _3198_ (.A(\u_ddc_top_level.i2s_rx_inst.bit_count[0] ),
    .B(\u_ddc_top_level.i2s_rx_inst.bit_count[1] ),
    .Y(_1402_));
 sg13g2_nor3_1 _3199_ (.A(_1400_),
    .B(_1401_),
    .C(_1402_),
    .Y(_0001_));
 sg13g2_a21oi_1 _3200_ (.A1(\u_ddc_top_level.i2s_rx_inst.bit_count[2] ),
    .A2(_1401_),
    .Y(_1403_),
    .B1(_1400_));
 sg13g2_o21ai_1 _3201_ (.B1(_1403_),
    .Y(_1404_),
    .A1(\u_ddc_top_level.i2s_rx_inst.bit_count[2] ),
    .A2(_1401_));
 sg13g2_inv_1 _3202_ (.Y(_0002_),
    .A(_1404_));
 sg13g2_a21oi_1 _3203_ (.A1(\u_ddc_top_level.i2s_rx_inst.bit_count[2] ),
    .A2(_1401_),
    .Y(_1405_),
    .B1(\u_ddc_top_level.i2s_rx_inst.bit_count[3] ));
 sg13g2_and3_1 _3204_ (.X(_1406_),
    .A(\u_ddc_top_level.i2s_rx_inst.bit_count[2] ),
    .B(\u_ddc_top_level.i2s_rx_inst.bit_count[3] ),
    .C(_1401_));
 sg13g2_nor3_1 _3205_ (.A(_1400_),
    .B(_1405_),
    .C(_1406_),
    .Y(_0003_));
 sg13g2_nor2_1 _3206_ (.A(\u_ddc_top_level.i2s_rx_inst.bit_count[4] ),
    .B(_1406_),
    .Y(_1407_));
 sg13g2_and2_1 _3207_ (.A(\u_ddc_top_level.i2s_rx_inst.bit_count[4] ),
    .B(_1406_),
    .X(_1408_));
 sg13g2_nor3_1 _3208_ (.A(_1400_),
    .B(_1407_),
    .C(_1408_),
    .Y(_0004_));
 sg13g2_a21oi_1 _3209_ (.A1(\u_ddc_top_level.i2s_rx_inst.bit_count[5] ),
    .A2(_1408_),
    .Y(_1409_),
    .B1(_1400_));
 sg13g2_o21ai_1 _3210_ (.B1(_1409_),
    .Y(_1410_),
    .A1(\u_ddc_top_level.i2s_rx_inst.bit_count[5] ),
    .A2(_1408_));
 sg13g2_inv_1 _3211_ (.Y(_0005_),
    .A(_1410_));
 sg13g2_nand2_1 _3212_ (.Y(_1411_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg2[0] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[0] ));
 sg13g2_xor2_1 _3213_ (.B(\u_ddc_top_level.cic_right_inst.int_reg1[0] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg2[0] ),
    .X(_0083_));
 sg13g2_nand2_1 _3214_ (.Y(_1412_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg2[1] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[1] ));
 sg13g2_nor2_1 _3215_ (.A(\u_ddc_top_level.cic_right_inst.int_reg2[1] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[1] ),
    .Y(_1413_));
 sg13g2_xor2_1 _3216_ (.B(\u_ddc_top_level.cic_right_inst.int_reg1[1] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg2[1] ),
    .X(_1414_));
 sg13g2_xnor2_1 _3217_ (.Y(_0094_),
    .A(_1411_),
    .B(_1414_));
 sg13g2_o21ai_1 _3218_ (.B1(_1412_),
    .Y(_1415_),
    .A1(_1411_),
    .A2(_1413_));
 sg13g2_and2_1 _3219_ (.A(\u_ddc_top_level.cic_right_inst.int_reg2[2] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[2] ),
    .X(_1416_));
 sg13g2_or2_1 _3220_ (.X(_1417_),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[2] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg2[2] ));
 sg13g2_nand2b_1 _3221_ (.Y(_1418_),
    .B(_1417_),
    .A_N(_1416_));
 sg13g2_xnor2_1 _3222_ (.Y(_0103_),
    .A(_1415_),
    .B(_1418_));
 sg13g2_a21o_1 _3223_ (.A2(_1417_),
    .A1(_1415_),
    .B1(_1416_),
    .X(_1419_));
 sg13g2_and2_1 _3224_ (.A(\u_ddc_top_level.cic_right_inst.int_reg2[3] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[3] ),
    .X(_1420_));
 sg13g2_or2_1 _3225_ (.X(_1421_),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[3] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg2[3] ));
 sg13g2_nand2b_1 _3226_ (.Y(_1422_),
    .B(_1421_),
    .A_N(_1420_));
 sg13g2_xnor2_1 _3227_ (.Y(_0104_),
    .A(_1419_),
    .B(_1422_));
 sg13g2_a21o_1 _3228_ (.A2(_1421_),
    .A1(_1419_),
    .B1(_1420_),
    .X(_1423_));
 sg13g2_xnor2_1 _3229_ (.Y(_1424_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg2[4] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[4] ));
 sg13g2_nor2b_1 _3230_ (.A(_1424_),
    .B_N(_1423_),
    .Y(_1425_));
 sg13g2_xnor2_1 _3231_ (.Y(_0105_),
    .A(_1423_),
    .B(_1424_));
 sg13g2_nor2_1 _3232_ (.A(\u_ddc_top_level.cic_right_inst.int_reg2[5] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[5] ),
    .Y(_1426_));
 sg13g2_xnor2_1 _3233_ (.Y(_1427_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg2[5] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[5] ));
 sg13g2_a21oi_1 _3234_ (.A1(\u_ddc_top_level.cic_right_inst.int_reg2[4] ),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg1[4] ),
    .Y(_1428_),
    .B1(_1425_));
 sg13g2_xor2_1 _3235_ (.B(_1428_),
    .A(_1427_),
    .X(_0106_));
 sg13g2_nor2_1 _3236_ (.A(\u_ddc_top_level.cic_right_inst.int_reg2[6] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[6] ),
    .Y(_1429_));
 sg13g2_xor2_1 _3237_ (.B(\u_ddc_top_level.cic_right_inst.int_reg1[6] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg2[6] ),
    .X(_1430_));
 sg13g2_a22oi_1 _3238_ (.Y(_1431_),
    .B1(\u_ddc_top_level.cic_right_inst.int_reg2[5] ),
    .B2(\u_ddc_top_level.cic_right_inst.int_reg1[5] ),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg1[4] ),
    .A1(\u_ddc_top_level.cic_right_inst.int_reg2[4] ));
 sg13g2_nor2_1 _3239_ (.A(_1424_),
    .B(_1427_),
    .Y(_1432_));
 sg13g2_nor2_1 _3240_ (.A(_1426_),
    .B(_1431_),
    .Y(_1433_));
 sg13g2_a21oi_1 _3241_ (.A1(_1423_),
    .A2(_1432_),
    .Y(_1434_),
    .B1(_1433_));
 sg13g2_xnor2_1 _3242_ (.Y(_0107_),
    .A(_1430_),
    .B(_1434_));
 sg13g2_nand2_1 _3243_ (.Y(_1435_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg2[7] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[7] ));
 sg13g2_nor2_1 _3244_ (.A(\u_ddc_top_level.cic_right_inst.int_reg2[7] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[7] ),
    .Y(_1436_));
 sg13g2_xnor2_1 _3245_ (.Y(_1437_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg2[7] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[7] ));
 sg13g2_a221oi_1 _3246_ (.B2(_1432_),
    .C1(_1433_),
    .B1(_1423_),
    .A1(\u_ddc_top_level.cic_right_inst.int_reg2[6] ),
    .Y(_1438_),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg1[6] ));
 sg13g2_nor2_1 _3247_ (.A(_1429_),
    .B(_1438_),
    .Y(_1439_));
 sg13g2_xnor2_1 _3248_ (.Y(_0108_),
    .A(_1437_),
    .B(_1439_));
 sg13g2_xnor2_1 _3249_ (.Y(_1440_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg2[8] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[8] ));
 sg13g2_or2_1 _3250_ (.X(_1441_),
    .B(_1436_),
    .A(_1429_));
 sg13g2_o21ai_1 _3251_ (.B1(_1435_),
    .Y(_1442_),
    .A1(_1438_),
    .A2(_1441_));
 sg13g2_nor2b_1 _3252_ (.A(_1440_),
    .B_N(_1442_),
    .Y(_1443_));
 sg13g2_xnor2_1 _3253_ (.Y(_0109_),
    .A(_1440_),
    .B(_1442_));
 sg13g2_nor2_1 _3254_ (.A(\u_ddc_top_level.cic_right_inst.int_reg2[9] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[9] ),
    .Y(_1444_));
 sg13g2_xnor2_1 _3255_ (.Y(_1445_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg2[9] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[9] ));
 sg13g2_a21oi_1 _3256_ (.A1(\u_ddc_top_level.cic_right_inst.int_reg2[8] ),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg1[8] ),
    .Y(_1446_),
    .B1(_1443_));
 sg13g2_xor2_1 _3257_ (.B(_1446_),
    .A(_1445_),
    .X(_0110_));
 sg13g2_nand2_1 _3258_ (.Y(_1447_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg2[10] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[10] ));
 sg13g2_xnor2_1 _3259_ (.Y(_1448_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg2[10] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[10] ));
 sg13g2_a22oi_1 _3260_ (.Y(_1449_),
    .B1(\u_ddc_top_level.cic_right_inst.int_reg2[9] ),
    .B2(\u_ddc_top_level.cic_right_inst.int_reg1[9] ),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg1[8] ),
    .A1(\u_ddc_top_level.cic_right_inst.int_reg2[8] ));
 sg13g2_nor2_1 _3261_ (.A(_1444_),
    .B(_1449_),
    .Y(_1450_));
 sg13g2_nor2_1 _3262_ (.A(_1440_),
    .B(_1445_),
    .Y(_1451_));
 sg13g2_a21oi_1 _3263_ (.A1(_1442_),
    .A2(_1451_),
    .Y(_1452_),
    .B1(_1450_));
 sg13g2_xor2_1 _3264_ (.B(_1452_),
    .A(_1448_),
    .X(_0084_));
 sg13g2_nor2_1 _3265_ (.A(\u_ddc_top_level.cic_right_inst.int_reg2[11] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[11] ),
    .Y(_1453_));
 sg13g2_nand2_1 _3266_ (.Y(_1454_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg2[11] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[11] ));
 sg13g2_nor2b_1 _3267_ (.A(_1453_),
    .B_N(_1454_),
    .Y(_1455_));
 sg13g2_o21ai_1 _3268_ (.B1(_1447_),
    .Y(_1456_),
    .A1(_1448_),
    .A2(_1452_));
 sg13g2_xor2_1 _3269_ (.B(_1456_),
    .A(_1455_),
    .X(_0085_));
 sg13g2_nor2b_1 _3270_ (.A(_1448_),
    .B_N(_1455_),
    .Y(_1457_));
 sg13g2_and2_1 _3271_ (.A(_1451_),
    .B(_1457_),
    .X(_1458_));
 sg13g2_o21ai_1 _3272_ (.B1(_1454_),
    .Y(_1459_),
    .A1(_1447_),
    .A2(_1453_));
 sg13g2_a21o_1 _3273_ (.A2(_1457_),
    .A1(_1450_),
    .B1(_1459_),
    .X(_1460_));
 sg13g2_a21o_2 _3274_ (.A2(_1458_),
    .A1(_1442_),
    .B1(_1460_),
    .X(_1461_));
 sg13g2_nand2_1 _3275_ (.Y(_1462_),
    .A(\u_ddc_top_level.cic_out_right[0] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[12] ));
 sg13g2_xor2_1 _3276_ (.B(\u_ddc_top_level.cic_right_inst.int_reg1[12] ),
    .A(\u_ddc_top_level.cic_out_right[0] ),
    .X(_1463_));
 sg13g2_nand2_1 _3277_ (.Y(_1464_),
    .A(_1461_),
    .B(_1463_));
 sg13g2_xor2_1 _3278_ (.B(_1463_),
    .A(_1461_),
    .X(_0086_));
 sg13g2_nor2_1 _3279_ (.A(\u_ddc_top_level.cic_out_right[1] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[13] ),
    .Y(_1465_));
 sg13g2_xor2_1 _3280_ (.B(\u_ddc_top_level.cic_right_inst.int_reg1[13] ),
    .A(\u_ddc_top_level.cic_out_right[1] ),
    .X(_1466_));
 sg13g2_and2_1 _3281_ (.A(_1462_),
    .B(_1464_),
    .X(_1467_));
 sg13g2_xnor2_1 _3282_ (.Y(_0087_),
    .A(_1466_),
    .B(_1467_));
 sg13g2_and2_1 _3283_ (.A(\u_ddc_top_level.cic_out_right[2] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[14] ),
    .X(_1468_));
 sg13g2_xor2_1 _3284_ (.B(\u_ddc_top_level.cic_right_inst.int_reg1[14] ),
    .A(\u_ddc_top_level.cic_out_right[2] ),
    .X(_1469_));
 sg13g2_a22oi_1 _3285_ (.Y(_1470_),
    .B1(\u_ddc_top_level.cic_out_right[1] ),
    .B2(\u_ddc_top_level.cic_right_inst.int_reg1[13] ),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg1[12] ),
    .A1(\u_ddc_top_level.cic_out_right[0] ));
 sg13g2_a21oi_1 _3286_ (.A1(_1464_),
    .A2(_1470_),
    .Y(_1471_),
    .B1(_1465_));
 sg13g2_xor2_1 _3287_ (.B(_1471_),
    .A(_1469_),
    .X(_0088_));
 sg13g2_nand2_1 _3288_ (.Y(_1472_),
    .A(\u_ddc_top_level.cic_out_right[3] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[15] ));
 sg13g2_xor2_1 _3289_ (.B(\u_ddc_top_level.cic_right_inst.int_reg1[15] ),
    .A(\u_ddc_top_level.cic_out_right[3] ),
    .X(_1473_));
 sg13g2_a21oi_1 _3290_ (.A1(_1469_),
    .A2(_1471_),
    .Y(_1474_),
    .B1(_1468_));
 sg13g2_xnor2_1 _3291_ (.Y(_0089_),
    .A(_1473_),
    .B(_1474_));
 sg13g2_and4_1 _3292_ (.A(_1463_),
    .B(_1466_),
    .C(_1469_),
    .D(_1473_),
    .X(_1475_));
 sg13g2_o21ai_1 _3293_ (.B1(_1468_),
    .Y(_1476_),
    .A1(\u_ddc_top_level.cic_out_right[3] ),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg1[15] ));
 sg13g2_nor2_1 _3294_ (.A(_1465_),
    .B(_1470_),
    .Y(_1477_));
 sg13g2_nand3_1 _3295_ (.B(_1473_),
    .C(_1477_),
    .A(_1469_),
    .Y(_1478_));
 sg13g2_nand3_1 _3296_ (.B(_1476_),
    .C(_1478_),
    .A(_1472_),
    .Y(_1479_));
 sg13g2_a21oi_2 _3297_ (.B1(_1479_),
    .Y(_1480_),
    .A2(_1475_),
    .A1(_1461_));
 sg13g2_a21o_1 _3298_ (.A2(_1475_),
    .A1(_1461_),
    .B1(_1479_),
    .X(_1481_));
 sg13g2_nand2_1 _3299_ (.Y(_1482_),
    .A(\u_ddc_top_level.cic_out_right[4] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[16] ));
 sg13g2_xnor2_1 _3300_ (.Y(_1483_),
    .A(\u_ddc_top_level.cic_out_right[4] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[16] ));
 sg13g2_xnor2_1 _3301_ (.Y(_0090_),
    .A(_1481_),
    .B(_1483_));
 sg13g2_nor2_1 _3302_ (.A(\u_ddc_top_level.cic_out_right[5] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[17] ),
    .Y(_1484_));
 sg13g2_nand2_1 _3303_ (.Y(_1485_),
    .A(\u_ddc_top_level.cic_out_right[5] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[17] ));
 sg13g2_nand2b_1 _3304_ (.Y(_1486_),
    .B(_1485_),
    .A_N(_1484_));
 sg13g2_o21ai_1 _3305_ (.B1(_1482_),
    .Y(_1487_),
    .A1(_1480_),
    .A2(_1483_));
 sg13g2_xnor2_1 _3306_ (.Y(_0091_),
    .A(_1486_),
    .B(_1487_));
 sg13g2_and2_1 _3307_ (.A(\u_ddc_top_level.cic_out_right[6] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[18] ),
    .X(_1488_));
 sg13g2_xor2_1 _3308_ (.B(\u_ddc_top_level.cic_right_inst.int_reg1[18] ),
    .A(\u_ddc_top_level.cic_out_right[6] ),
    .X(_1489_));
 sg13g2_inv_1 _3309_ (.Y(_1490_),
    .A(_1489_));
 sg13g2_o21ai_1 _3310_ (.B1(_1485_),
    .Y(_1491_),
    .A1(_1482_),
    .A2(_1484_));
 sg13g2_or2_1 _3311_ (.X(_1492_),
    .B(_1486_),
    .A(_1483_));
 sg13g2_nor2_1 _3312_ (.A(_1480_),
    .B(_1492_),
    .Y(_1493_));
 sg13g2_or2_1 _3313_ (.X(_1494_),
    .B(_1493_),
    .A(_1491_));
 sg13g2_xnor2_1 _3314_ (.Y(_0092_),
    .A(_1490_),
    .B(_1494_));
 sg13g2_or2_1 _3315_ (.X(_1495_),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[19] ),
    .A(\u_ddc_top_level.cic_out_right[7] ));
 sg13g2_and2_1 _3316_ (.A(\u_ddc_top_level.cic_out_right[7] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[19] ),
    .X(_1496_));
 sg13g2_xnor2_1 _3317_ (.Y(_1497_),
    .A(\u_ddc_top_level.cic_out_right[7] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[19] ));
 sg13g2_a21oi_1 _3318_ (.A1(_1489_),
    .A2(_1494_),
    .Y(_1498_),
    .B1(_1488_));
 sg13g2_xor2_1 _3319_ (.B(_1498_),
    .A(_1497_),
    .X(_0093_));
 sg13g2_xnor2_1 _3320_ (.Y(_1499_),
    .A(\u_ddc_top_level.cic_out_right[8] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[20] ));
 sg13g2_nor2_1 _3321_ (.A(_1490_),
    .B(_1497_),
    .Y(_1500_));
 sg13g2_a221oi_1 _3322_ (.B2(_1491_),
    .C1(_1496_),
    .B1(_1500_),
    .A1(_1488_),
    .Y(_1501_),
    .A2(_1495_));
 sg13g2_nand2b_1 _3323_ (.Y(_1502_),
    .B(_1500_),
    .A_N(_1492_));
 sg13g2_o21ai_1 _3324_ (.B1(_1501_),
    .Y(_1503_),
    .A1(_1480_),
    .A2(_1502_));
 sg13g2_nor2b_1 _3325_ (.A(_1499_),
    .B_N(_1503_),
    .Y(_1504_));
 sg13g2_xnor2_1 _3326_ (.Y(_0095_),
    .A(_1499_),
    .B(_1503_));
 sg13g2_nor2_1 _3327_ (.A(\u_ddc_top_level.cic_out_right[9] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[21] ),
    .Y(_1505_));
 sg13g2_xor2_1 _3328_ (.B(\u_ddc_top_level.cic_right_inst.int_reg1[21] ),
    .A(\u_ddc_top_level.cic_out_right[9] ),
    .X(_1506_));
 sg13g2_a21oi_1 _3329_ (.A1(\u_ddc_top_level.cic_out_right[8] ),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg1[20] ),
    .Y(_1507_),
    .B1(_1504_));
 sg13g2_xnor2_1 _3330_ (.Y(_0096_),
    .A(_1506_),
    .B(_1507_));
 sg13g2_nand2_1 _3331_ (.Y(_1508_),
    .A(\u_ddc_top_level.cic_out_right[10] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[22] ));
 sg13g2_xnor2_1 _3332_ (.Y(_1509_),
    .A(\u_ddc_top_level.cic_out_right[10] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg1[22] ));
 sg13g2_nor2b_1 _3333_ (.A(_1499_),
    .B_N(_1506_),
    .Y(_1510_));
 sg13g2_a22oi_1 _3334_ (.Y(_1511_),
    .B1(\u_ddc_top_level.cic_out_right[9] ),
    .B2(\u_ddc_top_level.cic_right_inst.int_reg1[21] ),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg1[20] ),
    .A1(\u_ddc_top_level.cic_out_right[8] ));
 sg13g2_nor2_1 _3335_ (.A(_1505_),
    .B(_1511_),
    .Y(_1512_));
 sg13g2_a21oi_1 _3336_ (.A1(_1503_),
    .A2(_1510_),
    .Y(_1513_),
    .B1(_1512_));
 sg13g2_xor2_1 _3337_ (.B(_1513_),
    .A(_1509_),
    .X(_0097_));
 sg13g2_nor2_1 _3338_ (.A(\u_ddc_top_level.cic_out_right[11] ),
    .B(net884),
    .Y(_1514_));
 sg13g2_xnor2_1 _3339_ (.Y(_1515_),
    .A(\u_ddc_top_level.cic_out_right[11] ),
    .B(net884));
 sg13g2_o21ai_1 _3340_ (.B1(_1508_),
    .Y(_1516_),
    .A1(_1509_),
    .A2(_1513_));
 sg13g2_xnor2_1 _3341_ (.Y(_0098_),
    .A(_1515_),
    .B(_1516_));
 sg13g2_nor2_1 _3342_ (.A(_1509_),
    .B(_1515_),
    .Y(_1517_));
 sg13g2_and2_1 _3343_ (.A(_1510_),
    .B(_1517_),
    .X(_1518_));
 sg13g2_inv_1 _3344_ (.Y(_1519_),
    .A(_1518_));
 sg13g2_nor2_1 _3345_ (.A(_1502_),
    .B(_1519_),
    .Y(_1520_));
 sg13g2_nor2_1 _3346_ (.A(_1508_),
    .B(_1514_),
    .Y(_1521_));
 sg13g2_a221oi_1 _3347_ (.B2(_1517_),
    .C1(_1521_),
    .B1(_1512_),
    .A1(\u_ddc_top_level.cic_out_right[11] ),
    .Y(_1522_),
    .A2(net884));
 sg13g2_o21ai_1 _3348_ (.B1(_1522_),
    .Y(_1523_),
    .A1(_1501_),
    .A2(_1519_));
 sg13g2_a21oi_2 _3349_ (.B1(_1523_),
    .Y(_1524_),
    .A2(_1520_),
    .A1(_1481_));
 sg13g2_xor2_1 _3350_ (.B(\u_ddc_top_level.cic_out_right[12] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[23] ),
    .X(_1525_));
 sg13g2_nor2b_1 _3351_ (.A(_1524_),
    .B_N(_1525_),
    .Y(_1526_));
 sg13g2_xnor2_1 _3352_ (.Y(_0099_),
    .A(_1524_),
    .B(_1525_));
 sg13g2_xor2_1 _3353_ (.B(\u_ddc_top_level.cic_out_right[13] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[23] ),
    .X(_1527_));
 sg13g2_a21oi_1 _3354_ (.A1(\u_ddc_top_level.cic_right_inst.int_reg1[23] ),
    .A2(\u_ddc_top_level.cic_out_right[12] ),
    .Y(_1528_),
    .B1(_1526_));
 sg13g2_xnor2_1 _3355_ (.Y(_0100_),
    .A(_1527_),
    .B(_1528_));
 sg13g2_nand2_1 _3356_ (.Y(_1529_),
    .A(_1525_),
    .B(_1527_));
 sg13g2_o21ai_1 _3357_ (.B1(net884),
    .Y(_1530_),
    .A1(\u_ddc_top_level.cic_out_right[12] ),
    .A2(\u_ddc_top_level.cic_out_right[13] ));
 sg13g2_o21ai_1 _3358_ (.B1(_1530_),
    .Y(_1531_),
    .A1(_1524_),
    .A2(_1529_));
 sg13g2_and2_1 _3359_ (.A(net884),
    .B(\u_ddc_top_level.cic_out_right[14] ),
    .X(_1532_));
 sg13g2_or2_1 _3360_ (.X(_1533_),
    .B(\u_ddc_top_level.cic_out_right[14] ),
    .A(net884));
 sg13g2_nand2b_1 _3361_ (.Y(_1534_),
    .B(_1533_),
    .A_N(_1532_));
 sg13g2_xnor2_1 _3362_ (.Y(_0101_),
    .A(_1531_),
    .B(_1534_));
 sg13g2_a21oi_1 _3363_ (.A1(_1531_),
    .A2(_1533_),
    .Y(_1535_),
    .B1(_1532_));
 sg13g2_xor2_1 _3364_ (.B(\u_ddc_top_level.cic_out_right[15] ),
    .A(net884),
    .X(_1536_));
 sg13g2_xnor2_1 _3365_ (.Y(_0102_),
    .A(_1535_),
    .B(_1536_));
 sg13g2_nand2_1 _3366_ (.Y(_1537_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[0] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[0] ));
 sg13g2_xor2_1 _3367_ (.B(\u_ddc_top_level.cic_right_inst.int_reg0[0] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[0] ),
    .X(_0059_));
 sg13g2_nand2_1 _3368_ (.Y(_1538_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[1] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[1] ));
 sg13g2_nor2_1 _3369_ (.A(\u_ddc_top_level.cic_right_inst.int_reg1[1] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[1] ),
    .Y(_1539_));
 sg13g2_xor2_1 _3370_ (.B(\u_ddc_top_level.cic_right_inst.int_reg0[1] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[1] ),
    .X(_1540_));
 sg13g2_xnor2_1 _3371_ (.Y(_0070_),
    .A(_1537_),
    .B(_1540_));
 sg13g2_o21ai_1 _3372_ (.B1(_1538_),
    .Y(_1541_),
    .A1(_1537_),
    .A2(_1539_));
 sg13g2_and2_1 _3373_ (.A(\u_ddc_top_level.cic_right_inst.int_reg1[2] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[2] ),
    .X(_1542_));
 sg13g2_or2_1 _3374_ (.X(_1543_),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[2] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[2] ));
 sg13g2_nand2b_1 _3375_ (.Y(_1544_),
    .B(_1543_),
    .A_N(_1542_));
 sg13g2_xnor2_1 _3376_ (.Y(_0075_),
    .A(_1541_),
    .B(_1544_));
 sg13g2_a21o_1 _3377_ (.A2(_1543_),
    .A1(_1541_),
    .B1(_1542_),
    .X(_1545_));
 sg13g2_and2_1 _3378_ (.A(\u_ddc_top_level.cic_right_inst.int_reg1[3] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[3] ),
    .X(_1546_));
 sg13g2_or2_1 _3379_ (.X(_1547_),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[3] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[3] ));
 sg13g2_nand2b_1 _3380_ (.Y(_1548_),
    .B(_1547_),
    .A_N(_1546_));
 sg13g2_xnor2_1 _3381_ (.Y(_0076_),
    .A(_1545_),
    .B(_1548_));
 sg13g2_a21o_1 _3382_ (.A2(_1547_),
    .A1(_1545_),
    .B1(_1546_),
    .X(_1549_));
 sg13g2_xnor2_1 _3383_ (.Y(_1550_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[4] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[4] ));
 sg13g2_nor2b_1 _3384_ (.A(_1550_),
    .B_N(_1549_),
    .Y(_1551_));
 sg13g2_xnor2_1 _3385_ (.Y(_0077_),
    .A(_1549_),
    .B(_1550_));
 sg13g2_nor2_1 _3386_ (.A(\u_ddc_top_level.cic_right_inst.int_reg1[5] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[5] ),
    .Y(_1552_));
 sg13g2_xnor2_1 _3387_ (.Y(_1553_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[5] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[5] ));
 sg13g2_a21oi_1 _3388_ (.A1(\u_ddc_top_level.cic_right_inst.int_reg1[4] ),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg0[4] ),
    .Y(_1554_),
    .B1(_1551_));
 sg13g2_xor2_1 _3389_ (.B(_1554_),
    .A(_1553_),
    .X(_0078_));
 sg13g2_nand2_1 _3390_ (.Y(_1555_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[6] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[6] ));
 sg13g2_nor2_1 _3391_ (.A(\u_ddc_top_level.cic_right_inst.int_reg1[6] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[6] ),
    .Y(_1556_));
 sg13g2_xor2_1 _3392_ (.B(\u_ddc_top_level.cic_right_inst.int_reg0[6] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[6] ),
    .X(_1557_));
 sg13g2_a22oi_1 _3393_ (.Y(_1558_),
    .B1(\u_ddc_top_level.cic_right_inst.int_reg0[5] ),
    .B2(\u_ddc_top_level.cic_right_inst.int_reg1[5] ),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg0[4] ),
    .A1(\u_ddc_top_level.cic_right_inst.int_reg1[4] ));
 sg13g2_nor2_1 _3394_ (.A(_1550_),
    .B(_1553_),
    .Y(_1559_));
 sg13g2_nor2_1 _3395_ (.A(_1552_),
    .B(_1558_),
    .Y(_1560_));
 sg13g2_a21oi_1 _3396_ (.A1(_1549_),
    .A2(_1559_),
    .Y(_1561_),
    .B1(_1560_));
 sg13g2_xnor2_1 _3397_ (.Y(_0079_),
    .A(_1557_),
    .B(_1561_));
 sg13g2_nor2_1 _3398_ (.A(\u_ddc_top_level.cic_right_inst.int_reg1[7] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[7] ),
    .Y(_1562_));
 sg13g2_nand2_1 _3399_ (.Y(_1563_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[7] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[7] ));
 sg13g2_nand2b_1 _3400_ (.Y(_1564_),
    .B(_1563_),
    .A_N(_1562_));
 sg13g2_o21ai_1 _3401_ (.B1(_1555_),
    .Y(_1565_),
    .A1(_1556_),
    .A2(_1561_));
 sg13g2_xnor2_1 _3402_ (.Y(_0080_),
    .A(_1564_),
    .B(_1565_));
 sg13g2_nand2_1 _3403_ (.Y(_1566_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[8] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[8] ));
 sg13g2_xor2_1 _3404_ (.B(\u_ddc_top_level.cic_right_inst.int_reg0[8] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[8] ),
    .X(_1567_));
 sg13g2_inv_1 _3405_ (.Y(_1568_),
    .A(_1567_));
 sg13g2_a21oi_1 _3406_ (.A1(_1556_),
    .A2(_1563_),
    .Y(_1569_),
    .B1(_1562_));
 sg13g2_o21ai_1 _3407_ (.B1(_1563_),
    .Y(_1570_),
    .A1(_1555_),
    .A2(_1562_));
 sg13g2_or2_1 _3408_ (.X(_1571_),
    .B(_1570_),
    .A(_1560_));
 sg13g2_a21oi_1 _3409_ (.A1(_1549_),
    .A2(_1559_),
    .Y(_1572_),
    .B1(_1571_));
 sg13g2_nor2b_1 _3410_ (.A(_1572_),
    .B_N(_1569_),
    .Y(_1573_));
 sg13g2_nand2_1 _3411_ (.Y(_1574_),
    .A(_1567_),
    .B(_1573_));
 sg13g2_xnor2_1 _3412_ (.Y(_0081_),
    .A(_1568_),
    .B(_1573_));
 sg13g2_nor2_1 _3413_ (.A(\u_ddc_top_level.cic_right_inst.int_reg1[9] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[9] ),
    .Y(_1575_));
 sg13g2_xnor2_1 _3414_ (.Y(_1576_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[9] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[9] ));
 sg13g2_nand2_1 _3415_ (.Y(_1577_),
    .A(_1566_),
    .B(_1574_));
 sg13g2_xnor2_1 _3416_ (.Y(_0082_),
    .A(_1576_),
    .B(_1577_));
 sg13g2_and2_1 _3417_ (.A(\u_ddc_top_level.cic_right_inst.int_reg1[10] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[10] ),
    .X(_1578_));
 sg13g2_xor2_1 _3418_ (.B(\u_ddc_top_level.cic_right_inst.int_reg0[10] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[10] ),
    .X(_1579_));
 sg13g2_a22oi_1 _3419_ (.Y(_1580_),
    .B1(\u_ddc_top_level.cic_right_inst.int_reg0[9] ),
    .B2(\u_ddc_top_level.cic_right_inst.int_reg1[9] ),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg0[8] ),
    .A1(\u_ddc_top_level.cic_right_inst.int_reg1[8] ));
 sg13g2_a21oi_1 _3420_ (.A1(_1574_),
    .A2(_1580_),
    .Y(_1581_),
    .B1(_1575_));
 sg13g2_xor2_1 _3421_ (.B(_1581_),
    .A(_1579_),
    .X(_0060_));
 sg13g2_nand2_1 _3422_ (.Y(_1582_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[11] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[11] ));
 sg13g2_xor2_1 _3423_ (.B(\u_ddc_top_level.cic_right_inst.int_reg0[11] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[11] ),
    .X(_1583_));
 sg13g2_a21oi_1 _3424_ (.A1(_1579_),
    .A2(_1581_),
    .Y(_1584_),
    .B1(_1578_));
 sg13g2_xnor2_1 _3425_ (.Y(_0061_),
    .A(_1583_),
    .B(_1584_));
 sg13g2_nand2_1 _3426_ (.Y(_1585_),
    .A(_1579_),
    .B(_1583_));
 sg13g2_nor3_1 _3427_ (.A(_1568_),
    .B(_1576_),
    .C(_1585_),
    .Y(_1586_));
 sg13g2_nand3b_1 _3428_ (.B(_1586_),
    .C(_1569_),
    .Y(_1587_),
    .A_N(_1572_));
 sg13g2_o21ai_1 _3429_ (.B1(_1578_),
    .Y(_1588_),
    .A1(\u_ddc_top_level.cic_right_inst.int_reg1[11] ),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg0[11] ));
 sg13g2_or3_1 _3430_ (.A(_1575_),
    .B(_1580_),
    .C(_1585_),
    .X(_1589_));
 sg13g2_nand3_1 _3431_ (.B(_1588_),
    .C(_1589_),
    .A(_1582_),
    .Y(_1590_));
 sg13g2_inv_1 _3432_ (.Y(_1591_),
    .A(_1590_));
 sg13g2_nand2_1 _3433_ (.Y(_1592_),
    .A(_1587_),
    .B(_1591_));
 sg13g2_nand2_1 _3434_ (.Y(_1593_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[12] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[12] ));
 sg13g2_xor2_1 _3435_ (.B(\u_ddc_top_level.cic_right_inst.int_reg0[12] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[12] ),
    .X(_1594_));
 sg13g2_nand2_1 _3436_ (.Y(_1595_),
    .A(_1592_),
    .B(_1594_));
 sg13g2_xor2_1 _3437_ (.B(_1594_),
    .A(_1592_),
    .X(_0062_));
 sg13g2_nor2_1 _3438_ (.A(\u_ddc_top_level.cic_right_inst.int_reg1[13] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[13] ),
    .Y(_1596_));
 sg13g2_xor2_1 _3439_ (.B(\u_ddc_top_level.cic_right_inst.int_reg0[13] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[13] ),
    .X(_1597_));
 sg13g2_nand2_1 _3440_ (.Y(_1598_),
    .A(_1593_),
    .B(_1595_));
 sg13g2_xor2_1 _3441_ (.B(_1598_),
    .A(_1597_),
    .X(_0063_));
 sg13g2_and2_1 _3442_ (.A(\u_ddc_top_level.cic_right_inst.int_reg1[14] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[14] ),
    .X(_1599_));
 sg13g2_xor2_1 _3443_ (.B(\u_ddc_top_level.cic_right_inst.int_reg0[14] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[14] ),
    .X(_1600_));
 sg13g2_a22oi_1 _3444_ (.Y(_1601_),
    .B1(\u_ddc_top_level.cic_right_inst.int_reg0[13] ),
    .B2(\u_ddc_top_level.cic_right_inst.int_reg1[13] ),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg0[12] ),
    .A1(\u_ddc_top_level.cic_right_inst.int_reg1[12] ));
 sg13g2_a21oi_1 _3445_ (.A1(_1595_),
    .A2(_1601_),
    .Y(_1602_),
    .B1(_1596_));
 sg13g2_xor2_1 _3446_ (.B(_1602_),
    .A(_1600_),
    .X(_0064_));
 sg13g2_nand2_1 _3447_ (.Y(_1603_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[15] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[15] ));
 sg13g2_xor2_1 _3448_ (.B(\u_ddc_top_level.cic_right_inst.int_reg0[15] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[15] ),
    .X(_1604_));
 sg13g2_a21oi_1 _3449_ (.A1(_1600_),
    .A2(_1602_),
    .Y(_1605_),
    .B1(_1599_));
 sg13g2_xnor2_1 _3450_ (.Y(_0065_),
    .A(_1604_),
    .B(_1605_));
 sg13g2_nand4_1 _3451_ (.B(_1597_),
    .C(_1600_),
    .A(_1594_),
    .Y(_1606_),
    .D(_1604_));
 sg13g2_a21oi_2 _3452_ (.B1(_1606_),
    .Y(_1607_),
    .A2(_1591_),
    .A1(_1587_));
 sg13g2_o21ai_1 _3453_ (.B1(_1599_),
    .Y(_1608_),
    .A1(\u_ddc_top_level.cic_right_inst.int_reg1[15] ),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg0[15] ));
 sg13g2_nor2_1 _3454_ (.A(_1596_),
    .B(_1601_),
    .Y(_1609_));
 sg13g2_nand3_1 _3455_ (.B(_1604_),
    .C(_1609_),
    .A(_1600_),
    .Y(_1610_));
 sg13g2_nand3_1 _3456_ (.B(_1608_),
    .C(_1610_),
    .A(_1603_),
    .Y(_1611_));
 sg13g2_nand2_1 _3457_ (.Y(_1612_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[16] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[16] ));
 sg13g2_xor2_1 _3458_ (.B(\u_ddc_top_level.cic_right_inst.int_reg0[16] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[16] ),
    .X(_1613_));
 sg13g2_o21ai_1 _3459_ (.B1(_1613_),
    .Y(_1614_),
    .A1(_1607_),
    .A2(_1611_));
 sg13g2_or3_1 _3460_ (.A(_1607_),
    .B(_1611_),
    .C(_1613_),
    .X(_1615_));
 sg13g2_and2_1 _3461_ (.A(_1614_),
    .B(_1615_),
    .X(_0066_));
 sg13g2_nor2_1 _3462_ (.A(\u_ddc_top_level.cic_right_inst.int_reg1[17] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[17] ),
    .Y(_1616_));
 sg13g2_xnor2_1 _3463_ (.Y(_1617_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[17] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[17] ));
 sg13g2_nand2_1 _3464_ (.Y(_1618_),
    .A(_1612_),
    .B(_1614_));
 sg13g2_xnor2_1 _3465_ (.Y(_0067_),
    .A(_1617_),
    .B(_1618_));
 sg13g2_and2_1 _3466_ (.A(\u_ddc_top_level.cic_right_inst.int_reg1[18] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[18] ),
    .X(_1619_));
 sg13g2_xor2_1 _3467_ (.B(\u_ddc_top_level.cic_right_inst.int_reg0[18] ),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[18] ),
    .X(_1620_));
 sg13g2_a22oi_1 _3468_ (.Y(_1621_),
    .B1(\u_ddc_top_level.cic_right_inst.int_reg0[17] ),
    .B2(\u_ddc_top_level.cic_right_inst.int_reg1[17] ),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg0[16] ),
    .A1(\u_ddc_top_level.cic_right_inst.int_reg1[16] ));
 sg13g2_a21oi_1 _3469_ (.A1(_1614_),
    .A2(_1621_),
    .Y(_1622_),
    .B1(_1616_));
 sg13g2_xor2_1 _3470_ (.B(_1622_),
    .A(_1620_),
    .X(_0068_));
 sg13g2_nand2_1 _3471_ (.Y(_1623_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[19] ),
    .B(net882));
 sg13g2_xor2_1 _3472_ (.B(net882),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[19] ),
    .X(_1624_));
 sg13g2_a21oi_1 _3473_ (.A1(_1620_),
    .A2(_1622_),
    .Y(_1625_),
    .B1(_1619_));
 sg13g2_xnor2_1 _3474_ (.Y(_0069_),
    .A(_1624_),
    .B(_1625_));
 sg13g2_nand3_1 _3475_ (.B(_1620_),
    .C(_1624_),
    .A(_1613_),
    .Y(_1626_));
 sg13g2_nor2_1 _3476_ (.A(_1617_),
    .B(_1626_),
    .Y(_1627_));
 sg13g2_o21ai_1 _3477_ (.B1(_1627_),
    .Y(_1628_),
    .A1(_1607_),
    .A2(_1611_));
 sg13g2_o21ai_1 _3478_ (.B1(_1619_),
    .Y(_1629_),
    .A1(\u_ddc_top_level.cic_right_inst.int_reg1[19] ),
    .A2(net882));
 sg13g2_nor2_1 _3479_ (.A(_1616_),
    .B(_1621_),
    .Y(_1630_));
 sg13g2_nand3_1 _3480_ (.B(_1624_),
    .C(_1630_),
    .A(_1620_),
    .Y(_1631_));
 sg13g2_and4_1 _3481_ (.A(_1623_),
    .B(_1628_),
    .C(_1629_),
    .D(_1631_),
    .X(_1632_));
 sg13g2_nand2_1 _3482_ (.Y(_1633_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[20] ),
    .B(net883));
 sg13g2_xnor2_1 _3483_ (.Y(_1634_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[20] ),
    .B(net883));
 sg13g2_xor2_1 _3484_ (.B(_1634_),
    .A(_1632_),
    .X(_0071_));
 sg13g2_xor2_1 _3485_ (.B(net883),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[21] ),
    .X(_1635_));
 sg13g2_o21ai_1 _3486_ (.B1(_1633_),
    .Y(_1636_),
    .A1(_1632_),
    .A2(_1634_));
 sg13g2_xor2_1 _3487_ (.B(_1636_),
    .A(_1635_),
    .X(_0072_));
 sg13g2_and2_1 _3488_ (.A(\u_ddc_top_level.cic_right_inst.int_reg1[22] ),
    .B(net883),
    .X(_1637_));
 sg13g2_or2_1 _3489_ (.X(_1638_),
    .B(net882),
    .A(\u_ddc_top_level.cic_right_inst.int_reg1[22] ));
 sg13g2_nand2b_1 _3490_ (.Y(_1639_),
    .B(_1638_),
    .A_N(_1637_));
 sg13g2_nand2b_1 _3491_ (.Y(_1640_),
    .B(_1635_),
    .A_N(_1634_));
 sg13g2_o21ai_1 _3492_ (.B1(net882),
    .Y(_1641_),
    .A1(\u_ddc_top_level.cic_right_inst.int_reg1[20] ),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg1[21] ));
 sg13g2_o21ai_1 _3493_ (.B1(_1641_),
    .Y(_1642_),
    .A1(_1632_),
    .A2(_1640_));
 sg13g2_xnor2_1 _3494_ (.Y(_0073_),
    .A(_1639_),
    .B(_1642_));
 sg13g2_a21oi_1 _3495_ (.A1(_1638_),
    .A2(_1642_),
    .Y(_1643_),
    .B1(_1637_));
 sg13g2_xor2_1 _3496_ (.B(net882),
    .A(net884),
    .X(_1644_));
 sg13g2_xnor2_1 _3497_ (.Y(_0074_),
    .A(_1643_),
    .B(_1644_));
 sg13g2_nand2_1 _3498_ (.Y(_1645_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[0] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[0] ));
 sg13g2_nand2_1 _3499_ (.Y(_1646_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[1] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[1] ));
 sg13g2_nor2_1 _3500_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[1] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[1] ),
    .Y(_1647_));
 sg13g2_xor2_1 _3501_ (.B(\u_ddc_top_level.cic_left_inst.int_reg0[1] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[1] ),
    .X(_1648_));
 sg13g2_xnor2_1 _3502_ (.Y(_0018_),
    .A(_1645_),
    .B(_1648_));
 sg13g2_o21ai_1 _3503_ (.B1(_1646_),
    .Y(_1649_),
    .A1(_1645_),
    .A2(_1647_));
 sg13g2_and2_1 _3504_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[2] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[2] ),
    .X(_1650_));
 sg13g2_or2_1 _3505_ (.X(_1651_),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[2] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[2] ));
 sg13g2_nand2b_1 _3506_ (.Y(_1652_),
    .B(_1651_),
    .A_N(_1650_));
 sg13g2_xnor2_1 _3507_ (.Y(_0023_),
    .A(_1649_),
    .B(_1652_));
 sg13g2_a21o_1 _3508_ (.A2(_1651_),
    .A1(_1649_),
    .B1(_1650_),
    .X(_1653_));
 sg13g2_and2_1 _3509_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[3] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[3] ),
    .X(_1654_));
 sg13g2_or2_1 _3510_ (.X(_1655_),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[3] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[3] ));
 sg13g2_nand2b_1 _3511_ (.Y(_1656_),
    .B(_1655_),
    .A_N(_1654_));
 sg13g2_xnor2_1 _3512_ (.Y(_0024_),
    .A(_1653_),
    .B(_1656_));
 sg13g2_a21o_1 _3513_ (.A2(_1655_),
    .A1(_1653_),
    .B1(_1654_),
    .X(_1657_));
 sg13g2_xnor2_1 _3514_ (.Y(_1658_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[4] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[4] ));
 sg13g2_nor2b_1 _3515_ (.A(_1658_),
    .B_N(_1657_),
    .Y(_1659_));
 sg13g2_xnor2_1 _3516_ (.Y(_0025_),
    .A(_1657_),
    .B(_1658_));
 sg13g2_nor2_1 _3517_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[5] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[5] ),
    .Y(_1660_));
 sg13g2_xnor2_1 _3518_ (.Y(_1661_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[5] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[5] ));
 sg13g2_a21oi_1 _3519_ (.A1(\u_ddc_top_level.cic_left_inst.int_reg1[4] ),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg0[4] ),
    .Y(_1662_),
    .B1(_1659_));
 sg13g2_xor2_1 _3520_ (.B(_1662_),
    .A(_1661_),
    .X(_0026_));
 sg13g2_nand2_1 _3521_ (.Y(_1663_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[6] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[6] ));
 sg13g2_nor2_1 _3522_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[6] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[6] ),
    .Y(_1664_));
 sg13g2_xor2_1 _3523_ (.B(\u_ddc_top_level.cic_left_inst.int_reg0[6] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[6] ),
    .X(_1665_));
 sg13g2_a22oi_1 _3524_ (.Y(_1666_),
    .B1(\u_ddc_top_level.cic_left_inst.int_reg1[5] ),
    .B2(\u_ddc_top_level.cic_left_inst.int_reg0[5] ),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg0[4] ),
    .A1(\u_ddc_top_level.cic_left_inst.int_reg1[4] ));
 sg13g2_nor2_1 _3525_ (.A(_1658_),
    .B(_1661_),
    .Y(_1667_));
 sg13g2_nor2_1 _3526_ (.A(_1660_),
    .B(_1666_),
    .Y(_1668_));
 sg13g2_a21oi_1 _3527_ (.A1(_1657_),
    .A2(_1667_),
    .Y(_1669_),
    .B1(_1668_));
 sg13g2_xnor2_1 _3528_ (.Y(_0027_),
    .A(_1665_),
    .B(_1669_));
 sg13g2_nand2_1 _3529_ (.Y(_1670_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[7] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[7] ));
 sg13g2_nor2_1 _3530_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[7] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[7] ),
    .Y(_1671_));
 sg13g2_xnor2_1 _3531_ (.Y(_1672_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[7] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[7] ));
 sg13g2_o21ai_1 _3532_ (.B1(_1663_),
    .Y(_1673_),
    .A1(_1664_),
    .A2(_1669_));
 sg13g2_xnor2_1 _3533_ (.Y(_0028_),
    .A(_1672_),
    .B(_1673_));
 sg13g2_nand2_1 _3534_ (.Y(_1674_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[8] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[8] ));
 sg13g2_xor2_1 _3535_ (.B(\u_ddc_top_level.cic_left_inst.int_reg0[8] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[8] ),
    .X(_1675_));
 sg13g2_a21o_1 _3536_ (.A2(_1670_),
    .A1(_1664_),
    .B1(_1671_),
    .X(_1676_));
 sg13g2_o21ai_1 _3537_ (.B1(_1670_),
    .Y(_1677_),
    .A1(_1663_),
    .A2(_1671_));
 sg13g2_or2_1 _3538_ (.X(_1678_),
    .B(_1677_),
    .A(_1668_));
 sg13g2_a21oi_1 _3539_ (.A1(_1657_),
    .A2(_1667_),
    .Y(_1679_),
    .B1(_1678_));
 sg13g2_nor2_1 _3540_ (.A(_1676_),
    .B(_1679_),
    .Y(_1680_));
 sg13g2_nand2_1 _3541_ (.Y(_1681_),
    .A(_1675_),
    .B(_1680_));
 sg13g2_xor2_1 _3542_ (.B(_1680_),
    .A(_1675_),
    .X(_0029_));
 sg13g2_nand2_1 _3543_ (.Y(_1682_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[9] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[9] ));
 sg13g2_nor2_1 _3544_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[9] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[9] ),
    .Y(_1683_));
 sg13g2_xnor2_1 _3545_ (.Y(_1684_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[9] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[9] ));
 sg13g2_nand2_1 _3546_ (.Y(_1685_),
    .A(_1674_),
    .B(_1681_));
 sg13g2_xnor2_1 _3547_ (.Y(_0030_),
    .A(_1684_),
    .B(_1685_));
 sg13g2_and2_1 _3548_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[10] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[10] ),
    .X(_1686_));
 sg13g2_xor2_1 _3549_ (.B(\u_ddc_top_level.cic_left_inst.int_reg0[10] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[10] ),
    .X(_1687_));
 sg13g2_and2_1 _3550_ (.A(_1674_),
    .B(_1682_),
    .X(_1688_));
 sg13g2_a21oi_1 _3551_ (.A1(_1681_),
    .A2(_1688_),
    .Y(_1689_),
    .B1(_1683_));
 sg13g2_xor2_1 _3552_ (.B(_1689_),
    .A(_1687_),
    .X(_0008_));
 sg13g2_nand2_1 _3553_ (.Y(_1690_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[11] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[11] ));
 sg13g2_xor2_1 _3554_ (.B(\u_ddc_top_level.cic_left_inst.int_reg0[11] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[11] ),
    .X(_1691_));
 sg13g2_a21oi_1 _3555_ (.A1(_1687_),
    .A2(_1689_),
    .Y(_1692_),
    .B1(_1686_));
 sg13g2_xnor2_1 _3556_ (.Y(_0009_),
    .A(_1691_),
    .B(_1692_));
 sg13g2_nand3b_1 _3557_ (.B(_1675_),
    .C(_1682_),
    .Y(_1693_),
    .A_N(_1683_));
 sg13g2_nand2_1 _3558_ (.Y(_1694_),
    .A(_1687_),
    .B(_1691_));
 sg13g2_or4_2 _3559_ (.A(_1676_),
    .B(_1679_),
    .C(_1693_),
    .D(_1694_),
    .X(_1695_));
 sg13g2_o21ai_1 _3560_ (.B1(_1686_),
    .Y(_1696_),
    .A1(\u_ddc_top_level.cic_left_inst.int_reg1[11] ),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg0[11] ));
 sg13g2_or3_1 _3561_ (.A(_1683_),
    .B(_1688_),
    .C(_1694_),
    .X(_1697_));
 sg13g2_nand3_1 _3562_ (.B(_1696_),
    .C(_1697_),
    .A(_1690_),
    .Y(_1698_));
 sg13g2_inv_1 _3563_ (.Y(_1699_),
    .A(_1698_));
 sg13g2_nand2_1 _3564_ (.Y(_1700_),
    .A(_1695_),
    .B(_1699_));
 sg13g2_nand2_1 _3565_ (.Y(_1701_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[12] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[12] ));
 sg13g2_xor2_1 _3566_ (.B(\u_ddc_top_level.cic_left_inst.int_reg0[12] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[12] ),
    .X(_1702_));
 sg13g2_nand2_1 _3567_ (.Y(_1703_),
    .A(_1700_),
    .B(_1702_));
 sg13g2_xor2_1 _3568_ (.B(_1702_),
    .A(_1700_),
    .X(_0010_));
 sg13g2_nor2_1 _3569_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[13] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[13] ),
    .Y(_1704_));
 sg13g2_xor2_1 _3570_ (.B(\u_ddc_top_level.cic_left_inst.int_reg0[13] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[13] ),
    .X(_1705_));
 sg13g2_and2_1 _3571_ (.A(_1701_),
    .B(_1703_),
    .X(_1706_));
 sg13g2_xnor2_1 _3572_ (.Y(_0011_),
    .A(_1705_),
    .B(_1706_));
 sg13g2_nand2_1 _3573_ (.Y(_1707_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[14] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[14] ));
 sg13g2_xor2_1 _3574_ (.B(\u_ddc_top_level.cic_left_inst.int_reg0[14] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[14] ),
    .X(_1708_));
 sg13g2_a22oi_1 _3575_ (.Y(_1709_),
    .B1(\u_ddc_top_level.cic_left_inst.int_reg1[13] ),
    .B2(\u_ddc_top_level.cic_left_inst.int_reg0[13] ),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg0[12] ),
    .A1(\u_ddc_top_level.cic_left_inst.int_reg1[12] ));
 sg13g2_a21oi_1 _3576_ (.A1(_1703_),
    .A2(_1709_),
    .Y(_1710_),
    .B1(_1704_));
 sg13g2_nand2_1 _3577_ (.Y(_1711_),
    .A(_1708_),
    .B(_1710_));
 sg13g2_xor2_1 _3578_ (.B(_1710_),
    .A(_1708_),
    .X(_0012_));
 sg13g2_nor2_1 _3579_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[15] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[15] ),
    .Y(_1712_));
 sg13g2_nand2_1 _3580_ (.Y(_1713_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[15] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[15] ));
 sg13g2_nor2b_2 _3581_ (.A(_1712_),
    .B_N(_1713_),
    .Y(_1714_));
 sg13g2_nand2_1 _3582_ (.Y(_1715_),
    .A(_1707_),
    .B(_1711_));
 sg13g2_xor2_1 _3583_ (.B(_1715_),
    .A(_1714_),
    .X(_0013_));
 sg13g2_nand2_1 _3584_ (.Y(_1716_),
    .A(_1708_),
    .B(_1714_));
 sg13g2_nand4_1 _3585_ (.B(_1705_),
    .C(_1708_),
    .A(_1702_),
    .Y(_1717_),
    .D(_1714_));
 sg13g2_a21oi_2 _3586_ (.B1(_1717_),
    .Y(_1718_),
    .A2(_1699_),
    .A1(_1695_));
 sg13g2_o21ai_1 _3587_ (.B1(_1713_),
    .Y(_1719_),
    .A1(_1707_),
    .A2(_1712_));
 sg13g2_nor3_1 _3588_ (.A(_1704_),
    .B(_1709_),
    .C(_1716_),
    .Y(_1720_));
 sg13g2_or2_1 _3589_ (.X(_1721_),
    .B(_1720_),
    .A(_1719_));
 sg13g2_nor2_1 _3590_ (.A(_1718_),
    .B(_1721_),
    .Y(_1722_));
 sg13g2_nand2_1 _3591_ (.Y(_1723_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[16] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[16] ));
 sg13g2_xnor2_1 _3592_ (.Y(_1724_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[16] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[16] ));
 sg13g2_inv_1 _3593_ (.Y(_1725_),
    .A(_1724_));
 sg13g2_o21ai_1 _3594_ (.B1(_1725_),
    .Y(_1726_),
    .A1(_1718_),
    .A2(_1721_));
 sg13g2_xnor2_1 _3595_ (.Y(_0014_),
    .A(_1722_),
    .B(_1725_));
 sg13g2_nor2_1 _3596_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[17] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[17] ),
    .Y(_1727_));
 sg13g2_xnor2_1 _3597_ (.Y(_1728_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[17] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[17] ));
 sg13g2_nand2_1 _3598_ (.Y(_1729_),
    .A(_1723_),
    .B(_1726_));
 sg13g2_xnor2_1 _3599_ (.Y(_0015_),
    .A(_1728_),
    .B(_1729_));
 sg13g2_and2_1 _3600_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[18] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[18] ),
    .X(_1730_));
 sg13g2_xor2_1 _3601_ (.B(\u_ddc_top_level.cic_left_inst.int_reg0[18] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[18] ),
    .X(_1731_));
 sg13g2_a22oi_1 _3602_ (.Y(_1732_),
    .B1(\u_ddc_top_level.cic_left_inst.int_reg1[17] ),
    .B2(\u_ddc_top_level.cic_left_inst.int_reg0[17] ),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg0[16] ),
    .A1(\u_ddc_top_level.cic_left_inst.int_reg1[16] ));
 sg13g2_a21oi_1 _3603_ (.A1(_1726_),
    .A2(_1732_),
    .Y(_1733_),
    .B1(_1727_));
 sg13g2_xor2_1 _3604_ (.B(_1733_),
    .A(_1731_),
    .X(_0016_));
 sg13g2_nand2_1 _3605_ (.Y(_1734_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[19] ),
    .B(net880));
 sg13g2_xor2_1 _3606_ (.B(net880),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[19] ),
    .X(_1735_));
 sg13g2_a21oi_1 _3607_ (.A1(_1731_),
    .A2(_1733_),
    .Y(_1736_),
    .B1(_1730_));
 sg13g2_xnor2_1 _3608_ (.Y(_0017_),
    .A(_1735_),
    .B(_1736_));
 sg13g2_nand2_1 _3609_ (.Y(_1737_),
    .A(_1731_),
    .B(_1735_));
 sg13g2_nor3_1 _3610_ (.A(_1724_),
    .B(_1728_),
    .C(_1737_),
    .Y(_1738_));
 sg13g2_o21ai_1 _3611_ (.B1(_1738_),
    .Y(_1739_),
    .A1(_1718_),
    .A2(_1721_));
 sg13g2_o21ai_1 _3612_ (.B1(_1730_),
    .Y(_1740_),
    .A1(\u_ddc_top_level.cic_left_inst.int_reg1[19] ),
    .A2(net880));
 sg13g2_or3_1 _3613_ (.A(_1727_),
    .B(_1732_),
    .C(_1737_),
    .X(_1741_));
 sg13g2_and4_2 _3614_ (.A(_1734_),
    .B(_1739_),
    .C(_1740_),
    .D(_1741_),
    .X(_1742_));
 sg13g2_nand2_1 _3615_ (.Y(_1743_),
    .A(net879),
    .B(\u_ddc_top_level.cic_left_inst.int_reg1[20] ));
 sg13g2_xnor2_1 _3616_ (.Y(_1744_),
    .A(net879),
    .B(\u_ddc_top_level.cic_left_inst.int_reg1[20] ));
 sg13g2_xor2_1 _3617_ (.B(_1744_),
    .A(_1742_),
    .X(_0019_));
 sg13g2_xor2_1 _3618_ (.B(\u_ddc_top_level.cic_left_inst.int_reg1[21] ),
    .A(net879),
    .X(_1745_));
 sg13g2_o21ai_1 _3619_ (.B1(_1743_),
    .Y(_1746_),
    .A1(_1742_),
    .A2(_1744_));
 sg13g2_xor2_1 _3620_ (.B(_1746_),
    .A(_1745_),
    .X(_0020_));
 sg13g2_and2_1 _3621_ (.A(net879),
    .B(\u_ddc_top_level.cic_left_inst.int_reg1[22] ),
    .X(_1747_));
 sg13g2_or2_1 _3622_ (.X(_1748_),
    .B(\u_ddc_top_level.cic_left_inst.int_reg1[22] ),
    .A(net879));
 sg13g2_nand2b_1 _3623_ (.Y(_1749_),
    .B(_1748_),
    .A_N(_1747_));
 sg13g2_nand2b_1 _3624_ (.Y(_1750_),
    .B(_1745_),
    .A_N(_1744_));
 sg13g2_o21ai_1 _3625_ (.B1(net879),
    .Y(_1751_),
    .A1(\u_ddc_top_level.cic_left_inst.int_reg1[20] ),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg1[21] ));
 sg13g2_o21ai_1 _3626_ (.B1(_1751_),
    .Y(_1752_),
    .A1(_1742_),
    .A2(_1750_));
 sg13g2_xnor2_1 _3627_ (.Y(_0021_),
    .A(_1749_),
    .B(_1752_));
 sg13g2_a21oi_1 _3628_ (.A1(_1748_),
    .A2(_1752_),
    .Y(_1753_),
    .B1(_1747_));
 sg13g2_xor2_1 _3629_ (.B(\u_ddc_top_level.cic_left_inst.int_reg1[23] ),
    .A(net879),
    .X(_1754_));
 sg13g2_xnor2_1 _3630_ (.Y(_0022_),
    .A(_1753_),
    .B(_1754_));
 sg13g2_xor2_1 _3631_ (.B(\u_ddc_top_level.cic_left_inst.int_reg0[0] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[0] ),
    .X(_0007_));
 sg13g2_nand2_1 _3632_ (.Y(_1755_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[0] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[0] ));
 sg13g2_nand2_1 _3633_ (.Y(_1756_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[1] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[1] ));
 sg13g2_nor2_1 _3634_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[1] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[1] ),
    .Y(_1757_));
 sg13g2_xor2_1 _3635_ (.B(\u_ddc_top_level.cic_left_inst.int_reg2[1] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[1] ),
    .X(_1758_));
 sg13g2_xnor2_1 _3636_ (.Y(_0042_),
    .A(_1755_),
    .B(_1758_));
 sg13g2_o21ai_1 _3637_ (.B1(_1756_),
    .Y(_1759_),
    .A1(_1755_),
    .A2(_1757_));
 sg13g2_and2_1 _3638_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[2] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[2] ),
    .X(_1760_));
 sg13g2_or2_1 _3639_ (.X(_1761_),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[2] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[2] ));
 sg13g2_nand2b_1 _3640_ (.Y(_1762_),
    .B(_1761_),
    .A_N(_1760_));
 sg13g2_xnor2_1 _3641_ (.Y(_0051_),
    .A(_1759_),
    .B(_1762_));
 sg13g2_a21o_1 _3642_ (.A2(_1761_),
    .A1(_1759_),
    .B1(_1760_),
    .X(_1763_));
 sg13g2_and2_1 _3643_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[3] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[3] ),
    .X(_1764_));
 sg13g2_or2_1 _3644_ (.X(_1765_),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[3] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[3] ));
 sg13g2_nand2b_1 _3645_ (.Y(_1766_),
    .B(_1765_),
    .A_N(_1764_));
 sg13g2_xnor2_1 _3646_ (.Y(_0052_),
    .A(_1763_),
    .B(_1766_));
 sg13g2_a21o_1 _3647_ (.A2(_1765_),
    .A1(_1763_),
    .B1(_1764_),
    .X(_1767_));
 sg13g2_xnor2_1 _3648_ (.Y(_1768_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[4] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[4] ));
 sg13g2_nor2b_1 _3649_ (.A(_1768_),
    .B_N(_1767_),
    .Y(_1769_));
 sg13g2_xnor2_1 _3650_ (.Y(_0053_),
    .A(_1767_),
    .B(_1768_));
 sg13g2_nor2_1 _3651_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[5] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[5] ),
    .Y(_1770_));
 sg13g2_xnor2_1 _3652_ (.Y(_1771_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[5] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[5] ));
 sg13g2_a21oi_1 _3653_ (.A1(\u_ddc_top_level.cic_left_inst.int_reg1[4] ),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg2[4] ),
    .Y(_1772_),
    .B1(_1769_));
 sg13g2_xor2_1 _3654_ (.B(_1772_),
    .A(_1771_),
    .X(_0054_));
 sg13g2_nor2_1 _3655_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[6] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[6] ),
    .Y(_1773_));
 sg13g2_xor2_1 _3656_ (.B(\u_ddc_top_level.cic_left_inst.int_reg2[6] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[6] ),
    .X(_1774_));
 sg13g2_a22oi_1 _3657_ (.Y(_1775_),
    .B1(\u_ddc_top_level.cic_left_inst.int_reg2[5] ),
    .B2(\u_ddc_top_level.cic_left_inst.int_reg1[5] ),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg2[4] ),
    .A1(\u_ddc_top_level.cic_left_inst.int_reg1[4] ));
 sg13g2_nor2_1 _3658_ (.A(_1768_),
    .B(_1771_),
    .Y(_1776_));
 sg13g2_nor2_1 _3659_ (.A(_1770_),
    .B(_1775_),
    .Y(_1777_));
 sg13g2_a21oi_1 _3660_ (.A1(_1767_),
    .A2(_1776_),
    .Y(_1778_),
    .B1(_1777_));
 sg13g2_xnor2_1 _3661_ (.Y(_0055_),
    .A(_1774_),
    .B(_1778_));
 sg13g2_nand2_1 _3662_ (.Y(_1779_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[7] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[7] ));
 sg13g2_nor2_1 _3663_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[7] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[7] ),
    .Y(_1780_));
 sg13g2_xnor2_1 _3664_ (.Y(_1781_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[7] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[7] ));
 sg13g2_a221oi_1 _3665_ (.B2(_1776_),
    .C1(_1777_),
    .B1(_1767_),
    .A1(\u_ddc_top_level.cic_left_inst.int_reg1[6] ),
    .Y(_1782_),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg2[6] ));
 sg13g2_nor2_1 _3666_ (.A(_1773_),
    .B(_1782_),
    .Y(_1783_));
 sg13g2_xnor2_1 _3667_ (.Y(_0056_),
    .A(_1781_),
    .B(_1783_));
 sg13g2_xnor2_1 _3668_ (.Y(_1784_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[8] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[8] ));
 sg13g2_or2_1 _3669_ (.X(_1785_),
    .B(_1780_),
    .A(_1773_));
 sg13g2_o21ai_1 _3670_ (.B1(_1779_),
    .Y(_1786_),
    .A1(_1782_),
    .A2(_1785_));
 sg13g2_nor2b_1 _3671_ (.A(_1784_),
    .B_N(_1786_),
    .Y(_1787_));
 sg13g2_xnor2_1 _3672_ (.Y(_0057_),
    .A(_1784_),
    .B(_1786_));
 sg13g2_nor2_1 _3673_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[9] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[9] ),
    .Y(_1788_));
 sg13g2_xnor2_1 _3674_ (.Y(_1789_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[9] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[9] ));
 sg13g2_a21oi_1 _3675_ (.A1(\u_ddc_top_level.cic_left_inst.int_reg1[8] ),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg2[8] ),
    .Y(_1790_),
    .B1(_1787_));
 sg13g2_xor2_1 _3676_ (.B(_1790_),
    .A(_1789_),
    .X(_0058_));
 sg13g2_nand2_1 _3677_ (.Y(_1791_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[10] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[10] ));
 sg13g2_xnor2_1 _3678_ (.Y(_1792_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[10] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[10] ));
 sg13g2_a22oi_1 _3679_ (.Y(_1793_),
    .B1(\u_ddc_top_level.cic_left_inst.int_reg2[9] ),
    .B2(\u_ddc_top_level.cic_left_inst.int_reg1[9] ),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg2[8] ),
    .A1(\u_ddc_top_level.cic_left_inst.int_reg1[8] ));
 sg13g2_nor2_1 _3680_ (.A(_1788_),
    .B(_1793_),
    .Y(_1794_));
 sg13g2_nor2_1 _3681_ (.A(_1784_),
    .B(_1789_),
    .Y(_1795_));
 sg13g2_a21oi_1 _3682_ (.A1(_1786_),
    .A2(_1795_),
    .Y(_1796_),
    .B1(_1794_));
 sg13g2_xor2_1 _3683_ (.B(_1796_),
    .A(_1792_),
    .X(_0032_));
 sg13g2_nor2_1 _3684_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[11] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[11] ),
    .Y(_1797_));
 sg13g2_nand2_1 _3685_ (.Y(_1798_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[11] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[11] ));
 sg13g2_nor2b_1 _3686_ (.A(_1797_),
    .B_N(_1798_),
    .Y(_1799_));
 sg13g2_o21ai_1 _3687_ (.B1(_1791_),
    .Y(_1800_),
    .A1(_1792_),
    .A2(_1796_));
 sg13g2_xor2_1 _3688_ (.B(_1800_),
    .A(_1799_),
    .X(_0033_));
 sg13g2_nor2b_1 _3689_ (.A(_1792_),
    .B_N(_1799_),
    .Y(_1801_));
 sg13g2_and2_1 _3690_ (.A(_1795_),
    .B(_1801_),
    .X(_1802_));
 sg13g2_o21ai_1 _3691_ (.B1(_1798_),
    .Y(_1803_),
    .A1(_1791_),
    .A2(_1797_));
 sg13g2_a21o_1 _3692_ (.A2(_1801_),
    .A1(_1794_),
    .B1(_1803_),
    .X(_1804_));
 sg13g2_a21o_2 _3693_ (.A2(_1802_),
    .A1(_1786_),
    .B1(_1804_),
    .X(_1805_));
 sg13g2_nand2_1 _3694_ (.Y(_1806_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[12] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[12] ));
 sg13g2_xor2_1 _3695_ (.B(\u_ddc_top_level.cic_left_inst.int_reg2[12] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[12] ),
    .X(_1807_));
 sg13g2_nand2_1 _3696_ (.Y(_1808_),
    .A(_1805_),
    .B(_1807_));
 sg13g2_xor2_1 _3697_ (.B(_1807_),
    .A(_1805_),
    .X(_0034_));
 sg13g2_nor2_1 _3698_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[13] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[13] ),
    .Y(_1809_));
 sg13g2_xor2_1 _3699_ (.B(\u_ddc_top_level.cic_left_inst.int_reg2[13] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[13] ),
    .X(_1810_));
 sg13g2_and2_1 _3700_ (.A(_1806_),
    .B(_1808_),
    .X(_1811_));
 sg13g2_xnor2_1 _3701_ (.Y(_0035_),
    .A(_1810_),
    .B(_1811_));
 sg13g2_nand2_1 _3702_ (.Y(_1812_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[14] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[14] ));
 sg13g2_xor2_1 _3703_ (.B(\u_ddc_top_level.cic_left_inst.int_reg2[14] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[14] ),
    .X(_1813_));
 sg13g2_a22oi_1 _3704_ (.Y(_1814_),
    .B1(\u_ddc_top_level.cic_left_inst.int_reg2[13] ),
    .B2(\u_ddc_top_level.cic_left_inst.int_reg1[13] ),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg2[12] ),
    .A1(\u_ddc_top_level.cic_left_inst.int_reg1[12] ));
 sg13g2_a21oi_1 _3705_ (.A1(_1808_),
    .A2(_1814_),
    .Y(_1815_),
    .B1(_1809_));
 sg13g2_nand2_1 _3706_ (.Y(_1816_),
    .A(_1813_),
    .B(_1815_));
 sg13g2_xor2_1 _3707_ (.B(_1815_),
    .A(_1813_),
    .X(_0036_));
 sg13g2_nor2_1 _3708_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[15] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[15] ),
    .Y(_1817_));
 sg13g2_nand2_1 _3709_ (.Y(_1818_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[15] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[15] ));
 sg13g2_nor2b_1 _3710_ (.A(_1817_),
    .B_N(_1818_),
    .Y(_1819_));
 sg13g2_nand2_1 _3711_ (.Y(_1820_),
    .A(_1812_),
    .B(_1816_));
 sg13g2_xor2_1 _3712_ (.B(_1820_),
    .A(_1819_),
    .X(_0037_));
 sg13g2_and4_1 _3713_ (.A(_1807_),
    .B(_1810_),
    .C(_1813_),
    .D(_1819_),
    .X(_1821_));
 sg13g2_o21ai_1 _3714_ (.B1(_1818_),
    .Y(_1822_),
    .A1(_1812_),
    .A2(_1817_));
 sg13g2_nor2_1 _3715_ (.A(_1809_),
    .B(_1814_),
    .Y(_1823_));
 sg13g2_nand3_1 _3716_ (.B(_1819_),
    .C(_1823_),
    .A(_1813_),
    .Y(_1824_));
 sg13g2_nand2b_1 _3717_ (.Y(_1825_),
    .B(_1824_),
    .A_N(_1822_));
 sg13g2_a21oi_2 _3718_ (.B1(_1825_),
    .Y(_1826_),
    .A2(_1821_),
    .A1(_1805_));
 sg13g2_a21o_2 _3719_ (.A2(_1821_),
    .A1(_1805_),
    .B1(_1825_),
    .X(_1827_));
 sg13g2_nand2_1 _3720_ (.Y(_1828_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[16] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[16] ));
 sg13g2_xnor2_1 _3721_ (.Y(_1829_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[16] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[16] ));
 sg13g2_xnor2_1 _3722_ (.Y(_0038_),
    .A(_1827_),
    .B(_1829_));
 sg13g2_nor2_1 _3723_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[17] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[17] ),
    .Y(_1830_));
 sg13g2_nand2_1 _3724_ (.Y(_1831_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[17] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[17] ));
 sg13g2_nand2b_1 _3725_ (.Y(_1832_),
    .B(_1831_),
    .A_N(_1830_));
 sg13g2_o21ai_1 _3726_ (.B1(_1828_),
    .Y(_1833_),
    .A1(_1826_),
    .A2(_1829_));
 sg13g2_xnor2_1 _3727_ (.Y(_0039_),
    .A(_1832_),
    .B(_1833_));
 sg13g2_xor2_1 _3728_ (.B(\u_ddc_top_level.cic_left_inst.int_reg2[18] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[18] ),
    .X(_1834_));
 sg13g2_o21ai_1 _3729_ (.B1(_1831_),
    .Y(_1835_),
    .A1(_1828_),
    .A2(_1830_));
 sg13g2_nor2_1 _3730_ (.A(_1829_),
    .B(_1832_),
    .Y(_1836_));
 sg13g2_a21oi_1 _3731_ (.A1(_1827_),
    .A2(_1836_),
    .Y(_1837_),
    .B1(_1835_));
 sg13g2_nor2b_1 _3732_ (.A(_1837_),
    .B_N(_1834_),
    .Y(_1838_));
 sg13g2_xnor2_1 _3733_ (.Y(_0040_),
    .A(_1834_),
    .B(_1837_));
 sg13g2_or2_1 _3734_ (.X(_1839_),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[19] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[19] ));
 sg13g2_xor2_1 _3735_ (.B(\u_ddc_top_level.cic_left_inst.int_reg2[19] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[19] ),
    .X(_1840_));
 sg13g2_a21oi_1 _3736_ (.A1(\u_ddc_top_level.cic_left_inst.int_reg1[18] ),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg2[18] ),
    .Y(_1841_),
    .B1(_1838_));
 sg13g2_xnor2_1 _3737_ (.Y(_0041_),
    .A(_1840_),
    .B(_1841_));
 sg13g2_and2_1 _3738_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[20] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[20] ),
    .X(_1842_));
 sg13g2_or2_1 _3739_ (.X(_1843_),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[20] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[20] ));
 sg13g2_nand2b_1 _3740_ (.Y(_1844_),
    .B(_1843_),
    .A_N(_1842_));
 sg13g2_nand2_1 _3741_ (.Y(_1845_),
    .A(_1834_),
    .B(_1840_));
 sg13g2_inv_1 _3742_ (.Y(_1846_),
    .A(_1845_));
 sg13g2_and3_1 _3743_ (.X(_1847_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[18] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[18] ),
    .C(_1839_));
 sg13g2_a221oi_1 _3744_ (.B2(_1846_),
    .C1(_1847_),
    .B1(_1835_),
    .A1(\u_ddc_top_level.cic_left_inst.int_reg1[19] ),
    .Y(_1848_),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg2[19] ));
 sg13g2_nand2_1 _3745_ (.Y(_1849_),
    .A(_1836_),
    .B(_1846_));
 sg13g2_o21ai_1 _3746_ (.B1(_1848_),
    .Y(_1850_),
    .A1(_1826_),
    .A2(_1849_));
 sg13g2_xnor2_1 _3747_ (.Y(_0043_),
    .A(_1844_),
    .B(_1850_));
 sg13g2_nor2_1 _3748_ (.A(\u_ddc_top_level.cic_left_inst.int_reg1[21] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[21] ),
    .Y(_1851_));
 sg13g2_xor2_1 _3749_ (.B(\u_ddc_top_level.cic_left_inst.int_reg2[21] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[21] ),
    .X(_1852_));
 sg13g2_a21oi_1 _3750_ (.A1(_1843_),
    .A2(_1850_),
    .Y(_1853_),
    .B1(_1842_));
 sg13g2_xnor2_1 _3751_ (.Y(_0044_),
    .A(_1852_),
    .B(_1853_));
 sg13g2_nand2_1 _3752_ (.Y(_1854_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[22] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[22] ));
 sg13g2_xnor2_1 _3753_ (.Y(_1855_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[22] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[22] ));
 sg13g2_nor2b_1 _3754_ (.A(_1844_),
    .B_N(_1852_),
    .Y(_1856_));
 sg13g2_a21oi_1 _3755_ (.A1(\u_ddc_top_level.cic_left_inst.int_reg1[21] ),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg2[21] ),
    .Y(_1857_),
    .B1(_1842_));
 sg13g2_nor2_1 _3756_ (.A(_1851_),
    .B(_1857_),
    .Y(_1858_));
 sg13g2_a21oi_1 _3757_ (.A1(_1850_),
    .A2(_1856_),
    .Y(_1859_),
    .B1(_1858_));
 sg13g2_xor2_1 _3758_ (.B(_1859_),
    .A(_1855_),
    .X(_0045_));
 sg13g2_nor2_1 _3759_ (.A(net881),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[23] ),
    .Y(_1860_));
 sg13g2_xnor2_1 _3760_ (.Y(_1861_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[23] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[23] ));
 sg13g2_o21ai_1 _3761_ (.B1(_1854_),
    .Y(_1862_),
    .A1(_1855_),
    .A2(_1859_));
 sg13g2_xnor2_1 _3762_ (.Y(_0046_),
    .A(_1861_),
    .B(_1862_));
 sg13g2_nor2_1 _3763_ (.A(_1855_),
    .B(_1861_),
    .Y(_1863_));
 sg13g2_and2_1 _3764_ (.A(_1856_),
    .B(_1863_),
    .X(_1864_));
 sg13g2_inv_1 _3765_ (.Y(_1865_),
    .A(_1864_));
 sg13g2_nor2_1 _3766_ (.A(_1849_),
    .B(_1865_),
    .Y(_1866_));
 sg13g2_nor2_1 _3767_ (.A(_1854_),
    .B(_1860_),
    .Y(_1867_));
 sg13g2_a221oi_1 _3768_ (.B2(_1863_),
    .C1(_1867_),
    .B1(_1858_),
    .A1(\u_ddc_top_level.cic_left_inst.int_reg1[23] ),
    .Y(_1868_),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg2[23] ));
 sg13g2_o21ai_1 _3769_ (.B1(_1868_),
    .Y(_1869_),
    .A1(_1848_),
    .A2(_1865_));
 sg13g2_a21oi_2 _3770_ (.B1(_1869_),
    .Y(_1870_),
    .A2(_1866_),
    .A1(_1827_));
 sg13g2_xor2_1 _3771_ (.B(\u_ddc_top_level.cic_left_inst.int_reg2[24] ),
    .A(net881),
    .X(_1871_));
 sg13g2_nor2b_1 _3772_ (.A(_1870_),
    .B_N(_1871_),
    .Y(_1872_));
 sg13g2_xnor2_1 _3773_ (.Y(_0047_),
    .A(_1870_),
    .B(_1871_));
 sg13g2_xor2_1 _3774_ (.B(\u_ddc_top_level.cic_left_inst.int_reg2[25] ),
    .A(net881),
    .X(_1873_));
 sg13g2_a21oi_1 _3775_ (.A1(net881),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg2[24] ),
    .Y(_1874_),
    .B1(_1872_));
 sg13g2_xnor2_1 _3776_ (.Y(_0048_),
    .A(_1873_),
    .B(_1874_));
 sg13g2_nand2_1 _3777_ (.Y(_1875_),
    .A(_1871_),
    .B(_1873_));
 sg13g2_o21ai_1 _3778_ (.B1(net881),
    .Y(_1876_),
    .A1(\u_ddc_top_level.cic_left_inst.int_reg2[24] ),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg2[25] ));
 sg13g2_o21ai_1 _3779_ (.B1(_1876_),
    .Y(_1877_),
    .A1(_1870_),
    .A2(_1875_));
 sg13g2_and2_1 _3780_ (.A(net881),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[26] ),
    .X(_1878_));
 sg13g2_or2_1 _3781_ (.X(_1879_),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[26] ),
    .A(net881));
 sg13g2_nand2b_1 _3782_ (.Y(_1880_),
    .B(_1879_),
    .A_N(_1878_));
 sg13g2_xnor2_1 _3783_ (.Y(_0049_),
    .A(_1877_),
    .B(_1880_));
 sg13g2_a21oi_1 _3784_ (.A1(_1877_),
    .A2(_1879_),
    .Y(_1881_),
    .B1(_1878_));
 sg13g2_xor2_1 _3785_ (.B(\u_ddc_top_level.cic_left_inst.int_reg2[27] ),
    .A(net881),
    .X(_1882_));
 sg13g2_xnor2_1 _3786_ (.Y(_0050_),
    .A(_1881_),
    .B(_1882_));
 sg13g2_xor2_1 _3787_ (.B(\u_ddc_top_level.cic_left_inst.int_reg2[0] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg1[0] ),
    .X(_0031_));
 sg13g2_nand2_1 _3788_ (.Y(_1883_),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[0] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[0] ));
 sg13g2_xor2_1 _3789_ (.B(\u_ddc_top_level.dsm_left_inst.integrator1[0] ),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[0] ),
    .X(_1884_));
 sg13g2_xnor2_1 _3790_ (.Y(_0169_),
    .A(_0006_),
    .B(_1884_));
 sg13g2_or2_1 _3791_ (.X(_1885_),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[1] ),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[1] ));
 sg13g2_xnor2_1 _3792_ (.Y(_1886_),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[1] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[1] ));
 sg13g2_o21ai_1 _3793_ (.B1(\u_ddc_top_level.dsm_left_inst.in_dither ),
    .Y(_1887_),
    .A1(\u_ddc_top_level.dsm_left_inst.integrator2[0] ),
    .A2(\u_ddc_top_level.dsm_left_inst.integrator1[0] ));
 sg13g2_nand2_1 _3794_ (.Y(_1888_),
    .A(_1883_),
    .B(_1887_));
 sg13g2_nand3b_1 _3795_ (.B(_1887_),
    .C(_1883_),
    .Y(_1889_),
    .A_N(_1886_));
 sg13g2_xnor2_1 _3796_ (.Y(_0179_),
    .A(_1886_),
    .B(_1888_));
 sg13g2_nor2_1 _3797_ (.A(\u_ddc_top_level.dsm_left_inst.integrator2[2] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[2] ),
    .Y(_1890_));
 sg13g2_xnor2_1 _3798_ (.Y(_1891_),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[2] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[2] ));
 sg13g2_and3_1 _3799_ (.X(_1892_),
    .A(_1885_),
    .B(_1889_),
    .C(_1891_));
 sg13g2_a21oi_1 _3800_ (.A1(_1885_),
    .A2(_1889_),
    .Y(_1893_),
    .B1(_1891_));
 sg13g2_or2_1 _3801_ (.X(_0180_),
    .B(_1893_),
    .A(_1892_));
 sg13g2_nor2_1 _3802_ (.A(\u_ddc_top_level.dsm_left_inst.integrator2[3] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[3] ),
    .Y(_1894_));
 sg13g2_xor2_1 _3803_ (.B(\u_ddc_top_level.dsm_left_inst.integrator1[3] ),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[3] ),
    .X(_1895_));
 sg13g2_o21ai_1 _3804_ (.B1(_1895_),
    .Y(_1896_),
    .A1(_1890_),
    .A2(_1893_));
 sg13g2_or3_1 _3805_ (.A(_1890_),
    .B(_1893_),
    .C(_1895_),
    .X(_1897_));
 sg13g2_nand2_1 _3806_ (.Y(_0181_),
    .A(_1896_),
    .B(_1897_));
 sg13g2_xor2_1 _3807_ (.B(\u_ddc_top_level.dsm_left_inst.integrator1[4] ),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[4] ),
    .X(_1898_));
 sg13g2_nor2_1 _3808_ (.A(_1894_),
    .B(_1898_),
    .Y(_1899_));
 sg13g2_xnor2_1 _3809_ (.Y(_1900_),
    .A(_1894_),
    .B(_1898_));
 sg13g2_xnor2_1 _3810_ (.Y(_0182_),
    .A(_1896_),
    .B(_1900_));
 sg13g2_nand2b_1 _3811_ (.Y(_1901_),
    .B(_0182_),
    .A_N(_1899_));
 sg13g2_nor2_1 _3812_ (.A(\u_ddc_top_level.dsm_left_inst.integrator2[5] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[5] ),
    .Y(_1902_));
 sg13g2_xnor2_1 _3813_ (.Y(_1903_),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[5] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[5] ));
 sg13g2_nor3_1 _3814_ (.A(\u_ddc_top_level.dsm_left_inst.integrator2[4] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[4] ),
    .C(_1903_),
    .Y(_1904_));
 sg13g2_o21ai_1 _3815_ (.B1(_1903_),
    .Y(_1905_),
    .A1(\u_ddc_top_level.dsm_left_inst.integrator2[4] ),
    .A2(\u_ddc_top_level.dsm_left_inst.integrator1[4] ));
 sg13g2_nand2b_1 _3816_ (.Y(_1906_),
    .B(_1905_),
    .A_N(_1904_));
 sg13g2_xnor2_1 _3817_ (.Y(_0183_),
    .A(_1901_),
    .B(_1906_));
 sg13g2_nor2_1 _3818_ (.A(\u_ddc_top_level.dsm_left_inst.integrator2[6] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[6] ),
    .Y(_1907_));
 sg13g2_xnor2_1 _3819_ (.Y(_1908_),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[6] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[6] ));
 sg13g2_nand2b_1 _3820_ (.Y(_1909_),
    .B(_1908_),
    .A_N(_1902_));
 sg13g2_xor2_1 _3821_ (.B(_1908_),
    .A(_1902_),
    .X(_1910_));
 sg13g2_nor2b_1 _3822_ (.A(_1899_),
    .B_N(_1905_),
    .Y(_1911_));
 sg13g2_o21ai_1 _3823_ (.B1(_0183_),
    .Y(_1912_),
    .A1(_1904_),
    .A2(_1911_));
 sg13g2_xnor2_1 _3824_ (.Y(_0184_),
    .A(_1910_),
    .B(_1912_));
 sg13g2_nor2_1 _3825_ (.A(\u_ddc_top_level.dsm_left_inst.integrator2[7] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[7] ),
    .Y(_1913_));
 sg13g2_xor2_1 _3826_ (.B(\u_ddc_top_level.dsm_left_inst.integrator1[7] ),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[7] ),
    .X(_1914_));
 sg13g2_nand2_1 _3827_ (.Y(_1915_),
    .A(_1907_),
    .B(_1914_));
 sg13g2_xnor2_1 _3828_ (.Y(_1916_),
    .A(_1907_),
    .B(_1914_));
 sg13g2_nand2_1 _3829_ (.Y(_1917_),
    .A(_1909_),
    .B(_0184_));
 sg13g2_xnor2_1 _3830_ (.Y(_0185_),
    .A(_1916_),
    .B(_1917_));
 sg13g2_nor4_1 _3831_ (.A(_1900_),
    .B(_1906_),
    .C(_1910_),
    .D(_1916_),
    .Y(_1918_));
 sg13g2_o21ai_1 _3832_ (.B1(_1909_),
    .Y(_1919_),
    .A1(_1907_),
    .A2(_1914_));
 sg13g2_nor4_1 _3833_ (.A(_1904_),
    .B(_1910_),
    .C(_1911_),
    .D(_1916_),
    .Y(_1920_));
 sg13g2_a221oi_1 _3834_ (.B2(_1915_),
    .C1(_1920_),
    .B1(_1919_),
    .A1(_1896_),
    .Y(_1921_),
    .A2(_1918_));
 sg13g2_xnor2_1 _3835_ (.Y(_1922_),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[8] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[8] ));
 sg13g2_nor2b_1 _3836_ (.A(_1913_),
    .B_N(_1922_),
    .Y(_1923_));
 sg13g2_xor2_1 _3837_ (.B(_1922_),
    .A(_1913_),
    .X(_1924_));
 sg13g2_xor2_1 _3838_ (.B(_1924_),
    .A(_1921_),
    .X(_0186_));
 sg13g2_nor2_1 _3839_ (.A(\u_ddc_top_level.dsm_left_inst.integrator2[9] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[9] ),
    .Y(_1925_));
 sg13g2_xnor2_1 _3840_ (.Y(_1926_),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[9] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[9] ));
 sg13g2_or3_1 _3841_ (.A(\u_ddc_top_level.dsm_left_inst.integrator2[8] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[8] ),
    .C(_1926_),
    .X(_1927_));
 sg13g2_o21ai_1 _3842_ (.B1(_1926_),
    .Y(_1928_),
    .A1(\u_ddc_top_level.dsm_left_inst.integrator2[8] ),
    .A2(\u_ddc_top_level.dsm_left_inst.integrator1[8] ));
 sg13g2_nand2_1 _3843_ (.Y(_1929_),
    .A(_1927_),
    .B(_1928_));
 sg13g2_nand2b_1 _3844_ (.Y(_1930_),
    .B(_0186_),
    .A_N(_1923_));
 sg13g2_xnor2_1 _3845_ (.Y(_0187_),
    .A(_1929_),
    .B(_1930_));
 sg13g2_xnor2_1 _3846_ (.Y(_1931_),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[10] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[10] ));
 sg13g2_nand2b_1 _3847_ (.Y(_1932_),
    .B(_1931_),
    .A_N(_1925_));
 sg13g2_xor2_1 _3848_ (.B(_1931_),
    .A(_1925_),
    .X(_1933_));
 sg13g2_nand2_1 _3849_ (.Y(_1934_),
    .A(_1923_),
    .B(_1927_));
 sg13g2_nand2_1 _3850_ (.Y(_1935_),
    .A(_1928_),
    .B(_1934_));
 sg13g2_nand3_1 _3851_ (.B(_0187_),
    .C(_1934_),
    .A(_1928_),
    .Y(_1936_));
 sg13g2_xnor2_1 _3852_ (.Y(_0170_),
    .A(_1933_),
    .B(_1936_));
 sg13g2_nor2_1 _3853_ (.A(\u_ddc_top_level.dsm_left_inst.integrator2[11] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[11] ),
    .Y(_1937_));
 sg13g2_xnor2_1 _3854_ (.Y(_1938_),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[11] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[11] ));
 sg13g2_o21ai_1 _3855_ (.B1(_1938_),
    .Y(_1939_),
    .A1(\u_ddc_top_level.dsm_left_inst.integrator2[10] ),
    .A2(\u_ddc_top_level.dsm_left_inst.integrator1[10] ));
 sg13g2_or3_1 _3856_ (.A(\u_ddc_top_level.dsm_left_inst.integrator2[10] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[10] ),
    .C(_1938_),
    .X(_1940_));
 sg13g2_nand2_1 _3857_ (.Y(_1941_),
    .A(_1939_),
    .B(_1940_));
 sg13g2_nand2_1 _3858_ (.Y(_1942_),
    .A(_1932_),
    .B(_0170_));
 sg13g2_xnor2_1 _3859_ (.Y(_0171_),
    .A(_1941_),
    .B(_1942_));
 sg13g2_nor2_1 _3860_ (.A(_1933_),
    .B(_1941_),
    .Y(_1943_));
 sg13g2_or4_1 _3861_ (.A(_1924_),
    .B(_1929_),
    .C(_1933_),
    .D(_1941_),
    .X(_1944_));
 sg13g2_nand2_1 _3862_ (.Y(_1945_),
    .A(_1932_),
    .B(_1939_));
 sg13g2_a22oi_1 _3863_ (.Y(_1946_),
    .B1(_1945_),
    .B2(_1940_),
    .A2(_1943_),
    .A1(_1935_));
 sg13g2_o21ai_1 _3864_ (.B1(_1946_),
    .Y(_1947_),
    .A1(_1921_),
    .A2(_1944_));
 sg13g2_nor2_1 _3865_ (.A(\u_ddc_top_level.dsm_left_inst.integrator2[12] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[12] ),
    .Y(_1948_));
 sg13g2_xnor2_1 _3866_ (.Y(_1949_),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[12] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[12] ));
 sg13g2_nor2b_1 _3867_ (.A(_1937_),
    .B_N(_1949_),
    .Y(_1950_));
 sg13g2_xor2_1 _3868_ (.B(_1949_),
    .A(_1937_),
    .X(_1951_));
 sg13g2_xnor2_1 _3869_ (.Y(_0172_),
    .A(_1947_),
    .B(_1951_));
 sg13g2_nand2b_1 _3870_ (.Y(_1952_),
    .B(_0172_),
    .A_N(_1950_));
 sg13g2_nor2_1 _3871_ (.A(\u_ddc_top_level.dsm_left_inst.integrator2[13] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[13] ),
    .Y(_1953_));
 sg13g2_xor2_1 _3872_ (.B(\u_ddc_top_level.dsm_left_inst.integrator1[13] ),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[13] ),
    .X(_1954_));
 sg13g2_nand2_1 _3873_ (.Y(_1955_),
    .A(_1948_),
    .B(_1954_));
 sg13g2_nor2_1 _3874_ (.A(_1948_),
    .B(_1954_),
    .Y(_1956_));
 sg13g2_xnor2_1 _3875_ (.Y(_1957_),
    .A(_1948_),
    .B(_1954_));
 sg13g2_xnor2_1 _3876_ (.Y(_0173_),
    .A(_1952_),
    .B(_1957_));
 sg13g2_nor2_1 _3877_ (.A(\u_ddc_top_level.dsm_left_inst.integrator2[14] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[14] ),
    .Y(_1958_));
 sg13g2_xnor2_1 _3878_ (.Y(_1959_),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[14] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[14] ));
 sg13g2_nor2b_1 _3879_ (.A(_1953_),
    .B_N(_1959_),
    .Y(_1960_));
 sg13g2_nor3_1 _3880_ (.A(\u_ddc_top_level.dsm_left_inst.integrator2[13] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[13] ),
    .C(_1959_),
    .Y(_1961_));
 sg13g2_nor2_1 _3881_ (.A(_1960_),
    .B(_1961_),
    .Y(_1962_));
 sg13g2_nor2_1 _3882_ (.A(_1951_),
    .B(_1957_),
    .Y(_1963_));
 sg13g2_o21ai_1 _3883_ (.B1(_1955_),
    .Y(_1964_),
    .A1(_1950_),
    .A2(_1956_));
 sg13g2_inv_1 _3884_ (.Y(_1965_),
    .A(_1964_));
 sg13g2_a21oi_1 _3885_ (.A1(_1947_),
    .A2(_1963_),
    .Y(_1966_),
    .B1(_1965_));
 sg13g2_xnor2_1 _3886_ (.Y(_0174_),
    .A(_1962_),
    .B(_1966_));
 sg13g2_nor2_1 _3887_ (.A(\u_ddc_top_level.dsm_left_inst.integrator2[15] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[15] ),
    .Y(_1967_));
 sg13g2_xor2_1 _3888_ (.B(\u_ddc_top_level.dsm_left_inst.integrator1[15] ),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[15] ),
    .X(_1968_));
 sg13g2_nand2_1 _3889_ (.Y(_1969_),
    .A(_1958_),
    .B(_1968_));
 sg13g2_or2_1 _3890_ (.X(_1970_),
    .B(_1968_),
    .A(_1958_));
 sg13g2_nand2_1 _3891_ (.Y(_1971_),
    .A(_1969_),
    .B(_1970_));
 sg13g2_nand2b_1 _3892_ (.Y(_1972_),
    .B(_0174_),
    .A_N(_1960_));
 sg13g2_xnor2_1 _3893_ (.Y(_0175_),
    .A(_1971_),
    .B(_1972_));
 sg13g2_nor2_1 _3894_ (.A(\u_ddc_top_level.dsm_left_inst.integrator2[16] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[16] ),
    .Y(_1973_));
 sg13g2_xor2_1 _3895_ (.B(\u_ddc_top_level.dsm_left_inst.integrator1[16] ),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[16] ),
    .X(_1974_));
 sg13g2_nor2_1 _3896_ (.A(_1967_),
    .B(_1974_),
    .Y(_1975_));
 sg13g2_xnor2_1 _3897_ (.Y(_1976_),
    .A(_1967_),
    .B(_1974_));
 sg13g2_nand2_1 _3898_ (.Y(_1977_),
    .A(_1960_),
    .B(_1969_));
 sg13g2_nand3_1 _3899_ (.B(_1970_),
    .C(_1977_),
    .A(_1964_),
    .Y(_1978_));
 sg13g2_a21o_1 _3900_ (.A2(_1963_),
    .A1(_1947_),
    .B1(_1978_),
    .X(_1979_));
 sg13g2_o21ai_1 _3901_ (.B1(_1968_),
    .Y(_1980_),
    .A1(_1958_),
    .A2(_1961_));
 sg13g2_a21o_1 _3902_ (.A2(_1980_),
    .A1(_1979_),
    .B1(_1976_),
    .X(_1981_));
 sg13g2_nand3_1 _3903_ (.B(_1979_),
    .C(_1980_),
    .A(_1976_),
    .Y(_1982_));
 sg13g2_nand2_1 _3904_ (.Y(_0176_),
    .A(_1981_),
    .B(_1982_));
 sg13g2_a21oi_1 _3905_ (.A1(_1981_),
    .A2(_1982_),
    .Y(_1983_),
    .B1(_1975_));
 sg13g2_nand2_1 _3906_ (.Y(_1984_),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[17] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[17] ));
 sg13g2_xor2_1 _3907_ (.B(\u_ddc_top_level.dsm_left_inst.integrator1[17] ),
    .A(\u_ddc_top_level.dsm_left_inst.integrator2[17] ),
    .X(_1985_));
 sg13g2_xnor2_1 _3908_ (.Y(_1986_),
    .A(_1973_),
    .B(_1985_));
 sg13g2_xnor2_1 _3909_ (.Y(_0177_),
    .A(_1983_),
    .B(_1986_));
 sg13g2_nand2b_1 _3910_ (.Y(_1987_),
    .B(_0177_),
    .A_N(_1985_));
 sg13g2_xnor2_1 _3911_ (.Y(_1988_),
    .A(\u_ddc_top_level.dsm_left_inst.integrator1[18] ),
    .B(_1984_));
 sg13g2_xnor2_1 _3912_ (.Y(_0178_),
    .A(_1987_),
    .B(_1988_));
 sg13g2_nand2_1 _3913_ (.Y(_1989_),
    .A(\u_ddc_top_level.cic_out_right[0] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[0] ));
 sg13g2_xor2_1 _3914_ (.B(\u_ddc_top_level.dsm_right_inst.integrator1[0] ),
    .A(\u_ddc_top_level.cic_out_right[0] ),
    .X(_0150_));
 sg13g2_nor2_1 _3915_ (.A(\u_ddc_top_level.cic_out_right[1] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[1] ),
    .Y(_1990_));
 sg13g2_xor2_1 _3916_ (.B(\u_ddc_top_level.dsm_right_inst.integrator1[1] ),
    .A(\u_ddc_top_level.cic_out_right[1] ),
    .X(_1991_));
 sg13g2_xnor2_1 _3917_ (.Y(_0160_),
    .A(_1989_),
    .B(_1991_));
 sg13g2_or2_1 _3918_ (.X(_1992_),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[2] ),
    .A(\u_ddc_top_level.cic_out_right[2] ));
 sg13g2_nand2_1 _3919_ (.Y(_1993_),
    .A(\u_ddc_top_level.cic_out_right[2] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[2] ));
 sg13g2_nand2_1 _3920_ (.Y(_1994_),
    .A(_1992_),
    .B(_1993_));
 sg13g2_a22oi_1 _3921_ (.Y(_1995_),
    .B1(\u_ddc_top_level.dsm_right_inst.integrator1[1] ),
    .B2(\u_ddc_top_level.cic_out_right[1] ),
    .A2(\u_ddc_top_level.dsm_right_inst.integrator1[0] ),
    .A1(\u_ddc_top_level.cic_out_right[0] ));
 sg13g2_nor2_1 _3922_ (.A(_1990_),
    .B(_1995_),
    .Y(_1996_));
 sg13g2_xnor2_1 _3923_ (.Y(_0161_),
    .A(_1994_),
    .B(_1996_));
 sg13g2_nor2_1 _3924_ (.A(\u_ddc_top_level.cic_out_right[3] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[3] ),
    .Y(_1997_));
 sg13g2_xnor2_1 _3925_ (.Y(_1998_),
    .A(\u_ddc_top_level.cic_out_right[3] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[3] ));
 sg13g2_o21ai_1 _3926_ (.B1(_1993_),
    .Y(_1999_),
    .A1(_1990_),
    .A2(_1995_));
 sg13g2_and3_1 _3927_ (.X(_2000_),
    .A(_1992_),
    .B(_1998_),
    .C(_1999_));
 sg13g2_a21oi_2 _3928_ (.B1(_1998_),
    .Y(_2001_),
    .A2(_1999_),
    .A1(_1992_));
 sg13g2_or2_1 _3929_ (.X(_0162_),
    .B(_2001_),
    .A(_2000_));
 sg13g2_nor2_1 _3930_ (.A(\u_ddc_top_level.cic_out_right[4] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[4] ),
    .Y(_2002_));
 sg13g2_xnor2_1 _3931_ (.Y(_2003_),
    .A(\u_ddc_top_level.cic_out_right[4] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[4] ));
 sg13g2_nor2b_1 _3932_ (.A(_1997_),
    .B_N(_2003_),
    .Y(_2004_));
 sg13g2_nand2b_1 _3933_ (.Y(_2005_),
    .B(_2003_),
    .A_N(_1997_));
 sg13g2_nor3_1 _3934_ (.A(\u_ddc_top_level.cic_out_right[3] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[3] ),
    .C(_2003_),
    .Y(_2006_));
 sg13g2_nor2_1 _3935_ (.A(_2001_),
    .B(_2006_),
    .Y(_2007_));
 sg13g2_a22oi_1 _3936_ (.Y(_0163_),
    .B1(_2005_),
    .B2(_2007_),
    .A2(_2003_),
    .A1(_2001_));
 sg13g2_nor2_1 _3937_ (.A(\u_ddc_top_level.cic_out_right[5] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[5] ),
    .Y(_2008_));
 sg13g2_xnor2_1 _3938_ (.Y(_2009_),
    .A(\u_ddc_top_level.cic_out_right[5] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[5] ));
 sg13g2_nor3_1 _3939_ (.A(\u_ddc_top_level.cic_out_right[4] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[4] ),
    .C(_2009_),
    .Y(_2010_));
 sg13g2_nand2b_1 _3940_ (.Y(_2011_),
    .B(_2009_),
    .A_N(_2002_));
 sg13g2_xor2_1 _3941_ (.B(_2009_),
    .A(_2002_),
    .X(_2012_));
 sg13g2_nand2_1 _3942_ (.Y(_2013_),
    .A(_2005_),
    .B(_0163_));
 sg13g2_xnor2_1 _3943_ (.Y(_0164_),
    .A(_2012_),
    .B(_2013_));
 sg13g2_nor2_1 _3944_ (.A(\u_ddc_top_level.cic_out_right[6] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[6] ),
    .Y(_2014_));
 sg13g2_xnor2_1 _3945_ (.Y(_2015_),
    .A(\u_ddc_top_level.cic_out_right[6] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[6] ));
 sg13g2_nand2b_1 _3946_ (.Y(_2016_),
    .B(_2015_),
    .A_N(_2008_));
 sg13g2_xor2_1 _3947_ (.B(_2015_),
    .A(_2008_),
    .X(_2017_));
 sg13g2_nand2b_1 _3948_ (.Y(_2018_),
    .B(_2004_),
    .A_N(_2010_));
 sg13g2_o21ai_1 _3949_ (.B1(_2011_),
    .Y(_2019_),
    .A1(_2005_),
    .A2(_2010_));
 sg13g2_nand3_1 _3950_ (.B(_0164_),
    .C(_2018_),
    .A(_2011_),
    .Y(_2020_));
 sg13g2_xnor2_1 _3951_ (.Y(_0165_),
    .A(_2017_),
    .B(_2020_));
 sg13g2_nor2_1 _3952_ (.A(\u_ddc_top_level.cic_out_right[7] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[7] ),
    .Y(_2021_));
 sg13g2_xor2_1 _3953_ (.B(\u_ddc_top_level.dsm_right_inst.integrator1[7] ),
    .A(\u_ddc_top_level.cic_out_right[7] ),
    .X(_2022_));
 sg13g2_nand2_1 _3954_ (.Y(_2023_),
    .A(_2014_),
    .B(_2022_));
 sg13g2_xnor2_1 _3955_ (.Y(_2024_),
    .A(_2014_),
    .B(_2022_));
 sg13g2_nand2_1 _3956_ (.Y(_2025_),
    .A(_2016_),
    .B(_0165_));
 sg13g2_xnor2_1 _3957_ (.Y(_0166_),
    .A(_2024_),
    .B(_2025_));
 sg13g2_nor2_1 _3958_ (.A(_2017_),
    .B(_2024_),
    .Y(_2026_));
 sg13g2_or3_1 _3959_ (.A(_2012_),
    .B(_2017_),
    .C(_2024_),
    .X(_2027_));
 sg13g2_nor4_1 _3960_ (.A(_2001_),
    .B(_2004_),
    .C(_2006_),
    .D(_2027_),
    .Y(_2028_));
 sg13g2_o21ai_1 _3961_ (.B1(_2016_),
    .Y(_2029_),
    .A1(_2014_),
    .A2(_2022_));
 sg13g2_a22oi_1 _3962_ (.Y(_2030_),
    .B1(_2029_),
    .B2(_2023_),
    .A2(_2026_),
    .A1(_2019_));
 sg13g2_nand2b_1 _3963_ (.Y(_2031_),
    .B(_2030_),
    .A_N(_2028_));
 sg13g2_nor2_1 _3964_ (.A(\u_ddc_top_level.cic_out_right[8] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[8] ),
    .Y(_2032_));
 sg13g2_xnor2_1 _3965_ (.Y(_2033_),
    .A(\u_ddc_top_level.cic_out_right[8] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[8] ));
 sg13g2_nor2b_1 _3966_ (.A(_2021_),
    .B_N(_2033_),
    .Y(_2034_));
 sg13g2_xor2_1 _3967_ (.B(_2033_),
    .A(_2021_),
    .X(_2035_));
 sg13g2_xnor2_1 _3968_ (.Y(_0167_),
    .A(_2031_),
    .B(_2035_));
 sg13g2_nand2b_1 _3969_ (.Y(_2036_),
    .B(_0167_),
    .A_N(_2034_));
 sg13g2_nor2_1 _3970_ (.A(\u_ddc_top_level.cic_out_right[9] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[9] ),
    .Y(_2037_));
 sg13g2_xor2_1 _3971_ (.B(\u_ddc_top_level.dsm_right_inst.integrator1[9] ),
    .A(\u_ddc_top_level.cic_out_right[9] ),
    .X(_2038_));
 sg13g2_nand2_1 _3972_ (.Y(_2039_),
    .A(_2032_),
    .B(_2038_));
 sg13g2_nor2_1 _3973_ (.A(_2032_),
    .B(_2038_),
    .Y(_2040_));
 sg13g2_xnor2_1 _3974_ (.Y(_2041_),
    .A(_2032_),
    .B(_2038_));
 sg13g2_xnor2_1 _3975_ (.Y(_0168_),
    .A(_2036_),
    .B(_2041_));
 sg13g2_xnor2_1 _3976_ (.Y(_2042_),
    .A(\u_ddc_top_level.cic_out_right[10] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[10] ));
 sg13g2_nand2b_1 _3977_ (.Y(_2043_),
    .B(_2042_),
    .A_N(_2037_));
 sg13g2_xor2_1 _3978_ (.B(_2042_),
    .A(_2037_),
    .X(_2044_));
 sg13g2_o21ai_1 _3979_ (.B1(_2039_),
    .Y(_2045_),
    .A1(_2034_),
    .A2(_2040_));
 sg13g2_nand2_1 _3980_ (.Y(_2046_),
    .A(_0168_),
    .B(_2045_));
 sg13g2_xnor2_1 _3981_ (.Y(_0151_),
    .A(_2044_),
    .B(_2046_));
 sg13g2_nor2_1 _3982_ (.A(\u_ddc_top_level.cic_out_right[11] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[11] ),
    .Y(_2047_));
 sg13g2_xnor2_1 _3983_ (.Y(_2048_),
    .A(\u_ddc_top_level.cic_out_right[11] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[11] ));
 sg13g2_o21ai_1 _3984_ (.B1(_2048_),
    .Y(_2049_),
    .A1(\u_ddc_top_level.cic_out_right[10] ),
    .A2(\u_ddc_top_level.dsm_right_inst.integrator1[10] ));
 sg13g2_or3_1 _3985_ (.A(\u_ddc_top_level.cic_out_right[10] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[10] ),
    .C(_2048_),
    .X(_2050_));
 sg13g2_nand2_1 _3986_ (.Y(_2051_),
    .A(_2049_),
    .B(_2050_));
 sg13g2_nand2_1 _3987_ (.Y(_2052_),
    .A(_2043_),
    .B(_0151_));
 sg13g2_xnor2_1 _3988_ (.Y(_0152_),
    .A(_2051_),
    .B(_2052_));
 sg13g2_xor2_1 _3989_ (.B(\u_ddc_top_level.dsm_right_inst.integrator1[12] ),
    .A(\u_ddc_top_level.cic_out_right[12] ),
    .X(_2053_));
 sg13g2_nor2_1 _3990_ (.A(_2047_),
    .B(_2053_),
    .Y(_2054_));
 sg13g2_xnor2_1 _3991_ (.Y(_2055_),
    .A(_2047_),
    .B(_2053_));
 sg13g2_nor3_1 _3992_ (.A(_2044_),
    .B(_2045_),
    .C(_2051_),
    .Y(_2056_));
 sg13g2_nor4_1 _3993_ (.A(_2035_),
    .B(_2041_),
    .C(_2044_),
    .D(_2051_),
    .Y(_2057_));
 sg13g2_nand2_1 _3994_ (.Y(_2058_),
    .A(_2043_),
    .B(_2049_));
 sg13g2_a221oi_1 _3995_ (.B2(_2050_),
    .C1(_2056_),
    .B1(_2058_),
    .A1(_2031_),
    .Y(_2059_),
    .A2(_2057_));
 sg13g2_xor2_1 _3996_ (.B(_2059_),
    .A(_2055_),
    .X(_0153_));
 sg13g2_nand2b_1 _3997_ (.Y(_2060_),
    .B(_0153_),
    .A_N(_2054_));
 sg13g2_nor2_1 _3998_ (.A(\u_ddc_top_level.cic_out_right[13] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[13] ),
    .Y(_2061_));
 sg13g2_xnor2_1 _3999_ (.Y(_2062_),
    .A(\u_ddc_top_level.cic_out_right[13] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[13] ));
 sg13g2_or3_1 _4000_ (.A(\u_ddc_top_level.cic_out_right[12] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[12] ),
    .C(_2062_),
    .X(_2063_));
 sg13g2_o21ai_1 _4001_ (.B1(_2062_),
    .Y(_2064_),
    .A1(\u_ddc_top_level.cic_out_right[12] ),
    .A2(\u_ddc_top_level.dsm_right_inst.integrator1[12] ));
 sg13g2_nand2_1 _4002_ (.Y(_2065_),
    .A(_2063_),
    .B(_2064_));
 sg13g2_xnor2_1 _4003_ (.Y(_0154_),
    .A(_2060_),
    .B(_2065_));
 sg13g2_nor2_1 _4004_ (.A(\u_ddc_top_level.cic_out_right[14] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[14] ),
    .Y(_2066_));
 sg13g2_xnor2_1 _4005_ (.Y(_2067_),
    .A(\u_ddc_top_level.cic_out_right[14] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[14] ));
 sg13g2_nor2b_1 _4006_ (.A(_2061_),
    .B_N(_2067_),
    .Y(_2068_));
 sg13g2_xnor2_1 _4007_ (.Y(_2069_),
    .A(_2061_),
    .B(_2067_));
 sg13g2_nor3_1 _4008_ (.A(_2055_),
    .B(_2059_),
    .C(_2065_),
    .Y(_2070_));
 sg13g2_nand2_1 _4009_ (.Y(_2071_),
    .A(_2054_),
    .B(_2063_));
 sg13g2_nand2_1 _4010_ (.Y(_2072_),
    .A(_2064_),
    .B(_2071_));
 sg13g2_nor2_1 _4011_ (.A(_2070_),
    .B(_2072_),
    .Y(_2073_));
 sg13g2_o21ai_1 _4012_ (.B1(_2069_),
    .Y(_2074_),
    .A1(_2070_),
    .A2(_2072_));
 sg13g2_xnor2_1 _4013_ (.Y(_0155_),
    .A(_2069_),
    .B(_2073_));
 sg13g2_or2_1 _4014_ (.X(_2075_),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[15] ),
    .A(\u_ddc_top_level.cic_out_right[15] ));
 sg13g2_nand2_1 _4015_ (.Y(_2076_),
    .A(\u_ddc_top_level.cic_out_right[15] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[15] ));
 sg13g2_nand3_1 _4016_ (.B(_2075_),
    .C(_2076_),
    .A(_2066_),
    .Y(_2077_));
 sg13g2_a21oi_1 _4017_ (.A1(_2075_),
    .A2(_2076_),
    .Y(_2078_),
    .B1(_2066_));
 sg13g2_a21o_1 _4018_ (.A2(_2076_),
    .A1(_2075_),
    .B1(_2066_),
    .X(_2079_));
 sg13g2_nand2_1 _4019_ (.Y(_2080_),
    .A(_2077_),
    .B(_2079_));
 sg13g2_nand2b_1 _4020_ (.Y(_2081_),
    .B(_0155_),
    .A_N(_2068_));
 sg13g2_xnor2_1 _4021_ (.Y(_0156_),
    .A(_2080_),
    .B(_2081_));
 sg13g2_nand2_1 _4022_ (.Y(_2082_),
    .A(\u_ddc_top_level.cic_out_right[15] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator1[16] ));
 sg13g2_a21oi_1 _4023_ (.A1(\u_ddc_top_level.dsm_right_inst.integrator1[15] ),
    .A2(\u_ddc_top_level.dsm_right_inst.integrator1[16] ),
    .Y(_2083_),
    .B1(\u_ddc_top_level.cic_out_right[15] ));
 sg13g2_nand2b_1 _4024_ (.Y(_2084_),
    .B(_2082_),
    .A_N(_2083_));
 sg13g2_o21ai_1 _4025_ (.B1(_2084_),
    .Y(_2085_),
    .A1(\u_ddc_top_level.dsm_right_inst.integrator1[16] ),
    .A2(_2075_));
 sg13g2_o21ai_1 _4026_ (.B1(_2077_),
    .Y(_2086_),
    .A1(_2068_),
    .A2(_2078_));
 sg13g2_o21ai_1 _4027_ (.B1(_2086_),
    .Y(_2087_),
    .A1(_2074_),
    .A2(_2080_));
 sg13g2_nand2b_1 _4028_ (.Y(_2088_),
    .B(_2087_),
    .A_N(_2085_));
 sg13g2_xnor2_1 _4029_ (.Y(_0157_),
    .A(_2085_),
    .B(_2087_));
 sg13g2_nand2_1 _4030_ (.Y(_2089_),
    .A(_2084_),
    .B(_0157_));
 sg13g2_nand2b_1 _4031_ (.Y(_2090_),
    .B(\u_ddc_top_level.cic_out_right[15] ),
    .A_N(\u_ddc_top_level.dsm_right_inst.feedback[17] ));
 sg13g2_nor2b_1 _4032_ (.A(\u_ddc_top_level.cic_out_right[15] ),
    .B_N(\u_ddc_top_level.dsm_right_inst.feedback[17] ),
    .Y(_2091_));
 sg13g2_xnor2_1 _4033_ (.Y(_2092_),
    .A(\u_ddc_top_level.dsm_right_inst.feedback[17] ),
    .B(\u_ddc_top_level.cic_out_right[15] ));
 sg13g2_xnor2_1 _4034_ (.Y(_2093_),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[17] ),
    .B(_2092_));
 sg13g2_xnor2_1 _4035_ (.Y(_2094_),
    .A(_2082_),
    .B(_2093_));
 sg13g2_xnor2_1 _4036_ (.Y(_0158_),
    .A(_2089_),
    .B(_2094_));
 sg13g2_or2_1 _4037_ (.X(_2095_),
    .B(_2093_),
    .A(_2083_));
 sg13g2_o21ai_1 _4038_ (.B1(_2095_),
    .Y(_2096_),
    .A1(_2088_),
    .A2(_2094_));
 sg13g2_o21ai_1 _4039_ (.B1(_2090_),
    .Y(_2097_),
    .A1(\u_ddc_top_level.dsm_right_inst.integrator1[17] ),
    .A2(_2091_));
 sg13g2_xnor2_1 _4040_ (.Y(_2098_),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[18] ),
    .B(_2097_));
 sg13g2_xnor2_1 _4041_ (.Y(_0159_),
    .A(_2096_),
    .B(_2098_));
 sg13g2_nand2_1 _4042_ (.Y(_2099_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg2[12] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[0] ));
 sg13g2_xor2_1 _4043_ (.B(\u_ddc_top_level.dsm_left_inst.integrator1[0] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg2[12] ),
    .X(_0131_));
 sg13g2_nor2_1 _4044_ (.A(\u_ddc_top_level.cic_left_inst.int_reg2[13] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[1] ),
    .Y(_2100_));
 sg13g2_xor2_1 _4045_ (.B(\u_ddc_top_level.dsm_left_inst.integrator1[1] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg2[13] ),
    .X(_2101_));
 sg13g2_xnor2_1 _4046_ (.Y(_0141_),
    .A(_2099_),
    .B(_2101_));
 sg13g2_nor2_1 _4047_ (.A(\u_ddc_top_level.cic_left_inst.int_reg2[14] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[2] ),
    .Y(_2102_));
 sg13g2_and2_1 _4048_ (.A(\u_ddc_top_level.cic_left_inst.int_reg2[14] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[2] ),
    .X(_2103_));
 sg13g2_or2_1 _4049_ (.X(_2104_),
    .B(_2103_),
    .A(_2102_));
 sg13g2_a22oi_1 _4050_ (.Y(_2105_),
    .B1(\u_ddc_top_level.dsm_left_inst.integrator1[1] ),
    .B2(\u_ddc_top_level.cic_left_inst.int_reg2[13] ),
    .A2(\u_ddc_top_level.dsm_left_inst.integrator1[0] ),
    .A1(\u_ddc_top_level.cic_left_inst.int_reg2[12] ));
 sg13g2_nor2_1 _4051_ (.A(_2100_),
    .B(_2105_),
    .Y(_2106_));
 sg13g2_xnor2_1 _4052_ (.Y(_0142_),
    .A(_2104_),
    .B(_2106_));
 sg13g2_nor2_1 _4053_ (.A(\u_ddc_top_level.cic_left_inst.int_reg2[15] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[3] ),
    .Y(_2107_));
 sg13g2_xnor2_1 _4054_ (.Y(_2108_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg2[15] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[3] ));
 sg13g2_nor3_2 _4055_ (.A(_2100_),
    .B(_2102_),
    .C(_2105_),
    .Y(_2109_));
 sg13g2_nor3_2 _4056_ (.A(_2103_),
    .B(_2108_),
    .C(_2109_),
    .Y(_2110_));
 sg13g2_o21ai_1 _4057_ (.B1(_2108_),
    .Y(_2111_),
    .A1(_2103_),
    .A2(_2109_));
 sg13g2_nand2b_1 _4058_ (.Y(_0143_),
    .B(_2111_),
    .A_N(_2110_));
 sg13g2_xnor2_1 _4059_ (.Y(_2112_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg2[16] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[4] ));
 sg13g2_nand2b_1 _4060_ (.Y(_2113_),
    .B(_2112_),
    .A_N(_2107_));
 sg13g2_xor2_1 _4061_ (.B(_2112_),
    .A(_2107_),
    .X(_2114_));
 sg13g2_nor2_1 _4062_ (.A(_2110_),
    .B(_2114_),
    .Y(_2115_));
 sg13g2_a21oi_1 _4063_ (.A1(_2110_),
    .A2(_2112_),
    .Y(_0144_),
    .B1(_2115_));
 sg13g2_nor2_1 _4064_ (.A(\u_ddc_top_level.cic_left_inst.int_reg2[17] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[5] ),
    .Y(_2116_));
 sg13g2_xnor2_1 _4065_ (.Y(_2117_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg2[17] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[5] ));
 sg13g2_nor3_1 _4066_ (.A(\u_ddc_top_level.cic_left_inst.int_reg2[16] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[4] ),
    .C(_2117_),
    .Y(_2118_));
 sg13g2_o21ai_1 _4067_ (.B1(_2117_),
    .Y(_2119_),
    .A1(\u_ddc_top_level.cic_left_inst.int_reg2[16] ),
    .A2(\u_ddc_top_level.dsm_left_inst.integrator1[4] ));
 sg13g2_nand2b_1 _4068_ (.Y(_2120_),
    .B(_2119_),
    .A_N(_2118_));
 sg13g2_nand2_1 _4069_ (.Y(_2121_),
    .A(_2113_),
    .B(_0144_));
 sg13g2_xnor2_1 _4070_ (.Y(_0145_),
    .A(_2120_),
    .B(_2121_));
 sg13g2_nor2_1 _4071_ (.A(\u_ddc_top_level.cic_left_inst.int_reg2[18] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[6] ),
    .Y(_2122_));
 sg13g2_xnor2_1 _4072_ (.Y(_2123_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg2[18] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[6] ));
 sg13g2_nand2b_1 _4073_ (.Y(_2124_),
    .B(_2123_),
    .A_N(_2116_));
 sg13g2_xor2_1 _4074_ (.B(_2123_),
    .A(_2116_),
    .X(_2125_));
 sg13g2_a21oi_1 _4075_ (.A1(_2113_),
    .A2(_2119_),
    .Y(_2126_),
    .B1(_2118_));
 sg13g2_nor2b_1 _4076_ (.A(_2126_),
    .B_N(_0145_),
    .Y(_2127_));
 sg13g2_xor2_1 _4077_ (.B(_2127_),
    .A(_2125_),
    .X(_0146_));
 sg13g2_nor2_1 _4078_ (.A(\u_ddc_top_level.cic_left_inst.int_reg2[19] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[7] ),
    .Y(_2128_));
 sg13g2_xnor2_1 _4079_ (.Y(_2129_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg2[19] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[7] ));
 sg13g2_nand2b_1 _4080_ (.Y(_2130_),
    .B(_2129_),
    .A_N(_2122_));
 sg13g2_nor3_1 _4081_ (.A(\u_ddc_top_level.cic_left_inst.int_reg2[18] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[6] ),
    .C(_2129_),
    .Y(_2131_));
 sg13g2_xor2_1 _4082_ (.B(_2129_),
    .A(_2122_),
    .X(_2132_));
 sg13g2_nand2_1 _4083_ (.Y(_2133_),
    .A(_2124_),
    .B(_0146_));
 sg13g2_xnor2_1 _4084_ (.Y(_0147_),
    .A(_2132_),
    .B(_2133_));
 sg13g2_or2_1 _4085_ (.X(_2134_),
    .B(_2132_),
    .A(_2125_));
 sg13g2_nor2b_1 _4086_ (.A(_2134_),
    .B_N(_2126_),
    .Y(_2135_));
 sg13g2_nor4_1 _4087_ (.A(_2110_),
    .B(_2114_),
    .C(_2120_),
    .D(_2134_),
    .Y(_2136_));
 sg13g2_a21oi_1 _4088_ (.A1(_2124_),
    .A2(_2130_),
    .Y(_2137_),
    .B1(_2131_));
 sg13g2_or3_1 _4089_ (.A(_2135_),
    .B(_2136_),
    .C(_2137_),
    .X(_2138_));
 sg13g2_xnor2_1 _4090_ (.Y(_2139_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg2[20] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[8] ));
 sg13g2_nand2b_1 _4091_ (.Y(_2140_),
    .B(_2139_),
    .A_N(_2128_));
 sg13g2_xor2_1 _4092_ (.B(_2139_),
    .A(_2128_),
    .X(_2141_));
 sg13g2_xnor2_1 _4093_ (.Y(_0148_),
    .A(_2138_),
    .B(_2141_));
 sg13g2_nor2_1 _4094_ (.A(\u_ddc_top_level.cic_left_inst.int_reg2[21] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[9] ),
    .Y(_2142_));
 sg13g2_xnor2_1 _4095_ (.Y(_2143_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg2[21] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[9] ));
 sg13g2_nor3_1 _4096_ (.A(\u_ddc_top_level.cic_left_inst.int_reg2[20] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[8] ),
    .C(_2143_),
    .Y(_2144_));
 sg13g2_o21ai_1 _4097_ (.B1(_2143_),
    .Y(_2145_),
    .A1(\u_ddc_top_level.cic_left_inst.int_reg2[20] ),
    .A2(\u_ddc_top_level.dsm_left_inst.integrator1[8] ));
 sg13g2_nand2b_1 _4098_ (.Y(_2146_),
    .B(_2145_),
    .A_N(_2144_));
 sg13g2_nand2_1 _4099_ (.Y(_2147_),
    .A(_2140_),
    .B(_0148_));
 sg13g2_xnor2_1 _4100_ (.Y(_0149_),
    .A(_2146_),
    .B(_2147_));
 sg13g2_nor2_1 _4101_ (.A(\u_ddc_top_level.cic_left_inst.int_reg2[22] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[10] ),
    .Y(_2148_));
 sg13g2_xor2_1 _4102_ (.B(\u_ddc_top_level.dsm_left_inst.integrator1[10] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg2[22] ),
    .X(_2149_));
 sg13g2_nor2_1 _4103_ (.A(_2142_),
    .B(_2149_),
    .Y(_2150_));
 sg13g2_xnor2_1 _4104_ (.Y(_2151_),
    .A(_2142_),
    .B(_2149_));
 sg13g2_or2_1 _4105_ (.X(_2152_),
    .B(_2144_),
    .A(_2140_));
 sg13g2_nand2_1 _4106_ (.Y(_2153_),
    .A(_2145_),
    .B(_2152_));
 sg13g2_nand3_1 _4107_ (.B(_0149_),
    .C(_2152_),
    .A(_2145_),
    .Y(_2154_));
 sg13g2_xnor2_1 _4108_ (.Y(_0132_),
    .A(_2151_),
    .B(_2154_));
 sg13g2_nor2_1 _4109_ (.A(\u_ddc_top_level.cic_left_inst.int_reg2[23] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[11] ),
    .Y(_2155_));
 sg13g2_xnor2_1 _4110_ (.Y(_2156_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg2[23] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[11] ));
 sg13g2_nor2b_1 _4111_ (.A(_2148_),
    .B_N(_2156_),
    .Y(_2157_));
 sg13g2_or3_1 _4112_ (.A(\u_ddc_top_level.cic_left_inst.int_reg2[22] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[10] ),
    .C(_2156_),
    .X(_2158_));
 sg13g2_nand2b_1 _4113_ (.Y(_2159_),
    .B(_2158_),
    .A_N(_2157_));
 sg13g2_nand2b_1 _4114_ (.Y(_2160_),
    .B(_0132_),
    .A_N(_2150_));
 sg13g2_xnor2_1 _4115_ (.Y(_0133_),
    .A(_2159_),
    .B(_2160_));
 sg13g2_nor2_1 _4116_ (.A(_2151_),
    .B(_2159_),
    .Y(_2161_));
 sg13g2_nor4_1 _4117_ (.A(_2141_),
    .B(_2146_),
    .C(_2151_),
    .D(_2159_),
    .Y(_2162_));
 sg13g2_a21o_1 _4118_ (.A2(_2158_),
    .A1(_2150_),
    .B1(_2157_),
    .X(_2163_));
 sg13g2_a221oi_1 _4119_ (.B2(_2138_),
    .C1(_2163_),
    .B1(_2162_),
    .A1(_2153_),
    .Y(_2164_),
    .A2(_2161_));
 sg13g2_xnor2_1 _4120_ (.Y(_2165_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg2[24] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[12] ));
 sg13g2_nand2b_1 _4121_ (.Y(_2166_),
    .B(_2165_),
    .A_N(_2155_));
 sg13g2_xor2_1 _4122_ (.B(_2165_),
    .A(_2155_),
    .X(_2167_));
 sg13g2_xor2_1 _4123_ (.B(_2167_),
    .A(_2164_),
    .X(_0134_));
 sg13g2_nor2_1 _4124_ (.A(\u_ddc_top_level.cic_left_inst.int_reg2[25] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[13] ),
    .Y(_2168_));
 sg13g2_xnor2_1 _4125_ (.Y(_2169_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg2[25] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[13] ));
 sg13g2_o21ai_1 _4126_ (.B1(_2169_),
    .Y(_2170_),
    .A1(\u_ddc_top_level.cic_left_inst.int_reg2[24] ),
    .A2(\u_ddc_top_level.dsm_left_inst.integrator1[12] ));
 sg13g2_or3_1 _4127_ (.A(\u_ddc_top_level.cic_left_inst.int_reg2[24] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[12] ),
    .C(_2169_),
    .X(_2171_));
 sg13g2_nand2_1 _4128_ (.Y(_2172_),
    .A(_2170_),
    .B(_2171_));
 sg13g2_nand2_1 _4129_ (.Y(_2173_),
    .A(_2166_),
    .B(_0134_));
 sg13g2_xnor2_1 _4130_ (.Y(_0135_),
    .A(_2172_),
    .B(_2173_));
 sg13g2_nor2_1 _4131_ (.A(\u_ddc_top_level.cic_left_inst.int_reg2[26] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[14] ),
    .Y(_2174_));
 sg13g2_xor2_1 _4132_ (.B(\u_ddc_top_level.dsm_left_inst.integrator1[14] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg2[26] ),
    .X(_2175_));
 sg13g2_nor2_1 _4133_ (.A(_2168_),
    .B(_2175_),
    .Y(_2176_));
 sg13g2_xnor2_1 _4134_ (.Y(_2177_),
    .A(_2168_),
    .B(_2175_));
 sg13g2_or2_1 _4135_ (.X(_2178_),
    .B(_2172_),
    .A(_2167_));
 sg13g2_nand2b_1 _4136_ (.Y(_2179_),
    .B(_2171_),
    .A_N(_2166_));
 sg13g2_and2_1 _4137_ (.A(_2170_),
    .B(_2179_),
    .X(_2180_));
 sg13g2_o21ai_1 _4138_ (.B1(_2180_),
    .Y(_2181_),
    .A1(_2164_),
    .A2(_2178_));
 sg13g2_nand2b_1 _4139_ (.Y(_2182_),
    .B(_2181_),
    .A_N(_2177_));
 sg13g2_xnor2_1 _4140_ (.Y(_0136_),
    .A(_2177_),
    .B(_2181_));
 sg13g2_xor2_1 _4141_ (.B(\u_ddc_top_level.dsm_left_inst.integrator1[15] ),
    .A(\u_ddc_top_level.cic_left_inst.int_reg2[27] ),
    .X(_2183_));
 sg13g2_nand2_1 _4142_ (.Y(_2184_),
    .A(_2174_),
    .B(_2183_));
 sg13g2_nor2_1 _4143_ (.A(_2174_),
    .B(_2183_),
    .Y(_2185_));
 sg13g2_xnor2_1 _4144_ (.Y(_2186_),
    .A(_2174_),
    .B(_2183_));
 sg13g2_nand2b_1 _4145_ (.Y(_2187_),
    .B(_0136_),
    .A_N(_2176_));
 sg13g2_xnor2_1 _4146_ (.Y(_0137_),
    .A(_2186_),
    .B(_2187_));
 sg13g2_nand2_1 _4147_ (.Y(_2188_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg2[27] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[16] ));
 sg13g2_a21oi_1 _4148_ (.A1(\u_ddc_top_level.dsm_left_inst.integrator1[15] ),
    .A2(\u_ddc_top_level.dsm_left_inst.integrator1[16] ),
    .Y(_2189_),
    .B1(\u_ddc_top_level.cic_left_inst.int_reg2[27] ));
 sg13g2_nor2b_1 _4149_ (.A(_2189_),
    .B_N(_2188_),
    .Y(_2190_));
 sg13g2_or3_1 _4150_ (.A(\u_ddc_top_level.cic_left_inst.int_reg2[27] ),
    .B(\u_ddc_top_level.dsm_left_inst.integrator1[15] ),
    .C(\u_ddc_top_level.dsm_left_inst.integrator1[16] ),
    .X(_2191_));
 sg13g2_nor2b_1 _4151_ (.A(_2190_),
    .B_N(_2191_),
    .Y(_2192_));
 sg13g2_a21oi_1 _4152_ (.A1(_2176_),
    .A2(_2184_),
    .Y(_2193_),
    .B1(_2185_));
 sg13g2_o21ai_1 _4153_ (.B1(_2193_),
    .Y(_2194_),
    .A1(_2182_),
    .A2(_2186_));
 sg13g2_xor2_1 _4154_ (.B(_2194_),
    .A(_2192_),
    .X(_0138_));
 sg13g2_nor2b_1 _4155_ (.A(_2190_),
    .B_N(_0138_),
    .Y(_2195_));
 sg13g2_nand2b_1 _4156_ (.Y(_2196_),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[27] ),
    .A_N(\u_ddc_top_level.dsm_left_inst.feedback[17] ));
 sg13g2_nor2b_1 _4157_ (.A(\u_ddc_top_level.cic_left_inst.int_reg2[27] ),
    .B_N(\u_ddc_top_level.dsm_left_inst.feedback[17] ),
    .Y(_2197_));
 sg13g2_xnor2_1 _4158_ (.Y(_2198_),
    .A(\u_ddc_top_level.dsm_left_inst.feedback[17] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg2[27] ));
 sg13g2_xnor2_1 _4159_ (.Y(_2199_),
    .A(\u_ddc_top_level.dsm_left_inst.integrator1[17] ),
    .B(_2198_));
 sg13g2_xor2_1 _4160_ (.B(_2199_),
    .A(_2188_),
    .X(_2200_));
 sg13g2_xnor2_1 _4161_ (.Y(_0139_),
    .A(_2195_),
    .B(_2200_));
 sg13g2_nand3_1 _4162_ (.B(_2194_),
    .C(_2200_),
    .A(_2192_),
    .Y(_2201_));
 sg13g2_o21ai_1 _4163_ (.B1(_2201_),
    .Y(_2202_),
    .A1(_2189_),
    .A2(_2199_));
 sg13g2_o21ai_1 _4164_ (.B1(_2196_),
    .Y(_2203_),
    .A1(\u_ddc_top_level.dsm_left_inst.integrator1[17] ),
    .A2(_2197_));
 sg13g2_xnor2_1 _4165_ (.Y(_2204_),
    .A(\u_ddc_top_level.dsm_left_inst.integrator1[18] ),
    .B(_2203_));
 sg13g2_xnor2_1 _4166_ (.Y(_0140_),
    .A(_2202_),
    .B(_2204_));
 sg13g2_nand2_1 _4167_ (.Y(_2205_),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[0] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[0] ));
 sg13g2_xor2_1 _4168_ (.B(\u_ddc_top_level.dsm_right_inst.integrator2[0] ),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[0] ),
    .X(_2206_));
 sg13g2_xnor2_1 _4169_ (.Y(_0112_),
    .A(_0006_),
    .B(_2206_));
 sg13g2_or2_1 _4170_ (.X(_2207_),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[1] ),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[1] ));
 sg13g2_nand2_1 _4171_ (.Y(_2208_),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[1] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[1] ));
 sg13g2_nand2_1 _4172_ (.Y(_2209_),
    .A(_2207_),
    .B(_2208_));
 sg13g2_o21ai_1 _4173_ (.B1(\u_ddc_top_level.dsm_left_inst.in_dither ),
    .Y(_2210_),
    .A1(\u_ddc_top_level.dsm_right_inst.integrator1[0] ),
    .A2(\u_ddc_top_level.dsm_right_inst.integrator2[0] ));
 sg13g2_nand2_1 _4174_ (.Y(_2211_),
    .A(_2205_),
    .B(_2210_));
 sg13g2_nand4_1 _4175_ (.B(_2207_),
    .C(_2208_),
    .A(_2205_),
    .Y(_2212_),
    .D(_2210_));
 sg13g2_xnor2_1 _4176_ (.Y(_0122_),
    .A(_2209_),
    .B(_2211_));
 sg13g2_nor2_1 _4177_ (.A(\u_ddc_top_level.dsm_right_inst.integrator1[2] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[2] ),
    .Y(_2213_));
 sg13g2_xnor2_1 _4178_ (.Y(_2214_),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[2] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[2] ));
 sg13g2_a21oi_1 _4179_ (.A1(_2207_),
    .A2(_2212_),
    .Y(_2215_),
    .B1(_2214_));
 sg13g2_nand3_1 _4180_ (.B(_2212_),
    .C(_2214_),
    .A(_2207_),
    .Y(_2216_));
 sg13g2_nand2b_1 _4181_ (.Y(_0123_),
    .B(_2216_),
    .A_N(_2215_));
 sg13g2_nor2_1 _4182_ (.A(\u_ddc_top_level.dsm_right_inst.integrator1[3] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[3] ),
    .Y(_2217_));
 sg13g2_xnor2_1 _4183_ (.Y(_2218_),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[3] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[3] ));
 sg13g2_inv_1 _4184_ (.Y(_2219_),
    .A(_2218_));
 sg13g2_o21ai_1 _4185_ (.B1(_2219_),
    .Y(_2220_),
    .A1(_2213_),
    .A2(_2215_));
 sg13g2_or3_1 _4186_ (.A(_2213_),
    .B(_2215_),
    .C(_2219_),
    .X(_2221_));
 sg13g2_nand2_1 _4187_ (.Y(_0124_),
    .A(_2220_),
    .B(_2221_));
 sg13g2_xor2_1 _4188_ (.B(\u_ddc_top_level.dsm_right_inst.integrator2[4] ),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[4] ),
    .X(_2222_));
 sg13g2_or2_1 _4189_ (.X(_2223_),
    .B(_2222_),
    .A(_2217_));
 sg13g2_xnor2_1 _4190_ (.Y(_2224_),
    .A(_2217_),
    .B(_2222_));
 sg13g2_xnor2_1 _4191_ (.Y(_0125_),
    .A(_2220_),
    .B(_2224_));
 sg13g2_nand2_1 _4192_ (.Y(_2225_),
    .A(_2223_),
    .B(_0125_));
 sg13g2_nor2_1 _4193_ (.A(\u_ddc_top_level.dsm_right_inst.integrator1[5] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[5] ),
    .Y(_2226_));
 sg13g2_xnor2_1 _4194_ (.Y(_2227_),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[5] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[5] ));
 sg13g2_nor3_1 _4195_ (.A(\u_ddc_top_level.dsm_right_inst.integrator1[4] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[4] ),
    .C(_2227_),
    .Y(_2228_));
 sg13g2_o21ai_1 _4196_ (.B1(_2227_),
    .Y(_2229_),
    .A1(\u_ddc_top_level.dsm_right_inst.integrator1[4] ),
    .A2(\u_ddc_top_level.dsm_right_inst.integrator2[4] ));
 sg13g2_nand2b_1 _4197_ (.Y(_2230_),
    .B(_2229_),
    .A_N(_2228_));
 sg13g2_xnor2_1 _4198_ (.Y(_0126_),
    .A(_2225_),
    .B(_2230_));
 sg13g2_nor2_1 _4199_ (.A(\u_ddc_top_level.dsm_right_inst.integrator1[6] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[6] ),
    .Y(_2231_));
 sg13g2_xnor2_1 _4200_ (.Y(_2232_),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[6] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[6] ));
 sg13g2_nand2b_1 _4201_ (.Y(_2233_),
    .B(_2232_),
    .A_N(_2226_));
 sg13g2_xor2_1 _4202_ (.B(_2232_),
    .A(_2226_),
    .X(_2234_));
 sg13g2_a21oi_1 _4203_ (.A1(_2223_),
    .A2(_2229_),
    .Y(_2235_),
    .B1(_2228_));
 sg13g2_inv_1 _4204_ (.Y(_2236_),
    .A(_2235_));
 sg13g2_nand2_1 _4205_ (.Y(_2237_),
    .A(_0126_),
    .B(_2236_));
 sg13g2_xnor2_1 _4206_ (.Y(_0127_),
    .A(_2234_),
    .B(_2237_));
 sg13g2_nor2_1 _4207_ (.A(\u_ddc_top_level.dsm_right_inst.integrator1[7] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[7] ),
    .Y(_2238_));
 sg13g2_xor2_1 _4208_ (.B(\u_ddc_top_level.dsm_right_inst.integrator2[7] ),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[7] ),
    .X(_2239_));
 sg13g2_xnor2_1 _4209_ (.Y(_2240_),
    .A(_2231_),
    .B(_2239_));
 sg13g2_nand2_1 _4210_ (.Y(_2241_),
    .A(_2233_),
    .B(_0127_));
 sg13g2_xnor2_1 _4211_ (.Y(_0128_),
    .A(_2240_),
    .B(_2241_));
 sg13g2_nor2_1 _4212_ (.A(_2234_),
    .B(_2240_),
    .Y(_2242_));
 sg13g2_nor4_1 _4213_ (.A(_2224_),
    .B(_2230_),
    .C(_2234_),
    .D(_2240_),
    .Y(_2243_));
 sg13g2_a21o_1 _4214_ (.A2(_2239_),
    .A1(_2231_),
    .B1(_2233_),
    .X(_2244_));
 sg13g2_o21ai_1 _4215_ (.B1(_2244_),
    .Y(_2245_),
    .A1(_2231_),
    .A2(_2239_));
 sg13g2_a221oi_1 _4216_ (.B2(_2220_),
    .C1(_2245_),
    .B1(_2243_),
    .A1(_2235_),
    .Y(_2246_),
    .A2(_2242_));
 sg13g2_xnor2_1 _4217_ (.Y(_2247_),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[8] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[8] ));
 sg13g2_nor2b_1 _4218_ (.A(_2238_),
    .B_N(_2247_),
    .Y(_2248_));
 sg13g2_xor2_1 _4219_ (.B(_2247_),
    .A(_2238_),
    .X(_2249_));
 sg13g2_xor2_1 _4220_ (.B(_2249_),
    .A(_2246_),
    .X(_0129_));
 sg13g2_nor2_1 _4221_ (.A(\u_ddc_top_level.dsm_right_inst.integrator1[9] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[9] ),
    .Y(_2250_));
 sg13g2_xnor2_1 _4222_ (.Y(_2251_),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[9] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[9] ));
 sg13g2_or3_1 _4223_ (.A(\u_ddc_top_level.dsm_right_inst.integrator1[8] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[8] ),
    .C(_2251_),
    .X(_2252_));
 sg13g2_o21ai_1 _4224_ (.B1(_2251_),
    .Y(_2253_),
    .A1(\u_ddc_top_level.dsm_right_inst.integrator1[8] ),
    .A2(\u_ddc_top_level.dsm_right_inst.integrator2[8] ));
 sg13g2_nand2_1 _4225_ (.Y(_2254_),
    .A(_2252_),
    .B(_2253_));
 sg13g2_nand2b_1 _4226_ (.Y(_2255_),
    .B(_0129_),
    .A_N(_2248_));
 sg13g2_xnor2_1 _4227_ (.Y(_0130_),
    .A(_2254_),
    .B(_2255_));
 sg13g2_xnor2_1 _4228_ (.Y(_2256_),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[10] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[10] ));
 sg13g2_nor2b_1 _4229_ (.A(_2250_),
    .B_N(_2256_),
    .Y(_2257_));
 sg13g2_xor2_1 _4230_ (.B(_2256_),
    .A(_2250_),
    .X(_2258_));
 sg13g2_nand2_1 _4231_ (.Y(_2259_),
    .A(_2248_),
    .B(_2252_));
 sg13g2_nand2_1 _4232_ (.Y(_2260_),
    .A(_2253_),
    .B(_2259_));
 sg13g2_nand3_1 _4233_ (.B(_0130_),
    .C(_2259_),
    .A(_2253_),
    .Y(_2261_));
 sg13g2_xnor2_1 _4234_ (.Y(_0113_),
    .A(_2258_),
    .B(_2261_));
 sg13g2_nor2_1 _4235_ (.A(\u_ddc_top_level.dsm_right_inst.integrator1[11] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[11] ),
    .Y(_2262_));
 sg13g2_xnor2_1 _4236_ (.Y(_2263_),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[11] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[11] ));
 sg13g2_o21ai_1 _4237_ (.B1(_2263_),
    .Y(_2264_),
    .A1(\u_ddc_top_level.dsm_right_inst.integrator1[10] ),
    .A2(\u_ddc_top_level.dsm_right_inst.integrator2[10] ));
 sg13g2_or3_1 _4238_ (.A(\u_ddc_top_level.dsm_right_inst.integrator1[10] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[10] ),
    .C(_2263_),
    .X(_2265_));
 sg13g2_nand2_1 _4239_ (.Y(_2266_),
    .A(_2264_),
    .B(_2265_));
 sg13g2_nand2b_1 _4240_ (.Y(_2267_),
    .B(_0113_),
    .A_N(_2257_));
 sg13g2_xnor2_1 _4241_ (.Y(_0114_),
    .A(_2266_),
    .B(_2267_));
 sg13g2_nor2_1 _4242_ (.A(_2258_),
    .B(_2266_),
    .Y(_2268_));
 sg13g2_or4_1 _4243_ (.A(_2249_),
    .B(_2254_),
    .C(_2258_),
    .D(_2266_),
    .X(_2269_));
 sg13g2_nand2b_1 _4244_ (.Y(_2270_),
    .B(_2264_),
    .A_N(_2257_));
 sg13g2_a22oi_1 _4245_ (.Y(_2271_),
    .B1(_2270_),
    .B2(_2265_),
    .A2(_2268_),
    .A1(_2260_));
 sg13g2_o21ai_1 _4246_ (.B1(_2271_),
    .Y(_2272_),
    .A1(_2246_),
    .A2(_2269_));
 sg13g2_xnor2_1 _4247_ (.Y(_2273_),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[12] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[12] ));
 sg13g2_nand2b_1 _4248_ (.Y(_2274_),
    .B(_2273_),
    .A_N(_2262_));
 sg13g2_xor2_1 _4249_ (.B(_2273_),
    .A(_2262_),
    .X(_2275_));
 sg13g2_xnor2_1 _4250_ (.Y(_0115_),
    .A(_2272_),
    .B(_2275_));
 sg13g2_nand2_1 _4251_ (.Y(_2276_),
    .A(_2274_),
    .B(_0115_));
 sg13g2_xnor2_1 _4252_ (.Y(_2277_),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[13] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[13] ));
 sg13g2_or3_1 _4253_ (.A(\u_ddc_top_level.dsm_right_inst.integrator1[12] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[12] ),
    .C(_2277_),
    .X(_2278_));
 sg13g2_o21ai_1 _4254_ (.B1(_2277_),
    .Y(_2279_),
    .A1(\u_ddc_top_level.dsm_right_inst.integrator1[12] ),
    .A2(\u_ddc_top_level.dsm_right_inst.integrator2[12] ));
 sg13g2_nand2_1 _4255_ (.Y(_2280_),
    .A(_2278_),
    .B(_2279_));
 sg13g2_xnor2_1 _4256_ (.Y(_0116_),
    .A(_2276_),
    .B(_2280_));
 sg13g2_xnor2_1 _4257_ (.Y(_2281_),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[14] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[14] ));
 sg13g2_o21ai_1 _4258_ (.B1(_2281_),
    .Y(_2282_),
    .A1(\u_ddc_top_level.dsm_right_inst.integrator1[13] ),
    .A2(\u_ddc_top_level.dsm_right_inst.integrator2[13] ));
 sg13g2_or3_1 _4259_ (.A(\u_ddc_top_level.dsm_right_inst.integrator1[13] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[13] ),
    .C(_2281_),
    .X(_2283_));
 sg13g2_nand2_1 _4260_ (.Y(_2284_),
    .A(_2282_),
    .B(_2283_));
 sg13g2_nor2_1 _4261_ (.A(_2275_),
    .B(_2280_),
    .Y(_2285_));
 sg13g2_nand2_1 _4262_ (.Y(_2286_),
    .A(_2274_),
    .B(_2279_));
 sg13g2_a22oi_1 _4263_ (.Y(_2287_),
    .B1(_2286_),
    .B2(_2278_),
    .A2(_2285_),
    .A1(_2272_));
 sg13g2_xor2_1 _4264_ (.B(_2287_),
    .A(_2284_),
    .X(_0117_));
 sg13g2_nor2_1 _4265_ (.A(\u_ddc_top_level.dsm_right_inst.integrator1[15] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[15] ),
    .Y(_2288_));
 sg13g2_xnor2_1 _4266_ (.Y(_2289_),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[15] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[15] ));
 sg13g2_or3_1 _4267_ (.A(\u_ddc_top_level.dsm_right_inst.integrator1[14] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[14] ),
    .C(_2289_),
    .X(_2290_));
 sg13g2_o21ai_1 _4268_ (.B1(_2289_),
    .Y(_2291_),
    .A1(\u_ddc_top_level.dsm_right_inst.integrator1[14] ),
    .A2(\u_ddc_top_level.dsm_right_inst.integrator2[14] ));
 sg13g2_nand2_1 _4269_ (.Y(_2292_),
    .A(_2290_),
    .B(_2291_));
 sg13g2_nand2_1 _4270_ (.Y(_2293_),
    .A(_2282_),
    .B(_0117_));
 sg13g2_xnor2_1 _4271_ (.Y(_0118_),
    .A(_2292_),
    .B(_2293_));
 sg13g2_nor2_1 _4272_ (.A(\u_ddc_top_level.dsm_right_inst.integrator1[16] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[16] ),
    .Y(_2294_));
 sg13g2_xor2_1 _4273_ (.B(\u_ddc_top_level.dsm_right_inst.integrator2[16] ),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[16] ),
    .X(_2295_));
 sg13g2_nor2_1 _4274_ (.A(_2288_),
    .B(_2295_),
    .Y(_2296_));
 sg13g2_xor2_1 _4275_ (.B(_2295_),
    .A(_2288_),
    .X(_2297_));
 sg13g2_nand2_1 _4276_ (.Y(_2298_),
    .A(_2282_),
    .B(_2291_));
 sg13g2_a221oi_1 _4277_ (.B2(_2278_),
    .C1(_2298_),
    .B1(_2286_),
    .A1(_2272_),
    .Y(_2299_),
    .A2(_2285_));
 sg13g2_o21ai_1 _4278_ (.B1(_2290_),
    .Y(_2300_),
    .A1(_2283_),
    .A2(_2289_));
 sg13g2_o21ai_1 _4279_ (.B1(_2297_),
    .Y(_2301_),
    .A1(_2299_),
    .A2(_2300_));
 sg13g2_or3_1 _4280_ (.A(_2297_),
    .B(_2299_),
    .C(_2300_),
    .X(_2302_));
 sg13g2_nand2_1 _4281_ (.Y(_0119_),
    .A(_2301_),
    .B(_2302_));
 sg13g2_a21oi_1 _4282_ (.A1(_2301_),
    .A2(_2302_),
    .Y(_2303_),
    .B1(_2296_));
 sg13g2_nand2_1 _4283_ (.Y(_2304_),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[17] ),
    .B(\u_ddc_top_level.dsm_right_inst.integrator2[17] ));
 sg13g2_xor2_1 _4284_ (.B(\u_ddc_top_level.dsm_right_inst.integrator2[17] ),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[17] ),
    .X(_2305_));
 sg13g2_xnor2_1 _4285_ (.Y(_2306_),
    .A(_2294_),
    .B(_2305_));
 sg13g2_xnor2_1 _4286_ (.Y(_0120_),
    .A(_2303_),
    .B(_2306_));
 sg13g2_nand2b_1 _4287_ (.Y(_2307_),
    .B(_0120_),
    .A_N(_2305_));
 sg13g2_xnor2_1 _4288_ (.Y(_2308_),
    .A(\u_ddc_top_level.dsm_right_inst.integrator1[18] ),
    .B(_2304_));
 sg13g2_xnor2_1 _4289_ (.Y(_0121_),
    .A(_2307_),
    .B(_2308_));
 sg13g2_nor2_1 _4290_ (.A(_0111_),
    .B(net885),
    .Y(_2309_));
 sg13g2_xor2_1 _4291_ (.B(\u_ddc_top_level.lsfr_inst.lfsr_reg[4] ),
    .A(\u_ddc_top_level.lsfr_inst.lfsr_reg[13] ),
    .X(_2310_));
 sg13g2_xor2_1 _4292_ (.B(\u_ddc_top_level.lsfr_inst.lfsr_reg[15] ),
    .A(\u_ddc_top_level.dsm_left_inst.in_dither ),
    .X(_2311_));
 sg13g2_xnor2_1 _4293_ (.Y(_2312_),
    .A(_2310_),
    .B(_2311_));
 sg13g2_a21oi_1 _4294_ (.A1(net885),
    .A2(_2312_),
    .Y(_0398_),
    .B1(_2309_));
 sg13g2_mux2_1 _4295_ (.A0(\u_ddc_top_level.lsfr_inst.lfsr_reg[1] ),
    .A1(\u_ddc_top_level.lsfr_inst.lfsr_reg[0] ),
    .S(net885),
    .X(_0399_));
 sg13g2_mux2_1 _4296_ (.A0(\u_ddc_top_level.lsfr_inst.lfsr_reg[2] ),
    .A1(\u_ddc_top_level.lsfr_inst.lfsr_reg[1] ),
    .S(net885),
    .X(_0400_));
 sg13g2_mux2_1 _4297_ (.A0(\u_ddc_top_level.lsfr_inst.lfsr_reg[3] ),
    .A1(\u_ddc_top_level.lsfr_inst.lfsr_reg[2] ),
    .S(net885),
    .X(_0401_));
 sg13g2_mux2_1 _4298_ (.A0(\u_ddc_top_level.lsfr_inst.lfsr_reg[4] ),
    .A1(\u_ddc_top_level.lsfr_inst.lfsr_reg[3] ),
    .S(net885),
    .X(_0402_));
 sg13g2_mux2_1 _4299_ (.A0(\u_ddc_top_level.lsfr_inst.lfsr_reg[5] ),
    .A1(\u_ddc_top_level.lsfr_inst.lfsr_reg[4] ),
    .S(net3),
    .X(_0403_));
 sg13g2_mux2_1 _4300_ (.A0(\u_ddc_top_level.lsfr_inst.lfsr_reg[6] ),
    .A1(\u_ddc_top_level.lsfr_inst.lfsr_reg[5] ),
    .S(net3),
    .X(_0404_));
 sg13g2_mux2_1 _4301_ (.A0(\u_ddc_top_level.lsfr_inst.lfsr_reg[7] ),
    .A1(\u_ddc_top_level.lsfr_inst.lfsr_reg[6] ),
    .S(net3),
    .X(_0405_));
 sg13g2_mux2_1 _4302_ (.A0(\u_ddc_top_level.lsfr_inst.lfsr_reg[8] ),
    .A1(\u_ddc_top_level.lsfr_inst.lfsr_reg[7] ),
    .S(net886),
    .X(_0406_));
 sg13g2_mux2_1 _4303_ (.A0(\u_ddc_top_level.lsfr_inst.lfsr_reg[9] ),
    .A1(\u_ddc_top_level.lsfr_inst.lfsr_reg[8] ),
    .S(net886),
    .X(_0407_));
 sg13g2_mux2_1 _4304_ (.A0(\u_ddc_top_level.lsfr_inst.lfsr_reg[10] ),
    .A1(\u_ddc_top_level.lsfr_inst.lfsr_reg[9] ),
    .S(net886),
    .X(_0408_));
 sg13g2_mux2_1 _4305_ (.A0(\u_ddc_top_level.lsfr_inst.lfsr_reg[11] ),
    .A1(\u_ddc_top_level.lsfr_inst.lfsr_reg[10] ),
    .S(net886),
    .X(_0409_));
 sg13g2_mux2_1 _4306_ (.A0(\u_ddc_top_level.lsfr_inst.lfsr_reg[12] ),
    .A1(\u_ddc_top_level.lsfr_inst.lfsr_reg[11] ),
    .S(net886),
    .X(_0410_));
 sg13g2_mux2_1 _4307_ (.A0(\u_ddc_top_level.lsfr_inst.lfsr_reg[13] ),
    .A1(\u_ddc_top_level.lsfr_inst.lfsr_reg[12] ),
    .S(net886),
    .X(_0411_));
 sg13g2_mux2_1 _4308_ (.A0(\u_ddc_top_level.lsfr_inst.lfsr_reg[14] ),
    .A1(\u_ddc_top_level.lsfr_inst.lfsr_reg[13] ),
    .S(net885),
    .X(_0412_));
 sg13g2_mux2_1 _4309_ (.A0(\u_ddc_top_level.lsfr_inst.lfsr_reg[15] ),
    .A1(\u_ddc_top_level.lsfr_inst.lfsr_reg[14] ),
    .S(net885),
    .X(_0413_));
 sg13g2_mux2_1 _4310_ (.A0(\u_ddc_top_level.dsm_left_inst.in_dither ),
    .A1(\u_ddc_top_level.lsfr_inst.lfsr_reg[15] ),
    .S(net886),
    .X(_0414_));
 sg13g2_or3_1 _4311_ (.A(\u_ddc_top_level.i2s_rx_inst.bit_count[5] ),
    .B(\u_ddc_top_level.i2s_rx_inst.bit_count[4] ),
    .C(_1400_),
    .X(_2313_));
 sg13g2_mux2_1 _4312_ (.A0(net2),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[0] ),
    .S(net806),
    .X(_0415_));
 sg13g2_mux2_1 _4313_ (.A0(\u_ddc_top_level.i2s_rx_inst.shift_reg[0] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[1] ),
    .S(net806),
    .X(_0416_));
 sg13g2_mux2_1 _4314_ (.A0(\u_ddc_top_level.i2s_rx_inst.shift_reg[1] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[2] ),
    .S(net806),
    .X(_0417_));
 sg13g2_mux2_1 _4315_ (.A0(\u_ddc_top_level.i2s_rx_inst.shift_reg[2] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[3] ),
    .S(net806),
    .X(_0418_));
 sg13g2_mux2_1 _4316_ (.A0(\u_ddc_top_level.i2s_rx_inst.shift_reg[3] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[4] ),
    .S(net806),
    .X(_0419_));
 sg13g2_mux2_1 _4317_ (.A0(\u_ddc_top_level.i2s_rx_inst.shift_reg[4] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[5] ),
    .S(net806),
    .X(_0420_));
 sg13g2_mux2_1 _4318_ (.A0(\u_ddc_top_level.i2s_rx_inst.shift_reg[5] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[6] ),
    .S(net806),
    .X(_0421_));
 sg13g2_mux2_1 _4319_ (.A0(\u_ddc_top_level.i2s_rx_inst.shift_reg[6] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[7] ),
    .S(net806),
    .X(_0422_));
 sg13g2_mux2_1 _4320_ (.A0(\u_ddc_top_level.i2s_rx_inst.shift_reg[7] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[8] ),
    .S(net807),
    .X(_0423_));
 sg13g2_mux2_1 _4321_ (.A0(\u_ddc_top_level.i2s_rx_inst.shift_reg[8] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[9] ),
    .S(net807),
    .X(_0424_));
 sg13g2_mux2_1 _4322_ (.A0(\u_ddc_top_level.i2s_rx_inst.shift_reg[9] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[10] ),
    .S(net807),
    .X(_0425_));
 sg13g2_mux2_1 _4323_ (.A0(\u_ddc_top_level.i2s_rx_inst.shift_reg[10] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[11] ),
    .S(net807),
    .X(_0426_));
 sg13g2_mux2_1 _4324_ (.A0(\u_ddc_top_level.i2s_rx_inst.shift_reg[11] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[12] ),
    .S(net807),
    .X(_0427_));
 sg13g2_mux2_1 _4325_ (.A0(\u_ddc_top_level.i2s_rx_inst.shift_reg[12] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[13] ),
    .S(net807),
    .X(_0428_));
 sg13g2_mux2_1 _4326_ (.A0(\u_ddc_top_level.i2s_rx_inst.shift_reg[13] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[14] ),
    .S(_2313_),
    .X(_0429_));
 sg13g2_mux2_1 _4327_ (.A0(\u_ddc_top_level.i2s_rx_inst.shift_reg[14] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[15] ),
    .S(net807),
    .X(_0430_));
 sg13g2_nand2_1 _4328_ (.Y(_2314_),
    .A(net852),
    .B(\u_ddc_top_level.cic_right_inst.comb_out2[0] ));
 sg13g2_xnor2_1 _4329_ (.Y(_0518_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg0[0] ),
    .B(_2314_));
 sg13g2_nand2_1 _4330_ (.Y(_2315_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[0] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[0] ));
 sg13g2_nand2_1 _4331_ (.Y(_2316_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[1] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[1] ));
 sg13g2_xnor2_1 _4332_ (.Y(_2317_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[1] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[1] ));
 sg13g2_nor2_1 _4333_ (.A(net852),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[1] ),
    .Y(_2318_));
 sg13g2_xnor2_1 _4334_ (.Y(_2319_),
    .A(_2315_),
    .B(_2317_));
 sg13g2_a21oi_1 _4335_ (.A1(net852),
    .A2(_2319_),
    .Y(_0519_),
    .B1(_2318_));
 sg13g2_nor2_1 _4336_ (.A(net853),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[2] ),
    .Y(_2320_));
 sg13g2_and2_1 _4337_ (.A(\u_ddc_top_level.cic_right_inst.comb_out2[2] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[2] ),
    .X(_2321_));
 sg13g2_xor2_1 _4338_ (.B(\u_ddc_top_level.cic_right_inst.int_reg0[2] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[2] ),
    .X(_2322_));
 sg13g2_o21ai_1 _4339_ (.B1(_2316_),
    .Y(_2323_),
    .A1(_2315_),
    .A2(_2317_));
 sg13g2_xnor2_1 _4340_ (.Y(_2324_),
    .A(_2322_),
    .B(_2323_));
 sg13g2_a21oi_1 _4341_ (.A1(net853),
    .A2(_2324_),
    .Y(_0520_),
    .B1(_2320_));
 sg13g2_nor2_1 _4342_ (.A(net853),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[3] ),
    .Y(_2325_));
 sg13g2_nand2_1 _4343_ (.Y(_2326_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[3] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[3] ));
 sg13g2_xnor2_1 _4344_ (.Y(_2327_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[3] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[3] ));
 sg13g2_a21oi_1 _4345_ (.A1(_2322_),
    .A2(_2323_),
    .Y(_2328_),
    .B1(_2321_));
 sg13g2_xnor2_1 _4346_ (.Y(_2329_),
    .A(_2327_),
    .B(_2328_));
 sg13g2_a21oi_1 _4347_ (.A1(net853),
    .A2(_2329_),
    .Y(_0521_),
    .B1(_2325_));
 sg13g2_o21ai_1 _4348_ (.B1(_2326_),
    .Y(_2330_),
    .A1(_2327_),
    .A2(_2328_));
 sg13g2_and2_1 _4349_ (.A(\u_ddc_top_level.cic_right_inst.comb_out2[4] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[4] ),
    .X(_2331_));
 sg13g2_xor2_1 _4350_ (.B(\u_ddc_top_level.cic_right_inst.int_reg0[4] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[4] ),
    .X(_2332_));
 sg13g2_inv_1 _4351_ (.Y(_2333_),
    .A(_2332_));
 sg13g2_o21ai_1 _4352_ (.B1(net856),
    .Y(_2334_),
    .A1(_2330_),
    .A2(_2332_));
 sg13g2_a21oi_1 _4353_ (.A1(_2330_),
    .A2(_2332_),
    .Y(_2335_),
    .B1(_2334_));
 sg13g2_a21o_1 _4354_ (.A2(\u_ddc_top_level.cic_right_inst.int_reg0[4] ),
    .A1(net813),
    .B1(_2335_),
    .X(_0522_));
 sg13g2_or2_1 _4355_ (.X(_2336_),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[5] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[5] ));
 sg13g2_and2_1 _4356_ (.A(\u_ddc_top_level.cic_right_inst.comb_out2[5] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[5] ),
    .X(_2337_));
 sg13g2_xnor2_1 _4357_ (.Y(_2338_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[5] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[5] ));
 sg13g2_a21oi_1 _4358_ (.A1(_2330_),
    .A2(_2332_),
    .Y(_2339_),
    .B1(_2331_));
 sg13g2_xnor2_1 _4359_ (.Y(_2340_),
    .A(_2338_),
    .B(_2339_));
 sg13g2_nor2_1 _4360_ (.A(net863),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[5] ),
    .Y(_2341_));
 sg13g2_a21oi_1 _4361_ (.A1(net853),
    .A2(_2340_),
    .Y(_0523_),
    .B1(_2341_));
 sg13g2_and2_1 _4362_ (.A(\u_ddc_top_level.cic_right_inst.comb_out2[6] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[6] ),
    .X(_2342_));
 sg13g2_nor2_1 _4363_ (.A(\u_ddc_top_level.cic_right_inst.comb_out2[6] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[6] ),
    .Y(_2343_));
 sg13g2_nor2_1 _4364_ (.A(_2342_),
    .B(_2343_),
    .Y(_2344_));
 sg13g2_nor2_1 _4365_ (.A(_2333_),
    .B(_2338_),
    .Y(_2345_));
 sg13g2_nand2_1 _4366_ (.Y(_2346_),
    .A(_2330_),
    .B(_2345_));
 sg13g2_a21oi_1 _4367_ (.A1(_2331_),
    .A2(_2336_),
    .Y(_2347_),
    .B1(_2337_));
 sg13g2_nand2_1 _4368_ (.Y(_2348_),
    .A(_2346_),
    .B(_2347_));
 sg13g2_o21ai_1 _4369_ (.B1(net856),
    .Y(_2349_),
    .A1(_2344_),
    .A2(_2348_));
 sg13g2_a21oi_1 _4370_ (.A1(_2344_),
    .A2(_2348_),
    .Y(_2350_),
    .B1(_2349_));
 sg13g2_a21o_1 _4371_ (.A2(\u_ddc_top_level.cic_right_inst.int_reg0[6] ),
    .A1(net813),
    .B1(_2350_),
    .X(_0524_));
 sg13g2_nand2_1 _4372_ (.Y(_2351_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[7] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[7] ));
 sg13g2_nor2_1 _4373_ (.A(\u_ddc_top_level.cic_right_inst.comb_out2[7] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[7] ),
    .Y(_2352_));
 sg13g2_xor2_1 _4374_ (.B(\u_ddc_top_level.cic_right_inst.int_reg0[7] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[7] ),
    .X(_2353_));
 sg13g2_a21o_1 _4375_ (.A2(_2348_),
    .A1(_2344_),
    .B1(_2342_),
    .X(_2354_));
 sg13g2_xnor2_1 _4376_ (.Y(_2355_),
    .A(_2353_),
    .B(_2354_));
 sg13g2_nor2_1 _4377_ (.A(net853),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[7] ),
    .Y(_2356_));
 sg13g2_a21oi_1 _4378_ (.A1(net856),
    .A2(_2355_),
    .Y(_0525_),
    .B1(_2356_));
 sg13g2_nand2b_1 _4379_ (.Y(_2357_),
    .B(_2342_),
    .A_N(_2352_));
 sg13g2_nand3_1 _4380_ (.B(_2351_),
    .C(_2357_),
    .A(_2347_),
    .Y(_2358_));
 sg13g2_a21oi_1 _4381_ (.A1(_2330_),
    .A2(_2345_),
    .Y(_2359_),
    .B1(_2358_));
 sg13g2_a21oi_1 _4382_ (.A1(_2343_),
    .A2(_2351_),
    .Y(_2360_),
    .B1(_2352_));
 sg13g2_inv_1 _4383_ (.Y(_2361_),
    .A(_2360_));
 sg13g2_nand2b_1 _4384_ (.Y(_2362_),
    .B(_2360_),
    .A_N(_2359_));
 sg13g2_nand2_1 _4385_ (.Y(_2363_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[8] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[8] ));
 sg13g2_xnor2_1 _4386_ (.Y(_2364_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[8] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[8] ));
 sg13g2_or2_1 _4387_ (.X(_2365_),
    .B(_2364_),
    .A(_2362_));
 sg13g2_nor2b_1 _4388_ (.A(net858),
    .B_N(\u_ddc_top_level.cic_right_inst.int_reg0[8] ),
    .Y(_2366_));
 sg13g2_a21oi_1 _4389_ (.A1(_2362_),
    .A2(_2364_),
    .Y(_2367_),
    .B1(net817));
 sg13g2_a21o_1 _4390_ (.A2(_2367_),
    .A1(_2365_),
    .B1(_2366_),
    .X(_0526_));
 sg13g2_nor2_1 _4391_ (.A(\u_ddc_top_level.cic_right_inst.comb_out2[9] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[9] ),
    .Y(_2368_));
 sg13g2_xor2_1 _4392_ (.B(\u_ddc_top_level.cic_right_inst.int_reg0[9] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[9] ),
    .X(_2369_));
 sg13g2_nand2_1 _4393_ (.Y(_2370_),
    .A(_2363_),
    .B(_2365_));
 sg13g2_xnor2_1 _4394_ (.Y(_2371_),
    .A(_2369_),
    .B(_2370_));
 sg13g2_nor2_1 _4395_ (.A(net858),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[9] ),
    .Y(_2372_));
 sg13g2_a21oi_1 _4396_ (.A1(net858),
    .A2(_2371_),
    .Y(_0527_),
    .B1(_2372_));
 sg13g2_and2_1 _4397_ (.A(\u_ddc_top_level.cic_right_inst.comb_out2[10] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[10] ),
    .X(_2373_));
 sg13g2_xnor2_1 _4398_ (.Y(_2374_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[10] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[10] ));
 sg13g2_a22oi_1 _4399_ (.Y(_2375_),
    .B1(\u_ddc_top_level.cic_right_inst.int_reg0[9] ),
    .B2(\u_ddc_top_level.cic_right_inst.comb_out2[9] ),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg0[8] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out2[8] ));
 sg13g2_and2_1 _4400_ (.A(_2365_),
    .B(_2375_),
    .X(_2376_));
 sg13g2_nor3_1 _4401_ (.A(_2368_),
    .B(_2374_),
    .C(_2376_),
    .Y(_2377_));
 sg13g2_o21ai_1 _4402_ (.B1(_2374_),
    .Y(_2378_),
    .A1(_2368_),
    .A2(_2376_));
 sg13g2_nand2_1 _4403_ (.Y(_2379_),
    .A(net817),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[10] ));
 sg13g2_nand2_1 _4404_ (.Y(_2380_),
    .A(net860),
    .B(_2378_));
 sg13g2_o21ai_1 _4405_ (.B1(_2379_),
    .Y(_0528_),
    .A1(_2377_),
    .A2(_2380_));
 sg13g2_nor2_1 _4406_ (.A(net858),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[11] ),
    .Y(_2381_));
 sg13g2_nand2_1 _4407_ (.Y(_2382_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[11] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[11] ));
 sg13g2_xnor2_1 _4408_ (.Y(_2383_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[11] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[11] ));
 sg13g2_nor2_1 _4409_ (.A(_2373_),
    .B(_2377_),
    .Y(_2384_));
 sg13g2_xnor2_1 _4410_ (.Y(_2385_),
    .A(_2383_),
    .B(_2384_));
 sg13g2_a21oi_1 _4411_ (.A1(net858),
    .A2(_2385_),
    .Y(_0529_),
    .B1(_2381_));
 sg13g2_nor2_1 _4412_ (.A(net858),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[12] ),
    .Y(_2386_));
 sg13g2_nor2_1 _4413_ (.A(_2374_),
    .B(_2383_),
    .Y(_2387_));
 sg13g2_nand2_1 _4414_ (.Y(_2388_),
    .A(_2369_),
    .B(_2387_));
 sg13g2_nor4_2 _4415_ (.A(_2359_),
    .B(_2361_),
    .C(_2364_),
    .Y(_2389_),
    .D(_2388_));
 sg13g2_o21ai_1 _4416_ (.B1(_2373_),
    .Y(_2390_),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out2[11] ),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg0[11] ));
 sg13g2_or4_1 _4417_ (.A(_2368_),
    .B(_2374_),
    .C(_2375_),
    .D(_2383_),
    .X(_2391_));
 sg13g2_nand3_1 _4418_ (.B(_2390_),
    .C(_2391_),
    .A(_2382_),
    .Y(_2392_));
 sg13g2_nor2_2 _4419_ (.A(_2389_),
    .B(_2392_),
    .Y(_2393_));
 sg13g2_nand2_1 _4420_ (.Y(_2394_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[12] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[12] ));
 sg13g2_xnor2_1 _4421_ (.Y(_2395_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[12] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[12] ));
 sg13g2_xnor2_1 _4422_ (.Y(_2396_),
    .A(_2393_),
    .B(_2395_));
 sg13g2_a21oi_1 _4423_ (.A1(net858),
    .A2(_2396_),
    .Y(_0530_),
    .B1(_2386_));
 sg13g2_nor2_1 _4424_ (.A(\u_ddc_top_level.cic_right_inst.comb_out2[13] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[13] ),
    .Y(_2397_));
 sg13g2_xor2_1 _4425_ (.B(\u_ddc_top_level.cic_right_inst.int_reg0[13] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[13] ),
    .X(_2398_));
 sg13g2_o21ai_1 _4426_ (.B1(_2394_),
    .Y(_2399_),
    .A1(_2393_),
    .A2(_2395_));
 sg13g2_xor2_1 _4427_ (.B(_2399_),
    .A(_2398_),
    .X(_2400_));
 sg13g2_mux2_1 _4428_ (.A0(\u_ddc_top_level.cic_right_inst.int_reg0[13] ),
    .A1(_2400_),
    .S(net860),
    .X(_0531_));
 sg13g2_nor2_1 _4429_ (.A(net861),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[14] ),
    .Y(_2401_));
 sg13g2_nand2_1 _4430_ (.Y(_2402_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[14] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[14] ));
 sg13g2_xnor2_1 _4431_ (.Y(_2403_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[14] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[14] ));
 sg13g2_a22oi_1 _4432_ (.Y(_2404_),
    .B1(\u_ddc_top_level.cic_right_inst.int_reg0[13] ),
    .B2(\u_ddc_top_level.cic_right_inst.comb_out2[13] ),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg0[12] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out2[12] ));
 sg13g2_nor2_1 _4433_ (.A(_2397_),
    .B(_2404_),
    .Y(_2405_));
 sg13g2_nand2b_1 _4434_ (.Y(_2406_),
    .B(_2398_),
    .A_N(_2395_));
 sg13g2_nor2_1 _4435_ (.A(_2393_),
    .B(_2406_),
    .Y(_2407_));
 sg13g2_nor2_1 _4436_ (.A(_2405_),
    .B(_2407_),
    .Y(_2408_));
 sg13g2_xnor2_1 _4437_ (.Y(_2409_),
    .A(_2403_),
    .B(_2408_));
 sg13g2_a21oi_1 _4438_ (.A1(net862),
    .A2(_2409_),
    .Y(_0532_),
    .B1(_2401_));
 sg13g2_nor2_1 _4439_ (.A(net861),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[15] ),
    .Y(_2410_));
 sg13g2_nor2_1 _4440_ (.A(\u_ddc_top_level.cic_right_inst.comb_out2[15] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[15] ),
    .Y(_2411_));
 sg13g2_xor2_1 _4441_ (.B(\u_ddc_top_level.cic_right_inst.int_reg0[15] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[15] ),
    .X(_2412_));
 sg13g2_o21ai_1 _4442_ (.B1(_2402_),
    .Y(_2413_),
    .A1(_2403_),
    .A2(_2408_));
 sg13g2_xnor2_1 _4443_ (.Y(_2414_),
    .A(_2412_),
    .B(_2413_));
 sg13g2_a21oi_1 _4444_ (.A1(net862),
    .A2(_2414_),
    .Y(_0533_),
    .B1(_2410_));
 sg13g2_nor2b_1 _4445_ (.A(_2403_),
    .B_N(_2412_),
    .Y(_2415_));
 sg13g2_nor2b_1 _4446_ (.A(_2406_),
    .B_N(_2415_),
    .Y(_2416_));
 sg13g2_o21ai_1 _4447_ (.B1(_2416_),
    .Y(_2417_),
    .A1(_2389_),
    .A2(_2392_));
 sg13g2_nor2_1 _4448_ (.A(_2402_),
    .B(_2411_),
    .Y(_2418_));
 sg13g2_a221oi_1 _4449_ (.B2(_2415_),
    .C1(_2418_),
    .B1(_2405_),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out2[15] ),
    .Y(_2419_),
    .A2(\u_ddc_top_level.cic_right_inst.int_reg0[15] ));
 sg13g2_nand2_1 _4450_ (.Y(_2420_),
    .A(_2417_),
    .B(_2419_));
 sg13g2_nand2_1 _4451_ (.Y(_2421_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[16] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[16] ));
 sg13g2_xor2_1 _4452_ (.B(\u_ddc_top_level.cic_right_inst.int_reg0[16] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[16] ),
    .X(_2422_));
 sg13g2_nand2_1 _4453_ (.Y(_2423_),
    .A(_2420_),
    .B(_2422_));
 sg13g2_o21ai_1 _4454_ (.B1(net859),
    .Y(_2424_),
    .A1(_2420_),
    .A2(_2422_));
 sg13g2_nor2b_1 _4455_ (.A(_2424_),
    .B_N(_2423_),
    .Y(_2425_));
 sg13g2_a21o_1 _4456_ (.A2(\u_ddc_top_level.cic_right_inst.int_reg0[16] ),
    .A1(net817),
    .B1(_2425_),
    .X(_0534_));
 sg13g2_nand2_1 _4457_ (.Y(_2426_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[17] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[17] ));
 sg13g2_nor2_1 _4458_ (.A(\u_ddc_top_level.cic_right_inst.comb_out2[17] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[17] ),
    .Y(_2427_));
 sg13g2_xnor2_1 _4459_ (.Y(_2428_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[17] ),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[17] ));
 sg13g2_and2_1 _4460_ (.A(_2421_),
    .B(_2423_),
    .X(_2429_));
 sg13g2_xnor2_1 _4461_ (.Y(_2430_),
    .A(_2428_),
    .B(_2429_));
 sg13g2_nor2_1 _4462_ (.A(net859),
    .B(\u_ddc_top_level.cic_right_inst.int_reg0[17] ),
    .Y(_2431_));
 sg13g2_a21oi_1 _4463_ (.A1(net859),
    .A2(_2430_),
    .Y(_0535_),
    .B1(_2431_));
 sg13g2_xor2_1 _4464_ (.B(\u_ddc_top_level.cic_right_inst.int_reg0[18] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[18] ),
    .X(_2432_));
 sg13g2_nand3b_1 _4465_ (.B(_2422_),
    .C(_2426_),
    .Y(_2433_),
    .A_N(_2427_));
 sg13g2_a21oi_1 _4466_ (.A1(_2417_),
    .A2(_2419_),
    .Y(_2434_),
    .B1(_2433_));
 sg13g2_o21ai_1 _4467_ (.B1(_2426_),
    .Y(_2435_),
    .A1(_2421_),
    .A2(_2427_));
 sg13g2_o21ai_1 _4468_ (.B1(_2432_),
    .Y(_2436_),
    .A1(_2434_),
    .A2(_2435_));
 sg13g2_or3_1 _4469_ (.A(_2432_),
    .B(_2434_),
    .C(_2435_),
    .X(_2437_));
 sg13g2_nand3_1 _4470_ (.B(_2436_),
    .C(_2437_),
    .A(net859),
    .Y(_2438_));
 sg13g2_o21ai_1 _4471_ (.B1(_2438_),
    .Y(_0536_),
    .A1(net859),
    .A2(_0744_));
 sg13g2_o21ai_1 _4472_ (.B1(_2436_),
    .Y(_2439_),
    .A1(_0740_),
    .A2(_0744_));
 sg13g2_xor2_1 _4473_ (.B(net882),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[18] ),
    .X(_2440_));
 sg13g2_xnor2_1 _4474_ (.Y(_2441_),
    .A(_2439_),
    .B(_2440_));
 sg13g2_nor2_1 _4475_ (.A(net858),
    .B(net882),
    .Y(_2442_));
 sg13g2_a21oi_1 _4476_ (.A1(net859),
    .A2(_2441_),
    .Y(_0537_),
    .B1(_2442_));
 sg13g2_nand2_1 _4477_ (.Y(_2443_),
    .A(net831),
    .B(\u_ddc_top_level.cic_left_inst.comb_out2[0] ));
 sg13g2_xnor2_1 _4478_ (.Y(_0626_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg0[0] ),
    .B(_2443_));
 sg13g2_and2_1 _4479_ (.A(\u_ddc_top_level.cic_left_inst.comb_out2[0] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[0] ),
    .X(_2444_));
 sg13g2_and2_1 _4480_ (.A(\u_ddc_top_level.cic_left_inst.comb_out2[1] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[1] ),
    .X(_2445_));
 sg13g2_xor2_1 _4481_ (.B(\u_ddc_top_level.cic_left_inst.int_reg0[1] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[1] ),
    .X(_2446_));
 sg13g2_nor2_1 _4482_ (.A(net831),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[1] ),
    .Y(_2447_));
 sg13g2_xnor2_1 _4483_ (.Y(_2448_),
    .A(_2444_),
    .B(_2446_));
 sg13g2_a21oi_1 _4484_ (.A1(net831),
    .A2(_2448_),
    .Y(_0627_),
    .B1(_2447_));
 sg13g2_nand2_1 _4485_ (.Y(_2449_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[2] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[2] ));
 sg13g2_xnor2_1 _4486_ (.Y(_2450_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[2] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[2] ));
 sg13g2_a21oi_1 _4487_ (.A1(_2444_),
    .A2(_2446_),
    .Y(_2451_),
    .B1(_2445_));
 sg13g2_xnor2_1 _4488_ (.Y(_2452_),
    .A(_2450_),
    .B(_2451_));
 sg13g2_nor2_1 _4489_ (.A(net832),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[2] ),
    .Y(_2453_));
 sg13g2_a21oi_1 _4490_ (.A1(net832),
    .A2(_2452_),
    .Y(_0628_),
    .B1(_2453_));
 sg13g2_and2_1 _4491_ (.A(\u_ddc_top_level.cic_left_inst.comb_out2[3] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[3] ),
    .X(_2454_));
 sg13g2_or2_1 _4492_ (.X(_2455_),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[3] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[3] ));
 sg13g2_nand2b_1 _4493_ (.Y(_2456_),
    .B(_2455_),
    .A_N(_2454_));
 sg13g2_o21ai_1 _4494_ (.B1(_2449_),
    .Y(_2457_),
    .A1(_2450_),
    .A2(_2451_));
 sg13g2_xnor2_1 _4495_ (.Y(_2458_),
    .A(_2456_),
    .B(_2457_));
 sg13g2_mux2_1 _4496_ (.A0(\u_ddc_top_level.cic_left_inst.int_reg0[3] ),
    .A1(_2458_),
    .S(net835),
    .X(_0629_));
 sg13g2_a21oi_2 _4497_ (.B1(_2454_),
    .Y(_2459_),
    .A2(_2457_),
    .A1(_2455_));
 sg13g2_nand2_1 _4498_ (.Y(_2460_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[4] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[4] ));
 sg13g2_xnor2_1 _4499_ (.Y(_2461_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[4] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[4] ));
 sg13g2_xnor2_1 _4500_ (.Y(_2462_),
    .A(_2459_),
    .B(_2461_));
 sg13g2_nor2_1 _4501_ (.A(net835),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[4] ),
    .Y(_2463_));
 sg13g2_a21oi_1 _4502_ (.A1(net835),
    .A2(_2462_),
    .Y(_0630_),
    .B1(_2463_));
 sg13g2_nor2_1 _4503_ (.A(\u_ddc_top_level.cic_left_inst.comb_out2[5] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[5] ),
    .Y(_2464_));
 sg13g2_nand2_1 _4504_ (.Y(_2465_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[5] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[5] ));
 sg13g2_nand2b_1 _4505_ (.Y(_2466_),
    .B(_2465_),
    .A_N(_2464_));
 sg13g2_o21ai_1 _4506_ (.B1(_2460_),
    .Y(_2467_),
    .A1(_2459_),
    .A2(_2461_));
 sg13g2_xnor2_1 _4507_ (.Y(_2468_),
    .A(_2466_),
    .B(_2467_));
 sg13g2_mux2_1 _4508_ (.A0(\u_ddc_top_level.cic_left_inst.int_reg0[5] ),
    .A1(_2468_),
    .S(net835),
    .X(_0631_));
 sg13g2_nor2_1 _4509_ (.A(net836),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[6] ),
    .Y(_2469_));
 sg13g2_nand2_1 _4510_ (.Y(_2470_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[6] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[6] ));
 sg13g2_inv_1 _4511_ (.Y(_2471_),
    .A(_2470_));
 sg13g2_nor2_1 _4512_ (.A(\u_ddc_top_level.cic_left_inst.comb_out2[6] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[6] ),
    .Y(_2472_));
 sg13g2_or2_1 _4513_ (.X(_2473_),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[6] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[6] ));
 sg13g2_nand2_1 _4514_ (.Y(_2474_),
    .A(_2470_),
    .B(_2473_));
 sg13g2_or2_1 _4515_ (.X(_2475_),
    .B(_2466_),
    .A(_2461_));
 sg13g2_nor2_1 _4516_ (.A(_2459_),
    .B(_2475_),
    .Y(_2476_));
 sg13g2_o21ai_1 _4517_ (.B1(_2465_),
    .Y(_2477_),
    .A1(_2460_),
    .A2(_2464_));
 sg13g2_or2_1 _4518_ (.X(_2478_),
    .B(_2477_),
    .A(_2476_));
 sg13g2_xor2_1 _4519_ (.B(_2478_),
    .A(_2474_),
    .X(_2479_));
 sg13g2_a21oi_1 _4520_ (.A1(net836),
    .A2(_2479_),
    .Y(_0632_),
    .B1(_2469_));
 sg13g2_nor2_1 _4521_ (.A(net836),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[7] ),
    .Y(_2480_));
 sg13g2_nor2_1 _4522_ (.A(\u_ddc_top_level.cic_left_inst.comb_out2[7] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[7] ),
    .Y(_2481_));
 sg13g2_nand2_1 _4523_ (.Y(_2482_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[7] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[7] ));
 sg13g2_nand2b_1 _4524_ (.Y(_2483_),
    .B(_2482_),
    .A_N(_2481_));
 sg13g2_a21oi_1 _4525_ (.A1(_2473_),
    .A2(_2478_),
    .Y(_2484_),
    .B1(_2471_));
 sg13g2_xnor2_1 _4526_ (.Y(_2485_),
    .A(_2483_),
    .B(_2484_));
 sg13g2_a21oi_1 _4527_ (.A1(net836),
    .A2(_2485_),
    .Y(_0633_),
    .B1(_2480_));
 sg13g2_nand2_1 _4528_ (.Y(_2486_),
    .A(net811),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[8] ));
 sg13g2_o21ai_1 _4529_ (.B1(_2482_),
    .Y(_2487_),
    .A1(_2470_),
    .A2(_2481_));
 sg13g2_nor2_1 _4530_ (.A(_2477_),
    .B(_2487_),
    .Y(_2488_));
 sg13g2_o21ai_1 _4531_ (.B1(_2488_),
    .Y(_2489_),
    .A1(_2459_),
    .A2(_2475_));
 sg13g2_a21oi_1 _4532_ (.A1(_2472_),
    .A2(_2482_),
    .Y(_2490_),
    .B1(_2481_));
 sg13g2_nand2_1 _4533_ (.Y(_2491_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[8] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[8] ));
 sg13g2_xor2_1 _4534_ (.B(\u_ddc_top_level.cic_left_inst.int_reg0[8] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[8] ),
    .X(_2492_));
 sg13g2_nand3_1 _4535_ (.B(_2490_),
    .C(_2492_),
    .A(_2489_),
    .Y(_2493_));
 sg13g2_a21oi_1 _4536_ (.A1(_2489_),
    .A2(_2490_),
    .Y(_2494_),
    .B1(_2492_));
 sg13g2_nand2_1 _4537_ (.Y(_2495_),
    .A(net844),
    .B(_2493_));
 sg13g2_o21ai_1 _4538_ (.B1(_2486_),
    .Y(_0634_),
    .A1(_2494_),
    .A2(_2495_));
 sg13g2_nor2_1 _4539_ (.A(\u_ddc_top_level.cic_left_inst.comb_out2[9] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[9] ),
    .Y(_2496_));
 sg13g2_xor2_1 _4540_ (.B(\u_ddc_top_level.cic_left_inst.int_reg0[9] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[9] ),
    .X(_2497_));
 sg13g2_and2_1 _4541_ (.A(_2491_),
    .B(_2493_),
    .X(_2498_));
 sg13g2_xor2_1 _4542_ (.B(_2498_),
    .A(_2497_),
    .X(_2499_));
 sg13g2_nor2_1 _4543_ (.A(net844),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[9] ),
    .Y(_2500_));
 sg13g2_a21oi_1 _4544_ (.A1(net844),
    .A2(_2499_),
    .Y(_0635_),
    .B1(_2500_));
 sg13g2_nor2_1 _4545_ (.A(net845),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[10] ),
    .Y(_2501_));
 sg13g2_nand2_1 _4546_ (.Y(_2502_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[10] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[10] ));
 sg13g2_xor2_1 _4547_ (.B(\u_ddc_top_level.cic_left_inst.int_reg0[10] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[10] ),
    .X(_2503_));
 sg13g2_inv_1 _4548_ (.Y(_2504_),
    .A(_2503_));
 sg13g2_a22oi_1 _4549_ (.Y(_2505_),
    .B1(\u_ddc_top_level.cic_left_inst.int_reg0[9] ),
    .B2(\u_ddc_top_level.cic_left_inst.comb_out2[9] ),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg0[8] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out2[8] ));
 sg13g2_a21oi_1 _4550_ (.A1(_2493_),
    .A2(_2505_),
    .Y(_2506_),
    .B1(_2496_));
 sg13g2_nand2_1 _4551_ (.Y(_2507_),
    .A(_2503_),
    .B(_2506_));
 sg13g2_xnor2_1 _4552_ (.Y(_2508_),
    .A(_2503_),
    .B(_2506_));
 sg13g2_a21oi_1 _4553_ (.A1(net845),
    .A2(_2508_),
    .Y(_0636_),
    .B1(_2501_));
 sg13g2_nor2_1 _4554_ (.A(net845),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[11] ),
    .Y(_2509_));
 sg13g2_nor2_1 _4555_ (.A(\u_ddc_top_level.cic_left_inst.comb_out2[11] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[11] ),
    .Y(_2510_));
 sg13g2_xnor2_1 _4556_ (.Y(_2511_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[11] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[11] ));
 sg13g2_nand2_1 _4557_ (.Y(_2512_),
    .A(_2502_),
    .B(_2507_));
 sg13g2_xor2_1 _4558_ (.B(_2512_),
    .A(_2511_),
    .X(_2513_));
 sg13g2_a21oi_1 _4559_ (.A1(net845),
    .A2(_2513_),
    .Y(_0637_),
    .B1(_2509_));
 sg13g2_nor2_1 _4560_ (.A(_2504_),
    .B(_2511_),
    .Y(_2514_));
 sg13g2_nand2_1 _4561_ (.Y(_2515_),
    .A(_2497_),
    .B(_2514_));
 sg13g2_nor2_1 _4562_ (.A(_2496_),
    .B(_2505_),
    .Y(_2516_));
 sg13g2_nor2_1 _4563_ (.A(_2502_),
    .B(_2510_),
    .Y(_2517_));
 sg13g2_a221oi_1 _4564_ (.B2(_2516_),
    .C1(_2517_),
    .B1(_2514_),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out2[11] ),
    .Y(_2518_),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg0[11] ));
 sg13g2_o21ai_1 _4565_ (.B1(_2518_),
    .Y(_2519_),
    .A1(_2493_),
    .A2(_2515_));
 sg13g2_nand2_1 _4566_ (.Y(_2520_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[12] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[12] ));
 sg13g2_xor2_1 _4567_ (.B(\u_ddc_top_level.cic_left_inst.int_reg0[12] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[12] ),
    .X(_2521_));
 sg13g2_nand2_1 _4568_ (.Y(_2522_),
    .A(_2519_),
    .B(_2521_));
 sg13g2_o21ai_1 _4569_ (.B1(net848),
    .Y(_2523_),
    .A1(_2519_),
    .A2(_2521_));
 sg13g2_nor2b_1 _4570_ (.A(_2523_),
    .B_N(_2522_),
    .Y(_2524_));
 sg13g2_a21o_1 _4571_ (.A2(\u_ddc_top_level.cic_left_inst.int_reg0[12] ),
    .A1(net811),
    .B1(_2524_),
    .X(_0638_));
 sg13g2_nor2_1 _4572_ (.A(\u_ddc_top_level.cic_left_inst.comb_out2[13] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[13] ),
    .Y(_2525_));
 sg13g2_xor2_1 _4573_ (.B(\u_ddc_top_level.cic_left_inst.int_reg0[13] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[13] ),
    .X(_2526_));
 sg13g2_nand2_1 _4574_ (.Y(_2527_),
    .A(_2520_),
    .B(_2522_));
 sg13g2_xor2_1 _4575_ (.B(_2527_),
    .A(_2526_),
    .X(_2528_));
 sg13g2_mux2_1 _4576_ (.A0(\u_ddc_top_level.cic_left_inst.int_reg0[13] ),
    .A1(_2528_),
    .S(net848),
    .X(_0639_));
 sg13g2_and2_1 _4577_ (.A(\u_ddc_top_level.cic_left_inst.comb_out2[14] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[14] ),
    .X(_2529_));
 sg13g2_xor2_1 _4578_ (.B(\u_ddc_top_level.cic_left_inst.int_reg0[14] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[14] ),
    .X(_2530_));
 sg13g2_a22oi_1 _4579_ (.Y(_2531_),
    .B1(\u_ddc_top_level.cic_left_inst.int_reg0[13] ),
    .B2(\u_ddc_top_level.cic_left_inst.comb_out2[13] ),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg0[12] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out2[12] ));
 sg13g2_nor2_1 _4580_ (.A(_2525_),
    .B(_2531_),
    .Y(_2532_));
 sg13g2_a21oi_2 _4581_ (.B1(_2525_),
    .Y(_2533_),
    .A2(_2531_),
    .A1(_2522_));
 sg13g2_o21ai_1 _4582_ (.B1(net848),
    .Y(_2534_),
    .A1(_2530_),
    .A2(_2533_));
 sg13g2_a21oi_1 _4583_ (.A1(_2530_),
    .A2(_2533_),
    .Y(_2535_),
    .B1(_2534_));
 sg13g2_a21o_1 _4584_ (.A2(\u_ddc_top_level.cic_left_inst.int_reg0[14] ),
    .A1(net810),
    .B1(_2535_),
    .X(_0640_));
 sg13g2_nor2_1 _4585_ (.A(net848),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[15] ),
    .Y(_2536_));
 sg13g2_nand2_1 _4586_ (.Y(_2537_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[15] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[15] ));
 sg13g2_xor2_1 _4587_ (.B(\u_ddc_top_level.cic_left_inst.int_reg0[15] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[15] ),
    .X(_2538_));
 sg13g2_a21oi_1 _4588_ (.A1(_2530_),
    .A2(_2533_),
    .Y(_2539_),
    .B1(_2529_));
 sg13g2_xor2_1 _4589_ (.B(_2539_),
    .A(_2538_),
    .X(_2540_));
 sg13g2_a21oi_1 _4590_ (.A1(net848),
    .A2(_2540_),
    .Y(_0641_),
    .B1(_2536_));
 sg13g2_and4_1 _4591_ (.A(_2521_),
    .B(_2526_),
    .C(_2530_),
    .D(_2538_),
    .X(_2541_));
 sg13g2_nand3_1 _4592_ (.B(_2532_),
    .C(_2538_),
    .A(_2530_),
    .Y(_2542_));
 sg13g2_o21ai_1 _4593_ (.B1(_2529_),
    .Y(_2543_),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out2[15] ),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg0[15] ));
 sg13g2_nand3_1 _4594_ (.B(_2542_),
    .C(_2543_),
    .A(_2537_),
    .Y(_2544_));
 sg13g2_a21o_1 _4595_ (.A2(_2541_),
    .A1(_2519_),
    .B1(_2544_),
    .X(_2545_));
 sg13g2_nand2_1 _4596_ (.Y(_2546_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[16] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[16] ));
 sg13g2_xor2_1 _4597_ (.B(\u_ddc_top_level.cic_left_inst.int_reg0[16] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[16] ),
    .X(_2547_));
 sg13g2_nand2_1 _4598_ (.Y(_2548_),
    .A(_2545_),
    .B(_2547_));
 sg13g2_o21ai_1 _4599_ (.B1(net849),
    .Y(_2549_),
    .A1(_2545_),
    .A2(_2547_));
 sg13g2_nor2b_1 _4600_ (.A(_2549_),
    .B_N(_2548_),
    .Y(_2550_));
 sg13g2_a21o_1 _4601_ (.A2(\u_ddc_top_level.cic_left_inst.int_reg0[16] ),
    .A1(net810),
    .B1(_2550_),
    .X(_0642_));
 sg13g2_nor2_1 _4602_ (.A(net849),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[17] ),
    .Y(_2551_));
 sg13g2_xor2_1 _4603_ (.B(\u_ddc_top_level.cic_left_inst.int_reg0[17] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[17] ),
    .X(_2552_));
 sg13g2_nand2_1 _4604_ (.Y(_2553_),
    .A(_2546_),
    .B(_2548_));
 sg13g2_xnor2_1 _4605_ (.Y(_2554_),
    .A(_2552_),
    .B(_2553_));
 sg13g2_a21oi_1 _4606_ (.A1(net849),
    .A2(_2554_),
    .Y(_0643_),
    .B1(_2551_));
 sg13g2_nor2_1 _4607_ (.A(net849),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[18] ),
    .Y(_2555_));
 sg13g2_nand2_1 _4608_ (.Y(_2556_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[18] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[18] ));
 sg13g2_nor2_1 _4609_ (.A(\u_ddc_top_level.cic_left_inst.comb_out2[18] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[18] ),
    .Y(_2557_));
 sg13g2_xnor2_1 _4610_ (.Y(_2558_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[18] ),
    .B(\u_ddc_top_level.cic_left_inst.int_reg0[18] ));
 sg13g2_and2_1 _4611_ (.A(_2547_),
    .B(_2552_),
    .X(_2559_));
 sg13g2_a21oi_1 _4612_ (.A1(_0730_),
    .A2(_0745_),
    .Y(_2560_),
    .B1(_2546_));
 sg13g2_a221oi_1 _4613_ (.B2(_2559_),
    .C1(_2560_),
    .B1(_2545_),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out2[17] ),
    .Y(_2561_),
    .A2(\u_ddc_top_level.cic_left_inst.int_reg0[17] ));
 sg13g2_xnor2_1 _4614_ (.Y(_2562_),
    .A(_2558_),
    .B(_2561_));
 sg13g2_a21oi_1 _4615_ (.A1(net849),
    .A2(_2562_),
    .Y(_0644_),
    .B1(_2555_));
 sg13g2_o21ai_1 _4616_ (.B1(_2556_),
    .Y(_2563_),
    .A1(_2557_),
    .A2(_2561_));
 sg13g2_xor2_1 _4617_ (.B(net879),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[18] ),
    .X(_2564_));
 sg13g2_xnor2_1 _4618_ (.Y(_2565_),
    .A(_2563_),
    .B(_2564_));
 sg13g2_nor2_1 _4619_ (.A(net847),
    .B(net880),
    .Y(_2566_));
 sg13g2_a21oi_1 _4620_ (.A1(net847),
    .A2(_2565_),
    .Y(_0645_),
    .B1(_2566_));
 sg13g2_mux2_1 _4621_ (.A0(net820),
    .A1(net876),
    .S(net823),
    .X(_0681_));
 sg13g2_mux2_1 _4622_ (.A0(\u_ddc_top_level.cic_left_inst.in_data[0] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[0] ),
    .S(net821),
    .X(_0682_));
 sg13g2_mux2_1 _4623_ (.A0(\u_ddc_top_level.cic_left_inst.in_data[1] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[1] ),
    .S(net821),
    .X(_0683_));
 sg13g2_mux2_1 _4624_ (.A0(\u_ddc_top_level.cic_left_inst.in_data[2] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[2] ),
    .S(net821),
    .X(_0684_));
 sg13g2_mux2_1 _4625_ (.A0(\u_ddc_top_level.cic_left_inst.in_data[3] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[3] ),
    .S(net821),
    .X(_0685_));
 sg13g2_mux2_1 _4626_ (.A0(\u_ddc_top_level.cic_left_inst.in_data[4] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[4] ),
    .S(net821),
    .X(_0686_));
 sg13g2_mux2_1 _4627_ (.A0(\u_ddc_top_level.cic_left_inst.in_data[5] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[5] ),
    .S(net821),
    .X(_0687_));
 sg13g2_mux2_1 _4628_ (.A0(\u_ddc_top_level.cic_left_inst.in_data[6] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[6] ),
    .S(net823),
    .X(_0688_));
 sg13g2_mux2_1 _4629_ (.A0(\u_ddc_top_level.cic_left_inst.in_data[7] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[7] ),
    .S(net821),
    .X(_0689_));
 sg13g2_mux2_1 _4630_ (.A0(\u_ddc_top_level.cic_left_inst.in_data[8] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[8] ),
    .S(net823),
    .X(_0690_));
 sg13g2_mux2_1 _4631_ (.A0(\u_ddc_top_level.cic_left_inst.in_data[9] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[9] ),
    .S(net823),
    .X(_0691_));
 sg13g2_nand2_1 _4632_ (.Y(_2567_),
    .A(\u_ddc_top_level.i2s_rx_inst.shift_reg[10] ),
    .B(net822));
 sg13g2_o21ai_1 _4633_ (.B1(_2567_),
    .Y(_0692_),
    .A1(_0728_),
    .A2(net822));
 sg13g2_mux2_1 _4634_ (.A0(\u_ddc_top_level.cic_left_inst.in_data[11] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[11] ),
    .S(net822),
    .X(_0693_));
 sg13g2_mux2_1 _4635_ (.A0(\u_ddc_top_level.cic_left_inst.in_data[12] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[12] ),
    .S(net822),
    .X(_0694_));
 sg13g2_mux2_1 _4636_ (.A0(\u_ddc_top_level.cic_left_inst.in_data[13] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[13] ),
    .S(net822),
    .X(_0695_));
 sg13g2_mux2_1 _4637_ (.A0(\u_ddc_top_level.cic_left_inst.in_data[14] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[14] ),
    .S(net822),
    .X(_0696_));
 sg13g2_mux2_1 _4638_ (.A0(\u_ddc_top_level.cic_left_inst.in_data[15] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[15] ),
    .S(net822),
    .X(_0697_));
 sg13g2_mux2_1 _4639_ (.A0(\u_ddc_top_level.cic_right_inst.in_data[0] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[0] ),
    .S(net818),
    .X(_0698_));
 sg13g2_mux2_1 _4640_ (.A0(\u_ddc_top_level.cic_right_inst.in_data[1] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[1] ),
    .S(net818),
    .X(_0699_));
 sg13g2_mux2_1 _4641_ (.A0(\u_ddc_top_level.cic_right_inst.in_data[2] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[2] ),
    .S(net818),
    .X(_0700_));
 sg13g2_mux2_1 _4642_ (.A0(\u_ddc_top_level.cic_right_inst.in_data[3] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[3] ),
    .S(net818),
    .X(_0701_));
 sg13g2_mux2_1 _4643_ (.A0(\u_ddc_top_level.cic_right_inst.in_data[4] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[4] ),
    .S(net818),
    .X(_0702_));
 sg13g2_mux2_1 _4644_ (.A0(\u_ddc_top_level.cic_right_inst.in_data[5] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[5] ),
    .S(net818),
    .X(_0703_));
 sg13g2_mux2_1 _4645_ (.A0(\u_ddc_top_level.cic_right_inst.in_data[6] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[6] ),
    .S(net818),
    .X(_0704_));
 sg13g2_mux2_1 _4646_ (.A0(\u_ddc_top_level.cic_right_inst.in_data[7] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[7] ),
    .S(net820),
    .X(_0705_));
 sg13g2_mux2_1 _4647_ (.A0(\u_ddc_top_level.cic_right_inst.in_data[8] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[8] ),
    .S(net820),
    .X(_0706_));
 sg13g2_mux2_1 _4648_ (.A0(\u_ddc_top_level.cic_right_inst.in_data[9] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[9] ),
    .S(net820),
    .X(_0707_));
 sg13g2_mux2_1 _4649_ (.A0(\u_ddc_top_level.cic_right_inst.in_data[10] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[10] ),
    .S(net819),
    .X(_0708_));
 sg13g2_mux2_1 _4650_ (.A0(\u_ddc_top_level.cic_right_inst.in_data[11] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[11] ),
    .S(net819),
    .X(_0709_));
 sg13g2_mux2_1 _4651_ (.A0(\u_ddc_top_level.cic_right_inst.in_data[12] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[12] ),
    .S(net819),
    .X(_0710_));
 sg13g2_nand2_1 _4652_ (.Y(_2568_),
    .A(\u_ddc_top_level.i2s_rx_inst.shift_reg[13] ),
    .B(net819));
 sg13g2_o21ai_1 _4653_ (.B1(_2568_),
    .Y(_0711_),
    .A1(_0739_),
    .A2(net819));
 sg13g2_mux2_1 _4654_ (.A0(\u_ddc_top_level.cic_right_inst.in_data[14] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[14] ),
    .S(net819),
    .X(_0712_));
 sg13g2_mux2_1 _4655_ (.A0(\u_ddc_top_level.cic_right_inst.in_data[15] ),
    .A1(\u_ddc_top_level.i2s_rx_inst.shift_reg[15] ),
    .S(net819),
    .X(_0713_));
 sg13g2_mux2_1 _4656_ (.A0(net821),
    .A1(net826),
    .S(net818),
    .X(_0714_));
 sg13g2_inv_1 _4657_ (.Y(_0189_),
    .A(net890));
 sg13g2_inv_1 _4658_ (.Y(_0190_),
    .A(net890));
 sg13g2_inv_1 _4659_ (.Y(_0191_),
    .A(net891));
 sg13g2_inv_1 _4660_ (.Y(_0192_),
    .A(net891));
 sg13g2_inv_1 _4661_ (.Y(_0193_),
    .A(net899));
 sg13g2_inv_1 _4662_ (.Y(_0194_),
    .A(net899));
 sg13g2_inv_1 _4663_ (.Y(_0195_),
    .A(net902));
 sg13g2_inv_1 _4664_ (.Y(_0196_),
    .A(net903));
 sg13g2_inv_1 _4665_ (.Y(_0197_),
    .A(net903));
 sg13g2_inv_1 _4666_ (.Y(_0198_),
    .A(net904));
 sg13g2_inv_1 _4667_ (.Y(_0199_),
    .A(net904));
 sg13g2_inv_1 _4668_ (.Y(_0200_),
    .A(net904));
 sg13g2_inv_1 _4669_ (.Y(_0201_),
    .A(net904));
 sg13g2_inv_1 _4670_ (.Y(_0202_),
    .A(net918));
 sg13g2_inv_1 _4671_ (.Y(_0203_),
    .A(net918));
 sg13g2_inv_1 _4672_ (.Y(_0204_),
    .A(net919));
 sg13g2_inv_1 _4673_ (.Y(_0205_),
    .A(net919));
 sg13g2_inv_1 _4674_ (.Y(_0206_),
    .A(net887));
 sg13g2_inv_1 _4675_ (.Y(_0207_),
    .A(net887));
 sg13g2_inv_1 _4676_ (.Y(_0208_),
    .A(net888));
 sg13g2_inv_1 _4677_ (.Y(_0209_),
    .A(net891));
 sg13g2_inv_1 _4678_ (.Y(_0210_),
    .A(net892));
 sg13g2_inv_1 _4679_ (.Y(_0211_),
    .A(net892));
 sg13g2_inv_1 _4680_ (.Y(_0212_),
    .A(net895));
 sg13g2_inv_1 _4681_ (.Y(_0213_),
    .A(net895));
 sg13g2_inv_1 _4682_ (.Y(_0214_),
    .A(net895));
 sg13g2_inv_1 _4683_ (.Y(_0215_),
    .A(net896));
 sg13g2_inv_1 _4684_ (.Y(_0216_),
    .A(net896));
 sg13g2_inv_1 _4685_ (.Y(_0217_),
    .A(net895));
 sg13g2_inv_1 _4686_ (.Y(_0218_),
    .A(net895));
 sg13g2_inv_1 _4687_ (.Y(_0219_),
    .A(net895));
 sg13g2_inv_1 _4688_ (.Y(_0220_),
    .A(net912));
 sg13g2_inv_1 _4689_ (.Y(_0221_),
    .A(net912));
 sg13g2_inv_1 _4690_ (.Y(_0222_),
    .A(net912));
 sg13g2_inv_1 _4691_ (.Y(_0223_),
    .A(net912));
 sg13g2_inv_1 _4692_ (.Y(_0224_),
    .A(net909));
 sg13g2_inv_1 _4693_ (.Y(_0225_),
    .A(net898));
 sg13g2_inv_1 _4694_ (.Y(_0226_),
    .A(net898));
 sg13g2_inv_1 _4695_ (.Y(_0227_),
    .A(net898));
 sg13g2_inv_1 _4696_ (.Y(_0228_),
    .A(net900));
 sg13g2_inv_1 _4697_ (.Y(_0229_),
    .A(net900));
 sg13g2_inv_1 _4698_ (.Y(_0230_),
    .A(net900));
 sg13g2_inv_1 _4699_ (.Y(_0231_),
    .A(net901));
 sg13g2_inv_1 _4700_ (.Y(_0232_),
    .A(net901));
 sg13g2_inv_1 _4701_ (.Y(_0233_),
    .A(net906));
 sg13g2_inv_1 _4702_ (.Y(_0234_),
    .A(net905));
 sg13g2_inv_1 _4703_ (.Y(_0235_),
    .A(net905));
 sg13g2_inv_1 _4704_ (.Y(_0236_),
    .A(net906));
 sg13g2_inv_1 _4705_ (.Y(_0237_),
    .A(net906));
 sg13g2_inv_1 _4706_ (.Y(_0238_),
    .A(net921));
 sg13g2_inv_1 _4707_ (.Y(_0239_),
    .A(net920));
 sg13g2_inv_1 _4708_ (.Y(_0240_),
    .A(net921));
 sg13g2_inv_1 _4709_ (.Y(_0241_),
    .A(net933));
 sg13g2_inv_1 _4710_ (.Y(_0242_),
    .A(net934));
 sg13g2_inv_1 _4711_ (.Y(_0243_),
    .A(net933));
 sg13g2_inv_1 _4712_ (.Y(_0244_),
    .A(net933));
 sg13g2_inv_1 _4713_ (.Y(_0245_),
    .A(net934));
 sg13g2_inv_1 _4714_ (.Y(_0246_),
    .A(net934));
 sg13g2_inv_1 _4715_ (.Y(_0247_),
    .A(net934));
 sg13g2_inv_1 _4716_ (.Y(_0248_),
    .A(net938));
 sg13g2_inv_1 _4717_ (.Y(_0249_),
    .A(net938));
 sg13g2_inv_1 _4718_ (.Y(_0250_),
    .A(net938));
 sg13g2_inv_1 _4719_ (.Y(_0251_),
    .A(net937));
 sg13g2_inv_1 _4720_ (.Y(_0252_),
    .A(net937));
 sg13g2_inv_1 _4721_ (.Y(_0253_),
    .A(net954));
 sg13g2_inv_1 _4722_ (.Y(_0254_),
    .A(net952));
 sg13g2_inv_1 _4723_ (.Y(_0255_),
    .A(net954));
 sg13g2_inv_1 _4724_ (.Y(_0256_),
    .A(net953));
 sg13g2_inv_1 _4725_ (.Y(_0257_),
    .A(net953));
 sg13g2_inv_1 _4726_ (.Y(_0258_),
    .A(net890));
 sg13g2_inv_1 _4727_ (.Y(_0259_),
    .A(net890));
 sg13g2_inv_1 _4728_ (.Y(_0260_),
    .A(net890));
 sg13g2_inv_1 _4729_ (.Y(_0261_),
    .A(net898));
 sg13g2_inv_1 _4730_ (.Y(_0262_),
    .A(net898));
 sg13g2_inv_1 _4731_ (.Y(_0263_),
    .A(net899));
 sg13g2_inv_1 _4732_ (.Y(_0264_),
    .A(net899));
 sg13g2_inv_1 _4733_ (.Y(_0265_),
    .A(net899));
 sg13g2_inv_1 _4734_ (.Y(_0266_),
    .A(net903));
 sg13g2_inv_1 _4735_ (.Y(_0267_),
    .A(net903));
 sg13g2_inv_1 _4736_ (.Y(_0268_),
    .A(net903));
 sg13g2_inv_1 _4737_ (.Y(_0269_),
    .A(net906));
 sg13g2_inv_1 _4738_ (.Y(_0270_),
    .A(net907));
 sg13g2_inv_1 _4739_ (.Y(_0271_),
    .A(net920));
 sg13g2_inv_1 _4740_ (.Y(_0272_),
    .A(net920));
 sg13g2_inv_1 _4741_ (.Y(_0273_),
    .A(net921));
 sg13g2_inv_1 _4742_ (.Y(_0274_),
    .A(net918));
 sg13g2_inv_1 _4743_ (.Y(_0275_),
    .A(net887));
 sg13g2_inv_1 _4744_ (.Y(_0276_),
    .A(net890));
 sg13g2_inv_1 _4745_ (.Y(_0277_),
    .A(net890));
 sg13g2_inv_1 _4746_ (.Y(_0278_),
    .A(net891));
 sg13g2_inv_1 _4747_ (.Y(_0279_),
    .A(net891));
 sg13g2_inv_1 _4748_ (.Y(_0280_),
    .A(net891));
 sg13g2_inv_1 _4749_ (.Y(_0281_),
    .A(net899));
 sg13g2_inv_1 _4750_ (.Y(_0282_),
    .A(net903));
 sg13g2_inv_1 _4751_ (.Y(_0283_),
    .A(net903));
 sg13g2_inv_1 _4752_ (.Y(_0284_),
    .A(net903));
 sg13g2_inv_1 _4753_ (.Y(_0285_),
    .A(net904));
 sg13g2_inv_1 _4754_ (.Y(_0286_),
    .A(net904));
 sg13g2_inv_1 _4755_ (.Y(_0287_),
    .A(net907));
 sg13g2_inv_1 _4756_ (.Y(_0288_),
    .A(net904));
 sg13g2_inv_1 _4757_ (.Y(_0289_),
    .A(net918));
 sg13g2_inv_1 _4758_ (.Y(_0290_),
    .A(net918));
 sg13g2_inv_1 _4759_ (.Y(_0291_),
    .A(net919));
 sg13g2_inv_1 _4760_ (.Y(_0292_),
    .A(net919));
 sg13g2_inv_1 _4761_ (.Y(_0293_),
    .A(net941));
 sg13g2_inv_1 _4762_ (.Y(_0294_),
    .A(net941));
 sg13g2_inv_1 _4763_ (.Y(_0295_),
    .A(net941));
 sg13g2_inv_1 _4764_ (.Y(_0296_),
    .A(net945));
 sg13g2_inv_1 _4765_ (.Y(_0297_),
    .A(net934));
 sg13g2_inv_1 _4766_ (.Y(_0298_),
    .A(net934));
 sg13g2_inv_1 _4767_ (.Y(_0299_),
    .A(net938));
 sg13g2_inv_1 _4768_ (.Y(_0300_),
    .A(net946));
 sg13g2_inv_1 _4769_ (.Y(_0301_),
    .A(net938));
 sg13g2_inv_1 _4770_ (.Y(_0302_),
    .A(net939));
 sg13g2_inv_1 _4771_ (.Y(_0303_),
    .A(net939));
 sg13g2_inv_1 _4772_ (.Y(_0304_),
    .A(net939));
 sg13g2_inv_1 _4773_ (.Y(_0305_),
    .A(net955));
 sg13g2_inv_1 _4774_ (.Y(_0306_),
    .A(net955));
 sg13g2_inv_1 _4775_ (.Y(_0307_),
    .A(net956));
 sg13g2_inv_1 _4776_ (.Y(_0308_),
    .A(net955));
 sg13g2_inv_1 _4777_ (.Y(_0309_),
    .A(net956));
 sg13g2_inv_1 _4778_ (.Y(_0310_),
    .A(net956));
 sg13g2_inv_1 _4779_ (.Y(_0311_),
    .A(net942));
 sg13g2_inv_1 _4780_ (.Y(_0312_),
    .A(net941));
 sg13g2_inv_1 _4781_ (.Y(_0313_),
    .A(net942));
 sg13g2_inv_1 _4782_ (.Y(_0314_),
    .A(net942));
 sg13g2_inv_1 _4783_ (.Y(_0315_),
    .A(net942));
 sg13g2_inv_1 _4784_ (.Y(_0316_),
    .A(net946));
 sg13g2_inv_1 _4785_ (.Y(_0317_),
    .A(net946));
 sg13g2_inv_1 _4786_ (.Y(_0318_),
    .A(net946));
 sg13g2_inv_1 _4787_ (.Y(_0319_),
    .A(net947));
 sg13g2_inv_1 _4788_ (.Y(_0320_),
    .A(net947));
 sg13g2_inv_1 _4789_ (.Y(_0321_),
    .A(net947));
 sg13g2_inv_1 _4790_ (.Y(_0322_),
    .A(net946));
 sg13g2_inv_1 _4791_ (.Y(_0323_),
    .A(net963));
 sg13g2_inv_1 _4792_ (.Y(_0324_),
    .A(net963));
 sg13g2_inv_1 _4793_ (.Y(_0325_),
    .A(net963));
 sg13g2_inv_1 _4794_ (.Y(_0326_),
    .A(net963));
 sg13g2_inv_1 _4795_ (.Y(_0327_),
    .A(net963));
 sg13g2_inv_1 _4796_ (.Y(_0328_),
    .A(net963));
 sg13g2_inv_1 _4797_ (.Y(_0329_),
    .A(net956));
 sg13g2_inv_1 _4798_ (.Y(_0330_),
    .A(net933));
 sg13g2_inv_1 _4799_ (.Y(_0331_),
    .A(net933));
 sg13g2_inv_1 _4800_ (.Y(_0332_),
    .A(net930));
 sg13g2_inv_1 _4801_ (.Y(_0333_),
    .A(net930));
 sg13g2_inv_1 _4802_ (.Y(_0334_),
    .A(net932));
 sg13g2_inv_1 _4803_ (.Y(_0335_),
    .A(net931));
 sg13g2_inv_1 _4804_ (.Y(_0336_),
    .A(net931));
 sg13g2_inv_1 _4805_ (.Y(_0337_),
    .A(net936));
 sg13g2_inv_1 _4806_ (.Y(_0338_),
    .A(net936));
 sg13g2_inv_1 _4807_ (.Y(_0339_),
    .A(net936));
 sg13g2_inv_1 _4808_ (.Y(_0340_),
    .A(net937));
 sg13g2_inv_1 _4809_ (.Y(_0341_),
    .A(net937));
 sg13g2_inv_1 _4810_ (.Y(_0342_),
    .A(net952));
 sg13g2_inv_1 _4811_ (.Y(_0343_),
    .A(net952));
 sg13g2_inv_1 _4812_ (.Y(_0344_),
    .A(net952));
 sg13g2_inv_1 _4813_ (.Y(_0345_),
    .A(net953));
 sg13g2_inv_1 _4814_ (.Y(_0346_),
    .A(net941));
 sg13g2_inv_1 _4815_ (.Y(_0347_),
    .A(net933));
 sg13g2_inv_1 _4816_ (.Y(_0348_),
    .A(net933));
 sg13g2_inv_1 _4817_ (.Y(_0349_),
    .A(net933));
 sg13g2_inv_1 _4818_ (.Y(_0350_),
    .A(net935));
 sg13g2_inv_1 _4819_ (.Y(_0351_),
    .A(net935));
 sg13g2_inv_1 _4820_ (.Y(_0352_),
    .A(net934));
 sg13g2_inv_1 _4821_ (.Y(_0353_),
    .A(net938));
 sg13g2_inv_1 _4822_ (.Y(_0354_),
    .A(net938));
 sg13g2_inv_1 _4823_ (.Y(_0355_),
    .A(net938));
 sg13g2_inv_1 _4824_ (.Y(_0356_),
    .A(net939));
 sg13g2_inv_1 _4825_ (.Y(_0357_),
    .A(net939));
 sg13g2_inv_1 _4826_ (.Y(_0358_),
    .A(net955));
 sg13g2_inv_1 _4827_ (.Y(_0359_),
    .A(net955));
 sg13g2_inv_1 _4828_ (.Y(_0360_),
    .A(net952));
 sg13g2_inv_1 _4829_ (.Y(_0361_),
    .A(net954));
 sg13g2_inv_1 _4830_ (.Y(_0362_),
    .A(net953));
 sg13g2_inv_1 _4831_ (.Y(_0363_),
    .A(net941));
 sg13g2_inv_1 _4832_ (.Y(_0364_),
    .A(net941));
 sg13g2_inv_1 _4833_ (.Y(_0365_),
    .A(net941));
 sg13g2_inv_1 _4834_ (.Y(_0366_),
    .A(net942));
 sg13g2_inv_1 _4835_ (.Y(_0367_),
    .A(net942));
 sg13g2_inv_1 _4836_ (.Y(_0368_),
    .A(net942));
 sg13g2_inv_1 _4837_ (.Y(_0369_),
    .A(net946));
 sg13g2_inv_1 _4838_ (.Y(_0370_),
    .A(net946));
 sg13g2_inv_1 _4839_ (.Y(_0371_),
    .A(net946));
 sg13g2_inv_1 _4840_ (.Y(_0372_),
    .A(net939));
 sg13g2_inv_1 _4841_ (.Y(_0373_),
    .A(net947));
 sg13g2_inv_1 _4842_ (.Y(_0374_),
    .A(net939));
 sg13g2_inv_1 _4843_ (.Y(_0375_),
    .A(net955));
 sg13g2_inv_1 _4844_ (.Y(_0376_),
    .A(net955));
 sg13g2_inv_1 _4845_ (.Y(_0377_),
    .A(net956));
 sg13g2_inv_1 _4846_ (.Y(_0378_),
    .A(net955));
 sg13g2_inv_1 _4847_ (.Y(_0379_),
    .A(net956));
 sg13g2_inv_1 _4848_ (.Y(_0380_),
    .A(net956));
 sg13g2_inv_1 _4849_ (.Y(_0381_),
    .A(net891));
 sg13g2_inv_1 _4850_ (.Y(_0382_),
    .A(net890));
 sg13g2_inv_1 _4851_ (.Y(_0383_),
    .A(net898));
 sg13g2_inv_1 _4852_ (.Y(_0384_),
    .A(net899));
 sg13g2_inv_1 _4853_ (.Y(_0385_),
    .A(net898));
 sg13g2_inv_1 _4854_ (.Y(_0386_),
    .A(net898));
 sg13g2_inv_1 _4855_ (.Y(_0387_),
    .A(net901));
 sg13g2_inv_1 _4856_ (.Y(_0388_),
    .A(net901));
 sg13g2_inv_1 _4857_ (.Y(_0389_),
    .A(net905));
 sg13g2_inv_1 _4858_ (.Y(_0390_),
    .A(net905));
 sg13g2_inv_1 _4859_ (.Y(_0391_),
    .A(net905));
 sg13g2_inv_1 _4860_ (.Y(_0392_),
    .A(net906));
 sg13g2_inv_1 _4861_ (.Y(_0393_),
    .A(net907));
 sg13g2_inv_1 _4862_ (.Y(_0394_),
    .A(net920));
 sg13g2_inv_1 _4863_ (.Y(_0395_),
    .A(net920));
 sg13g2_inv_1 _4864_ (.Y(_0396_),
    .A(net922));
 sg13g2_inv_1 _4865_ (.Y(_0397_),
    .A(net922));
 sg13g2_inv_2 _4866_ (.Y(_0715_),
    .A(net869));
 sg13g2_inv_1 _4867_ (.Y(_0716_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out0[13] ));
 sg13g2_inv_1 _4868_ (.Y(_0717_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out0[10] ));
 sg13g2_inv_1 _4869_ (.Y(_0718_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out0[0] ));
 sg13g2_inv_1 _4870_ (.Y(_0719_),
    .A(net829));
 sg13g2_inv_1 _4871_ (.Y(_0720_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out1[13] ));
 sg13g2_inv_1 _4872_ (.Y(_0721_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out1[11] ));
 sg13g2_inv_1 _4873_ (.Y(_0722_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out1[7] ));
 sg13g2_inv_1 _4874_ (.Y(_0723_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out1[2] ));
 sg13g2_inv_1 _4875_ (.Y(_0724_),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg1[13] ));
 sg13g2_inv_1 _4876_ (.Y(_0725_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out0[13] ));
 sg13g2_inv_1 _4877_ (.Y(_0726_),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg1[7] ));
 sg13g2_inv_1 _4878_ (.Y(_0727_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out0[7] ));
 sg13g2_inv_1 _4879_ (.Y(_0728_),
    .A(\u_ddc_top_level.cic_left_inst.in_data[10] ));
 sg13g2_inv_1 _4880_ (.Y(_0729_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[18] ));
 sg13g2_inv_1 _4881_ (.Y(_0730_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[17] ));
 sg13g2_inv_1 _4882_ (.Y(_0731_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[16] ));
 sg13g2_inv_1 _4883_ (.Y(_0732_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out2[0] ));
 sg13g2_inv_1 _4884_ (.Y(_0733_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out1[13] ));
 sg13g2_inv_1 _4885_ (.Y(_0734_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out1[9] ));
 sg13g2_inv_1 _4886_ (.Y(_0735_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out1[7] ));
 sg13g2_inv_1 _4887_ (.Y(_0736_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out1[0] ));
 sg13g2_inv_1 _4888_ (.Y(_0737_),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg1[13] ));
 sg13g2_inv_1 _4889_ (.Y(_0738_),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg0[13] ));
 sg13g2_inv_1 _4890_ (.Y(_0739_),
    .A(\u_ddc_top_level.cic_right_inst.in_data[13] ));
 sg13g2_inv_1 _4891_ (.Y(_0740_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[18] ));
 sg13g2_inv_1 _4892_ (.Y(_0741_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[17] ));
 sg13g2_inv_1 _4893_ (.Y(_0742_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[16] ));
 sg13g2_inv_1 _4894_ (.Y(_0743_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out2[0] ));
 sg13g2_inv_1 _4895_ (.Y(_0744_),
    .A(\u_ddc_top_level.cic_right_inst.int_reg0[18] ));
 sg13g2_inv_1 _4896_ (.Y(_0745_),
    .A(\u_ddc_top_level.cic_left_inst.int_reg0[17] ));
 sg13g2_inv_1 _4897_ (.Y(_0188_),
    .A(net887));
 sg13g2_nand2_1 _4898_ (.Y(_0746_),
    .A(\u_ddc_top_level.cic_right_inst.comb_out0[16] ),
    .B(net815));
 sg13g2_nor2b_1 _4899_ (.A(\u_ddc_top_level.cic_right_inst.comb_reg0[15] ),
    .B_N(\u_ddc_top_level.cic_right_inst.in_data[15] ),
    .Y(_0747_));
 sg13g2_xor2_1 _4900_ (.B(\u_ddc_top_level.cic_right_inst.in_data[15] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg0[15] ),
    .X(_0748_));
 sg13g2_nor2b_1 _4901_ (.A(\u_ddc_top_level.cic_right_inst.in_data[14] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg0[14] ),
    .Y(_0749_));
 sg13g2_xnor2_1 _4902_ (.Y(_0750_),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg0[14] ),
    .B(\u_ddc_top_level.cic_right_inst.in_data[14] ));
 sg13g2_nand2b_1 _4903_ (.Y(_0751_),
    .B(\u_ddc_top_level.cic_right_inst.in_data[7] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_reg0[7] ));
 sg13g2_nand2b_1 _4904_ (.Y(_0752_),
    .B(\u_ddc_top_level.cic_right_inst.in_data[5] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_reg0[5] ));
 sg13g2_nor2b_1 _4905_ (.A(\u_ddc_top_level.cic_right_inst.in_data[5] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg0[5] ),
    .Y(_0753_));
 sg13g2_nor2b_1 _4906_ (.A(\u_ddc_top_level.cic_right_inst.in_data[4] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg0[4] ),
    .Y(_0754_));
 sg13g2_nand2b_1 _4907_ (.Y(_0755_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg0[3] ),
    .A_N(\u_ddc_top_level.cic_right_inst.in_data[3] ));
 sg13g2_xor2_1 _4908_ (.B(\u_ddc_top_level.cic_right_inst.in_data[3] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg0[3] ),
    .X(_0756_));
 sg13g2_nor2b_1 _4909_ (.A(\u_ddc_top_level.cic_right_inst.in_data[2] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg0[2] ),
    .Y(_0757_));
 sg13g2_nand2b_1 _4910_ (.Y(_0758_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg0[1] ),
    .A_N(\u_ddc_top_level.cic_right_inst.in_data[1] ));
 sg13g2_nor2b_2 _4911_ (.A(\u_ddc_top_level.cic_right_inst.comb_reg0[0] ),
    .B_N(\u_ddc_top_level.cic_right_inst.in_data[0] ),
    .Y(_0759_));
 sg13g2_nor2b_1 _4912_ (.A(\u_ddc_top_level.cic_right_inst.comb_reg0[1] ),
    .B_N(\u_ddc_top_level.cic_right_inst.in_data[1] ),
    .Y(_0760_));
 sg13g2_xnor2_1 _4913_ (.Y(_0761_),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg0[1] ),
    .B(\u_ddc_top_level.cic_right_inst.in_data[1] ));
 sg13g2_o21ai_1 _4914_ (.B1(_0758_),
    .Y(_0762_),
    .A1(_0759_),
    .A2(_0760_));
 sg13g2_xnor2_1 _4915_ (.Y(_0763_),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg0[2] ),
    .B(\u_ddc_top_level.cic_right_inst.in_data[2] ));
 sg13g2_a21oi_1 _4916_ (.A1(_0762_),
    .A2(_0763_),
    .Y(_0764_),
    .B1(_0757_));
 sg13g2_o21ai_1 _4917_ (.B1(_0755_),
    .Y(_0765_),
    .A1(_0756_),
    .A2(_0764_));
 sg13g2_xnor2_1 _4918_ (.Y(_0766_),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg0[4] ),
    .B(\u_ddc_top_level.cic_right_inst.in_data[4] ));
 sg13g2_a21oi_1 _4919_ (.A1(_0765_),
    .A2(_0766_),
    .Y(_0767_),
    .B1(_0754_));
 sg13g2_xnor2_1 _4920_ (.Y(_0768_),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg0[5] ),
    .B(\u_ddc_top_level.cic_right_inst.in_data[5] ));
 sg13g2_and2_1 _4921_ (.A(_0766_),
    .B(_0768_),
    .X(_0769_));
 sg13g2_a221oi_1 _4922_ (.B2(_0769_),
    .C1(_0753_),
    .B1(_0765_),
    .A1(_0752_),
    .Y(_0770_),
    .A2(_0754_));
 sg13g2_nor2b_1 _4923_ (.A(\u_ddc_top_level.cic_right_inst.in_data[6] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg0[6] ),
    .Y(_0771_));
 sg13g2_xor2_1 _4924_ (.B(\u_ddc_top_level.cic_right_inst.in_data[6] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg0[6] ),
    .X(_0772_));
 sg13g2_nor2_1 _4925_ (.A(_0770_),
    .B(_0772_),
    .Y(_0773_));
 sg13g2_nor2b_1 _4926_ (.A(\u_ddc_top_level.cic_right_inst.in_data[7] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg0[7] ),
    .Y(_0774_));
 sg13g2_a21oi_1 _4927_ (.A1(_0751_),
    .A2(_0771_),
    .Y(_0775_),
    .B1(_0774_));
 sg13g2_xnor2_1 _4928_ (.Y(_0776_),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg0[7] ),
    .B(\u_ddc_top_level.cic_right_inst.in_data[7] ));
 sg13g2_nand2b_1 _4929_ (.Y(_0777_),
    .B(_0776_),
    .A_N(_0772_));
 sg13g2_o21ai_1 _4930_ (.B1(_0775_),
    .Y(_0778_),
    .A1(_0770_),
    .A2(_0777_));
 sg13g2_nand2b_1 _4931_ (.Y(_0779_),
    .B(\u_ddc_top_level.cic_right_inst.in_data[9] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_reg0[9] ));
 sg13g2_nor2b_1 _4932_ (.A(\u_ddc_top_level.cic_right_inst.in_data[9] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg0[9] ),
    .Y(_0780_));
 sg13g2_xnor2_1 _4933_ (.Y(_0781_),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg0[9] ),
    .B(\u_ddc_top_level.cic_right_inst.in_data[9] ));
 sg13g2_nor2b_1 _4934_ (.A(\u_ddc_top_level.cic_right_inst.in_data[8] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg0[8] ),
    .Y(_0782_));
 sg13g2_xnor2_1 _4935_ (.Y(_0783_),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg0[8] ),
    .B(\u_ddc_top_level.cic_right_inst.in_data[8] ));
 sg13g2_and3_1 _4936_ (.X(_0784_),
    .A(_0778_),
    .B(_0781_),
    .C(_0783_));
 sg13g2_inv_1 _4937_ (.Y(_0785_),
    .A(_0784_));
 sg13g2_a21oi_1 _4938_ (.A1(_0779_),
    .A2(_0782_),
    .Y(_0786_),
    .B1(_0780_));
 sg13g2_nor2b_1 _4939_ (.A(\u_ddc_top_level.cic_right_inst.in_data[10] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg0[10] ),
    .Y(_0787_));
 sg13g2_nor2b_1 _4940_ (.A(\u_ddc_top_level.cic_right_inst.comb_reg0[11] ),
    .B_N(\u_ddc_top_level.cic_right_inst.in_data[11] ),
    .Y(_0788_));
 sg13g2_nand2b_1 _4941_ (.Y(_0789_),
    .B(_0787_),
    .A_N(_0788_));
 sg13g2_nand2b_1 _4942_ (.Y(_0790_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg0[11] ),
    .A_N(\u_ddc_top_level.cic_right_inst.in_data[11] ));
 sg13g2_nand3_1 _4943_ (.B(_0789_),
    .C(_0790_),
    .A(_0786_),
    .Y(_0791_));
 sg13g2_nor2b_1 _4944_ (.A(\u_ddc_top_level.cic_right_inst.comb_reg0[10] ),
    .B_N(\u_ddc_top_level.cic_right_inst.in_data[10] ),
    .Y(_0792_));
 sg13g2_o21ai_1 _4945_ (.B1(_0790_),
    .Y(_0793_),
    .A1(_0788_),
    .A2(_0792_));
 sg13g2_o21ai_1 _4946_ (.B1(_0793_),
    .Y(_0794_),
    .A1(_0784_),
    .A2(_0791_));
 sg13g2_xnor2_1 _4947_ (.Y(_0795_),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg0[13] ),
    .B(\u_ddc_top_level.cic_right_inst.in_data[13] ));
 sg13g2_nand2b_1 _4948_ (.Y(_0796_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg0[12] ),
    .A_N(\u_ddc_top_level.cic_right_inst.in_data[12] ));
 sg13g2_xor2_1 _4949_ (.B(\u_ddc_top_level.cic_right_inst.in_data[12] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg0[12] ),
    .X(_0797_));
 sg13g2_inv_1 _4950_ (.Y(_0798_),
    .A(_0797_));
 sg13g2_nand2_1 _4951_ (.Y(_0799_),
    .A(_0795_),
    .B(_0798_));
 sg13g2_a21oi_1 _4952_ (.A1(_0738_),
    .A2(\u_ddc_top_level.cic_right_inst.in_data[13] ),
    .Y(_0800_),
    .B1(_0796_));
 sg13g2_a21oi_1 _4953_ (.A1(\u_ddc_top_level.cic_right_inst.comb_reg0[13] ),
    .A2(_0739_),
    .Y(_0801_),
    .B1(_0800_));
 sg13g2_o21ai_1 _4954_ (.B1(_0801_),
    .Y(_0802_),
    .A1(_0794_),
    .A2(_0799_));
 sg13g2_a21oi_1 _4955_ (.A1(_0750_),
    .A2(_0802_),
    .Y(_0803_),
    .B1(_0749_));
 sg13g2_o21ai_1 _4956_ (.B1(net876),
    .Y(_0804_),
    .A1(_0748_),
    .A2(_0803_));
 sg13g2_o21ai_1 _4957_ (.B1(_0746_),
    .Y(_0680_),
    .A1(_0747_),
    .A2(_0804_));
 sg13g2_nand2_1 _4958_ (.Y(_0805_),
    .A(net815),
    .B(\u_ddc_top_level.cic_right_inst.comb_out0[15] ));
 sg13g2_and2_1 _4959_ (.A(_0748_),
    .B(_0803_),
    .X(_0806_));
 sg13g2_o21ai_1 _4960_ (.B1(_0805_),
    .Y(_0679_),
    .A1(_0804_),
    .A2(_0806_));
 sg13g2_nor2_1 _4961_ (.A(net877),
    .B(\u_ddc_top_level.cic_right_inst.comb_out0[14] ),
    .Y(_0807_));
 sg13g2_xnor2_1 _4962_ (.Y(_0808_),
    .A(_0750_),
    .B(_0802_));
 sg13g2_a21oi_1 _4963_ (.A1(net877),
    .A2(_0808_),
    .Y(_0678_),
    .B1(_0807_));
 sg13g2_o21ai_1 _4964_ (.B1(_0796_),
    .Y(_0809_),
    .A1(_0794_),
    .A2(_0797_));
 sg13g2_o21ai_1 _4965_ (.B1(net875),
    .Y(_0810_),
    .A1(_0795_),
    .A2(_0809_));
 sg13g2_a21o_1 _4966_ (.A2(_0809_),
    .A1(_0795_),
    .B1(_0810_),
    .X(_0811_));
 sg13g2_o21ai_1 _4967_ (.B1(_0811_),
    .Y(_0677_),
    .A1(net874),
    .A2(_0716_));
 sg13g2_o21ai_1 _4968_ (.B1(net875),
    .Y(_0812_),
    .A1(_0794_),
    .A2(_0797_));
 sg13g2_a21oi_1 _4969_ (.A1(_0794_),
    .A2(_0797_),
    .Y(_0813_),
    .B1(_0812_));
 sg13g2_a21o_1 _4970_ (.A2(\u_ddc_top_level.cic_right_inst.comb_out0[12] ),
    .A1(net816),
    .B1(_0813_),
    .X(_0676_));
 sg13g2_nor2b_1 _4971_ (.A(_0788_),
    .B_N(_0790_),
    .Y(_0814_));
 sg13g2_or2_1 _4972_ (.X(_0815_),
    .B(_0792_),
    .A(_0787_));
 sg13g2_a21oi_1 _4973_ (.A1(_0785_),
    .A2(_0786_),
    .Y(_0816_),
    .B1(_0815_));
 sg13g2_nor2_1 _4974_ (.A(_0787_),
    .B(_0816_),
    .Y(_0817_));
 sg13g2_xnor2_1 _4975_ (.Y(_0818_),
    .A(_0814_),
    .B(_0817_));
 sg13g2_mux2_1 _4976_ (.A0(\u_ddc_top_level.cic_right_inst.comb_out0[11] ),
    .A1(_0818_),
    .S(net874),
    .X(_0675_));
 sg13g2_nand3_1 _4977_ (.B(_0786_),
    .C(_0815_),
    .A(_0785_),
    .Y(_0819_));
 sg13g2_nand3b_1 _4978_ (.B(_0819_),
    .C(net875),
    .Y(_0820_),
    .A_N(_0816_));
 sg13g2_o21ai_1 _4979_ (.B1(_0820_),
    .Y(_0674_),
    .A1(net874),
    .A2(_0717_));
 sg13g2_a21oi_1 _4980_ (.A1(_0778_),
    .A2(_0783_),
    .Y(_0821_),
    .B1(_0782_));
 sg13g2_xnor2_1 _4981_ (.Y(_0822_),
    .A(_0781_),
    .B(_0821_));
 sg13g2_mux2_1 _4982_ (.A0(\u_ddc_top_level.cic_right_inst.comb_out0[9] ),
    .A1(_0822_),
    .S(net870),
    .X(_0673_));
 sg13g2_nor2_1 _4983_ (.A(net870),
    .B(\u_ddc_top_level.cic_right_inst.comb_out0[8] ),
    .Y(_0823_));
 sg13g2_xnor2_1 _4984_ (.Y(_0824_),
    .A(_0778_),
    .B(_0783_));
 sg13g2_a21oi_1 _4985_ (.A1(net870),
    .A2(_0824_),
    .Y(_0672_),
    .B1(_0823_));
 sg13g2_nor2_1 _4986_ (.A(_0771_),
    .B(_0773_),
    .Y(_0825_));
 sg13g2_xnor2_1 _4987_ (.Y(_0826_),
    .A(_0776_),
    .B(_0825_));
 sg13g2_mux2_1 _4988_ (.A0(\u_ddc_top_level.cic_right_inst.comb_out0[7] ),
    .A1(_0826_),
    .S(net870),
    .X(_0671_));
 sg13g2_o21ai_1 _4989_ (.B1(net871),
    .Y(_0827_),
    .A1(_0770_),
    .A2(_0772_));
 sg13g2_a21oi_1 _4990_ (.A1(_0770_),
    .A2(_0772_),
    .Y(_0828_),
    .B1(_0827_));
 sg13g2_a21o_1 _4991_ (.A2(\u_ddc_top_level.cic_right_inst.comb_out0[6] ),
    .A1(net813),
    .B1(_0828_),
    .X(_0670_));
 sg13g2_xor2_1 _4992_ (.B(_0768_),
    .A(_0767_),
    .X(_0829_));
 sg13g2_nor2_1 _4993_ (.A(net869),
    .B(\u_ddc_top_level.cic_right_inst.comb_out0[5] ),
    .Y(_0830_));
 sg13g2_a21oi_1 _4994_ (.A1(net869),
    .A2(_0829_),
    .Y(_0669_),
    .B1(_0830_));
 sg13g2_xnor2_1 _4995_ (.Y(_0831_),
    .A(_0765_),
    .B(_0766_));
 sg13g2_nor2_1 _4996_ (.A(net869),
    .B(\u_ddc_top_level.cic_right_inst.comb_out0[4] ),
    .Y(_0832_));
 sg13g2_a21oi_1 _4997_ (.A1(net869),
    .A2(_0831_),
    .Y(_0668_),
    .B1(_0832_));
 sg13g2_nor2_1 _4998_ (.A(net865),
    .B(\u_ddc_top_level.cic_right_inst.comb_out0[3] ),
    .Y(_0833_));
 sg13g2_xnor2_1 _4999_ (.Y(_0834_),
    .A(_0756_),
    .B(_0764_));
 sg13g2_a21oi_1 _5000_ (.A1(net865),
    .A2(_0834_),
    .Y(_0667_),
    .B1(_0833_));
 sg13g2_nor2_1 _5001_ (.A(net864),
    .B(\u_ddc_top_level.cic_right_inst.comb_out0[2] ),
    .Y(_0835_));
 sg13g2_xnor2_1 _5002_ (.Y(_0836_),
    .A(_0762_),
    .B(_0763_));
 sg13g2_a21oi_1 _5003_ (.A1(net864),
    .A2(_0836_),
    .Y(_0666_),
    .B1(_0835_));
 sg13g2_xnor2_1 _5004_ (.Y(_0837_),
    .A(_0759_),
    .B(_0761_));
 sg13g2_mux2_1 _5005_ (.A0(\u_ddc_top_level.cic_right_inst.comb_out0[1] ),
    .A1(_0837_),
    .S(net855),
    .X(_0665_));
 sg13g2_nand2b_1 _5006_ (.Y(_0838_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg0[0] ),
    .A_N(\u_ddc_top_level.cic_right_inst.in_data[0] ));
 sg13g2_nor2_1 _5007_ (.A(net814),
    .B(_0759_),
    .Y(_0839_));
 sg13g2_a22oi_1 _5008_ (.Y(_0664_),
    .B1(_0838_),
    .B2(_0839_),
    .A2(_0718_),
    .A1(net814));
 sg13g2_mux2_1 _5009_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg2[17] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out1[17] ),
    .S(net843),
    .X(_0663_));
 sg13g2_mux2_1 _5010_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg2[16] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out1[16] ),
    .S(net843),
    .X(_0662_));
 sg13g2_mux2_1 _5011_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg2[15] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out1[15] ),
    .S(net847),
    .X(_0661_));
 sg13g2_mux2_1 _5012_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg2[14] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out1[14] ),
    .S(net847),
    .X(_0660_));
 sg13g2_nor2_1 _5013_ (.A(net847),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg2[13] ),
    .Y(_0840_));
 sg13g2_a21oi_1 _5014_ (.A1(net847),
    .A2(_0720_),
    .Y(_0659_),
    .B1(_0840_));
 sg13g2_mux2_1 _5015_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg2[12] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out1[12] ),
    .S(net846),
    .X(_0658_));
 sg13g2_nor2_1 _5016_ (.A(net846),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg2[11] ),
    .Y(_0841_));
 sg13g2_a21oi_1 _5017_ (.A1(net846),
    .A2(_0721_),
    .Y(_0657_),
    .B1(_0841_));
 sg13g2_mux2_1 _5018_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg2[10] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out1[10] ),
    .S(net846),
    .X(_0656_));
 sg13g2_mux2_1 _5019_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg2[9] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out1[9] ),
    .S(net846),
    .X(_0655_));
 sg13g2_mux2_1 _5020_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg2[8] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out1[8] ),
    .S(net846),
    .X(_0654_));
 sg13g2_nor2_1 _5021_ (.A(net834),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg2[7] ),
    .Y(_0842_));
 sg13g2_a21oi_1 _5022_ (.A1(net834),
    .A2(_0722_),
    .Y(_0653_),
    .B1(_0842_));
 sg13g2_mux2_1 _5023_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg2[6] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out1[6] ),
    .S(net834),
    .X(_0652_));
 sg13g2_mux2_1 _5024_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg2[5] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out1[5] ),
    .S(net834),
    .X(_0651_));
 sg13g2_mux2_1 _5025_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg2[4] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out1[4] ),
    .S(net834),
    .X(_0650_));
 sg13g2_mux2_1 _5026_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg2[3] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out1[3] ),
    .S(net830),
    .X(_0649_));
 sg13g2_nor2_1 _5027_ (.A(net830),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg2[2] ),
    .Y(_0843_));
 sg13g2_a21oi_1 _5028_ (.A1(net830),
    .A2(_0723_),
    .Y(_0648_),
    .B1(_0843_));
 sg13g2_mux2_1 _5029_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg2[1] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out1[1] ),
    .S(net831),
    .X(_0647_));
 sg13g2_mux2_1 _5030_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg2[0] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out1[0] ),
    .S(net831),
    .X(_0646_));
 sg13g2_mux2_1 _5031_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg1[16] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out0[16] ),
    .S(net842),
    .X(_0625_));
 sg13g2_mux2_1 _5032_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg1[15] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out0[15] ),
    .S(net842),
    .X(_0624_));
 sg13g2_mux2_1 _5033_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg1[14] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out0[14] ),
    .S(net842),
    .X(_0623_));
 sg13g2_nor2_1 _5034_ (.A(net851),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg1[13] ),
    .Y(_0844_));
 sg13g2_a21oi_1 _5035_ (.A1(net843),
    .A2(_0725_),
    .Y(_0622_),
    .B1(_0844_));
 sg13g2_mux2_1 _5036_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg1[12] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out0[12] ),
    .S(net841),
    .X(_0621_));
 sg13g2_mux2_1 _5037_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg1[11] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out0[11] ),
    .S(net840),
    .X(_0620_));
 sg13g2_mux2_1 _5038_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg1[10] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out0[10] ),
    .S(net840),
    .X(_0619_));
 sg13g2_mux2_1 _5039_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg1[9] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out0[9] ),
    .S(net827),
    .X(_0618_));
 sg13g2_mux2_1 _5040_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg1[8] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out0[8] ),
    .S(net827),
    .X(_0617_));
 sg13g2_nor2_1 _5041_ (.A(net827),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg1[7] ),
    .Y(_0845_));
 sg13g2_a21oi_1 _5042_ (.A1(net827),
    .A2(_0727_),
    .Y(_0616_),
    .B1(_0845_));
 sg13g2_mux2_1 _5043_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg1[6] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out0[6] ),
    .S(net827),
    .X(_0615_));
 sg13g2_mux2_1 _5044_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg1[5] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out0[5] ),
    .S(net827),
    .X(_0614_));
 sg13g2_mux2_1 _5045_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg1[4] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out0[4] ),
    .S(net825),
    .X(_0613_));
 sg13g2_mux2_1 _5046_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg1[3] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out0[3] ),
    .S(net825),
    .X(_0612_));
 sg13g2_mux2_1 _5047_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg1[2] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out0[2] ),
    .S(net824),
    .X(_0611_));
 sg13g2_mux2_1 _5048_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg1[1] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out0[1] ),
    .S(net829),
    .X(_0610_));
 sg13g2_mux2_1 _5049_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg1[0] ),
    .A1(\u_ddc_top_level.cic_left_inst.comb_out0[0] ),
    .S(net829),
    .X(_0609_));
 sg13g2_mux2_1 _5050_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg0[15] ),
    .A1(\u_ddc_top_level.cic_left_inst.in_data[15] ),
    .S(net843),
    .X(_0608_));
 sg13g2_mux2_1 _5051_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg0[14] ),
    .A1(\u_ddc_top_level.cic_left_inst.in_data[14] ),
    .S(net842),
    .X(_0607_));
 sg13g2_mux2_1 _5052_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg0[13] ),
    .A1(\u_ddc_top_level.cic_left_inst.in_data[13] ),
    .S(net842),
    .X(_0606_));
 sg13g2_mux2_1 _5053_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg0[12] ),
    .A1(\u_ddc_top_level.cic_left_inst.in_data[12] ),
    .S(net841),
    .X(_0605_));
 sg13g2_mux2_1 _5054_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg0[11] ),
    .A1(\u_ddc_top_level.cic_left_inst.in_data[11] ),
    .S(net839),
    .X(_0604_));
 sg13g2_nor2_1 _5055_ (.A(net839),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg0[10] ),
    .Y(_0846_));
 sg13g2_a21oi_1 _5056_ (.A1(net839),
    .A2(_0728_),
    .Y(_0603_),
    .B1(_0846_));
 sg13g2_mux2_1 _5057_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg0[9] ),
    .A1(\u_ddc_top_level.cic_left_inst.in_data[9] ),
    .S(net828),
    .X(_0602_));
 sg13g2_mux2_1 _5058_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg0[8] ),
    .A1(\u_ddc_top_level.cic_left_inst.in_data[8] ),
    .S(net828),
    .X(_0601_));
 sg13g2_mux2_1 _5059_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg0[7] ),
    .A1(\u_ddc_top_level.cic_left_inst.in_data[7] ),
    .S(net828),
    .X(_0600_));
 sg13g2_mux2_1 _5060_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg0[6] ),
    .A1(\u_ddc_top_level.cic_left_inst.in_data[6] ),
    .S(net828),
    .X(_0599_));
 sg13g2_mux2_1 _5061_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg0[5] ),
    .A1(\u_ddc_top_level.cic_left_inst.in_data[5] ),
    .S(net826),
    .X(_0598_));
 sg13g2_mux2_1 _5062_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg0[4] ),
    .A1(\u_ddc_top_level.cic_left_inst.in_data[4] ),
    .S(net826),
    .X(_0597_));
 sg13g2_mux2_1 _5063_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg0[3] ),
    .A1(\u_ddc_top_level.cic_left_inst.in_data[3] ),
    .S(net826),
    .X(_0596_));
 sg13g2_mux2_1 _5064_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg0[2] ),
    .A1(\u_ddc_top_level.cic_left_inst.in_data[2] ),
    .S(net826),
    .X(_0595_));
 sg13g2_mux2_1 _5065_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg0[1] ),
    .A1(\u_ddc_top_level.cic_left_inst.in_data[1] ),
    .S(net824),
    .X(_0594_));
 sg13g2_mux2_1 _5066_ (.A0(\u_ddc_top_level.cic_left_inst.comb_reg0[0] ),
    .A1(\u_ddc_top_level.cic_left_inst.in_data[0] ),
    .S(net824),
    .X(_0593_));
 sg13g2_nand2b_1 _5067_ (.Y(_0847_),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg2[17] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_out1[17] ));
 sg13g2_xnor2_1 _5068_ (.Y(_0848_),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg2[17] ),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[17] ));
 sg13g2_nand2b_1 _5069_ (.Y(_0849_),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg2[16] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_out1[16] ));
 sg13g2_nor2_1 _5070_ (.A(\u_ddc_top_level.cic_left_inst.comb_reg2[7] ),
    .B(_0722_),
    .Y(_0850_));
 sg13g2_nor2b_1 _5071_ (.A(\u_ddc_top_level.cic_left_inst.comb_out1[6] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg2[6] ),
    .Y(_0851_));
 sg13g2_xnor2_1 _5072_ (.Y(_0852_),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg2[6] ),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[6] ));
 sg13g2_nor2b_1 _5073_ (.A(\u_ddc_top_level.cic_left_inst.comb_reg2[5] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_out1[5] ),
    .Y(_0853_));
 sg13g2_nand2b_1 _5074_ (.Y(_0854_),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg2[5] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_out1[5] ));
 sg13g2_nand2b_1 _5075_ (.Y(_0855_),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg2[4] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_out1[4] ));
 sg13g2_nand2b_1 _5076_ (.Y(_0856_),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg2[3] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_out1[3] ));
 sg13g2_xor2_1 _5077_ (.B(\u_ddc_top_level.cic_left_inst.comb_out1[3] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg2[3] ),
    .X(_0857_));
 sg13g2_nor2b_1 _5078_ (.A(\u_ddc_top_level.cic_left_inst.comb_out1[2] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg2[2] ),
    .Y(_0858_));
 sg13g2_nand2b_1 _5079_ (.Y(_0859_),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg2[1] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_out1[1] ));
 sg13g2_nor2b_1 _5080_ (.A(\u_ddc_top_level.cic_left_inst.comb_reg2[0] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_out1[0] ),
    .Y(_0860_));
 sg13g2_nor2b_1 _5081_ (.A(\u_ddc_top_level.cic_left_inst.comb_reg2[1] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_out1[1] ),
    .Y(_0861_));
 sg13g2_xnor2_1 _5082_ (.Y(_0862_),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg2[1] ),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[1] ));
 sg13g2_o21ai_1 _5083_ (.B1(_0859_),
    .Y(_0863_),
    .A1(_0860_),
    .A2(_0861_));
 sg13g2_xnor2_1 _5084_ (.Y(_0864_),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg2[2] ),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[2] ));
 sg13g2_a21oi_1 _5085_ (.A1(_0863_),
    .A2(_0864_),
    .Y(_0865_),
    .B1(_0858_));
 sg13g2_o21ai_1 _5086_ (.B1(_0856_),
    .Y(_0866_),
    .A1(_0857_),
    .A2(_0865_));
 sg13g2_xnor2_1 _5087_ (.Y(_0867_),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg2[4] ),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[4] ));
 sg13g2_nand2_1 _5088_ (.Y(_0868_),
    .A(_0866_),
    .B(_0867_));
 sg13g2_and2_1 _5089_ (.A(_0855_),
    .B(_0868_),
    .X(_0869_));
 sg13g2_o21ai_1 _5090_ (.B1(_0854_),
    .Y(_0870_),
    .A1(_0853_),
    .A2(_0855_));
 sg13g2_nor2b_1 _5091_ (.A(_0853_),
    .B_N(_0854_),
    .Y(_0871_));
 sg13g2_and2_1 _5092_ (.A(_0867_),
    .B(_0871_),
    .X(_0872_));
 sg13g2_a21o_1 _5093_ (.A2(_0872_),
    .A1(_0866_),
    .B1(_0870_),
    .X(_0873_));
 sg13g2_a21oi_1 _5094_ (.A1(_0852_),
    .A2(_0873_),
    .Y(_0874_),
    .B1(_0851_));
 sg13g2_a221oi_1 _5095_ (.B2(_0873_),
    .C1(_0851_),
    .B1(_0852_),
    .A1(\u_ddc_top_level.cic_left_inst.comb_reg2[7] ),
    .Y(_0875_),
    .A2(_0722_));
 sg13g2_nor2_1 _5096_ (.A(_0850_),
    .B(_0875_),
    .Y(_0876_));
 sg13g2_nor2b_1 _5097_ (.A(\u_ddc_top_level.cic_left_inst.comb_out1[11] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg2[11] ),
    .Y(_0877_));
 sg13g2_nand2b_1 _5098_ (.Y(_0878_),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[11] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_reg2[11] ));
 sg13g2_nor2b_1 _5099_ (.A(_0877_),
    .B_N(_0878_),
    .Y(_0879_));
 sg13g2_nor2b_1 _5100_ (.A(\u_ddc_top_level.cic_left_inst.comb_out1[10] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg2[10] ),
    .Y(_0880_));
 sg13g2_xor2_1 _5101_ (.B(\u_ddc_top_level.cic_left_inst.comb_out1[10] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg2[10] ),
    .X(_0881_));
 sg13g2_inv_1 _5102_ (.Y(_0882_),
    .A(_0881_));
 sg13g2_nand2_1 _5103_ (.Y(_0883_),
    .A(_0879_),
    .B(_0882_));
 sg13g2_nor2b_1 _5104_ (.A(\u_ddc_top_level.cic_left_inst.comb_out1[9] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg2[9] ),
    .Y(_0884_));
 sg13g2_nand2b_1 _5105_ (.Y(_0885_),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[9] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_reg2[9] ));
 sg13g2_nand2b_1 _5106_ (.Y(_0886_),
    .B(_0885_),
    .A_N(_0884_));
 sg13g2_nor2b_1 _5107_ (.A(\u_ddc_top_level.cic_left_inst.comb_out1[8] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg2[8] ),
    .Y(_0887_));
 sg13g2_xnor2_1 _5108_ (.Y(_0888_),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg2[8] ),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[8] ));
 sg13g2_nor2b_1 _5109_ (.A(_0886_),
    .B_N(_0888_),
    .Y(_0889_));
 sg13g2_inv_1 _5110_ (.Y(_0890_),
    .A(_0889_));
 sg13g2_nor4_2 _5111_ (.A(_0850_),
    .B(_0875_),
    .C(_0883_),
    .Y(_0891_),
    .D(_0890_));
 sg13g2_a21oi_2 _5112_ (.B1(_0884_),
    .Y(_0892_),
    .A2(_0887_),
    .A1(_0885_));
 sg13g2_a21oi_1 _5113_ (.A1(_0878_),
    .A2(_0880_),
    .Y(_0893_),
    .B1(_0877_));
 sg13g2_o21ai_1 _5114_ (.B1(_0893_),
    .Y(_0894_),
    .A1(_0883_),
    .A2(_0892_));
 sg13g2_nor2_2 _5115_ (.A(_0891_),
    .B(_0894_),
    .Y(_0895_));
 sg13g2_nand2b_1 _5116_ (.Y(_0896_),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg2[15] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_out1[15] ));
 sg13g2_nand2b_1 _5117_ (.Y(_0897_),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[15] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_reg2[15] ));
 sg13g2_and2_1 _5118_ (.A(_0896_),
    .B(_0897_),
    .X(_0898_));
 sg13g2_nor2b_1 _5119_ (.A(\u_ddc_top_level.cic_left_inst.comb_out1[14] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg2[14] ),
    .Y(_0899_));
 sg13g2_xor2_1 _5120_ (.B(\u_ddc_top_level.cic_left_inst.comb_out1[14] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg2[14] ),
    .X(_0900_));
 sg13g2_inv_1 _5121_ (.Y(_0901_),
    .A(_0900_));
 sg13g2_nand2_1 _5122_ (.Y(_0902_),
    .A(_0898_),
    .B(_0901_));
 sg13g2_nor2b_1 _5123_ (.A(\u_ddc_top_level.cic_left_inst.comb_out1[13] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg2[13] ),
    .Y(_0903_));
 sg13g2_nand2b_1 _5124_ (.Y(_0904_),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[13] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_reg2[13] ));
 sg13g2_nand2b_1 _5125_ (.Y(_0905_),
    .B(_0904_),
    .A_N(_0903_));
 sg13g2_nor2b_1 _5126_ (.A(\u_ddc_top_level.cic_left_inst.comb_out1[12] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg2[12] ),
    .Y(_0906_));
 sg13g2_xor2_1 _5127_ (.B(\u_ddc_top_level.cic_left_inst.comb_out1[12] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg2[12] ),
    .X(_0907_));
 sg13g2_or2_1 _5128_ (.X(_0908_),
    .B(_0907_),
    .A(_0905_));
 sg13g2_nor2_1 _5129_ (.A(_0902_),
    .B(_0908_),
    .Y(_0909_));
 sg13g2_o21ai_1 _5130_ (.B1(_0909_),
    .Y(_0910_),
    .A1(_0891_),
    .A2(_0894_));
 sg13g2_a21oi_1 _5131_ (.A1(_0904_),
    .A2(_0906_),
    .Y(_0911_),
    .B1(_0903_));
 sg13g2_o21ai_1 _5132_ (.B1(_0896_),
    .Y(_0912_),
    .A1(_0902_),
    .A2(_0911_));
 sg13g2_a21oi_1 _5133_ (.A1(_0897_),
    .A2(_0899_),
    .Y(_0913_),
    .B1(_0912_));
 sg13g2_xor2_1 _5134_ (.B(\u_ddc_top_level.cic_left_inst.comb_out1[16] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg2[16] ),
    .X(_0914_));
 sg13g2_a21o_1 _5135_ (.A2(_0913_),
    .A1(_0910_),
    .B1(_0914_),
    .X(_0915_));
 sg13g2_nand3_1 _5136_ (.B(_0849_),
    .C(_0915_),
    .A(_0848_),
    .Y(_0916_));
 sg13g2_and2_1 _5137_ (.A(net847),
    .B(_0916_),
    .X(_0917_));
 sg13g2_a22oi_1 _5138_ (.Y(_0592_),
    .B1(_0847_),
    .B2(_0917_),
    .A2(_0729_),
    .A1(net808));
 sg13g2_a21o_1 _5139_ (.A2(_0915_),
    .A1(_0849_),
    .B1(_0848_),
    .X(_0918_));
 sg13g2_a22oi_1 _5140_ (.Y(_0591_),
    .B1(_0917_),
    .B2(_0918_),
    .A2(_0730_),
    .A1(net810));
 sg13g2_nand3_1 _5141_ (.B(_0913_),
    .C(_0914_),
    .A(_0910_),
    .Y(_0919_));
 sg13g2_a21oi_1 _5142_ (.A1(_0915_),
    .A2(_0919_),
    .Y(_0920_),
    .B1(net810));
 sg13g2_a21oi_1 _5143_ (.A1(net810),
    .A2(_0731_),
    .Y(_0590_),
    .B1(_0920_));
 sg13g2_o21ai_1 _5144_ (.B1(_0911_),
    .Y(_0921_),
    .A1(_0895_),
    .A2(_0908_));
 sg13g2_a21oi_1 _5145_ (.A1(_0901_),
    .A2(_0921_),
    .Y(_0922_),
    .B1(_0899_));
 sg13g2_nand2_1 _5146_ (.Y(_0923_),
    .A(net810),
    .B(\u_ddc_top_level.cic_left_inst.comb_out2[15] ));
 sg13g2_xor2_1 _5147_ (.B(_0922_),
    .A(_0898_),
    .X(_0924_));
 sg13g2_o21ai_1 _5148_ (.B1(_0923_),
    .Y(_0589_),
    .A1(net810),
    .A2(_0924_));
 sg13g2_nor2_1 _5149_ (.A(net848),
    .B(\u_ddc_top_level.cic_left_inst.comb_out2[14] ),
    .Y(_0925_));
 sg13g2_xnor2_1 _5150_ (.Y(_0926_),
    .A(_0901_),
    .B(_0921_));
 sg13g2_a21oi_1 _5151_ (.A1(net847),
    .A2(_0926_),
    .Y(_0588_),
    .B1(_0925_));
 sg13g2_nor2_1 _5152_ (.A(_0895_),
    .B(_0907_),
    .Y(_0927_));
 sg13g2_nor2_1 _5153_ (.A(_0906_),
    .B(_0927_),
    .Y(_0928_));
 sg13g2_nor2_1 _5154_ (.A(net848),
    .B(\u_ddc_top_level.cic_left_inst.comb_out2[13] ),
    .Y(_0929_));
 sg13g2_xnor2_1 _5155_ (.Y(_0930_),
    .A(_0905_),
    .B(_0928_));
 sg13g2_a21oi_1 _5156_ (.A1(net848),
    .A2(_0930_),
    .Y(_0587_),
    .B1(_0929_));
 sg13g2_o21ai_1 _5157_ (.B1(net846),
    .Y(_0931_),
    .A1(_0895_),
    .A2(_0907_));
 sg13g2_a21oi_1 _5158_ (.A1(_0895_),
    .A2(_0907_),
    .Y(_0932_),
    .B1(_0931_));
 sg13g2_a21o_1 _5159_ (.A2(\u_ddc_top_level.cic_left_inst.comb_out2[12] ),
    .A1(net810),
    .B1(_0932_),
    .X(_0586_));
 sg13g2_nand2_1 _5160_ (.Y(_0933_),
    .A(_0876_),
    .B(_0889_));
 sg13g2_a21oi_1 _5161_ (.A1(_0892_),
    .A2(_0933_),
    .Y(_0934_),
    .B1(_0881_));
 sg13g2_nor2_1 _5162_ (.A(_0880_),
    .B(_0934_),
    .Y(_0935_));
 sg13g2_xnor2_1 _5163_ (.Y(_0936_),
    .A(_0879_),
    .B(_0935_));
 sg13g2_mux2_1 _5164_ (.A0(\u_ddc_top_level.cic_left_inst.comb_out2[11] ),
    .A1(_0936_),
    .S(net844),
    .X(_0585_));
 sg13g2_nor2_1 _5165_ (.A(net845),
    .B(\u_ddc_top_level.cic_left_inst.comb_out2[10] ),
    .Y(_0937_));
 sg13g2_nand3_1 _5166_ (.B(_0892_),
    .C(_0933_),
    .A(_0881_),
    .Y(_0938_));
 sg13g2_nand2b_1 _5167_ (.Y(_0939_),
    .B(_0938_),
    .A_N(_0934_));
 sg13g2_a21oi_1 _5168_ (.A1(net845),
    .A2(_0939_),
    .Y(_0584_),
    .B1(_0937_));
 sg13g2_a21oi_1 _5169_ (.A1(_0876_),
    .A2(_0888_),
    .Y(_0940_),
    .B1(_0887_));
 sg13g2_nor2_1 _5170_ (.A(net844),
    .B(\u_ddc_top_level.cic_left_inst.comb_out2[9] ),
    .Y(_0941_));
 sg13g2_xnor2_1 _5171_ (.Y(_0942_),
    .A(_0886_),
    .B(_0940_));
 sg13g2_a21oi_1 _5172_ (.A1(net844),
    .A2(_0942_),
    .Y(_0583_),
    .B1(_0941_));
 sg13g2_nor2_1 _5173_ (.A(net844),
    .B(\u_ddc_top_level.cic_left_inst.comb_out2[8] ),
    .Y(_0943_));
 sg13g2_xnor2_1 _5174_ (.Y(_0944_),
    .A(_0876_),
    .B(_0888_));
 sg13g2_a21oi_1 _5175_ (.A1(net844),
    .A2(_0944_),
    .Y(_0582_),
    .B1(_0943_));
 sg13g2_xnor2_1 _5176_ (.Y(_0945_),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg2[7] ),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[7] ));
 sg13g2_xnor2_1 _5177_ (.Y(_0946_),
    .A(_0874_),
    .B(_0945_));
 sg13g2_mux2_1 _5178_ (.A0(\u_ddc_top_level.cic_left_inst.comb_out2[7] ),
    .A1(_0946_),
    .S(net836),
    .X(_0581_));
 sg13g2_xnor2_1 _5179_ (.Y(_0947_),
    .A(_0852_),
    .B(_0873_));
 sg13g2_nor2_1 _5180_ (.A(net836),
    .B(\u_ddc_top_level.cic_left_inst.comb_out2[6] ),
    .Y(_0948_));
 sg13g2_a21oi_1 _5181_ (.A1(net836),
    .A2(_0947_),
    .Y(_0580_),
    .B1(_0948_));
 sg13g2_nor2_1 _5182_ (.A(net835),
    .B(\u_ddc_top_level.cic_left_inst.comb_out2[5] ),
    .Y(_0949_));
 sg13g2_xor2_1 _5183_ (.B(_0871_),
    .A(_0869_),
    .X(_0950_));
 sg13g2_a21oi_1 _5184_ (.A1(net835),
    .A2(_0950_),
    .Y(_0579_),
    .B1(_0949_));
 sg13g2_nor2_1 _5185_ (.A(net835),
    .B(\u_ddc_top_level.cic_left_inst.comb_out2[4] ),
    .Y(_0951_));
 sg13g2_xnor2_1 _5186_ (.Y(_0952_),
    .A(_0866_),
    .B(_0867_));
 sg13g2_a21oi_1 _5187_ (.A1(net835),
    .A2(_0952_),
    .Y(_0578_),
    .B1(_0951_));
 sg13g2_nor2_1 _5188_ (.A(net832),
    .B(\u_ddc_top_level.cic_left_inst.comb_out2[3] ),
    .Y(_0953_));
 sg13g2_xnor2_1 _5189_ (.Y(_0954_),
    .A(_0857_),
    .B(_0865_));
 sg13g2_a21oi_1 _5190_ (.A1(net831),
    .A2(_0954_),
    .Y(_0577_),
    .B1(_0953_));
 sg13g2_nor2_1 _5191_ (.A(net832),
    .B(\u_ddc_top_level.cic_left_inst.comb_out2[2] ),
    .Y(_0955_));
 sg13g2_xnor2_1 _5192_ (.Y(_0956_),
    .A(_0863_),
    .B(_0864_));
 sg13g2_a21oi_1 _5193_ (.A1(net831),
    .A2(_0956_),
    .Y(_0576_),
    .B1(_0955_));
 sg13g2_xnor2_1 _5194_ (.Y(_0957_),
    .A(_0860_),
    .B(_0862_));
 sg13g2_mux2_1 _5195_ (.A0(\u_ddc_top_level.cic_left_inst.comb_out2[1] ),
    .A1(_0957_),
    .S(net831),
    .X(_0575_));
 sg13g2_nand2b_1 _5196_ (.Y(_0958_),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg2[0] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_out1[0] ));
 sg13g2_nor2_1 _5197_ (.A(net812),
    .B(_0860_),
    .Y(_0959_));
 sg13g2_a22oi_1 _5198_ (.Y(_0574_),
    .B1(_0958_),
    .B2(_0959_),
    .A2(_0732_),
    .A1(net812));
 sg13g2_nand2_1 _5199_ (.Y(_0960_),
    .A(\u_ddc_top_level.cic_left_inst.comb_out1[17] ),
    .B(net809));
 sg13g2_nor2b_1 _5200_ (.A(\u_ddc_top_level.cic_left_inst.comb_reg1[16] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_out0[16] ),
    .Y(_0961_));
 sg13g2_xor2_1 _5201_ (.B(\u_ddc_top_level.cic_left_inst.comb_out0[16] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg1[16] ),
    .X(_0962_));
 sg13g2_nand2b_1 _5202_ (.Y(_0963_),
    .B(\u_ddc_top_level.cic_left_inst.comb_out0[5] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_reg1[5] ));
 sg13g2_nand2b_1 _5203_ (.Y(_0964_),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg1[5] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_out0[5] ));
 sg13g2_nor2b_1 _5204_ (.A(\u_ddc_top_level.cic_left_inst.comb_out0[4] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg1[4] ),
    .Y(_0965_));
 sg13g2_nand2b_1 _5205_ (.Y(_0966_),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg1[3] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_out0[3] ));
 sg13g2_xor2_1 _5206_ (.B(\u_ddc_top_level.cic_left_inst.comb_out0[3] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg1[3] ),
    .X(_0967_));
 sg13g2_nand2b_1 _5207_ (.Y(_0968_),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg1[2] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_out0[2] ));
 sg13g2_nand2b_1 _5208_ (.Y(_0969_),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg1[1] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_out0[1] ));
 sg13g2_nand2b_1 _5209_ (.Y(_0970_),
    .B(\u_ddc_top_level.cic_left_inst.comb_out0[0] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_reg1[0] ));
 sg13g2_xnor2_1 _5210_ (.Y(_0971_),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg1[1] ),
    .B(\u_ddc_top_level.cic_left_inst.comb_out0[1] ));
 sg13g2_nand2_1 _5211_ (.Y(_0972_),
    .A(_0970_),
    .B(_0971_));
 sg13g2_xor2_1 _5212_ (.B(\u_ddc_top_level.cic_left_inst.comb_out0[2] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg1[2] ),
    .X(_0973_));
 sg13g2_a21o_1 _5213_ (.A2(_0972_),
    .A1(_0969_),
    .B1(_0973_),
    .X(_0974_));
 sg13g2_a21o_1 _5214_ (.A2(_0974_),
    .A1(_0968_),
    .B1(_0967_),
    .X(_0975_));
 sg13g2_nand2_1 _5215_ (.Y(_0976_),
    .A(_0966_),
    .B(_0975_));
 sg13g2_xnor2_1 _5216_ (.Y(_0977_),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg1[4] ),
    .B(\u_ddc_top_level.cic_left_inst.comb_out0[4] ));
 sg13g2_a21oi_1 _5217_ (.A1(_0976_),
    .A2(_0977_),
    .Y(_0978_),
    .B1(_0965_));
 sg13g2_nand2_1 _5218_ (.Y(_0979_),
    .A(_0963_),
    .B(_0965_));
 sg13g2_nand2_1 _5219_ (.Y(_0980_),
    .A(_0964_),
    .B(_0979_));
 sg13g2_and2_1 _5220_ (.A(_0963_),
    .B(_0964_),
    .X(_0981_));
 sg13g2_nand2_1 _5221_ (.Y(_0982_),
    .A(_0977_),
    .B(_0981_));
 sg13g2_a21oi_1 _5222_ (.A1(_0966_),
    .A2(_0975_),
    .Y(_0983_),
    .B1(_0982_));
 sg13g2_nor2b_1 _5223_ (.A(\u_ddc_top_level.cic_left_inst.comb_out0[6] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg1[6] ),
    .Y(_0984_));
 sg13g2_xnor2_1 _5224_ (.Y(_0985_),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg1[6] ),
    .B(\u_ddc_top_level.cic_left_inst.comb_out0[6] ));
 sg13g2_o21ai_1 _5225_ (.B1(_0985_),
    .Y(_0986_),
    .A1(_0980_),
    .A2(_0983_));
 sg13g2_a21oi_1 _5226_ (.A1(\u_ddc_top_level.cic_left_inst.comb_reg1[7] ),
    .A2(_0727_),
    .Y(_0987_),
    .B1(_0984_));
 sg13g2_xor2_1 _5227_ (.B(\u_ddc_top_level.cic_left_inst.comb_out0[7] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg1[7] ),
    .X(_0988_));
 sg13g2_a22oi_1 _5228_ (.Y(_0989_),
    .B1(_0986_),
    .B2(_0987_),
    .A2(\u_ddc_top_level.cic_left_inst.comb_out0[7] ),
    .A1(_0726_));
 sg13g2_nand2b_1 _5229_ (.Y(_0990_),
    .B(\u_ddc_top_level.cic_left_inst.comb_out0[9] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_reg1[9] ));
 sg13g2_nor2b_1 _5230_ (.A(\u_ddc_top_level.cic_left_inst.comb_out0[9] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg1[9] ),
    .Y(_0991_));
 sg13g2_xor2_1 _5231_ (.B(\u_ddc_top_level.cic_left_inst.comb_out0[9] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg1[9] ),
    .X(_0992_));
 sg13g2_nor2b_1 _5232_ (.A(\u_ddc_top_level.cic_left_inst.comb_out0[8] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg1[8] ),
    .Y(_0993_));
 sg13g2_nand2b_1 _5233_ (.Y(_0994_),
    .B(\u_ddc_top_level.cic_left_inst.comb_out0[8] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_reg1[8] ));
 sg13g2_nand2b_1 _5234_ (.Y(_0995_),
    .B(_0994_),
    .A_N(_0993_));
 sg13g2_or2_1 _5235_ (.X(_0996_),
    .B(_0995_),
    .A(_0992_));
 sg13g2_a221oi_1 _5236_ (.B2(_0987_),
    .C1(_0996_),
    .B1(_0986_),
    .A1(_0726_),
    .Y(_0997_),
    .A2(\u_ddc_top_level.cic_left_inst.comb_out0[7] ));
 sg13g2_a21o_1 _5237_ (.A2(_0993_),
    .A1(_0990_),
    .B1(_0991_),
    .X(_0998_));
 sg13g2_nor2b_1 _5238_ (.A(\u_ddc_top_level.cic_left_inst.comb_reg1[11] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_out0[11] ),
    .Y(_0999_));
 sg13g2_nand2b_1 _5239_ (.Y(_1000_),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg1[11] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_out0[11] ));
 sg13g2_nor2b_1 _5240_ (.A(\u_ddc_top_level.cic_left_inst.comb_out0[10] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg1[10] ),
    .Y(_1001_));
 sg13g2_inv_1 _5241_ (.Y(_1002_),
    .A(_1001_));
 sg13g2_o21ai_1 _5242_ (.B1(_1000_),
    .Y(_1003_),
    .A1(_0999_),
    .A2(_1002_));
 sg13g2_or2_1 _5243_ (.X(_1004_),
    .B(_1003_),
    .A(_0998_));
 sg13g2_nor2b_1 _5244_ (.A(\u_ddc_top_level.cic_left_inst.comb_reg1[10] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_out0[10] ),
    .Y(_1005_));
 sg13g2_o21ai_1 _5245_ (.B1(_1000_),
    .Y(_1006_),
    .A1(_0999_),
    .A2(_1005_));
 sg13g2_o21ai_1 _5246_ (.B1(_1006_),
    .Y(_1007_),
    .A1(_0997_),
    .A2(_1004_));
 sg13g2_xor2_1 _5247_ (.B(\u_ddc_top_level.cic_left_inst.comb_out0[13] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg1[13] ),
    .X(_1008_));
 sg13g2_nand2b_1 _5248_ (.Y(_1009_),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg1[12] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_out0[12] ));
 sg13g2_xor2_1 _5249_ (.B(\u_ddc_top_level.cic_left_inst.comb_out0[12] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg1[12] ),
    .X(_1010_));
 sg13g2_or2_1 _5250_ (.X(_1011_),
    .B(_1010_),
    .A(_1008_));
 sg13g2_a21oi_1 _5251_ (.A1(_0724_),
    .A2(\u_ddc_top_level.cic_left_inst.comb_out0[13] ),
    .Y(_1012_),
    .B1(_1009_));
 sg13g2_a21oi_1 _5252_ (.A1(\u_ddc_top_level.cic_left_inst.comb_reg1[13] ),
    .A2(_0725_),
    .Y(_1013_),
    .B1(_1012_));
 sg13g2_o21ai_1 _5253_ (.B1(_1013_),
    .Y(_1014_),
    .A1(_1007_),
    .A2(_1011_));
 sg13g2_nor2b_1 _5254_ (.A(\u_ddc_top_level.cic_left_inst.comb_out0[15] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg1[15] ),
    .Y(_1015_));
 sg13g2_nand2b_1 _5255_ (.Y(_1016_),
    .B(\u_ddc_top_level.cic_left_inst.comb_out0[15] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_reg1[15] ));
 sg13g2_nand2b_1 _5256_ (.Y(_1017_),
    .B(_1016_),
    .A_N(_1015_));
 sg13g2_nor2b_1 _5257_ (.A(\u_ddc_top_level.cic_left_inst.comb_out0[14] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg1[14] ),
    .Y(_1018_));
 sg13g2_nand2b_1 _5258_ (.Y(_1019_),
    .B(\u_ddc_top_level.cic_left_inst.comb_out0[14] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_reg1[14] ));
 sg13g2_nand2b_1 _5259_ (.Y(_1020_),
    .B(_1019_),
    .A_N(_1018_));
 sg13g2_nor2_1 _5260_ (.A(_1017_),
    .B(_1020_),
    .Y(_1021_));
 sg13g2_a221oi_1 _5261_ (.B2(_1014_),
    .C1(_1015_),
    .B1(_1021_),
    .A1(_1016_),
    .Y(_1022_),
    .A2(_1018_));
 sg13g2_o21ai_1 _5262_ (.B1(net843),
    .Y(_1023_),
    .A1(_0962_),
    .A2(_1022_));
 sg13g2_o21ai_1 _5263_ (.B1(_0960_),
    .Y(_0573_),
    .A1(_0961_),
    .A2(_1023_));
 sg13g2_nand2_1 _5264_ (.Y(_1024_),
    .A(net809),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[16] ));
 sg13g2_and2_1 _5265_ (.A(_0962_),
    .B(_1022_),
    .X(_1025_));
 sg13g2_o21ai_1 _5266_ (.B1(_1024_),
    .Y(_0572_),
    .A1(_1023_),
    .A2(_1025_));
 sg13g2_a21oi_1 _5267_ (.A1(_1014_),
    .A2(_1019_),
    .Y(_1026_),
    .B1(_1018_));
 sg13g2_nand2_1 _5268_ (.Y(_1027_),
    .A(net808),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[15] ));
 sg13g2_xnor2_1 _5269_ (.Y(_1028_),
    .A(_1017_),
    .B(_1026_));
 sg13g2_o21ai_1 _5270_ (.B1(_1027_),
    .Y(_0571_),
    .A1(net809),
    .A2(_1028_));
 sg13g2_nor2_1 _5271_ (.A(net843),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[14] ),
    .Y(_1029_));
 sg13g2_xor2_1 _5272_ (.B(_1020_),
    .A(_1014_),
    .X(_1030_));
 sg13g2_a21oi_1 _5273_ (.A1(net843),
    .A2(_1030_),
    .Y(_0570_),
    .B1(_1029_));
 sg13g2_o21ai_1 _5274_ (.B1(_1009_),
    .Y(_1031_),
    .A1(_1007_),
    .A2(_1010_));
 sg13g2_o21ai_1 _5275_ (.B1(net840),
    .Y(_1032_),
    .A1(_1008_),
    .A2(_1031_));
 sg13g2_a21oi_1 _5276_ (.A1(_1008_),
    .A2(_1031_),
    .Y(_1033_),
    .B1(_1032_));
 sg13g2_a21oi_1 _5277_ (.A1(net809),
    .A2(_0720_),
    .Y(_0569_),
    .B1(_1033_));
 sg13g2_o21ai_1 _5278_ (.B1(net840),
    .Y(_1034_),
    .A1(_1007_),
    .A2(_1010_));
 sg13g2_a21oi_1 _5279_ (.A1(_1007_),
    .A2(_1010_),
    .Y(_1035_),
    .B1(_1034_));
 sg13g2_a21o_1 _5280_ (.A2(\u_ddc_top_level.cic_left_inst.comb_out1[12] ),
    .A1(net808),
    .B1(_1035_),
    .X(_0568_));
 sg13g2_nand2b_1 _5281_ (.Y(_1036_),
    .B(_1000_),
    .A_N(_0999_));
 sg13g2_nor2_1 _5282_ (.A(_1001_),
    .B(_1005_),
    .Y(_1037_));
 sg13g2_nor2_1 _5283_ (.A(_0997_),
    .B(_0998_),
    .Y(_1038_));
 sg13g2_o21ai_1 _5284_ (.B1(_1002_),
    .Y(_1039_),
    .A1(_1005_),
    .A2(_1038_));
 sg13g2_o21ai_1 _5285_ (.B1(net840),
    .Y(_1040_),
    .A1(_1036_),
    .A2(_1039_));
 sg13g2_a21oi_1 _5286_ (.A1(_1036_),
    .A2(_1039_),
    .Y(_1041_),
    .B1(_1040_));
 sg13g2_a21oi_1 _5287_ (.A1(net808),
    .A2(_0721_),
    .Y(_0567_),
    .B1(_1041_));
 sg13g2_nor2_1 _5288_ (.A(net846),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[10] ),
    .Y(_1042_));
 sg13g2_xor2_1 _5289_ (.B(_1038_),
    .A(_1037_),
    .X(_1043_));
 sg13g2_a21oi_1 _5290_ (.A1(net840),
    .A2(_1043_),
    .Y(_0566_),
    .B1(_1042_));
 sg13g2_a21oi_1 _5291_ (.A1(_0989_),
    .A2(_0994_),
    .Y(_1044_),
    .B1(_0993_));
 sg13g2_nand2_1 _5292_ (.Y(_1045_),
    .A(net808),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[9] ));
 sg13g2_xnor2_1 _5293_ (.Y(_1046_),
    .A(_0992_),
    .B(_1044_));
 sg13g2_o21ai_1 _5294_ (.B1(_1045_),
    .Y(_0565_),
    .A1(net812),
    .A2(_1046_));
 sg13g2_xor2_1 _5295_ (.B(_0995_),
    .A(_0989_),
    .X(_1047_));
 sg13g2_nor2_1 _5296_ (.A(net834),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[8] ),
    .Y(_1048_));
 sg13g2_a21oi_1 _5297_ (.A1(net837),
    .A2(_1047_),
    .Y(_0564_),
    .B1(_1048_));
 sg13g2_nand2b_1 _5298_ (.Y(_1049_),
    .B(_0986_),
    .A_N(_0984_));
 sg13g2_o21ai_1 _5299_ (.B1(net837),
    .Y(_1050_),
    .A1(_0988_),
    .A2(_1049_));
 sg13g2_a21oi_1 _5300_ (.A1(_0988_),
    .A2(_1049_),
    .Y(_1051_),
    .B1(_1050_));
 sg13g2_a21oi_1 _5301_ (.A1(net812),
    .A2(_0722_),
    .Y(_0563_),
    .B1(_1051_));
 sg13g2_nor3_1 _5302_ (.A(_0980_),
    .B(_0983_),
    .C(_0985_),
    .Y(_1052_));
 sg13g2_nand2_1 _5303_ (.Y(_1053_),
    .A(net812),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[6] ));
 sg13g2_nand2_1 _5304_ (.Y(_1054_),
    .A(net834),
    .B(_0986_));
 sg13g2_o21ai_1 _5305_ (.B1(_1053_),
    .Y(_0562_),
    .A1(_1052_),
    .A2(_1054_));
 sg13g2_xnor2_1 _5306_ (.Y(_1055_),
    .A(_0978_),
    .B(_0981_));
 sg13g2_mux2_1 _5307_ (.A0(\u_ddc_top_level.cic_left_inst.comb_out1[5] ),
    .A1(_1055_),
    .S(net834),
    .X(_0561_));
 sg13g2_xnor2_1 _5308_ (.Y(_1056_),
    .A(_0976_),
    .B(_0977_));
 sg13g2_nor2_1 _5309_ (.A(net830),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[4] ),
    .Y(_1057_));
 sg13g2_a21oi_1 _5310_ (.A1(net830),
    .A2(_1056_),
    .Y(_0560_),
    .B1(_1057_));
 sg13g2_nand2_1 _5311_ (.Y(_1058_),
    .A(net812),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[3] ));
 sg13g2_and3_1 _5312_ (.X(_1059_),
    .A(_0967_),
    .B(_0968_),
    .C(_0974_));
 sg13g2_nand2_1 _5313_ (.Y(_1060_),
    .A(net830),
    .B(_0975_));
 sg13g2_o21ai_1 _5314_ (.B1(_1058_),
    .Y(_0559_),
    .A1(_1059_),
    .A2(_1060_));
 sg13g2_nand3_1 _5315_ (.B(_0972_),
    .C(_0973_),
    .A(_0969_),
    .Y(_1061_));
 sg13g2_nand3_1 _5316_ (.B(_0974_),
    .C(_1061_),
    .A(net829),
    .Y(_1062_));
 sg13g2_o21ai_1 _5317_ (.B1(_1062_),
    .Y(_0558_),
    .A1(net830),
    .A2(_0723_));
 sg13g2_nor2_1 _5318_ (.A(net829),
    .B(\u_ddc_top_level.cic_left_inst.comb_out1[1] ),
    .Y(_1063_));
 sg13g2_xnor2_1 _5319_ (.Y(_1064_),
    .A(_0970_),
    .B(_0971_));
 sg13g2_a21oi_1 _5320_ (.A1(net829),
    .A2(_1064_),
    .Y(_0557_),
    .B1(_1063_));
 sg13g2_xor2_1 _5321_ (.B(\u_ddc_top_level.cic_left_inst.comb_out0[0] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg1[0] ),
    .X(_1065_));
 sg13g2_mux2_1 _5322_ (.A0(\u_ddc_top_level.cic_left_inst.comb_out1[0] ),
    .A1(_1065_),
    .S(net829),
    .X(_0556_));
 sg13g2_mux2_1 _5323_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg2[17] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out1[17] ),
    .S(net861),
    .X(_0555_));
 sg13g2_mux2_1 _5324_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg2[16] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out1[16] ),
    .S(net873),
    .X(_0554_));
 sg13g2_mux2_1 _5325_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg2[15] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out1[15] ),
    .S(net873),
    .X(_0553_));
 sg13g2_mux2_1 _5326_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg2[14] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out1[14] ),
    .S(net873),
    .X(_0552_));
 sg13g2_nor2_1 _5327_ (.A(net872),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg2[13] ),
    .Y(_1066_));
 sg13g2_a21oi_1 _5328_ (.A1(net872),
    .A2(_0733_),
    .Y(_0551_),
    .B1(_1066_));
 sg13g2_mux2_1 _5329_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg2[12] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out1[12] ),
    .S(net872),
    .X(_0550_));
 sg13g2_mux2_1 _5330_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg2[11] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out1[11] ),
    .S(net872),
    .X(_0549_));
 sg13g2_mux2_1 _5331_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg2[10] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out1[10] ),
    .S(net872),
    .X(_0548_));
 sg13g2_nor2_1 _5332_ (.A(net866),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg2[9] ),
    .Y(_1067_));
 sg13g2_a21oi_1 _5333_ (.A1(net866),
    .A2(_0734_),
    .Y(_0547_),
    .B1(_1067_));
 sg13g2_mux2_1 _5334_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg2[8] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out1[8] ),
    .S(net866),
    .X(_0546_));
 sg13g2_nor2_1 _5335_ (.A(net866),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg2[7] ),
    .Y(_1068_));
 sg13g2_a21oi_1 _5336_ (.A1(net866),
    .A2(_0735_),
    .Y(_0545_),
    .B1(_1068_));
 sg13g2_mux2_1 _5337_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg2[6] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out1[6] ),
    .S(net866),
    .X(_0544_));
 sg13g2_mux2_1 _5338_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg2[5] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out1[5] ),
    .S(net856),
    .X(_0543_));
 sg13g2_mux2_1 _5339_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg2[4] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out1[4] ),
    .S(net855),
    .X(_0542_));
 sg13g2_mux2_1 _5340_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg2[3] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out1[3] ),
    .S(net854),
    .X(_0541_));
 sg13g2_mux2_1 _5341_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg2[2] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out1[2] ),
    .S(net854),
    .X(_0540_));
 sg13g2_mux2_1 _5342_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg2[1] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out1[1] ),
    .S(net852),
    .X(_0539_));
 sg13g2_nor2_1 _5343_ (.A(net852),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg2[0] ),
    .Y(_1069_));
 sg13g2_a21oi_1 _5344_ (.A1(net852),
    .A2(_0736_),
    .Y(_0538_),
    .B1(_1069_));
 sg13g2_mux2_1 _5345_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg1[16] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out0[16] ),
    .S(net872),
    .X(_0517_));
 sg13g2_mux2_1 _5346_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg1[15] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out0[15] ),
    .S(net876),
    .X(_0516_));
 sg13g2_mux2_1 _5347_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg1[14] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out0[14] ),
    .S(net876),
    .X(_0515_));
 sg13g2_nor2_1 _5348_ (.A(net874),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg1[13] ),
    .Y(_1070_));
 sg13g2_a21oi_1 _5349_ (.A1(net875),
    .A2(_0716_),
    .Y(_0514_),
    .B1(_1070_));
 sg13g2_mux2_1 _5350_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg1[12] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out0[12] ),
    .S(net875),
    .X(_0513_));
 sg13g2_mux2_1 _5351_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg1[11] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out0[11] ),
    .S(net874),
    .X(_0512_));
 sg13g2_nor2_1 _5352_ (.A(net870),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg1[10] ),
    .Y(_1071_));
 sg13g2_a21oi_1 _5353_ (.A1(net870),
    .A2(_0717_),
    .Y(_0511_),
    .B1(_1071_));
 sg13g2_mux2_1 _5354_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg1[9] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out0[9] ),
    .S(net870),
    .X(_0510_));
 sg13g2_mux2_1 _5355_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg1[8] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out0[8] ),
    .S(net867),
    .X(_0509_));
 sg13g2_mux2_1 _5356_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg1[7] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out0[7] ),
    .S(net867),
    .X(_0508_));
 sg13g2_mux2_1 _5357_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg1[6] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out0[6] ),
    .S(net865),
    .X(_0507_));
 sg13g2_mux2_1 _5358_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg1[5] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out0[5] ),
    .S(net865),
    .X(_0506_));
 sg13g2_mux2_1 _5359_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg1[4] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out0[4] ),
    .S(net865),
    .X(_0505_));
 sg13g2_mux2_1 _5360_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg1[3] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out0[3] ),
    .S(net864),
    .X(_0504_));
 sg13g2_mux2_1 _5361_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg1[2] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out0[2] ),
    .S(net854),
    .X(_0503_));
 sg13g2_mux2_1 _5362_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg1[1] ),
    .A1(\u_ddc_top_level.cic_right_inst.comb_out0[1] ),
    .S(net854),
    .X(_0502_));
 sg13g2_nor2_1 _5363_ (.A(net855),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg1[0] ),
    .Y(_1072_));
 sg13g2_a21oi_1 _5364_ (.A1(net854),
    .A2(_0718_),
    .Y(_0501_),
    .B1(_1072_));
 sg13g2_nand2_1 _5365_ (.Y(_1073_),
    .A(net808),
    .B(\u_ddc_top_level.cic_left_inst.comb_out0[16] ));
 sg13g2_nor2b_1 _5366_ (.A(\u_ddc_top_level.cic_left_inst.comb_reg0[15] ),
    .B_N(\u_ddc_top_level.cic_left_inst.in_data[15] ),
    .Y(_1074_));
 sg13g2_xor2_1 _5367_ (.B(\u_ddc_top_level.cic_left_inst.in_data[15] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg0[15] ),
    .X(_1075_));
 sg13g2_nand2b_1 _5368_ (.Y(_1076_),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg0[14] ),
    .A_N(\u_ddc_top_level.cic_left_inst.in_data[14] ));
 sg13g2_xor2_1 _5369_ (.B(\u_ddc_top_level.cic_left_inst.in_data[14] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg0[14] ),
    .X(_1077_));
 sg13g2_inv_1 _5370_ (.Y(_1078_),
    .A(_1077_));
 sg13g2_nand2b_1 _5371_ (.Y(_1079_),
    .B(\u_ddc_top_level.cic_left_inst.in_data[7] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_reg0[7] ));
 sg13g2_nand2b_1 _5372_ (.Y(_1080_),
    .B(\u_ddc_top_level.cic_left_inst.in_data[5] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_reg0[5] ));
 sg13g2_nor2b_1 _5373_ (.A(\u_ddc_top_level.cic_left_inst.in_data[5] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg0[5] ),
    .Y(_1081_));
 sg13g2_nor2b_1 _5374_ (.A(\u_ddc_top_level.cic_left_inst.in_data[4] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg0[4] ),
    .Y(_1082_));
 sg13g2_nand2b_1 _5375_ (.Y(_1083_),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg0[3] ),
    .A_N(\u_ddc_top_level.cic_left_inst.in_data[3] ));
 sg13g2_xor2_1 _5376_ (.B(\u_ddc_top_level.cic_left_inst.in_data[3] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg0[3] ),
    .X(_1084_));
 sg13g2_nor2b_1 _5377_ (.A(\u_ddc_top_level.cic_left_inst.in_data[2] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg0[2] ),
    .Y(_1085_));
 sg13g2_nand2b_1 _5378_ (.Y(_1086_),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg0[1] ),
    .A_N(\u_ddc_top_level.cic_left_inst.in_data[1] ));
 sg13g2_nor2b_1 _5379_ (.A(\u_ddc_top_level.cic_left_inst.comb_reg0[0] ),
    .B_N(\u_ddc_top_level.cic_left_inst.in_data[0] ),
    .Y(_1087_));
 sg13g2_nor2b_1 _5380_ (.A(\u_ddc_top_level.cic_left_inst.comb_reg0[1] ),
    .B_N(\u_ddc_top_level.cic_left_inst.in_data[1] ),
    .Y(_1088_));
 sg13g2_xnor2_1 _5381_ (.Y(_1089_),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg0[1] ),
    .B(\u_ddc_top_level.cic_left_inst.in_data[1] ));
 sg13g2_o21ai_1 _5382_ (.B1(_1086_),
    .Y(_1090_),
    .A1(_1087_),
    .A2(_1088_));
 sg13g2_nand2b_1 _5383_ (.Y(_1091_),
    .B(\u_ddc_top_level.cic_left_inst.in_data[2] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_reg0[2] ));
 sg13g2_nand2b_1 _5384_ (.Y(_1092_),
    .B(_1091_),
    .A_N(_1085_));
 sg13g2_a21oi_1 _5385_ (.A1(_1090_),
    .A2(_1091_),
    .Y(_1093_),
    .B1(_1085_));
 sg13g2_o21ai_1 _5386_ (.B1(_1083_),
    .Y(_1094_),
    .A1(_1084_),
    .A2(_1093_));
 sg13g2_xnor2_1 _5387_ (.Y(_1095_),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg0[4] ),
    .B(\u_ddc_top_level.cic_left_inst.in_data[4] ));
 sg13g2_a21oi_1 _5388_ (.A1(_1094_),
    .A2(_1095_),
    .Y(_1096_),
    .B1(_1082_));
 sg13g2_xnor2_1 _5389_ (.Y(_1097_),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg0[5] ),
    .B(\u_ddc_top_level.cic_left_inst.in_data[5] ));
 sg13g2_and2_1 _5390_ (.A(_1095_),
    .B(_1097_),
    .X(_1098_));
 sg13g2_a221oi_1 _5391_ (.B2(_1098_),
    .C1(_1081_),
    .B1(_1094_),
    .A1(_1080_),
    .Y(_1099_),
    .A2(_1082_));
 sg13g2_nor2b_1 _5392_ (.A(\u_ddc_top_level.cic_left_inst.in_data[6] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg0[6] ),
    .Y(_1100_));
 sg13g2_xor2_1 _5393_ (.B(\u_ddc_top_level.cic_left_inst.in_data[6] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg0[6] ),
    .X(_1101_));
 sg13g2_nor2_1 _5394_ (.A(_1099_),
    .B(_1101_),
    .Y(_1102_));
 sg13g2_nor2b_1 _5395_ (.A(\u_ddc_top_level.cic_left_inst.in_data[7] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg0[7] ),
    .Y(_1103_));
 sg13g2_a21oi_1 _5396_ (.A1(_1079_),
    .A2(_1100_),
    .Y(_1104_),
    .B1(_1103_));
 sg13g2_xnor2_1 _5397_ (.Y(_1105_),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg0[7] ),
    .B(\u_ddc_top_level.cic_left_inst.in_data[7] ));
 sg13g2_nand2b_1 _5398_ (.Y(_1106_),
    .B(_1105_),
    .A_N(_1101_));
 sg13g2_o21ai_1 _5399_ (.B1(_1104_),
    .Y(_1107_),
    .A1(_1099_),
    .A2(_1106_));
 sg13g2_nand2b_1 _5400_ (.Y(_1108_),
    .B(\u_ddc_top_level.cic_left_inst.in_data[9] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_reg0[9] ));
 sg13g2_nor2b_1 _5401_ (.A(\u_ddc_top_level.cic_left_inst.in_data[9] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg0[9] ),
    .Y(_1109_));
 sg13g2_xnor2_1 _5402_ (.Y(_1110_),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg0[9] ),
    .B(\u_ddc_top_level.cic_left_inst.in_data[9] ));
 sg13g2_nor2b_1 _5403_ (.A(\u_ddc_top_level.cic_left_inst.in_data[8] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg0[8] ),
    .Y(_1111_));
 sg13g2_xnor2_1 _5404_ (.Y(_1112_),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg0[8] ),
    .B(\u_ddc_top_level.cic_left_inst.in_data[8] ));
 sg13g2_and2_1 _5405_ (.A(_1110_),
    .B(_1112_),
    .X(_1113_));
 sg13g2_nand2_1 _5406_ (.Y(_1114_),
    .A(_1107_),
    .B(_1113_));
 sg13g2_a21oi_1 _5407_ (.A1(_1108_),
    .A2(_1111_),
    .Y(_1115_),
    .B1(_1109_));
 sg13g2_nand2b_1 _5408_ (.Y(_1116_),
    .B(\u_ddc_top_level.cic_left_inst.in_data[11] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_reg0[11] ));
 sg13g2_nand2b_1 _5409_ (.Y(_1117_),
    .B(\u_ddc_top_level.cic_left_inst.comb_reg0[11] ),
    .A_N(\u_ddc_top_level.cic_left_inst.in_data[11] ));
 sg13g2_nor2b_1 _5410_ (.A(\u_ddc_top_level.cic_left_inst.in_data[10] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg0[10] ),
    .Y(_1118_));
 sg13g2_nand2_1 _5411_ (.Y(_1119_),
    .A(_1116_),
    .B(_1118_));
 sg13g2_and3_1 _5412_ (.X(_1120_),
    .A(_1115_),
    .B(_1117_),
    .C(_1119_));
 sg13g2_inv_1 _5413_ (.Y(_1121_),
    .A(_1120_));
 sg13g2_a21oi_2 _5414_ (.B1(_1121_),
    .Y(_1122_),
    .A2(_1113_),
    .A1(_1107_));
 sg13g2_o21ai_1 _5415_ (.B1(_1116_),
    .Y(_1123_),
    .A1(\u_ddc_top_level.cic_left_inst.comb_reg0[10] ),
    .A2(_0728_));
 sg13g2_and2_1 _5416_ (.A(_1117_),
    .B(_1123_),
    .X(_1124_));
 sg13g2_nor2_1 _5417_ (.A(_1122_),
    .B(_1124_),
    .Y(_1125_));
 sg13g2_or2_1 _5418_ (.X(_1126_),
    .B(_1124_),
    .A(_1122_));
 sg13g2_nor2b_1 _5419_ (.A(\u_ddc_top_level.cic_left_inst.in_data[13] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg0[13] ),
    .Y(_1127_));
 sg13g2_nand2b_1 _5420_ (.Y(_1128_),
    .B(\u_ddc_top_level.cic_left_inst.in_data[13] ),
    .A_N(\u_ddc_top_level.cic_left_inst.comb_reg0[13] ));
 sg13g2_nor2b_1 _5421_ (.A(_1127_),
    .B_N(_1128_),
    .Y(_1129_));
 sg13g2_nor2b_1 _5422_ (.A(\u_ddc_top_level.cic_left_inst.in_data[12] ),
    .B_N(\u_ddc_top_level.cic_left_inst.comb_reg0[12] ),
    .Y(_1130_));
 sg13g2_xor2_1 _5423_ (.B(\u_ddc_top_level.cic_left_inst.in_data[12] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg0[12] ),
    .X(_1131_));
 sg13g2_inv_1 _5424_ (.Y(_1132_),
    .A(_1131_));
 sg13g2_nand2_1 _5425_ (.Y(_1133_),
    .A(_1129_),
    .B(_1132_));
 sg13g2_nor3_1 _5426_ (.A(_1122_),
    .B(_1124_),
    .C(_1133_),
    .Y(_1134_));
 sg13g2_a21oi_1 _5427_ (.A1(_1128_),
    .A2(_1130_),
    .Y(_1135_),
    .B1(_1127_));
 sg13g2_inv_1 _5428_ (.Y(_1136_),
    .A(_1135_));
 sg13g2_nor2_1 _5429_ (.A(_1134_),
    .B(_1136_),
    .Y(_1137_));
 sg13g2_o21ai_1 _5430_ (.B1(_1078_),
    .Y(_1138_),
    .A1(_1134_),
    .A2(_1136_));
 sg13g2_and2_1 _5431_ (.A(_1076_),
    .B(_1138_),
    .X(_1139_));
 sg13g2_o21ai_1 _5432_ (.B1(net842),
    .Y(_1140_),
    .A1(_1075_),
    .A2(_1139_));
 sg13g2_o21ai_1 _5433_ (.B1(_1073_),
    .Y(_0500_),
    .A1(_1074_),
    .A2(_1140_));
 sg13g2_nand2_1 _5434_ (.Y(_1141_),
    .A(net808),
    .B(\u_ddc_top_level.cic_left_inst.comb_out0[15] ));
 sg13g2_and2_1 _5435_ (.A(_1075_),
    .B(_1139_),
    .X(_1142_));
 sg13g2_o21ai_1 _5436_ (.B1(_1141_),
    .Y(_0499_),
    .A1(_1140_),
    .A2(_1142_));
 sg13g2_nor2_1 _5437_ (.A(net842),
    .B(\u_ddc_top_level.cic_left_inst.comb_out0[14] ),
    .Y(_1143_));
 sg13g2_xnor2_1 _5438_ (.Y(_1144_),
    .A(_1077_),
    .B(_1137_));
 sg13g2_a21oi_1 _5439_ (.A1(net842),
    .A2(_1144_),
    .Y(_0498_),
    .B1(_1143_));
 sg13g2_a21oi_1 _5440_ (.A1(_1125_),
    .A2(_1132_),
    .Y(_1145_),
    .B1(_1130_));
 sg13g2_xnor2_1 _5441_ (.Y(_1146_),
    .A(_1129_),
    .B(_1145_));
 sg13g2_nand2_1 _5442_ (.Y(_1147_),
    .A(net839),
    .B(_1146_));
 sg13g2_o21ai_1 _5443_ (.B1(_1147_),
    .Y(_0497_),
    .A1(net839),
    .A2(_0725_));
 sg13g2_o21ai_1 _5444_ (.B1(net839),
    .Y(_1148_),
    .A1(_1126_),
    .A2(_1131_));
 sg13g2_a21oi_1 _5445_ (.A1(_1126_),
    .A2(_1131_),
    .Y(_1149_),
    .B1(_1148_));
 sg13g2_a21o_1 _5446_ (.A2(\u_ddc_top_level.cic_left_inst.comb_out0[12] ),
    .A1(net808),
    .B1(_1149_),
    .X(_0496_));
 sg13g2_nor2_1 _5447_ (.A(net840),
    .B(\u_ddc_top_level.cic_left_inst.comb_out0[11] ),
    .Y(_1150_));
 sg13g2_nand2_1 _5448_ (.Y(_1151_),
    .A(_1116_),
    .B(_1117_));
 sg13g2_xnor2_1 _5449_ (.Y(_1152_),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg0[10] ),
    .B(\u_ddc_top_level.cic_left_inst.in_data[10] ));
 sg13g2_nand2_1 _5450_ (.Y(_1153_),
    .A(_1114_),
    .B(_1115_));
 sg13g2_a21oi_1 _5451_ (.A1(_1152_),
    .A2(_1153_),
    .Y(_1154_),
    .B1(_1118_));
 sg13g2_xnor2_1 _5452_ (.Y(_1155_),
    .A(_1151_),
    .B(_1154_));
 sg13g2_a21oi_1 _5453_ (.A1(net839),
    .A2(_1155_),
    .Y(_0495_),
    .B1(_1150_));
 sg13g2_nor2_1 _5454_ (.A(net840),
    .B(\u_ddc_top_level.cic_left_inst.comb_out0[10] ),
    .Y(_1156_));
 sg13g2_xnor2_1 _5455_ (.Y(_1157_),
    .A(_1152_),
    .B(_1153_));
 sg13g2_a21oi_1 _5456_ (.A1(net839),
    .A2(_1157_),
    .Y(_0494_),
    .B1(_1156_));
 sg13g2_a21oi_1 _5457_ (.A1(_1107_),
    .A2(_1112_),
    .Y(_1158_),
    .B1(_1111_));
 sg13g2_xnor2_1 _5458_ (.Y(_1159_),
    .A(_1110_),
    .B(_1158_));
 sg13g2_mux2_1 _5459_ (.A0(\u_ddc_top_level.cic_left_inst.comb_out0[9] ),
    .A1(_1159_),
    .S(net838),
    .X(_0493_));
 sg13g2_xnor2_1 _5460_ (.Y(_1160_),
    .A(_1107_),
    .B(_1112_));
 sg13g2_nor2_1 _5461_ (.A(net828),
    .B(\u_ddc_top_level.cic_left_inst.comb_out0[8] ),
    .Y(_1161_));
 sg13g2_a21oi_1 _5462_ (.A1(net828),
    .A2(_1160_),
    .Y(_0492_),
    .B1(_1161_));
 sg13g2_nor2_1 _5463_ (.A(_1100_),
    .B(_1102_),
    .Y(_1162_));
 sg13g2_xnor2_1 _5464_ (.Y(_1163_),
    .A(_1105_),
    .B(_1162_));
 sg13g2_nand2_1 _5465_ (.Y(_1164_),
    .A(net827),
    .B(_1163_));
 sg13g2_o21ai_1 _5466_ (.B1(_1164_),
    .Y(_0491_),
    .A1(net827),
    .A2(_0727_));
 sg13g2_o21ai_1 _5467_ (.B1(net828),
    .Y(_1165_),
    .A1(_1099_),
    .A2(_1101_));
 sg13g2_a21oi_1 _5468_ (.A1(_1099_),
    .A2(_1101_),
    .Y(_1166_),
    .B1(_1165_));
 sg13g2_a21o_1 _5469_ (.A2(\u_ddc_top_level.cic_left_inst.comb_out0[6] ),
    .A1(net812),
    .B1(_1166_),
    .X(_0490_));
 sg13g2_nor2_1 _5470_ (.A(net825),
    .B(\u_ddc_top_level.cic_left_inst.comb_out0[5] ),
    .Y(_1167_));
 sg13g2_xor2_1 _5471_ (.B(_1097_),
    .A(_1096_),
    .X(_1168_));
 sg13g2_a21oi_1 _5472_ (.A1(net825),
    .A2(_1168_),
    .Y(_0489_),
    .B1(_1167_));
 sg13g2_nor2_1 _5473_ (.A(net825),
    .B(\u_ddc_top_level.cic_left_inst.comb_out0[4] ),
    .Y(_1169_));
 sg13g2_xnor2_1 _5474_ (.Y(_1170_),
    .A(_1094_),
    .B(_1095_));
 sg13g2_a21oi_1 _5475_ (.A1(net824),
    .A2(_1170_),
    .Y(_0488_),
    .B1(_1169_));
 sg13g2_nor2_1 _5476_ (.A(net824),
    .B(\u_ddc_top_level.cic_left_inst.comb_out0[3] ),
    .Y(_1171_));
 sg13g2_xnor2_1 _5477_ (.Y(_1172_),
    .A(_1084_),
    .B(_1093_));
 sg13g2_a21oi_1 _5478_ (.A1(net825),
    .A2(_1172_),
    .Y(_0487_),
    .B1(_1171_));
 sg13g2_xor2_1 _5479_ (.B(_1092_),
    .A(_1090_),
    .X(_1173_));
 sg13g2_nor2_1 _5480_ (.A(net824),
    .B(\u_ddc_top_level.cic_left_inst.comb_out0[2] ),
    .Y(_1174_));
 sg13g2_a21oi_1 _5481_ (.A1(net824),
    .A2(_1173_),
    .Y(_0486_),
    .B1(_1174_));
 sg13g2_xnor2_1 _5482_ (.Y(_1175_),
    .A(_1087_),
    .B(_1089_));
 sg13g2_mux2_1 _5483_ (.A0(\u_ddc_top_level.cic_left_inst.comb_out0[1] ),
    .A1(_1175_),
    .S(net824),
    .X(_0485_));
 sg13g2_xor2_1 _5484_ (.B(\u_ddc_top_level.cic_left_inst.in_data[0] ),
    .A(\u_ddc_top_level.cic_left_inst.comb_reg0[0] ),
    .X(_1176_));
 sg13g2_mux2_1 _5485_ (.A0(\u_ddc_top_level.cic_left_inst.comb_out0[0] ),
    .A1(_1176_),
    .S(net829),
    .X(_0484_));
 sg13g2_mux2_1 _5486_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg0[15] ),
    .A1(\u_ddc_top_level.cic_right_inst.in_data[15] ),
    .S(net876),
    .X(_0483_));
 sg13g2_mux2_1 _5487_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg0[14] ),
    .A1(\u_ddc_top_level.cic_right_inst.in_data[14] ),
    .S(net876),
    .X(_0482_));
 sg13g2_nor2_1 _5488_ (.A(net876),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg0[13] ),
    .Y(_1177_));
 sg13g2_a21oi_1 _5489_ (.A1(net876),
    .A2(_0739_),
    .Y(_0481_),
    .B1(_1177_));
 sg13g2_mux2_1 _5490_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg0[12] ),
    .A1(\u_ddc_top_level.cic_right_inst.in_data[12] ),
    .S(net875),
    .X(_0480_));
 sg13g2_mux2_1 _5491_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg0[11] ),
    .A1(\u_ddc_top_level.cic_right_inst.in_data[11] ),
    .S(net877),
    .X(_0479_));
 sg13g2_mux2_1 _5492_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg0[10] ),
    .A1(\u_ddc_top_level.cic_right_inst.in_data[10] ),
    .S(net875),
    .X(_0478_));
 sg13g2_mux2_1 _5493_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg0[9] ),
    .A1(\u_ddc_top_level.cic_right_inst.in_data[9] ),
    .S(net871),
    .X(_0477_));
 sg13g2_mux2_1 _5494_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg0[8] ),
    .A1(\u_ddc_top_level.cic_right_inst.in_data[8] ),
    .S(net870),
    .X(_0476_));
 sg13g2_mux2_1 _5495_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg0[7] ),
    .A1(\u_ddc_top_level.cic_right_inst.in_data[7] ),
    .S(net871),
    .X(_0475_));
 sg13g2_mux2_1 _5496_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg0[6] ),
    .A1(\u_ddc_top_level.cic_right_inst.in_data[6] ),
    .S(net871),
    .X(_0474_));
 sg13g2_mux2_1 _5497_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg0[5] ),
    .A1(\u_ddc_top_level.cic_right_inst.in_data[5] ),
    .S(net869),
    .X(_0473_));
 sg13g2_mux2_1 _5498_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg0[4] ),
    .A1(\u_ddc_top_level.cic_right_inst.in_data[4] ),
    .S(net869),
    .X(_0472_));
 sg13g2_mux2_1 _5499_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg0[3] ),
    .A1(\u_ddc_top_level.cic_right_inst.in_data[3] ),
    .S(net869),
    .X(_0471_));
 sg13g2_mux2_1 _5500_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg0[2] ),
    .A1(\u_ddc_top_level.cic_right_inst.in_data[2] ),
    .S(net864),
    .X(_0470_));
 sg13g2_mux2_1 _5501_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg0[1] ),
    .A1(\u_ddc_top_level.cic_right_inst.in_data[1] ),
    .S(net864),
    .X(_0469_));
 sg13g2_mux2_1 _5502_ (.A0(\u_ddc_top_level.cic_right_inst.comb_reg0[0] ),
    .A1(\u_ddc_top_level.cic_right_inst.in_data[0] ),
    .S(net864),
    .X(_0468_));
 sg13g2_nand2b_1 _5503_ (.Y(_1178_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg2[17] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_out1[17] ));
 sg13g2_xnor2_1 _5504_ (.Y(_1179_),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg2[17] ),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[17] ));
 sg13g2_nand2b_1 _5505_ (.Y(_1180_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg2[16] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_out1[16] ));
 sg13g2_nor2_1 _5506_ (.A(\u_ddc_top_level.cic_right_inst.comb_reg2[7] ),
    .B(_0735_),
    .Y(_1181_));
 sg13g2_nand2b_1 _5507_ (.Y(_1182_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg2[6] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_out1[6] ));
 sg13g2_inv_1 _5508_ (.Y(_1183_),
    .A(_1182_));
 sg13g2_nand2b_1 _5509_ (.Y(_1184_),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[6] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_reg2[6] ));
 sg13g2_nand2b_1 _5510_ (.Y(_1185_),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[5] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_reg2[5] ));
 sg13g2_nand2b_1 _5511_ (.Y(_1186_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg2[5] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_out1[5] ));
 sg13g2_nand2b_1 _5512_ (.Y(_1187_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg2[4] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_out1[4] ));
 sg13g2_nor2b_1 _5513_ (.A(\u_ddc_top_level.cic_right_inst.comb_out1[3] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg2[3] ),
    .Y(_1188_));
 sg13g2_xnor2_1 _5514_ (.Y(_1189_),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg2[3] ),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[3] ));
 sg13g2_nor2b_1 _5515_ (.A(\u_ddc_top_level.cic_right_inst.comb_out1[2] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg2[2] ),
    .Y(_1190_));
 sg13g2_nand2b_1 _5516_ (.Y(_1191_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg2[1] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_out1[1] ));
 sg13g2_nor2b_1 _5517_ (.A(\u_ddc_top_level.cic_right_inst.comb_reg2[0] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_out1[0] ),
    .Y(_1192_));
 sg13g2_nor2b_1 _5518_ (.A(\u_ddc_top_level.cic_right_inst.comb_reg2[1] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_out1[1] ),
    .Y(_1193_));
 sg13g2_xnor2_1 _5519_ (.Y(_1194_),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg2[1] ),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[1] ));
 sg13g2_o21ai_1 _5520_ (.B1(_1191_),
    .Y(_1195_),
    .A1(_1192_),
    .A2(_1193_));
 sg13g2_xnor2_1 _5521_ (.Y(_1196_),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg2[2] ),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[2] ));
 sg13g2_a21o_1 _5522_ (.A2(_1196_),
    .A1(_1195_),
    .B1(_1190_),
    .X(_1197_));
 sg13g2_a21oi_2 _5523_ (.B1(_1188_),
    .Y(_1198_),
    .A2(_1197_),
    .A1(_1189_));
 sg13g2_xnor2_1 _5524_ (.Y(_1199_),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg2[4] ),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[4] ));
 sg13g2_nand2b_1 _5525_ (.Y(_1200_),
    .B(_1199_),
    .A_N(_1198_));
 sg13g2_nand2_1 _5526_ (.Y(_1201_),
    .A(_1187_),
    .B(_1200_));
 sg13g2_nand2b_1 _5527_ (.Y(_1202_),
    .B(_1185_),
    .A_N(_1187_));
 sg13g2_and2_1 _5528_ (.A(_1186_),
    .B(_1202_),
    .X(_1203_));
 sg13g2_nand2_1 _5529_ (.Y(_1204_),
    .A(_1185_),
    .B(_1186_));
 sg13g2_nand3_1 _5530_ (.B(_1186_),
    .C(_1199_),
    .A(_1185_),
    .Y(_1205_));
 sg13g2_o21ai_1 _5531_ (.B1(_1203_),
    .Y(_1206_),
    .A1(_1198_),
    .A2(_1205_));
 sg13g2_nand3_1 _5532_ (.B(_1184_),
    .C(_1206_),
    .A(_1182_),
    .Y(_1207_));
 sg13g2_nand2_1 _5533_ (.Y(_1208_),
    .A(_1182_),
    .B(_1207_));
 sg13g2_a221oi_1 _5534_ (.B2(_1206_),
    .C1(_1183_),
    .B1(_1184_),
    .A1(\u_ddc_top_level.cic_right_inst.comb_reg2[7] ),
    .Y(_1209_),
    .A2(_0735_));
 sg13g2_nor2_1 _5535_ (.A(_1181_),
    .B(_1209_),
    .Y(_1210_));
 sg13g2_nor2b_1 _5536_ (.A(\u_ddc_top_level.cic_right_inst.comb_out1[11] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg2[11] ),
    .Y(_1211_));
 sg13g2_nand2b_1 _5537_ (.Y(_1212_),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[11] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_reg2[11] ));
 sg13g2_nand2b_1 _5538_ (.Y(_1213_),
    .B(_1212_),
    .A_N(_1211_));
 sg13g2_nor2b_1 _5539_ (.A(\u_ddc_top_level.cic_right_inst.comb_out1[10] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg2[10] ),
    .Y(_1214_));
 sg13g2_nand2b_1 _5540_ (.Y(_1215_),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[10] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_reg2[10] ));
 sg13g2_nand2b_1 _5541_ (.Y(_1216_),
    .B(_1215_),
    .A_N(_1214_));
 sg13g2_nor2_1 _5542_ (.A(_1213_),
    .B(_1216_),
    .Y(_1217_));
 sg13g2_nand2_1 _5543_ (.Y(_1218_),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg2[9] ),
    .B(_0734_));
 sg13g2_nor2_1 _5544_ (.A(\u_ddc_top_level.cic_right_inst.comb_reg2[9] ),
    .B(_0734_),
    .Y(_1219_));
 sg13g2_xnor2_1 _5545_ (.Y(_1220_),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg2[9] ),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[9] ));
 sg13g2_nor2b_1 _5546_ (.A(\u_ddc_top_level.cic_right_inst.comb_out1[8] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg2[8] ),
    .Y(_1221_));
 sg13g2_nand2b_1 _5547_ (.Y(_1222_),
    .B(\u_ddc_top_level.cic_right_inst.comb_reg2[8] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_out1[8] ));
 sg13g2_xnor2_1 _5548_ (.Y(_1223_),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg2[8] ),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[8] ));
 sg13g2_nand3_1 _5549_ (.B(_1220_),
    .C(_1223_),
    .A(_1217_),
    .Y(_1224_));
 sg13g2_nor3_2 _5550_ (.A(_1181_),
    .B(_1209_),
    .C(_1224_),
    .Y(_1225_));
 sg13g2_a21oi_1 _5551_ (.A1(_1212_),
    .A2(_1214_),
    .Y(_1226_),
    .B1(_1211_));
 sg13g2_o21ai_1 _5552_ (.B1(_1218_),
    .Y(_1227_),
    .A1(_1219_),
    .A2(_1222_));
 sg13g2_nand2_1 _5553_ (.Y(_1228_),
    .A(_1217_),
    .B(_1227_));
 sg13g2_nand2_1 _5554_ (.Y(_1229_),
    .A(_1226_),
    .B(_1228_));
 sg13g2_nor2_2 _5555_ (.A(_1225_),
    .B(_1229_),
    .Y(_1230_));
 sg13g2_nor2b_1 _5556_ (.A(\u_ddc_top_level.cic_right_inst.comb_out1[15] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg2[15] ),
    .Y(_1231_));
 sg13g2_nand2b_1 _5557_ (.Y(_1232_),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[15] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_reg2[15] ));
 sg13g2_nand2b_1 _5558_ (.Y(_1233_),
    .B(_1232_),
    .A_N(_1231_));
 sg13g2_nor2b_1 _5559_ (.A(\u_ddc_top_level.cic_right_inst.comb_out1[14] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg2[14] ),
    .Y(_1234_));
 sg13g2_nand2b_1 _5560_ (.Y(_1235_),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[14] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_reg2[14] ));
 sg13g2_nand2b_1 _5561_ (.Y(_1236_),
    .B(_1235_),
    .A_N(_1234_));
 sg13g2_nor2_1 _5562_ (.A(_1233_),
    .B(_1236_),
    .Y(_1237_));
 sg13g2_nor2b_1 _5563_ (.A(\u_ddc_top_level.cic_right_inst.comb_out1[13] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg2[13] ),
    .Y(_1238_));
 sg13g2_nand2b_1 _5564_ (.Y(_1239_),
    .B(\u_ddc_top_level.cic_right_inst.comb_out1[13] ),
    .A_N(\u_ddc_top_level.cic_right_inst.comb_reg2[13] ));
 sg13g2_nand2b_1 _5565_ (.Y(_1240_),
    .B(_1239_),
    .A_N(_1238_));
 sg13g2_nor2b_1 _5566_ (.A(\u_ddc_top_level.cic_right_inst.comb_out1[12] ),
    .B_N(\u_ddc_top_level.cic_right_inst.comb_reg2[12] ),
    .Y(_1241_));
 sg13g2_xor2_1 _5567_ (.B(\u_ddc_top_level.cic_right_inst.comb_out1[12] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg2[12] ),
    .X(_1242_));
 sg13g2_nor2_1 _5568_ (.A(_1240_),
    .B(_1242_),
    .Y(_1243_));
 sg13g2_inv_1 _5569_ (.Y(_1244_),
    .A(_1243_));
 sg13g2_and2_1 _5570_ (.A(_1237_),
    .B(_1243_),
    .X(_1245_));
 sg13g2_o21ai_1 _5571_ (.B1(_1245_),
    .Y(_1246_),
    .A1(_1225_),
    .A2(_1229_));
 sg13g2_a21oi_1 _5572_ (.A1(_1239_),
    .A2(_1241_),
    .Y(_1247_),
    .B1(_1238_));
 sg13g2_inv_1 _5573_ (.Y(_1248_),
    .A(_1247_));
 sg13g2_a221oi_1 _5574_ (.B2(_1248_),
    .C1(_1231_),
    .B1(_1237_),
    .A1(_1232_),
    .Y(_1249_),
    .A2(_1234_));
 sg13g2_xor2_1 _5575_ (.B(\u_ddc_top_level.cic_right_inst.comb_out1[16] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg2[16] ),
    .X(_1250_));
 sg13g2_a21o_1 _5576_ (.A2(_1249_),
    .A1(_1246_),
    .B1(_1250_),
    .X(_1251_));
 sg13g2_nand3_1 _5577_ (.B(_1180_),
    .C(_1251_),
    .A(_1179_),
    .Y(_1252_));
 sg13g2_and2_1 _5578_ (.A(net861),
    .B(_1252_),
    .X(_1253_));
 sg13g2_a22oi_1 _5579_ (.Y(_0467_),
    .B1(_1178_),
    .B2(_1253_),
    .A2(_0740_),
    .A1(net817));
 sg13g2_a21o_1 _5580_ (.A2(_1251_),
    .A1(_1180_),
    .B1(_1179_),
    .X(_1254_));
 sg13g2_a22oi_1 _5581_ (.Y(_0466_),
    .B1(_1253_),
    .B2(_1254_),
    .A2(_0741_),
    .A1(net817));
 sg13g2_nand3_1 _5582_ (.B(_1249_),
    .C(_1250_),
    .A(_1246_),
    .Y(_1255_));
 sg13g2_a21oi_1 _5583_ (.A1(_1251_),
    .A2(_1255_),
    .Y(_1256_),
    .B1(net815));
 sg13g2_a21oi_1 _5584_ (.A1(net815),
    .A2(_0742_),
    .Y(_0465_),
    .B1(_1256_));
 sg13g2_o21ai_1 _5585_ (.B1(_1247_),
    .Y(_1257_),
    .A1(_1230_),
    .A2(_1244_));
 sg13g2_a21oi_1 _5586_ (.A1(_1235_),
    .A2(_1257_),
    .Y(_1258_),
    .B1(_1234_));
 sg13g2_nand2_1 _5587_ (.Y(_1259_),
    .A(net815),
    .B(\u_ddc_top_level.cic_right_inst.comb_out2[15] ));
 sg13g2_xnor2_1 _5588_ (.Y(_1260_),
    .A(_1233_),
    .B(_1258_));
 sg13g2_o21ai_1 _5589_ (.B1(_1259_),
    .Y(_0464_),
    .A1(net815),
    .A2(_1260_));
 sg13g2_nor2_1 _5590_ (.A(net861),
    .B(\u_ddc_top_level.cic_right_inst.comb_out2[14] ),
    .Y(_1261_));
 sg13g2_xor2_1 _5591_ (.B(_1257_),
    .A(_1236_),
    .X(_1262_));
 sg13g2_a21oi_1 _5592_ (.A1(net862),
    .A2(_1262_),
    .Y(_0463_),
    .B1(_1261_));
 sg13g2_nor2_1 _5593_ (.A(_1230_),
    .B(_1242_),
    .Y(_1263_));
 sg13g2_nor2_1 _5594_ (.A(_1241_),
    .B(_1263_),
    .Y(_1264_));
 sg13g2_nor2_1 _5595_ (.A(net860),
    .B(\u_ddc_top_level.cic_right_inst.comb_out2[13] ),
    .Y(_1265_));
 sg13g2_xnor2_1 _5596_ (.Y(_1266_),
    .A(_1240_),
    .B(_1264_));
 sg13g2_a21oi_1 _5597_ (.A1(net860),
    .A2(_1266_),
    .Y(_0462_),
    .B1(_1265_));
 sg13g2_o21ai_1 _5598_ (.B1(net872),
    .Y(_1267_),
    .A1(_1230_),
    .A2(_1242_));
 sg13g2_a21oi_1 _5599_ (.A1(_1230_),
    .A2(_1242_),
    .Y(_1268_),
    .B1(_1267_));
 sg13g2_a21o_1 _5600_ (.A2(\u_ddc_top_level.cic_right_inst.comb_out2[12] ),
    .A1(net817),
    .B1(_1268_),
    .X(_0461_));
 sg13g2_a21oi_1 _5601_ (.A1(_1210_),
    .A2(_1223_),
    .Y(_1269_),
    .B1(_1221_));
 sg13g2_o21ai_1 _5602_ (.B1(_1218_),
    .Y(_1270_),
    .A1(_1219_),
    .A2(_1269_));
 sg13g2_a21oi_1 _5603_ (.A1(_1215_),
    .A2(_1270_),
    .Y(_1271_),
    .B1(_1214_));
 sg13g2_xnor2_1 _5604_ (.Y(_1272_),
    .A(_1213_),
    .B(_1271_));
 sg13g2_nor2_1 _5605_ (.A(net860),
    .B(\u_ddc_top_level.cic_right_inst.comb_out2[11] ),
    .Y(_1273_));
 sg13g2_a21oi_1 _5606_ (.A1(net860),
    .A2(_1272_),
    .Y(_0460_),
    .B1(_1273_));
 sg13g2_xnor2_1 _5607_ (.Y(_1274_),
    .A(_1216_),
    .B(_1270_));
 sg13g2_mux2_1 _5608_ (.A0(\u_ddc_top_level.cic_right_inst.comb_out2[10] ),
    .A1(_1274_),
    .S(net860),
    .X(_0459_));
 sg13g2_xnor2_1 _5609_ (.Y(_1275_),
    .A(_1220_),
    .B(_1269_));
 sg13g2_mux2_1 _5610_ (.A0(\u_ddc_top_level.cic_right_inst.comb_out2[9] ),
    .A1(_1275_),
    .S(net861),
    .X(_0458_));
 sg13g2_xnor2_1 _5611_ (.Y(_1276_),
    .A(_1210_),
    .B(_1223_));
 sg13g2_nor2_1 _5612_ (.A(net861),
    .B(\u_ddc_top_level.cic_right_inst.comb_out2[8] ),
    .Y(_1277_));
 sg13g2_a21oi_1 _5613_ (.A1(net860),
    .A2(_1276_),
    .Y(_0457_),
    .B1(_1277_));
 sg13g2_xor2_1 _5614_ (.B(\u_ddc_top_level.cic_right_inst.comb_out1[7] ),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg2[7] ),
    .X(_1278_));
 sg13g2_xnor2_1 _5615_ (.Y(_1279_),
    .A(_1208_),
    .B(_1278_));
 sg13g2_mux2_1 _5616_ (.A0(\u_ddc_top_level.cic_right_inst.comb_out2[7] ),
    .A1(_1279_),
    .S(net857),
    .X(_0456_));
 sg13g2_a21oi_1 _5617_ (.A1(_1182_),
    .A2(_1184_),
    .Y(_1280_),
    .B1(_1206_));
 sg13g2_nand2_1 _5618_ (.Y(_1281_),
    .A(net813),
    .B(\u_ddc_top_level.cic_right_inst.comb_out2[6] ));
 sg13g2_nand2_1 _5619_ (.Y(_1282_),
    .A(net856),
    .B(_1207_));
 sg13g2_o21ai_1 _5620_ (.B1(_1281_),
    .Y(_0455_),
    .A1(_1280_),
    .A2(_1282_));
 sg13g2_nor2_1 _5621_ (.A(net856),
    .B(\u_ddc_top_level.cic_right_inst.comb_out2[5] ),
    .Y(_1283_));
 sg13g2_xor2_1 _5622_ (.B(_1204_),
    .A(_1201_),
    .X(_1284_));
 sg13g2_a21oi_1 _5623_ (.A1(net857),
    .A2(_1284_),
    .Y(_0454_),
    .B1(_1283_));
 sg13g2_xnor2_1 _5624_ (.Y(_1285_),
    .A(_1198_),
    .B(_1199_));
 sg13g2_mux2_1 _5625_ (.A0(\u_ddc_top_level.cic_right_inst.comb_out2[4] ),
    .A1(_1285_),
    .S(net856),
    .X(_0453_));
 sg13g2_nor2_1 _5626_ (.A(net856),
    .B(\u_ddc_top_level.cic_right_inst.comb_out2[3] ),
    .Y(_1286_));
 sg13g2_xnor2_1 _5627_ (.Y(_1287_),
    .A(_1189_),
    .B(_1197_));
 sg13g2_a21oi_1 _5628_ (.A1(net854),
    .A2(_1287_),
    .Y(_0452_),
    .B1(_1286_));
 sg13g2_nor2_1 _5629_ (.A(net853),
    .B(\u_ddc_top_level.cic_right_inst.comb_out2[2] ),
    .Y(_1288_));
 sg13g2_xnor2_1 _5630_ (.Y(_1289_),
    .A(_1195_),
    .B(_1196_));
 sg13g2_a21oi_1 _5631_ (.A1(net852),
    .A2(_1289_),
    .Y(_0451_),
    .B1(_1288_));
 sg13g2_xnor2_1 _5632_ (.Y(_1290_),
    .A(_1192_),
    .B(_1194_));
 sg13g2_mux2_1 _5633_ (.A0(\u_ddc_top_level.cic_right_inst.comb_out2[1] ),
    .A1(_1290_),
    .S(net852),
    .X(_0450_));
 sg13g2_nand2_1 _5634_ (.Y(_1291_),
    .A(\u_ddc_top_level.cic_right_inst.comb_reg2[0] ),
    .B(_0736_));
 sg13g2_nor2_1 _5635_ (.A(net813),
    .B(_1192_),
    .Y(_1292_));
 sg13g2_dfrbp_1 _5636_ (.CLK(net925),
    .RESET_B(net1012),
    .D(_0398_),
    .Q_N(\u_ddc_top_level.lsfr_inst.lfsr_reg[0] ),
    .Q(_0111_));
 sg13g2_dfrbp_1 _5637_ (.CLK(net925),
    .RESET_B(net1012),
    .D(_0399_),
    .Q_N(_2883_),
    .Q(\u_ddc_top_level.lsfr_inst.lfsr_reg[1] ));
 sg13g2_dfrbp_1 _5638_ (.CLK(net925),
    .RESET_B(net1012),
    .D(_0400_),
    .Q_N(_2882_),
    .Q(\u_ddc_top_level.lsfr_inst.lfsr_reg[2] ));
 sg13g2_dfrbp_1 _5639_ (.CLK(net925),
    .RESET_B(net1012),
    .D(_0401_),
    .Q_N(_2881_),
    .Q(\u_ddc_top_level.lsfr_inst.lfsr_reg[3] ));
 sg13g2_dfrbp_1 _5640_ (.CLK(net925),
    .RESET_B(net1012),
    .D(_0402_),
    .Q_N(_2880_),
    .Q(\u_ddc_top_level.lsfr_inst.lfsr_reg[4] ));
 sg13g2_dfrbp_1 _5641_ (.CLK(net925),
    .RESET_B(net1012),
    .D(_0403_),
    .Q_N(_2879_),
    .Q(\u_ddc_top_level.lsfr_inst.lfsr_reg[5] ));
 sg13g2_dfrbp_1 _5642_ (.CLK(net927),
    .RESET_B(net1015),
    .D(_0404_),
    .Q_N(_2878_),
    .Q(\u_ddc_top_level.lsfr_inst.lfsr_reg[6] ));
 sg13g2_dfrbp_1 _5643_ (.CLK(net927),
    .RESET_B(net1014),
    .D(_0405_),
    .Q_N(_2877_),
    .Q(\u_ddc_top_level.lsfr_inst.lfsr_reg[7] ));
 sg13g2_dfrbp_1 _5644_ (.CLK(net927),
    .RESET_B(net1014),
    .D(_0406_),
    .Q_N(_2876_),
    .Q(\u_ddc_top_level.lsfr_inst.lfsr_reg[8] ));
 sg13g2_dfrbp_1 _5645_ (.CLK(net927),
    .RESET_B(net1014),
    .D(_0407_),
    .Q_N(_2875_),
    .Q(\u_ddc_top_level.lsfr_inst.lfsr_reg[9] ));
 sg13g2_dfrbp_1 _5646_ (.CLK(net926),
    .RESET_B(net1014),
    .D(_0408_),
    .Q_N(_2874_),
    .Q(\u_ddc_top_level.lsfr_inst.lfsr_reg[10] ));
 sg13g2_dfrbp_1 _5647_ (.CLK(net926),
    .RESET_B(net1013),
    .D(_0409_),
    .Q_N(_2873_),
    .Q(\u_ddc_top_level.lsfr_inst.lfsr_reg[11] ));
 sg13g2_dfrbp_1 _5648_ (.CLK(net925),
    .RESET_B(net1013),
    .D(_0410_),
    .Q_N(_2872_),
    .Q(\u_ddc_top_level.lsfr_inst.lfsr_reg[12] ));
 sg13g2_dfrbp_1 _5649_ (.CLK(net926),
    .RESET_B(net1013),
    .D(_0411_),
    .Q_N(_2871_),
    .Q(\u_ddc_top_level.lsfr_inst.lfsr_reg[13] ));
 sg13g2_dfrbp_1 _5650_ (.CLK(net926),
    .RESET_B(net1012),
    .D(_0412_),
    .Q_N(_2870_),
    .Q(\u_ddc_top_level.lsfr_inst.lfsr_reg[14] ));
 sg13g2_dfrbp_1 _5651_ (.CLK(net926),
    .RESET_B(net1013),
    .D(_0413_),
    .Q_N(_2869_),
    .Q(\u_ddc_top_level.lsfr_inst.lfsr_reg[15] ));
 sg13g2_dfrbp_1 _5652_ (.CLK(net925),
    .RESET_B(net1012),
    .D(_0414_),
    .Q_N(_0006_),
    .Q(\u_ddc_top_level.dsm_left_inst.in_dither ));
 sg13g2_dfrbp_1 _5653_ (.CLK(net900),
    .RESET_B(net987),
    .D(_0415_),
    .Q_N(_2868_),
    .Q(\u_ddc_top_level.i2s_rx_inst.shift_reg[0] ));
 sg13g2_dfrbp_1 _5654_ (.CLK(net929),
    .RESET_B(net1017),
    .D(_0416_),
    .Q_N(_2867_),
    .Q(\u_ddc_top_level.i2s_rx_inst.shift_reg[1] ));
 sg13g2_dfrbp_1 _5655_ (.CLK(net929),
    .RESET_B(net1017),
    .D(_0417_),
    .Q_N(_2866_),
    .Q(\u_ddc_top_level.i2s_rx_inst.shift_reg[2] ));
 sg13g2_dfrbp_1 _5656_ (.CLK(net929),
    .RESET_B(net1017),
    .D(_0418_),
    .Q_N(_2865_),
    .Q(\u_ddc_top_level.i2s_rx_inst.shift_reg[3] ));
 sg13g2_dfrbp_1 _5657_ (.CLK(net929),
    .RESET_B(net1017),
    .D(_0419_),
    .Q_N(_2864_),
    .Q(\u_ddc_top_level.i2s_rx_inst.shift_reg[4] ));
 sg13g2_dfrbp_1 _5658_ (.CLK(net931),
    .RESET_B(net1019),
    .D(_0420_),
    .Q_N(_2863_),
    .Q(\u_ddc_top_level.i2s_rx_inst.shift_reg[5] ));
 sg13g2_dfrbp_1 _5659_ (.CLK(net931),
    .RESET_B(net1022),
    .D(_0421_),
    .Q_N(_2862_),
    .Q(\u_ddc_top_level.i2s_rx_inst.shift_reg[6] ));
 sg13g2_dfrbp_1 _5660_ (.CLK(net931),
    .RESET_B(net1022),
    .D(_0422_),
    .Q_N(_2861_),
    .Q(\u_ddc_top_level.i2s_rx_inst.shift_reg[7] ));
 sg13g2_dfrbp_1 _5661_ (.CLK(net936),
    .RESET_B(net1023),
    .D(_0423_),
    .Q_N(_2860_),
    .Q(\u_ddc_top_level.i2s_rx_inst.shift_reg[8] ));
 sg13g2_dfrbp_1 _5662_ (.CLK(net936),
    .RESET_B(net1023),
    .D(_0424_),
    .Q_N(_2859_),
    .Q(\u_ddc_top_level.i2s_rx_inst.shift_reg[9] ));
 sg13g2_dfrbp_1 _5663_ (.CLK(net936),
    .RESET_B(net1024),
    .D(_0425_),
    .Q_N(_2858_),
    .Q(\u_ddc_top_level.i2s_rx_inst.shift_reg[10] ));
 sg13g2_dfrbp_1 _5664_ (.CLK(net937),
    .RESET_B(net1024),
    .D(_0426_),
    .Q_N(_2857_),
    .Q(\u_ddc_top_level.i2s_rx_inst.shift_reg[11] ));
 sg13g2_dfrbp_1 _5665_ (.CLK(net937),
    .RESET_B(net1024),
    .D(_0427_),
    .Q_N(_2856_),
    .Q(\u_ddc_top_level.i2s_rx_inst.shift_reg[12] ));
 sg13g2_dfrbp_1 _5666_ (.CLK(net920),
    .RESET_B(net1007),
    .D(_0428_),
    .Q_N(_2855_),
    .Q(\u_ddc_top_level.i2s_rx_inst.shift_reg[13] ));
 sg13g2_dfrbp_1 _5667_ (.CLK(net920),
    .RESET_B(net1007),
    .D(_0429_),
    .Q_N(_2854_),
    .Q(\u_ddc_top_level.i2s_rx_inst.shift_reg[14] ));
 sg13g2_dfrbp_1 _5668_ (.CLK(net953),
    .RESET_B(net1041),
    .D(_0430_),
    .Q_N(_2884_),
    .Q(\u_ddc_top_level.i2s_rx_inst.shift_reg[15] ));
 sg13g2_dfrbp_1 _5669_ (.CLK(net921),
    .RESET_B(net1008),
    .D(_0112_),
    .Q_N(_2885_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator2[0] ));
 sg13g2_dfrbp_1 _5670_ (.CLK(net918),
    .RESET_B(net1006),
    .D(_0122_),
    .Q_N(_2886_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator2[1] ));
 sg13g2_dfrbp_1 _5671_ (.CLK(net918),
    .RESET_B(net1005),
    .D(_0123_),
    .Q_N(_2887_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator2[2] ));
 sg13g2_dfrbp_1 _5672_ (.CLK(net918),
    .RESET_B(net1005),
    .D(_0124_),
    .Q_N(_2888_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator2[3] ));
 sg13g2_dfrbp_1 _5673_ (.CLK(net913),
    .RESET_B(net998),
    .D(_0125_),
    .Q_N(_2889_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator2[4] ));
 sg13g2_dfrbp_1 _5674_ (.CLK(net916),
    .RESET_B(net1002),
    .D(_0126_),
    .Q_N(_2890_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator2[5] ));
 sg13g2_dfrbp_1 _5675_ (.CLK(net924),
    .RESET_B(net1011),
    .D(_0127_),
    .Q_N(_2891_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator2[6] ));
 sg13g2_dfrbp_1 _5676_ (.CLK(net924),
    .RESET_B(net1011),
    .D(_0128_),
    .Q_N(_2892_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator2[7] ));
 sg13g2_dfrbp_1 _5677_ (.CLK(net916),
    .RESET_B(net1002),
    .D(_0129_),
    .Q_N(_2893_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator2[8] ));
 sg13g2_dfrbp_1 _5678_ (.CLK(net916),
    .RESET_B(net1002),
    .D(_0130_),
    .Q_N(_2894_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator2[9] ));
 sg13g2_dfrbp_1 _5679_ (.CLK(net916),
    .RESET_B(net1001),
    .D(_0113_),
    .Q_N(_2895_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator2[10] ));
 sg13g2_dfrbp_1 _5680_ (.CLK(net915),
    .RESET_B(net1001),
    .D(_0114_),
    .Q_N(_2896_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator2[11] ));
 sg13g2_dfrbp_1 _5681_ (.CLK(net924),
    .RESET_B(net1011),
    .D(_0115_),
    .Q_N(_2897_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator2[12] ));
 sg13g2_dfrbp_1 _5682_ (.CLK(net924),
    .RESET_B(net1011),
    .D(_0116_),
    .Q_N(_2898_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator2[13] ));
 sg13g2_dfrbp_1 _5683_ (.CLK(net923),
    .RESET_B(net1010),
    .D(_0117_),
    .Q_N(_2899_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator2[14] ));
 sg13g2_dfrbp_1 _5684_ (.CLK(net924),
    .RESET_B(net1011),
    .D(_0118_),
    .Q_N(_2900_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator2[15] ));
 sg13g2_dfrbp_1 _5685_ (.CLK(net924),
    .RESET_B(net1010),
    .D(_0119_),
    .Q_N(_2901_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator2[16] ));
 sg13g2_dfrbp_1 _5686_ (.CLK(net927),
    .RESET_B(net1014),
    .D(_0120_),
    .Q_N(_2902_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator2[17] ));
 sg13g2_dfrbp_1 _5687_ (.CLK(net923),
    .RESET_B(net1010),
    .D(_0121_),
    .Q_N(\u_ddc_top_level.dsm_right_inst.out_bitstream ),
    .Q(\u_ddc_top_level.dsm_right_inst.feedback[17] ));
 sg13g2_dfrbp_1 _5688_ (.CLK(net911),
    .RESET_B(net998),
    .D(_0150_),
    .Q_N(_2903_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator1[0] ));
 sg13g2_dfrbp_1 _5689_ (.CLK(net911),
    .RESET_B(net998),
    .D(_0160_),
    .Q_N(_2904_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator1[1] ));
 sg13g2_dfrbp_1 _5690_ (.CLK(net911),
    .RESET_B(net998),
    .D(_0161_),
    .Q_N(_2905_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator1[2] ));
 sg13g2_dfrbp_1 _5691_ (.CLK(net913),
    .RESET_B(net999),
    .D(_0162_),
    .Q_N(_2906_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator1[3] ));
 sg13g2_dfrbp_1 _5692_ (.CLK(net911),
    .RESET_B(net998),
    .D(_0163_),
    .Q_N(_2907_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator1[4] ));
 sg13g2_dfrbp_1 _5693_ (.CLK(net911),
    .RESET_B(net1002),
    .D(_0164_),
    .Q_N(_2908_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator1[5] ));
 sg13g2_dfrbp_1 _5694_ (.CLK(net916),
    .RESET_B(net1002),
    .D(_0165_),
    .Q_N(_2909_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator1[6] ));
 sg13g2_dfrbp_1 _5695_ (.CLK(net916),
    .RESET_B(net1002),
    .D(_0166_),
    .Q_N(_2910_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator1[7] ));
 sg13g2_dfrbp_1 _5696_ (.CLK(net916),
    .RESET_B(net1002),
    .D(_0167_),
    .Q_N(_2911_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator1[8] ));
 sg13g2_dfrbp_1 _5697_ (.CLK(net916),
    .RESET_B(net1002),
    .D(_0168_),
    .Q_N(_2912_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator1[9] ));
 sg13g2_dfrbp_1 _5698_ (.CLK(net915),
    .RESET_B(net1001),
    .D(_0151_),
    .Q_N(_2913_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator1[10] ));
 sg13g2_dfrbp_1 _5699_ (.CLK(net915),
    .RESET_B(net1001),
    .D(_0152_),
    .Q_N(_2914_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator1[11] ));
 sg13g2_dfrbp_1 _5700_ (.CLK(net917),
    .RESET_B(net1001),
    .D(_0153_),
    .Q_N(_2915_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator1[12] ));
 sg13g2_dfrbp_1 _5701_ (.CLK(net915),
    .RESET_B(net1003),
    .D(_0154_),
    .Q_N(_2916_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator1[13] ));
 sg13g2_dfrbp_1 _5702_ (.CLK(net923),
    .RESET_B(net1010),
    .D(_0155_),
    .Q_N(_2917_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator1[14] ));
 sg13g2_dfrbp_1 _5703_ (.CLK(net923),
    .RESET_B(net1010),
    .D(_0156_),
    .Q_N(_2918_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator1[15] ));
 sg13g2_dfrbp_1 _5704_ (.CLK(net923),
    .RESET_B(net1010),
    .D(_0157_),
    .Q_N(_2919_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator1[16] ));
 sg13g2_dfrbp_1 _5705_ (.CLK(net923),
    .RESET_B(net1010),
    .D(_0158_),
    .Q_N(_2920_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator1[17] ));
 sg13g2_dfrbp_1 _5706_ (.CLK(net923),
    .RESET_B(net1010),
    .D(_0159_),
    .Q_N(_2921_),
    .Q(\u_ddc_top_level.dsm_right_inst.integrator1[18] ));
 sg13g2_dfrbp_1 _5707_ (.CLK(net970),
    .RESET_B(net1057),
    .D(_0169_),
    .Q_N(_2922_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator2[0] ));
 sg13g2_dfrbp_1 _5708_ (.CLK(net971),
    .RESET_B(net1058),
    .D(_0179_),
    .Q_N(_2923_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator2[1] ));
 sg13g2_dfrbp_1 _5709_ (.CLK(net970),
    .RESET_B(net1057),
    .D(_0180_),
    .Q_N(_2924_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator2[2] ));
 sg13g2_dfrbp_1 _5710_ (.CLK(net971),
    .RESET_B(net1058),
    .D(_0181_),
    .Q_N(_2925_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator2[3] ));
 sg13g2_dfrbp_1 _5711_ (.CLK(net971),
    .RESET_B(net1059),
    .D(_0182_),
    .Q_N(_2926_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator2[4] ));
 sg13g2_dfrbp_1 _5712_ (.CLK(net971),
    .RESET_B(net1058),
    .D(_0183_),
    .Q_N(_2927_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator2[5] ));
 sg13g2_dfrbp_1 _5713_ (.CLK(net971),
    .RESET_B(net1058),
    .D(_0184_),
    .Q_N(_2928_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator2[6] ));
 sg13g2_dfrbp_1 _5714_ (.CLK(net968),
    .RESET_B(net1056),
    .D(_0185_),
    .Q_N(_2929_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator2[7] ));
 sg13g2_dfrbp_1 _5715_ (.CLK(net969),
    .RESET_B(net1056),
    .D(_0186_),
    .Q_N(_2930_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator2[8] ));
 sg13g2_dfrbp_1 _5716_ (.CLK(net969),
    .RESET_B(net1056),
    .D(_0187_),
    .Q_N(_2931_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator2[9] ));
 sg13g2_dfrbp_1 _5717_ (.CLK(net959),
    .RESET_B(net1047),
    .D(_0170_),
    .Q_N(_2932_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator2[10] ));
 sg13g2_dfrbp_1 _5718_ (.CLK(net960),
    .RESET_B(net1048),
    .D(_0171_),
    .Q_N(_2933_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator2[11] ));
 sg13g2_dfrbp_1 _5719_ (.CLK(net960),
    .RESET_B(net1048),
    .D(_0172_),
    .Q_N(_2934_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator2[12] ));
 sg13g2_dfrbp_1 _5720_ (.CLK(net960),
    .RESET_B(net1048),
    .D(_0173_),
    .Q_N(_2935_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator2[13] ));
 sg13g2_dfrbp_1 _5721_ (.CLK(net958),
    .RESET_B(net1046),
    .D(_0174_),
    .Q_N(_2936_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator2[14] ));
 sg13g2_dfrbp_1 _5722_ (.CLK(net958),
    .RESET_B(net1046),
    .D(_0175_),
    .Q_N(_2937_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator2[15] ));
 sg13g2_dfrbp_1 _5723_ (.CLK(net958),
    .RESET_B(net1046),
    .D(_0176_),
    .Q_N(_2938_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator2[16] ));
 sg13g2_dfrbp_1 _5724_ (.CLK(net958),
    .RESET_B(net1046),
    .D(_0177_),
    .Q_N(_2939_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator2[17] ));
 sg13g2_dfrbp_1 _5725_ (.CLK(net927),
    .RESET_B(net1014),
    .D(_0178_),
    .Q_N(\u_ddc_top_level.dsm_left_inst.out_bitstream ),
    .Q(\u_ddc_top_level.dsm_left_inst.feedback[17] ));
 sg13g2_dfrbp_1 _5726_ (.CLK(net966),
    .RESET_B(net1057),
    .D(_0131_),
    .Q_N(_2940_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator1[0] ));
 sg13g2_dfrbp_1 _5727_ (.CLK(net970),
    .RESET_B(net1057),
    .D(_0141_),
    .Q_N(_2941_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator1[1] ));
 sg13g2_dfrbp_1 _5728_ (.CLK(net970),
    .RESET_B(net1057),
    .D(_0142_),
    .Q_N(_2942_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator1[2] ));
 sg13g2_dfrbp_1 _5729_ (.CLK(net970),
    .RESET_B(net1057),
    .D(_0143_),
    .Q_N(_2943_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator1[3] ));
 sg13g2_dfrbp_1 _5730_ (.CLK(net970),
    .RESET_B(net1058),
    .D(_0144_),
    .Q_N(_2944_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator1[4] ));
 sg13g2_dfrbp_1 _5731_ (.CLK(net971),
    .RESET_B(net1058),
    .D(_0145_),
    .Q_N(_2945_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator1[5] ));
 sg13g2_dfrbp_1 _5732_ (.CLK(net971),
    .RESET_B(net1058),
    .D(_0146_),
    .Q_N(_2946_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator1[6] ));
 sg13g2_dfrbp_1 _5733_ (.CLK(net969),
    .RESET_B(net1055),
    .D(_0147_),
    .Q_N(_2947_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator1[7] ));
 sg13g2_dfrbp_1 _5734_ (.CLK(net969),
    .RESET_B(net1056),
    .D(_0148_),
    .Q_N(_2948_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator1[8] ));
 sg13g2_dfrbp_1 _5735_ (.CLK(net968),
    .RESET_B(net1056),
    .D(_0149_),
    .Q_N(_2949_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator1[9] ));
 sg13g2_dfrbp_1 _5736_ (.CLK(net960),
    .RESET_B(net1048),
    .D(_0132_),
    .Q_N(_2950_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator1[10] ));
 sg13g2_dfrbp_1 _5737_ (.CLK(net960),
    .RESET_B(net1048),
    .D(_0133_),
    .Q_N(_2951_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator1[11] ));
 sg13g2_dfrbp_1 _5738_ (.CLK(net960),
    .RESET_B(net1048),
    .D(_0134_),
    .Q_N(_2952_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator1[12] ));
 sg13g2_dfrbp_1 _5739_ (.CLK(net960),
    .RESET_B(net1048),
    .D(_0135_),
    .Q_N(_2953_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator1[13] ));
 sg13g2_dfrbp_1 _5740_ (.CLK(net957),
    .RESET_B(net1045),
    .D(_0136_),
    .Q_N(_2954_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator1[14] ));
 sg13g2_dfrbp_1 _5741_ (.CLK(net958),
    .RESET_B(net1046),
    .D(_0137_),
    .Q_N(_2955_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator1[15] ));
 sg13g2_dfrbp_1 _5742_ (.CLK(net958),
    .RESET_B(net1046),
    .D(_0138_),
    .Q_N(_2956_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator1[16] ));
 sg13g2_dfrbp_1 _5743_ (.CLK(net958),
    .RESET_B(net1046),
    .D(_0139_),
    .Q_N(_2957_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator1[17] ));
 sg13g2_dfrbp_1 _5744_ (.CLK(net958),
    .RESET_B(net1046),
    .D(_0140_),
    .Q_N(_2853_),
    .Q(\u_ddc_top_level.dsm_left_inst.integrator1[18] ));
 sg13g2_dfrbp_1 _5745_ (.CLK(_0188_),
    .RESET_B(net974),
    .D(_0431_),
    .Q_N(_2852_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out1[0] ));
 sg13g2_dfrbp_1 _5746_ (.CLK(_0189_),
    .RESET_B(net976),
    .D(_0432_),
    .Q_N(_2851_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out1[1] ));
 sg13g2_dfrbp_1 _5747_ (.CLK(_0190_),
    .RESET_B(net976),
    .D(_0433_),
    .Q_N(_2850_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out1[2] ));
 sg13g2_dfrbp_1 _5748_ (.CLK(_0191_),
    .RESET_B(net977),
    .D(_0434_),
    .Q_N(_2849_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out1[3] ));
 sg13g2_dfrbp_1 _5749_ (.CLK(_0192_),
    .RESET_B(net986),
    .D(_0435_),
    .Q_N(_2848_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out1[4] ));
 sg13g2_dfrbp_1 _5750_ (.CLK(_0193_),
    .RESET_B(net986),
    .D(_0436_),
    .Q_N(_2847_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out1[5] ));
 sg13g2_dfrbp_1 _5751_ (.CLK(_0194_),
    .RESET_B(net989),
    .D(_0437_),
    .Q_N(_2846_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out1[6] ));
 sg13g2_dfrbp_1 _5752_ (.CLK(_0195_),
    .RESET_B(net989),
    .D(_0438_),
    .Q_N(_2845_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out1[7] ));
 sg13g2_dfrbp_1 _5753_ (.CLK(_0196_),
    .RESET_B(net990),
    .D(_0439_),
    .Q_N(_2844_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out1[8] ));
 sg13g2_dfrbp_1 _5754_ (.CLK(_0197_),
    .RESET_B(net990),
    .D(_0440_),
    .Q_N(_2843_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out1[9] ));
 sg13g2_dfrbp_1 _5755_ (.CLK(_0198_),
    .RESET_B(net991),
    .D(_0441_),
    .Q_N(_2842_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out1[10] ));
 sg13g2_dfrbp_1 _5756_ (.CLK(_0199_),
    .RESET_B(net991),
    .D(_0442_),
    .Q_N(_2841_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out1[11] ));
 sg13g2_dfrbp_1 _5757_ (.CLK(_0200_),
    .RESET_B(net991),
    .D(_0443_),
    .Q_N(_2840_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out1[12] ));
 sg13g2_dfrbp_1 _5758_ (.CLK(_0201_),
    .RESET_B(net1005),
    .D(_0444_),
    .Q_N(_2839_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out1[13] ));
 sg13g2_dfrbp_1 _5759_ (.CLK(_0202_),
    .RESET_B(net1005),
    .D(_0445_),
    .Q_N(_2838_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out1[14] ));
 sg13g2_dfrbp_1 _5760_ (.CLK(_0203_),
    .RESET_B(net1005),
    .D(_0446_),
    .Q_N(_2837_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out1[15] ));
 sg13g2_dfrbp_1 _5761_ (.CLK(_0204_),
    .RESET_B(net1006),
    .D(_0447_),
    .Q_N(_2836_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out1[16] ));
 sg13g2_dfrbp_1 _5762_ (.CLK(_0205_),
    .RESET_B(net1006),
    .D(_0448_),
    .Q_N(_2835_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out1[17] ));
 sg13g2_dfrbp_1 _5763_ (.CLK(_0206_),
    .RESET_B(net974),
    .D(_0449_),
    .Q_N(_2834_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out2[0] ));
 sg13g2_dfrbp_1 _5764_ (.CLK(_0207_),
    .RESET_B(net974),
    .D(_0450_),
    .Q_N(_2833_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out2[1] ));
 sg13g2_dfrbp_1 _5765_ (.CLK(_0208_),
    .RESET_B(net977),
    .D(_0451_),
    .Q_N(_2832_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out2[2] ));
 sg13g2_dfrbp_1 _5766_ (.CLK(_0209_),
    .RESET_B(net977),
    .D(_0452_),
    .Q_N(_2831_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out2[3] ));
 sg13g2_dfrbp_1 _5767_ (.CLK(_0210_),
    .RESET_B(net978),
    .D(_0453_),
    .Q_N(_2830_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out2[4] ));
 sg13g2_dfrbp_1 _5768_ (.CLK(_0211_),
    .RESET_B(net978),
    .D(_0454_),
    .Q_N(_2829_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out2[5] ));
 sg13g2_dfrbp_1 _5769_ (.CLK(_0212_),
    .RESET_B(net982),
    .D(_0455_),
    .Q_N(_2828_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out2[6] ));
 sg13g2_dfrbp_1 _5770_ (.CLK(_0213_),
    .RESET_B(net982),
    .D(_0456_),
    .Q_N(_2827_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out2[7] ));
 sg13g2_dfrbp_1 _5771_ (.CLK(_0214_),
    .RESET_B(net982),
    .D(_0457_),
    .Q_N(_2826_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out2[8] ));
 sg13g2_dfrbp_1 _5772_ (.CLK(_0215_),
    .RESET_B(net983),
    .D(_0458_),
    .Q_N(_2825_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out2[9] ));
 sg13g2_dfrbp_1 _5773_ (.CLK(_0216_),
    .RESET_B(net983),
    .D(_0459_),
    .Q_N(_2824_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out2[10] ));
 sg13g2_dfrbp_1 _5774_ (.CLK(_0217_),
    .RESET_B(net982),
    .D(_0460_),
    .Q_N(_2823_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out2[11] ));
 sg13g2_dfrbp_1 _5775_ (.CLK(_0218_),
    .RESET_B(net982),
    .D(_0461_),
    .Q_N(_2822_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out2[12] ));
 sg13g2_dfrbp_1 _5776_ (.CLK(_0219_),
    .RESET_B(net999),
    .D(_0462_),
    .Q_N(_2821_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out2[13] ));
 sg13g2_dfrbp_1 _5777_ (.CLK(_0220_),
    .RESET_B(net997),
    .D(_0463_),
    .Q_N(_2820_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out2[14] ));
 sg13g2_dfrbp_1 _5778_ (.CLK(_0221_),
    .RESET_B(net997),
    .D(_0464_),
    .Q_N(_2819_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out2[15] ));
 sg13g2_dfrbp_1 _5779_ (.CLK(_0222_),
    .RESET_B(net997),
    .D(_0465_),
    .Q_N(_2818_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out2[16] ));
 sg13g2_dfrbp_1 _5780_ (.CLK(_0223_),
    .RESET_B(net997),
    .D(_0466_),
    .Q_N(_2817_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out2[17] ));
 sg13g2_dfrbp_1 _5781_ (.CLK(_0224_),
    .RESET_B(net995),
    .D(_0467_),
    .Q_N(_2816_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out2[18] ));
 sg13g2_dfrbp_1 _5782_ (.CLK(_0225_),
    .RESET_B(net985),
    .D(_0468_),
    .Q_N(_2815_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg0[0] ));
 sg13g2_dfrbp_1 _5783_ (.CLK(_0226_),
    .RESET_B(net985),
    .D(_0469_),
    .Q_N(_2814_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg0[1] ));
 sg13g2_dfrbp_1 _5784_ (.CLK(_0227_),
    .RESET_B(net985),
    .D(_0470_),
    .Q_N(_2813_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg0[2] ));
 sg13g2_dfrbp_1 _5785_ (.CLK(_0228_),
    .RESET_B(net987),
    .D(_0471_),
    .Q_N(_2812_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg0[3] ));
 sg13g2_dfrbp_1 _5786_ (.CLK(_0229_),
    .RESET_B(net987),
    .D(_0472_),
    .Q_N(_2811_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg0[4] ));
 sg13g2_dfrbp_1 _5787_ (.CLK(_0230_),
    .RESET_B(net988),
    .D(_0473_),
    .Q_N(_2810_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg0[5] ));
 sg13g2_dfrbp_1 _5788_ (.CLK(_0231_),
    .RESET_B(net988),
    .D(_0474_),
    .Q_N(_2809_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg0[6] ));
 sg13g2_dfrbp_1 _5789_ (.CLK(_0232_),
    .RESET_B(net988),
    .D(_0475_),
    .Q_N(_2808_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg0[7] ));
 sg13g2_dfrbp_1 _5790_ (.CLK(_0233_),
    .RESET_B(net992),
    .D(_0476_),
    .Q_N(_2807_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg0[8] ));
 sg13g2_dfrbp_1 _5791_ (.CLK(_0234_),
    .RESET_B(net992),
    .D(_0477_),
    .Q_N(_2806_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg0[9] ));
 sg13g2_dfrbp_1 _5792_ (.CLK(_0235_),
    .RESET_B(net992),
    .D(_0478_),
    .Q_N(_2805_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg0[10] ));
 sg13g2_dfrbp_1 _5793_ (.CLK(_0236_),
    .RESET_B(net993),
    .D(_0479_),
    .Q_N(_2804_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg0[11] ));
 sg13g2_dfrbp_1 _5794_ (.CLK(_0237_),
    .RESET_B(net993),
    .D(_0480_),
    .Q_N(_2803_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg0[12] ));
 sg13g2_dfrbp_1 _5795_ (.CLK(_0238_),
    .RESET_B(net1009),
    .D(_0481_),
    .Q_N(_2802_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg0[13] ));
 sg13g2_dfrbp_1 _5796_ (.CLK(_0239_),
    .RESET_B(net1008),
    .D(_0482_),
    .Q_N(_2801_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg0[14] ));
 sg13g2_dfrbp_1 _5797_ (.CLK(_0240_),
    .RESET_B(net1008),
    .D(_0483_),
    .Q_N(_2958_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg0[15] ));
 sg13g2_dfrbp_1 _5798_ (.CLK(net887),
    .RESET_B(net974),
    .D(_0059_),
    .Q_N(_2959_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[0] ));
 sg13g2_dfrbp_1 _5799_ (.CLK(net887),
    .RESET_B(net974),
    .D(_0070_),
    .Q_N(_2960_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[1] ));
 sg13g2_dfrbp_1 _5800_ (.CLK(net888),
    .RESET_B(net975),
    .D(_0075_),
    .Q_N(_2961_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[2] ));
 sg13g2_dfrbp_1 _5801_ (.CLK(net888),
    .RESET_B(net975),
    .D(_0076_),
    .Q_N(_2962_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[3] ));
 sg13g2_dfrbp_1 _5802_ (.CLK(net888),
    .RESET_B(net979),
    .D(_0077_),
    .Q_N(_2963_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[4] ));
 sg13g2_dfrbp_1 _5803_ (.CLK(net894),
    .RESET_B(net981),
    .D(_0078_),
    .Q_N(_2964_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[5] ));
 sg13g2_dfrbp_1 _5804_ (.CLK(net894),
    .RESET_B(net979),
    .D(_0079_),
    .Q_N(_2965_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[6] ));
 sg13g2_dfrbp_1 _5805_ (.CLK(net894),
    .RESET_B(net979),
    .D(_0080_),
    .Q_N(_2966_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[7] ));
 sg13g2_dfrbp_1 _5806_ (.CLK(net893),
    .RESET_B(net980),
    .D(_0081_),
    .Q_N(_2967_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[8] ));
 sg13g2_dfrbp_1 _5807_ (.CLK(net897),
    .RESET_B(net980),
    .D(_0082_),
    .Q_N(_2968_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[9] ));
 sg13g2_dfrbp_1 _5808_ (.CLK(net893),
    .RESET_B(net980),
    .D(_0060_),
    .Q_N(_2969_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[10] ));
 sg13g2_dfrbp_1 _5809_ (.CLK(net893),
    .RESET_B(net980),
    .D(_0061_),
    .Q_N(_2970_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[11] ));
 sg13g2_dfrbp_1 _5810_ (.CLK(net909),
    .RESET_B(net995),
    .D(_0062_),
    .Q_N(_2971_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[12] ));
 sg13g2_dfrbp_1 _5811_ (.CLK(net909),
    .RESET_B(net995),
    .D(_0063_),
    .Q_N(_2972_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[13] ));
 sg13g2_dfrbp_1 _5812_ (.CLK(net912),
    .RESET_B(net997),
    .D(_0064_),
    .Q_N(_2973_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[14] ));
 sg13g2_dfrbp_1 _5813_ (.CLK(net909),
    .RESET_B(net995),
    .D(_0065_),
    .Q_N(_2974_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[15] ));
 sg13g2_dfrbp_1 _5814_ (.CLK(net910),
    .RESET_B(net996),
    .D(_0066_),
    .Q_N(_2975_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[16] ));
 sg13g2_dfrbp_1 _5815_ (.CLK(net910),
    .RESET_B(net996),
    .D(_0067_),
    .Q_N(_2976_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[17] ));
 sg13g2_dfrbp_1 _5816_ (.CLK(net910),
    .RESET_B(net996),
    .D(_0068_),
    .Q_N(_2977_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[18] ));
 sg13g2_dfrbp_1 _5817_ (.CLK(net910),
    .RESET_B(net996),
    .D(_0069_),
    .Q_N(_2978_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[19] ));
 sg13g2_dfrbp_1 _5818_ (.CLK(net914),
    .RESET_B(net1000),
    .D(_0071_),
    .Q_N(_2979_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[20] ));
 sg13g2_dfrbp_1 _5819_ (.CLK(net914),
    .RESET_B(net1000),
    .D(_0072_),
    .Q_N(_2980_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[21] ));
 sg13g2_dfrbp_1 _5820_ (.CLK(net917),
    .RESET_B(net1003),
    .D(_0073_),
    .Q_N(_2981_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[22] ));
 sg13g2_dfrbp_1 _5821_ (.CLK(net917),
    .RESET_B(net1003),
    .D(_0074_),
    .Q_N(_2800_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg1[23] ));
 sg13g2_dfrbp_1 _5822_ (.CLK(_0241_),
    .RESET_B(net1020),
    .D(_0484_),
    .Q_N(_2799_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out0[0] ));
 sg13g2_dfrbp_1 _5823_ (.CLK(_0242_),
    .RESET_B(net1020),
    .D(_0485_),
    .Q_N(_2798_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out0[1] ));
 sg13g2_dfrbp_1 _5824_ (.CLK(_0243_),
    .RESET_B(net1020),
    .D(_0486_),
    .Q_N(_2797_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out0[2] ));
 sg13g2_dfrbp_1 _5825_ (.CLK(_0244_),
    .RESET_B(net1020),
    .D(_0487_),
    .Q_N(_2796_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out0[3] ));
 sg13g2_dfrbp_1 _5826_ (.CLK(_0245_),
    .RESET_B(net1021),
    .D(_0488_),
    .Q_N(_2795_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out0[4] ));
 sg13g2_dfrbp_1 _5827_ (.CLK(_0246_),
    .RESET_B(net1021),
    .D(_0489_),
    .Q_N(_2794_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out0[5] ));
 sg13g2_dfrbp_1 _5828_ (.CLK(_0247_),
    .RESET_B(net1021),
    .D(_0490_),
    .Q_N(_2793_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out0[6] ));
 sg13g2_dfrbp_1 _5829_ (.CLK(_0248_),
    .RESET_B(net1026),
    .D(_0491_),
    .Q_N(_2792_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out0[7] ));
 sg13g2_dfrbp_1 _5830_ (.CLK(_0249_),
    .RESET_B(net1026),
    .D(_0492_),
    .Q_N(_2791_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out0[8] ));
 sg13g2_dfrbp_1 _5831_ (.CLK(_0250_),
    .RESET_B(net1026),
    .D(_0493_),
    .Q_N(_2790_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out0[9] ));
 sg13g2_dfrbp_1 _5832_ (.CLK(_0251_),
    .RESET_B(net1025),
    .D(_0494_),
    .Q_N(_2789_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out0[10] ));
 sg13g2_dfrbp_1 _5833_ (.CLK(_0252_),
    .RESET_B(net1024),
    .D(_0495_),
    .Q_N(_2788_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out0[11] ));
 sg13g2_dfrbp_1 _5834_ (.CLK(_0253_),
    .RESET_B(net1042),
    .D(_0496_),
    .Q_N(_2787_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out0[12] ));
 sg13g2_dfrbp_1 _5835_ (.CLK(_0254_),
    .RESET_B(net1040),
    .D(_0497_),
    .Q_N(_2786_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out0[13] ));
 sg13g2_dfrbp_1 _5836_ (.CLK(_0255_),
    .RESET_B(net1042),
    .D(_0498_),
    .Q_N(_2785_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out0[14] ));
 sg13g2_dfrbp_1 _5837_ (.CLK(_0256_),
    .RESET_B(net1041),
    .D(_0499_),
    .Q_N(_2784_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out0[15] ));
 sg13g2_dfrbp_1 _5838_ (.CLK(_0257_),
    .RESET_B(net1041),
    .D(_0500_),
    .Q_N(_2982_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out0[16] ));
 sg13g2_dfrbp_1 _5839_ (.CLK(net887),
    .RESET_B(net974),
    .D(_0083_),
    .Q_N(_2983_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg2[0] ));
 sg13g2_dfrbp_1 _5840_ (.CLK(net888),
    .RESET_B(net975),
    .D(_0094_),
    .Q_N(_2984_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg2[1] ));
 sg13g2_dfrbp_1 _5841_ (.CLK(net888),
    .RESET_B(net975),
    .D(_0103_),
    .Q_N(_2985_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg2[2] ));
 sg13g2_dfrbp_1 _5842_ (.CLK(net888),
    .RESET_B(net975),
    .D(_0104_),
    .Q_N(_2986_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg2[3] ));
 sg13g2_dfrbp_1 _5843_ (.CLK(net888),
    .RESET_B(net979),
    .D(_0105_),
    .Q_N(_2987_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg2[4] ));
 sg13g2_dfrbp_1 _5844_ (.CLK(net894),
    .RESET_B(net979),
    .D(_0106_),
    .Q_N(_2988_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg2[5] ));
 sg13g2_dfrbp_1 _5845_ (.CLK(net894),
    .RESET_B(net979),
    .D(_0107_),
    .Q_N(_2989_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg2[6] ));
 sg13g2_dfrbp_1 _5846_ (.CLK(net894),
    .RESET_B(net979),
    .D(_0108_),
    .Q_N(_2990_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg2[7] ));
 sg13g2_dfrbp_1 _5847_ (.CLK(net893),
    .RESET_B(net980),
    .D(_0109_),
    .Q_N(_2991_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg2[8] ));
 sg13g2_dfrbp_1 _5848_ (.CLK(net893),
    .RESET_B(net980),
    .D(_0110_),
    .Q_N(_2992_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg2[9] ));
 sg13g2_dfrbp_1 _5849_ (.CLK(net893),
    .RESET_B(net980),
    .D(_0084_),
    .Q_N(_2993_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg2[10] ));
 sg13g2_dfrbp_1 _5850_ (.CLK(net893),
    .RESET_B(net980),
    .D(_0085_),
    .Q_N(_2994_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg2[11] ));
 sg13g2_dfrbp_1 _5851_ (.CLK(net909),
    .RESET_B(net996),
    .D(_0086_),
    .Q_N(_2995_),
    .Q(\u_ddc_top_level.cic_out_right[0] ));
 sg13g2_dfrbp_1 _5852_ (.CLK(net911),
    .RESET_B(net998),
    .D(_0087_),
    .Q_N(_2996_),
    .Q(\u_ddc_top_level.cic_out_right[1] ));
 sg13g2_dfrbp_1 _5853_ (.CLK(net911),
    .RESET_B(net998),
    .D(_0088_),
    .Q_N(_2997_),
    .Q(\u_ddc_top_level.cic_out_right[2] ));
 sg13g2_dfrbp_1 _5854_ (.CLK(net911),
    .RESET_B(net998),
    .D(_0089_),
    .Q_N(_2998_),
    .Q(\u_ddc_top_level.cic_out_right[3] ));
 sg13g2_dfrbp_1 _5855_ (.CLK(net910),
    .RESET_B(net996),
    .D(_0090_),
    .Q_N(_2999_),
    .Q(\u_ddc_top_level.cic_out_right[4] ));
 sg13g2_dfrbp_1 _5856_ (.CLK(net910),
    .RESET_B(net996),
    .D(_0091_),
    .Q_N(_3000_),
    .Q(\u_ddc_top_level.cic_out_right[5] ));
 sg13g2_dfrbp_1 _5857_ (.CLK(net914),
    .RESET_B(net1000),
    .D(_0092_),
    .Q_N(_3001_),
    .Q(\u_ddc_top_level.cic_out_right[6] ));
 sg13g2_dfrbp_1 _5858_ (.CLK(net914),
    .RESET_B(net1000),
    .D(_0093_),
    .Q_N(_3002_),
    .Q(\u_ddc_top_level.cic_out_right[7] ));
 sg13g2_dfrbp_1 _5859_ (.CLK(net914),
    .RESET_B(net1000),
    .D(_0095_),
    .Q_N(_3003_),
    .Q(\u_ddc_top_level.cic_out_right[8] ));
 sg13g2_dfrbp_1 _5860_ (.CLK(net914),
    .RESET_B(net1000),
    .D(_0096_),
    .Q_N(_3004_),
    .Q(\u_ddc_top_level.cic_out_right[9] ));
 sg13g2_dfrbp_1 _5861_ (.CLK(net917),
    .RESET_B(net1000),
    .D(_0097_),
    .Q_N(_3005_),
    .Q(\u_ddc_top_level.cic_out_right[10] ));
 sg13g2_dfrbp_1 _5862_ (.CLK(net914),
    .RESET_B(net1003),
    .D(_0098_),
    .Q_N(_3006_),
    .Q(\u_ddc_top_level.cic_out_right[11] ));
 sg13g2_dfrbp_1 _5863_ (.CLK(net914),
    .RESET_B(net1000),
    .D(_0099_),
    .Q_N(_3007_),
    .Q(\u_ddc_top_level.cic_out_right[12] ));
 sg13g2_dfrbp_1 _5864_ (.CLK(net915),
    .RESET_B(net1001),
    .D(_0100_),
    .Q_N(_3008_),
    .Q(\u_ddc_top_level.cic_out_right[13] ));
 sg13g2_dfrbp_1 _5865_ (.CLK(net915),
    .RESET_B(net1001),
    .D(_0101_),
    .Q_N(_3009_),
    .Q(\u_ddc_top_level.cic_out_right[14] ));
 sg13g2_dfrbp_1 _5866_ (.CLK(net915),
    .RESET_B(net1001),
    .D(_0102_),
    .Q_N(_2783_),
    .Q(\u_ddc_top_level.cic_out_right[15] ));
 sg13g2_dfrbp_1 _5867_ (.CLK(_0258_),
    .RESET_B(net976),
    .D(_0501_),
    .Q_N(_2782_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg1[0] ));
 sg13g2_dfrbp_1 _5868_ (.CLK(_0259_),
    .RESET_B(net976),
    .D(_0502_),
    .Q_N(_2781_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg1[1] ));
 sg13g2_dfrbp_1 _5869_ (.CLK(_0260_),
    .RESET_B(net976),
    .D(_0503_),
    .Q_N(_2780_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg1[2] ));
 sg13g2_dfrbp_1 _5870_ (.CLK(_0261_),
    .RESET_B(net985),
    .D(_0504_),
    .Q_N(_2779_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg1[3] ));
 sg13g2_dfrbp_1 _5871_ (.CLK(_0262_),
    .RESET_B(net986),
    .D(_0505_),
    .Q_N(_2778_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg1[4] ));
 sg13g2_dfrbp_1 _5872_ (.CLK(_0263_),
    .RESET_B(net985),
    .D(_0506_),
    .Q_N(_2777_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg1[5] ));
 sg13g2_dfrbp_1 _5873_ (.CLK(_0264_),
    .RESET_B(net986),
    .D(_0507_),
    .Q_N(_2776_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg1[6] ));
 sg13g2_dfrbp_1 _5874_ (.CLK(_0265_),
    .RESET_B(net986),
    .D(_0508_),
    .Q_N(_2775_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg1[7] ));
 sg13g2_dfrbp_1 _5875_ (.CLK(_0266_),
    .RESET_B(net990),
    .D(_0509_),
    .Q_N(_2774_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg1[8] ));
 sg13g2_dfrbp_1 _5876_ (.CLK(_0267_),
    .RESET_B(net990),
    .D(_0510_),
    .Q_N(_2773_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg1[9] ));
 sg13g2_dfrbp_1 _5877_ (.CLK(_0268_),
    .RESET_B(net990),
    .D(_0511_),
    .Q_N(_2772_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg1[10] ));
 sg13g2_dfrbp_1 _5878_ (.CLK(_0269_),
    .RESET_B(net993),
    .D(_0512_),
    .Q_N(_2771_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg1[11] ));
 sg13g2_dfrbp_1 _5879_ (.CLK(_0270_),
    .RESET_B(net993),
    .D(_0513_),
    .Q_N(_2770_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg1[12] ));
 sg13g2_dfrbp_1 _5880_ (.CLK(_0271_),
    .RESET_B(net1007),
    .D(_0514_),
    .Q_N(_2769_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg1[13] ));
 sg13g2_dfrbp_1 _5881_ (.CLK(_0272_),
    .RESET_B(net1007),
    .D(_0515_),
    .Q_N(_2768_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg1[14] ));
 sg13g2_dfrbp_1 _5882_ (.CLK(_0273_),
    .RESET_B(net1008),
    .D(_0516_),
    .Q_N(_2767_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg1[15] ));
 sg13g2_dfrbp_1 _5883_ (.CLK(_0274_),
    .RESET_B(net1006),
    .D(_0517_),
    .Q_N(_2766_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg1[16] ));
 sg13g2_dfrbp_1 _5884_ (.CLK(net887),
    .RESET_B(net974),
    .D(_0518_),
    .Q_N(_2765_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg0[0] ));
 sg13g2_dfrbp_1 _5885_ (.CLK(net889),
    .RESET_B(net975),
    .D(_0519_),
    .Q_N(_2764_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg0[1] ));
 sg13g2_dfrbp_1 _5886_ (.CLK(net889),
    .RESET_B(net975),
    .D(_0520_),
    .Q_N(_2763_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg0[2] ));
 sg13g2_dfrbp_1 _5887_ (.CLK(net889),
    .RESET_B(net978),
    .D(_0521_),
    .Q_N(_2762_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg0[3] ));
 sg13g2_dfrbp_1 _5888_ (.CLK(net889),
    .RESET_B(net978),
    .D(_0522_),
    .Q_N(_2761_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg0[4] ));
 sg13g2_dfrbp_1 _5889_ (.CLK(net895),
    .RESET_B(net982),
    .D(_0523_),
    .Q_N(_2760_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg0[5] ));
 sg13g2_dfrbp_1 _5890_ (.CLK(net894),
    .RESET_B(net979),
    .D(_0524_),
    .Q_N(_2759_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg0[6] ));
 sg13g2_dfrbp_1 _5891_ (.CLK(net895),
    .RESET_B(net982),
    .D(_0525_),
    .Q_N(_2758_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg0[7] ));
 sg13g2_dfrbp_1 _5892_ (.CLK(net896),
    .RESET_B(net983),
    .D(_0526_),
    .Q_N(_2757_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg0[8] ));
 sg13g2_dfrbp_1 _5893_ (.CLK(net897),
    .RESET_B(net981),
    .D(_0527_),
    .Q_N(_2756_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg0[9] ));
 sg13g2_dfrbp_1 _5894_ (.CLK(net896),
    .RESET_B(net983),
    .D(_0528_),
    .Q_N(_2755_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg0[10] ));
 sg13g2_dfrbp_1 _5895_ (.CLK(net896),
    .RESET_B(net982),
    .D(_0529_),
    .Q_N(_2754_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg0[11] ));
 sg13g2_dfrbp_1 _5896_ (.CLK(net893),
    .RESET_B(net995),
    .D(_0530_),
    .Q_N(_2753_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg0[12] ));
 sg13g2_dfrbp_1 _5897_ (.CLK(net912),
    .RESET_B(net997),
    .D(_0531_),
    .Q_N(_2752_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg0[13] ));
 sg13g2_dfrbp_1 _5898_ (.CLK(net912),
    .RESET_B(net997),
    .D(_0532_),
    .Q_N(_2751_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg0[14] ));
 sg13g2_dfrbp_1 _5899_ (.CLK(net912),
    .RESET_B(net997),
    .D(_0533_),
    .Q_N(_2750_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg0[15] ));
 sg13g2_dfrbp_1 _5900_ (.CLK(net909),
    .RESET_B(net995),
    .D(_0534_),
    .Q_N(_2749_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg0[16] ));
 sg13g2_dfrbp_1 _5901_ (.CLK(net909),
    .RESET_B(net995),
    .D(_0535_),
    .Q_N(_2748_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg0[17] ));
 sg13g2_dfrbp_1 _5902_ (.CLK(net909),
    .RESET_B(net995),
    .D(_0536_),
    .Q_N(_2747_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg0[18] ));
 sg13g2_dfrbp_1 _5903_ (.CLK(net910),
    .RESET_B(net996),
    .D(_0537_),
    .Q_N(_2746_),
    .Q(\u_ddc_top_level.cic_right_inst.int_reg0[19] ));
 sg13g2_dfrbp_1 _5904_ (.CLK(_0275_),
    .RESET_B(net974),
    .D(_0538_),
    .Q_N(_2745_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg2[0] ));
 sg13g2_dfrbp_1 _5905_ (.CLK(_0276_),
    .RESET_B(net976),
    .D(_0539_),
    .Q_N(_2744_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg2[1] ));
 sg13g2_dfrbp_1 _5906_ (.CLK(_0277_),
    .RESET_B(net976),
    .D(_0540_),
    .Q_N(_2743_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg2[2] ));
 sg13g2_dfrbp_1 _5907_ (.CLK(_0278_),
    .RESET_B(net977),
    .D(_0541_),
    .Q_N(_2742_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg2[3] ));
 sg13g2_dfrbp_1 _5908_ (.CLK(_0279_),
    .RESET_B(net977),
    .D(_0542_),
    .Q_N(_2741_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg2[4] ));
 sg13g2_dfrbp_1 _5909_ (.CLK(_0280_),
    .RESET_B(net977),
    .D(_0543_),
    .Q_N(_2740_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg2[5] ));
 sg13g2_dfrbp_1 _5910_ (.CLK(_0281_),
    .RESET_B(net986),
    .D(_0544_),
    .Q_N(_2739_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg2[6] ));
 sg13g2_dfrbp_1 _5911_ (.CLK(_0282_),
    .RESET_B(net990),
    .D(_0545_),
    .Q_N(_2738_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg2[7] ));
 sg13g2_dfrbp_1 _5912_ (.CLK(_0283_),
    .RESET_B(net990),
    .D(_0546_),
    .Q_N(_2737_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg2[8] ));
 sg13g2_dfrbp_1 _5913_ (.CLK(_0284_),
    .RESET_B(net990),
    .D(_0547_),
    .Q_N(_2736_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg2[9] ));
 sg13g2_dfrbp_1 _5914_ (.CLK(_0285_),
    .RESET_B(net991),
    .D(_0548_),
    .Q_N(_2735_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg2[10] ));
 sg13g2_dfrbp_1 _5915_ (.CLK(_0286_),
    .RESET_B(net991),
    .D(_0549_),
    .Q_N(_2734_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg2[11] ));
 sg13g2_dfrbp_1 _5916_ (.CLK(_0287_),
    .RESET_B(net991),
    .D(_0550_),
    .Q_N(_2733_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg2[12] ));
 sg13g2_dfrbp_1 _5917_ (.CLK(_0288_),
    .RESET_B(net1005),
    .D(_0551_),
    .Q_N(_2732_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg2[13] ));
 sg13g2_dfrbp_1 _5918_ (.CLK(_0289_),
    .RESET_B(net1005),
    .D(_0552_),
    .Q_N(_2731_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg2[14] ));
 sg13g2_dfrbp_1 _5919_ (.CLK(_0290_),
    .RESET_B(net1005),
    .D(_0553_),
    .Q_N(_2730_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg2[15] ));
 sg13g2_dfrbp_1 _5920_ (.CLK(_0291_),
    .RESET_B(net1006),
    .D(_0554_),
    .Q_N(_2729_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg2[16] ));
 sg13g2_dfrbp_1 _5921_ (.CLK(_0292_),
    .RESET_B(net1006),
    .D(_0555_),
    .Q_N(_2728_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_reg2[17] ));
 sg13g2_dfrbp_1 _5922_ (.CLK(_0293_),
    .RESET_B(net1028),
    .D(_0556_),
    .Q_N(_2727_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out1[0] ));
 sg13g2_dfrbp_1 _5923_ (.CLK(_0294_),
    .RESET_B(net1028),
    .D(_0557_),
    .Q_N(_2726_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out1[1] ));
 sg13g2_dfrbp_1 _5924_ (.CLK(_0295_),
    .RESET_B(net1028),
    .D(_0558_),
    .Q_N(_2725_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out1[2] ));
 sg13g2_dfrbp_1 _5925_ (.CLK(_0296_),
    .RESET_B(net1032),
    .D(_0559_),
    .Q_N(_2724_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out1[3] ));
 sg13g2_dfrbp_1 _5926_ (.CLK(_0297_),
    .RESET_B(net1032),
    .D(_0560_),
    .Q_N(_2723_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out1[4] ));
 sg13g2_dfrbp_1 _5927_ (.CLK(_0298_),
    .RESET_B(net1021),
    .D(_0561_),
    .Q_N(_2722_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out1[5] ));
 sg13g2_dfrbp_1 _5928_ (.CLK(_0299_),
    .RESET_B(net1026),
    .D(_0562_),
    .Q_N(_2721_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out1[6] ));
 sg13g2_dfrbp_1 _5929_ (.CLK(_0300_),
    .RESET_B(net1033),
    .D(_0563_),
    .Q_N(_2720_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out1[7] ));
 sg13g2_dfrbp_1 _5930_ (.CLK(_0301_),
    .RESET_B(net1026),
    .D(_0564_),
    .Q_N(_2719_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out1[8] ));
 sg13g2_dfrbp_1 _5931_ (.CLK(_0302_),
    .RESET_B(net1027),
    .D(_0565_),
    .Q_N(_2718_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out1[9] ));
 sg13g2_dfrbp_1 _5932_ (.CLK(_0303_),
    .RESET_B(net1025),
    .D(_0566_),
    .Q_N(_2717_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out1[10] ));
 sg13g2_dfrbp_1 _5933_ (.CLK(_0304_),
    .RESET_B(net1025),
    .D(_0567_),
    .Q_N(_2716_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out1[11] ));
 sg13g2_dfrbp_1 _5934_ (.CLK(_0305_),
    .RESET_B(net1043),
    .D(_0568_),
    .Q_N(_2715_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out1[12] ));
 sg13g2_dfrbp_1 _5935_ (.CLK(_0306_),
    .RESET_B(net1043),
    .D(_0569_),
    .Q_N(_2714_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out1[13] ));
 sg13g2_dfrbp_1 _5936_ (.CLK(_0307_),
    .RESET_B(net1044),
    .D(_0570_),
    .Q_N(_2713_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out1[14] ));
 sg13g2_dfrbp_1 _5937_ (.CLK(_0308_),
    .RESET_B(net1043),
    .D(_0571_),
    .Q_N(_2712_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out1[15] ));
 sg13g2_dfrbp_1 _5938_ (.CLK(_0309_),
    .RESET_B(net1044),
    .D(_0572_),
    .Q_N(_2711_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out1[16] ));
 sg13g2_dfrbp_1 _5939_ (.CLK(_0310_),
    .RESET_B(net1044),
    .D(_0573_),
    .Q_N(_2710_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out1[17] ));
 sg13g2_dfrbp_1 _5940_ (.CLK(_0311_),
    .RESET_B(net1029),
    .D(_0574_),
    .Q_N(_2709_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out2[0] ));
 sg13g2_dfrbp_1 _5941_ (.CLK(_0312_),
    .RESET_B(net1028),
    .D(_0575_),
    .Q_N(_2708_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out2[1] ));
 sg13g2_dfrbp_1 _5942_ (.CLK(_0313_),
    .RESET_B(net1029),
    .D(_0576_),
    .Q_N(_2707_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out2[2] ));
 sg13g2_dfrbp_1 _5943_ (.CLK(_0314_),
    .RESET_B(net1029),
    .D(_0577_),
    .Q_N(_2706_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out2[3] ));
 sg13g2_dfrbp_1 _5944_ (.CLK(_0315_),
    .RESET_B(net1029),
    .D(_0578_),
    .Q_N(_2705_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out2[4] ));
 sg13g2_dfrbp_1 _5945_ (.CLK(_0316_),
    .RESET_B(net1033),
    .D(_0579_),
    .Q_N(_2704_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out2[5] ));
 sg13g2_dfrbp_1 _5946_ (.CLK(_0317_),
    .RESET_B(net1033),
    .D(_0580_),
    .Q_N(_2703_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out2[6] ));
 sg13g2_dfrbp_1 _5947_ (.CLK(_0318_),
    .RESET_B(net1033),
    .D(_0581_),
    .Q_N(_2702_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out2[7] ));
 sg13g2_dfrbp_1 _5948_ (.CLK(_0319_),
    .RESET_B(net1033),
    .D(_0582_),
    .Q_N(_2701_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out2[8] ));
 sg13g2_dfrbp_1 _5949_ (.CLK(_0320_),
    .RESET_B(net1033),
    .D(_0583_),
    .Q_N(_2700_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out2[9] ));
 sg13g2_dfrbp_1 _5950_ (.CLK(_0321_),
    .RESET_B(net1034),
    .D(_0584_),
    .Q_N(_2699_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out2[10] ));
 sg13g2_dfrbp_1 _5951_ (.CLK(_0322_),
    .RESET_B(net1034),
    .D(_0585_),
    .Q_N(_2698_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out2[11] ));
 sg13g2_dfrbp_1 _5952_ (.CLK(_0323_),
    .RESET_B(net1051),
    .D(_0586_),
    .Q_N(_2697_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out2[12] ));
 sg13g2_dfrbp_1 _5953_ (.CLK(_0324_),
    .RESET_B(net1051),
    .D(_0587_),
    .Q_N(_2696_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out2[13] ));
 sg13g2_dfrbp_1 _5954_ (.CLK(_0325_),
    .RESET_B(net1051),
    .D(_0588_),
    .Q_N(_2695_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out2[14] ));
 sg13g2_dfrbp_1 _5955_ (.CLK(_0326_),
    .RESET_B(net1051),
    .D(_0589_),
    .Q_N(_2694_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out2[15] ));
 sg13g2_dfrbp_1 _5956_ (.CLK(_0327_),
    .RESET_B(net1051),
    .D(_0590_),
    .Q_N(_2693_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out2[16] ));
 sg13g2_dfrbp_1 _5957_ (.CLK(_0328_),
    .RESET_B(net1051),
    .D(_0591_),
    .Q_N(_2692_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out2[17] ));
 sg13g2_dfrbp_1 _5958_ (.CLK(_0329_),
    .RESET_B(net1054),
    .D(_0592_),
    .Q_N(_2691_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_out2[18] ));
 sg13g2_dfrbp_1 _5959_ (.CLK(_0330_),
    .RESET_B(net1020),
    .D(_0593_),
    .Q_N(_2690_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg0[0] ));
 sg13g2_dfrbp_1 _5960_ (.CLK(_0331_),
    .RESET_B(net1020),
    .D(_0594_),
    .Q_N(_2689_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg0[1] ));
 sg13g2_dfrbp_1 _5961_ (.CLK(_0332_),
    .RESET_B(net1018),
    .D(_0595_),
    .Q_N(_2688_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg0[2] ));
 sg13g2_dfrbp_1 _5962_ (.CLK(_0333_),
    .RESET_B(net1018),
    .D(_0596_),
    .Q_N(_2687_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg0[3] ));
 sg13g2_dfrbp_1 _5963_ (.CLK(_0334_),
    .RESET_B(net1019),
    .D(_0597_),
    .Q_N(_2686_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg0[4] ));
 sg13g2_dfrbp_1 _5964_ (.CLK(_0335_),
    .RESET_B(net1019),
    .D(_0598_),
    .Q_N(_2685_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg0[5] ));
 sg13g2_dfrbp_1 _5965_ (.CLK(_0336_),
    .RESET_B(net1019),
    .D(_0599_),
    .Q_N(_2684_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg0[6] ));
 sg13g2_dfrbp_1 _5966_ (.CLK(_0337_),
    .RESET_B(net1023),
    .D(_0600_),
    .Q_N(_2683_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg0[7] ));
 sg13g2_dfrbp_1 _5967_ (.CLK(_0338_),
    .RESET_B(net1023),
    .D(_0601_),
    .Q_N(_2682_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg0[8] ));
 sg13g2_dfrbp_1 _5968_ (.CLK(_0339_),
    .RESET_B(net1023),
    .D(_0602_),
    .Q_N(_2681_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg0[9] ));
 sg13g2_dfrbp_1 _5969_ (.CLK(_0340_),
    .RESET_B(net1024),
    .D(_0603_),
    .Q_N(_2680_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg0[10] ));
 sg13g2_dfrbp_1 _5970_ (.CLK(_0341_),
    .RESET_B(net1024),
    .D(_0604_),
    .Q_N(_2679_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg0[11] ));
 sg13g2_dfrbp_1 _5971_ (.CLK(_0342_),
    .RESET_B(net1040),
    .D(_0605_),
    .Q_N(_2678_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg0[12] ));
 sg13g2_dfrbp_1 _5972_ (.CLK(_0343_),
    .RESET_B(net1040),
    .D(_0606_),
    .Q_N(_2677_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg0[13] ));
 sg13g2_dfrbp_1 _5973_ (.CLK(_0344_),
    .RESET_B(net1040),
    .D(_0607_),
    .Q_N(_2676_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg0[14] ));
 sg13g2_dfrbp_1 _5974_ (.CLK(_0345_),
    .RESET_B(net1042),
    .D(_0608_),
    .Q_N(_3010_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg0[15] ));
 sg13g2_dfrbp_1 _5975_ (.CLK(net943),
    .RESET_B(net1030),
    .D(_0007_),
    .Q_N(_3011_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[0] ));
 sg13g2_dfrbp_1 _5976_ (.CLK(net943),
    .RESET_B(net1030),
    .D(_0018_),
    .Q_N(_3012_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[1] ));
 sg13g2_dfrbp_1 _5977_ (.CLK(net943),
    .RESET_B(net1030),
    .D(_0023_),
    .Q_N(_3013_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[2] ));
 sg13g2_dfrbp_1 _5978_ (.CLK(net944),
    .RESET_B(net1031),
    .D(_0024_),
    .Q_N(_3014_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[3] ));
 sg13g2_dfrbp_1 _5979_ (.CLK(net950),
    .RESET_B(net1036),
    .D(_0025_),
    .Q_N(_3015_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[4] ));
 sg13g2_dfrbp_1 _5980_ (.CLK(net950),
    .RESET_B(net1036),
    .D(_0026_),
    .Q_N(_3016_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[5] ));
 sg13g2_dfrbp_1 _5981_ (.CLK(net948),
    .RESET_B(net1035),
    .D(_0027_),
    .Q_N(_3017_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[6] ));
 sg13g2_dfrbp_1 _5982_ (.CLK(net948),
    .RESET_B(net1035),
    .D(_0028_),
    .Q_N(_3018_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[7] ));
 sg13g2_dfrbp_1 _5983_ (.CLK(net950),
    .RESET_B(net1038),
    .D(_0029_),
    .Q_N(_3019_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[8] ));
 sg13g2_dfrbp_1 _5984_ (.CLK(net949),
    .RESET_B(net1037),
    .D(_0030_),
    .Q_N(_3020_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[9] ));
 sg13g2_dfrbp_1 _5985_ (.CLK(net949),
    .RESET_B(net1037),
    .D(_0008_),
    .Q_N(_3021_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[10] ));
 sg13g2_dfrbp_1 _5986_ (.CLK(net966),
    .RESET_B(net1053),
    .D(_0009_),
    .Q_N(_3022_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[11] ));
 sg13g2_dfrbp_1 _5987_ (.CLK(net964),
    .RESET_B(net1053),
    .D(_0010_),
    .Q_N(_3023_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[12] ));
 sg13g2_dfrbp_1 _5988_ (.CLK(net964),
    .RESET_B(net1053),
    .D(_0011_),
    .Q_N(_3024_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[13] ));
 sg13g2_dfrbp_1 _5989_ (.CLK(net964),
    .RESET_B(net1054),
    .D(_0012_),
    .Q_N(_3025_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[14] ));
 sg13g2_dfrbp_1 _5990_ (.CLK(net965),
    .RESET_B(net1052),
    .D(_0013_),
    .Q_N(_3026_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[15] ));
 sg13g2_dfrbp_1 _5991_ (.CLK(net965),
    .RESET_B(net1052),
    .D(_0014_),
    .Q_N(_3027_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[16] ));
 sg13g2_dfrbp_1 _5992_ (.CLK(net965),
    .RESET_B(net1052),
    .D(_0015_),
    .Q_N(_3028_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[17] ));
 sg13g2_dfrbp_1 _5993_ (.CLK(net968),
    .RESET_B(net1055),
    .D(_0016_),
    .Q_N(_3029_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[18] ));
 sg13g2_dfrbp_1 _5994_ (.CLK(net968),
    .RESET_B(net1055),
    .D(_0017_),
    .Q_N(_3030_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[19] ));
 sg13g2_dfrbp_1 _5995_ (.CLK(net959),
    .RESET_B(net1047),
    .D(_0019_),
    .Q_N(_3031_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[20] ));
 sg13g2_dfrbp_1 _5996_ (.CLK(net959),
    .RESET_B(net1047),
    .D(_0020_),
    .Q_N(_3032_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[21] ));
 sg13g2_dfrbp_1 _5997_ (.CLK(net959),
    .RESET_B(net1047),
    .D(_0021_),
    .Q_N(_3033_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[22] ));
 sg13g2_dfrbp_1 _5998_ (.CLK(net959),
    .RESET_B(net1047),
    .D(_0022_),
    .Q_N(_3034_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg1[23] ));
 sg13g2_dfrbp_1 _5999_ (.CLK(net943),
    .RESET_B(net1030),
    .D(_0031_),
    .Q_N(_3035_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[0] ));
 sg13g2_dfrbp_1 _6000_ (.CLK(net943),
    .RESET_B(net1030),
    .D(_0042_),
    .Q_N(_3036_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[1] ));
 sg13g2_dfrbp_1 _6001_ (.CLK(net943),
    .RESET_B(net1030),
    .D(_0051_),
    .Q_N(_3037_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[2] ));
 sg13g2_dfrbp_1 _6002_ (.CLK(net944),
    .RESET_B(net1031),
    .D(_0052_),
    .Q_N(_3038_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[3] ));
 sg13g2_dfrbp_1 _6003_ (.CLK(net950),
    .RESET_B(net1036),
    .D(_0053_),
    .Q_N(_3039_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[4] ));
 sg13g2_dfrbp_1 _6004_ (.CLK(net948),
    .RESET_B(net1035),
    .D(_0054_),
    .Q_N(_3040_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[5] ));
 sg13g2_dfrbp_1 _6005_ (.CLK(net948),
    .RESET_B(net1036),
    .D(_0055_),
    .Q_N(_3041_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[6] ));
 sg13g2_dfrbp_1 _6006_ (.CLK(net948),
    .RESET_B(net1035),
    .D(_0056_),
    .Q_N(_3042_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[7] ));
 sg13g2_dfrbp_1 _6007_ (.CLK(net949),
    .RESET_B(net1037),
    .D(_0057_),
    .Q_N(_3043_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[8] ));
 sg13g2_dfrbp_1 _6008_ (.CLK(net949),
    .RESET_B(net1037),
    .D(_0058_),
    .Q_N(_3044_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[9] ));
 sg13g2_dfrbp_1 _6009_ (.CLK(net949),
    .RESET_B(net1037),
    .D(_0032_),
    .Q_N(_3045_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[10] ));
 sg13g2_dfrbp_1 _6010_ (.CLK(net964),
    .RESET_B(net1053),
    .D(_0033_),
    .Q_N(_3046_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[11] ));
 sg13g2_dfrbp_1 _6011_ (.CLK(net965),
    .RESET_B(net1052),
    .D(_0034_),
    .Q_N(_3047_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[12] ));
 sg13g2_dfrbp_1 _6012_ (.CLK(net965),
    .RESET_B(net1052),
    .D(_0035_),
    .Q_N(_3048_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[13] ));
 sg13g2_dfrbp_1 _6013_ (.CLK(net965),
    .RESET_B(net1052),
    .D(_0036_),
    .Q_N(_3049_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[14] ));
 sg13g2_dfrbp_1 _6014_ (.CLK(net965),
    .RESET_B(net1052),
    .D(_0037_),
    .Q_N(_3050_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[15] ));
 sg13g2_dfrbp_1 _6015_ (.CLK(net970),
    .RESET_B(net1057),
    .D(_0038_),
    .Q_N(_3051_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[16] ));
 sg13g2_dfrbp_1 _6016_ (.CLK(net970),
    .RESET_B(net1057),
    .D(_0039_),
    .Q_N(_3052_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[17] ));
 sg13g2_dfrbp_1 _6017_ (.CLK(net968),
    .RESET_B(net1055),
    .D(_0040_),
    .Q_N(_3053_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[18] ));
 sg13g2_dfrbp_1 _6018_ (.CLK(net968),
    .RESET_B(net1055),
    .D(_0041_),
    .Q_N(_3054_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[19] ));
 sg13g2_dfrbp_1 _6019_ (.CLK(net968),
    .RESET_B(net1055),
    .D(_0043_),
    .Q_N(_3055_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[20] ));
 sg13g2_dfrbp_1 _6020_ (.CLK(net968),
    .RESET_B(net1055),
    .D(_0044_),
    .Q_N(_3056_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[21] ));
 sg13g2_dfrbp_1 _6021_ (.CLK(net959),
    .RESET_B(net1047),
    .D(_0045_),
    .Q_N(_3057_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[22] ));
 sg13g2_dfrbp_1 _6022_ (.CLK(net959),
    .RESET_B(net1047),
    .D(_0046_),
    .Q_N(_3058_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[23] ));
 sg13g2_dfrbp_1 _6023_ (.CLK(net959),
    .RESET_B(net1047),
    .D(_0047_),
    .Q_N(_3059_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[24] ));
 sg13g2_dfrbp_1 _6024_ (.CLK(net957),
    .RESET_B(net1045),
    .D(_0048_),
    .Q_N(_3060_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[25] ));
 sg13g2_dfrbp_1 _6025_ (.CLK(net957),
    .RESET_B(net1045),
    .D(_0049_),
    .Q_N(_3061_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[26] ));
 sg13g2_dfrbp_1 _6026_ (.CLK(net957),
    .RESET_B(net1045),
    .D(_0050_),
    .Q_N(_2675_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg2[27] ));
 sg13g2_dfrbp_1 _6027_ (.CLK(_0346_),
    .RESET_B(net1028),
    .D(_0609_),
    .Q_N(_2674_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg1[0] ));
 sg13g2_dfrbp_1 _6028_ (.CLK(_0347_),
    .RESET_B(net1020),
    .D(_0610_),
    .Q_N(_2673_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg1[1] ));
 sg13g2_dfrbp_1 _6029_ (.CLK(_0348_),
    .RESET_B(net1020),
    .D(_0611_),
    .Q_N(_2672_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg1[2] ));
 sg13g2_dfrbp_1 _6030_ (.CLK(_0349_),
    .RESET_B(net1021),
    .D(_0612_),
    .Q_N(_2671_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg1[3] ));
 sg13g2_dfrbp_1 _6031_ (.CLK(_0350_),
    .RESET_B(net1021),
    .D(_0613_),
    .Q_N(_2670_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg1[4] ));
 sg13g2_dfrbp_1 _6032_ (.CLK(_0351_),
    .RESET_B(net1021),
    .D(_0614_),
    .Q_N(_2669_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg1[5] ));
 sg13g2_dfrbp_1 _6033_ (.CLK(_0352_),
    .RESET_B(net1026),
    .D(_0615_),
    .Q_N(_2668_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg1[6] ));
 sg13g2_dfrbp_1 _6034_ (.CLK(_0353_),
    .RESET_B(net1026),
    .D(_0616_),
    .Q_N(_2667_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg1[7] ));
 sg13g2_dfrbp_1 _6035_ (.CLK(_0354_),
    .RESET_B(net1026),
    .D(_0617_),
    .Q_N(_2666_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg1[8] ));
 sg13g2_dfrbp_1 _6036_ (.CLK(_0355_),
    .RESET_B(net1025),
    .D(_0618_),
    .Q_N(_2665_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg1[9] ));
 sg13g2_dfrbp_1 _6037_ (.CLK(_0356_),
    .RESET_B(net1025),
    .D(_0619_),
    .Q_N(_2664_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg1[10] ));
 sg13g2_dfrbp_1 _6038_ (.CLK(_0357_),
    .RESET_B(net1025),
    .D(_0620_),
    .Q_N(_2663_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg1[11] ));
 sg13g2_dfrbp_1 _6039_ (.CLK(_0358_),
    .RESET_B(net1043),
    .D(_0621_),
    .Q_N(_2662_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg1[12] ));
 sg13g2_dfrbp_1 _6040_ (.CLK(_0359_),
    .RESET_B(net1043),
    .D(_0622_),
    .Q_N(_2661_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg1[13] ));
 sg13g2_dfrbp_1 _6041_ (.CLK(_0360_),
    .RESET_B(net1040),
    .D(_0623_),
    .Q_N(_2660_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg1[14] ));
 sg13g2_dfrbp_1 _6042_ (.CLK(_0361_),
    .RESET_B(net1041),
    .D(_0624_),
    .Q_N(_2659_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg1[15] ));
 sg13g2_dfrbp_1 _6043_ (.CLK(_0362_),
    .RESET_B(net1041),
    .D(_0625_),
    .Q_N(_2658_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg1[16] ));
 sg13g2_dfrbp_1 _6044_ (.CLK(net943),
    .RESET_B(net1030),
    .D(_0626_),
    .Q_N(_2657_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg0[0] ));
 sg13g2_dfrbp_1 _6045_ (.CLK(net943),
    .RESET_B(net1030),
    .D(_0627_),
    .Q_N(_2656_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg0[1] ));
 sg13g2_dfrbp_1 _6046_ (.CLK(net944),
    .RESET_B(net1031),
    .D(_0628_),
    .Q_N(_2655_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg0[2] ));
 sg13g2_dfrbp_1 _6047_ (.CLK(net944),
    .RESET_B(net1031),
    .D(_0629_),
    .Q_N(_2654_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg0[3] ));
 sg13g2_dfrbp_1 _6048_ (.CLK(net944),
    .RESET_B(net1035),
    .D(_0630_),
    .Q_N(_2653_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg0[4] ));
 sg13g2_dfrbp_1 _6049_ (.CLK(net948),
    .RESET_B(net1035),
    .D(_0631_),
    .Q_N(_2652_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg0[5] ));
 sg13g2_dfrbp_1 _6050_ (.CLK(net948),
    .RESET_B(net1035),
    .D(_0632_),
    .Q_N(_2651_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg0[6] ));
 sg13g2_dfrbp_1 _6051_ (.CLK(net948),
    .RESET_B(net1035),
    .D(_0633_),
    .Q_N(_2650_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg0[7] ));
 sg13g2_dfrbp_1 _6052_ (.CLK(net949),
    .RESET_B(net1037),
    .D(_0634_),
    .Q_N(_2649_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg0[8] ));
 sg13g2_dfrbp_1 _6053_ (.CLK(net949),
    .RESET_B(net1037),
    .D(_0635_),
    .Q_N(_2648_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg0[9] ));
 sg13g2_dfrbp_1 _6054_ (.CLK(net949),
    .RESET_B(net1037),
    .D(_0636_),
    .Q_N(_2647_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg0[10] ));
 sg13g2_dfrbp_1 _6055_ (.CLK(net964),
    .RESET_B(net1053),
    .D(_0637_),
    .Q_N(_2646_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg0[11] ));
 sg13g2_dfrbp_1 _6056_ (.CLK(net964),
    .RESET_B(net1053),
    .D(_0638_),
    .Q_N(_2645_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg0[12] ));
 sg13g2_dfrbp_1 _6057_ (.CLK(net964),
    .RESET_B(net1053),
    .D(_0639_),
    .Q_N(_2644_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg0[13] ));
 sg13g2_dfrbp_1 _6058_ (.CLK(net965),
    .RESET_B(net1052),
    .D(_0640_),
    .Q_N(_2643_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg0[14] ));
 sg13g2_dfrbp_1 _6059_ (.CLK(net964),
    .RESET_B(net1053),
    .D(_0641_),
    .Q_N(_2642_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg0[15] ));
 sg13g2_dfrbp_1 _6060_ (.CLK(net963),
    .RESET_B(net1051),
    .D(_0642_),
    .Q_N(_2641_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg0[16] ));
 sg13g2_dfrbp_1 _6061_ (.CLK(net967),
    .RESET_B(net1054),
    .D(_0643_),
    .Q_N(_2640_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg0[17] ));
 sg13g2_dfrbp_1 _6062_ (.CLK(net963),
    .RESET_B(net1051),
    .D(_0644_),
    .Q_N(_2639_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg0[18] ));
 sg13g2_dfrbp_1 _6063_ (.CLK(net967),
    .RESET_B(net1055),
    .D(_0645_),
    .Q_N(_2638_),
    .Q(\u_ddc_top_level.cic_left_inst.int_reg0[19] ));
 sg13g2_dfrbp_1 _6064_ (.CLK(_0363_),
    .RESET_B(net1028),
    .D(_0646_),
    .Q_N(_2637_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg2[0] ));
 sg13g2_dfrbp_1 _6065_ (.CLK(_0364_),
    .RESET_B(net1028),
    .D(_0647_),
    .Q_N(_2636_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg2[1] ));
 sg13g2_dfrbp_1 _6066_ (.CLK(_0365_),
    .RESET_B(net1028),
    .D(_0648_),
    .Q_N(_2635_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg2[2] ));
 sg13g2_dfrbp_1 _6067_ (.CLK(_0366_),
    .RESET_B(net1029),
    .D(_0649_),
    .Q_N(_2634_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg2[3] ));
 sg13g2_dfrbp_1 _6068_ (.CLK(_0367_),
    .RESET_B(net1029),
    .D(_0650_),
    .Q_N(_2633_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg2[4] ));
 sg13g2_dfrbp_1 _6069_ (.CLK(_0368_),
    .RESET_B(net1029),
    .D(_0651_),
    .Q_N(_2632_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg2[5] ));
 sg13g2_dfrbp_1 _6070_ (.CLK(_0369_),
    .RESET_B(net1033),
    .D(_0652_),
    .Q_N(_2631_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg2[6] ));
 sg13g2_dfrbp_1 _6071_ (.CLK(_0370_),
    .RESET_B(net1033),
    .D(_0653_),
    .Q_N(_2630_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg2[7] ));
 sg13g2_dfrbp_1 _6072_ (.CLK(_0371_),
    .RESET_B(net1034),
    .D(_0654_),
    .Q_N(_2629_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg2[8] ));
 sg13g2_dfrbp_1 _6073_ (.CLK(_0372_),
    .RESET_B(net1025),
    .D(_0655_),
    .Q_N(_2628_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg2[9] ));
 sg13g2_dfrbp_1 _6074_ (.CLK(_0373_),
    .RESET_B(net1034),
    .D(_0656_),
    .Q_N(_2627_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg2[10] ));
 sg13g2_dfrbp_1 _6075_ (.CLK(_0374_),
    .RESET_B(net1025),
    .D(_0657_),
    .Q_N(_2626_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg2[11] ));
 sg13g2_dfrbp_1 _6076_ (.CLK(_0375_),
    .RESET_B(net1043),
    .D(_0658_),
    .Q_N(_2625_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg2[12] ));
 sg13g2_dfrbp_1 _6077_ (.CLK(_0376_),
    .RESET_B(net1043),
    .D(_0659_),
    .Q_N(_2624_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg2[13] ));
 sg13g2_dfrbp_1 _6078_ (.CLK(_0377_),
    .RESET_B(net1044),
    .D(_0660_),
    .Q_N(_2623_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg2[14] ));
 sg13g2_dfrbp_1 _6079_ (.CLK(_0378_),
    .RESET_B(net1043),
    .D(_0661_),
    .Q_N(_2622_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg2[15] ));
 sg13g2_dfrbp_1 _6080_ (.CLK(_0379_),
    .RESET_B(net1044),
    .D(_0662_),
    .Q_N(_2621_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg2[16] ));
 sg13g2_dfrbp_1 _6081_ (.CLK(_0380_),
    .RESET_B(net1044),
    .D(_0663_),
    .Q_N(_3062_),
    .Q(\u_ddc_top_level.cic_left_inst.comb_reg2[17] ));
 sg13g2_dfrbp_1 _6082_ (.CLK(net921),
    .RESET_B(net1008),
    .D(net1),
    .Q_N(_2620_),
    .Q(\u_ddc_top_level.i2s_rx_inst.lrclk_prev ));
 sg13g2_dfrbp_1 _6083_ (.CLK(_0381_),
    .RESET_B(net977),
    .D(_0664_),
    .Q_N(_2619_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out0[0] ));
 sg13g2_dfrbp_1 _6084_ (.CLK(_0382_),
    .RESET_B(net976),
    .D(_0665_),
    .Q_N(_2618_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out0[1] ));
 sg13g2_dfrbp_1 _6085_ (.CLK(_0383_),
    .RESET_B(net985),
    .D(_0666_),
    .Q_N(_2617_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out0[2] ));
 sg13g2_dfrbp_1 _6086_ (.CLK(_0384_),
    .RESET_B(net986),
    .D(_0667_),
    .Q_N(_2616_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out0[3] ));
 sg13g2_dfrbp_1 _6087_ (.CLK(_0385_),
    .RESET_B(net985),
    .D(_0668_),
    .Q_N(_2615_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out0[4] ));
 sg13g2_dfrbp_1 _6088_ (.CLK(_0386_),
    .RESET_B(net985),
    .D(_0669_),
    .Q_N(_2614_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out0[5] ));
 sg13g2_dfrbp_1 _6089_ (.CLK(_0387_),
    .RESET_B(net988),
    .D(_0670_),
    .Q_N(_2613_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out0[6] ));
 sg13g2_dfrbp_1 _6090_ (.CLK(_0388_),
    .RESET_B(net988),
    .D(_0671_),
    .Q_N(_2612_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out0[7] ));
 sg13g2_dfrbp_1 _6091_ (.CLK(_0389_),
    .RESET_B(net992),
    .D(_0672_),
    .Q_N(_2611_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out0[8] ));
 sg13g2_dfrbp_1 _6092_ (.CLK(_0390_),
    .RESET_B(net992),
    .D(_0673_),
    .Q_N(_2610_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out0[9] ));
 sg13g2_dfrbp_1 _6093_ (.CLK(_0391_),
    .RESET_B(net992),
    .D(_0674_),
    .Q_N(_2609_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out0[10] ));
 sg13g2_dfrbp_1 _6094_ (.CLK(_0392_),
    .RESET_B(net993),
    .D(_0675_),
    .Q_N(_2608_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out0[11] ));
 sg13g2_dfrbp_1 _6095_ (.CLK(_0393_),
    .RESET_B(net993),
    .D(_0676_),
    .Q_N(_2607_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out0[12] ));
 sg13g2_dfrbp_1 _6096_ (.CLK(_0394_),
    .RESET_B(net1007),
    .D(_0677_),
    .Q_N(_2606_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out0[13] ));
 sg13g2_dfrbp_1 _6097_ (.CLK(_0395_),
    .RESET_B(net1007),
    .D(_0678_),
    .Q_N(_2605_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out0[14] ));
 sg13g2_dfrbp_1 _6098_ (.CLK(_0396_),
    .RESET_B(net1008),
    .D(_0679_),
    .Q_N(_2604_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out0[15] ));
 sg13g2_dfrbp_1 _6099_ (.CLK(_0397_),
    .RESET_B(net1008),
    .D(_0680_),
    .Q_N(_2603_),
    .Q(\u_ddc_top_level.cic_right_inst.comb_out0[16] ));
 sg13g2_dfrbp_1 _6100_ (.CLK(net922),
    .RESET_B(net1009),
    .D(_0681_),
    .Q_N(_2602_),
    .Q(\u_ddc_top_level.cic_right_inst.in_valid ));
 sg13g2_dfrbp_1 _6101_ (.CLK(net929),
    .RESET_B(net1017),
    .D(_0682_),
    .Q_N(_2601_),
    .Q(\u_ddc_top_level.cic_left_inst.in_data[0] ));
 sg13g2_dfrbp_1 _6102_ (.CLK(net930),
    .RESET_B(net1018),
    .D(_0683_),
    .Q_N(_2600_),
    .Q(\u_ddc_top_level.cic_left_inst.in_data[1] ));
 sg13g2_dfrbp_1 _6103_ (.CLK(net930),
    .RESET_B(net1018),
    .D(_0684_),
    .Q_N(_2599_),
    .Q(\u_ddc_top_level.cic_left_inst.in_data[2] ));
 sg13g2_dfrbp_1 _6104_ (.CLK(net929),
    .RESET_B(net1017),
    .D(_0685_),
    .Q_N(_2598_),
    .Q(\u_ddc_top_level.cic_left_inst.in_data[3] ));
 sg13g2_dfrbp_1 _6105_ (.CLK(net929),
    .RESET_B(net1017),
    .D(_0686_),
    .Q_N(_2597_),
    .Q(\u_ddc_top_level.cic_left_inst.in_data[4] ));
 sg13g2_dfrbp_1 _6106_ (.CLK(net931),
    .RESET_B(net1019),
    .D(_0687_),
    .Q_N(_2596_),
    .Q(\u_ddc_top_level.cic_left_inst.in_data[5] ));
 sg13g2_dfrbp_1 _6107_ (.CLK(net931),
    .RESET_B(net1019),
    .D(_0688_),
    .Q_N(_2595_),
    .Q(\u_ddc_top_level.cic_left_inst.in_data[6] ));
 sg13g2_dfrbp_1 _6108_ (.CLK(net931),
    .RESET_B(net1023),
    .D(_0689_),
    .Q_N(_2594_),
    .Q(\u_ddc_top_level.cic_left_inst.in_data[7] ));
 sg13g2_dfrbp_1 _6109_ (.CLK(net936),
    .RESET_B(net1023),
    .D(_0690_),
    .Q_N(_2593_),
    .Q(\u_ddc_top_level.cic_left_inst.in_data[8] ));
 sg13g2_dfrbp_1 _6110_ (.CLK(net936),
    .RESET_B(net1023),
    .D(_0691_),
    .Q_N(_2592_),
    .Q(\u_ddc_top_level.cic_left_inst.in_data[9] ));
 sg13g2_dfrbp_1 _6111_ (.CLK(net937),
    .RESET_B(net1024),
    .D(_0692_),
    .Q_N(_2591_),
    .Q(\u_ddc_top_level.cic_left_inst.in_data[10] ));
 sg13g2_dfrbp_1 _6112_ (.CLK(net937),
    .RESET_B(net1024),
    .D(_0693_),
    .Q_N(_2590_),
    .Q(\u_ddc_top_level.cic_left_inst.in_data[11] ));
 sg13g2_dfrbp_1 _6113_ (.CLK(net952),
    .RESET_B(net1040),
    .D(_0694_),
    .Q_N(_2589_),
    .Q(\u_ddc_top_level.cic_left_inst.in_data[12] ));
 sg13g2_dfrbp_1 _6114_ (.CLK(net952),
    .RESET_B(net1040),
    .D(_0695_),
    .Q_N(_2588_),
    .Q(\u_ddc_top_level.cic_left_inst.in_data[13] ));
 sg13g2_dfrbp_1 _6115_ (.CLK(net952),
    .RESET_B(net1040),
    .D(_0696_),
    .Q_N(_2587_),
    .Q(\u_ddc_top_level.cic_left_inst.in_data[14] ));
 sg13g2_dfrbp_1 _6116_ (.CLK(net953),
    .RESET_B(net1041),
    .D(_0697_),
    .Q_N(_3063_),
    .Q(\u_ddc_top_level.cic_left_inst.in_data[15] ));
 sg13g2_dfrbp_1 _6117_ (.CLK(net957),
    .RESET_B(net1045),
    .D(_0000_),
    .Q_N(_3064_),
    .Q(\u_ddc_top_level.i2s_rx_inst.bit_count[0] ));
 sg13g2_dfrbp_1 _6118_ (.CLK(net957),
    .RESET_B(net1045),
    .D(_0001_),
    .Q_N(_3065_),
    .Q(\u_ddc_top_level.i2s_rx_inst.bit_count[1] ));
 sg13g2_dfrbp_1 _6119_ (.CLK(net957),
    .RESET_B(net1045),
    .D(_0002_),
    .Q_N(_3066_),
    .Q(\u_ddc_top_level.i2s_rx_inst.bit_count[2] ));
 sg13g2_dfrbp_1 _6120_ (.CLK(net957),
    .RESET_B(net1045),
    .D(_0003_),
    .Q_N(_3067_),
    .Q(\u_ddc_top_level.i2s_rx_inst.bit_count[3] ));
 sg13g2_dfrbp_1 _6121_ (.CLK(net953),
    .RESET_B(net1041),
    .D(_0004_),
    .Q_N(_3068_),
    .Q(\u_ddc_top_level.i2s_rx_inst.bit_count[4] ));
 sg13g2_dfrbp_1 _6122_ (.CLK(net953),
    .RESET_B(net1041),
    .D(_0005_),
    .Q_N(_2586_),
    .Q(\u_ddc_top_level.i2s_rx_inst.bit_count[5] ));
 sg13g2_dfrbp_1 _6123_ (.CLK(net900),
    .RESET_B(net987),
    .D(_0698_),
    .Q_N(_2585_),
    .Q(\u_ddc_top_level.cic_right_inst.in_data[0] ));
 sg13g2_dfrbp_1 _6124_ (.CLK(net900),
    .RESET_B(net987),
    .D(_0699_),
    .Q_N(_2584_),
    .Q(\u_ddc_top_level.cic_right_inst.in_data[1] ));
 sg13g2_dfrbp_1 _6125_ (.CLK(net900),
    .RESET_B(net987),
    .D(_0700_),
    .Q_N(_2583_),
    .Q(\u_ddc_top_level.cic_right_inst.in_data[2] ));
 sg13g2_dfrbp_1 _6126_ (.CLK(net901),
    .RESET_B(net987),
    .D(_0701_),
    .Q_N(_2582_),
    .Q(\u_ddc_top_level.cic_right_inst.in_data[3] ));
 sg13g2_dfrbp_1 _6127_ (.CLK(net900),
    .RESET_B(net987),
    .D(_0702_),
    .Q_N(_2581_),
    .Q(\u_ddc_top_level.cic_right_inst.in_data[4] ));
 sg13g2_dfrbp_1 _6128_ (.CLK(net902),
    .RESET_B(net988),
    .D(_0703_),
    .Q_N(_2580_),
    .Q(\u_ddc_top_level.cic_right_inst.in_data[5] ));
 sg13g2_dfrbp_1 _6129_ (.CLK(net901),
    .RESET_B(net988),
    .D(_0704_),
    .Q_N(_2579_),
    .Q(\u_ddc_top_level.cic_right_inst.in_data[6] ));
 sg13g2_dfrbp_1 _6130_ (.CLK(net901),
    .RESET_B(net988),
    .D(_0705_),
    .Q_N(_2578_),
    .Q(\u_ddc_top_level.cic_right_inst.in_data[7] ));
 sg13g2_dfrbp_1 _6131_ (.CLK(net905),
    .RESET_B(net992),
    .D(_0706_),
    .Q_N(_2577_),
    .Q(\u_ddc_top_level.cic_right_inst.in_data[8] ));
 sg13g2_dfrbp_1 _6132_ (.CLK(net905),
    .RESET_B(net992),
    .D(_0707_),
    .Q_N(_2576_),
    .Q(\u_ddc_top_level.cic_right_inst.in_data[9] ));
 sg13g2_dfrbp_1 _6133_ (.CLK(net905),
    .RESET_B(net993),
    .D(_0708_),
    .Q_N(_2575_),
    .Q(\u_ddc_top_level.cic_right_inst.in_data[10] ));
 sg13g2_dfrbp_1 _6134_ (.CLK(net906),
    .RESET_B(net993),
    .D(_0709_),
    .Q_N(_2574_),
    .Q(\u_ddc_top_level.cic_right_inst.in_data[11] ));
 sg13g2_dfrbp_1 _6135_ (.CLK(net906),
    .RESET_B(net1007),
    .D(_0710_),
    .Q_N(_2573_),
    .Q(\u_ddc_top_level.cic_right_inst.in_data[12] ));
 sg13g2_dfrbp_1 _6136_ (.CLK(net920),
    .RESET_B(net1007),
    .D(_0711_),
    .Q_N(_2572_),
    .Q(\u_ddc_top_level.cic_right_inst.in_data[13] ));
 sg13g2_dfrbp_1 _6137_ (.CLK(net921),
    .RESET_B(net1009),
    .D(_0712_),
    .Q_N(_2571_),
    .Q(\u_ddc_top_level.cic_right_inst.in_data[14] ));
 sg13g2_dfrbp_1 _6138_ (.CLK(net921),
    .RESET_B(net1008),
    .D(_0713_),
    .Q_N(_2570_),
    .Q(\u_ddc_top_level.cic_right_inst.in_data[15] ));
 sg13g2_dfrbp_1 _6139_ (.CLK(net929),
    .RESET_B(net1017),
    .D(_0714_),
    .Q_N(_2569_),
    .Q(\u_ddc_top_level.cic_left_inst.in_valid ));
 sg13g2_tielo tt_um_ddc_arghunter_5 (.L_LO(net5));
 sg13g2_tielo tt_um_ddc_arghunter_6 (.L_LO(net6));
 sg13g2_tielo tt_um_ddc_arghunter_7 (.L_LO(net7));
 sg13g2_tielo tt_um_ddc_arghunter_8 (.L_LO(net8));
 sg13g2_tielo tt_um_ddc_arghunter_9 (.L_LO(net9));
 sg13g2_tielo tt_um_ddc_arghunter_10 (.L_LO(net10));
 sg13g2_tielo tt_um_ddc_arghunter_11 (.L_LO(net11));
 sg13g2_tielo tt_um_ddc_arghunter_12 (.L_LO(net12));
 sg13g2_tielo tt_um_ddc_arghunter_13 (.L_LO(net13));
 sg13g2_tielo tt_um_ddc_arghunter_14 (.L_LO(net14));
 sg13g2_tielo tt_um_ddc_arghunter_15 (.L_LO(net15));
 sg13g2_tielo tt_um_ddc_arghunter_16 (.L_LO(net16));
 sg13g2_tielo tt_um_ddc_arghunter_17 (.L_LO(net17));
 sg13g2_tielo tt_um_ddc_arghunter_18 (.L_LO(net18));
 sg13g2_tielo tt_um_ddc_arghunter_19 (.L_LO(net19));
 sg13g2_tielo tt_um_ddc_arghunter_20 (.L_LO(net20));
 sg13g2_tielo tt_um_ddc_arghunter_21 (.L_LO(net21));
 sg13g2_tielo tt_um_ddc_arghunter_22 (.L_LO(net22));
 sg13g2_tielo tt_um_ddc_arghunter_23 (.L_LO(net23));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_buf_2 _6160_ (.A(\u_ddc_top_level.dsm_left_inst.out_bitstream ),
    .X(uo_out[0]));
 sg13g2_buf_1 _6161_ (.A(\u_ddc_top_level.dsm_right_inst.out_bitstream ),
    .X(uo_out[1]));
 sg13g2_buf_1 _6162_ (.A(net923),
    .X(uo_out[2]));
 sg13g2_buf_1 _6163_ (.A(net915),
    .X(uo_out[3]));
 sg13g2_buf_4 fanout806 (.X(net806),
    .A(net807));
 sg13g2_buf_4 fanout807 (.X(net807),
    .A(_2313_));
 sg13g2_buf_4 fanout808 (.X(net808),
    .A(net811));
 sg13g2_buf_1 fanout809 (.A(net811),
    .X(net809));
 sg13g2_buf_2 fanout810 (.A(net811),
    .X(net810));
 sg13g2_buf_2 fanout811 (.A(net812),
    .X(net811));
 sg13g2_buf_4 fanout812 (.X(net812),
    .A(_0719_));
 sg13g2_buf_4 fanout813 (.X(net813),
    .A(_0715_));
 sg13g2_buf_2 fanout814 (.A(_0715_),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(net816),
    .X(net815));
 sg13g2_buf_2 fanout816 (.A(net817),
    .X(net816));
 sg13g2_buf_4 fanout817 (.X(net817),
    .A(_0715_));
 sg13g2_buf_4 fanout818 (.X(net818),
    .A(net820));
 sg13g2_buf_4 fanout819 (.X(net819),
    .A(net820));
 sg13g2_buf_2 fanout820 (.A(_1399_),
    .X(net820));
 sg13g2_buf_4 fanout821 (.X(net821),
    .A(net823));
 sg13g2_buf_4 fanout822 (.X(net822),
    .A(net823));
 sg13g2_buf_4 fanout823 (.X(net823),
    .A(_1398_));
 sg13g2_buf_4 fanout824 (.X(net824),
    .A(net826));
 sg13g2_buf_2 fanout825 (.A(net826),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(net838),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(net828),
    .X(net827));
 sg13g2_buf_4 fanout828 (.X(net828),
    .A(net838));
 sg13g2_buf_2 fanout829 (.A(net833),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(net833),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(net833),
    .X(net831));
 sg13g2_buf_1 fanout832 (.A(net833),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(net838),
    .X(net833));
 sg13g2_buf_4 fanout834 (.X(net834),
    .A(net837));
 sg13g2_buf_2 fanout835 (.A(net837),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(net837),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(net838),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(\u_ddc_top_level.cic_left_inst.in_valid ),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(net841),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(net841),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(net851),
    .X(net841));
 sg13g2_buf_4 fanout842 (.X(net842),
    .A(net843));
 sg13g2_buf_4 fanout843 (.X(net843),
    .A(net851));
 sg13g2_buf_2 fanout844 (.A(net850),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(net850),
    .X(net845));
 sg13g2_buf_4 fanout846 (.X(net846),
    .A(net850));
 sg13g2_buf_2 fanout847 (.A(net849),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(net849),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(net850),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(net851),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(\u_ddc_top_level.cic_left_inst.in_valid ),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(net853),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(net863),
    .X(net853));
 sg13g2_buf_4 fanout854 (.X(net854),
    .A(net857));
 sg13g2_buf_2 fanout855 (.A(net857),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(net857),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(net863),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(net862),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(net862),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(net861),
    .X(net860));
 sg13g2_buf_4 fanout861 (.X(net861),
    .A(net862));
 sg13g2_buf_2 fanout862 (.A(net863),
    .X(net862));
 sg13g2_buf_2 fanout863 (.A(\u_ddc_top_level.cic_right_inst.in_valid ),
    .X(net863));
 sg13g2_buf_4 fanout864 (.X(net864),
    .A(net868));
 sg13g2_buf_2 fanout865 (.A(net868),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(net868),
    .X(net866));
 sg13g2_buf_1 fanout867 (.A(net868),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(net878),
    .X(net868));
 sg13g2_buf_4 fanout869 (.X(net869),
    .A(net871));
 sg13g2_buf_2 fanout870 (.A(net871),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(net878),
    .X(net871));
 sg13g2_buf_4 fanout872 (.X(net872),
    .A(net878));
 sg13g2_buf_2 fanout873 (.A(net878),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(net875),
    .X(net874));
 sg13g2_buf_4 fanout875 (.X(net875),
    .A(net877));
 sg13g2_buf_4 fanout876 (.X(net876),
    .A(net877));
 sg13g2_buf_2 fanout877 (.A(net878),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(\u_ddc_top_level.cic_right_inst.in_valid ),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(\u_ddc_top_level.cic_left_inst.int_reg0[19] ),
    .X(net879));
 sg13g2_buf_1 fanout880 (.A(\u_ddc_top_level.cic_left_inst.int_reg0[19] ),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(\u_ddc_top_level.cic_left_inst.int_reg1[23] ),
    .X(net881));
 sg13g2_buf_4 fanout882 (.X(net882),
    .A(\u_ddc_top_level.cic_right_inst.int_reg0[19] ));
 sg13g2_buf_1 fanout883 (.A(\u_ddc_top_level.cic_right_inst.int_reg0[19] ),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(\u_ddc_top_level.cic_right_inst.int_reg1[23] ),
    .X(net884));
 sg13g2_buf_4 fanout885 (.X(net885),
    .A(net886));
 sg13g2_buf_4 fanout886 (.X(net886),
    .A(net3));
 sg13g2_buf_2 fanout887 (.A(net889),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(net889),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(net892),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(net891),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(net892),
    .X(net891));
 sg13g2_buf_1 fanout892 (.A(net908),
    .X(net892));
 sg13g2_buf_2 fanout893 (.A(net894),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(net897),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(net897),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(net897),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(net908),
    .X(net897));
 sg13g2_buf_2 fanout898 (.A(net899),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(net902),
    .X(net899));
 sg13g2_buf_2 fanout900 (.A(net901),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(net902),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(net908),
    .X(net902));
 sg13g2_buf_2 fanout903 (.A(net904),
    .X(net903));
 sg13g2_buf_2 fanout904 (.A(net907),
    .X(net904));
 sg13g2_buf_2 fanout905 (.A(net906),
    .X(net905));
 sg13g2_buf_2 fanout906 (.A(net907),
    .X(net906));
 sg13g2_buf_2 fanout907 (.A(net908),
    .X(net907));
 sg13g2_buf_2 fanout908 (.A(ui_in[0]),
    .X(net908));
 sg13g2_buf_2 fanout909 (.A(net913),
    .X(net909));
 sg13g2_buf_2 fanout910 (.A(net913),
    .X(net910));
 sg13g2_buf_2 fanout911 (.A(net913),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(net913),
    .X(net912));
 sg13g2_buf_2 fanout913 (.A(net928),
    .X(net913));
 sg13g2_buf_2 fanout914 (.A(net917),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(net917),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(net917),
    .X(net916));
 sg13g2_buf_2 fanout917 (.A(net928),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(net922),
    .X(net918));
 sg13g2_buf_1 fanout919 (.A(net922),
    .X(net919));
 sg13g2_buf_2 fanout920 (.A(net921),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(net922),
    .X(net921));
 sg13g2_buf_2 fanout922 (.A(net928),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(net924),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(net928),
    .X(net924));
 sg13g2_buf_2 fanout925 (.A(net927),
    .X(net925));
 sg13g2_buf_2 fanout926 (.A(net927),
    .X(net926));
 sg13g2_buf_2 fanout927 (.A(net928),
    .X(net927));
 sg13g2_buf_2 fanout928 (.A(ui_in[0]),
    .X(net928));
 sg13g2_buf_2 fanout929 (.A(net932),
    .X(net929));
 sg13g2_buf_1 fanout930 (.A(net932),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(net932),
    .X(net931));
 sg13g2_buf_1 fanout932 (.A(net935),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(net934),
    .X(net933));
 sg13g2_buf_2 fanout934 (.A(net935),
    .X(net934));
 sg13g2_buf_1 fanout935 (.A(net973),
    .X(net935));
 sg13g2_buf_2 fanout936 (.A(net940),
    .X(net936));
 sg13g2_buf_2 fanout937 (.A(net940),
    .X(net937));
 sg13g2_buf_2 fanout938 (.A(net940),
    .X(net938));
 sg13g2_buf_2 fanout939 (.A(net940),
    .X(net939));
 sg13g2_buf_1 fanout940 (.A(net973),
    .X(net940));
 sg13g2_buf_2 fanout941 (.A(net942),
    .X(net941));
 sg13g2_buf_2 fanout942 (.A(net945),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(net945),
    .X(net943));
 sg13g2_buf_1 fanout944 (.A(net945),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(net951),
    .X(net945));
 sg13g2_buf_2 fanout946 (.A(net951),
    .X(net946));
 sg13g2_buf_1 fanout947 (.A(net951),
    .X(net947));
 sg13g2_buf_2 fanout948 (.A(net950),
    .X(net948));
 sg13g2_buf_2 fanout949 (.A(net950),
    .X(net949));
 sg13g2_buf_2 fanout950 (.A(net951),
    .X(net950));
 sg13g2_buf_2 fanout951 (.A(net973),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(net954),
    .X(net952));
 sg13g2_buf_2 fanout953 (.A(net954),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(net962),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(net962),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(net962),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(net961),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(net961),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(net961),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(net961),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(net962),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(net973),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(net967),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(net966),
    .X(net964));
 sg13g2_buf_2 fanout965 (.A(net966),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(net967),
    .X(net966));
 sg13g2_buf_1 fanout967 (.A(net972),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(net972),
    .X(net968));
 sg13g2_buf_1 fanout969 (.A(net972),
    .X(net969));
 sg13g2_buf_2 fanout970 (.A(net971),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(net972),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(net973),
    .X(net972));
 sg13g2_buf_4 fanout973 (.X(net973),
    .A(ui_in[0]));
 sg13g2_buf_4 fanout974 (.X(net974),
    .A(net975));
 sg13g2_buf_4 fanout975 (.X(net975),
    .A(net978));
 sg13g2_buf_4 fanout976 (.X(net976),
    .A(net977));
 sg13g2_buf_4 fanout977 (.X(net977),
    .A(net978));
 sg13g2_buf_4 fanout978 (.X(net978),
    .A(net984));
 sg13g2_buf_4 fanout979 (.X(net979),
    .A(net981));
 sg13g2_buf_4 fanout980 (.X(net980),
    .A(net981));
 sg13g2_buf_2 fanout981 (.A(net984),
    .X(net981));
 sg13g2_buf_4 fanout982 (.X(net982),
    .A(net984));
 sg13g2_buf_2 fanout983 (.A(net984),
    .X(net983));
 sg13g2_buf_2 fanout984 (.A(net1016),
    .X(net984));
 sg13g2_buf_4 fanout985 (.X(net985),
    .A(net986));
 sg13g2_buf_4 fanout986 (.X(net986),
    .A(net989));
 sg13g2_buf_4 fanout987 (.X(net987),
    .A(net989));
 sg13g2_buf_4 fanout988 (.X(net988),
    .A(net989));
 sg13g2_buf_2 fanout989 (.A(net994),
    .X(net989));
 sg13g2_buf_4 fanout990 (.X(net990),
    .A(net991));
 sg13g2_buf_4 fanout991 (.X(net991),
    .A(net994));
 sg13g2_buf_4 fanout992 (.X(net992),
    .A(net994));
 sg13g2_buf_4 fanout993 (.X(net993),
    .A(net994));
 sg13g2_buf_2 fanout994 (.A(net1016),
    .X(net994));
 sg13g2_buf_4 fanout995 (.X(net995),
    .A(net1004));
 sg13g2_buf_4 fanout996 (.X(net996),
    .A(net1004));
 sg13g2_buf_4 fanout997 (.X(net997),
    .A(net999));
 sg13g2_buf_4 fanout998 (.X(net998),
    .A(net999));
 sg13g2_buf_2 fanout999 (.A(net1004),
    .X(net999));
 sg13g2_buf_4 fanout1000 (.X(net1000),
    .A(net1003));
 sg13g2_buf_4 fanout1001 (.X(net1001),
    .A(net1003));
 sg13g2_buf_4 fanout1002 (.X(net1002),
    .A(net1003));
 sg13g2_buf_4 fanout1003 (.X(net1003),
    .A(net1004));
 sg13g2_buf_2 fanout1004 (.A(net1016),
    .X(net1004));
 sg13g2_buf_4 fanout1005 (.X(net1005),
    .A(net1015));
 sg13g2_buf_4 fanout1006 (.X(net1006),
    .A(net1015));
 sg13g2_buf_4 fanout1007 (.X(net1007),
    .A(net1009));
 sg13g2_buf_4 fanout1008 (.X(net1008),
    .A(net1009));
 sg13g2_buf_2 fanout1009 (.A(net1015),
    .X(net1009));
 sg13g2_buf_4 fanout1010 (.X(net1010),
    .A(net1011));
 sg13g2_buf_4 fanout1011 (.X(net1011),
    .A(net1015));
 sg13g2_buf_4 fanout1012 (.X(net1012),
    .A(net1014));
 sg13g2_buf_2 fanout1013 (.A(net1014),
    .X(net1013));
 sg13g2_buf_4 fanout1014 (.X(net1014),
    .A(net1015));
 sg13g2_buf_2 fanout1015 (.A(net1016),
    .X(net1015));
 sg13g2_buf_4 fanout1016 (.X(net1016),
    .A(rst_n));
 sg13g2_buf_4 fanout1017 (.X(net1017),
    .A(net1019));
 sg13g2_buf_2 fanout1018 (.A(net1019),
    .X(net1018));
 sg13g2_buf_4 fanout1019 (.X(net1019),
    .A(net1022));
 sg13g2_buf_4 fanout1020 (.X(net1020),
    .A(net1022));
 sg13g2_buf_4 fanout1021 (.X(net1021),
    .A(net1022));
 sg13g2_buf_2 fanout1022 (.A(net1060),
    .X(net1022));
 sg13g2_buf_4 fanout1023 (.X(net1023),
    .A(net1027));
 sg13g2_buf_4 fanout1024 (.X(net1024),
    .A(net1027));
 sg13g2_buf_4 fanout1025 (.X(net1025),
    .A(net1027));
 sg13g2_buf_4 fanout1026 (.X(net1026),
    .A(net1027));
 sg13g2_buf_2 fanout1027 (.A(net1060),
    .X(net1027));
 sg13g2_buf_4 fanout1028 (.X(net1028),
    .A(net1029));
 sg13g2_buf_4 fanout1029 (.X(net1029),
    .A(net1032));
 sg13g2_buf_4 fanout1030 (.X(net1030),
    .A(net1032));
 sg13g2_buf_2 fanout1031 (.A(net1032),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(net1039),
    .X(net1032));
 sg13g2_buf_4 fanout1033 (.X(net1033),
    .A(net1039));
 sg13g2_buf_2 fanout1034 (.A(net1039),
    .X(net1034));
 sg13g2_buf_4 fanout1035 (.X(net1035),
    .A(net1038));
 sg13g2_buf_2 fanout1036 (.A(net1038),
    .X(net1036));
 sg13g2_buf_4 fanout1037 (.X(net1037),
    .A(net1038));
 sg13g2_buf_2 fanout1038 (.A(net1039),
    .X(net1038));
 sg13g2_buf_2 fanout1039 (.A(net1060),
    .X(net1039));
 sg13g2_buf_4 fanout1040 (.X(net1040),
    .A(net1042));
 sg13g2_buf_4 fanout1041 (.X(net1041),
    .A(net1042));
 sg13g2_buf_2 fanout1042 (.A(net1050),
    .X(net1042));
 sg13g2_buf_4 fanout1043 (.X(net1043),
    .A(net1050));
 sg13g2_buf_4 fanout1044 (.X(net1044),
    .A(net1050));
 sg13g2_buf_4 fanout1045 (.X(net1045),
    .A(net1049));
 sg13g2_buf_4 fanout1046 (.X(net1046),
    .A(net1049));
 sg13g2_buf_4 fanout1047 (.X(net1047),
    .A(net1049));
 sg13g2_buf_4 fanout1048 (.X(net1048),
    .A(net1049));
 sg13g2_buf_2 fanout1049 (.A(net1050),
    .X(net1049));
 sg13g2_buf_2 fanout1050 (.A(net1060),
    .X(net1050));
 sg13g2_buf_4 fanout1051 (.X(net1051),
    .A(net1054));
 sg13g2_buf_4 fanout1052 (.X(net1052),
    .A(net1054));
 sg13g2_buf_4 fanout1053 (.X(net1053),
    .A(net1054));
 sg13g2_buf_4 fanout1054 (.X(net1054),
    .A(net1060));
 sg13g2_buf_4 fanout1055 (.X(net1055),
    .A(net1059));
 sg13g2_buf_2 fanout1056 (.A(net1059),
    .X(net1056));
 sg13g2_buf_4 fanout1057 (.X(net1057),
    .A(net1058));
 sg13g2_buf_4 fanout1058 (.X(net1058),
    .A(net1059));
 sg13g2_buf_2 fanout1059 (.A(net1060),
    .X(net1059));
 sg13g2_buf_4 fanout1060 (.X(net1060),
    .A(rst_n));
 sg13g2_buf_2 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_tielo tt_um_ddc_arghunter_4 (.L_LO(net4));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_decap_8 FILLER_13_588 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_decap_8 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_637 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_8 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_decap_8 FILLER_13_798 ();
 sg13g2_decap_8 FILLER_13_805 ();
 sg13g2_decap_8 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_833 ();
 sg13g2_decap_8 FILLER_13_840 ();
 sg13g2_decap_8 FILLER_13_847 ();
 sg13g2_decap_8 FILLER_13_854 ();
 sg13g2_fill_1 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_8 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_511 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_574 ();
 sg13g2_decap_8 FILLER_14_581 ();
 sg13g2_decap_8 FILLER_14_588 ();
 sg13g2_decap_8 FILLER_14_595 ();
 sg13g2_decap_8 FILLER_14_602 ();
 sg13g2_decap_8 FILLER_14_609 ();
 sg13g2_decap_8 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_623 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_decap_8 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_decap_8 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_658 ();
 sg13g2_decap_8 FILLER_14_665 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_decap_8 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_decap_8 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_14_840 ();
 sg13g2_decap_8 FILLER_14_847 ();
 sg13g2_decap_8 FILLER_14_854 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_434 ();
 sg13g2_decap_8 FILLER_15_441 ();
 sg13g2_decap_8 FILLER_15_448 ();
 sg13g2_decap_8 FILLER_15_455 ();
 sg13g2_decap_8 FILLER_15_462 ();
 sg13g2_decap_8 FILLER_15_469 ();
 sg13g2_decap_8 FILLER_15_476 ();
 sg13g2_decap_8 FILLER_15_483 ();
 sg13g2_decap_8 FILLER_15_490 ();
 sg13g2_decap_8 FILLER_15_497 ();
 sg13g2_decap_8 FILLER_15_504 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_518 ();
 sg13g2_decap_8 FILLER_15_525 ();
 sg13g2_decap_8 FILLER_15_532 ();
 sg13g2_decap_8 FILLER_15_539 ();
 sg13g2_decap_8 FILLER_15_546 ();
 sg13g2_decap_8 FILLER_15_553 ();
 sg13g2_decap_8 FILLER_15_560 ();
 sg13g2_decap_8 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_574 ();
 sg13g2_decap_8 FILLER_15_581 ();
 sg13g2_decap_8 FILLER_15_588 ();
 sg13g2_decap_8 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_602 ();
 sg13g2_decap_8 FILLER_15_609 ();
 sg13g2_decap_8 FILLER_15_616 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_8 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_644 ();
 sg13g2_decap_8 FILLER_15_651 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_decap_8 FILLER_15_665 ();
 sg13g2_decap_8 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_679 ();
 sg13g2_decap_8 FILLER_15_686 ();
 sg13g2_decap_8 FILLER_15_693 ();
 sg13g2_decap_8 FILLER_15_700 ();
 sg13g2_decap_8 FILLER_15_707 ();
 sg13g2_decap_8 FILLER_15_714 ();
 sg13g2_decap_8 FILLER_15_721 ();
 sg13g2_decap_8 FILLER_15_728 ();
 sg13g2_decap_8 FILLER_15_735 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_decap_8 FILLER_15_749 ();
 sg13g2_decap_8 FILLER_15_756 ();
 sg13g2_decap_8 FILLER_15_763 ();
 sg13g2_decap_8 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_777 ();
 sg13g2_decap_8 FILLER_15_784 ();
 sg13g2_decap_8 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_798 ();
 sg13g2_decap_8 FILLER_15_805 ();
 sg13g2_decap_8 FILLER_15_812 ();
 sg13g2_decap_8 FILLER_15_819 ();
 sg13g2_decap_8 FILLER_15_826 ();
 sg13g2_decap_8 FILLER_15_833 ();
 sg13g2_decap_8 FILLER_15_840 ();
 sg13g2_decap_8 FILLER_15_847 ();
 sg13g2_decap_8 FILLER_15_854 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_8 FILLER_16_455 ();
 sg13g2_decap_8 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_469 ();
 sg13g2_decap_8 FILLER_16_476 ();
 sg13g2_decap_8 FILLER_16_483 ();
 sg13g2_decap_8 FILLER_16_490 ();
 sg13g2_decap_8 FILLER_16_497 ();
 sg13g2_decap_8 FILLER_16_504 ();
 sg13g2_decap_8 FILLER_16_511 ();
 sg13g2_decap_8 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_525 ();
 sg13g2_decap_8 FILLER_16_532 ();
 sg13g2_decap_8 FILLER_16_539 ();
 sg13g2_decap_8 FILLER_16_546 ();
 sg13g2_decap_8 FILLER_16_553 ();
 sg13g2_decap_8 FILLER_16_560 ();
 sg13g2_decap_8 FILLER_16_567 ();
 sg13g2_decap_8 FILLER_16_574 ();
 sg13g2_decap_8 FILLER_16_581 ();
 sg13g2_decap_8 FILLER_16_588 ();
 sg13g2_decap_8 FILLER_16_595 ();
 sg13g2_decap_8 FILLER_16_602 ();
 sg13g2_decap_8 FILLER_16_609 ();
 sg13g2_decap_8 FILLER_16_616 ();
 sg13g2_decap_8 FILLER_16_623 ();
 sg13g2_decap_8 FILLER_16_630 ();
 sg13g2_decap_8 FILLER_16_637 ();
 sg13g2_decap_8 FILLER_16_644 ();
 sg13g2_decap_8 FILLER_16_651 ();
 sg13g2_decap_8 FILLER_16_658 ();
 sg13g2_decap_8 FILLER_16_665 ();
 sg13g2_decap_8 FILLER_16_672 ();
 sg13g2_decap_8 FILLER_16_679 ();
 sg13g2_decap_8 FILLER_16_686 ();
 sg13g2_decap_8 FILLER_16_693 ();
 sg13g2_decap_8 FILLER_16_700 ();
 sg13g2_decap_8 FILLER_16_707 ();
 sg13g2_decap_8 FILLER_16_714 ();
 sg13g2_decap_8 FILLER_16_721 ();
 sg13g2_decap_8 FILLER_16_728 ();
 sg13g2_decap_8 FILLER_16_735 ();
 sg13g2_decap_8 FILLER_16_742 ();
 sg13g2_decap_8 FILLER_16_749 ();
 sg13g2_decap_8 FILLER_16_756 ();
 sg13g2_decap_8 FILLER_16_763 ();
 sg13g2_decap_8 FILLER_16_770 ();
 sg13g2_decap_8 FILLER_16_777 ();
 sg13g2_decap_8 FILLER_16_784 ();
 sg13g2_decap_8 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_798 ();
 sg13g2_decap_8 FILLER_16_805 ();
 sg13g2_decap_8 FILLER_16_812 ();
 sg13g2_decap_8 FILLER_16_819 ();
 sg13g2_decap_8 FILLER_16_826 ();
 sg13g2_decap_8 FILLER_16_833 ();
 sg13g2_decap_8 FILLER_16_840 ();
 sg13g2_decap_8 FILLER_16_847 ();
 sg13g2_decap_8 FILLER_16_854 ();
 sg13g2_fill_1 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_427 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_448 ();
 sg13g2_decap_8 FILLER_17_455 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_497 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_fill_1 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_decap_8 FILLER_18_427 ();
 sg13g2_decap_8 FILLER_18_434 ();
 sg13g2_decap_8 FILLER_18_441 ();
 sg13g2_decap_8 FILLER_18_448 ();
 sg13g2_decap_8 FILLER_18_455 ();
 sg13g2_decap_8 FILLER_18_462 ();
 sg13g2_decap_8 FILLER_18_469 ();
 sg13g2_decap_8 FILLER_18_476 ();
 sg13g2_decap_8 FILLER_18_483 ();
 sg13g2_decap_8 FILLER_18_490 ();
 sg13g2_decap_8 FILLER_18_497 ();
 sg13g2_decap_8 FILLER_18_504 ();
 sg13g2_decap_8 FILLER_18_511 ();
 sg13g2_decap_8 FILLER_18_518 ();
 sg13g2_decap_8 FILLER_18_525 ();
 sg13g2_decap_8 FILLER_18_532 ();
 sg13g2_decap_8 FILLER_18_539 ();
 sg13g2_decap_8 FILLER_18_546 ();
 sg13g2_decap_8 FILLER_18_553 ();
 sg13g2_decap_8 FILLER_18_560 ();
 sg13g2_decap_8 FILLER_18_567 ();
 sg13g2_decap_8 FILLER_18_574 ();
 sg13g2_decap_8 FILLER_18_581 ();
 sg13g2_decap_8 FILLER_18_588 ();
 sg13g2_decap_8 FILLER_18_595 ();
 sg13g2_decap_8 FILLER_18_602 ();
 sg13g2_decap_8 FILLER_18_609 ();
 sg13g2_decap_8 FILLER_18_616 ();
 sg13g2_decap_8 FILLER_18_623 ();
 sg13g2_decap_8 FILLER_18_630 ();
 sg13g2_decap_8 FILLER_18_637 ();
 sg13g2_decap_8 FILLER_18_644 ();
 sg13g2_decap_8 FILLER_18_651 ();
 sg13g2_decap_8 FILLER_18_658 ();
 sg13g2_decap_8 FILLER_18_665 ();
 sg13g2_decap_8 FILLER_18_672 ();
 sg13g2_decap_8 FILLER_18_679 ();
 sg13g2_decap_8 FILLER_18_686 ();
 sg13g2_decap_8 FILLER_18_693 ();
 sg13g2_decap_8 FILLER_18_700 ();
 sg13g2_decap_8 FILLER_18_707 ();
 sg13g2_decap_8 FILLER_18_714 ();
 sg13g2_decap_8 FILLER_18_721 ();
 sg13g2_decap_8 FILLER_18_728 ();
 sg13g2_decap_8 FILLER_18_735 ();
 sg13g2_decap_8 FILLER_18_742 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_decap_8 FILLER_18_756 ();
 sg13g2_decap_8 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_770 ();
 sg13g2_decap_8 FILLER_18_777 ();
 sg13g2_decap_8 FILLER_18_784 ();
 sg13g2_decap_8 FILLER_18_791 ();
 sg13g2_decap_8 FILLER_18_798 ();
 sg13g2_decap_8 FILLER_18_805 ();
 sg13g2_decap_8 FILLER_18_812 ();
 sg13g2_decap_8 FILLER_18_819 ();
 sg13g2_decap_8 FILLER_18_826 ();
 sg13g2_decap_8 FILLER_18_833 ();
 sg13g2_decap_8 FILLER_18_840 ();
 sg13g2_decap_8 FILLER_18_847 ();
 sg13g2_decap_8 FILLER_18_854 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_decap_8 FILLER_19_427 ();
 sg13g2_decap_8 FILLER_19_434 ();
 sg13g2_decap_8 FILLER_19_441 ();
 sg13g2_decap_8 FILLER_19_448 ();
 sg13g2_decap_8 FILLER_19_455 ();
 sg13g2_decap_8 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_490 ();
 sg13g2_decap_8 FILLER_19_497 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_532 ();
 sg13g2_decap_8 FILLER_19_539 ();
 sg13g2_decap_8 FILLER_19_546 ();
 sg13g2_decap_8 FILLER_19_553 ();
 sg13g2_decap_8 FILLER_19_560 ();
 sg13g2_decap_8 FILLER_19_567 ();
 sg13g2_decap_8 FILLER_19_574 ();
 sg13g2_decap_8 FILLER_19_581 ();
 sg13g2_decap_8 FILLER_19_588 ();
 sg13g2_decap_8 FILLER_19_595 ();
 sg13g2_decap_8 FILLER_19_602 ();
 sg13g2_decap_8 FILLER_19_609 ();
 sg13g2_decap_8 FILLER_19_616 ();
 sg13g2_decap_8 FILLER_19_623 ();
 sg13g2_decap_8 FILLER_19_630 ();
 sg13g2_decap_8 FILLER_19_637 ();
 sg13g2_decap_8 FILLER_19_644 ();
 sg13g2_decap_8 FILLER_19_651 ();
 sg13g2_decap_8 FILLER_19_658 ();
 sg13g2_decap_8 FILLER_19_665 ();
 sg13g2_decap_8 FILLER_19_672 ();
 sg13g2_decap_8 FILLER_19_679 ();
 sg13g2_decap_8 FILLER_19_686 ();
 sg13g2_decap_8 FILLER_19_693 ();
 sg13g2_decap_8 FILLER_19_700 ();
 sg13g2_decap_8 FILLER_19_707 ();
 sg13g2_decap_8 FILLER_19_714 ();
 sg13g2_decap_8 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_784 ();
 sg13g2_decap_8 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_798 ();
 sg13g2_decap_8 FILLER_19_805 ();
 sg13g2_decap_8 FILLER_19_812 ();
 sg13g2_decap_8 FILLER_19_819 ();
 sg13g2_decap_8 FILLER_19_826 ();
 sg13g2_decap_8 FILLER_19_833 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_decap_8 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_854 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_decap_8 FILLER_20_427 ();
 sg13g2_decap_8 FILLER_20_434 ();
 sg13g2_decap_8 FILLER_20_441 ();
 sg13g2_decap_8 FILLER_20_448 ();
 sg13g2_decap_8 FILLER_20_455 ();
 sg13g2_decap_8 FILLER_20_462 ();
 sg13g2_decap_8 FILLER_20_469 ();
 sg13g2_decap_8 FILLER_20_476 ();
 sg13g2_decap_8 FILLER_20_483 ();
 sg13g2_decap_8 FILLER_20_490 ();
 sg13g2_decap_8 FILLER_20_497 ();
 sg13g2_decap_8 FILLER_20_504 ();
 sg13g2_decap_8 FILLER_20_511 ();
 sg13g2_decap_8 FILLER_20_518 ();
 sg13g2_decap_8 FILLER_20_525 ();
 sg13g2_decap_8 FILLER_20_532 ();
 sg13g2_decap_8 FILLER_20_539 ();
 sg13g2_decap_8 FILLER_20_546 ();
 sg13g2_decap_8 FILLER_20_553 ();
 sg13g2_decap_8 FILLER_20_560 ();
 sg13g2_decap_8 FILLER_20_567 ();
 sg13g2_decap_8 FILLER_20_574 ();
 sg13g2_decap_8 FILLER_20_581 ();
 sg13g2_decap_8 FILLER_20_588 ();
 sg13g2_decap_8 FILLER_20_595 ();
 sg13g2_decap_8 FILLER_20_602 ();
 sg13g2_decap_8 FILLER_20_609 ();
 sg13g2_decap_8 FILLER_20_616 ();
 sg13g2_decap_8 FILLER_20_623 ();
 sg13g2_decap_8 FILLER_20_630 ();
 sg13g2_decap_8 FILLER_20_637 ();
 sg13g2_decap_8 FILLER_20_644 ();
 sg13g2_decap_8 FILLER_20_651 ();
 sg13g2_decap_8 FILLER_20_658 ();
 sg13g2_decap_8 FILLER_20_665 ();
 sg13g2_decap_8 FILLER_20_672 ();
 sg13g2_decap_8 FILLER_20_679 ();
 sg13g2_decap_8 FILLER_20_686 ();
 sg13g2_decap_8 FILLER_20_693 ();
 sg13g2_decap_8 FILLER_20_700 ();
 sg13g2_decap_8 FILLER_20_707 ();
 sg13g2_decap_8 FILLER_20_714 ();
 sg13g2_decap_8 FILLER_20_721 ();
 sg13g2_decap_8 FILLER_20_728 ();
 sg13g2_decap_8 FILLER_20_735 ();
 sg13g2_decap_8 FILLER_20_742 ();
 sg13g2_decap_8 FILLER_20_749 ();
 sg13g2_decap_8 FILLER_20_756 ();
 sg13g2_decap_8 FILLER_20_763 ();
 sg13g2_decap_8 FILLER_20_770 ();
 sg13g2_decap_8 FILLER_20_777 ();
 sg13g2_decap_8 FILLER_20_784 ();
 sg13g2_decap_8 FILLER_20_791 ();
 sg13g2_decap_8 FILLER_20_798 ();
 sg13g2_decap_8 FILLER_20_805 ();
 sg13g2_decap_8 FILLER_20_812 ();
 sg13g2_decap_8 FILLER_20_819 ();
 sg13g2_decap_8 FILLER_20_826 ();
 sg13g2_decap_8 FILLER_20_833 ();
 sg13g2_decap_8 FILLER_20_840 ();
 sg13g2_decap_8 FILLER_20_847 ();
 sg13g2_decap_8 FILLER_20_854 ();
 sg13g2_fill_1 FILLER_20_861 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_decap_8 FILLER_21_427 ();
 sg13g2_decap_8 FILLER_21_434 ();
 sg13g2_decap_8 FILLER_21_441 ();
 sg13g2_decap_8 FILLER_21_448 ();
 sg13g2_decap_8 FILLER_21_455 ();
 sg13g2_decap_8 FILLER_21_462 ();
 sg13g2_decap_8 FILLER_21_469 ();
 sg13g2_decap_8 FILLER_21_476 ();
 sg13g2_decap_8 FILLER_21_483 ();
 sg13g2_decap_8 FILLER_21_490 ();
 sg13g2_decap_8 FILLER_21_497 ();
 sg13g2_decap_8 FILLER_21_504 ();
 sg13g2_decap_8 FILLER_21_511 ();
 sg13g2_decap_8 FILLER_21_518 ();
 sg13g2_decap_8 FILLER_21_525 ();
 sg13g2_decap_8 FILLER_21_532 ();
 sg13g2_decap_8 FILLER_21_539 ();
 sg13g2_decap_8 FILLER_21_546 ();
 sg13g2_decap_8 FILLER_21_553 ();
 sg13g2_decap_8 FILLER_21_560 ();
 sg13g2_decap_8 FILLER_21_567 ();
 sg13g2_decap_8 FILLER_21_574 ();
 sg13g2_decap_8 FILLER_21_581 ();
 sg13g2_decap_8 FILLER_21_588 ();
 sg13g2_decap_8 FILLER_21_595 ();
 sg13g2_decap_8 FILLER_21_602 ();
 sg13g2_decap_8 FILLER_21_609 ();
 sg13g2_decap_8 FILLER_21_616 ();
 sg13g2_decap_8 FILLER_21_623 ();
 sg13g2_decap_8 FILLER_21_630 ();
 sg13g2_decap_8 FILLER_21_637 ();
 sg13g2_decap_8 FILLER_21_644 ();
 sg13g2_decap_8 FILLER_21_651 ();
 sg13g2_decap_8 FILLER_21_658 ();
 sg13g2_decap_8 FILLER_21_665 ();
 sg13g2_decap_8 FILLER_21_672 ();
 sg13g2_decap_8 FILLER_21_679 ();
 sg13g2_decap_8 FILLER_21_686 ();
 sg13g2_decap_8 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_700 ();
 sg13g2_decap_8 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_714 ();
 sg13g2_decap_8 FILLER_21_721 ();
 sg13g2_decap_8 FILLER_21_728 ();
 sg13g2_decap_8 FILLER_21_735 ();
 sg13g2_decap_8 FILLER_21_742 ();
 sg13g2_decap_8 FILLER_21_749 ();
 sg13g2_decap_8 FILLER_21_756 ();
 sg13g2_decap_8 FILLER_21_763 ();
 sg13g2_decap_8 FILLER_21_770 ();
 sg13g2_decap_8 FILLER_21_777 ();
 sg13g2_decap_8 FILLER_21_784 ();
 sg13g2_decap_8 FILLER_21_791 ();
 sg13g2_decap_8 FILLER_21_798 ();
 sg13g2_decap_8 FILLER_21_805 ();
 sg13g2_decap_8 FILLER_21_812 ();
 sg13g2_decap_8 FILLER_21_819 ();
 sg13g2_decap_8 FILLER_21_826 ();
 sg13g2_decap_8 FILLER_21_833 ();
 sg13g2_decap_8 FILLER_21_840 ();
 sg13g2_decap_8 FILLER_21_847 ();
 sg13g2_decap_8 FILLER_21_854 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_22_406 ();
 sg13g2_decap_8 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_decap_8 FILLER_22_427 ();
 sg13g2_decap_8 FILLER_22_434 ();
 sg13g2_decap_8 FILLER_22_441 ();
 sg13g2_decap_8 FILLER_22_448 ();
 sg13g2_decap_8 FILLER_22_455 ();
 sg13g2_decap_8 FILLER_22_462 ();
 sg13g2_decap_8 FILLER_22_469 ();
 sg13g2_decap_8 FILLER_22_476 ();
 sg13g2_decap_8 FILLER_22_483 ();
 sg13g2_decap_8 FILLER_22_490 ();
 sg13g2_decap_8 FILLER_22_497 ();
 sg13g2_decap_8 FILLER_22_504 ();
 sg13g2_decap_8 FILLER_22_511 ();
 sg13g2_decap_8 FILLER_22_518 ();
 sg13g2_decap_8 FILLER_22_525 ();
 sg13g2_decap_8 FILLER_22_532 ();
 sg13g2_decap_8 FILLER_22_539 ();
 sg13g2_decap_8 FILLER_22_546 ();
 sg13g2_decap_8 FILLER_22_553 ();
 sg13g2_decap_8 FILLER_22_560 ();
 sg13g2_decap_8 FILLER_22_567 ();
 sg13g2_decap_8 FILLER_22_574 ();
 sg13g2_decap_8 FILLER_22_581 ();
 sg13g2_decap_8 FILLER_22_588 ();
 sg13g2_decap_8 FILLER_22_595 ();
 sg13g2_decap_8 FILLER_22_602 ();
 sg13g2_decap_8 FILLER_22_609 ();
 sg13g2_decap_8 FILLER_22_616 ();
 sg13g2_decap_8 FILLER_22_623 ();
 sg13g2_decap_8 FILLER_22_630 ();
 sg13g2_decap_8 FILLER_22_637 ();
 sg13g2_decap_8 FILLER_22_644 ();
 sg13g2_decap_8 FILLER_22_651 ();
 sg13g2_decap_8 FILLER_22_658 ();
 sg13g2_decap_8 FILLER_22_665 ();
 sg13g2_decap_8 FILLER_22_672 ();
 sg13g2_decap_8 FILLER_22_679 ();
 sg13g2_decap_8 FILLER_22_686 ();
 sg13g2_decap_8 FILLER_22_693 ();
 sg13g2_decap_8 FILLER_22_700 ();
 sg13g2_decap_8 FILLER_22_707 ();
 sg13g2_decap_8 FILLER_22_714 ();
 sg13g2_decap_8 FILLER_22_721 ();
 sg13g2_decap_8 FILLER_22_728 ();
 sg13g2_decap_8 FILLER_22_735 ();
 sg13g2_decap_8 FILLER_22_742 ();
 sg13g2_decap_8 FILLER_22_749 ();
 sg13g2_decap_8 FILLER_22_756 ();
 sg13g2_decap_8 FILLER_22_763 ();
 sg13g2_decap_8 FILLER_22_770 ();
 sg13g2_decap_8 FILLER_22_777 ();
 sg13g2_decap_8 FILLER_22_784 ();
 sg13g2_decap_8 FILLER_22_791 ();
 sg13g2_decap_8 FILLER_22_798 ();
 sg13g2_decap_8 FILLER_22_805 ();
 sg13g2_decap_8 FILLER_22_812 ();
 sg13g2_decap_8 FILLER_22_819 ();
 sg13g2_decap_8 FILLER_22_826 ();
 sg13g2_decap_8 FILLER_22_833 ();
 sg13g2_decap_8 FILLER_22_840 ();
 sg13g2_decap_8 FILLER_22_847 ();
 sg13g2_decap_8 FILLER_22_854 ();
 sg13g2_fill_1 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_decap_8 FILLER_23_406 ();
 sg13g2_decap_8 FILLER_23_413 ();
 sg13g2_decap_8 FILLER_23_420 ();
 sg13g2_decap_8 FILLER_23_427 ();
 sg13g2_decap_8 FILLER_23_434 ();
 sg13g2_decap_8 FILLER_23_441 ();
 sg13g2_decap_8 FILLER_23_448 ();
 sg13g2_decap_8 FILLER_23_455 ();
 sg13g2_decap_8 FILLER_23_462 ();
 sg13g2_decap_8 FILLER_23_469 ();
 sg13g2_decap_8 FILLER_23_476 ();
 sg13g2_decap_8 FILLER_23_483 ();
 sg13g2_decap_8 FILLER_23_490 ();
 sg13g2_decap_8 FILLER_23_497 ();
 sg13g2_decap_8 FILLER_23_504 ();
 sg13g2_decap_8 FILLER_23_511 ();
 sg13g2_decap_8 FILLER_23_518 ();
 sg13g2_decap_8 FILLER_23_525 ();
 sg13g2_decap_8 FILLER_23_532 ();
 sg13g2_decap_8 FILLER_23_539 ();
 sg13g2_decap_8 FILLER_23_546 ();
 sg13g2_decap_8 FILLER_23_553 ();
 sg13g2_decap_8 FILLER_23_560 ();
 sg13g2_decap_8 FILLER_23_567 ();
 sg13g2_decap_8 FILLER_23_574 ();
 sg13g2_decap_8 FILLER_23_581 ();
 sg13g2_decap_8 FILLER_23_588 ();
 sg13g2_decap_8 FILLER_23_595 ();
 sg13g2_decap_8 FILLER_23_602 ();
 sg13g2_decap_8 FILLER_23_609 ();
 sg13g2_decap_8 FILLER_23_616 ();
 sg13g2_decap_8 FILLER_23_623 ();
 sg13g2_decap_8 FILLER_23_630 ();
 sg13g2_decap_8 FILLER_23_637 ();
 sg13g2_decap_8 FILLER_23_644 ();
 sg13g2_decap_8 FILLER_23_651 ();
 sg13g2_decap_8 FILLER_23_658 ();
 sg13g2_decap_8 FILLER_23_665 ();
 sg13g2_decap_8 FILLER_23_672 ();
 sg13g2_decap_8 FILLER_23_679 ();
 sg13g2_decap_8 FILLER_23_686 ();
 sg13g2_decap_8 FILLER_23_693 ();
 sg13g2_decap_8 FILLER_23_700 ();
 sg13g2_decap_8 FILLER_23_707 ();
 sg13g2_decap_8 FILLER_23_714 ();
 sg13g2_decap_8 FILLER_23_721 ();
 sg13g2_decap_8 FILLER_23_728 ();
 sg13g2_decap_8 FILLER_23_735 ();
 sg13g2_decap_8 FILLER_23_742 ();
 sg13g2_decap_8 FILLER_23_749 ();
 sg13g2_decap_8 FILLER_23_756 ();
 sg13g2_decap_8 FILLER_23_763 ();
 sg13g2_decap_8 FILLER_23_770 ();
 sg13g2_decap_8 FILLER_23_777 ();
 sg13g2_decap_8 FILLER_23_784 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_798 ();
 sg13g2_decap_8 FILLER_23_805 ();
 sg13g2_decap_8 FILLER_23_812 ();
 sg13g2_decap_8 FILLER_23_819 ();
 sg13g2_decap_8 FILLER_23_826 ();
 sg13g2_decap_8 FILLER_23_833 ();
 sg13g2_decap_8 FILLER_23_840 ();
 sg13g2_decap_8 FILLER_23_847 ();
 sg13g2_decap_8 FILLER_23_854 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_decap_8 FILLER_24_406 ();
 sg13g2_decap_8 FILLER_24_413 ();
 sg13g2_decap_8 FILLER_24_420 ();
 sg13g2_decap_8 FILLER_24_427 ();
 sg13g2_decap_8 FILLER_24_434 ();
 sg13g2_decap_8 FILLER_24_441 ();
 sg13g2_decap_8 FILLER_24_448 ();
 sg13g2_decap_8 FILLER_24_455 ();
 sg13g2_decap_8 FILLER_24_462 ();
 sg13g2_decap_8 FILLER_24_469 ();
 sg13g2_decap_8 FILLER_24_476 ();
 sg13g2_decap_8 FILLER_24_483 ();
 sg13g2_decap_8 FILLER_24_490 ();
 sg13g2_decap_8 FILLER_24_497 ();
 sg13g2_decap_8 FILLER_24_504 ();
 sg13g2_decap_8 FILLER_24_511 ();
 sg13g2_decap_8 FILLER_24_518 ();
 sg13g2_decap_8 FILLER_24_525 ();
 sg13g2_decap_8 FILLER_24_532 ();
 sg13g2_decap_8 FILLER_24_539 ();
 sg13g2_decap_8 FILLER_24_546 ();
 sg13g2_decap_8 FILLER_24_553 ();
 sg13g2_decap_8 FILLER_24_560 ();
 sg13g2_decap_8 FILLER_24_567 ();
 sg13g2_decap_8 FILLER_24_574 ();
 sg13g2_decap_8 FILLER_24_581 ();
 sg13g2_decap_8 FILLER_24_588 ();
 sg13g2_decap_8 FILLER_24_595 ();
 sg13g2_decap_8 FILLER_24_602 ();
 sg13g2_decap_8 FILLER_24_609 ();
 sg13g2_decap_8 FILLER_24_616 ();
 sg13g2_decap_8 FILLER_24_623 ();
 sg13g2_decap_8 FILLER_24_630 ();
 sg13g2_decap_8 FILLER_24_637 ();
 sg13g2_decap_8 FILLER_24_644 ();
 sg13g2_decap_8 FILLER_24_651 ();
 sg13g2_decap_8 FILLER_24_658 ();
 sg13g2_decap_8 FILLER_24_665 ();
 sg13g2_decap_8 FILLER_24_672 ();
 sg13g2_decap_8 FILLER_24_679 ();
 sg13g2_decap_8 FILLER_24_686 ();
 sg13g2_decap_8 FILLER_24_693 ();
 sg13g2_decap_8 FILLER_24_700 ();
 sg13g2_decap_8 FILLER_24_707 ();
 sg13g2_decap_8 FILLER_24_714 ();
 sg13g2_decap_8 FILLER_24_721 ();
 sg13g2_decap_8 FILLER_24_728 ();
 sg13g2_decap_8 FILLER_24_735 ();
 sg13g2_decap_8 FILLER_24_742 ();
 sg13g2_decap_8 FILLER_24_749 ();
 sg13g2_decap_8 FILLER_24_756 ();
 sg13g2_decap_8 FILLER_24_763 ();
 sg13g2_decap_8 FILLER_24_770 ();
 sg13g2_decap_8 FILLER_24_777 ();
 sg13g2_decap_8 FILLER_24_784 ();
 sg13g2_decap_8 FILLER_24_791 ();
 sg13g2_decap_8 FILLER_24_798 ();
 sg13g2_decap_8 FILLER_24_805 ();
 sg13g2_decap_8 FILLER_24_812 ();
 sg13g2_decap_8 FILLER_24_819 ();
 sg13g2_decap_8 FILLER_24_826 ();
 sg13g2_decap_8 FILLER_24_833 ();
 sg13g2_decap_8 FILLER_24_840 ();
 sg13g2_decap_8 FILLER_24_847 ();
 sg13g2_decap_8 FILLER_24_854 ();
 sg13g2_fill_1 FILLER_24_861 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_fill_1 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_125 ();
 sg13g2_decap_8 FILLER_25_132 ();
 sg13g2_decap_8 FILLER_25_139 ();
 sg13g2_decap_8 FILLER_25_146 ();
 sg13g2_decap_8 FILLER_25_153 ();
 sg13g2_decap_8 FILLER_25_160 ();
 sg13g2_decap_8 FILLER_25_167 ();
 sg13g2_decap_8 FILLER_25_174 ();
 sg13g2_decap_8 FILLER_25_181 ();
 sg13g2_decap_8 FILLER_25_188 ();
 sg13g2_decap_8 FILLER_25_195 ();
 sg13g2_decap_8 FILLER_25_202 ();
 sg13g2_decap_8 FILLER_25_209 ();
 sg13g2_decap_8 FILLER_25_216 ();
 sg13g2_decap_8 FILLER_25_223 ();
 sg13g2_decap_8 FILLER_25_230 ();
 sg13g2_decap_8 FILLER_25_237 ();
 sg13g2_decap_8 FILLER_25_244 ();
 sg13g2_decap_8 FILLER_25_251 ();
 sg13g2_decap_8 FILLER_25_258 ();
 sg13g2_decap_8 FILLER_25_265 ();
 sg13g2_decap_8 FILLER_25_272 ();
 sg13g2_decap_8 FILLER_25_279 ();
 sg13g2_decap_8 FILLER_25_286 ();
 sg13g2_decap_8 FILLER_25_293 ();
 sg13g2_decap_8 FILLER_25_300 ();
 sg13g2_decap_8 FILLER_25_307 ();
 sg13g2_decap_8 FILLER_25_314 ();
 sg13g2_decap_8 FILLER_25_321 ();
 sg13g2_decap_8 FILLER_25_328 ();
 sg13g2_decap_8 FILLER_25_335 ();
 sg13g2_decap_8 FILLER_25_342 ();
 sg13g2_decap_8 FILLER_25_349 ();
 sg13g2_decap_8 FILLER_25_356 ();
 sg13g2_decap_8 FILLER_25_363 ();
 sg13g2_decap_8 FILLER_25_370 ();
 sg13g2_decap_8 FILLER_25_377 ();
 sg13g2_decap_8 FILLER_25_384 ();
 sg13g2_decap_8 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_8 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_25_412 ();
 sg13g2_decap_8 FILLER_25_419 ();
 sg13g2_decap_8 FILLER_25_426 ();
 sg13g2_decap_8 FILLER_25_433 ();
 sg13g2_decap_8 FILLER_25_440 ();
 sg13g2_decap_8 FILLER_25_447 ();
 sg13g2_decap_8 FILLER_25_454 ();
 sg13g2_decap_8 FILLER_25_461 ();
 sg13g2_decap_8 FILLER_25_468 ();
 sg13g2_decap_8 FILLER_25_475 ();
 sg13g2_decap_8 FILLER_25_482 ();
 sg13g2_decap_8 FILLER_25_489 ();
 sg13g2_decap_8 FILLER_25_496 ();
 sg13g2_decap_8 FILLER_25_503 ();
 sg13g2_decap_8 FILLER_25_510 ();
 sg13g2_decap_8 FILLER_25_517 ();
 sg13g2_decap_8 FILLER_25_524 ();
 sg13g2_decap_8 FILLER_25_531 ();
 sg13g2_decap_8 FILLER_25_538 ();
 sg13g2_decap_8 FILLER_25_545 ();
 sg13g2_decap_8 FILLER_25_552 ();
 sg13g2_decap_8 FILLER_25_559 ();
 sg13g2_decap_8 FILLER_25_566 ();
 sg13g2_decap_8 FILLER_25_573 ();
 sg13g2_decap_8 FILLER_25_580 ();
 sg13g2_decap_8 FILLER_25_587 ();
 sg13g2_decap_8 FILLER_25_594 ();
 sg13g2_decap_8 FILLER_25_601 ();
 sg13g2_decap_8 FILLER_25_608 ();
 sg13g2_decap_8 FILLER_25_615 ();
 sg13g2_decap_8 FILLER_25_622 ();
 sg13g2_decap_8 FILLER_25_629 ();
 sg13g2_decap_8 FILLER_25_636 ();
 sg13g2_decap_8 FILLER_25_643 ();
 sg13g2_decap_8 FILLER_25_650 ();
 sg13g2_decap_8 FILLER_25_657 ();
 sg13g2_decap_8 FILLER_25_664 ();
 sg13g2_decap_8 FILLER_25_671 ();
 sg13g2_decap_8 FILLER_25_678 ();
 sg13g2_decap_8 FILLER_25_685 ();
 sg13g2_decap_8 FILLER_25_692 ();
 sg13g2_decap_8 FILLER_25_699 ();
 sg13g2_decap_8 FILLER_25_706 ();
 sg13g2_decap_8 FILLER_25_713 ();
 sg13g2_decap_8 FILLER_25_720 ();
 sg13g2_decap_8 FILLER_25_727 ();
 sg13g2_decap_8 FILLER_25_734 ();
 sg13g2_decap_8 FILLER_25_741 ();
 sg13g2_decap_8 FILLER_25_748 ();
 sg13g2_decap_8 FILLER_25_755 ();
 sg13g2_decap_8 FILLER_25_762 ();
 sg13g2_decap_8 FILLER_25_769 ();
 sg13g2_decap_8 FILLER_25_776 ();
 sg13g2_decap_8 FILLER_25_783 ();
 sg13g2_decap_8 FILLER_25_790 ();
 sg13g2_decap_8 FILLER_25_797 ();
 sg13g2_decap_8 FILLER_25_804 ();
 sg13g2_decap_8 FILLER_25_811 ();
 sg13g2_decap_8 FILLER_25_818 ();
 sg13g2_decap_8 FILLER_25_825 ();
 sg13g2_decap_8 FILLER_25_832 ();
 sg13g2_decap_8 FILLER_25_839 ();
 sg13g2_decap_8 FILLER_25_846 ();
 sg13g2_decap_8 FILLER_25_853 ();
 sg13g2_fill_2 FILLER_25_860 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_fill_2 FILLER_26_28 ();
 sg13g2_fill_1 FILLER_26_30 ();
 sg13g2_decap_8 FILLER_26_57 ();
 sg13g2_decap_8 FILLER_26_90 ();
 sg13g2_fill_2 FILLER_26_97 ();
 sg13g2_decap_8 FILLER_26_131 ();
 sg13g2_decap_8 FILLER_26_138 ();
 sg13g2_fill_2 FILLER_26_145 ();
 sg13g2_fill_1 FILLER_26_147 ();
 sg13g2_fill_2 FILLER_26_174 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_218 ();
 sg13g2_decap_8 FILLER_26_225 ();
 sg13g2_decap_4 FILLER_26_232 ();
 sg13g2_decap_8 FILLER_26_239 ();
 sg13g2_decap_8 FILLER_26_246 ();
 sg13g2_decap_8 FILLER_26_253 ();
 sg13g2_decap_8 FILLER_26_260 ();
 sg13g2_decap_8 FILLER_26_267 ();
 sg13g2_decap_8 FILLER_26_274 ();
 sg13g2_decap_8 FILLER_26_281 ();
 sg13g2_decap_8 FILLER_26_288 ();
 sg13g2_decap_8 FILLER_26_295 ();
 sg13g2_decap_8 FILLER_26_302 ();
 sg13g2_decap_8 FILLER_26_309 ();
 sg13g2_decap_8 FILLER_26_316 ();
 sg13g2_decap_8 FILLER_26_323 ();
 sg13g2_decap_8 FILLER_26_330 ();
 sg13g2_decap_8 FILLER_26_337 ();
 sg13g2_decap_8 FILLER_26_344 ();
 sg13g2_decap_8 FILLER_26_351 ();
 sg13g2_decap_8 FILLER_26_358 ();
 sg13g2_decap_8 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_26_372 ();
 sg13g2_decap_8 FILLER_26_379 ();
 sg13g2_decap_8 FILLER_26_386 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_decap_8 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_26_414 ();
 sg13g2_decap_8 FILLER_26_421 ();
 sg13g2_decap_8 FILLER_26_428 ();
 sg13g2_decap_8 FILLER_26_435 ();
 sg13g2_decap_8 FILLER_26_442 ();
 sg13g2_decap_8 FILLER_26_449 ();
 sg13g2_decap_8 FILLER_26_456 ();
 sg13g2_decap_8 FILLER_26_463 ();
 sg13g2_decap_8 FILLER_26_470 ();
 sg13g2_decap_8 FILLER_26_477 ();
 sg13g2_decap_8 FILLER_26_484 ();
 sg13g2_decap_8 FILLER_26_491 ();
 sg13g2_decap_8 FILLER_26_498 ();
 sg13g2_decap_8 FILLER_26_505 ();
 sg13g2_decap_8 FILLER_26_512 ();
 sg13g2_decap_8 FILLER_26_519 ();
 sg13g2_decap_8 FILLER_26_526 ();
 sg13g2_decap_8 FILLER_26_533 ();
 sg13g2_decap_8 FILLER_26_540 ();
 sg13g2_decap_8 FILLER_26_547 ();
 sg13g2_decap_8 FILLER_26_554 ();
 sg13g2_decap_8 FILLER_26_561 ();
 sg13g2_decap_8 FILLER_26_568 ();
 sg13g2_decap_8 FILLER_26_575 ();
 sg13g2_decap_8 FILLER_26_582 ();
 sg13g2_decap_8 FILLER_26_589 ();
 sg13g2_decap_8 FILLER_26_596 ();
 sg13g2_decap_8 FILLER_26_603 ();
 sg13g2_decap_8 FILLER_26_610 ();
 sg13g2_decap_8 FILLER_26_617 ();
 sg13g2_decap_8 FILLER_26_624 ();
 sg13g2_decap_8 FILLER_26_631 ();
 sg13g2_decap_8 FILLER_26_638 ();
 sg13g2_decap_8 FILLER_26_645 ();
 sg13g2_decap_8 FILLER_26_652 ();
 sg13g2_decap_8 FILLER_26_659 ();
 sg13g2_decap_8 FILLER_26_666 ();
 sg13g2_decap_8 FILLER_26_673 ();
 sg13g2_decap_8 FILLER_26_680 ();
 sg13g2_decap_8 FILLER_26_687 ();
 sg13g2_decap_8 FILLER_26_694 ();
 sg13g2_decap_8 FILLER_26_701 ();
 sg13g2_decap_8 FILLER_26_708 ();
 sg13g2_decap_8 FILLER_26_715 ();
 sg13g2_decap_8 FILLER_26_722 ();
 sg13g2_decap_8 FILLER_26_729 ();
 sg13g2_decap_8 FILLER_26_736 ();
 sg13g2_decap_8 FILLER_26_743 ();
 sg13g2_decap_8 FILLER_26_750 ();
 sg13g2_decap_8 FILLER_26_757 ();
 sg13g2_decap_8 FILLER_26_764 ();
 sg13g2_decap_8 FILLER_26_771 ();
 sg13g2_decap_8 FILLER_26_778 ();
 sg13g2_decap_8 FILLER_26_785 ();
 sg13g2_decap_8 FILLER_26_792 ();
 sg13g2_decap_8 FILLER_26_799 ();
 sg13g2_decap_8 FILLER_26_806 ();
 sg13g2_decap_8 FILLER_26_813 ();
 sg13g2_decap_8 FILLER_26_820 ();
 sg13g2_decap_8 FILLER_26_827 ();
 sg13g2_decap_8 FILLER_26_834 ();
 sg13g2_decap_8 FILLER_26_841 ();
 sg13g2_decap_8 FILLER_26_848 ();
 sg13g2_decap_8 FILLER_26_855 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_4 FILLER_27_14 ();
 sg13g2_fill_1 FILLER_27_18 ();
 sg13g2_decap_4 FILLER_27_57 ();
 sg13g2_fill_2 FILLER_27_61 ();
 sg13g2_fill_2 FILLER_27_71 ();
 sg13g2_fill_2 FILLER_27_103 ();
 sg13g2_decap_4 FILLER_27_132 ();
 sg13g2_fill_2 FILLER_27_136 ();
 sg13g2_decap_4 FILLER_27_148 ();
 sg13g2_fill_2 FILLER_27_152 ();
 sg13g2_fill_1 FILLER_27_157 ();
 sg13g2_fill_2 FILLER_27_215 ();
 sg13g2_decap_8 FILLER_27_261 ();
 sg13g2_decap_8 FILLER_27_268 ();
 sg13g2_decap_8 FILLER_27_275 ();
 sg13g2_decap_8 FILLER_27_282 ();
 sg13g2_decap_8 FILLER_27_289 ();
 sg13g2_decap_8 FILLER_27_296 ();
 sg13g2_decap_8 FILLER_27_303 ();
 sg13g2_decap_8 FILLER_27_310 ();
 sg13g2_decap_8 FILLER_27_317 ();
 sg13g2_decap_8 FILLER_27_324 ();
 sg13g2_decap_8 FILLER_27_331 ();
 sg13g2_decap_8 FILLER_27_338 ();
 sg13g2_decap_8 FILLER_27_345 ();
 sg13g2_decap_8 FILLER_27_352 ();
 sg13g2_decap_8 FILLER_27_359 ();
 sg13g2_decap_8 FILLER_27_366 ();
 sg13g2_decap_8 FILLER_27_373 ();
 sg13g2_decap_8 FILLER_27_380 ();
 sg13g2_decap_8 FILLER_27_387 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_decap_8 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_27_415 ();
 sg13g2_decap_8 FILLER_27_422 ();
 sg13g2_decap_8 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_27_436 ();
 sg13g2_decap_8 FILLER_27_443 ();
 sg13g2_decap_8 FILLER_27_450 ();
 sg13g2_decap_8 FILLER_27_457 ();
 sg13g2_decap_8 FILLER_27_464 ();
 sg13g2_decap_8 FILLER_27_471 ();
 sg13g2_decap_8 FILLER_27_478 ();
 sg13g2_decap_8 FILLER_27_485 ();
 sg13g2_decap_8 FILLER_27_492 ();
 sg13g2_decap_8 FILLER_27_499 ();
 sg13g2_decap_8 FILLER_27_506 ();
 sg13g2_decap_8 FILLER_27_513 ();
 sg13g2_decap_8 FILLER_27_520 ();
 sg13g2_decap_8 FILLER_27_527 ();
 sg13g2_decap_8 FILLER_27_534 ();
 sg13g2_decap_8 FILLER_27_541 ();
 sg13g2_decap_8 FILLER_27_548 ();
 sg13g2_decap_8 FILLER_27_555 ();
 sg13g2_decap_8 FILLER_27_562 ();
 sg13g2_decap_8 FILLER_27_569 ();
 sg13g2_decap_8 FILLER_27_576 ();
 sg13g2_decap_8 FILLER_27_583 ();
 sg13g2_decap_8 FILLER_27_590 ();
 sg13g2_decap_8 FILLER_27_597 ();
 sg13g2_decap_8 FILLER_27_604 ();
 sg13g2_decap_8 FILLER_27_611 ();
 sg13g2_decap_8 FILLER_27_618 ();
 sg13g2_decap_8 FILLER_27_625 ();
 sg13g2_decap_8 FILLER_27_632 ();
 sg13g2_decap_8 FILLER_27_639 ();
 sg13g2_decap_8 FILLER_27_646 ();
 sg13g2_decap_8 FILLER_27_653 ();
 sg13g2_decap_8 FILLER_27_660 ();
 sg13g2_decap_8 FILLER_27_667 ();
 sg13g2_decap_8 FILLER_27_674 ();
 sg13g2_decap_8 FILLER_27_681 ();
 sg13g2_decap_8 FILLER_27_688 ();
 sg13g2_decap_8 FILLER_27_695 ();
 sg13g2_decap_8 FILLER_27_702 ();
 sg13g2_decap_8 FILLER_27_709 ();
 sg13g2_decap_8 FILLER_27_716 ();
 sg13g2_decap_8 FILLER_27_723 ();
 sg13g2_decap_8 FILLER_27_730 ();
 sg13g2_decap_8 FILLER_27_737 ();
 sg13g2_decap_8 FILLER_27_744 ();
 sg13g2_decap_8 FILLER_27_751 ();
 sg13g2_decap_8 FILLER_27_758 ();
 sg13g2_decap_8 FILLER_27_765 ();
 sg13g2_decap_8 FILLER_27_772 ();
 sg13g2_decap_8 FILLER_27_779 ();
 sg13g2_decap_8 FILLER_27_786 ();
 sg13g2_decap_8 FILLER_27_793 ();
 sg13g2_decap_8 FILLER_27_800 ();
 sg13g2_decap_8 FILLER_27_807 ();
 sg13g2_decap_8 FILLER_27_814 ();
 sg13g2_decap_8 FILLER_27_821 ();
 sg13g2_decap_8 FILLER_27_828 ();
 sg13g2_decap_8 FILLER_27_835 ();
 sg13g2_decap_8 FILLER_27_842 ();
 sg13g2_decap_8 FILLER_27_849 ();
 sg13g2_decap_4 FILLER_27_856 ();
 sg13g2_fill_2 FILLER_27_860 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_4 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_33 ();
 sg13g2_fill_2 FILLER_28_40 ();
 sg13g2_decap_8 FILLER_28_54 ();
 sg13g2_decap_8 FILLER_28_61 ();
 sg13g2_decap_4 FILLER_28_68 ();
 sg13g2_fill_2 FILLER_28_72 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_fill_1 FILLER_28_91 ();
 sg13g2_decap_4 FILLER_28_96 ();
 sg13g2_decap_8 FILLER_28_103 ();
 sg13g2_fill_2 FILLER_28_110 ();
 sg13g2_fill_1 FILLER_28_112 ();
 sg13g2_decap_4 FILLER_28_122 ();
 sg13g2_fill_2 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_4 FILLER_28_161 ();
 sg13g2_fill_2 FILLER_28_165 ();
 sg13g2_decap_8 FILLER_28_170 ();
 sg13g2_decap_8 FILLER_28_177 ();
 sg13g2_decap_8 FILLER_28_184 ();
 sg13g2_decap_8 FILLER_28_191 ();
 sg13g2_fill_2 FILLER_28_198 ();
 sg13g2_fill_2 FILLER_28_215 ();
 sg13g2_fill_1 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_264 ();
 sg13g2_decap_8 FILLER_28_271 ();
 sg13g2_decap_8 FILLER_28_278 ();
 sg13g2_decap_8 FILLER_28_285 ();
 sg13g2_decap_8 FILLER_28_292 ();
 sg13g2_decap_8 FILLER_28_299 ();
 sg13g2_decap_8 FILLER_28_306 ();
 sg13g2_decap_8 FILLER_28_313 ();
 sg13g2_decap_8 FILLER_28_320 ();
 sg13g2_decap_8 FILLER_28_327 ();
 sg13g2_decap_8 FILLER_28_334 ();
 sg13g2_decap_8 FILLER_28_341 ();
 sg13g2_decap_8 FILLER_28_348 ();
 sg13g2_decap_8 FILLER_28_355 ();
 sg13g2_decap_8 FILLER_28_362 ();
 sg13g2_decap_8 FILLER_28_369 ();
 sg13g2_decap_8 FILLER_28_376 ();
 sg13g2_decap_8 FILLER_28_383 ();
 sg13g2_decap_8 FILLER_28_390 ();
 sg13g2_decap_8 FILLER_28_397 ();
 sg13g2_decap_8 FILLER_28_404 ();
 sg13g2_decap_8 FILLER_28_411 ();
 sg13g2_decap_8 FILLER_28_418 ();
 sg13g2_decap_8 FILLER_28_425 ();
 sg13g2_decap_8 FILLER_28_432 ();
 sg13g2_decap_8 FILLER_28_439 ();
 sg13g2_decap_8 FILLER_28_446 ();
 sg13g2_decap_8 FILLER_28_453 ();
 sg13g2_decap_8 FILLER_28_460 ();
 sg13g2_decap_8 FILLER_28_467 ();
 sg13g2_decap_8 FILLER_28_474 ();
 sg13g2_decap_8 FILLER_28_481 ();
 sg13g2_decap_8 FILLER_28_488 ();
 sg13g2_decap_4 FILLER_28_495 ();
 sg13g2_decap_8 FILLER_28_502 ();
 sg13g2_decap_8 FILLER_28_509 ();
 sg13g2_decap_8 FILLER_28_516 ();
 sg13g2_decap_8 FILLER_28_523 ();
 sg13g2_decap_8 FILLER_28_530 ();
 sg13g2_decap_8 FILLER_28_537 ();
 sg13g2_decap_4 FILLER_28_544 ();
 sg13g2_decap_8 FILLER_28_558 ();
 sg13g2_decap_8 FILLER_28_565 ();
 sg13g2_decap_8 FILLER_28_572 ();
 sg13g2_fill_1 FILLER_28_579 ();
 sg13g2_fill_2 FILLER_28_588 ();
 sg13g2_fill_1 FILLER_28_590 ();
 sg13g2_decap_8 FILLER_28_601 ();
 sg13g2_fill_1 FILLER_28_608 ();
 sg13g2_decap_8 FILLER_28_612 ();
 sg13g2_decap_8 FILLER_28_619 ();
 sg13g2_decap_4 FILLER_28_626 ();
 sg13g2_fill_1 FILLER_28_630 ();
 sg13g2_decap_8 FILLER_28_654 ();
 sg13g2_decap_8 FILLER_28_661 ();
 sg13g2_decap_8 FILLER_28_668 ();
 sg13g2_decap_8 FILLER_28_675 ();
 sg13g2_decap_8 FILLER_28_682 ();
 sg13g2_decap_8 FILLER_28_689 ();
 sg13g2_decap_8 FILLER_28_696 ();
 sg13g2_decap_8 FILLER_28_703 ();
 sg13g2_decap_8 FILLER_28_710 ();
 sg13g2_decap_8 FILLER_28_717 ();
 sg13g2_decap_8 FILLER_28_724 ();
 sg13g2_decap_8 FILLER_28_731 ();
 sg13g2_decap_8 FILLER_28_738 ();
 sg13g2_decap_8 FILLER_28_745 ();
 sg13g2_decap_8 FILLER_28_752 ();
 sg13g2_decap_8 FILLER_28_759 ();
 sg13g2_decap_8 FILLER_28_766 ();
 sg13g2_decap_8 FILLER_28_773 ();
 sg13g2_decap_8 FILLER_28_780 ();
 sg13g2_decap_8 FILLER_28_787 ();
 sg13g2_decap_8 FILLER_28_794 ();
 sg13g2_decap_8 FILLER_28_801 ();
 sg13g2_decap_8 FILLER_28_808 ();
 sg13g2_decap_8 FILLER_28_815 ();
 sg13g2_decap_8 FILLER_28_822 ();
 sg13g2_decap_8 FILLER_28_829 ();
 sg13g2_decap_8 FILLER_28_836 ();
 sg13g2_decap_8 FILLER_28_843 ();
 sg13g2_decap_8 FILLER_28_850 ();
 sg13g2_decap_4 FILLER_28_857 ();
 sg13g2_fill_1 FILLER_28_861 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_11 ();
 sg13g2_fill_2 FILLER_29_34 ();
 sg13g2_decap_8 FILLER_29_83 ();
 sg13g2_decap_4 FILLER_29_90 ();
 sg13g2_fill_1 FILLER_29_141 ();
 sg13g2_fill_1 FILLER_29_147 ();
 sg13g2_decap_4 FILLER_29_187 ();
 sg13g2_fill_1 FILLER_29_191 ();
 sg13g2_decap_4 FILLER_29_200 ();
 sg13g2_fill_2 FILLER_29_208 ();
 sg13g2_decap_8 FILLER_29_228 ();
 sg13g2_decap_8 FILLER_29_241 ();
 sg13g2_decap_8 FILLER_29_248 ();
 sg13g2_fill_1 FILLER_29_255 ();
 sg13g2_decap_8 FILLER_29_271 ();
 sg13g2_decap_4 FILLER_29_278 ();
 sg13g2_fill_1 FILLER_29_282 ();
 sg13g2_fill_2 FILLER_29_291 ();
 sg13g2_fill_1 FILLER_29_293 ();
 sg13g2_decap_8 FILLER_29_322 ();
 sg13g2_decap_8 FILLER_29_329 ();
 sg13g2_decap_8 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_343 ();
 sg13g2_decap_8 FILLER_29_350 ();
 sg13g2_decap_8 FILLER_29_357 ();
 sg13g2_decap_4 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_decap_8 FILLER_29_406 ();
 sg13g2_decap_8 FILLER_29_413 ();
 sg13g2_decap_8 FILLER_29_420 ();
 sg13g2_decap_8 FILLER_29_427 ();
 sg13g2_decap_8 FILLER_29_434 ();
 sg13g2_decap_8 FILLER_29_441 ();
 sg13g2_decap_8 FILLER_29_448 ();
 sg13g2_decap_8 FILLER_29_455 ();
 sg13g2_decap_8 FILLER_29_462 ();
 sg13g2_decap_8 FILLER_29_469 ();
 sg13g2_decap_8 FILLER_29_476 ();
 sg13g2_decap_8 FILLER_29_483 ();
 sg13g2_fill_2 FILLER_29_490 ();
 sg13g2_fill_2 FILLER_29_518 ();
 sg13g2_fill_1 FILLER_29_520 ();
 sg13g2_decap_8 FILLER_29_524 ();
 sg13g2_decap_8 FILLER_29_531 ();
 sg13g2_decap_4 FILLER_29_538 ();
 sg13g2_fill_2 FILLER_29_542 ();
 sg13g2_decap_4 FILLER_29_573 ();
 sg13g2_fill_1 FILLER_29_587 ();
 sg13g2_decap_8 FILLER_29_666 ();
 sg13g2_decap_8 FILLER_29_673 ();
 sg13g2_decap_8 FILLER_29_680 ();
 sg13g2_decap_8 FILLER_29_687 ();
 sg13g2_decap_8 FILLER_29_694 ();
 sg13g2_decap_8 FILLER_29_701 ();
 sg13g2_decap_8 FILLER_29_708 ();
 sg13g2_decap_8 FILLER_29_715 ();
 sg13g2_decap_8 FILLER_29_722 ();
 sg13g2_fill_1 FILLER_29_729 ();
 sg13g2_decap_8 FILLER_29_738 ();
 sg13g2_decap_8 FILLER_29_745 ();
 sg13g2_fill_2 FILLER_29_752 ();
 sg13g2_decap_8 FILLER_29_762 ();
 sg13g2_decap_8 FILLER_29_769 ();
 sg13g2_decap_8 FILLER_29_776 ();
 sg13g2_decap_8 FILLER_29_783 ();
 sg13g2_decap_8 FILLER_29_790 ();
 sg13g2_decap_8 FILLER_29_797 ();
 sg13g2_decap_8 FILLER_29_804 ();
 sg13g2_decap_8 FILLER_29_811 ();
 sg13g2_decap_8 FILLER_29_818 ();
 sg13g2_decap_8 FILLER_29_825 ();
 sg13g2_decap_8 FILLER_29_832 ();
 sg13g2_decap_8 FILLER_29_839 ();
 sg13g2_decap_8 FILLER_29_846 ();
 sg13g2_decap_8 FILLER_29_853 ();
 sg13g2_fill_2 FILLER_29_860 ();
 sg13g2_decap_8 FILLER_30_34 ();
 sg13g2_decap_4 FILLER_30_62 ();
 sg13g2_fill_2 FILLER_30_66 ();
 sg13g2_fill_2 FILLER_30_111 ();
 sg13g2_fill_1 FILLER_30_113 ();
 sg13g2_decap_8 FILLER_30_117 ();
 sg13g2_decap_8 FILLER_30_129 ();
 sg13g2_decap_8 FILLER_30_136 ();
 sg13g2_fill_2 FILLER_30_143 ();
 sg13g2_fill_1 FILLER_30_145 ();
 sg13g2_decap_4 FILLER_30_156 ();
 sg13g2_fill_1 FILLER_30_160 ();
 sg13g2_fill_2 FILLER_30_217 ();
 sg13g2_fill_2 FILLER_30_320 ();
 sg13g2_fill_1 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_decap_8 FILLER_30_442 ();
 sg13g2_decap_8 FILLER_30_449 ();
 sg13g2_decap_8 FILLER_30_456 ();
 sg13g2_decap_8 FILLER_30_463 ();
 sg13g2_decap_8 FILLER_30_470 ();
 sg13g2_decap_4 FILLER_30_477 ();
 sg13g2_fill_2 FILLER_30_501 ();
 sg13g2_fill_2 FILLER_30_552 ();
 sg13g2_fill_1 FILLER_30_554 ();
 sg13g2_decap_8 FILLER_30_565 ();
 sg13g2_decap_4 FILLER_30_572 ();
 sg13g2_fill_2 FILLER_30_576 ();
 sg13g2_decap_8 FILLER_30_583 ();
 sg13g2_fill_1 FILLER_30_590 ();
 sg13g2_decap_8 FILLER_30_601 ();
 sg13g2_decap_4 FILLER_30_608 ();
 sg13g2_fill_2 FILLER_30_612 ();
 sg13g2_decap_8 FILLER_30_617 ();
 sg13g2_decap_4 FILLER_30_624 ();
 sg13g2_fill_1 FILLER_30_638 ();
 sg13g2_fill_1 FILLER_30_644 ();
 sg13g2_decap_8 FILLER_30_689 ();
 sg13g2_fill_1 FILLER_30_696 ();
 sg13g2_fill_2 FILLER_30_731 ();
 sg13g2_fill_1 FILLER_30_733 ();
 sg13g2_decap_8 FILLER_30_786 ();
 sg13g2_decap_8 FILLER_30_793 ();
 sg13g2_decap_8 FILLER_30_800 ();
 sg13g2_decap_8 FILLER_30_807 ();
 sg13g2_decap_8 FILLER_30_814 ();
 sg13g2_decap_8 FILLER_30_821 ();
 sg13g2_decap_8 FILLER_30_828 ();
 sg13g2_decap_8 FILLER_30_835 ();
 sg13g2_decap_8 FILLER_30_842 ();
 sg13g2_decap_8 FILLER_30_849 ();
 sg13g2_decap_4 FILLER_30_856 ();
 sg13g2_fill_2 FILLER_30_860 ();
 sg13g2_decap_4 FILLER_31_39 ();
 sg13g2_fill_2 FILLER_31_43 ();
 sg13g2_decap_8 FILLER_31_71 ();
 sg13g2_decap_8 FILLER_31_78 ();
 sg13g2_decap_8 FILLER_31_85 ();
 sg13g2_fill_2 FILLER_31_101 ();
 sg13g2_fill_1 FILLER_31_103 ();
 sg13g2_fill_2 FILLER_31_143 ();
 sg13g2_fill_1 FILLER_31_145 ();
 sg13g2_fill_2 FILLER_31_166 ();
 sg13g2_fill_1 FILLER_31_168 ();
 sg13g2_decap_4 FILLER_31_201 ();
 sg13g2_fill_2 FILLER_31_205 ();
 sg13g2_decap_4 FILLER_31_211 ();
 sg13g2_fill_1 FILLER_31_215 ();
 sg13g2_decap_8 FILLER_31_239 ();
 sg13g2_fill_1 FILLER_31_246 ();
 sg13g2_decap_4 FILLER_31_273 ();
 sg13g2_fill_2 FILLER_31_277 ();
 sg13g2_decap_4 FILLER_31_288 ();
 sg13g2_decap_8 FILLER_31_295 ();
 sg13g2_decap_8 FILLER_31_302 ();
 sg13g2_decap_4 FILLER_31_309 ();
 sg13g2_fill_2 FILLER_31_313 ();
 sg13g2_decap_4 FILLER_31_325 ();
 sg13g2_fill_2 FILLER_31_329 ();
 sg13g2_decap_8 FILLER_31_357 ();
 sg13g2_decap_4 FILLER_31_364 ();
 sg13g2_fill_2 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_416 ();
 sg13g2_fill_2 FILLER_31_423 ();
 sg13g2_fill_2 FILLER_31_435 ();
 sg13g2_fill_1 FILLER_31_437 ();
 sg13g2_decap_4 FILLER_31_464 ();
 sg13g2_fill_2 FILLER_31_468 ();
 sg13g2_fill_1 FILLER_31_490 ();
 sg13g2_fill_2 FILLER_31_499 ();
 sg13g2_fill_1 FILLER_31_501 ();
 sg13g2_fill_1 FILLER_31_510 ();
 sg13g2_decap_8 FILLER_31_521 ();
 sg13g2_decap_8 FILLER_31_528 ();
 sg13g2_decap_4 FILLER_31_535 ();
 sg13g2_fill_1 FILLER_31_576 ();
 sg13g2_fill_1 FILLER_31_585 ();
 sg13g2_fill_1 FILLER_31_661 ();
 sg13g2_decap_8 FILLER_31_665 ();
 sg13g2_decap_8 FILLER_31_672 ();
 sg13g2_fill_2 FILLER_31_679 ();
 sg13g2_decap_8 FILLER_31_684 ();
 sg13g2_fill_2 FILLER_31_691 ();
 sg13g2_decap_8 FILLER_31_710 ();
 sg13g2_decap_8 FILLER_31_717 ();
 sg13g2_decap_4 FILLER_31_724 ();
 sg13g2_fill_1 FILLER_31_728 ();
 sg13g2_decap_8 FILLER_31_745 ();
 sg13g2_decap_8 FILLER_31_752 ();
 sg13g2_fill_2 FILLER_31_759 ();
 sg13g2_fill_1 FILLER_31_761 ();
 sg13g2_decap_8 FILLER_31_779 ();
 sg13g2_decap_8 FILLER_31_786 ();
 sg13g2_decap_8 FILLER_31_793 ();
 sg13g2_decap_8 FILLER_31_800 ();
 sg13g2_decap_8 FILLER_31_807 ();
 sg13g2_decap_8 FILLER_31_814 ();
 sg13g2_decap_8 FILLER_31_821 ();
 sg13g2_decap_8 FILLER_31_828 ();
 sg13g2_decap_8 FILLER_31_835 ();
 sg13g2_decap_8 FILLER_31_842 ();
 sg13g2_decap_8 FILLER_31_849 ();
 sg13g2_decap_4 FILLER_31_856 ();
 sg13g2_fill_2 FILLER_31_860 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_4 FILLER_32_38 ();
 sg13g2_fill_1 FILLER_32_42 ();
 sg13g2_decap_4 FILLER_32_65 ();
 sg13g2_fill_1 FILLER_32_69 ();
 sg13g2_fill_2 FILLER_32_117 ();
 sg13g2_fill_1 FILLER_32_119 ();
 sg13g2_fill_1 FILLER_32_125 ();
 sg13g2_decap_8 FILLER_32_129 ();
 sg13g2_decap_4 FILLER_32_136 ();
 sg13g2_fill_1 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_149 ();
 sg13g2_decap_4 FILLER_32_179 ();
 sg13g2_fill_2 FILLER_32_183 ();
 sg13g2_fill_1 FILLER_32_219 ();
 sg13g2_decap_4 FILLER_32_228 ();
 sg13g2_decap_8 FILLER_32_237 ();
 sg13g2_decap_8 FILLER_32_244 ();
 sg13g2_fill_2 FILLER_32_251 ();
 sg13g2_fill_1 FILLER_32_253 ();
 sg13g2_fill_2 FILLER_32_257 ();
 sg13g2_fill_1 FILLER_32_259 ();
 sg13g2_decap_8 FILLER_32_289 ();
 sg13g2_fill_2 FILLER_32_296 ();
 sg13g2_fill_1 FILLER_32_298 ();
 sg13g2_fill_1 FILLER_32_309 ();
 sg13g2_fill_2 FILLER_32_326 ();
 sg13g2_fill_1 FILLER_32_328 ();
 sg13g2_decap_8 FILLER_32_342 ();
 sg13g2_fill_1 FILLER_32_349 ();
 sg13g2_decap_4 FILLER_32_376 ();
 sg13g2_decap_8 FILLER_32_416 ();
 sg13g2_fill_2 FILLER_32_433 ();
 sg13g2_decap_4 FILLER_32_487 ();
 sg13g2_fill_1 FILLER_32_504 ();
 sg13g2_decap_8 FILLER_32_512 ();
 sg13g2_decap_8 FILLER_32_545 ();
 sg13g2_decap_8 FILLER_32_552 ();
 sg13g2_decap_8 FILLER_32_559 ();
 sg13g2_decap_4 FILLER_32_571 ();
 sg13g2_fill_2 FILLER_32_579 ();
 sg13g2_decap_8 FILLER_32_597 ();
 sg13g2_decap_8 FILLER_32_604 ();
 sg13g2_decap_4 FILLER_32_611 ();
 sg13g2_decap_8 FILLER_32_621 ();
 sg13g2_decap_8 FILLER_32_628 ();
 sg13g2_decap_4 FILLER_32_635 ();
 sg13g2_fill_1 FILLER_32_639 ();
 sg13g2_decap_8 FILLER_32_650 ();
 sg13g2_fill_1 FILLER_32_686 ();
 sg13g2_fill_2 FILLER_32_762 ();
 sg13g2_decap_8 FILLER_32_798 ();
 sg13g2_decap_8 FILLER_32_805 ();
 sg13g2_decap_8 FILLER_32_812 ();
 sg13g2_decap_8 FILLER_32_819 ();
 sg13g2_decap_8 FILLER_32_826 ();
 sg13g2_decap_8 FILLER_32_833 ();
 sg13g2_decap_8 FILLER_32_840 ();
 sg13g2_decap_8 FILLER_32_847 ();
 sg13g2_decap_8 FILLER_32_854 ();
 sg13g2_fill_1 FILLER_32_861 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_14 ();
 sg13g2_decap_4 FILLER_33_29 ();
 sg13g2_fill_1 FILLER_33_33 ();
 sg13g2_decap_8 FILLER_33_39 ();
 sg13g2_decap_4 FILLER_33_46 ();
 sg13g2_fill_1 FILLER_33_50 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_4 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_89 ();
 sg13g2_decap_4 FILLER_33_96 ();
 sg13g2_fill_1 FILLER_33_100 ();
 sg13g2_fill_2 FILLER_33_106 ();
 sg13g2_fill_2 FILLER_33_118 ();
 sg13g2_fill_1 FILLER_33_120 ();
 sg13g2_fill_1 FILLER_33_152 ();
 sg13g2_fill_1 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_4 FILLER_33_217 ();
 sg13g2_fill_2 FILLER_33_221 ();
 sg13g2_decap_8 FILLER_33_246 ();
 sg13g2_decap_8 FILLER_33_253 ();
 sg13g2_fill_1 FILLER_33_260 ();
 sg13g2_fill_2 FILLER_33_264 ();
 sg13g2_fill_1 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_275 ();
 sg13g2_fill_2 FILLER_33_282 ();
 sg13g2_decap_4 FILLER_33_318 ();
 sg13g2_fill_1 FILLER_33_322 ();
 sg13g2_decap_8 FILLER_33_359 ();
 sg13g2_decap_8 FILLER_33_366 ();
 sg13g2_fill_2 FILLER_33_373 ();
 sg13g2_fill_2 FILLER_33_411 ();
 sg13g2_fill_1 FILLER_33_413 ();
 sg13g2_decap_8 FILLER_33_440 ();
 sg13g2_fill_2 FILLER_33_447 ();
 sg13g2_decap_8 FILLER_33_455 ();
 sg13g2_decap_8 FILLER_33_462 ();
 sg13g2_decap_4 FILLER_33_469 ();
 sg13g2_fill_2 FILLER_33_473 ();
 sg13g2_fill_1 FILLER_33_480 ();
 sg13g2_fill_2 FILLER_33_496 ();
 sg13g2_decap_8 FILLER_33_532 ();
 sg13g2_decap_8 FILLER_33_547 ();
 sg13g2_decap_8 FILLER_33_554 ();
 sg13g2_fill_1 FILLER_33_589 ();
 sg13g2_decap_4 FILLER_33_642 ();
 sg13g2_decap_4 FILLER_33_651 ();
 sg13g2_fill_1 FILLER_33_655 ();
 sg13g2_fill_2 FILLER_33_661 ();
 sg13g2_fill_1 FILLER_33_663 ();
 sg13g2_fill_1 FILLER_33_667 ();
 sg13g2_fill_2 FILLER_33_676 ();
 sg13g2_fill_1 FILLER_33_678 ();
 sg13g2_decap_8 FILLER_33_683 ();
 sg13g2_decap_4 FILLER_33_690 ();
 sg13g2_fill_1 FILLER_33_694 ();
 sg13g2_decap_8 FILLER_33_709 ();
 sg13g2_decap_8 FILLER_33_716 ();
 sg13g2_decap_8 FILLER_33_723 ();
 sg13g2_fill_1 FILLER_33_730 ();
 sg13g2_decap_8 FILLER_33_743 ();
 sg13g2_decap_8 FILLER_33_750 ();
 sg13g2_decap_8 FILLER_33_757 ();
 sg13g2_fill_1 FILLER_33_764 ();
 sg13g2_fill_1 FILLER_33_773 ();
 sg13g2_decap_8 FILLER_33_792 ();
 sg13g2_decap_8 FILLER_33_799 ();
 sg13g2_decap_8 FILLER_33_806 ();
 sg13g2_decap_8 FILLER_33_813 ();
 sg13g2_decap_8 FILLER_33_820 ();
 sg13g2_decap_8 FILLER_33_827 ();
 sg13g2_decap_8 FILLER_33_834 ();
 sg13g2_decap_8 FILLER_33_841 ();
 sg13g2_decap_8 FILLER_33_848 ();
 sg13g2_decap_8 FILLER_33_855 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_fill_2 FILLER_34_14 ();
 sg13g2_fill_2 FILLER_34_42 ();
 sg13g2_fill_1 FILLER_34_78 ();
 sg13g2_fill_1 FILLER_34_105 ();
 sg13g2_fill_2 FILLER_34_126 ();
 sg13g2_decap_4 FILLER_34_136 ();
 sg13g2_fill_2 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_146 ();
 sg13g2_decap_8 FILLER_34_153 ();
 sg13g2_fill_2 FILLER_34_160 ();
 sg13g2_decap_8 FILLER_34_167 ();
 sg13g2_fill_1 FILLER_34_174 ();
 sg13g2_decap_8 FILLER_34_201 ();
 sg13g2_fill_2 FILLER_34_234 ();
 sg13g2_fill_1 FILLER_34_236 ();
 sg13g2_fill_2 FILLER_34_246 ();
 sg13g2_fill_1 FILLER_34_284 ();
 sg13g2_fill_1 FILLER_34_311 ();
 sg13g2_fill_1 FILLER_34_338 ();
 sg13g2_fill_2 FILLER_34_365 ();
 sg13g2_fill_1 FILLER_34_367 ();
 sg13g2_decap_8 FILLER_34_388 ();
 sg13g2_decap_8 FILLER_34_395 ();
 sg13g2_decap_4 FILLER_34_402 ();
 sg13g2_fill_1 FILLER_34_406 ();
 sg13g2_decap_8 FILLER_34_427 ();
 sg13g2_decap_4 FILLER_34_434 ();
 sg13g2_fill_1 FILLER_34_438 ();
 sg13g2_decap_8 FILLER_34_491 ();
 sg13g2_fill_1 FILLER_34_506 ();
 sg13g2_decap_8 FILLER_34_514 ();
 sg13g2_decap_4 FILLER_34_521 ();
 sg13g2_fill_1 FILLER_34_525 ();
 sg13g2_fill_1 FILLER_34_562 ();
 sg13g2_decap_8 FILLER_34_568 ();
 sg13g2_decap_8 FILLER_34_575 ();
 sg13g2_fill_2 FILLER_34_582 ();
 sg13g2_fill_1 FILLER_34_584 ();
 sg13g2_decap_8 FILLER_34_603 ();
 sg13g2_decap_4 FILLER_34_610 ();
 sg13g2_decap_8 FILLER_34_626 ();
 sg13g2_fill_2 FILLER_34_633 ();
 sg13g2_fill_2 FILLER_34_656 ();
 sg13g2_fill_2 FILLER_34_689 ();
 sg13g2_decap_4 FILLER_34_711 ();
 sg13g2_fill_1 FILLER_34_715 ();
 sg13g2_decap_8 FILLER_34_724 ();
 sg13g2_decap_4 FILLER_34_770 ();
 sg13g2_decap_8 FILLER_34_800 ();
 sg13g2_decap_8 FILLER_34_807 ();
 sg13g2_decap_8 FILLER_34_814 ();
 sg13g2_decap_8 FILLER_34_821 ();
 sg13g2_decap_8 FILLER_34_828 ();
 sg13g2_decap_8 FILLER_34_835 ();
 sg13g2_decap_8 FILLER_34_842 ();
 sg13g2_decap_8 FILLER_34_849 ();
 sg13g2_decap_4 FILLER_34_856 ();
 sg13g2_fill_2 FILLER_34_860 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_4 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_25 ();
 sg13g2_fill_2 FILLER_35_32 ();
 sg13g2_decap_8 FILLER_35_39 ();
 sg13g2_decap_4 FILLER_35_46 ();
 sg13g2_decap_8 FILLER_35_68 ();
 sg13g2_fill_2 FILLER_35_75 ();
 sg13g2_fill_1 FILLER_35_77 ();
 sg13g2_decap_4 FILLER_35_83 ();
 sg13g2_fill_1 FILLER_35_87 ();
 sg13g2_decap_4 FILLER_35_95 ();
 sg13g2_decap_4 FILLER_35_116 ();
 sg13g2_decap_4 FILLER_35_123 ();
 sg13g2_fill_2 FILLER_35_132 ();
 sg13g2_decap_8 FILLER_35_163 ();
 sg13g2_decap_8 FILLER_35_183 ();
 sg13g2_fill_2 FILLER_35_224 ();
 sg13g2_fill_2 FILLER_35_251 ();
 sg13g2_fill_1 FILLER_35_253 ();
 sg13g2_decap_8 FILLER_35_269 ();
 sg13g2_decap_4 FILLER_35_276 ();
 sg13g2_fill_2 FILLER_35_280 ();
 sg13g2_fill_2 FILLER_35_285 ();
 sg13g2_fill_2 FILLER_35_290 ();
 sg13g2_decap_8 FILLER_35_297 ();
 sg13g2_fill_1 FILLER_35_304 ();
 sg13g2_fill_1 FILLER_35_314 ();
 sg13g2_decap_8 FILLER_35_333 ();
 sg13g2_fill_2 FILLER_35_340 ();
 sg13g2_decap_4 FILLER_35_345 ();
 sg13g2_fill_2 FILLER_35_349 ();
 sg13g2_fill_2 FILLER_35_382 ();
 sg13g2_fill_1 FILLER_35_384 ();
 sg13g2_fill_2 FILLER_35_411 ();
 sg13g2_fill_1 FILLER_35_413 ();
 sg13g2_fill_1 FILLER_35_440 ();
 sg13g2_fill_2 FILLER_35_445 ();
 sg13g2_fill_1 FILLER_35_447 ();
 sg13g2_decap_8 FILLER_35_453 ();
 sg13g2_fill_2 FILLER_35_470 ();
 sg13g2_fill_1 FILLER_35_472 ();
 sg13g2_decap_8 FILLER_35_478 ();
 sg13g2_decap_4 FILLER_35_485 ();
 sg13g2_fill_2 FILLER_35_497 ();
 sg13g2_fill_2 FILLER_35_618 ();
 sg13g2_fill_2 FILLER_35_646 ();
 sg13g2_fill_1 FILLER_35_648 ();
 sg13g2_decap_4 FILLER_35_657 ();
 sg13g2_fill_1 FILLER_35_661 ();
 sg13g2_fill_2 FILLER_35_676 ();
 sg13g2_fill_1 FILLER_35_678 ();
 sg13g2_decap_8 FILLER_35_683 ();
 sg13g2_fill_2 FILLER_35_690 ();
 sg13g2_fill_1 FILLER_35_692 ();
 sg13g2_fill_1 FILLER_35_702 ();
 sg13g2_fill_2 FILLER_35_734 ();
 sg13g2_fill_1 FILLER_35_736 ();
 sg13g2_decap_8 FILLER_35_754 ();
 sg13g2_decap_8 FILLER_35_761 ();
 sg13g2_decap_8 FILLER_35_768 ();
 sg13g2_decap_4 FILLER_35_775 ();
 sg13g2_decap_8 FILLER_35_791 ();
 sg13g2_decap_8 FILLER_35_798 ();
 sg13g2_decap_8 FILLER_35_805 ();
 sg13g2_decap_8 FILLER_35_812 ();
 sg13g2_decap_8 FILLER_35_819 ();
 sg13g2_decap_8 FILLER_35_826 ();
 sg13g2_decap_8 FILLER_35_833 ();
 sg13g2_decap_8 FILLER_35_840 ();
 sg13g2_decap_8 FILLER_35_847 ();
 sg13g2_decap_8 FILLER_35_854 ();
 sg13g2_fill_1 FILLER_35_861 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_77 ();
 sg13g2_fill_1 FILLER_36_79 ();
 sg13g2_fill_1 FILLER_36_106 ();
 sg13g2_decap_8 FILLER_36_143 ();
 sg13g2_decap_4 FILLER_36_150 ();
 sg13g2_fill_1 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_183 ();
 sg13g2_fill_1 FILLER_36_190 ();
 sg13g2_decap_8 FILLER_36_194 ();
 sg13g2_decap_8 FILLER_36_201 ();
 sg13g2_fill_1 FILLER_36_208 ();
 sg13g2_decap_4 FILLER_36_212 ();
 sg13g2_decap_4 FILLER_36_220 ();
 sg13g2_fill_1 FILLER_36_248 ();
 sg13g2_decap_8 FILLER_36_306 ();
 sg13g2_fill_1 FILLER_36_313 ();
 sg13g2_fill_1 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_341 ();
 sg13g2_decap_8 FILLER_36_348 ();
 sg13g2_decap_8 FILLER_36_355 ();
 sg13g2_decap_8 FILLER_36_362 ();
 sg13g2_decap_4 FILLER_36_369 ();
 sg13g2_decap_8 FILLER_36_383 ();
 sg13g2_decap_8 FILLER_36_390 ();
 sg13g2_fill_2 FILLER_36_405 ();
 sg13g2_fill_1 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_36_418 ();
 sg13g2_decap_4 FILLER_36_425 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_decap_8 FILLER_36_435 ();
 sg13g2_fill_1 FILLER_36_442 ();
 sg13g2_fill_2 FILLER_36_480 ();
 sg13g2_decap_8 FILLER_36_500 ();
 sg13g2_fill_2 FILLER_36_507 ();
 sg13g2_decap_8 FILLER_36_521 ();
 sg13g2_fill_2 FILLER_36_528 ();
 sg13g2_fill_1 FILLER_36_530 ();
 sg13g2_fill_1 FILLER_36_541 ();
 sg13g2_decap_8 FILLER_36_545 ();
 sg13g2_decap_4 FILLER_36_552 ();
 sg13g2_fill_2 FILLER_36_556 ();
 sg13g2_fill_2 FILLER_36_563 ();
 sg13g2_fill_1 FILLER_36_565 ();
 sg13g2_fill_2 FILLER_36_571 ();
 sg13g2_decap_8 FILLER_36_577 ();
 sg13g2_fill_1 FILLER_36_584 ();
 sg13g2_fill_2 FILLER_36_594 ();
 sg13g2_fill_1 FILLER_36_596 ();
 sg13g2_decap_8 FILLER_36_601 ();
 sg13g2_decap_4 FILLER_36_608 ();
 sg13g2_fill_2 FILLER_36_612 ();
 sg13g2_decap_8 FILLER_36_624 ();
 sg13g2_decap_8 FILLER_36_631 ();
 sg13g2_fill_2 FILLER_36_638 ();
 sg13g2_fill_1 FILLER_36_640 ();
 sg13g2_fill_2 FILLER_36_688 ();
 sg13g2_decap_8 FILLER_36_703 ();
 sg13g2_fill_2 FILLER_36_714 ();
 sg13g2_fill_1 FILLER_36_716 ();
 sg13g2_decap_8 FILLER_36_722 ();
 sg13g2_decap_8 FILLER_36_729 ();
 sg13g2_decap_4 FILLER_36_736 ();
 sg13g2_fill_2 FILLER_36_745 ();
 sg13g2_fill_1 FILLER_36_747 ();
 sg13g2_decap_8 FILLER_36_774 ();
 sg13g2_fill_2 FILLER_36_781 ();
 sg13g2_fill_1 FILLER_36_783 ();
 sg13g2_decap_8 FILLER_36_794 ();
 sg13g2_decap_8 FILLER_36_801 ();
 sg13g2_decap_8 FILLER_36_808 ();
 sg13g2_decap_8 FILLER_36_815 ();
 sg13g2_decap_8 FILLER_36_822 ();
 sg13g2_decap_8 FILLER_36_829 ();
 sg13g2_decap_8 FILLER_36_836 ();
 sg13g2_decap_8 FILLER_36_843 ();
 sg13g2_decap_8 FILLER_36_850 ();
 sg13g2_decap_4 FILLER_36_857 ();
 sg13g2_fill_1 FILLER_36_861 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_25 ();
 sg13g2_decap_4 FILLER_37_32 ();
 sg13g2_fill_1 FILLER_37_36 ();
 sg13g2_decap_8 FILLER_37_47 ();
 sg13g2_decap_4 FILLER_37_54 ();
 sg13g2_fill_1 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_69 ();
 sg13g2_decap_8 FILLER_37_76 ();
 sg13g2_fill_2 FILLER_37_83 ();
 sg13g2_fill_1 FILLER_37_85 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_4 FILLER_37_98 ();
 sg13g2_fill_1 FILLER_37_102 ();
 sg13g2_decap_8 FILLER_37_118 ();
 sg13g2_decap_4 FILLER_37_125 ();
 sg13g2_fill_1 FILLER_37_129 ();
 sg13g2_decap_8 FILLER_37_137 ();
 sg13g2_fill_2 FILLER_37_144 ();
 sg13g2_fill_1 FILLER_37_146 ();
 sg13g2_fill_1 FILLER_37_151 ();
 sg13g2_fill_2 FILLER_37_169 ();
 sg13g2_fill_1 FILLER_37_171 ();
 sg13g2_decap_8 FILLER_37_220 ();
 sg13g2_fill_1 FILLER_37_227 ();
 sg13g2_decap_8 FILLER_37_248 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_fill_2 FILLER_37_290 ();
 sg13g2_decap_4 FILLER_37_296 ();
 sg13g2_decap_4 FILLER_37_308 ();
 sg13g2_fill_1 FILLER_37_312 ();
 sg13g2_decap_8 FILLER_37_339 ();
 sg13g2_decap_8 FILLER_37_349 ();
 sg13g2_fill_1 FILLER_37_356 ();
 sg13g2_decap_8 FILLER_37_383 ();
 sg13g2_decap_8 FILLER_37_390 ();
 sg13g2_fill_2 FILLER_37_397 ();
 sg13g2_fill_1 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_444 ();
 sg13g2_decap_8 FILLER_37_456 ();
 sg13g2_decap_8 FILLER_37_463 ();
 sg13g2_decap_4 FILLER_37_470 ();
 sg13g2_fill_1 FILLER_37_479 ();
 sg13g2_decap_8 FILLER_37_490 ();
 sg13g2_fill_2 FILLER_37_497 ();
 sg13g2_fill_2 FILLER_37_508 ();
 sg13g2_fill_1 FILLER_37_570 ();
 sg13g2_fill_1 FILLER_37_615 ();
 sg13g2_decap_8 FILLER_37_645 ();
 sg13g2_fill_2 FILLER_37_652 ();
 sg13g2_fill_1 FILLER_37_654 ();
 sg13g2_fill_2 FILLER_37_660 ();
 sg13g2_decap_8 FILLER_37_670 ();
 sg13g2_decap_8 FILLER_37_677 ();
 sg13g2_fill_2 FILLER_37_684 ();
 sg13g2_fill_1 FILLER_37_686 ();
 sg13g2_fill_1 FILLER_37_756 ();
 sg13g2_fill_1 FILLER_37_783 ();
 sg13g2_decap_8 FILLER_37_804 ();
 sg13g2_decap_8 FILLER_37_811 ();
 sg13g2_decap_8 FILLER_37_818 ();
 sg13g2_decap_8 FILLER_37_825 ();
 sg13g2_decap_8 FILLER_37_832 ();
 sg13g2_decap_8 FILLER_37_839 ();
 sg13g2_decap_8 FILLER_37_846 ();
 sg13g2_decap_8 FILLER_37_853 ();
 sg13g2_fill_2 FILLER_37_860 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_4 ();
 sg13g2_fill_1 FILLER_38_14 ();
 sg13g2_fill_1 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_76 ();
 sg13g2_decap_8 FILLER_38_83 ();
 sg13g2_decap_8 FILLER_38_90 ();
 sg13g2_fill_2 FILLER_38_118 ();
 sg13g2_fill_2 FILLER_38_125 ();
 sg13g2_fill_1 FILLER_38_153 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_fill_1 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_219 ();
 sg13g2_decap_8 FILLER_38_226 ();
 sg13g2_fill_1 FILLER_38_233 ();
 sg13g2_fill_1 FILLER_38_244 ();
 sg13g2_decap_8 FILLER_38_307 ();
 sg13g2_decap_8 FILLER_38_314 ();
 sg13g2_fill_1 FILLER_38_321 ();
 sg13g2_decap_4 FILLER_38_327 ();
 sg13g2_fill_1 FILLER_38_331 ();
 sg13g2_decap_8 FILLER_38_368 ();
 sg13g2_fill_2 FILLER_38_375 ();
 sg13g2_fill_1 FILLER_38_413 ();
 sg13g2_decap_4 FILLER_38_471 ();
 sg13g2_decap_8 FILLER_38_531 ();
 sg13g2_decap_8 FILLER_38_538 ();
 sg13g2_decap_8 FILLER_38_545 ();
 sg13g2_decap_8 FILLER_38_552 ();
 sg13g2_decap_4 FILLER_38_559 ();
 sg13g2_fill_1 FILLER_38_563 ();
 sg13g2_fill_1 FILLER_38_568 ();
 sg13g2_fill_2 FILLER_38_586 ();
 sg13g2_fill_1 FILLER_38_588 ();
 sg13g2_decap_8 FILLER_38_592 ();
 sg13g2_decap_8 FILLER_38_599 ();
 sg13g2_decap_4 FILLER_38_606 ();
 sg13g2_fill_1 FILLER_38_610 ();
 sg13g2_decap_8 FILLER_38_624 ();
 sg13g2_decap_4 FILLER_38_631 ();
 sg13g2_fill_1 FILLER_38_635 ();
 sg13g2_fill_2 FILLER_38_649 ();
 sg13g2_fill_1 FILLER_38_651 ();
 sg13g2_decap_4 FILLER_38_660 ();
 sg13g2_fill_1 FILLER_38_664 ();
 sg13g2_decap_8 FILLER_38_673 ();
 sg13g2_decap_4 FILLER_38_689 ();
 sg13g2_fill_1 FILLER_38_693 ();
 sg13g2_fill_1 FILLER_38_703 ();
 sg13g2_decap_8 FILLER_38_708 ();
 sg13g2_decap_4 FILLER_38_715 ();
 sg13g2_decap_8 FILLER_38_724 ();
 sg13g2_decap_8 FILLER_38_731 ();
 sg13g2_decap_4 FILLER_38_738 ();
 sg13g2_decap_4 FILLER_38_747 ();
 sg13g2_fill_1 FILLER_38_759 ();
 sg13g2_decap_8 FILLER_38_765 ();
 sg13g2_decap_8 FILLER_38_772 ();
 sg13g2_decap_8 FILLER_38_779 ();
 sg13g2_fill_2 FILLER_38_786 ();
 sg13g2_decap_4 FILLER_38_796 ();
 sg13g2_decap_8 FILLER_38_808 ();
 sg13g2_decap_8 FILLER_38_815 ();
 sg13g2_decap_8 FILLER_38_822 ();
 sg13g2_decap_8 FILLER_38_829 ();
 sg13g2_decap_8 FILLER_38_836 ();
 sg13g2_decap_8 FILLER_38_843 ();
 sg13g2_decap_8 FILLER_38_850 ();
 sg13g2_decap_4 FILLER_38_857 ();
 sg13g2_fill_1 FILLER_38_861 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_20 ();
 sg13g2_decap_8 FILLER_39_27 ();
 sg13g2_fill_2 FILLER_39_34 ();
 sg13g2_fill_2 FILLER_39_40 ();
 sg13g2_decap_4 FILLER_39_50 ();
 sg13g2_fill_2 FILLER_39_64 ();
 sg13g2_fill_1 FILLER_39_66 ();
 sg13g2_fill_2 FILLER_39_101 ();
 sg13g2_fill_1 FILLER_39_103 ();
 sg13g2_fill_2 FILLER_39_117 ();
 sg13g2_fill_1 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_146 ();
 sg13g2_fill_2 FILLER_39_153 ();
 sg13g2_fill_2 FILLER_39_168 ();
 sg13g2_fill_1 FILLER_39_170 ();
 sg13g2_fill_2 FILLER_39_175 ();
 sg13g2_fill_1 FILLER_39_177 ();
 sg13g2_decap_8 FILLER_39_183 ();
 sg13g2_decap_4 FILLER_39_193 ();
 sg13g2_fill_1 FILLER_39_197 ();
 sg13g2_fill_1 FILLER_39_227 ();
 sg13g2_fill_2 FILLER_39_243 ();
 sg13g2_fill_1 FILLER_39_245 ();
 sg13g2_decap_8 FILLER_39_259 ();
 sg13g2_decap_8 FILLER_39_266 ();
 sg13g2_decap_8 FILLER_39_273 ();
 sg13g2_fill_1 FILLER_39_280 ();
 sg13g2_decap_8 FILLER_39_288 ();
 sg13g2_decap_4 FILLER_39_295 ();
 sg13g2_decap_4 FILLER_39_325 ();
 sg13g2_fill_2 FILLER_39_329 ();
 sg13g2_fill_2 FILLER_39_341 ();
 sg13g2_fill_1 FILLER_39_343 ();
 sg13g2_decap_8 FILLER_39_370 ();
 sg13g2_fill_2 FILLER_39_385 ();
 sg13g2_fill_1 FILLER_39_387 ();
 sg13g2_decap_8 FILLER_39_398 ();
 sg13g2_decap_8 FILLER_39_405 ();
 sg13g2_decap_8 FILLER_39_422 ();
 sg13g2_decap_8 FILLER_39_429 ();
 sg13g2_decap_4 FILLER_39_436 ();
 sg13g2_fill_1 FILLER_39_440 ();
 sg13g2_fill_2 FILLER_39_447 ();
 sg13g2_fill_1 FILLER_39_453 ();
 sg13g2_decap_8 FILLER_39_464 ();
 sg13g2_decap_4 FILLER_39_471 ();
 sg13g2_fill_1 FILLER_39_475 ();
 sg13g2_decap_8 FILLER_39_481 ();
 sg13g2_decap_8 FILLER_39_488 ();
 sg13g2_decap_4 FILLER_39_495 ();
 sg13g2_fill_2 FILLER_39_507 ();
 sg13g2_decap_8 FILLER_39_517 ();
 sg13g2_decap_4 FILLER_39_524 ();
 sg13g2_fill_2 FILLER_39_528 ();
 sg13g2_decap_4 FILLER_39_578 ();
 sg13g2_decap_8 FILLER_39_592 ();
 sg13g2_decap_4 FILLER_39_599 ();
 sg13g2_fill_2 FILLER_39_639 ();
 sg13g2_fill_1 FILLER_39_641 ();
 sg13g2_fill_2 FILLER_39_647 ();
 sg13g2_decap_4 FILLER_39_658 ();
 sg13g2_fill_2 FILLER_39_662 ();
 sg13g2_fill_2 FILLER_39_690 ();
 sg13g2_fill_1 FILLER_39_692 ();
 sg13g2_fill_1 FILLER_39_740 ();
 sg13g2_fill_2 FILLER_39_759 ();
 sg13g2_fill_1 FILLER_39_787 ();
 sg13g2_decap_8 FILLER_39_814 ();
 sg13g2_decap_8 FILLER_39_821 ();
 sg13g2_decap_8 FILLER_39_828 ();
 sg13g2_decap_8 FILLER_39_835 ();
 sg13g2_decap_8 FILLER_39_842 ();
 sg13g2_decap_8 FILLER_39_849 ();
 sg13g2_decap_4 FILLER_39_856 ();
 sg13g2_fill_2 FILLER_39_860 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_75 ();
 sg13g2_decap_8 FILLER_40_82 ();
 sg13g2_decap_8 FILLER_40_89 ();
 sg13g2_fill_1 FILLER_40_96 ();
 sg13g2_decap_4 FILLER_40_119 ();
 sg13g2_fill_1 FILLER_40_123 ();
 sg13g2_decap_4 FILLER_40_128 ();
 sg13g2_fill_2 FILLER_40_132 ();
 sg13g2_fill_1 FILLER_40_163 ();
 sg13g2_fill_2 FILLER_40_210 ();
 sg13g2_fill_1 FILLER_40_212 ();
 sg13g2_fill_1 FILLER_40_257 ();
 sg13g2_decap_4 FILLER_40_291 ();
 sg13g2_fill_2 FILLER_40_295 ();
 sg13g2_decap_8 FILLER_40_302 ();
 sg13g2_fill_2 FILLER_40_309 ();
 sg13g2_fill_1 FILLER_40_311 ();
 sg13g2_decap_8 FILLER_40_351 ();
 sg13g2_fill_2 FILLER_40_358 ();
 sg13g2_fill_2 FILLER_40_386 ();
 sg13g2_fill_1 FILLER_40_388 ();
 sg13g2_fill_2 FILLER_40_467 ();
 sg13g2_fill_2 FILLER_40_477 ();
 sg13g2_fill_1 FILLER_40_479 ();
 sg13g2_fill_2 FILLER_40_495 ();
 sg13g2_fill_2 FILLER_40_540 ();
 sg13g2_fill_1 FILLER_40_542 ();
 sg13g2_decap_8 FILLER_40_546 ();
 sg13g2_decap_8 FILLER_40_553 ();
 sg13g2_fill_2 FILLER_40_560 ();
 sg13g2_fill_1 FILLER_40_562 ();
 sg13g2_fill_1 FILLER_40_581 ();
 sg13g2_fill_2 FILLER_40_611 ();
 sg13g2_fill_1 FILLER_40_613 ();
 sg13g2_decap_8 FILLER_40_617 ();
 sg13g2_decap_8 FILLER_40_624 ();
 sg13g2_fill_2 FILLER_40_631 ();
 sg13g2_fill_2 FILLER_40_643 ();
 sg13g2_fill_1 FILLER_40_652 ();
 sg13g2_fill_2 FILLER_40_661 ();
 sg13g2_decap_4 FILLER_40_668 ();
 sg13g2_fill_1 FILLER_40_672 ();
 sg13g2_decap_8 FILLER_40_677 ();
 sg13g2_decap_8 FILLER_40_684 ();
 sg13g2_decap_8 FILLER_40_708 ();
 sg13g2_decap_8 FILLER_40_715 ();
 sg13g2_decap_8 FILLER_40_722 ();
 sg13g2_decap_8 FILLER_40_729 ();
 sg13g2_decap_4 FILLER_40_736 ();
 sg13g2_fill_1 FILLER_40_740 ();
 sg13g2_fill_1 FILLER_40_761 ();
 sg13g2_decap_4 FILLER_40_788 ();
 sg13g2_fill_1 FILLER_40_810 ();
 sg13g2_decap_8 FILLER_40_837 ();
 sg13g2_decap_8 FILLER_40_844 ();
 sg13g2_decap_8 FILLER_40_851 ();
 sg13g2_decap_4 FILLER_40_858 ();
 sg13g2_decap_4 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_4 ();
 sg13g2_fill_2 FILLER_41_14 ();
 sg13g2_fill_1 FILLER_41_16 ();
 sg13g2_decap_8 FILLER_41_30 ();
 sg13g2_decap_4 FILLER_41_37 ();
 sg13g2_fill_2 FILLER_41_49 ();
 sg13g2_fill_1 FILLER_41_51 ();
 sg13g2_fill_1 FILLER_41_103 ();
 sg13g2_decap_4 FILLER_41_118 ();
 sg13g2_fill_2 FILLER_41_122 ();
 sg13g2_decap_8 FILLER_41_129 ();
 sg13g2_decap_8 FILLER_41_136 ();
 sg13g2_decap_8 FILLER_41_143 ();
 sg13g2_decap_4 FILLER_41_150 ();
 sg13g2_fill_2 FILLER_41_154 ();
 sg13g2_fill_2 FILLER_41_161 ();
 sg13g2_decap_8 FILLER_41_186 ();
 sg13g2_decap_8 FILLER_41_193 ();
 sg13g2_fill_2 FILLER_41_200 ();
 sg13g2_fill_1 FILLER_41_228 ();
 sg13g2_decap_8 FILLER_41_264 ();
 sg13g2_decap_8 FILLER_41_271 ();
 sg13g2_fill_2 FILLER_41_286 ();
 sg13g2_fill_1 FILLER_41_288 ();
 sg13g2_decap_4 FILLER_41_292 ();
 sg13g2_fill_1 FILLER_41_296 ();
 sg13g2_decap_8 FILLER_41_305 ();
 sg13g2_fill_2 FILLER_41_312 ();
 sg13g2_fill_2 FILLER_41_327 ();
 sg13g2_fill_1 FILLER_41_334 ();
 sg13g2_decap_4 FILLER_41_340 ();
 sg13g2_decap_8 FILLER_41_370 ();
 sg13g2_fill_1 FILLER_41_377 ();
 sg13g2_decap_8 FILLER_41_398 ();
 sg13g2_fill_2 FILLER_41_405 ();
 sg13g2_decap_8 FILLER_41_415 ();
 sg13g2_decap_8 FILLER_41_432 ();
 sg13g2_decap_8 FILLER_41_439 ();
 sg13g2_decap_8 FILLER_41_446 ();
 sg13g2_decap_8 FILLER_41_453 ();
 sg13g2_decap_8 FILLER_41_460 ();
 sg13g2_fill_2 FILLER_41_467 ();
 sg13g2_decap_4 FILLER_41_497 ();
 sg13g2_fill_1 FILLER_41_501 ();
 sg13g2_decap_8 FILLER_41_505 ();
 sg13g2_fill_2 FILLER_41_512 ();
 sg13g2_fill_1 FILLER_41_514 ();
 sg13g2_decap_8 FILLER_41_519 ();
 sg13g2_fill_1 FILLER_41_526 ();
 sg13g2_decap_4 FILLER_41_573 ();
 sg13g2_fill_2 FILLER_41_577 ();
 sg13g2_decap_8 FILLER_41_588 ();
 sg13g2_fill_2 FILLER_41_595 ();
 sg13g2_fill_1 FILLER_41_597 ();
 sg13g2_decap_4 FILLER_41_638 ();
 sg13g2_fill_1 FILLER_41_642 ();
 sg13g2_fill_1 FILLER_41_648 ();
 sg13g2_decap_4 FILLER_41_654 ();
 sg13g2_fill_1 FILLER_41_658 ();
 sg13g2_fill_2 FILLER_41_688 ();
 sg13g2_fill_1 FILLER_41_690 ();
 sg13g2_fill_2 FILLER_41_706 ();
 sg13g2_fill_2 FILLER_41_744 ();
 sg13g2_fill_1 FILLER_41_746 ();
 sg13g2_decap_8 FILLER_41_766 ();
 sg13g2_decap_4 FILLER_41_773 ();
 sg13g2_fill_2 FILLER_41_777 ();
 sg13g2_decap_8 FILLER_41_784 ();
 sg13g2_decap_8 FILLER_41_817 ();
 sg13g2_decap_8 FILLER_41_824 ();
 sg13g2_decap_8 FILLER_41_831 ();
 sg13g2_decap_8 FILLER_41_838 ();
 sg13g2_decap_8 FILLER_41_845 ();
 sg13g2_decap_8 FILLER_41_852 ();
 sg13g2_fill_2 FILLER_41_859 ();
 sg13g2_fill_1 FILLER_41_861 ();
 sg13g2_decap_4 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_33 ();
 sg13g2_fill_2 FILLER_42_40 ();
 sg13g2_decap_8 FILLER_42_64 ();
 sg13g2_fill_2 FILLER_42_71 ();
 sg13g2_fill_1 FILLER_42_73 ();
 sg13g2_decap_8 FILLER_42_82 ();
 sg13g2_fill_2 FILLER_42_89 ();
 sg13g2_fill_1 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_4 FILLER_42_164 ();
 sg13g2_fill_1 FILLER_42_168 ();
 sg13g2_decap_8 FILLER_42_194 ();
 sg13g2_decap_4 FILLER_42_201 ();
 sg13g2_fill_2 FILLER_42_205 ();
 sg13g2_decap_8 FILLER_42_210 ();
 sg13g2_decap_8 FILLER_42_217 ();
 sg13g2_fill_2 FILLER_42_229 ();
 sg13g2_fill_1 FILLER_42_231 ();
 sg13g2_decap_8 FILLER_42_241 ();
 sg13g2_decap_8 FILLER_42_248 ();
 sg13g2_fill_2 FILLER_42_255 ();
 sg13g2_decap_8 FILLER_42_267 ();
 sg13g2_fill_1 FILLER_42_274 ();
 sg13g2_decap_4 FILLER_42_311 ();
 sg13g2_fill_1 FILLER_42_336 ();
 sg13g2_decap_8 FILLER_42_350 ();
 sg13g2_fill_2 FILLER_42_357 ();
 sg13g2_decap_4 FILLER_42_385 ();
 sg13g2_fill_1 FILLER_42_389 ();
 sg13g2_decap_8 FILLER_42_452 ();
 sg13g2_decap_4 FILLER_42_459 ();
 sg13g2_fill_1 FILLER_42_463 ();
 sg13g2_decap_4 FILLER_42_477 ();
 sg13g2_fill_1 FILLER_42_489 ();
 sg13g2_decap_8 FILLER_42_551 ();
 sg13g2_fill_1 FILLER_42_558 ();
 sg13g2_decap_4 FILLER_42_564 ();
 sg13g2_fill_2 FILLER_42_568 ();
 sg13g2_fill_2 FILLER_42_575 ();
 sg13g2_fill_2 FILLER_42_606 ();
 sg13g2_fill_1 FILLER_42_608 ();
 sg13g2_decap_8 FILLER_42_612 ();
 sg13g2_decap_8 FILLER_42_619 ();
 sg13g2_decap_4 FILLER_42_626 ();
 sg13g2_fill_2 FILLER_42_630 ();
 sg13g2_fill_1 FILLER_42_645 ();
 sg13g2_decap_4 FILLER_42_656 ();
 sg13g2_fill_1 FILLER_42_660 ();
 sg13g2_fill_2 FILLER_42_666 ();
 sg13g2_fill_1 FILLER_42_668 ();
 sg13g2_decap_8 FILLER_42_677 ();
 sg13g2_decap_8 FILLER_42_684 ();
 sg13g2_fill_1 FILLER_42_698 ();
 sg13g2_fill_2 FILLER_42_713 ();
 sg13g2_decap_8 FILLER_42_720 ();
 sg13g2_decap_8 FILLER_42_727 ();
 sg13g2_decap_8 FILLER_42_734 ();
 sg13g2_decap_4 FILLER_42_741 ();
 sg13g2_fill_2 FILLER_42_789 ();
 sg13g2_fill_1 FILLER_42_791 ();
 sg13g2_decap_8 FILLER_42_813 ();
 sg13g2_decap_8 FILLER_42_820 ();
 sg13g2_decap_8 FILLER_42_827 ();
 sg13g2_decap_8 FILLER_42_834 ();
 sg13g2_decap_8 FILLER_42_841 ();
 sg13g2_decap_8 FILLER_42_848 ();
 sg13g2_decap_8 FILLER_42_855 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_fill_2 FILLER_43_14 ();
 sg13g2_fill_1 FILLER_43_16 ();
 sg13g2_decap_8 FILLER_43_43 ();
 sg13g2_decap_8 FILLER_43_90 ();
 sg13g2_decap_4 FILLER_43_97 ();
 sg13g2_fill_1 FILLER_43_114 ();
 sg13g2_decap_4 FILLER_43_132 ();
 sg13g2_decap_8 FILLER_43_165 ();
 sg13g2_fill_2 FILLER_43_172 ();
 sg13g2_fill_1 FILLER_43_174 ();
 sg13g2_fill_2 FILLER_43_179 ();
 sg13g2_fill_1 FILLER_43_181 ();
 sg13g2_decap_4 FILLER_43_211 ();
 sg13g2_fill_1 FILLER_43_215 ();
 sg13g2_fill_1 FILLER_43_223 ();
 sg13g2_fill_2 FILLER_43_232 ();
 sg13g2_fill_2 FILLER_43_276 ();
 sg13g2_fill_1 FILLER_43_278 ();
 sg13g2_decap_4 FILLER_43_284 ();
 sg13g2_fill_2 FILLER_43_288 ();
 sg13g2_decap_8 FILLER_43_293 ();
 sg13g2_decap_4 FILLER_43_300 ();
 sg13g2_fill_2 FILLER_43_304 ();
 sg13g2_decap_4 FILLER_43_310 ();
 sg13g2_fill_1 FILLER_43_314 ();
 sg13g2_fill_1 FILLER_43_320 ();
 sg13g2_fill_2 FILLER_43_326 ();
 sg13g2_decap_4 FILLER_43_338 ();
 sg13g2_fill_2 FILLER_43_342 ();
 sg13g2_decap_8 FILLER_43_370 ();
 sg13g2_fill_2 FILLER_43_377 ();
 sg13g2_decap_8 FILLER_43_397 ();
 sg13g2_decap_8 FILLER_43_404 ();
 sg13g2_decap_8 FILLER_43_411 ();
 sg13g2_decap_8 FILLER_43_418 ();
 sg13g2_decap_8 FILLER_43_425 ();
 sg13g2_fill_2 FILLER_43_432 ();
 sg13g2_fill_1 FILLER_43_434 ();
 sg13g2_fill_2 FILLER_43_440 ();
 sg13g2_fill_1 FILLER_43_442 ();
 sg13g2_fill_1 FILLER_43_477 ();
 sg13g2_decap_4 FILLER_43_483 ();
 sg13g2_fill_1 FILLER_43_496 ();
 sg13g2_decap_8 FILLER_43_500 ();
 sg13g2_decap_8 FILLER_43_507 ();
 sg13g2_decap_4 FILLER_43_514 ();
 sg13g2_fill_1 FILLER_43_518 ();
 sg13g2_decap_8 FILLER_43_539 ();
 sg13g2_fill_2 FILLER_43_546 ();
 sg13g2_fill_1 FILLER_43_548 ();
 sg13g2_fill_2 FILLER_43_574 ();
 sg13g2_fill_1 FILLER_43_576 ();
 sg13g2_decap_4 FILLER_43_587 ();
 sg13g2_fill_1 FILLER_43_591 ();
 sg13g2_decap_4 FILLER_43_631 ();
 sg13g2_fill_2 FILLER_43_656 ();
 sg13g2_fill_2 FILLER_43_745 ();
 sg13g2_decap_4 FILLER_43_768 ();
 sg13g2_fill_1 FILLER_43_772 ();
 sg13g2_decap_8 FILLER_43_778 ();
 sg13g2_decap_4 FILLER_43_785 ();
 sg13g2_fill_1 FILLER_43_789 ();
 sg13g2_decap_8 FILLER_43_828 ();
 sg13g2_decap_8 FILLER_43_835 ();
 sg13g2_decap_8 FILLER_43_842 ();
 sg13g2_decap_8 FILLER_43_849 ();
 sg13g2_decap_4 FILLER_43_856 ();
 sg13g2_fill_2 FILLER_43_860 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_fill_2 FILLER_44_28 ();
 sg13g2_fill_1 FILLER_44_30 ();
 sg13g2_decap_8 FILLER_44_36 ();
 sg13g2_decap_8 FILLER_44_43 ();
 sg13g2_decap_8 FILLER_44_50 ();
 sg13g2_decap_4 FILLER_44_57 ();
 sg13g2_fill_2 FILLER_44_61 ();
 sg13g2_decap_8 FILLER_44_76 ();
 sg13g2_decap_8 FILLER_44_83 ();
 sg13g2_fill_2 FILLER_44_90 ();
 sg13g2_fill_1 FILLER_44_92 ();
 sg13g2_decap_8 FILLER_44_113 ();
 sg13g2_fill_2 FILLER_44_120 ();
 sg13g2_fill_2 FILLER_44_130 ();
 sg13g2_fill_1 FILLER_44_132 ();
 sg13g2_decap_4 FILLER_44_136 ();
 sg13g2_fill_1 FILLER_44_140 ();
 sg13g2_decap_8 FILLER_44_146 ();
 sg13g2_decap_8 FILLER_44_153 ();
 sg13g2_decap_4 FILLER_44_160 ();
 sg13g2_fill_2 FILLER_44_164 ();
 sg13g2_fill_2 FILLER_44_179 ();
 sg13g2_fill_1 FILLER_44_181 ();
 sg13g2_fill_2 FILLER_44_234 ();
 sg13g2_decap_4 FILLER_44_246 ();
 sg13g2_decap_4 FILLER_44_255 ();
 sg13g2_fill_1 FILLER_44_259 ();
 sg13g2_decap_4 FILLER_44_275 ();
 sg13g2_fill_1 FILLER_44_279 ();
 sg13g2_decap_4 FILLER_44_319 ();
 sg13g2_decap_8 FILLER_44_331 ();
 sg13g2_fill_1 FILLER_44_338 ();
 sg13g2_decap_8 FILLER_44_352 ();
 sg13g2_fill_1 FILLER_44_359 ();
 sg13g2_decap_8 FILLER_44_422 ();
 sg13g2_decap_8 FILLER_44_429 ();
 sg13g2_decap_4 FILLER_44_436 ();
 sg13g2_fill_2 FILLER_44_440 ();
 sg13g2_fill_2 FILLER_44_445 ();
 sg13g2_fill_1 FILLER_44_447 ();
 sg13g2_decap_4 FILLER_44_458 ();
 sg13g2_fill_2 FILLER_44_462 ();
 sg13g2_decap_8 FILLER_44_469 ();
 sg13g2_fill_2 FILLER_44_518 ();
 sg13g2_decap_4 FILLER_44_554 ();
 sg13g2_decap_8 FILLER_44_571 ();
 sg13g2_fill_1 FILLER_44_578 ();
 sg13g2_fill_1 FILLER_44_582 ();
 sg13g2_decap_8 FILLER_44_588 ();
 sg13g2_decap_8 FILLER_44_595 ();
 sg13g2_decap_4 FILLER_44_602 ();
 sg13g2_decap_8 FILLER_44_615 ();
 sg13g2_decap_8 FILLER_44_622 ();
 sg13g2_fill_2 FILLER_44_629 ();
 sg13g2_decap_8 FILLER_44_650 ();
 sg13g2_fill_2 FILLER_44_657 ();
 sg13g2_decap_8 FILLER_44_676 ();
 sg13g2_decap_8 FILLER_44_683 ();
 sg13g2_decap_4 FILLER_44_690 ();
 sg13g2_decap_8 FILLER_44_719 ();
 sg13g2_decap_4 FILLER_44_726 ();
 sg13g2_fill_2 FILLER_44_730 ();
 sg13g2_decap_4 FILLER_44_740 ();
 sg13g2_fill_1 FILLER_44_744 ();
 sg13g2_fill_2 FILLER_44_765 ();
 sg13g2_fill_2 FILLER_44_793 ();
 sg13g2_fill_1 FILLER_44_795 ();
 sg13g2_decap_8 FILLER_44_813 ();
 sg13g2_decap_8 FILLER_44_820 ();
 sg13g2_decap_8 FILLER_44_827 ();
 sg13g2_decap_8 FILLER_44_834 ();
 sg13g2_decap_8 FILLER_44_841 ();
 sg13g2_decap_8 FILLER_44_848 ();
 sg13g2_decap_8 FILLER_44_855 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_fill_2 FILLER_45_14 ();
 sg13g2_fill_1 FILLER_45_16 ();
 sg13g2_fill_2 FILLER_45_63 ();
 sg13g2_decap_4 FILLER_45_91 ();
 sg13g2_fill_2 FILLER_45_99 ();
 sg13g2_decap_4 FILLER_45_114 ();
 sg13g2_fill_2 FILLER_45_118 ();
 sg13g2_fill_2 FILLER_45_177 ();
 sg13g2_fill_1 FILLER_45_179 ();
 sg13g2_decap_8 FILLER_45_193 ();
 sg13g2_decap_8 FILLER_45_200 ();
 sg13g2_fill_2 FILLER_45_207 ();
 sg13g2_fill_1 FILLER_45_209 ();
 sg13g2_decap_8 FILLER_45_218 ();
 sg13g2_fill_1 FILLER_45_225 ();
 sg13g2_decap_4 FILLER_45_272 ();
 sg13g2_decap_4 FILLER_45_312 ();
 sg13g2_fill_1 FILLER_45_316 ();
 sg13g2_fill_2 FILLER_45_340 ();
 sg13g2_decap_8 FILLER_45_350 ();
 sg13g2_decap_8 FILLER_45_357 ();
 sg13g2_decap_8 FILLER_45_364 ();
 sg13g2_decap_8 FILLER_45_371 ();
 sg13g2_decap_8 FILLER_45_474 ();
 sg13g2_decap_4 FILLER_45_481 ();
 sg13g2_decap_8 FILLER_45_493 ();
 sg13g2_fill_1 FILLER_45_500 ();
 sg13g2_decap_8 FILLER_45_504 ();
 sg13g2_decap_8 FILLER_45_511 ();
 sg13g2_decap_8 FILLER_45_518 ();
 sg13g2_decap_8 FILLER_45_525 ();
 sg13g2_decap_8 FILLER_45_532 ();
 sg13g2_decap_8 FILLER_45_539 ();
 sg13g2_fill_1 FILLER_45_546 ();
 sg13g2_decap_4 FILLER_45_552 ();
 sg13g2_decap_4 FILLER_45_569 ();
 sg13g2_fill_1 FILLER_45_604 ();
 sg13g2_decap_8 FILLER_45_635 ();
 sg13g2_decap_8 FILLER_45_642 ();
 sg13g2_fill_2 FILLER_45_649 ();
 sg13g2_fill_1 FILLER_45_651 ();
 sg13g2_fill_2 FILLER_45_692 ();
 sg13g2_fill_1 FILLER_45_694 ();
 sg13g2_fill_2 FILLER_45_709 ();
 sg13g2_fill_1 FILLER_45_711 ();
 sg13g2_fill_1 FILLER_45_717 ();
 sg13g2_decap_8 FILLER_45_765 ();
 sg13g2_decap_8 FILLER_45_772 ();
 sg13g2_fill_2 FILLER_45_779 ();
 sg13g2_fill_2 FILLER_45_786 ();
 sg13g2_fill_1 FILLER_45_788 ();
 sg13g2_fill_2 FILLER_45_806 ();
 sg13g2_fill_1 FILLER_45_808 ();
 sg13g2_decap_8 FILLER_45_835 ();
 sg13g2_decap_8 FILLER_45_842 ();
 sg13g2_decap_8 FILLER_45_849 ();
 sg13g2_decap_4 FILLER_45_856 ();
 sg13g2_fill_2 FILLER_45_860 ();
 sg13g2_decap_8 FILLER_46_26 ();
 sg13g2_decap_8 FILLER_46_33 ();
 sg13g2_fill_2 FILLER_46_40 ();
 sg13g2_decap_8 FILLER_46_62 ();
 sg13g2_fill_1 FILLER_46_69 ();
 sg13g2_decap_4 FILLER_46_79 ();
 sg13g2_fill_1 FILLER_46_83 ();
 sg13g2_fill_2 FILLER_46_96 ();
 sg13g2_fill_1 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_132 ();
 sg13g2_fill_1 FILLER_46_139 ();
 sg13g2_decap_8 FILLER_46_144 ();
 sg13g2_decap_8 FILLER_46_151 ();
 sg13g2_decap_8 FILLER_46_158 ();
 sg13g2_fill_1 FILLER_46_165 ();
 sg13g2_decap_4 FILLER_46_197 ();
 sg13g2_fill_1 FILLER_46_201 ();
 sg13g2_decap_4 FILLER_46_236 ();
 sg13g2_fill_1 FILLER_46_240 ();
 sg13g2_decap_8 FILLER_46_244 ();
 sg13g2_decap_8 FILLER_46_251 ();
 sg13g2_fill_2 FILLER_46_258 ();
 sg13g2_fill_1 FILLER_46_260 ();
 sg13g2_decap_8 FILLER_46_276 ();
 sg13g2_decap_4 FILLER_46_283 ();
 sg13g2_fill_2 FILLER_46_287 ();
 sg13g2_decap_8 FILLER_46_292 ();
 sg13g2_decap_8 FILLER_46_299 ();
 sg13g2_decap_4 FILLER_46_306 ();
 sg13g2_fill_1 FILLER_46_313 ();
 sg13g2_decap_4 FILLER_46_324 ();
 sg13g2_fill_1 FILLER_46_328 ();
 sg13g2_fill_2 FILLER_46_339 ();
 sg13g2_fill_1 FILLER_46_341 ();
 sg13g2_fill_1 FILLER_46_357 ();
 sg13g2_decap_4 FILLER_46_384 ();
 sg13g2_decap_8 FILLER_46_398 ();
 sg13g2_decap_8 FILLER_46_405 ();
 sg13g2_fill_2 FILLER_46_412 ();
 sg13g2_fill_1 FILLER_46_414 ();
 sg13g2_decap_8 FILLER_46_425 ();
 sg13g2_fill_2 FILLER_46_432 ();
 sg13g2_fill_1 FILLER_46_434 ();
 sg13g2_decap_8 FILLER_46_438 ();
 sg13g2_decap_8 FILLER_46_445 ();
 sg13g2_decap_4 FILLER_46_467 ();
 sg13g2_fill_2 FILLER_46_471 ();
 sg13g2_fill_2 FILLER_46_486 ();
 sg13g2_decap_8 FILLER_46_534 ();
 sg13g2_fill_1 FILLER_46_541 ();
 sg13g2_fill_2 FILLER_46_555 ();
 sg13g2_fill_1 FILLER_46_562 ();
 sg13g2_fill_1 FILLER_46_568 ();
 sg13g2_decap_8 FILLER_46_577 ();
 sg13g2_decap_8 FILLER_46_591 ();
 sg13g2_fill_1 FILLER_46_598 ();
 sg13g2_decap_4 FILLER_46_612 ();
 sg13g2_fill_1 FILLER_46_616 ();
 sg13g2_decap_4 FILLER_46_661 ();
 sg13g2_fill_1 FILLER_46_665 ();
 sg13g2_decap_8 FILLER_46_674 ();
 sg13g2_decap_8 FILLER_46_681 ();
 sg13g2_decap_8 FILLER_46_688 ();
 sg13g2_fill_2 FILLER_46_695 ();
 sg13g2_decap_8 FILLER_46_715 ();
 sg13g2_decap_8 FILLER_46_722 ();
 sg13g2_fill_2 FILLER_46_729 ();
 sg13g2_fill_1 FILLER_46_731 ();
 sg13g2_decap_8 FILLER_46_740 ();
 sg13g2_decap_4 FILLER_46_747 ();
 sg13g2_fill_2 FILLER_46_751 ();
 sg13g2_decap_4 FILLER_46_791 ();
 sg13g2_decap_8 FILLER_46_807 ();
 sg13g2_decap_8 FILLER_46_814 ();
 sg13g2_decap_8 FILLER_46_821 ();
 sg13g2_decap_8 FILLER_46_828 ();
 sg13g2_decap_8 FILLER_46_835 ();
 sg13g2_decap_8 FILLER_46_842 ();
 sg13g2_decap_8 FILLER_46_849 ();
 sg13g2_decap_4 FILLER_46_856 ();
 sg13g2_fill_2 FILLER_46_860 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_7 ();
 sg13g2_decap_4 FILLER_47_17 ();
 sg13g2_decap_8 FILLER_47_29 ();
 sg13g2_fill_2 FILLER_47_82 ();
 sg13g2_decap_8 FILLER_47_107 ();
 sg13g2_fill_2 FILLER_47_114 ();
 sg13g2_fill_2 FILLER_47_211 ();
 sg13g2_decap_8 FILLER_47_219 ();
 sg13g2_decap_4 FILLER_47_226 ();
 sg13g2_fill_2 FILLER_47_230 ();
 sg13g2_decap_8 FILLER_47_333 ();
 sg13g2_decap_8 FILLER_47_345 ();
 sg13g2_fill_2 FILLER_47_352 ();
 sg13g2_fill_1 FILLER_47_354 ();
 sg13g2_fill_2 FILLER_47_384 ();
 sg13g2_fill_2 FILLER_47_458 ();
 sg13g2_fill_1 FILLER_47_460 ();
 sg13g2_decap_4 FILLER_47_479 ();
 sg13g2_fill_1 FILLER_47_488 ();
 sg13g2_fill_2 FILLER_47_502 ();
 sg13g2_decap_8 FILLER_47_512 ();
 sg13g2_fill_1 FILLER_47_560 ();
 sg13g2_fill_2 FILLER_47_623 ();
 sg13g2_fill_1 FILLER_47_625 ();
 sg13g2_decap_8 FILLER_47_650 ();
 sg13g2_fill_2 FILLER_47_657 ();
 sg13g2_fill_1 FILLER_47_697 ();
 sg13g2_fill_2 FILLER_47_706 ();
 sg13g2_fill_1 FILLER_47_717 ();
 sg13g2_decap_8 FILLER_47_772 ();
 sg13g2_decap_8 FILLER_47_779 ();
 sg13g2_fill_2 FILLER_47_786 ();
 sg13g2_fill_1 FILLER_47_788 ();
 sg13g2_decap_8 FILLER_47_828 ();
 sg13g2_decap_8 FILLER_47_835 ();
 sg13g2_decap_8 FILLER_47_842 ();
 sg13g2_decap_8 FILLER_47_849 ();
 sg13g2_decap_4 FILLER_47_856 ();
 sg13g2_fill_2 FILLER_47_860 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_7 ();
 sg13g2_fill_1 FILLER_48_9 ();
 sg13g2_decap_8 FILLER_48_34 ();
 sg13g2_decap_4 FILLER_48_41 ();
 sg13g2_decap_8 FILLER_48_64 ();
 sg13g2_decap_8 FILLER_48_71 ();
 sg13g2_fill_2 FILLER_48_78 ();
 sg13g2_fill_1 FILLER_48_103 ();
 sg13g2_decap_8 FILLER_48_108 ();
 sg13g2_decap_8 FILLER_48_115 ();
 sg13g2_decap_8 FILLER_48_122 ();
 sg13g2_fill_1 FILLER_48_129 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_4 FILLER_48_140 ();
 sg13g2_fill_1 FILLER_48_144 ();
 sg13g2_decap_8 FILLER_48_155 ();
 sg13g2_decap_4 FILLER_48_162 ();
 sg13g2_fill_2 FILLER_48_166 ();
 sg13g2_fill_2 FILLER_48_177 ();
 sg13g2_fill_2 FILLER_48_188 ();
 sg13g2_fill_2 FILLER_48_200 ();
 sg13g2_decap_8 FILLER_48_205 ();
 sg13g2_fill_2 FILLER_48_212 ();
 sg13g2_decap_8 FILLER_48_222 ();
 sg13g2_decap_8 FILLER_48_229 ();
 sg13g2_decap_4 FILLER_48_236 ();
 sg13g2_fill_1 FILLER_48_243 ();
 sg13g2_decap_8 FILLER_48_252 ();
 sg13g2_fill_1 FILLER_48_293 ();
 sg13g2_decap_4 FILLER_48_299 ();
 sg13g2_fill_1 FILLER_48_303 ();
 sg13g2_decap_4 FILLER_48_307 ();
 sg13g2_fill_1 FILLER_48_311 ();
 sg13g2_decap_8 FILLER_48_317 ();
 sg13g2_decap_4 FILLER_48_324 ();
 sg13g2_decap_8 FILLER_48_368 ();
 sg13g2_decap_8 FILLER_48_375 ();
 sg13g2_decap_8 FILLER_48_382 ();
 sg13g2_fill_2 FILLER_48_389 ();
 sg13g2_fill_1 FILLER_48_417 ();
 sg13g2_decap_8 FILLER_48_434 ();
 sg13g2_decap_8 FILLER_48_441 ();
 sg13g2_decap_4 FILLER_48_458 ();
 sg13g2_fill_2 FILLER_48_462 ();
 sg13g2_decap_4 FILLER_48_469 ();
 sg13g2_fill_1 FILLER_48_485 ();
 sg13g2_decap_4 FILLER_48_491 ();
 sg13g2_fill_1 FILLER_48_495 ();
 sg13g2_decap_8 FILLER_48_520 ();
 sg13g2_decap_4 FILLER_48_527 ();
 sg13g2_fill_2 FILLER_48_531 ();
 sg13g2_decap_4 FILLER_48_538 ();
 sg13g2_fill_2 FILLER_48_545 ();
 sg13g2_fill_1 FILLER_48_547 ();
 sg13g2_decap_8 FILLER_48_552 ();
 sg13g2_decap_4 FILLER_48_559 ();
 sg13g2_fill_1 FILLER_48_563 ();
 sg13g2_decap_8 FILLER_48_576 ();
 sg13g2_fill_2 FILLER_48_583 ();
 sg13g2_fill_2 FILLER_48_588 ();
 sg13g2_fill_1 FILLER_48_590 ();
 sg13g2_decap_8 FILLER_48_601 ();
 sg13g2_decap_8 FILLER_48_608 ();
 sg13g2_fill_1 FILLER_48_615 ();
 sg13g2_fill_1 FILLER_48_629 ();
 sg13g2_fill_2 FILLER_48_650 ();
 sg13g2_decap_8 FILLER_48_683 ();
 sg13g2_decap_8 FILLER_48_690 ();
 sg13g2_fill_2 FILLER_48_703 ();
 sg13g2_fill_1 FILLER_48_705 ();
 sg13g2_fill_2 FILLER_48_715 ();
 sg13g2_decap_8 FILLER_48_722 ();
 sg13g2_decap_8 FILLER_48_729 ();
 sg13g2_decap_8 FILLER_48_736 ();
 sg13g2_fill_2 FILLER_48_743 ();
 sg13g2_decap_8 FILLER_48_772 ();
 sg13g2_decap_8 FILLER_48_779 ();
 sg13g2_fill_1 FILLER_48_786 ();
 sg13g2_decap_8 FILLER_48_814 ();
 sg13g2_decap_8 FILLER_48_821 ();
 sg13g2_decap_8 FILLER_48_828 ();
 sg13g2_decap_8 FILLER_48_835 ();
 sg13g2_decap_8 FILLER_48_842 ();
 sg13g2_decap_8 FILLER_48_849 ();
 sg13g2_decap_4 FILLER_48_856 ();
 sg13g2_fill_2 FILLER_48_860 ();
 sg13g2_decap_8 FILLER_49_34 ();
 sg13g2_decap_8 FILLER_49_41 ();
 sg13g2_fill_2 FILLER_49_48 ();
 sg13g2_fill_1 FILLER_49_50 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_fill_2 FILLER_49_77 ();
 sg13g2_fill_2 FILLER_49_95 ();
 sg13g2_fill_1 FILLER_49_97 ();
 sg13g2_fill_2 FILLER_49_155 ();
 sg13g2_fill_1 FILLER_49_157 ();
 sg13g2_fill_2 FILLER_49_174 ();
 sg13g2_fill_1 FILLER_49_176 ();
 sg13g2_decap_8 FILLER_49_254 ();
 sg13g2_fill_2 FILLER_49_261 ();
 sg13g2_decap_8 FILLER_49_278 ();
 sg13g2_decap_4 FILLER_49_285 ();
 sg13g2_fill_2 FILLER_49_289 ();
 sg13g2_fill_2 FILLER_49_327 ();
 sg13g2_fill_1 FILLER_49_329 ();
 sg13g2_fill_2 FILLER_49_338 ();
 sg13g2_fill_1 FILLER_49_355 ();
 sg13g2_decap_8 FILLER_49_397 ();
 sg13g2_decap_8 FILLER_49_404 ();
 sg13g2_fill_1 FILLER_49_411 ();
 sg13g2_fill_1 FILLER_49_438 ();
 sg13g2_decap_8 FILLER_49_451 ();
 sg13g2_decap_4 FILLER_49_458 ();
 sg13g2_fill_1 FILLER_49_462 ();
 sg13g2_decap_4 FILLER_49_482 ();
 sg13g2_decap_4 FILLER_49_616 ();
 sg13g2_fill_2 FILLER_49_620 ();
 sg13g2_fill_1 FILLER_49_638 ();
 sg13g2_decap_8 FILLER_49_648 ();
 sg13g2_fill_2 FILLER_49_655 ();
 sg13g2_decap_8 FILLER_49_672 ();
 sg13g2_decap_8 FILLER_49_679 ();
 sg13g2_fill_2 FILLER_49_686 ();
 sg13g2_fill_1 FILLER_49_688 ();
 sg13g2_fill_2 FILLER_49_718 ();
 sg13g2_fill_1 FILLER_49_764 ();
 sg13g2_fill_2 FILLER_49_791 ();
 sg13g2_fill_1 FILLER_49_793 ();
 sg13g2_fill_1 FILLER_49_807 ();
 sg13g2_decap_8 FILLER_49_834 ();
 sg13g2_decap_8 FILLER_49_841 ();
 sg13g2_decap_8 FILLER_49_848 ();
 sg13g2_decap_8 FILLER_49_855 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_fill_1 FILLER_50_14 ();
 sg13g2_fill_2 FILLER_50_27 ();
 sg13g2_fill_2 FILLER_50_55 ();
 sg13g2_fill_1 FILLER_50_57 ();
 sg13g2_decap_4 FILLER_50_76 ();
 sg13g2_fill_1 FILLER_50_80 ();
 sg13g2_fill_2 FILLER_50_98 ();
 sg13g2_fill_1 FILLER_50_100 ();
 sg13g2_decap_8 FILLER_50_109 ();
 sg13g2_decap_8 FILLER_50_116 ();
 sg13g2_decap_4 FILLER_50_123 ();
 sg13g2_fill_2 FILLER_50_127 ();
 sg13g2_decap_8 FILLER_50_132 ();
 sg13g2_decap_4 FILLER_50_139 ();
 sg13g2_fill_1 FILLER_50_143 ();
 sg13g2_decap_8 FILLER_50_153 ();
 sg13g2_decap_4 FILLER_50_160 ();
 sg13g2_fill_1 FILLER_50_164 ();
 sg13g2_fill_2 FILLER_50_178 ();
 sg13g2_decap_8 FILLER_50_190 ();
 sg13g2_decap_4 FILLER_50_197 ();
 sg13g2_decap_8 FILLER_50_204 ();
 sg13g2_decap_8 FILLER_50_211 ();
 sg13g2_decap_8 FILLER_50_218 ();
 sg13g2_decap_4 FILLER_50_225 ();
 sg13g2_decap_4 FILLER_50_232 ();
 sg13g2_fill_2 FILLER_50_236 ();
 sg13g2_decap_8 FILLER_50_245 ();
 sg13g2_fill_2 FILLER_50_274 ();
 sg13g2_decap_4 FILLER_50_296 ();
 sg13g2_fill_1 FILLER_50_300 ();
 sg13g2_decap_8 FILLER_50_304 ();
 sg13g2_decap_8 FILLER_50_311 ();
 sg13g2_decap_4 FILLER_50_318 ();
 sg13g2_fill_2 FILLER_50_322 ();
 sg13g2_fill_2 FILLER_50_327 ();
 sg13g2_decap_8 FILLER_50_358 ();
 sg13g2_decap_8 FILLER_50_365 ();
 sg13g2_decap_8 FILLER_50_372 ();
 sg13g2_fill_2 FILLER_50_379 ();
 sg13g2_fill_1 FILLER_50_381 ();
 sg13g2_fill_1 FILLER_50_427 ();
 sg13g2_fill_2 FILLER_50_454 ();
 sg13g2_fill_1 FILLER_50_456 ();
 sg13g2_fill_2 FILLER_50_470 ();
 sg13g2_fill_1 FILLER_50_472 ();
 sg13g2_fill_1 FILLER_50_481 ();
 sg13g2_decap_8 FILLER_50_497 ();
 sg13g2_decap_8 FILLER_50_521 ();
 sg13g2_decap_4 FILLER_50_528 ();
 sg13g2_fill_2 FILLER_50_532 ();
 sg13g2_fill_2 FILLER_50_566 ();
 sg13g2_fill_1 FILLER_50_568 ();
 sg13g2_decap_8 FILLER_50_572 ();
 sg13g2_decap_8 FILLER_50_579 ();
 sg13g2_decap_4 FILLER_50_586 ();
 sg13g2_fill_1 FILLER_50_590 ();
 sg13g2_decap_4 FILLER_50_594 ();
 sg13g2_fill_2 FILLER_50_598 ();
 sg13g2_decap_4 FILLER_50_604 ();
 sg13g2_fill_2 FILLER_50_608 ();
 sg13g2_fill_1 FILLER_50_635 ();
 sg13g2_decap_8 FILLER_50_685 ();
 sg13g2_fill_1 FILLER_50_692 ();
 sg13g2_fill_2 FILLER_50_714 ();
 sg13g2_fill_1 FILLER_50_716 ();
 sg13g2_decap_8 FILLER_50_721 ();
 sg13g2_decap_8 FILLER_50_728 ();
 sg13g2_decap_8 FILLER_50_735 ();
 sg13g2_decap_4 FILLER_50_742 ();
 sg13g2_fill_1 FILLER_50_746 ();
 sg13g2_decap_8 FILLER_50_768 ();
 sg13g2_decap_8 FILLER_50_775 ();
 sg13g2_decap_4 FILLER_50_782 ();
 sg13g2_fill_2 FILLER_50_786 ();
 sg13g2_fill_2 FILLER_50_800 ();
 sg13g2_fill_1 FILLER_50_802 ();
 sg13g2_decap_8 FILLER_50_815 ();
 sg13g2_decap_8 FILLER_50_822 ();
 sg13g2_decap_8 FILLER_50_829 ();
 sg13g2_decap_8 FILLER_50_836 ();
 sg13g2_decap_8 FILLER_50_843 ();
 sg13g2_decap_8 FILLER_50_850 ();
 sg13g2_decap_4 FILLER_50_857 ();
 sg13g2_fill_1 FILLER_50_861 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_7 ();
 sg13g2_fill_2 FILLER_51_34 ();
 sg13g2_fill_1 FILLER_51_36 ();
 sg13g2_decap_4 FILLER_51_45 ();
 sg13g2_fill_2 FILLER_51_75 ();
 sg13g2_fill_1 FILLER_51_77 ();
 sg13g2_fill_2 FILLER_51_96 ();
 sg13g2_fill_2 FILLER_51_103 ();
 sg13g2_decap_4 FILLER_51_131 ();
 sg13g2_fill_1 FILLER_51_135 ();
 sg13g2_decap_8 FILLER_51_165 ();
 sg13g2_decap_4 FILLER_51_172 ();
 sg13g2_fill_1 FILLER_51_176 ();
 sg13g2_decap_4 FILLER_51_182 ();
 sg13g2_fill_1 FILLER_51_222 ();
 sg13g2_fill_1 FILLER_51_228 ();
 sg13g2_decap_4 FILLER_51_255 ();
 sg13g2_fill_2 FILLER_51_259 ();
 sg13g2_decap_8 FILLER_51_276 ();
 sg13g2_decap_8 FILLER_51_283 ();
 sg13g2_decap_4 FILLER_51_290 ();
 sg13g2_fill_1 FILLER_51_294 ();
 sg13g2_fill_1 FILLER_51_321 ();
 sg13g2_decap_8 FILLER_51_348 ();
 sg13g2_fill_2 FILLER_51_355 ();
 sg13g2_fill_1 FILLER_51_357 ();
 sg13g2_decap_8 FILLER_51_394 ();
 sg13g2_decap_8 FILLER_51_401 ();
 sg13g2_fill_2 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_51_420 ();
 sg13g2_fill_2 FILLER_51_427 ();
 sg13g2_fill_1 FILLER_51_429 ();
 sg13g2_decap_8 FILLER_51_433 ();
 sg13g2_decap_4 FILLER_51_450 ();
 sg13g2_fill_2 FILLER_51_454 ();
 sg13g2_fill_1 FILLER_51_465 ();
 sg13g2_fill_2 FILLER_51_470 ();
 sg13g2_fill_2 FILLER_51_480 ();
 sg13g2_fill_1 FILLER_51_512 ();
 sg13g2_decap_4 FILLER_51_549 ();
 sg13g2_fill_2 FILLER_51_553 ();
 sg13g2_fill_2 FILLER_51_565 ();
 sg13g2_decap_4 FILLER_51_597 ();
 sg13g2_decap_8 FILLER_51_609 ();
 sg13g2_decap_4 FILLER_51_616 ();
 sg13g2_fill_2 FILLER_51_620 ();
 sg13g2_decap_4 FILLER_51_644 ();
 sg13g2_fill_1 FILLER_51_648 ();
 sg13g2_decap_8 FILLER_51_652 ();
 sg13g2_decap_4 FILLER_51_659 ();
 sg13g2_fill_1 FILLER_51_663 ();
 sg13g2_fill_2 FILLER_51_669 ();
 sg13g2_fill_1 FILLER_51_671 ();
 sg13g2_decap_8 FILLER_51_676 ();
 sg13g2_decap_4 FILLER_51_683 ();
 sg13g2_fill_1 FILLER_51_687 ();
 sg13g2_fill_1 FILLER_51_746 ();
 sg13g2_fill_2 FILLER_51_760 ();
 sg13g2_fill_1 FILLER_51_788 ();
 sg13g2_decap_8 FILLER_51_836 ();
 sg13g2_decap_8 FILLER_51_843 ();
 sg13g2_decap_8 FILLER_51_850 ();
 sg13g2_decap_4 FILLER_51_857 ();
 sg13g2_fill_1 FILLER_51_861 ();
 sg13g2_decap_8 FILLER_52_69 ();
 sg13g2_decap_4 FILLER_52_76 ();
 sg13g2_fill_1 FILLER_52_80 ();
 sg13g2_fill_1 FILLER_52_96 ();
 sg13g2_decap_8 FILLER_52_101 ();
 sg13g2_fill_1 FILLER_52_108 ();
 sg13g2_fill_1 FILLER_52_114 ();
 sg13g2_fill_1 FILLER_52_144 ();
 sg13g2_decap_8 FILLER_52_153 ();
 sg13g2_decap_8 FILLER_52_160 ();
 sg13g2_fill_1 FILLER_52_167 ();
 sg13g2_fill_1 FILLER_52_232 ();
 sg13g2_decap_4 FILLER_52_264 ();
 sg13g2_fill_2 FILLER_52_268 ();
 sg13g2_decap_8 FILLER_52_328 ();
 sg13g2_decap_8 FILLER_52_335 ();
 sg13g2_decap_8 FILLER_52_342 ();
 sg13g2_fill_2 FILLER_52_349 ();
 sg13g2_fill_1 FILLER_52_351 ();
 sg13g2_decap_8 FILLER_52_381 ();
 sg13g2_decap_4 FILLER_52_479 ();
 sg13g2_fill_1 FILLER_52_483 ();
 sg13g2_decap_8 FILLER_52_487 ();
 sg13g2_decap_8 FILLER_52_494 ();
 sg13g2_decap_8 FILLER_52_501 ();
 sg13g2_decap_8 FILLER_52_508 ();
 sg13g2_fill_1 FILLER_52_518 ();
 sg13g2_decap_8 FILLER_52_523 ();
 sg13g2_decap_8 FILLER_52_530 ();
 sg13g2_decap_4 FILLER_52_537 ();
 sg13g2_fill_2 FILLER_52_541 ();
 sg13g2_decap_4 FILLER_52_548 ();
 sg13g2_fill_2 FILLER_52_552 ();
 sg13g2_decap_8 FILLER_52_557 ();
 sg13g2_fill_2 FILLER_52_564 ();
 sg13g2_fill_1 FILLER_52_566 ();
 sg13g2_fill_2 FILLER_52_575 ();
 sg13g2_fill_1 FILLER_52_577 ();
 sg13g2_decap_8 FILLER_52_581 ();
 sg13g2_decap_8 FILLER_52_588 ();
 sg13g2_decap_4 FILLER_52_595 ();
 sg13g2_decap_4 FILLER_52_604 ();
 sg13g2_decap_8 FILLER_52_613 ();
 sg13g2_fill_1 FILLER_52_620 ();
 sg13g2_fill_2 FILLER_52_631 ();
 sg13g2_fill_1 FILLER_52_633 ();
 sg13g2_fill_2 FILLER_52_660 ();
 sg13g2_fill_2 FILLER_52_688 ();
 sg13g2_fill_1 FILLER_52_690 ();
 sg13g2_fill_2 FILLER_52_711 ();
 sg13g2_fill_1 FILLER_52_713 ();
 sg13g2_decap_8 FILLER_52_727 ();
 sg13g2_decap_8 FILLER_52_734 ();
 sg13g2_decap_4 FILLER_52_741 ();
 sg13g2_decap_4 FILLER_52_770 ();
 sg13g2_decap_8 FILLER_52_815 ();
 sg13g2_decap_8 FILLER_52_822 ();
 sg13g2_decap_8 FILLER_52_829 ();
 sg13g2_decap_8 FILLER_52_836 ();
 sg13g2_decap_8 FILLER_52_843 ();
 sg13g2_decap_8 FILLER_52_850 ();
 sg13g2_decap_4 FILLER_52_857 ();
 sg13g2_fill_1 FILLER_52_861 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_45 ();
 sg13g2_decap_8 FILLER_53_52 ();
 sg13g2_decap_8 FILLER_53_59 ();
 sg13g2_decap_4 FILLER_53_66 ();
 sg13g2_fill_2 FILLER_53_78 ();
 sg13g2_decap_8 FILLER_53_112 ();
 sg13g2_fill_2 FILLER_53_119 ();
 sg13g2_fill_1 FILLER_53_121 ();
 sg13g2_decap_8 FILLER_53_129 ();
 sg13g2_fill_2 FILLER_53_166 ();
 sg13g2_fill_1 FILLER_53_168 ();
 sg13g2_decap_8 FILLER_53_190 ();
 sg13g2_decap_8 FILLER_53_197 ();
 sg13g2_fill_1 FILLER_53_204 ();
 sg13g2_decap_4 FILLER_53_210 ();
 sg13g2_fill_2 FILLER_53_214 ();
 sg13g2_decap_4 FILLER_53_222 ();
 sg13g2_decap_8 FILLER_53_234 ();
 sg13g2_decap_8 FILLER_53_241 ();
 sg13g2_fill_1 FILLER_53_248 ();
 sg13g2_decap_4 FILLER_53_256 ();
 sg13g2_fill_2 FILLER_53_260 ();
 sg13g2_fill_1 FILLER_53_272 ();
 sg13g2_decap_8 FILLER_53_288 ();
 sg13g2_decap_8 FILLER_53_310 ();
 sg13g2_decap_8 FILLER_53_317 ();
 sg13g2_fill_1 FILLER_53_324 ();
 sg13g2_decap_8 FILLER_53_330 ();
 sg13g2_fill_1 FILLER_53_347 ();
 sg13g2_decap_8 FILLER_53_399 ();
 sg13g2_decap_8 FILLER_53_406 ();
 sg13g2_decap_8 FILLER_53_413 ();
 sg13g2_decap_8 FILLER_53_420 ();
 sg13g2_decap_8 FILLER_53_427 ();
 sg13g2_decap_8 FILLER_53_434 ();
 sg13g2_decap_8 FILLER_53_441 ();
 sg13g2_decap_8 FILLER_53_448 ();
 sg13g2_decap_8 FILLER_53_455 ();
 sg13g2_decap_8 FILLER_53_467 ();
 sg13g2_decap_8 FILLER_53_474 ();
 sg13g2_fill_2 FILLER_53_481 ();
 sg13g2_fill_1 FILLER_53_487 ();
 sg13g2_decap_4 FILLER_53_506 ();
 sg13g2_fill_1 FILLER_53_539 ();
 sg13g2_decap_8 FILLER_53_637 ();
 sg13g2_decap_8 FILLER_53_644 ();
 sg13g2_decap_4 FILLER_53_656 ();
 sg13g2_fill_1 FILLER_53_660 ();
 sg13g2_fill_2 FILLER_53_669 ();
 sg13g2_fill_1 FILLER_53_671 ();
 sg13g2_fill_1 FILLER_53_676 ();
 sg13g2_decap_8 FILLER_53_682 ();
 sg13g2_fill_1 FILLER_53_689 ();
 sg13g2_fill_1 FILLER_53_706 ();
 sg13g2_decap_4 FILLER_53_714 ();
 sg13g2_decap_8 FILLER_53_744 ();
 sg13g2_fill_2 FILLER_53_751 ();
 sg13g2_fill_2 FILLER_53_758 ();
 sg13g2_fill_1 FILLER_53_760 ();
 sg13g2_fill_2 FILLER_53_787 ();
 sg13g2_fill_1 FILLER_53_789 ();
 sg13g2_decap_8 FILLER_53_810 ();
 sg13g2_decap_8 FILLER_53_817 ();
 sg13g2_decap_8 FILLER_53_824 ();
 sg13g2_decap_8 FILLER_53_831 ();
 sg13g2_decap_8 FILLER_53_838 ();
 sg13g2_decap_8 FILLER_53_845 ();
 sg13g2_decap_8 FILLER_53_852 ();
 sg13g2_fill_2 FILLER_53_859 ();
 sg13g2_fill_1 FILLER_53_861 ();
 sg13g2_decap_8 FILLER_54_30 ();
 sg13g2_decap_8 FILLER_54_37 ();
 sg13g2_decap_4 FILLER_54_44 ();
 sg13g2_fill_2 FILLER_54_53 ();
 sg13g2_fill_1 FILLER_54_55 ();
 sg13g2_fill_1 FILLER_54_73 ();
 sg13g2_decap_8 FILLER_54_97 ();
 sg13g2_decap_4 FILLER_54_104 ();
 sg13g2_decap_8 FILLER_54_138 ();
 sg13g2_fill_2 FILLER_54_145 ();
 sg13g2_decap_8 FILLER_54_155 ();
 sg13g2_fill_2 FILLER_54_162 ();
 sg13g2_fill_1 FILLER_54_164 ();
 sg13g2_fill_1 FILLER_54_198 ();
 sg13g2_decap_4 FILLER_54_251 ();
 sg13g2_fill_2 FILLER_54_255 ();
 sg13g2_decap_4 FILLER_54_262 ();
 sg13g2_fill_1 FILLER_54_266 ();
 sg13g2_fill_2 FILLER_54_282 ();
 sg13g2_fill_1 FILLER_54_284 ();
 sg13g2_fill_2 FILLER_54_288 ();
 sg13g2_fill_1 FILLER_54_290 ();
 sg13g2_fill_2 FILLER_54_294 ();
 sg13g2_fill_1 FILLER_54_296 ();
 sg13g2_fill_2 FILLER_54_346 ();
 sg13g2_decap_8 FILLER_54_361 ();
 sg13g2_decap_8 FILLER_54_368 ();
 sg13g2_decap_4 FILLER_54_375 ();
 sg13g2_fill_2 FILLER_54_379 ();
 sg13g2_decap_4 FILLER_54_401 ();
 sg13g2_decap_8 FILLER_54_441 ();
 sg13g2_fill_2 FILLER_54_448 ();
 sg13g2_fill_1 FILLER_54_450 ();
 sg13g2_fill_1 FILLER_54_456 ();
 sg13g2_fill_2 FILLER_54_526 ();
 sg13g2_fill_2 FILLER_54_561 ();
 sg13g2_decap_8 FILLER_54_567 ();
 sg13g2_fill_2 FILLER_54_574 ();
 sg13g2_fill_1 FILLER_54_576 ();
 sg13g2_decap_4 FILLER_54_580 ();
 sg13g2_fill_1 FILLER_54_584 ();
 sg13g2_fill_2 FILLER_54_590 ();
 sg13g2_fill_1 FILLER_54_592 ();
 sg13g2_decap_8 FILLER_54_597 ();
 sg13g2_decap_8 FILLER_54_604 ();
 sg13g2_fill_1 FILLER_54_611 ();
 sg13g2_fill_1 FILLER_54_706 ();
 sg13g2_fill_1 FILLER_54_720 ();
 sg13g2_decap_8 FILLER_54_747 ();
 sg13g2_decap_8 FILLER_54_762 ();
 sg13g2_decap_8 FILLER_54_769 ();
 sg13g2_decap_8 FILLER_54_776 ();
 sg13g2_decap_8 FILLER_54_783 ();
 sg13g2_decap_8 FILLER_54_790 ();
 sg13g2_decap_8 FILLER_54_797 ();
 sg13g2_decap_8 FILLER_54_804 ();
 sg13g2_decap_8 FILLER_54_811 ();
 sg13g2_decap_8 FILLER_54_818 ();
 sg13g2_decap_8 FILLER_54_825 ();
 sg13g2_decap_8 FILLER_54_832 ();
 sg13g2_decap_8 FILLER_54_839 ();
 sg13g2_decap_8 FILLER_54_846 ();
 sg13g2_decap_8 FILLER_54_853 ();
 sg13g2_fill_2 FILLER_54_860 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_fill_2 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_66 ();
 sg13g2_decap_4 FILLER_55_73 ();
 sg13g2_fill_1 FILLER_55_77 ();
 sg13g2_fill_1 FILLER_55_90 ();
 sg13g2_fill_1 FILLER_55_109 ();
 sg13g2_fill_1 FILLER_55_122 ();
 sg13g2_fill_2 FILLER_55_159 ();
 sg13g2_fill_2 FILLER_55_166 ();
 sg13g2_fill_1 FILLER_55_168 ();
 sg13g2_decap_8 FILLER_55_190 ();
 sg13g2_decap_4 FILLER_55_197 ();
 sg13g2_fill_2 FILLER_55_201 ();
 sg13g2_decap_8 FILLER_55_210 ();
 sg13g2_decap_8 FILLER_55_217 ();
 sg13g2_fill_2 FILLER_55_224 ();
 sg13g2_fill_1 FILLER_55_226 ();
 sg13g2_decap_8 FILLER_55_230 ();
 sg13g2_decap_4 FILLER_55_237 ();
 sg13g2_decap_4 FILLER_55_249 ();
 sg13g2_fill_1 FILLER_55_253 ();
 sg13g2_fill_2 FILLER_55_267 ();
 sg13g2_fill_1 FILLER_55_269 ();
 sg13g2_fill_2 FILLER_55_302 ();
 sg13g2_fill_1 FILLER_55_304 ();
 sg13g2_decap_8 FILLER_55_308 ();
 sg13g2_decap_8 FILLER_55_315 ();
 sg13g2_fill_2 FILLER_55_322 ();
 sg13g2_fill_1 FILLER_55_324 ();
 sg13g2_decap_8 FILLER_55_330 ();
 sg13g2_decap_4 FILLER_55_337 ();
 sg13g2_decap_4 FILLER_55_367 ();
 sg13g2_fill_2 FILLER_55_371 ();
 sg13g2_fill_1 FILLER_55_376 ();
 sg13g2_decap_8 FILLER_55_415 ();
 sg13g2_fill_2 FILLER_55_422 ();
 sg13g2_fill_1 FILLER_55_424 ();
 sg13g2_fill_2 FILLER_55_469 ();
 sg13g2_fill_2 FILLER_55_483 ();
 sg13g2_fill_1 FILLER_55_485 ();
 sg13g2_decap_4 FILLER_55_496 ();
 sg13g2_fill_1 FILLER_55_500 ();
 sg13g2_fill_1 FILLER_55_516 ();
 sg13g2_decap_8 FILLER_55_520 ();
 sg13g2_fill_2 FILLER_55_527 ();
 sg13g2_fill_1 FILLER_55_529 ();
 sg13g2_decap_4 FILLER_55_543 ();
 sg13g2_fill_1 FILLER_55_547 ();
 sg13g2_fill_1 FILLER_55_553 ();
 sg13g2_fill_1 FILLER_55_624 ();
 sg13g2_decap_4 FILLER_55_640 ();
 sg13g2_decap_8 FILLER_55_647 ();
 sg13g2_decap_4 FILLER_55_654 ();
 sg13g2_fill_1 FILLER_55_658 ();
 sg13g2_fill_1 FILLER_55_662 ();
 sg13g2_decap_8 FILLER_55_668 ();
 sg13g2_decap_8 FILLER_55_675 ();
 sg13g2_fill_2 FILLER_55_682 ();
 sg13g2_fill_2 FILLER_55_710 ();
 sg13g2_fill_2 FILLER_55_748 ();
 sg13g2_fill_2 FILLER_55_762 ();
 sg13g2_decap_8 FILLER_55_798 ();
 sg13g2_decap_8 FILLER_55_805 ();
 sg13g2_decap_8 FILLER_55_812 ();
 sg13g2_decap_8 FILLER_55_819 ();
 sg13g2_decap_8 FILLER_55_826 ();
 sg13g2_decap_8 FILLER_55_833 ();
 sg13g2_decap_8 FILLER_55_840 ();
 sg13g2_decap_8 FILLER_55_847 ();
 sg13g2_decap_8 FILLER_55_854 ();
 sg13g2_fill_1 FILLER_55_861 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_4 FILLER_56_28 ();
 sg13g2_fill_2 FILLER_56_37 ();
 sg13g2_fill_1 FILLER_56_39 ();
 sg13g2_fill_2 FILLER_56_49 ();
 sg13g2_decap_4 FILLER_56_71 ();
 sg13g2_fill_2 FILLER_56_75 ();
 sg13g2_fill_2 FILLER_56_93 ();
 sg13g2_fill_2 FILLER_56_103 ();
 sg13g2_decap_4 FILLER_56_123 ();
 sg13g2_decap_8 FILLER_56_138 ();
 sg13g2_decap_8 FILLER_56_145 ();
 sg13g2_decap_8 FILLER_56_152 ();
 sg13g2_decap_4 FILLER_56_159 ();
 sg13g2_fill_1 FILLER_56_163 ();
 sg13g2_fill_1 FILLER_56_176 ();
 sg13g2_fill_2 FILLER_56_231 ();
 sg13g2_fill_1 FILLER_56_233 ();
 sg13g2_fill_1 FILLER_56_238 ();
 sg13g2_decap_8 FILLER_56_244 ();
 sg13g2_fill_1 FILLER_56_251 ();
 sg13g2_decap_8 FILLER_56_255 ();
 sg13g2_fill_1 FILLER_56_262 ();
 sg13g2_fill_2 FILLER_56_273 ();
 sg13g2_fill_1 FILLER_56_275 ();
 sg13g2_decap_4 FILLER_56_281 ();
 sg13g2_fill_2 FILLER_56_345 ();
 sg13g2_fill_2 FILLER_56_365 ();
 sg13g2_fill_2 FILLER_56_377 ();
 sg13g2_decap_8 FILLER_56_420 ();
 sg13g2_decap_8 FILLER_56_427 ();
 sg13g2_decap_8 FILLER_56_437 ();
 sg13g2_decap_8 FILLER_56_444 ();
 sg13g2_decap_8 FILLER_56_451 ();
 sg13g2_fill_1 FILLER_56_458 ();
 sg13g2_decap_4 FILLER_56_479 ();
 sg13g2_fill_2 FILLER_56_483 ();
 sg13g2_fill_2 FILLER_56_511 ();
 sg13g2_fill_2 FILLER_56_547 ();
 sg13g2_fill_2 FILLER_56_554 ();
 sg13g2_decap_8 FILLER_56_561 ();
 sg13g2_decap_8 FILLER_56_568 ();
 sg13g2_fill_1 FILLER_56_575 ();
 sg13g2_decap_4 FILLER_56_579 ();
 sg13g2_decap_4 FILLER_56_586 ();
 sg13g2_fill_1 FILLER_56_590 ();
 sg13g2_decap_8 FILLER_56_601 ();
 sg13g2_decap_4 FILLER_56_608 ();
 sg13g2_fill_1 FILLER_56_612 ();
 sg13g2_fill_1 FILLER_56_622 ();
 sg13g2_decap_4 FILLER_56_632 ();
 sg13g2_fill_2 FILLER_56_636 ();
 sg13g2_fill_1 FILLER_56_643 ();
 sg13g2_decap_4 FILLER_56_647 ();
 sg13g2_fill_1 FILLER_56_651 ();
 sg13g2_decap_8 FILLER_56_681 ();
 sg13g2_fill_1 FILLER_56_688 ();
 sg13g2_decap_8 FILLER_56_710 ();
 sg13g2_decap_8 FILLER_56_717 ();
 sg13g2_decap_8 FILLER_56_724 ();
 sg13g2_decap_8 FILLER_56_731 ();
 sg13g2_decap_8 FILLER_56_738 ();
 sg13g2_decap_4 FILLER_56_745 ();
 sg13g2_fill_1 FILLER_56_749 ();
 sg13g2_decap_8 FILLER_56_776 ();
 sg13g2_decap_8 FILLER_56_783 ();
 sg13g2_decap_8 FILLER_56_790 ();
 sg13g2_decap_8 FILLER_56_797 ();
 sg13g2_decap_8 FILLER_56_804 ();
 sg13g2_decap_8 FILLER_56_811 ();
 sg13g2_decap_8 FILLER_56_818 ();
 sg13g2_decap_8 FILLER_56_825 ();
 sg13g2_decap_8 FILLER_56_832 ();
 sg13g2_decap_8 FILLER_56_839 ();
 sg13g2_decap_8 FILLER_56_846 ();
 sg13g2_decap_8 FILLER_56_853 ();
 sg13g2_fill_2 FILLER_56_860 ();
 sg13g2_fill_2 FILLER_57_26 ();
 sg13g2_fill_1 FILLER_57_28 ();
 sg13g2_fill_2 FILLER_57_36 ();
 sg13g2_fill_1 FILLER_57_38 ();
 sg13g2_fill_1 FILLER_57_53 ();
 sg13g2_decap_8 FILLER_57_92 ();
 sg13g2_decap_4 FILLER_57_99 ();
 sg13g2_decap_4 FILLER_57_129 ();
 sg13g2_decap_4 FILLER_57_171 ();
 sg13g2_fill_2 FILLER_57_175 ();
 sg13g2_fill_1 FILLER_57_182 ();
 sg13g2_fill_2 FILLER_57_188 ();
 sg13g2_fill_1 FILLER_57_190 ();
 sg13g2_decap_8 FILLER_57_201 ();
 sg13g2_decap_8 FILLER_57_211 ();
 sg13g2_decap_8 FILLER_57_218 ();
 sg13g2_fill_2 FILLER_57_285 ();
 sg13g2_decap_4 FILLER_57_292 ();
 sg13g2_fill_2 FILLER_57_296 ();
 sg13g2_decap_8 FILLER_57_304 ();
 sg13g2_decap_8 FILLER_57_311 ();
 sg13g2_decap_4 FILLER_57_318 ();
 sg13g2_fill_1 FILLER_57_330 ();
 sg13g2_fill_2 FILLER_57_334 ();
 sg13g2_fill_1 FILLER_57_336 ();
 sg13g2_decap_8 FILLER_57_366 ();
 sg13g2_decap_8 FILLER_57_373 ();
 sg13g2_decap_8 FILLER_57_393 ();
 sg13g2_decap_8 FILLER_57_400 ();
 sg13g2_decap_4 FILLER_57_474 ();
 sg13g2_decap_8 FILLER_57_494 ();
 sg13g2_decap_8 FILLER_57_501 ();
 sg13g2_decap_8 FILLER_57_508 ();
 sg13g2_decap_4 FILLER_57_515 ();
 sg13g2_fill_1 FILLER_57_519 ();
 sg13g2_decap_8 FILLER_57_525 ();
 sg13g2_decap_4 FILLER_57_532 ();
 sg13g2_fill_1 FILLER_57_544 ();
 sg13g2_fill_1 FILLER_57_574 ();
 sg13g2_decap_4 FILLER_57_601 ();
 sg13g2_fill_1 FILLER_57_605 ();
 sg13g2_fill_1 FILLER_57_616 ();
 sg13g2_fill_2 FILLER_57_622 ();
 sg13g2_fill_1 FILLER_57_640 ();
 sg13g2_fill_1 FILLER_57_671 ();
 sg13g2_decap_8 FILLER_57_676 ();
 sg13g2_fill_1 FILLER_57_683 ();
 sg13g2_fill_2 FILLER_57_704 ();
 sg13g2_fill_1 FILLER_57_706 ();
 sg13g2_decap_4 FILLER_57_724 ();
 sg13g2_decap_4 FILLER_57_736 ();
 sg13g2_fill_1 FILLER_57_740 ();
 sg13g2_decap_8 FILLER_57_799 ();
 sg13g2_decap_8 FILLER_57_806 ();
 sg13g2_decap_8 FILLER_57_813 ();
 sg13g2_decap_8 FILLER_57_820 ();
 sg13g2_decap_8 FILLER_57_827 ();
 sg13g2_decap_8 FILLER_57_834 ();
 sg13g2_decap_8 FILLER_57_841 ();
 sg13g2_decap_8 FILLER_57_848 ();
 sg13g2_decap_8 FILLER_57_855 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_fill_1 FILLER_58_21 ();
 sg13g2_fill_2 FILLER_58_27 ();
 sg13g2_decap_8 FILLER_58_48 ();
 sg13g2_decap_4 FILLER_58_55 ();
 sg13g2_fill_2 FILLER_58_59 ();
 sg13g2_decap_4 FILLER_58_73 ();
 sg13g2_fill_2 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_97 ();
 sg13g2_fill_1 FILLER_58_130 ();
 sg13g2_fill_1 FILLER_58_163 ();
 sg13g2_decap_8 FILLER_58_189 ();
 sg13g2_fill_2 FILLER_58_196 ();
 sg13g2_fill_2 FILLER_58_227 ();
 sg13g2_fill_1 FILLER_58_229 ();
 sg13g2_fill_1 FILLER_58_235 ();
 sg13g2_decap_8 FILLER_58_244 ();
 sg13g2_decap_8 FILLER_58_251 ();
 sg13g2_decap_4 FILLER_58_258 ();
 sg13g2_fill_1 FILLER_58_262 ();
 sg13g2_fill_2 FILLER_58_280 ();
 sg13g2_fill_2 FILLER_58_323 ();
 sg13g2_fill_2 FILLER_58_355 ();
 sg13g2_fill_1 FILLER_58_393 ();
 sg13g2_decap_4 FILLER_58_404 ();
 sg13g2_decap_8 FILLER_58_442 ();
 sg13g2_decap_4 FILLER_58_449 ();
 sg13g2_fill_2 FILLER_58_453 ();
 sg13g2_fill_1 FILLER_58_463 ();
 sg13g2_fill_1 FILLER_58_481 ();
 sg13g2_decap_4 FILLER_58_486 ();
 sg13g2_fill_2 FILLER_58_490 ();
 sg13g2_decap_8 FILLER_58_512 ();
 sg13g2_decap_4 FILLER_58_519 ();
 sg13g2_fill_1 FILLER_58_523 ();
 sg13g2_decap_4 FILLER_58_529 ();
 sg13g2_decap_8 FILLER_58_542 ();
 sg13g2_fill_2 FILLER_58_549 ();
 sg13g2_fill_1 FILLER_58_551 ();
 sg13g2_decap_8 FILLER_58_561 ();
 sg13g2_decap_8 FILLER_58_568 ();
 sg13g2_decap_4 FILLER_58_575 ();
 sg13g2_decap_8 FILLER_58_582 ();
 sg13g2_decap_4 FILLER_58_589 ();
 sg13g2_fill_1 FILLER_58_593 ();
 sg13g2_decap_4 FILLER_58_604 ();
 sg13g2_decap_4 FILLER_58_634 ();
 sg13g2_fill_1 FILLER_58_646 ();
 sg13g2_decap_8 FILLER_58_660 ();
 sg13g2_decap_8 FILLER_58_667 ();
 sg13g2_fill_2 FILLER_58_674 ();
 sg13g2_fill_2 FILLER_58_715 ();
 sg13g2_fill_1 FILLER_58_717 ();
 sg13g2_decap_4 FILLER_58_744 ();
 sg13g2_fill_2 FILLER_58_748 ();
 sg13g2_fill_1 FILLER_58_754 ();
 sg13g2_decap_8 FILLER_58_768 ();
 sg13g2_decap_8 FILLER_58_775 ();
 sg13g2_decap_8 FILLER_58_782 ();
 sg13g2_decap_8 FILLER_58_789 ();
 sg13g2_decap_8 FILLER_58_796 ();
 sg13g2_decap_8 FILLER_58_803 ();
 sg13g2_decap_8 FILLER_58_810 ();
 sg13g2_decap_8 FILLER_58_817 ();
 sg13g2_decap_8 FILLER_58_824 ();
 sg13g2_decap_8 FILLER_58_831 ();
 sg13g2_decap_8 FILLER_58_838 ();
 sg13g2_decap_8 FILLER_58_845 ();
 sg13g2_decap_8 FILLER_58_852 ();
 sg13g2_fill_2 FILLER_58_859 ();
 sg13g2_fill_1 FILLER_58_861 ();
 sg13g2_fill_2 FILLER_59_26 ();
 sg13g2_fill_2 FILLER_59_53 ();
 sg13g2_fill_1 FILLER_59_55 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_4 FILLER_59_77 ();
 sg13g2_fill_2 FILLER_59_81 ();
 sg13g2_decap_8 FILLER_59_101 ();
 sg13g2_fill_2 FILLER_59_108 ();
 sg13g2_fill_1 FILLER_59_110 ();
 sg13g2_decap_8 FILLER_59_119 ();
 sg13g2_decap_4 FILLER_59_126 ();
 sg13g2_fill_2 FILLER_59_130 ();
 sg13g2_decap_8 FILLER_59_135 ();
 sg13g2_fill_2 FILLER_59_142 ();
 sg13g2_decap_8 FILLER_59_150 ();
 sg13g2_fill_2 FILLER_59_157 ();
 sg13g2_fill_2 FILLER_59_164 ();
 sg13g2_decap_4 FILLER_59_212 ();
 sg13g2_decap_8 FILLER_59_253 ();
 sg13g2_decap_8 FILLER_59_260 ();
 sg13g2_fill_2 FILLER_59_267 ();
 sg13g2_decap_4 FILLER_59_291 ();
 sg13g2_fill_2 FILLER_59_295 ();
 sg13g2_decap_4 FILLER_59_300 ();
 sg13g2_fill_1 FILLER_59_304 ();
 sg13g2_decap_8 FILLER_59_310 ();
 sg13g2_decap_8 FILLER_59_317 ();
 sg13g2_decap_8 FILLER_59_324 ();
 sg13g2_fill_1 FILLER_59_331 ();
 sg13g2_decap_8 FILLER_59_337 ();
 sg13g2_fill_1 FILLER_59_344 ();
 sg13g2_decap_8 FILLER_59_353 ();
 sg13g2_decap_4 FILLER_59_360 ();
 sg13g2_fill_2 FILLER_59_364 ();
 sg13g2_decap_8 FILLER_59_369 ();
 sg13g2_decap_4 FILLER_59_376 ();
 sg13g2_fill_2 FILLER_59_380 ();
 sg13g2_decap_4 FILLER_59_387 ();
 sg13g2_fill_1 FILLER_59_391 ();
 sg13g2_fill_1 FILLER_59_428 ();
 sg13g2_fill_1 FILLER_59_465 ();
 sg13g2_fill_2 FILLER_59_550 ();
 sg13g2_decap_4 FILLER_59_604 ();
 sg13g2_fill_1 FILLER_59_608 ();
 sg13g2_fill_2 FILLER_59_617 ();
 sg13g2_fill_1 FILLER_59_619 ();
 sg13g2_fill_1 FILLER_59_697 ();
 sg13g2_decap_8 FILLER_59_715 ();
 sg13g2_decap_8 FILLER_59_722 ();
 sg13g2_decap_8 FILLER_59_729 ();
 sg13g2_decap_4 FILLER_59_736 ();
 sg13g2_fill_2 FILLER_59_760 ();
 sg13g2_fill_1 FILLER_59_762 ();
 sg13g2_decap_8 FILLER_59_789 ();
 sg13g2_decap_8 FILLER_59_796 ();
 sg13g2_decap_8 FILLER_59_803 ();
 sg13g2_decap_8 FILLER_59_810 ();
 sg13g2_decap_8 FILLER_59_817 ();
 sg13g2_decap_8 FILLER_59_824 ();
 sg13g2_decap_8 FILLER_59_831 ();
 sg13g2_decap_8 FILLER_59_838 ();
 sg13g2_decap_8 FILLER_59_845 ();
 sg13g2_decap_8 FILLER_59_852 ();
 sg13g2_fill_2 FILLER_59_859 ();
 sg13g2_fill_1 FILLER_59_861 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_11 ();
 sg13g2_decap_4 FILLER_60_18 ();
 sg13g2_fill_1 FILLER_60_22 ();
 sg13g2_decap_4 FILLER_60_27 ();
 sg13g2_fill_1 FILLER_60_31 ();
 sg13g2_decap_8 FILLER_60_46 ();
 sg13g2_fill_1 FILLER_60_79 ();
 sg13g2_fill_1 FILLER_60_93 ();
 sg13g2_fill_1 FILLER_60_102 ();
 sg13g2_fill_1 FILLER_60_129 ();
 sg13g2_fill_1 FILLER_60_161 ();
 sg13g2_decap_8 FILLER_60_174 ();
 sg13g2_decap_4 FILLER_60_181 ();
 sg13g2_fill_1 FILLER_60_188 ();
 sg13g2_decap_8 FILLER_60_192 ();
 sg13g2_fill_2 FILLER_60_199 ();
 sg13g2_fill_1 FILLER_60_201 ();
 sg13g2_fill_2 FILLER_60_231 ();
 sg13g2_fill_2 FILLER_60_282 ();
 sg13g2_fill_2 FILLER_60_294 ();
 sg13g2_decap_4 FILLER_60_322 ();
 sg13g2_decap_4 FILLER_60_330 ();
 sg13g2_fill_2 FILLER_60_339 ();
 sg13g2_decap_4 FILLER_60_390 ();
 sg13g2_decap_8 FILLER_60_402 ();
 sg13g2_decap_8 FILLER_60_409 ();
 sg13g2_decap_8 FILLER_60_416 ();
 sg13g2_decap_8 FILLER_60_423 ();
 sg13g2_decap_8 FILLER_60_433 ();
 sg13g2_decap_8 FILLER_60_440 ();
 sg13g2_decap_8 FILLER_60_447 ();
 sg13g2_fill_2 FILLER_60_454 ();
 sg13g2_fill_2 FILLER_60_461 ();
 sg13g2_decap_8 FILLER_60_468 ();
 sg13g2_decap_8 FILLER_60_475 ();
 sg13g2_decap_8 FILLER_60_485 ();
 sg13g2_fill_2 FILLER_60_499 ();
 sg13g2_fill_1 FILLER_60_501 ();
 sg13g2_decap_8 FILLER_60_505 ();
 sg13g2_decap_8 FILLER_60_512 ();
 sg13g2_decap_4 FILLER_60_519 ();
 sg13g2_fill_1 FILLER_60_523 ();
 sg13g2_decap_8 FILLER_60_547 ();
 sg13g2_fill_2 FILLER_60_561 ();
 sg13g2_decap_8 FILLER_60_599 ();
 sg13g2_decap_4 FILLER_60_606 ();
 sg13g2_fill_2 FILLER_60_610 ();
 sg13g2_decap_8 FILLER_60_625 ();
 sg13g2_fill_2 FILLER_60_632 ();
 sg13g2_fill_1 FILLER_60_634 ();
 sg13g2_fill_1 FILLER_60_640 ();
 sg13g2_decap_8 FILLER_60_644 ();
 sg13g2_decap_8 FILLER_60_651 ();
 sg13g2_decap_8 FILLER_60_658 ();
 sg13g2_decap_8 FILLER_60_665 ();
 sg13g2_decap_4 FILLER_60_672 ();
 sg13g2_fill_1 FILLER_60_676 ();
 sg13g2_fill_1 FILLER_60_685 ();
 sg13g2_decap_4 FILLER_60_705 ();
 sg13g2_fill_2 FILLER_60_735 ();
 sg13g2_decap_4 FILLER_60_766 ();
 sg13g2_fill_1 FILLER_60_770 ();
 sg13g2_decap_8 FILLER_60_805 ();
 sg13g2_decap_8 FILLER_60_812 ();
 sg13g2_decap_8 FILLER_60_819 ();
 sg13g2_decap_8 FILLER_60_826 ();
 sg13g2_decap_8 FILLER_60_833 ();
 sg13g2_decap_8 FILLER_60_840 ();
 sg13g2_decap_8 FILLER_60_847 ();
 sg13g2_decap_8 FILLER_60_854 ();
 sg13g2_fill_1 FILLER_60_861 ();
 sg13g2_fill_1 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_27 ();
 sg13g2_decap_8 FILLER_61_52 ();
 sg13g2_fill_1 FILLER_61_59 ();
 sg13g2_fill_2 FILLER_61_86 ();
 sg13g2_fill_1 FILLER_61_88 ();
 sg13g2_decap_8 FILLER_61_103 ();
 sg13g2_fill_1 FILLER_61_110 ();
 sg13g2_fill_2 FILLER_61_116 ();
 sg13g2_fill_1 FILLER_61_118 ();
 sg13g2_decap_8 FILLER_61_124 ();
 sg13g2_fill_2 FILLER_61_131 ();
 sg13g2_fill_1 FILLER_61_133 ();
 sg13g2_decap_4 FILLER_61_140 ();
 sg13g2_decap_4 FILLER_61_152 ();
 sg13g2_fill_1 FILLER_61_156 ();
 sg13g2_fill_2 FILLER_61_175 ();
 sg13g2_fill_1 FILLER_61_177 ();
 sg13g2_decap_8 FILLER_61_204 ();
 sg13g2_decap_4 FILLER_61_211 ();
 sg13g2_fill_2 FILLER_61_215 ();
 sg13g2_decap_8 FILLER_61_250 ();
 sg13g2_fill_2 FILLER_61_257 ();
 sg13g2_decap_8 FILLER_61_267 ();
 sg13g2_decap_8 FILLER_61_274 ();
 sg13g2_fill_1 FILLER_61_281 ();
 sg13g2_decap_8 FILLER_61_292 ();
 sg13g2_decap_8 FILLER_61_299 ();
 sg13g2_fill_2 FILLER_61_349 ();
 sg13g2_decap_8 FILLER_61_364 ();
 sg13g2_fill_2 FILLER_61_371 ();
 sg13g2_fill_1 FILLER_61_373 ();
 sg13g2_decap_8 FILLER_61_420 ();
 sg13g2_decap_8 FILLER_61_427 ();
 sg13g2_fill_2 FILLER_61_437 ();
 sg13g2_decap_8 FILLER_61_447 ();
 sg13g2_decap_4 FILLER_61_454 ();
 sg13g2_fill_1 FILLER_61_458 ();
 sg13g2_fill_1 FILLER_61_467 ();
 sg13g2_fill_2 FILLER_61_488 ();
 sg13g2_fill_1 FILLER_61_490 ();
 sg13g2_fill_1 FILLER_61_537 ();
 sg13g2_decap_4 FILLER_61_571 ();
 sg13g2_fill_1 FILLER_61_575 ();
 sg13g2_decap_8 FILLER_61_579 ();
 sg13g2_fill_2 FILLER_61_597 ();
 sg13g2_decap_8 FILLER_61_602 ();
 sg13g2_decap_4 FILLER_61_609 ();
 sg13g2_fill_1 FILLER_61_613 ();
 sg13g2_decap_8 FILLER_61_640 ();
 sg13g2_fill_2 FILLER_61_647 ();
 sg13g2_fill_1 FILLER_61_686 ();
 sg13g2_fill_2 FILLER_61_695 ();
 sg13g2_decap_4 FILLER_61_723 ();
 sg13g2_fill_2 FILLER_61_727 ();
 sg13g2_fill_2 FILLER_61_759 ();
 sg13g2_decap_8 FILLER_61_787 ();
 sg13g2_decap_8 FILLER_61_794 ();
 sg13g2_decap_8 FILLER_61_801 ();
 sg13g2_decap_8 FILLER_61_808 ();
 sg13g2_decap_8 FILLER_61_815 ();
 sg13g2_decap_8 FILLER_61_822 ();
 sg13g2_decap_8 FILLER_61_829 ();
 sg13g2_decap_8 FILLER_61_836 ();
 sg13g2_decap_8 FILLER_61_843 ();
 sg13g2_decap_8 FILLER_61_850 ();
 sg13g2_decap_4 FILLER_61_857 ();
 sg13g2_fill_1 FILLER_61_861 ();
 sg13g2_fill_1 FILLER_62_0 ();
 sg13g2_decap_4 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_73 ();
 sg13g2_decap_8 FILLER_62_80 ();
 sg13g2_decap_4 FILLER_62_87 ();
 sg13g2_fill_1 FILLER_62_91 ();
 sg13g2_fill_2 FILLER_62_104 ();
 sg13g2_fill_2 FILLER_62_114 ();
 sg13g2_decap_4 FILLER_62_150 ();
 sg13g2_fill_2 FILLER_62_162 ();
 sg13g2_fill_1 FILLER_62_164 ();
 sg13g2_decap_8 FILLER_62_170 ();
 sg13g2_decap_8 FILLER_62_177 ();
 sg13g2_decap_8 FILLER_62_184 ();
 sg13g2_decap_4 FILLER_62_233 ();
 sg13g2_fill_2 FILLER_62_237 ();
 sg13g2_decap_8 FILLER_62_243 ();
 sg13g2_fill_1 FILLER_62_250 ();
 sg13g2_decap_8 FILLER_62_277 ();
 sg13g2_decap_4 FILLER_62_284 ();
 sg13g2_fill_1 FILLER_62_324 ();
 sg13g2_fill_1 FILLER_62_330 ();
 sg13g2_decap_4 FILLER_62_349 ();
 sg13g2_fill_2 FILLER_62_353 ();
 sg13g2_decap_8 FILLER_62_381 ();
 sg13g2_decap_8 FILLER_62_388 ();
 sg13g2_decap_4 FILLER_62_395 ();
 sg13g2_fill_2 FILLER_62_399 ();
 sg13g2_decap_8 FILLER_62_503 ();
 sg13g2_decap_8 FILLER_62_510 ();
 sg13g2_decap_8 FILLER_62_517 ();
 sg13g2_fill_2 FILLER_62_524 ();
 sg13g2_fill_1 FILLER_62_541 ();
 sg13g2_decap_4 FILLER_62_550 ();
 sg13g2_fill_1 FILLER_62_594 ();
 sg13g2_fill_1 FILLER_62_626 ();
 sg13g2_decap_8 FILLER_62_665 ();
 sg13g2_decap_4 FILLER_62_672 ();
 sg13g2_fill_2 FILLER_62_676 ();
 sg13g2_decap_8 FILLER_62_701 ();
 sg13g2_decap_4 FILLER_62_708 ();
 sg13g2_fill_1 FILLER_62_712 ();
 sg13g2_decap_8 FILLER_62_717 ();
 sg13g2_fill_2 FILLER_62_724 ();
 sg13g2_decap_4 FILLER_62_734 ();
 sg13g2_decap_4 FILLER_62_748 ();
 sg13g2_fill_2 FILLER_62_752 ();
 sg13g2_fill_2 FILLER_62_784 ();
 sg13g2_decap_8 FILLER_62_812 ();
 sg13g2_decap_8 FILLER_62_819 ();
 sg13g2_decap_8 FILLER_62_826 ();
 sg13g2_decap_8 FILLER_62_833 ();
 sg13g2_decap_8 FILLER_62_840 ();
 sg13g2_decap_8 FILLER_62_847 ();
 sg13g2_decap_8 FILLER_62_854 ();
 sg13g2_fill_1 FILLER_62_861 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_4 FILLER_63_28 ();
 sg13g2_fill_2 FILLER_63_32 ();
 sg13g2_decap_8 FILLER_63_39 ();
 sg13g2_fill_2 FILLER_63_92 ();
 sg13g2_fill_1 FILLER_63_100 ();
 sg13g2_fill_2 FILLER_63_115 ();
 sg13g2_fill_1 FILLER_63_117 ();
 sg13g2_decap_8 FILLER_63_123 ();
 sg13g2_decap_8 FILLER_63_130 ();
 sg13g2_fill_2 FILLER_63_137 ();
 sg13g2_decap_8 FILLER_63_144 ();
 sg13g2_fill_1 FILLER_63_151 ();
 sg13g2_fill_2 FILLER_63_178 ();
 sg13g2_fill_1 FILLER_63_180 ();
 sg13g2_fill_1 FILLER_63_190 ();
 sg13g2_decap_8 FILLER_63_235 ();
 sg13g2_decap_8 FILLER_63_242 ();
 sg13g2_decap_8 FILLER_63_249 ();
 sg13g2_fill_2 FILLER_63_256 ();
 sg13g2_decap_4 FILLER_63_266 ();
 sg13g2_fill_2 FILLER_63_270 ();
 sg13g2_fill_2 FILLER_63_293 ();
 sg13g2_fill_2 FILLER_63_300 ();
 sg13g2_fill_1 FILLER_63_302 ();
 sg13g2_decap_8 FILLER_63_306 ();
 sg13g2_decap_8 FILLER_63_313 ();
 sg13g2_decap_8 FILLER_63_320 ();
 sg13g2_decap_4 FILLER_63_327 ();
 sg13g2_fill_1 FILLER_63_331 ();
 sg13g2_decap_4 FILLER_63_399 ();
 sg13g2_fill_2 FILLER_63_403 ();
 sg13g2_decap_8 FILLER_63_424 ();
 sg13g2_decap_8 FILLER_63_431 ();
 sg13g2_decap_8 FILLER_63_438 ();
 sg13g2_decap_8 FILLER_63_445 ();
 sg13g2_decap_4 FILLER_63_452 ();
 sg13g2_fill_2 FILLER_63_456 ();
 sg13g2_decap_8 FILLER_63_466 ();
 sg13g2_fill_1 FILLER_63_473 ();
 sg13g2_decap_8 FILLER_63_479 ();
 sg13g2_decap_4 FILLER_63_486 ();
 sg13g2_fill_1 FILLER_63_490 ();
 sg13g2_decap_8 FILLER_63_505 ();
 sg13g2_decap_8 FILLER_63_512 ();
 sg13g2_fill_1 FILLER_63_519 ();
 sg13g2_decap_4 FILLER_63_564 ();
 sg13g2_fill_2 FILLER_63_568 ();
 sg13g2_decap_8 FILLER_63_573 ();
 sg13g2_decap_8 FILLER_63_580 ();
 sg13g2_fill_1 FILLER_63_587 ();
 sg13g2_decap_8 FILLER_63_599 ();
 sg13g2_fill_1 FILLER_63_606 ();
 sg13g2_fill_2 FILLER_63_615 ();
 sg13g2_fill_2 FILLER_63_621 ();
 sg13g2_fill_1 FILLER_63_623 ();
 sg13g2_fill_2 FILLER_63_637 ();
 sg13g2_decap_8 FILLER_63_644 ();
 sg13g2_fill_1 FILLER_63_651 ();
 sg13g2_fill_2 FILLER_63_657 ();
 sg13g2_decap_8 FILLER_63_671 ();
 sg13g2_decap_8 FILLER_63_678 ();
 sg13g2_fill_2 FILLER_63_685 ();
 sg13g2_fill_1 FILLER_63_693 ();
 sg13g2_fill_2 FILLER_63_702 ();
 sg13g2_decap_8 FILLER_63_743 ();
 sg13g2_fill_1 FILLER_63_750 ();
 sg13g2_decap_4 FILLER_63_760 ();
 sg13g2_fill_1 FILLER_63_764 ();
 sg13g2_fill_2 FILLER_63_773 ();
 sg13g2_fill_1 FILLER_63_775 ();
 sg13g2_decap_8 FILLER_63_792 ();
 sg13g2_decap_8 FILLER_63_799 ();
 sg13g2_decap_8 FILLER_63_806 ();
 sg13g2_decap_8 FILLER_63_813 ();
 sg13g2_decap_8 FILLER_63_820 ();
 sg13g2_decap_8 FILLER_63_827 ();
 sg13g2_decap_8 FILLER_63_834 ();
 sg13g2_decap_8 FILLER_63_841 ();
 sg13g2_decap_8 FILLER_63_848 ();
 sg13g2_decap_8 FILLER_63_855 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_4 FILLER_64_21 ();
 sg13g2_fill_2 FILLER_64_25 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_4 FILLER_64_84 ();
 sg13g2_fill_1 FILLER_64_88 ();
 sg13g2_fill_2 FILLER_64_106 ();
 sg13g2_fill_2 FILLER_64_129 ();
 sg13g2_fill_1 FILLER_64_131 ();
 sg13g2_decap_4 FILLER_64_158 ();
 sg13g2_fill_1 FILLER_64_162 ();
 sg13g2_fill_2 FILLER_64_186 ();
 sg13g2_decap_8 FILLER_64_200 ();
 sg13g2_decap_8 FILLER_64_207 ();
 sg13g2_decap_4 FILLER_64_214 ();
 sg13g2_fill_1 FILLER_64_218 ();
 sg13g2_fill_2 FILLER_64_289 ();
 sg13g2_decap_4 FILLER_64_333 ();
 sg13g2_decap_8 FILLER_64_345 ();
 sg13g2_decap_8 FILLER_64_352 ();
 sg13g2_decap_8 FILLER_64_359 ();
 sg13g2_decap_8 FILLER_64_366 ();
 sg13g2_decap_8 FILLER_64_373 ();
 sg13g2_decap_8 FILLER_64_380 ();
 sg13g2_fill_2 FILLER_64_416 ();
 sg13g2_decap_8 FILLER_64_444 ();
 sg13g2_fill_1 FILLER_64_451 ();
 sg13g2_decap_8 FILLER_64_543 ();
 sg13g2_decap_8 FILLER_64_550 ();
 sg13g2_decap_8 FILLER_64_557 ();
 sg13g2_fill_2 FILLER_64_564 ();
 sg13g2_decap_8 FILLER_64_582 ();
 sg13g2_decap_8 FILLER_64_589 ();
 sg13g2_decap_4 FILLER_64_596 ();
 sg13g2_fill_1 FILLER_64_600 ();
 sg13g2_fill_2 FILLER_64_639 ();
 sg13g2_fill_2 FILLER_64_646 ();
 sg13g2_fill_1 FILLER_64_648 ();
 sg13g2_fill_1 FILLER_64_657 ();
 sg13g2_decap_4 FILLER_64_676 ();
 sg13g2_fill_2 FILLER_64_687 ();
 sg13g2_fill_1 FILLER_64_689 ();
 sg13g2_fill_1 FILLER_64_698 ();
 sg13g2_decap_8 FILLER_64_720 ();
 sg13g2_decap_8 FILLER_64_727 ();
 sg13g2_decap_8 FILLER_64_734 ();
 sg13g2_fill_2 FILLER_64_741 ();
 sg13g2_fill_1 FILLER_64_743 ();
 sg13g2_fill_2 FILLER_64_770 ();
 sg13g2_fill_2 FILLER_64_784 ();
 sg13g2_decap_8 FILLER_64_812 ();
 sg13g2_decap_8 FILLER_64_819 ();
 sg13g2_decap_8 FILLER_64_826 ();
 sg13g2_decap_8 FILLER_64_833 ();
 sg13g2_decap_8 FILLER_64_840 ();
 sg13g2_decap_8 FILLER_64_847 ();
 sg13g2_decap_8 FILLER_64_854 ();
 sg13g2_fill_1 FILLER_64_861 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_fill_2 FILLER_65_21 ();
 sg13g2_fill_1 FILLER_65_23 ();
 sg13g2_fill_1 FILLER_65_32 ();
 sg13g2_fill_2 FILLER_65_54 ();
 sg13g2_fill_1 FILLER_65_56 ();
 sg13g2_decap_4 FILLER_65_83 ();
 sg13g2_fill_2 FILLER_65_87 ();
 sg13g2_fill_2 FILLER_65_124 ();
 sg13g2_decap_8 FILLER_65_157 ();
 sg13g2_fill_2 FILLER_65_164 ();
 sg13g2_fill_1 FILLER_65_166 ();
 sg13g2_fill_2 FILLER_65_180 ();
 sg13g2_fill_2 FILLER_65_195 ();
 sg13g2_decap_8 FILLER_65_223 ();
 sg13g2_decap_8 FILLER_65_230 ();
 sg13g2_decap_8 FILLER_65_237 ();
 sg13g2_fill_1 FILLER_65_272 ();
 sg13g2_decap_4 FILLER_65_288 ();
 sg13g2_decap_8 FILLER_65_296 ();
 sg13g2_decap_4 FILLER_65_303 ();
 sg13g2_fill_2 FILLER_65_307 ();
 sg13g2_decap_8 FILLER_65_319 ();
 sg13g2_decap_8 FILLER_65_326 ();
 sg13g2_decap_4 FILLER_65_333 ();
 sg13g2_decap_4 FILLER_65_363 ();
 sg13g2_fill_2 FILLER_65_367 ();
 sg13g2_decap_8 FILLER_65_395 ();
 sg13g2_fill_1 FILLER_65_402 ();
 sg13g2_decap_4 FILLER_65_425 ();
 sg13g2_fill_1 FILLER_65_429 ();
 sg13g2_decap_4 FILLER_65_469 ();
 sg13g2_fill_1 FILLER_65_473 ();
 sg13g2_fill_2 FILLER_65_477 ();
 sg13g2_decap_4 FILLER_65_484 ();
 sg13g2_fill_2 FILLER_65_488 ();
 sg13g2_decap_8 FILLER_65_493 ();
 sg13g2_fill_2 FILLER_65_500 ();
 sg13g2_fill_1 FILLER_65_502 ();
 sg13g2_decap_8 FILLER_65_513 ();
 sg13g2_decap_8 FILLER_65_520 ();
 sg13g2_fill_1 FILLER_65_527 ();
 sg13g2_decap_4 FILLER_65_551 ();
 sg13g2_fill_1 FILLER_65_555 ();
 sg13g2_fill_2 FILLER_65_601 ();
 sg13g2_fill_1 FILLER_65_603 ();
 sg13g2_fill_2 FILLER_65_609 ();
 sg13g2_decap_8 FILLER_65_616 ();
 sg13g2_decap_8 FILLER_65_623 ();
 sg13g2_decap_8 FILLER_65_630 ();
 sg13g2_decap_4 FILLER_65_637 ();
 sg13g2_fill_1 FILLER_65_641 ();
 sg13g2_decap_4 FILLER_65_646 ();
 sg13g2_fill_2 FILLER_65_650 ();
 sg13g2_decap_4 FILLER_65_678 ();
 sg13g2_fill_1 FILLER_65_682 ();
 sg13g2_decap_8 FILLER_65_692 ();
 sg13g2_fill_2 FILLER_65_699 ();
 sg13g2_fill_2 FILLER_65_709 ();
 sg13g2_decap_8 FILLER_65_737 ();
 sg13g2_decap_8 FILLER_65_744 ();
 sg13g2_fill_2 FILLER_65_751 ();
 sg13g2_fill_2 FILLER_65_770 ();
 sg13g2_fill_2 FILLER_65_780 ();
 sg13g2_fill_1 FILLER_65_782 ();
 sg13g2_decap_8 FILLER_65_809 ();
 sg13g2_decap_8 FILLER_65_816 ();
 sg13g2_decap_8 FILLER_65_823 ();
 sg13g2_decap_8 FILLER_65_830 ();
 sg13g2_decap_8 FILLER_65_837 ();
 sg13g2_decap_8 FILLER_65_844 ();
 sg13g2_decap_8 FILLER_65_851 ();
 sg13g2_decap_4 FILLER_65_858 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_4 FILLER_66_14 ();
 sg13g2_fill_2 FILLER_66_18 ();
 sg13g2_fill_1 FILLER_66_34 ();
 sg13g2_fill_2 FILLER_66_45 ();
 sg13g2_fill_1 FILLER_66_73 ();
 sg13g2_decap_8 FILLER_66_79 ();
 sg13g2_decap_8 FILLER_66_86 ();
 sg13g2_fill_2 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_110 ();
 sg13g2_decap_8 FILLER_66_117 ();
 sg13g2_decap_8 FILLER_66_124 ();
 sg13g2_decap_8 FILLER_66_131 ();
 sg13g2_decap_8 FILLER_66_138 ();
 sg13g2_fill_1 FILLER_66_145 ();
 sg13g2_decap_4 FILLER_66_154 ();
 sg13g2_fill_1 FILLER_66_158 ();
 sg13g2_fill_2 FILLER_66_180 ();
 sg13g2_fill_1 FILLER_66_182 ();
 sg13g2_fill_1 FILLER_66_209 ();
 sg13g2_decap_8 FILLER_66_241 ();
 sg13g2_fill_2 FILLER_66_265 ();
 sg13g2_decap_8 FILLER_66_271 ();
 sg13g2_decap_8 FILLER_66_278 ();
 sg13g2_decap_4 FILLER_66_311 ();
 sg13g2_fill_1 FILLER_66_315 ();
 sg13g2_fill_1 FILLER_66_342 ();
 sg13g2_fill_2 FILLER_66_352 ();
 sg13g2_fill_1 FILLER_66_354 ();
 sg13g2_fill_2 FILLER_66_383 ();
 sg13g2_decap_8 FILLER_66_411 ();
 sg13g2_fill_2 FILLER_66_418 ();
 sg13g2_fill_1 FILLER_66_420 ();
 sg13g2_decap_8 FILLER_66_443 ();
 sg13g2_fill_1 FILLER_66_450 ();
 sg13g2_fill_2 FILLER_66_482 ();
 sg13g2_decap_8 FILLER_66_531 ();
 sg13g2_fill_2 FILLER_66_564 ();
 sg13g2_decap_8 FILLER_66_587 ();
 sg13g2_decap_4 FILLER_66_594 ();
 sg13g2_fill_1 FILLER_66_598 ();
 sg13g2_decap_4 FILLER_66_604 ();
 sg13g2_fill_2 FILLER_66_660 ();
 sg13g2_fill_1 FILLER_66_662 ();
 sg13g2_decap_4 FILLER_66_689 ();
 sg13g2_fill_1 FILLER_66_693 ();
 sg13g2_decap_8 FILLER_66_707 ();
 sg13g2_decap_8 FILLER_66_714 ();
 sg13g2_decap_8 FILLER_66_721 ();
 sg13g2_fill_1 FILLER_66_728 ();
 sg13g2_decap_8 FILLER_66_737 ();
 sg13g2_decap_8 FILLER_66_744 ();
 sg13g2_fill_2 FILLER_66_751 ();
 sg13g2_fill_2 FILLER_66_761 ();
 sg13g2_fill_1 FILLER_66_763 ();
 sg13g2_decap_8 FILLER_66_798 ();
 sg13g2_decap_8 FILLER_66_805 ();
 sg13g2_decap_8 FILLER_66_812 ();
 sg13g2_decap_8 FILLER_66_819 ();
 sg13g2_decap_8 FILLER_66_826 ();
 sg13g2_decap_8 FILLER_66_833 ();
 sg13g2_decap_8 FILLER_66_840 ();
 sg13g2_decap_8 FILLER_66_847 ();
 sg13g2_decap_8 FILLER_66_854 ();
 sg13g2_fill_1 FILLER_66_861 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_4 FILLER_67_21 ();
 sg13g2_fill_1 FILLER_67_25 ();
 sg13g2_fill_2 FILLER_67_34 ();
 sg13g2_fill_2 FILLER_67_75 ();
 sg13g2_fill_1 FILLER_67_105 ();
 sg13g2_decap_4 FILLER_67_132 ();
 sg13g2_fill_2 FILLER_67_136 ();
 sg13g2_fill_1 FILLER_67_155 ();
 sg13g2_decap_8 FILLER_67_184 ();
 sg13g2_decap_8 FILLER_67_191 ();
 sg13g2_decap_8 FILLER_67_198 ();
 sg13g2_decap_8 FILLER_67_205 ();
 sg13g2_decap_8 FILLER_67_217 ();
 sg13g2_decap_4 FILLER_67_224 ();
 sg13g2_fill_1 FILLER_67_228 ();
 sg13g2_fill_2 FILLER_67_242 ();
 sg13g2_fill_1 FILLER_67_244 ();
 sg13g2_decap_8 FILLER_67_272 ();
 sg13g2_decap_8 FILLER_67_279 ();
 sg13g2_decap_8 FILLER_67_322 ();
 sg13g2_decap_8 FILLER_67_339 ();
 sg13g2_decap_4 FILLER_67_346 ();
 sg13g2_decap_8 FILLER_67_394 ();
 sg13g2_fill_2 FILLER_67_427 ();
 sg13g2_fill_2 FILLER_67_458 ();
 sg13g2_decap_8 FILLER_67_465 ();
 sg13g2_decap_8 FILLER_67_472 ();
 sg13g2_decap_8 FILLER_67_479 ();
 sg13g2_fill_1 FILLER_67_486 ();
 sg13g2_fill_2 FILLER_67_495 ();
 sg13g2_decap_8 FILLER_67_515 ();
 sg13g2_decap_8 FILLER_67_522 ();
 sg13g2_fill_2 FILLER_67_529 ();
 sg13g2_fill_1 FILLER_67_531 ();
 sg13g2_decap_8 FILLER_67_556 ();
 sg13g2_decap_8 FILLER_67_563 ();
 sg13g2_fill_1 FILLER_67_596 ();
 sg13g2_decap_8 FILLER_67_615 ();
 sg13g2_decap_8 FILLER_67_622 ();
 sg13g2_decap_4 FILLER_67_629 ();
 sg13g2_fill_1 FILLER_67_633 ();
 sg13g2_decap_4 FILLER_67_639 ();
 sg13g2_decap_8 FILLER_67_675 ();
 sg13g2_decap_4 FILLER_67_682 ();
 sg13g2_fill_2 FILLER_67_772 ();
 sg13g2_fill_1 FILLER_67_774 ();
 sg13g2_decap_4 FILLER_67_781 ();
 sg13g2_decap_8 FILLER_67_815 ();
 sg13g2_decap_8 FILLER_67_822 ();
 sg13g2_decap_8 FILLER_67_829 ();
 sg13g2_decap_8 FILLER_67_836 ();
 sg13g2_decap_8 FILLER_67_843 ();
 sg13g2_decap_8 FILLER_67_850 ();
 sg13g2_decap_4 FILLER_67_857 ();
 sg13g2_fill_1 FILLER_67_861 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_fill_1 FILLER_68_28 ();
 sg13g2_fill_1 FILLER_68_34 ();
 sg13g2_decap_8 FILLER_68_48 ();
 sg13g2_decap_8 FILLER_68_55 ();
 sg13g2_decap_8 FILLER_68_62 ();
 sg13g2_decap_8 FILLER_68_69 ();
 sg13g2_fill_2 FILLER_68_76 ();
 sg13g2_fill_1 FILLER_68_78 ();
 sg13g2_decap_4 FILLER_68_102 ();
 sg13g2_fill_2 FILLER_68_132 ();
 sg13g2_fill_1 FILLER_68_134 ();
 sg13g2_fill_2 FILLER_68_147 ();
 sg13g2_decap_8 FILLER_68_154 ();
 sg13g2_decap_4 FILLER_68_161 ();
 sg13g2_decap_4 FILLER_68_185 ();
 sg13g2_fill_1 FILLER_68_189 ();
 sg13g2_decap_8 FILLER_68_216 ();
 sg13g2_decap_8 FILLER_68_223 ();
 sg13g2_fill_2 FILLER_68_238 ();
 sg13g2_fill_1 FILLER_68_240 ();
 sg13g2_decap_4 FILLER_68_249 ();
 sg13g2_fill_2 FILLER_68_258 ();
 sg13g2_decap_8 FILLER_68_282 ();
 sg13g2_decap_8 FILLER_68_289 ();
 sg13g2_decap_8 FILLER_68_296 ();
 sg13g2_decap_8 FILLER_68_303 ();
 sg13g2_fill_2 FILLER_68_310 ();
 sg13g2_fill_2 FILLER_68_348 ();
 sg13g2_decap_8 FILLER_68_358 ();
 sg13g2_decap_4 FILLER_68_365 ();
 sg13g2_decap_8 FILLER_68_374 ();
 sg13g2_decap_8 FILLER_68_381 ();
 sg13g2_fill_2 FILLER_68_388 ();
 sg13g2_fill_1 FILLER_68_390 ();
 sg13g2_decap_8 FILLER_68_406 ();
 sg13g2_decap_8 FILLER_68_413 ();
 sg13g2_decap_8 FILLER_68_420 ();
 sg13g2_decap_4 FILLER_68_427 ();
 sg13g2_fill_1 FILLER_68_431 ();
 sg13g2_decap_8 FILLER_68_447 ();
 sg13g2_decap_8 FILLER_68_454 ();
 sg13g2_decap_4 FILLER_68_461 ();
 sg13g2_fill_1 FILLER_68_465 ();
 sg13g2_fill_1 FILLER_68_505 ();
 sg13g2_fill_2 FILLER_68_537 ();
 sg13g2_decap_8 FILLER_68_571 ();
 sg13g2_fill_2 FILLER_68_578 ();
 sg13g2_fill_1 FILLER_68_598 ();
 sg13g2_decap_4 FILLER_68_617 ();
 sg13g2_decap_4 FILLER_68_641 ();
 sg13g2_fill_1 FILLER_68_645 ();
 sg13g2_fill_2 FILLER_68_658 ();
 sg13g2_decap_8 FILLER_68_668 ();
 sg13g2_decap_8 FILLER_68_675 ();
 sg13g2_decap_8 FILLER_68_682 ();
 sg13g2_fill_2 FILLER_68_689 ();
 sg13g2_fill_1 FILLER_68_691 ();
 sg13g2_fill_1 FILLER_68_701 ();
 sg13g2_decap_8 FILLER_68_736 ();
 sg13g2_fill_1 FILLER_68_748 ();
 sg13g2_decap_8 FILLER_68_762 ();
 sg13g2_decap_4 FILLER_68_769 ();
 sg13g2_fill_1 FILLER_68_773 ();
 sg13g2_fill_1 FILLER_68_778 ();
 sg13g2_fill_2 FILLER_68_787 ();
 sg13g2_decap_8 FILLER_68_797 ();
 sg13g2_decap_8 FILLER_68_804 ();
 sg13g2_decap_8 FILLER_68_811 ();
 sg13g2_decap_8 FILLER_68_818 ();
 sg13g2_decap_8 FILLER_68_825 ();
 sg13g2_decap_8 FILLER_68_832 ();
 sg13g2_decap_8 FILLER_68_839 ();
 sg13g2_decap_8 FILLER_68_846 ();
 sg13g2_decap_8 FILLER_68_853 ();
 sg13g2_fill_2 FILLER_68_860 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_4 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_72 ();
 sg13g2_fill_2 FILLER_69_79 ();
 sg13g2_fill_1 FILLER_69_81 ();
 sg13g2_fill_1 FILLER_69_95 ();
 sg13g2_decap_8 FILLER_69_109 ();
 sg13g2_fill_2 FILLER_69_116 ();
 sg13g2_fill_1 FILLER_69_118 ();
 sg13g2_fill_2 FILLER_69_135 ();
 sg13g2_decap_8 FILLER_69_158 ();
 sg13g2_fill_2 FILLER_69_175 ();
 sg13g2_decap_4 FILLER_69_181 ();
 sg13g2_fill_1 FILLER_69_237 ();
 sg13g2_fill_2 FILLER_69_251 ();
 sg13g2_fill_1 FILLER_69_253 ();
 sg13g2_decap_4 FILLER_69_285 ();
 sg13g2_fill_1 FILLER_69_289 ();
 sg13g2_decap_4 FILLER_69_326 ();
 sg13g2_fill_2 FILLER_69_330 ();
 sg13g2_decap_8 FILLER_69_358 ();
 sg13g2_fill_2 FILLER_69_373 ();
 sg13g2_fill_1 FILLER_69_427 ();
 sg13g2_fill_1 FILLER_69_436 ();
 sg13g2_decap_8 FILLER_69_471 ();
 sg13g2_decap_8 FILLER_69_478 ();
 sg13g2_decap_4 FILLER_69_485 ();
 sg13g2_fill_2 FILLER_69_489 ();
 sg13g2_decap_8 FILLER_69_513 ();
 sg13g2_decap_8 FILLER_69_520 ();
 sg13g2_decap_8 FILLER_69_527 ();
 sg13g2_decap_4 FILLER_69_555 ();
 sg13g2_fill_1 FILLER_69_559 ();
 sg13g2_decap_8 FILLER_69_586 ();
 sg13g2_decap_8 FILLER_69_632 ();
 sg13g2_decap_4 FILLER_69_639 ();
 sg13g2_fill_2 FILLER_69_643 ();
 sg13g2_fill_2 FILLER_69_653 ();
 sg13g2_fill_1 FILLER_69_655 ();
 sg13g2_decap_4 FILLER_69_690 ();
 sg13g2_fill_2 FILLER_69_712 ();
 sg13g2_fill_1 FILLER_69_714 ();
 sg13g2_decap_4 FILLER_69_719 ();
 sg13g2_decap_8 FILLER_69_731 ();
 sg13g2_fill_2 FILLER_69_738 ();
 sg13g2_fill_1 FILLER_69_784 ();
 sg13g2_decap_8 FILLER_69_811 ();
 sg13g2_decap_8 FILLER_69_818 ();
 sg13g2_decap_8 FILLER_69_825 ();
 sg13g2_decap_8 FILLER_69_832 ();
 sg13g2_decap_8 FILLER_69_839 ();
 sg13g2_decap_8 FILLER_69_846 ();
 sg13g2_decap_8 FILLER_69_853 ();
 sg13g2_fill_2 FILLER_69_860 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_4 FILLER_70_28 ();
 sg13g2_fill_2 FILLER_70_32 ();
 sg13g2_decap_4 FILLER_70_38 ();
 sg13g2_decap_4 FILLER_70_68 ();
 sg13g2_fill_2 FILLER_70_103 ();
 sg13g2_fill_2 FILLER_70_113 ();
 sg13g2_decap_8 FILLER_70_141 ();
 sg13g2_fill_2 FILLER_70_173 ();
 sg13g2_fill_1 FILLER_70_175 ();
 sg13g2_fill_1 FILLER_70_184 ();
 sg13g2_decap_8 FILLER_70_211 ();
 sg13g2_fill_2 FILLER_70_218 ();
 sg13g2_decap_4 FILLER_70_228 ();
 sg13g2_fill_2 FILLER_70_232 ();
 sg13g2_decap_8 FILLER_70_238 ();
 sg13g2_fill_2 FILLER_70_245 ();
 sg13g2_fill_1 FILLER_70_247 ();
 sg13g2_decap_8 FILLER_70_252 ();
 sg13g2_fill_2 FILLER_70_272 ();
 sg13g2_fill_1 FILLER_70_278 ();
 sg13g2_fill_2 FILLER_70_305 ();
 sg13g2_decap_4 FILLER_70_343 ();
 sg13g2_fill_1 FILLER_70_373 ();
 sg13g2_decap_8 FILLER_70_379 ();
 sg13g2_decap_8 FILLER_70_406 ();
 sg13g2_decap_8 FILLER_70_413 ();
 sg13g2_decap_4 FILLER_70_420 ();
 sg13g2_decap_4 FILLER_70_458 ();
 sg13g2_fill_2 FILLER_70_462 ();
 sg13g2_fill_1 FILLER_70_472 ();
 sg13g2_decap_4 FILLER_70_499 ();
 sg13g2_fill_2 FILLER_70_503 ();
 sg13g2_decap_4 FILLER_70_521 ();
 sg13g2_decap_4 FILLER_70_533 ();
 sg13g2_decap_8 FILLER_70_563 ();
 sg13g2_decap_4 FILLER_70_591 ();
 sg13g2_fill_2 FILLER_70_595 ();
 sg13g2_decap_8 FILLER_70_601 ();
 sg13g2_decap_4 FILLER_70_608 ();
 sg13g2_decap_8 FILLER_70_617 ();
 sg13g2_decap_4 FILLER_70_624 ();
 sg13g2_fill_1 FILLER_70_628 ();
 sg13g2_fill_1 FILLER_70_655 ();
 sg13g2_fill_2 FILLER_70_670 ();
 sg13g2_fill_2 FILLER_70_677 ();
 sg13g2_fill_1 FILLER_70_679 ();
 sg13g2_fill_2 FILLER_70_694 ();
 sg13g2_fill_1 FILLER_70_696 ();
 sg13g2_fill_2 FILLER_70_707 ();
 sg13g2_fill_2 FILLER_70_715 ();
 sg13g2_fill_1 FILLER_70_717 ();
 sg13g2_decap_8 FILLER_70_736 ();
 sg13g2_decap_8 FILLER_70_743 ();
 sg13g2_fill_2 FILLER_70_750 ();
 sg13g2_fill_2 FILLER_70_760 ();
 sg13g2_fill_2 FILLER_70_769 ();
 sg13g2_fill_1 FILLER_70_771 ();
 sg13g2_fill_2 FILLER_70_777 ();
 sg13g2_decap_8 FILLER_70_793 ();
 sg13g2_decap_8 FILLER_70_800 ();
 sg13g2_decap_8 FILLER_70_807 ();
 sg13g2_decap_8 FILLER_70_814 ();
 sg13g2_decap_8 FILLER_70_821 ();
 sg13g2_decap_8 FILLER_70_828 ();
 sg13g2_decap_8 FILLER_70_835 ();
 sg13g2_decap_8 FILLER_70_842 ();
 sg13g2_decap_8 FILLER_70_849 ();
 sg13g2_decap_4 FILLER_70_856 ();
 sg13g2_fill_2 FILLER_70_860 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_4 FILLER_71_42 ();
 sg13g2_decap_4 FILLER_71_54 ();
 sg13g2_fill_1 FILLER_71_58 ();
 sg13g2_decap_8 FILLER_71_114 ();
 sg13g2_decap_8 FILLER_71_121 ();
 sg13g2_fill_2 FILLER_71_128 ();
 sg13g2_decap_8 FILLER_71_138 ();
 sg13g2_decap_8 FILLER_71_145 ();
 sg13g2_decap_4 FILLER_71_152 ();
 sg13g2_fill_1 FILLER_71_156 ();
 sg13g2_fill_1 FILLER_71_170 ();
 sg13g2_decap_8 FILLER_71_176 ();
 sg13g2_decap_8 FILLER_71_183 ();
 sg13g2_decap_8 FILLER_71_190 ();
 sg13g2_decap_8 FILLER_71_197 ();
 sg13g2_decap_8 FILLER_71_204 ();
 sg13g2_fill_2 FILLER_71_211 ();
 sg13g2_decap_4 FILLER_71_247 ();
 sg13g2_fill_2 FILLER_71_251 ();
 sg13g2_decap_8 FILLER_71_270 ();
 sg13g2_fill_2 FILLER_71_277 ();
 sg13g2_decap_8 FILLER_71_305 ();
 sg13g2_fill_2 FILLER_71_312 ();
 sg13g2_decap_4 FILLER_71_322 ();
 sg13g2_fill_1 FILLER_71_326 ();
 sg13g2_decap_4 FILLER_71_335 ();
 sg13g2_fill_2 FILLER_71_339 ();
 sg13g2_decap_8 FILLER_71_361 ();
 sg13g2_decap_4 FILLER_71_368 ();
 sg13g2_fill_1 FILLER_71_372 ();
 sg13g2_decap_8 FILLER_71_409 ();
 sg13g2_fill_2 FILLER_71_416 ();
 sg13g2_fill_1 FILLER_71_418 ();
 sg13g2_decap_4 FILLER_71_424 ();
 sg13g2_fill_2 FILLER_71_433 ();
 sg13g2_decap_8 FILLER_71_440 ();
 sg13g2_decap_8 FILLER_71_447 ();
 sg13g2_decap_4 FILLER_71_454 ();
 sg13g2_fill_2 FILLER_71_458 ();
 sg13g2_fill_1 FILLER_71_468 ();
 sg13g2_decap_4 FILLER_71_489 ();
 sg13g2_fill_1 FILLER_71_497 ();
 sg13g2_fill_2 FILLER_71_524 ();
 sg13g2_fill_1 FILLER_71_526 ();
 sg13g2_decap_8 FILLER_71_540 ();
 sg13g2_fill_1 FILLER_71_547 ();
 sg13g2_decap_8 FILLER_71_552 ();
 sg13g2_fill_2 FILLER_71_567 ();
 sg13g2_fill_1 FILLER_71_569 ();
 sg13g2_fill_2 FILLER_71_584 ();
 sg13g2_fill_2 FILLER_71_602 ();
 sg13g2_decap_4 FILLER_71_609 ();
 sg13g2_fill_2 FILLER_71_626 ();
 sg13g2_fill_1 FILLER_71_628 ();
 sg13g2_decap_4 FILLER_71_645 ();
 sg13g2_fill_2 FILLER_71_649 ();
 sg13g2_fill_2 FILLER_71_663 ();
 sg13g2_fill_1 FILLER_71_665 ();
 sg13g2_fill_1 FILLER_71_676 ();
 sg13g2_fill_2 FILLER_71_705 ();
 sg13g2_fill_2 FILLER_71_720 ();
 sg13g2_fill_1 FILLER_71_722 ();
 sg13g2_decap_8 FILLER_71_727 ();
 sg13g2_decap_8 FILLER_71_734 ();
 sg13g2_fill_1 FILLER_71_775 ();
 sg13g2_decap_8 FILLER_71_787 ();
 sg13g2_decap_8 FILLER_71_794 ();
 sg13g2_decap_8 FILLER_71_801 ();
 sg13g2_decap_8 FILLER_71_808 ();
 sg13g2_decap_8 FILLER_71_815 ();
 sg13g2_decap_8 FILLER_71_822 ();
 sg13g2_decap_8 FILLER_71_829 ();
 sg13g2_decap_8 FILLER_71_836 ();
 sg13g2_decap_8 FILLER_71_843 ();
 sg13g2_decap_8 FILLER_71_850 ();
 sg13g2_decap_4 FILLER_71_857 ();
 sg13g2_fill_1 FILLER_71_861 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_4 FILLER_72_35 ();
 sg13g2_decap_4 FILLER_72_85 ();
 sg13g2_fill_2 FILLER_72_89 ();
 sg13g2_fill_2 FILLER_72_116 ();
 sg13g2_fill_2 FILLER_72_144 ();
 sg13g2_fill_1 FILLER_72_158 ();
 sg13g2_fill_2 FILLER_72_167 ();
 sg13g2_fill_2 FILLER_72_177 ();
 sg13g2_fill_1 FILLER_72_179 ();
 sg13g2_fill_2 FILLER_72_247 ();
 sg13g2_fill_1 FILLER_72_249 ();
 sg13g2_decap_4 FILLER_72_275 ();
 sg13g2_decap_8 FILLER_72_305 ();
 sg13g2_decap_4 FILLER_72_312 ();
 sg13g2_fill_1 FILLER_72_326 ();
 sg13g2_fill_2 FILLER_72_353 ();
 sg13g2_fill_1 FILLER_72_355 ();
 sg13g2_decap_8 FILLER_72_382 ();
 sg13g2_decap_8 FILLER_72_389 ();
 sg13g2_fill_2 FILLER_72_396 ();
 sg13g2_fill_1 FILLER_72_398 ();
 sg13g2_fill_2 FILLER_72_425 ();
 sg13g2_decap_8 FILLER_72_440 ();
 sg13g2_fill_2 FILLER_72_447 ();
 sg13g2_fill_1 FILLER_72_449 ();
 sg13g2_decap_8 FILLER_72_482 ();
 sg13g2_decap_8 FILLER_72_489 ();
 sg13g2_decap_8 FILLER_72_496 ();
 sg13g2_fill_2 FILLER_72_503 ();
 sg13g2_fill_1 FILLER_72_513 ();
 sg13g2_decap_8 FILLER_72_528 ();
 sg13g2_decap_4 FILLER_72_535 ();
 sg13g2_fill_1 FILLER_72_539 ();
 sg13g2_decap_8 FILLER_72_566 ();
 sg13g2_fill_1 FILLER_72_573 ();
 sg13g2_fill_2 FILLER_72_587 ();
 sg13g2_fill_1 FILLER_72_603 ();
 sg13g2_fill_2 FILLER_72_612 ();
 sg13g2_fill_1 FILLER_72_614 ();
 sg13g2_decap_4 FILLER_72_627 ();
 sg13g2_fill_1 FILLER_72_631 ();
 sg13g2_decap_4 FILLER_72_637 ();
 sg13g2_fill_1 FILLER_72_641 ();
 sg13g2_decap_8 FILLER_72_652 ();
 sg13g2_decap_4 FILLER_72_659 ();
 sg13g2_fill_1 FILLER_72_663 ();
 sg13g2_decap_4 FILLER_72_684 ();
 sg13g2_fill_2 FILLER_72_688 ();
 sg13g2_fill_1 FILLER_72_698 ();
 sg13g2_fill_2 FILLER_72_768 ();
 sg13g2_decap_8 FILLER_72_809 ();
 sg13g2_decap_8 FILLER_72_816 ();
 sg13g2_decap_8 FILLER_72_823 ();
 sg13g2_decap_8 FILLER_72_830 ();
 sg13g2_decap_8 FILLER_72_837 ();
 sg13g2_decap_8 FILLER_72_844 ();
 sg13g2_decap_8 FILLER_72_851 ();
 sg13g2_decap_4 FILLER_72_858 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_4 FILLER_73_42 ();
 sg13g2_fill_2 FILLER_73_46 ();
 sg13g2_decap_8 FILLER_73_57 ();
 sg13g2_decap_8 FILLER_73_64 ();
 sg13g2_decap_8 FILLER_73_71 ();
 sg13g2_decap_8 FILLER_73_78 ();
 sg13g2_decap_8 FILLER_73_85 ();
 sg13g2_decap_4 FILLER_73_92 ();
 sg13g2_fill_1 FILLER_73_96 ();
 sg13g2_fill_1 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_121 ();
 sg13g2_decap_8 FILLER_73_128 ();
 sg13g2_decap_8 FILLER_73_135 ();
 sg13g2_fill_2 FILLER_73_142 ();
 sg13g2_fill_2 FILLER_73_152 ();
 sg13g2_fill_2 FILLER_73_180 ();
 sg13g2_fill_1 FILLER_73_182 ();
 sg13g2_decap_8 FILLER_73_209 ();
 sg13g2_decap_8 FILLER_73_216 ();
 sg13g2_decap_4 FILLER_73_223 ();
 sg13g2_fill_2 FILLER_73_227 ();
 sg13g2_decap_4 FILLER_73_233 ();
 sg13g2_fill_2 FILLER_73_237 ();
 sg13g2_fill_2 FILLER_73_244 ();
 sg13g2_fill_1 FILLER_73_251 ();
 sg13g2_fill_2 FILLER_73_256 ();
 sg13g2_decap_8 FILLER_73_270 ();
 sg13g2_decap_8 FILLER_73_277 ();
 sg13g2_fill_2 FILLER_73_284 ();
 sg13g2_fill_1 FILLER_73_286 ();
 sg13g2_decap_4 FILLER_73_313 ();
 sg13g2_fill_1 FILLER_73_317 ();
 sg13g2_decap_8 FILLER_73_331 ();
 sg13g2_decap_4 FILLER_73_338 ();
 sg13g2_fill_2 FILLER_73_342 ();
 sg13g2_decap_8 FILLER_73_348 ();
 sg13g2_decap_8 FILLER_73_355 ();
 sg13g2_decap_8 FILLER_73_362 ();
 sg13g2_decap_4 FILLER_73_369 ();
 sg13g2_decap_8 FILLER_73_399 ();
 sg13g2_decap_8 FILLER_73_406 ();
 sg13g2_decap_8 FILLER_73_413 ();
 sg13g2_decap_8 FILLER_73_420 ();
 sg13g2_fill_1 FILLER_73_440 ();
 sg13g2_fill_2 FILLER_73_463 ();
 sg13g2_decap_4 FILLER_73_473 ();
 sg13g2_fill_1 FILLER_73_477 ();
 sg13g2_fill_1 FILLER_73_483 ();
 sg13g2_fill_2 FILLER_73_492 ();
 sg13g2_fill_1 FILLER_73_494 ();
 sg13g2_decap_8 FILLER_73_555 ();
 sg13g2_decap_8 FILLER_73_562 ();
 sg13g2_decap_8 FILLER_73_569 ();
 sg13g2_fill_1 FILLER_73_576 ();
 sg13g2_decap_8 FILLER_73_582 ();
 sg13g2_decap_4 FILLER_73_589 ();
 sg13g2_decap_8 FILLER_73_597 ();
 sg13g2_decap_8 FILLER_73_670 ();
 sg13g2_decap_4 FILLER_73_677 ();
 sg13g2_fill_1 FILLER_73_681 ();
 sg13g2_decap_8 FILLER_73_690 ();
 sg13g2_decap_8 FILLER_73_697 ();
 sg13g2_decap_8 FILLER_73_704 ();
 sg13g2_decap_8 FILLER_73_711 ();
 sg13g2_decap_8 FILLER_73_748 ();
 sg13g2_fill_1 FILLER_73_755 ();
 sg13g2_fill_2 FILLER_73_760 ();
 sg13g2_fill_1 FILLER_73_762 ();
 sg13g2_decap_4 FILLER_73_775 ();
 sg13g2_decap_8 FILLER_73_784 ();
 sg13g2_decap_8 FILLER_73_791 ();
 sg13g2_decap_8 FILLER_73_798 ();
 sg13g2_decap_8 FILLER_73_805 ();
 sg13g2_decap_8 FILLER_73_812 ();
 sg13g2_decap_8 FILLER_73_819 ();
 sg13g2_decap_8 FILLER_73_826 ();
 sg13g2_decap_8 FILLER_73_833 ();
 sg13g2_decap_8 FILLER_73_840 ();
 sg13g2_decap_8 FILLER_73_847 ();
 sg13g2_decap_8 FILLER_73_854 ();
 sg13g2_fill_1 FILLER_73_861 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_fill_2 FILLER_74_35 ();
 sg13g2_fill_2 FILLER_74_58 ();
 sg13g2_fill_1 FILLER_74_60 ();
 sg13g2_fill_2 FILLER_74_87 ();
 sg13g2_fill_2 FILLER_74_107 ();
 sg13g2_fill_1 FILLER_74_109 ();
 sg13g2_fill_2 FILLER_74_144 ();
 sg13g2_fill_2 FILLER_74_150 ();
 sg13g2_decap_8 FILLER_74_183 ();
 sg13g2_decap_4 FILLER_74_190 ();
 sg13g2_fill_2 FILLER_74_194 ();
 sg13g2_decap_8 FILLER_74_201 ();
 sg13g2_fill_2 FILLER_74_208 ();
 sg13g2_decap_8 FILLER_74_215 ();
 sg13g2_decap_4 FILLER_74_222 ();
 sg13g2_fill_1 FILLER_74_226 ();
 sg13g2_fill_2 FILLER_74_248 ();
 sg13g2_fill_2 FILLER_74_270 ();
 sg13g2_decap_8 FILLER_74_292 ();
 sg13g2_decap_8 FILLER_74_299 ();
 sg13g2_fill_2 FILLER_74_306 ();
 sg13g2_fill_2 FILLER_74_312 ();
 sg13g2_fill_1 FILLER_74_366 ();
 sg13g2_fill_2 FILLER_74_388 ();
 sg13g2_decap_4 FILLER_74_398 ();
 sg13g2_fill_2 FILLER_74_402 ();
 sg13g2_fill_2 FILLER_74_466 ();
 sg13g2_fill_1 FILLER_74_468 ();
 sg13g2_decap_4 FILLER_74_495 ();
 sg13g2_fill_2 FILLER_74_499 ();
 sg13g2_decap_8 FILLER_74_510 ();
 sg13g2_decap_8 FILLER_74_517 ();
 sg13g2_decap_8 FILLER_74_524 ();
 sg13g2_decap_8 FILLER_74_531 ();
 sg13g2_decap_8 FILLER_74_538 ();
 sg13g2_decap_4 FILLER_74_597 ();
 sg13g2_fill_2 FILLER_74_601 ();
 sg13g2_decap_8 FILLER_74_629 ();
 sg13g2_decap_4 FILLER_74_636 ();
 sg13g2_fill_1 FILLER_74_640 ();
 sg13g2_decap_8 FILLER_74_645 ();
 sg13g2_fill_2 FILLER_74_652 ();
 sg13g2_fill_1 FILLER_74_654 ();
 sg13g2_fill_2 FILLER_74_738 ();
 sg13g2_decap_8 FILLER_74_774 ();
 sg13g2_decap_8 FILLER_74_781 ();
 sg13g2_decap_8 FILLER_74_788 ();
 sg13g2_decap_8 FILLER_74_795 ();
 sg13g2_decap_8 FILLER_74_802 ();
 sg13g2_decap_8 FILLER_74_809 ();
 sg13g2_decap_8 FILLER_74_816 ();
 sg13g2_decap_8 FILLER_74_823 ();
 sg13g2_decap_8 FILLER_74_830 ();
 sg13g2_decap_8 FILLER_74_837 ();
 sg13g2_decap_8 FILLER_74_844 ();
 sg13g2_decap_8 FILLER_74_851 ();
 sg13g2_decap_4 FILLER_74_858 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_62 ();
 sg13g2_decap_8 FILLER_75_69 ();
 sg13g2_decap_8 FILLER_75_76 ();
 sg13g2_fill_1 FILLER_75_83 ();
 sg13g2_fill_2 FILLER_75_92 ();
 sg13g2_decap_8 FILLER_75_107 ();
 sg13g2_decap_8 FILLER_75_114 ();
 sg13g2_decap_8 FILLER_75_121 ();
 sg13g2_decap_8 FILLER_75_128 ();
 sg13g2_decap_8 FILLER_75_135 ();
 sg13g2_decap_4 FILLER_75_247 ();
 sg13g2_decap_4 FILLER_75_267 ();
 sg13g2_fill_1 FILLER_75_271 ();
 sg13g2_fill_1 FILLER_75_280 ();
 sg13g2_decap_8 FILLER_75_292 ();
 sg13g2_fill_2 FILLER_75_299 ();
 sg13g2_fill_2 FILLER_75_310 ();
 sg13g2_fill_1 FILLER_75_312 ();
 sg13g2_fill_2 FILLER_75_321 ();
 sg13g2_fill_1 FILLER_75_328 ();
 sg13g2_fill_2 FILLER_75_334 ();
 sg13g2_fill_1 FILLER_75_336 ();
 sg13g2_fill_2 FILLER_75_354 ();
 sg13g2_fill_1 FILLER_75_364 ();
 sg13g2_decap_8 FILLER_75_369 ();
 sg13g2_fill_2 FILLER_75_384 ();
 sg13g2_fill_1 FILLER_75_386 ();
 sg13g2_decap_8 FILLER_75_399 ();
 sg13g2_decap_8 FILLER_75_432 ();
 sg13g2_fill_2 FILLER_75_439 ();
 sg13g2_fill_1 FILLER_75_441 ();
 sg13g2_decap_8 FILLER_75_468 ();
 sg13g2_decap_8 FILLER_75_475 ();
 sg13g2_decap_8 FILLER_75_482 ();
 sg13g2_fill_2 FILLER_75_489 ();
 sg13g2_fill_2 FILLER_75_499 ();
 sg13g2_fill_1 FILLER_75_501 ();
 sg13g2_decap_8 FILLER_75_554 ();
 sg13g2_decap_4 FILLER_75_569 ();
 sg13g2_fill_1 FILLER_75_573 ();
 sg13g2_decap_4 FILLER_75_594 ();
 sg13g2_fill_2 FILLER_75_598 ();
 sg13g2_fill_1 FILLER_75_612 ();
 sg13g2_decap_8 FILLER_75_639 ();
 sg13g2_decap_8 FILLER_75_646 ();
 sg13g2_decap_4 FILLER_75_653 ();
 sg13g2_fill_2 FILLER_75_657 ();
 sg13g2_fill_2 FILLER_75_663 ();
 sg13g2_decap_8 FILLER_75_673 ();
 sg13g2_decap_8 FILLER_75_680 ();
 sg13g2_decap_8 FILLER_75_695 ();
 sg13g2_decap_8 FILLER_75_702 ();
 sg13g2_decap_4 FILLER_75_709 ();
 sg13g2_fill_1 FILLER_75_721 ();
 sg13g2_fill_2 FILLER_75_728 ();
 sg13g2_decap_8 FILLER_75_743 ();
 sg13g2_decap_8 FILLER_75_750 ();
 sg13g2_decap_8 FILLER_75_757 ();
 sg13g2_decap_8 FILLER_75_768 ();
 sg13g2_decap_8 FILLER_75_775 ();
 sg13g2_decap_8 FILLER_75_782 ();
 sg13g2_decap_8 FILLER_75_789 ();
 sg13g2_decap_8 FILLER_75_796 ();
 sg13g2_decap_8 FILLER_75_803 ();
 sg13g2_decap_8 FILLER_75_810 ();
 sg13g2_decap_8 FILLER_75_817 ();
 sg13g2_decap_8 FILLER_75_824 ();
 sg13g2_decap_8 FILLER_75_831 ();
 sg13g2_decap_8 FILLER_75_838 ();
 sg13g2_decap_8 FILLER_75_845 ();
 sg13g2_decap_8 FILLER_75_852 ();
 sg13g2_fill_2 FILLER_75_859 ();
 sg13g2_fill_1 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_fill_2 FILLER_76_35 ();
 sg13g2_fill_1 FILLER_76_58 ();
 sg13g2_fill_2 FILLER_76_85 ();
 sg13g2_fill_1 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_139 ();
 sg13g2_decap_4 FILLER_76_146 ();
 sg13g2_fill_1 FILLER_76_150 ();
 sg13g2_decap_4 FILLER_76_179 ();
 sg13g2_fill_2 FILLER_76_191 ();
 sg13g2_fill_1 FILLER_76_193 ();
 sg13g2_decap_4 FILLER_76_198 ();
 sg13g2_fill_1 FILLER_76_202 ();
 sg13g2_decap_8 FILLER_76_219 ();
 sg13g2_decap_8 FILLER_76_226 ();
 sg13g2_decap_4 FILLER_76_233 ();
 sg13g2_fill_2 FILLER_76_237 ();
 sg13g2_decap_8 FILLER_76_244 ();
 sg13g2_fill_1 FILLER_76_251 ();
 sg13g2_decap_8 FILLER_76_260 ();
 sg13g2_fill_2 FILLER_76_267 ();
 sg13g2_fill_1 FILLER_76_269 ();
 sg13g2_fill_2 FILLER_76_278 ();
 sg13g2_fill_1 FILLER_76_317 ();
 sg13g2_fill_2 FILLER_76_333 ();
 sg13g2_fill_1 FILLER_76_335 ();
 sg13g2_fill_2 FILLER_76_344 ();
 sg13g2_decap_8 FILLER_76_358 ();
 sg13g2_decap_8 FILLER_76_365 ();
 sg13g2_decap_4 FILLER_76_372 ();
 sg13g2_decap_8 FILLER_76_406 ();
 sg13g2_decap_8 FILLER_76_413 ();
 sg13g2_decap_4 FILLER_76_420 ();
 sg13g2_fill_2 FILLER_76_424 ();
 sg13g2_decap_8 FILLER_76_442 ();
 sg13g2_fill_1 FILLER_76_449 ();
 sg13g2_decap_8 FILLER_76_455 ();
 sg13g2_decap_8 FILLER_76_462 ();
 sg13g2_decap_8 FILLER_76_509 ();
 sg13g2_decap_8 FILLER_76_516 ();
 sg13g2_fill_1 FILLER_76_523 ();
 sg13g2_decap_4 FILLER_76_532 ();
 sg13g2_fill_1 FILLER_76_536 ();
 sg13g2_fill_1 FILLER_76_541 ();
 sg13g2_fill_2 FILLER_76_568 ();
 sg13g2_fill_1 FILLER_76_570 ();
 sg13g2_fill_1 FILLER_76_584 ();
 sg13g2_decap_4 FILLER_76_605 ();
 sg13g2_fill_1 FILLER_76_609 ();
 sg13g2_decap_4 FILLER_76_622 ();
 sg13g2_fill_1 FILLER_76_709 ();
 sg13g2_fill_2 FILLER_76_725 ();
 sg13g2_fill_1 FILLER_76_727 ();
 sg13g2_decap_8 FILLER_76_762 ();
 sg13g2_decap_8 FILLER_76_769 ();
 sg13g2_decap_8 FILLER_76_776 ();
 sg13g2_decap_8 FILLER_76_783 ();
 sg13g2_decap_8 FILLER_76_790 ();
 sg13g2_decap_8 FILLER_76_797 ();
 sg13g2_decap_8 FILLER_76_804 ();
 sg13g2_decap_8 FILLER_76_811 ();
 sg13g2_decap_8 FILLER_76_818 ();
 sg13g2_decap_8 FILLER_76_825 ();
 sg13g2_decap_8 FILLER_76_832 ();
 sg13g2_decap_8 FILLER_76_839 ();
 sg13g2_decap_8 FILLER_76_846 ();
 sg13g2_decap_8 FILLER_76_853 ();
 sg13g2_fill_2 FILLER_76_860 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_fill_1 FILLER_77_49 ();
 sg13g2_decap_4 FILLER_77_63 ();
 sg13g2_fill_2 FILLER_77_67 ();
 sg13g2_decap_8 FILLER_77_74 ();
 sg13g2_decap_4 FILLER_77_81 ();
 sg13g2_decap_8 FILLER_77_109 ();
 sg13g2_decap_4 FILLER_77_150 ();
 sg13g2_fill_2 FILLER_77_154 ();
 sg13g2_decap_4 FILLER_77_164 ();
 sg13g2_fill_2 FILLER_77_199 ();
 sg13g2_fill_1 FILLER_77_201 ();
 sg13g2_decap_8 FILLER_77_262 ();
 sg13g2_decap_4 FILLER_77_269 ();
 sg13g2_fill_2 FILLER_77_278 ();
 sg13g2_fill_1 FILLER_77_280 ();
 sg13g2_decap_4 FILLER_77_294 ();
 sg13g2_fill_2 FILLER_77_298 ();
 sg13g2_decap_8 FILLER_77_334 ();
 sg13g2_fill_1 FILLER_77_341 ();
 sg13g2_decap_8 FILLER_77_346 ();
 sg13g2_decap_4 FILLER_77_353 ();
 sg13g2_decap_4 FILLER_77_399 ();
 sg13g2_fill_2 FILLER_77_403 ();
 sg13g2_fill_2 FILLER_77_444 ();
 sg13g2_decap_4 FILLER_77_472 ();
 sg13g2_decap_8 FILLER_77_480 ();
 sg13g2_decap_4 FILLER_77_487 ();
 sg13g2_fill_1 FILLER_77_491 ();
 sg13g2_fill_1 FILLER_77_497 ();
 sg13g2_fill_2 FILLER_77_515 ();
 sg13g2_fill_2 FILLER_77_520 ();
 sg13g2_fill_1 FILLER_77_522 ();
 sg13g2_fill_2 FILLER_77_544 ();
 sg13g2_decap_8 FILLER_77_563 ();
 sg13g2_decap_8 FILLER_77_570 ();
 sg13g2_fill_1 FILLER_77_577 ();
 sg13g2_fill_2 FILLER_77_634 ();
 sg13g2_decap_8 FILLER_77_652 ();
 sg13g2_decap_8 FILLER_77_659 ();
 sg13g2_decap_8 FILLER_77_666 ();
 sg13g2_decap_8 FILLER_77_673 ();
 sg13g2_decap_8 FILLER_77_680 ();
 sg13g2_fill_2 FILLER_77_707 ();
 sg13g2_decap_8 FILLER_77_738 ();
 sg13g2_decap_8 FILLER_77_745 ();
 sg13g2_decap_8 FILLER_77_752 ();
 sg13g2_decap_8 FILLER_77_759 ();
 sg13g2_decap_8 FILLER_77_766 ();
 sg13g2_decap_8 FILLER_77_773 ();
 sg13g2_decap_8 FILLER_77_780 ();
 sg13g2_decap_8 FILLER_77_787 ();
 sg13g2_decap_8 FILLER_77_794 ();
 sg13g2_decap_8 FILLER_77_801 ();
 sg13g2_decap_8 FILLER_77_808 ();
 sg13g2_decap_8 FILLER_77_815 ();
 sg13g2_decap_8 FILLER_77_822 ();
 sg13g2_decap_8 FILLER_77_829 ();
 sg13g2_decap_8 FILLER_77_836 ();
 sg13g2_decap_8 FILLER_77_843 ();
 sg13g2_decap_8 FILLER_77_850 ();
 sg13g2_decap_4 FILLER_77_857 ();
 sg13g2_fill_1 FILLER_77_861 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_fill_2 FILLER_78_56 ();
 sg13g2_fill_1 FILLER_78_58 ();
 sg13g2_decap_8 FILLER_78_90 ();
 sg13g2_fill_2 FILLER_78_123 ();
 sg13g2_fill_1 FILLER_78_125 ();
 sg13g2_decap_8 FILLER_78_148 ();
 sg13g2_decap_4 FILLER_78_155 ();
 sg13g2_fill_2 FILLER_78_167 ();
 sg13g2_fill_1 FILLER_78_169 ();
 sg13g2_decap_8 FILLER_78_196 ();
 sg13g2_decap_4 FILLER_78_203 ();
 sg13g2_fill_1 FILLER_78_207 ();
 sg13g2_decap_8 FILLER_78_226 ();
 sg13g2_fill_2 FILLER_78_233 ();
 sg13g2_decap_8 FILLER_78_259 ();
 sg13g2_fill_1 FILLER_78_276 ();
 sg13g2_decap_8 FILLER_78_281 ();
 sg13g2_fill_1 FILLER_78_288 ();
 sg13g2_decap_8 FILLER_78_303 ();
 sg13g2_decap_8 FILLER_78_310 ();
 sg13g2_decap_8 FILLER_78_317 ();
 sg13g2_decap_8 FILLER_78_324 ();
 sg13g2_decap_4 FILLER_78_331 ();
 sg13g2_fill_2 FILLER_78_340 ();
 sg13g2_decap_8 FILLER_78_374 ();
 sg13g2_decap_8 FILLER_78_381 ();
 sg13g2_fill_1 FILLER_78_388 ();
 sg13g2_decap_8 FILLER_78_404 ();
 sg13g2_decap_8 FILLER_78_411 ();
 sg13g2_decap_8 FILLER_78_418 ();
 sg13g2_fill_2 FILLER_78_425 ();
 sg13g2_fill_1 FILLER_78_427 ();
 sg13g2_decap_8 FILLER_78_432 ();
 sg13g2_fill_1 FILLER_78_439 ();
 sg13g2_decap_4 FILLER_78_456 ();
 sg13g2_fill_2 FILLER_78_507 ();
 sg13g2_fill_1 FILLER_78_526 ();
 sg13g2_fill_1 FILLER_78_535 ();
 sg13g2_fill_1 FILLER_78_541 ();
 sg13g2_fill_2 FILLER_78_550 ();
 sg13g2_fill_1 FILLER_78_552 ();
 sg13g2_decap_8 FILLER_78_561 ();
 sg13g2_decap_8 FILLER_78_568 ();
 sg13g2_decap_8 FILLER_78_575 ();
 sg13g2_decap_4 FILLER_78_582 ();
 sg13g2_fill_2 FILLER_78_586 ();
 sg13g2_decap_8 FILLER_78_593 ();
 sg13g2_decap_8 FILLER_78_600 ();
 sg13g2_fill_2 FILLER_78_607 ();
 sg13g2_decap_8 FILLER_78_617 ();
 sg13g2_decap_8 FILLER_78_624 ();
 sg13g2_decap_8 FILLER_78_631 ();
 sg13g2_decap_8 FILLER_78_643 ();
 sg13g2_decap_8 FILLER_78_650 ();
 sg13g2_decap_8 FILLER_78_657 ();
 sg13g2_decap_8 FILLER_78_664 ();
 sg13g2_decap_8 FILLER_78_671 ();
 sg13g2_decap_8 FILLER_78_678 ();
 sg13g2_decap_8 FILLER_78_685 ();
 sg13g2_fill_1 FILLER_78_692 ();
 sg13g2_fill_2 FILLER_78_697 ();
 sg13g2_fill_1 FILLER_78_699 ();
 sg13g2_decap_8 FILLER_78_709 ();
 sg13g2_decap_8 FILLER_78_716 ();
 sg13g2_decap_8 FILLER_78_723 ();
 sg13g2_decap_8 FILLER_78_730 ();
 sg13g2_decap_8 FILLER_78_737 ();
 sg13g2_decap_8 FILLER_78_744 ();
 sg13g2_decap_8 FILLER_78_751 ();
 sg13g2_decap_8 FILLER_78_758 ();
 sg13g2_decap_8 FILLER_78_765 ();
 sg13g2_decap_8 FILLER_78_772 ();
 sg13g2_decap_8 FILLER_78_779 ();
 sg13g2_decap_8 FILLER_78_786 ();
 sg13g2_decap_8 FILLER_78_793 ();
 sg13g2_decap_8 FILLER_78_800 ();
 sg13g2_decap_8 FILLER_78_807 ();
 sg13g2_decap_8 FILLER_78_814 ();
 sg13g2_decap_8 FILLER_78_821 ();
 sg13g2_decap_8 FILLER_78_828 ();
 sg13g2_decap_8 FILLER_78_835 ();
 sg13g2_decap_8 FILLER_78_842 ();
 sg13g2_decap_8 FILLER_78_849 ();
 sg13g2_decap_4 FILLER_78_856 ();
 sg13g2_fill_2 FILLER_78_860 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_fill_1 FILLER_79_126 ();
 sg13g2_fill_2 FILLER_79_143 ();
 sg13g2_fill_1 FILLER_79_166 ();
 sg13g2_fill_1 FILLER_79_219 ();
 sg13g2_fill_2 FILLER_79_254 ();
 sg13g2_fill_2 FILLER_79_301 ();
 sg13g2_fill_1 FILLER_79_303 ();
 sg13g2_fill_1 FILLER_79_334 ();
 sg13g2_decap_8 FILLER_79_370 ();
 sg13g2_decap_8 FILLER_79_377 ();
 sg13g2_decap_4 FILLER_79_384 ();
 sg13g2_fill_1 FILLER_79_388 ();
 sg13g2_decap_8 FILLER_79_405 ();
 sg13g2_decap_8 FILLER_79_412 ();
 sg13g2_decap_8 FILLER_79_419 ();
 sg13g2_fill_2 FILLER_79_452 ();
 sg13g2_decap_8 FILLER_79_487 ();
 sg13g2_decap_8 FILLER_79_506 ();
 sg13g2_decap_8 FILLER_79_513 ();
 sg13g2_decap_8 FILLER_79_520 ();
 sg13g2_fill_2 FILLER_79_527 ();
 sg13g2_fill_1 FILLER_79_529 ();
 sg13g2_decap_8 FILLER_79_534 ();
 sg13g2_decap_8 FILLER_79_541 ();
 sg13g2_decap_8 FILLER_79_548 ();
 sg13g2_decap_8 FILLER_79_555 ();
 sg13g2_decap_8 FILLER_79_562 ();
 sg13g2_decap_8 FILLER_79_569 ();
 sg13g2_decap_8 FILLER_79_576 ();
 sg13g2_decap_8 FILLER_79_583 ();
 sg13g2_decap_8 FILLER_79_590 ();
 sg13g2_decap_8 FILLER_79_597 ();
 sg13g2_decap_8 FILLER_79_604 ();
 sg13g2_decap_8 FILLER_79_611 ();
 sg13g2_decap_8 FILLER_79_618 ();
 sg13g2_decap_8 FILLER_79_625 ();
 sg13g2_decap_8 FILLER_79_632 ();
 sg13g2_decap_8 FILLER_79_639 ();
 sg13g2_decap_8 FILLER_79_646 ();
 sg13g2_decap_8 FILLER_79_653 ();
 sg13g2_decap_8 FILLER_79_660 ();
 sg13g2_decap_8 FILLER_79_667 ();
 sg13g2_decap_8 FILLER_79_674 ();
 sg13g2_decap_8 FILLER_79_681 ();
 sg13g2_decap_8 FILLER_79_688 ();
 sg13g2_decap_8 FILLER_79_695 ();
 sg13g2_decap_8 FILLER_79_702 ();
 sg13g2_decap_8 FILLER_79_709 ();
 sg13g2_decap_8 FILLER_79_716 ();
 sg13g2_decap_8 FILLER_79_723 ();
 sg13g2_decap_8 FILLER_79_730 ();
 sg13g2_decap_8 FILLER_79_737 ();
 sg13g2_decap_8 FILLER_79_744 ();
 sg13g2_decap_8 FILLER_79_751 ();
 sg13g2_decap_8 FILLER_79_758 ();
 sg13g2_decap_8 FILLER_79_765 ();
 sg13g2_decap_8 FILLER_79_772 ();
 sg13g2_decap_8 FILLER_79_779 ();
 sg13g2_decap_8 FILLER_79_786 ();
 sg13g2_decap_8 FILLER_79_793 ();
 sg13g2_decap_8 FILLER_79_800 ();
 sg13g2_decap_8 FILLER_79_807 ();
 sg13g2_decap_8 FILLER_79_814 ();
 sg13g2_decap_8 FILLER_79_821 ();
 sg13g2_decap_8 FILLER_79_828 ();
 sg13g2_decap_8 FILLER_79_835 ();
 sg13g2_decap_8 FILLER_79_842 ();
 sg13g2_decap_8 FILLER_79_849 ();
 sg13g2_decap_4 FILLER_79_856 ();
 sg13g2_fill_2 FILLER_79_860 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_fill_2 FILLER_80_124 ();
 sg13g2_fill_1 FILLER_80_175 ();
 sg13g2_decap_4 FILLER_80_180 ();
 sg13g2_decap_4 FILLER_80_188 ();
 sg13g2_decap_4 FILLER_80_196 ();
 sg13g2_decap_4 FILLER_80_204 ();
 sg13g2_fill_2 FILLER_80_212 ();
 sg13g2_decap_8 FILLER_80_222 ();
 sg13g2_decap_8 FILLER_80_229 ();
 sg13g2_decap_8 FILLER_80_236 ();
 sg13g2_decap_8 FILLER_80_243 ();
 sg13g2_decap_8 FILLER_80_250 ();
 sg13g2_decap_8 FILLER_80_257 ();
 sg13g2_decap_8 FILLER_80_268 ();
 sg13g2_decap_8 FILLER_80_275 ();
 sg13g2_fill_2 FILLER_80_282 ();
 sg13g2_fill_1 FILLER_80_284 ();
 sg13g2_decap_4 FILLER_80_302 ();
 sg13g2_fill_2 FILLER_80_332 ();
 sg13g2_fill_1 FILLER_80_334 ();
 sg13g2_fill_1 FILLER_80_371 ();
 sg13g2_decap_8 FILLER_80_398 ();
 sg13g2_decap_8 FILLER_80_405 ();
 sg13g2_decap_8 FILLER_80_412 ();
 sg13g2_decap_8 FILLER_80_419 ();
 sg13g2_decap_8 FILLER_80_426 ();
 sg13g2_decap_8 FILLER_80_433 ();
 sg13g2_decap_8 FILLER_80_440 ();
 sg13g2_fill_1 FILLER_80_447 ();
 sg13g2_decap_8 FILLER_80_452 ();
 sg13g2_decap_8 FILLER_80_459 ();
 sg13g2_fill_1 FILLER_80_466 ();
 sg13g2_decap_8 FILLER_80_475 ();
 sg13g2_decap_8 FILLER_80_482 ();
 sg13g2_decap_8 FILLER_80_489 ();
 sg13g2_decap_8 FILLER_80_496 ();
 sg13g2_decap_8 FILLER_80_503 ();
 sg13g2_decap_8 FILLER_80_510 ();
 sg13g2_decap_8 FILLER_80_517 ();
 sg13g2_decap_8 FILLER_80_524 ();
 sg13g2_decap_8 FILLER_80_531 ();
 sg13g2_decap_8 FILLER_80_538 ();
 sg13g2_decap_8 FILLER_80_545 ();
 sg13g2_decap_8 FILLER_80_552 ();
 sg13g2_decap_8 FILLER_80_559 ();
 sg13g2_decap_8 FILLER_80_566 ();
 sg13g2_decap_8 FILLER_80_573 ();
 sg13g2_decap_8 FILLER_80_580 ();
 sg13g2_decap_8 FILLER_80_587 ();
 sg13g2_decap_8 FILLER_80_594 ();
 sg13g2_decap_8 FILLER_80_601 ();
 sg13g2_decap_8 FILLER_80_608 ();
 sg13g2_decap_8 FILLER_80_615 ();
 sg13g2_decap_8 FILLER_80_622 ();
 sg13g2_decap_8 FILLER_80_629 ();
 sg13g2_decap_8 FILLER_80_636 ();
 sg13g2_decap_8 FILLER_80_643 ();
 sg13g2_decap_8 FILLER_80_650 ();
 sg13g2_decap_8 FILLER_80_657 ();
 sg13g2_decap_8 FILLER_80_664 ();
 sg13g2_decap_8 FILLER_80_671 ();
 sg13g2_decap_8 FILLER_80_678 ();
 sg13g2_decap_8 FILLER_80_685 ();
 sg13g2_decap_8 FILLER_80_692 ();
 sg13g2_decap_8 FILLER_80_699 ();
 sg13g2_decap_8 FILLER_80_706 ();
 sg13g2_decap_8 FILLER_80_713 ();
 sg13g2_decap_8 FILLER_80_720 ();
 sg13g2_decap_8 FILLER_80_727 ();
 sg13g2_decap_8 FILLER_80_734 ();
 sg13g2_decap_8 FILLER_80_741 ();
 sg13g2_decap_8 FILLER_80_748 ();
 sg13g2_decap_8 FILLER_80_755 ();
 sg13g2_decap_8 FILLER_80_762 ();
 sg13g2_decap_8 FILLER_80_769 ();
 sg13g2_decap_8 FILLER_80_776 ();
 sg13g2_decap_8 FILLER_80_783 ();
 sg13g2_decap_8 FILLER_80_790 ();
 sg13g2_decap_8 FILLER_80_797 ();
 sg13g2_decap_8 FILLER_80_804 ();
 sg13g2_decap_8 FILLER_80_811 ();
 sg13g2_decap_8 FILLER_80_818 ();
 sg13g2_decap_8 FILLER_80_825 ();
 sg13g2_decap_8 FILLER_80_832 ();
 sg13g2_decap_8 FILLER_80_839 ();
 sg13g2_decap_8 FILLER_80_846 ();
 sg13g2_decap_8 FILLER_80_853 ();
 sg13g2_fill_2 FILLER_80_860 ();
 assign uio_oe[0] = net4;
 assign uio_oe[1] = net5;
 assign uio_oe[2] = net6;
 assign uio_oe[3] = net7;
 assign uio_oe[4] = net8;
 assign uio_oe[5] = net9;
 assign uio_oe[6] = net10;
 assign uio_oe[7] = net11;
 assign uio_out[0] = net12;
 assign uio_out[1] = net13;
 assign uio_out[2] = net14;
 assign uio_out[3] = net15;
 assign uio_out[4] = net16;
 assign uio_out[5] = net17;
 assign uio_out[6] = net18;
 assign uio_out[7] = net19;
 assign uo_out[4] = net20;
 assign uo_out[5] = net21;
 assign uo_out[6] = net22;
 assign uo_out[7] = net23;
endmodule

module tt_um_meriac_play_tune (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \db_entry[0] ;
 wire \db_entry[10] ;
 wire \db_entry[11] ;
 wire \db_entry[1] ;
 wire \db_entry[2] ;
 wire \db_entry[3] ;
 wire \db_entry[4] ;
 wire \db_entry[5] ;
 wire \db_entry[6] ;
 wire \db_entry[7] ;
 wire \db_entry[8] ;
 wire \db_entry[9] ;
 wire \freq[0] ;
 wire \freq[1] ;
 wire \freq[2] ;
 wire \freq[3] ;
 wire \freq[4] ;
 wire \freq[5] ;
 wire \freq[6] ;
 wire \freq[7] ;
 wire \meriac_tune_db.address[0] ;
 wire \meriac_tune_db.address[1] ;
 wire \meriac_tune_db.address[2] ;
 wire \meriac_tune_db.address[3] ;
 wire \meriac_tune_db.address[4] ;
 wire \meriac_tune_db.address[5] ;
 wire \meriac_tune_db.address[6] ;
 wire speaker;
 wire \ticks[0] ;
 wire \ticks[10] ;
 wire \ticks[11] ;
 wire \ticks[12] ;
 wire \ticks[13] ;
 wire \ticks[14] ;
 wire \ticks[15] ;
 wire \ticks[1] ;
 wire \ticks[2] ;
 wire \ticks[3] ;
 wire \ticks[4] ;
 wire \ticks[5] ;
 wire \ticks[6] ;
 wire \ticks[7] ;
 wire \ticks[8] ;
 wire \ticks[9] ;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire clknet_0_clk;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net1;
 wire net2;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;

 sg13g2_inv_1 _478_ (.Y(_062_),
    .A(\freq[7] ));
 sg13g2_inv_1 _479_ (.Y(_063_),
    .A(net82));
 sg13g2_inv_1 _480_ (.Y(_064_),
    .A(net110));
 sg13g2_inv_1 _481_ (.Y(_065_),
    .A(net122));
 sg13g2_inv_1 _482_ (.Y(_066_),
    .A(net76));
 sg13g2_inv_1 _483_ (.Y(_067_),
    .A(\freq[2] ));
 sg13g2_inv_1 _484_ (.Y(_068_),
    .A(net100));
 sg13g2_inv_1 _485_ (.Y(_069_),
    .A(net83));
 sg13g2_inv_1 _486_ (.Y(_070_),
    .A(net77));
 sg13g2_inv_1 _487_ (.Y(_071_),
    .A(net124));
 sg13g2_inv_1 _488_ (.Y(_072_),
    .A(\meriac_tune_db.address[4] ));
 sg13g2_inv_1 _489_ (.Y(_073_),
    .A(net120));
 sg13g2_inv_1 _490_ (.Y(_074_),
    .A(net111));
 sg13g2_inv_1 _491_ (.Y(_075_),
    .A(net179));
 sg13g2_inv_2 _492_ (.Y(_076_),
    .A(net166));
 sg13g2_inv_1 _493_ (.Y(_077_),
    .A(_011_));
 sg13g2_inv_1 _494_ (.Y(_078_),
    .A(_017_));
 sg13g2_inv_1 _495_ (.Y(_079_),
    .A(\counter[4] ));
 sg13g2_inv_1 _496_ (.Y(_080_),
    .A(\counter[3] ));
 sg13g2_nor3_1 _497_ (.A(\ticks[0] ),
    .B(net182),
    .C(net171),
    .Y(_081_));
 sg13g2_nor4_2 _498_ (.A(\ticks[0] ),
    .B(net106),
    .C(\ticks[2] ),
    .Y(_082_),
    .D(\ticks[1] ));
 sg13g2_nand2b_1 _499_ (.Y(_083_),
    .B(_081_),
    .A_N(net106));
 sg13g2_nor2_1 _500_ (.A(\ticks[4] ),
    .B(net90),
    .Y(_084_));
 sg13g2_nand2_1 _501_ (.Y(_085_),
    .A(_082_),
    .B(_084_));
 sg13g2_nor2_1 _502_ (.A(net85),
    .B(\ticks[6] ),
    .Y(_086_));
 sg13g2_nand3_1 _503_ (.B(_084_),
    .C(_086_),
    .A(_082_),
    .Y(_087_));
 sg13g2_nor4_1 _504_ (.A(\ticks[10] ),
    .B(net79),
    .C(\ticks[9] ),
    .D(\ticks[8] ),
    .Y(_088_));
 sg13g2_nand4_1 _505_ (.B(_084_),
    .C(_086_),
    .A(_082_),
    .Y(_089_),
    .D(_088_));
 sg13g2_nor3_1 _506_ (.A(net117),
    .B(\ticks[12] ),
    .C(_089_),
    .Y(_090_));
 sg13g2_or2_1 _507_ (.X(_091_),
    .B(\ticks[14] ),
    .A(\ticks[15] ));
 sg13g2_nor4_1 _508_ (.A(\ticks[13] ),
    .B(\ticks[12] ),
    .C(_089_),
    .D(_091_),
    .Y(_092_));
 sg13g2_or4_1 _509_ (.A(\ticks[13] ),
    .B(\ticks[12] ),
    .C(_089_),
    .D(_091_),
    .X(_093_));
 sg13g2_nor3_1 _510_ (.A(_071_),
    .B(\meriac_tune_db.address[4] ),
    .C(\meriac_tune_db.address[3] ),
    .Y(_094_));
 sg13g2_or2_1 _511_ (.X(_095_),
    .B(\meriac_tune_db.address[0] ),
    .A(\meriac_tune_db.address[1] ));
 sg13g2_o21ai_1 _512_ (.B1(\meriac_tune_db.address[2] ),
    .Y(_096_),
    .A1(\meriac_tune_db.address[1] ),
    .A2(\meriac_tune_db.address[0] ));
 sg13g2_nand4_1 _513_ (.B(_072_),
    .C(_073_),
    .A(\meriac_tune_db.address[5] ),
    .Y(_097_),
    .D(_096_));
 sg13g2_nor2_1 _514_ (.A(_070_),
    .B(_011_),
    .Y(_098_));
 sg13g2_nor3_1 _515_ (.A(_074_),
    .B(_010_),
    .C(_095_),
    .Y(_099_));
 sg13g2_a22oi_1 _516_ (.Y(_100_),
    .B1(_099_),
    .B2(_094_),
    .A2(_098_),
    .A1(_097_));
 sg13g2_and3_1 _517_ (.X(_101_),
    .A(net168),
    .B(net163),
    .C(_100_));
 sg13g2_nand2_2 _518_ (.Y(_102_),
    .A(\meriac_tune_db.address[1] ),
    .B(\meriac_tune_db.address[0] ));
 sg13g2_nand4_1 _519_ (.B(\meriac_tune_db.address[2] ),
    .C(\meriac_tune_db.address[1] ),
    .A(\meriac_tune_db.address[3] ),
    .Y(_103_),
    .D(\meriac_tune_db.address[0] ));
 sg13g2_or3_1 _520_ (.A(_071_),
    .B(_072_),
    .C(_103_),
    .X(_104_));
 sg13g2_xor2_1 _521_ (.B(_104_),
    .A(_010_),
    .X(_105_));
 sg13g2_nand2_1 _522_ (.Y(_106_),
    .A(_101_),
    .B(_105_));
 sg13g2_nor2_1 _523_ (.A(_076_),
    .B(net162),
    .Y(_107_));
 sg13g2_nand2_1 _524_ (.Y(_108_),
    .A(net167),
    .B(net161));
 sg13g2_o21ai_1 _525_ (.B1(_106_),
    .Y(_109_),
    .A1(_010_),
    .A2(net155));
 sg13g2_inv_1 _526_ (.Y(_110_),
    .A(net127));
 sg13g2_nor2_1 _527_ (.A(_017_),
    .B(_103_),
    .Y(_111_));
 sg13g2_xnor2_1 _528_ (.Y(_112_),
    .A(_078_),
    .B(_103_));
 sg13g2_and4_1 _529_ (.A(net168),
    .B(net163),
    .C(net159),
    .D(_112_),
    .X(_113_));
 sg13g2_a21oi_1 _530_ (.A1(_078_),
    .A2(net158),
    .Y(_114_),
    .B1(_113_));
 sg13g2_a21o_1 _531_ (.A2(net158),
    .A1(_078_),
    .B1(_113_),
    .X(_115_));
 sg13g2_nor2_1 _532_ (.A(_015_),
    .B(_102_),
    .Y(_116_));
 sg13g2_xnor2_1 _533_ (.Y(_117_),
    .A(_016_),
    .B(_116_));
 sg13g2_nand4_1 _534_ (.B(net163),
    .C(net159),
    .A(net168),
    .Y(_118_),
    .D(_117_));
 sg13g2_nand3b_1 _535_ (.B(net161),
    .C(net166),
    .Y(_119_),
    .A_N(_016_));
 sg13g2_and2_1 _536_ (.A(_118_),
    .B(_119_),
    .X(_120_));
 sg13g2_nand2_1 _537_ (.Y(_121_),
    .A(_118_),
    .B(_119_));
 sg13g2_nor2_1 _538_ (.A(net147),
    .B(net141),
    .Y(_122_));
 sg13g2_nand2_2 _539_ (.Y(_123_),
    .A(net149),
    .B(net143));
 sg13g2_nor2_1 _540_ (.A(\meriac_tune_db.address[0] ),
    .B(_076_),
    .Y(_124_));
 sg13g2_a22oi_1 _541_ (.Y(_125_),
    .B1(net159),
    .B2(_124_),
    .A2(net160),
    .A1(net167));
 sg13g2_and2_1 _542_ (.A(_013_),
    .B(net160),
    .X(_126_));
 sg13g2_nor2_1 _543_ (.A(_125_),
    .B(_126_),
    .Y(_127_));
 sg13g2_or2_1 _544_ (.X(_128_),
    .B(_126_),
    .A(_125_));
 sg13g2_xor2_1 _545_ (.B(_102_),
    .A(_015_),
    .X(_129_));
 sg13g2_and4_1 _546_ (.A(net166),
    .B(net162),
    .C(net159),
    .D(_129_),
    .X(_130_));
 sg13g2_nand4_1 _547_ (.B(net162),
    .C(net159),
    .A(net166),
    .Y(_131_),
    .D(_129_));
 sg13g2_nor3_2 _548_ (.A(_076_),
    .B(_015_),
    .C(net162),
    .Y(_132_));
 sg13g2_nand3b_1 _549_ (.B(net160),
    .C(net166),
    .Y(_133_),
    .A_N(_015_));
 sg13g2_nor2_2 _550_ (.A(_130_),
    .B(_132_),
    .Y(_134_));
 sg13g2_nand2_2 _551_ (.Y(_135_),
    .A(_131_),
    .B(_133_));
 sg13g2_and4_1 _552_ (.A(net162),
    .B(_095_),
    .C(net159),
    .D(_102_),
    .X(_136_));
 sg13g2_nand4_1 _553_ (.B(_095_),
    .C(net159),
    .A(net162),
    .Y(_137_),
    .D(_102_));
 sg13g2_nor2_1 _554_ (.A(_014_),
    .B(net162),
    .Y(_138_));
 sg13g2_nand2b_1 _555_ (.Y(_139_),
    .B(net160),
    .A_N(_014_));
 sg13g2_a21oi_1 _556_ (.A1(_137_),
    .A2(_139_),
    .Y(_140_),
    .B1(_076_));
 sg13g2_o21ai_1 _557_ (.B1(net166),
    .Y(_141_),
    .A1(_136_),
    .A2(_138_));
 sg13g2_a221oi_1 _558_ (.B2(_139_),
    .C1(_076_),
    .B1(_137_),
    .A1(_131_),
    .Y(_142_),
    .A2(_133_));
 sg13g2_nand2_1 _559_ (.Y(_143_),
    .A(net135),
    .B(net133));
 sg13g2_nand2_1 _560_ (.Y(_144_),
    .A(net137),
    .B(net133));
 sg13g2_and2_2 _561_ (.A(net138),
    .B(_142_),
    .X(_145_));
 sg13g2_nand2_2 _562_ (.Y(_146_),
    .A(net139),
    .B(net132));
 sg13g2_nor4_2 _563_ (.A(_125_),
    .B(_126_),
    .C(_130_),
    .Y(_147_),
    .D(_132_));
 sg13g2_xnor2_1 _564_ (.Y(_148_),
    .A(net139),
    .B(_142_));
 sg13g2_nor2_2 _565_ (.A(net147),
    .B(net144),
    .Y(_149_));
 sg13g2_nand2_1 _566_ (.Y(_150_),
    .A(net149),
    .B(net142));
 sg13g2_nand2_1 _567_ (.Y(_151_),
    .A(net137),
    .B(net135));
 sg13g2_nand2_1 _568_ (.Y(_152_),
    .A(_134_),
    .B(net132));
 sg13g2_a221oi_1 _569_ (.B2(_133_),
    .C1(_125_),
    .B1(_131_),
    .A1(_013_),
    .Y(_153_),
    .A2(net160));
 sg13g2_nand2_1 _570_ (.Y(_154_),
    .A(net139),
    .B(net135));
 sg13g2_nand4_1 _571_ (.B(_149_),
    .C(_151_),
    .A(_143_),
    .Y(_155_),
    .D(_152_));
 sg13g2_xnor2_1 _572_ (.Y(_156_),
    .A(_011_),
    .B(_111_));
 sg13g2_nand4_1 _573_ (.B(net163),
    .C(net159),
    .A(net168),
    .Y(_157_),
    .D(_156_));
 sg13g2_a22oi_1 _574_ (.Y(_158_),
    .B1(_156_),
    .B2(_101_),
    .A2(net158),
    .A1(_077_));
 sg13g2_o21ai_1 _575_ (.B1(_157_),
    .Y(_159_),
    .A1(_011_),
    .A2(net155));
 sg13g2_nand3_1 _576_ (.B(_134_),
    .C(net133),
    .A(net145),
    .Y(_160_));
 sg13g2_a221oi_1 _577_ (.B2(net148),
    .C1(net130),
    .B1(_160_),
    .A1(_122_),
    .Y(_161_),
    .A2(_148_));
 sg13g2_a21oi_1 _578_ (.A1(_155_),
    .A2(_161_),
    .Y(_162_),
    .B1(net127));
 sg13g2_nor2_2 _579_ (.A(net139),
    .B(net135),
    .Y(_163_));
 sg13g2_nor3_2 _580_ (.A(net140),
    .B(net136),
    .C(net131),
    .Y(_164_));
 sg13g2_nor2_1 _581_ (.A(net144),
    .B(_164_),
    .Y(_165_));
 sg13g2_a21oi_2 _582_ (.B1(_153_),
    .Y(_166_),
    .A2(net131),
    .A1(net139));
 sg13g2_o21ai_1 _583_ (.B1(net144),
    .Y(_167_),
    .A1(net136),
    .A2(net134));
 sg13g2_nor2_2 _584_ (.A(net138),
    .B(net131),
    .Y(_168_));
 sg13g2_nor2_2 _585_ (.A(net140),
    .B(net134),
    .Y(_169_));
 sg13g2_nand2_1 _586_ (.Y(_170_),
    .A(net137),
    .B(net132));
 sg13g2_or3_1 _587_ (.A(_167_),
    .B(_168_),
    .C(_169_),
    .X(_171_));
 sg13g2_nor2_2 _588_ (.A(net149),
    .B(_159_),
    .Y(_172_));
 sg13g2_nand2_1 _589_ (.Y(_173_),
    .A(net147),
    .B(net129));
 sg13g2_a21oi_1 _590_ (.A1(_165_),
    .A2(_166_),
    .Y(_174_),
    .B1(_173_));
 sg13g2_a21oi_2 _591_ (.B1(_153_),
    .Y(_175_),
    .A2(net134),
    .A1(net139));
 sg13g2_nand2b_1 _592_ (.Y(_176_),
    .B(net141),
    .A_N(_175_));
 sg13g2_nor2_2 _593_ (.A(net141),
    .B(net134),
    .Y(_177_));
 sg13g2_nand2_1 _594_ (.Y(_178_),
    .A(_154_),
    .B(_177_));
 sg13g2_nand2_1 _595_ (.Y(_179_),
    .A(net149),
    .B(net129));
 sg13g2_nor2b_1 _596_ (.A(_179_),
    .B_N(_176_),
    .Y(_180_));
 sg13g2_a22oi_1 _597_ (.Y(_181_),
    .B1(_178_),
    .B2(_180_),
    .A2(_174_),
    .A1(_171_));
 sg13g2_nand2_1 _598_ (.Y(_182_),
    .A(net141),
    .B(_153_));
 sg13g2_nand2_1 _599_ (.Y(_183_),
    .A(net143),
    .B(_164_));
 sg13g2_nor2_1 _600_ (.A(net145),
    .B(net139),
    .Y(_184_));
 sg13g2_nand2_2 _601_ (.Y(_185_),
    .A(net141),
    .B(_145_));
 sg13g2_a21oi_1 _602_ (.A1(net144),
    .A2(_164_),
    .Y(_186_),
    .B1(_179_));
 sg13g2_a22oi_1 _603_ (.Y(_187_),
    .B1(_185_),
    .B2(_186_),
    .A2(_182_),
    .A1(_172_));
 sg13g2_nand3_1 _604_ (.B(_159_),
    .C(_163_),
    .A(net126),
    .Y(_188_));
 sg13g2_and4_2 _605_ (.A(net127),
    .B(net126),
    .C(_159_),
    .D(_163_),
    .X(_189_));
 sg13g2_a21oi_1 _606_ (.A1(_187_),
    .A2(_188_),
    .Y(_190_),
    .B1(_110_));
 sg13g2_a21o_1 _607_ (.A2(_181_),
    .A1(_162_),
    .B1(_190_),
    .X(_000_));
 sg13g2_nand4_1 _608_ (.B(_147_),
    .C(_149_),
    .A(net131),
    .Y(_191_),
    .D(_159_));
 sg13g2_nand3_1 _609_ (.B(net138),
    .C(net135),
    .A(net145),
    .Y(_192_));
 sg13g2_nand4_1 _610_ (.B(net136),
    .C(_172_),
    .A(net138),
    .Y(_193_),
    .D(_177_));
 sg13g2_nand3_1 _611_ (.B(_191_),
    .C(_193_),
    .A(_110_),
    .Y(_194_));
 sg13g2_nor3_1 _612_ (.A(_123_),
    .B(net136),
    .C(_168_),
    .Y(_195_));
 sg13g2_nor2_1 _613_ (.A(_179_),
    .B(_185_),
    .Y(_196_));
 sg13g2_o21ai_1 _614_ (.B1(net127),
    .Y(_197_),
    .A1(net129),
    .A2(_195_));
 sg13g2_o21ai_1 _615_ (.B1(_194_),
    .Y(_002_),
    .A1(_196_),
    .A2(_197_));
 sg13g2_nor2_2 _616_ (.A(net142),
    .B(_142_),
    .Y(_198_));
 sg13g2_nand2_1 _617_ (.Y(_199_),
    .A(_175_),
    .B(_198_));
 sg13g2_a22oi_1 _618_ (.Y(_200_),
    .B1(_180_),
    .B2(_199_),
    .A2(_174_),
    .A1(_171_));
 sg13g2_a21oi_1 _619_ (.A1(net126),
    .A2(_147_),
    .Y(_201_),
    .B1(net129));
 sg13g2_nand2b_1 _620_ (.Y(_202_),
    .B(_187_),
    .A_N(_201_));
 sg13g2_a22oi_1 _621_ (.Y(_003_),
    .B1(_202_),
    .B2(net127),
    .A2(_200_),
    .A1(_162_));
 sg13g2_nand2_1 _622_ (.Y(_203_),
    .A(net135),
    .B(net131));
 sg13g2_a21oi_1 _623_ (.A1(net136),
    .A2(net131),
    .Y(_204_),
    .B1(net143));
 sg13g2_a22oi_1 _624_ (.Y(_205_),
    .B1(_204_),
    .B2(_166_),
    .A2(_168_),
    .A1(net143));
 sg13g2_a21o_1 _625_ (.A2(net131),
    .A1(net139),
    .B1(_142_),
    .X(_206_));
 sg13g2_nand2b_1 _626_ (.Y(_207_),
    .B(net150),
    .A_N(_206_));
 sg13g2_nand2b_1 _627_ (.Y(_208_),
    .B(net149),
    .A_N(_205_));
 sg13g2_a21oi_1 _628_ (.A1(_205_),
    .A2(_207_),
    .Y(_209_),
    .B1(net129));
 sg13g2_a21oi_1 _629_ (.A1(net145),
    .A2(_134_),
    .Y(_210_),
    .B1(net140));
 sg13g2_nor2_1 _630_ (.A(_159_),
    .B(_210_),
    .Y(_211_));
 sg13g2_nand2_1 _631_ (.Y(_212_),
    .A(_144_),
    .B(_198_));
 sg13g2_or2_1 _632_ (.X(_213_),
    .B(_211_),
    .A(_172_));
 sg13g2_a21o_1 _633_ (.A2(_212_),
    .A1(_211_),
    .B1(_172_),
    .X(_214_));
 sg13g2_nand3_1 _634_ (.B(net136),
    .C(_168_),
    .A(net143),
    .Y(_215_));
 sg13g2_nand3_1 _635_ (.B(_185_),
    .C(_215_),
    .A(net147),
    .Y(_216_));
 sg13g2_a221oi_1 _636_ (.B2(_216_),
    .C1(net128),
    .B1(_214_),
    .A1(_208_),
    .Y(_217_),
    .A2(_209_));
 sg13g2_nand2_2 _637_ (.Y(_218_),
    .A(net128),
    .B(net130));
 sg13g2_a221oi_1 _638_ (.B2(_142_),
    .C1(_147_),
    .B1(net137),
    .A1(_118_),
    .Y(_219_),
    .A2(_119_));
 sg13g2_a21oi_1 _639_ (.A1(_144_),
    .A2(_198_),
    .Y(_220_),
    .B1(_219_));
 sg13g2_nor2_1 _640_ (.A(net151),
    .B(_175_),
    .Y(_221_));
 sg13g2_xor2_1 _641_ (.B(_221_),
    .A(_220_),
    .X(_222_));
 sg13g2_nor2_1 _642_ (.A(_218_),
    .B(_222_),
    .Y(_223_));
 sg13g2_or3_1 _643_ (.A(_189_),
    .B(_217_),
    .C(_223_),
    .X(_004_));
 sg13g2_a21oi_2 _644_ (.B1(_134_),
    .Y(_224_),
    .A2(net134),
    .A1(net140));
 sg13g2_o21ai_1 _645_ (.B1(_167_),
    .Y(_225_),
    .A1(net143),
    .A2(_224_));
 sg13g2_a21oi_1 _646_ (.A1(net143),
    .A2(_168_),
    .Y(_226_),
    .B1(net149));
 sg13g2_nand2_1 _647_ (.Y(_227_),
    .A(_225_),
    .B(_226_));
 sg13g2_a21oi_1 _648_ (.A1(net142),
    .A2(_146_),
    .Y(_228_),
    .B1(net150));
 sg13g2_nor3_1 _649_ (.A(net141),
    .B(_169_),
    .C(_224_),
    .Y(_229_));
 sg13g2_nand2b_1 _650_ (.Y(_230_),
    .B(_228_),
    .A_N(_229_));
 sg13g2_nor2_1 _651_ (.A(net147),
    .B(_169_),
    .Y(_231_));
 sg13g2_a21oi_1 _652_ (.A1(_171_),
    .A2(_231_),
    .Y(_232_),
    .B1(net129));
 sg13g2_a221oi_1 _653_ (.B2(_232_),
    .C1(net128),
    .B1(_230_),
    .A1(_214_),
    .Y(_233_),
    .A2(_227_));
 sg13g2_a21o_1 _654_ (.A2(_147_),
    .A1(net131),
    .B1(_220_),
    .X(_234_));
 sg13g2_a21oi_2 _655_ (.B1(net135),
    .Y(_235_),
    .A2(_140_),
    .A1(net137));
 sg13g2_nand3_1 _656_ (.B(_146_),
    .C(_235_),
    .A(net142),
    .Y(_236_));
 sg13g2_a21oi_1 _657_ (.A1(_154_),
    .A2(_177_),
    .Y(_237_),
    .B1(net151));
 sg13g2_a221oi_1 _658_ (.B2(_237_),
    .C1(_218_),
    .B1(_236_),
    .A1(net151),
    .Y(_238_),
    .A2(_234_));
 sg13g2_nand2_1 _659_ (.Y(_239_),
    .A(net133),
    .B(_189_));
 sg13g2_inv_1 _660_ (.Y(_240_),
    .A(_239_));
 sg13g2_or3_1 _661_ (.A(_233_),
    .B(_238_),
    .C(_240_),
    .X(_005_));
 sg13g2_a21oi_2 _662_ (.B1(net146),
    .Y(_241_),
    .A2(net133),
    .A1(net137));
 sg13g2_a22oi_1 _663_ (.Y(_242_),
    .B1(_241_),
    .B2(_166_),
    .A2(_177_),
    .A1(_147_));
 sg13g2_or2_1 _664_ (.X(_243_),
    .B(_242_),
    .A(net151));
 sg13g2_a21o_1 _665_ (.A2(_224_),
    .A1(_170_),
    .B1(net142),
    .X(_244_));
 sg13g2_nor3_1 _666_ (.A(net148),
    .B(_145_),
    .C(_235_),
    .Y(_245_));
 sg13g2_and2_1 _667_ (.A(net126),
    .B(_235_),
    .X(_246_));
 sg13g2_a21oi_1 _668_ (.A1(_244_),
    .A2(_245_),
    .Y(_247_),
    .B1(_246_));
 sg13g2_a21oi_1 _669_ (.A1(_243_),
    .A2(_247_),
    .Y(_248_),
    .B1(_218_));
 sg13g2_nor4_1 _670_ (.A(net145),
    .B(_136_),
    .C(_138_),
    .D(_175_),
    .Y(_249_));
 sg13g2_a21o_1 _671_ (.A2(_175_),
    .A1(net145),
    .B1(net151),
    .X(_250_));
 sg13g2_a22oi_1 _672_ (.Y(_251_),
    .B1(_153_),
    .B2(net126),
    .A2(_148_),
    .A1(net151));
 sg13g2_o21ai_1 _673_ (.B1(_251_),
    .Y(_252_),
    .A1(_249_),
    .A2(_250_));
 sg13g2_o21ai_1 _674_ (.B1(_192_),
    .Y(_253_),
    .A1(net135),
    .A2(_146_));
 sg13g2_o21ai_1 _675_ (.B1(net148),
    .Y(_254_),
    .A1(_241_),
    .A2(_253_));
 sg13g2_a221oi_1 _676_ (.B2(_213_),
    .C1(net128),
    .B1(_254_),
    .A1(_159_),
    .Y(_255_),
    .A2(_252_));
 sg13g2_or3_1 _677_ (.A(_189_),
    .B(_248_),
    .C(_255_),
    .X(_006_));
 sg13g2_or3_1 _678_ (.A(net145),
    .B(net137),
    .C(_142_),
    .X(_256_));
 sg13g2_nand3_1 _679_ (.B(net137),
    .C(net132),
    .A(net145),
    .Y(_257_));
 sg13g2_nand3_1 _680_ (.B(_256_),
    .C(_257_),
    .A(net147),
    .Y(_258_));
 sg13g2_nor3_1 _681_ (.A(net147),
    .B(net133),
    .C(_147_),
    .Y(_259_));
 sg13g2_a22oi_1 _682_ (.Y(_260_),
    .B1(_259_),
    .B2(_151_),
    .A2(_166_),
    .A1(_122_));
 sg13g2_a21oi_1 _683_ (.A1(_258_),
    .A2(_260_),
    .Y(_261_),
    .B1(net130));
 sg13g2_nor3_1 _684_ (.A(net143),
    .B(_169_),
    .C(_224_),
    .Y(_262_));
 sg13g2_o21ai_1 _685_ (.B1(_172_),
    .Y(_263_),
    .A1(net141),
    .A2(_235_));
 sg13g2_o21ai_1 _686_ (.B1(_110_),
    .Y(_264_),
    .A1(_262_),
    .A2(_263_));
 sg13g2_a221oi_1 _687_ (.B2(_144_),
    .C1(_159_),
    .B1(_198_),
    .A1(_143_),
    .Y(_265_),
    .A2(_184_));
 sg13g2_and3_1 _688_ (.X(_266_),
    .A(net152),
    .B(_192_),
    .C(_265_));
 sg13g2_nor3_1 _689_ (.A(_261_),
    .B(_264_),
    .C(_266_),
    .Y(_267_));
 sg13g2_a21o_1 _690_ (.A2(_236_),
    .A1(_192_),
    .B1(net151),
    .X(_268_));
 sg13g2_a22oi_1 _691_ (.Y(_269_),
    .B1(_246_),
    .B2(_146_),
    .A2(_219_),
    .A1(net152));
 sg13g2_a21oi_1 _692_ (.A1(_268_),
    .A2(_269_),
    .Y(_270_),
    .B1(_218_));
 sg13g2_or3_1 _693_ (.A(_240_),
    .B(_267_),
    .C(_270_),
    .X(_007_));
 sg13g2_and2_1 _694_ (.A(_152_),
    .B(_241_),
    .X(_271_));
 sg13g2_a221oi_1 _695_ (.B2(_224_),
    .C1(net142),
    .B1(_170_),
    .A1(_134_),
    .Y(_272_),
    .A2(net133));
 sg13g2_o21ai_1 _696_ (.B1(net148),
    .Y(_273_),
    .A1(_271_),
    .A2(_272_));
 sg13g2_nor3_1 _697_ (.A(_150_),
    .B(_153_),
    .C(_164_),
    .Y(_274_));
 sg13g2_nor3_1 _698_ (.A(_123_),
    .B(net138),
    .C(_142_),
    .Y(_275_));
 sg13g2_nor3_1 _699_ (.A(net130),
    .B(_274_),
    .C(_275_),
    .Y(_276_));
 sg13g2_o21ai_1 _700_ (.B1(net142),
    .Y(_277_),
    .A1(net140),
    .A2(_135_));
 sg13g2_a21oi_1 _701_ (.A1(_170_),
    .A2(_224_),
    .Y(_278_),
    .B1(_277_));
 sg13g2_o21ai_1 _702_ (.B1(net144),
    .Y(_279_),
    .A1(net138),
    .A2(net134));
 sg13g2_nor2_1 _703_ (.A(_164_),
    .B(_279_),
    .Y(_280_));
 sg13g2_o21ai_1 _704_ (.B1(net148),
    .Y(_281_),
    .A1(_278_),
    .A2(_280_));
 sg13g2_a221oi_1 _705_ (.B2(_213_),
    .C1(net128),
    .B1(_281_),
    .A1(_273_),
    .Y(_282_),
    .A2(_276_));
 sg13g2_or2_1 _706_ (.X(_283_),
    .B(_166_),
    .A(net146));
 sg13g2_a21oi_1 _707_ (.A1(_212_),
    .A2(_283_),
    .Y(_284_),
    .B1(net150));
 sg13g2_nor3_1 _708_ (.A(_123_),
    .B(_145_),
    .C(_235_),
    .Y(_285_));
 sg13g2_a21oi_1 _709_ (.A1(net136),
    .A2(_168_),
    .Y(_286_),
    .B1(_150_));
 sg13g2_nor4_1 _710_ (.A(_218_),
    .B(_284_),
    .C(_285_),
    .D(_286_),
    .Y(_287_));
 sg13g2_or3_1 _711_ (.A(_189_),
    .B(_282_),
    .C(_287_),
    .X(_008_));
 sg13g2_o21ai_1 _712_ (.B1(net147),
    .Y(_288_),
    .A1(_165_),
    .A2(_198_));
 sg13g2_o21ai_1 _713_ (.B1(_149_),
    .Y(_289_),
    .A1(_145_),
    .A2(_235_));
 sg13g2_nand2_1 _714_ (.Y(_290_),
    .A(net134),
    .B(_147_));
 sg13g2_a21oi_1 _715_ (.A1(net126),
    .A2(_290_),
    .Y(_291_),
    .B1(_218_));
 sg13g2_nand3_1 _716_ (.B(_289_),
    .C(_291_),
    .A(_288_),
    .Y(_292_));
 sg13g2_a22oi_1 _717_ (.Y(_293_),
    .B1(_169_),
    .B2(net136),
    .A2(_168_),
    .A1(net141));
 sg13g2_a21oi_1 _718_ (.A1(_183_),
    .A2(_293_),
    .Y(_294_),
    .B1(net149));
 sg13g2_a21o_1 _719_ (.A2(_206_),
    .A1(net126),
    .B1(net129),
    .X(_295_));
 sg13g2_nor3_1 _720_ (.A(_274_),
    .B(_294_),
    .C(_295_),
    .Y(_296_));
 sg13g2_nand2_1 _721_ (.Y(_297_),
    .A(_153_),
    .B(_177_));
 sg13g2_a21oi_1 _722_ (.A1(_149_),
    .A2(_169_),
    .Y(_298_),
    .B1(_159_));
 sg13g2_a22oi_1 _723_ (.Y(_299_),
    .B1(_228_),
    .B2(_297_),
    .A2(_145_),
    .A1(net126));
 sg13g2_a21o_1 _724_ (.A2(_299_),
    .A1(_298_),
    .B1(net127),
    .X(_300_));
 sg13g2_o21ai_1 _725_ (.B1(_292_),
    .Y(_009_),
    .A1(_296_),
    .A2(_300_));
 sg13g2_a21o_1 _726_ (.A2(_199_),
    .A1(_176_),
    .B1(net149),
    .X(_301_));
 sg13g2_nand2b_1 _727_ (.Y(_302_),
    .B(_166_),
    .A_N(_163_));
 sg13g2_a21o_1 _728_ (.A2(_257_),
    .A1(_160_),
    .B1(_163_),
    .X(_303_));
 sg13g2_a21oi_1 _729_ (.A1(_184_),
    .A2(_203_),
    .Y(_304_),
    .B1(net150));
 sg13g2_a221oi_1 _730_ (.B2(_304_),
    .C1(_295_),
    .B1(_303_),
    .A1(_149_),
    .Y(_305_),
    .A2(_302_));
 sg13g2_a21o_1 _731_ (.A2(_301_),
    .A1(_265_),
    .B1(net127),
    .X(_306_));
 sg13g2_nand2b_1 _732_ (.Y(_307_),
    .B(_198_),
    .A_N(_175_));
 sg13g2_a21o_1 _733_ (.A2(_307_),
    .A1(_283_),
    .B1(net151),
    .X(_308_));
 sg13g2_o21ai_1 _734_ (.B1(net133),
    .Y(_309_),
    .A1(net140),
    .A2(_134_));
 sg13g2_a21oi_1 _735_ (.A1(_277_),
    .A2(_309_),
    .Y(_310_),
    .B1(net148));
 sg13g2_nor2_1 _736_ (.A(_218_),
    .B(_310_),
    .Y(_311_));
 sg13g2_a21oi_1 _737_ (.A1(_308_),
    .A2(_311_),
    .Y(_312_),
    .B1(_189_));
 sg13g2_o21ai_1 _738_ (.B1(_312_),
    .Y(_001_),
    .A1(_305_),
    .A2(_306_));
 sg13g2_nor3_1 _739_ (.A(_123_),
    .B(net129),
    .C(_290_),
    .Y(_313_));
 sg13g2_nor2_1 _740_ (.A(_196_),
    .B(_313_),
    .Y(_314_));
 sg13g2_nor2_1 _741_ (.A(_110_),
    .B(_314_),
    .Y(_020_));
 sg13g2_nor2_1 _742_ (.A(net127),
    .B(_314_),
    .Y(_021_));
 sg13g2_and2_1 _743_ (.A(net67),
    .B(net158),
    .X(_022_));
 sg13g2_xor2_1 _744_ (.B(net171),
    .A(\ticks[0] ),
    .X(_315_));
 sg13g2_nor2_1 _745_ (.A(net154),
    .B(net172),
    .Y(_023_));
 sg13g2_o21ai_1 _746_ (.B1(net182),
    .Y(_316_),
    .A1(\ticks[0] ),
    .A2(net171));
 sg13g2_nor2b_1 _747_ (.A(net183),
    .B_N(_316_),
    .Y(_317_));
 sg13g2_nor2_1 _748_ (.A(net154),
    .B(net184),
    .Y(_024_));
 sg13g2_nand2b_1 _749_ (.Y(_318_),
    .B(net106),
    .A_N(_081_));
 sg13g2_a21oi_1 _750_ (.A1(_083_),
    .A2(_318_),
    .Y(_025_),
    .B1(net154));
 sg13g2_xnor2_1 _751_ (.Y(_319_),
    .A(net115),
    .B(_082_));
 sg13g2_nor2_1 _752_ (.A(net153),
    .B(net116),
    .Y(_026_));
 sg13g2_o21ai_1 _753_ (.B1(net90),
    .Y(_320_),
    .A1(\ticks[4] ),
    .A2(_083_));
 sg13g2_a21oi_1 _754_ (.A1(_085_),
    .A2(net91),
    .Y(_027_),
    .B1(net153));
 sg13g2_xor2_1 _755_ (.B(_085_),
    .A(net176),
    .X(_321_));
 sg13g2_nor2_1 _756_ (.A(net153),
    .B(net177),
    .Y(_028_));
 sg13g2_o21ai_1 _757_ (.B1(net85),
    .Y(_322_),
    .A1(\ticks[6] ),
    .A2(_085_));
 sg13g2_a21oi_1 _758_ (.A1(_087_),
    .A2(net86),
    .Y(_029_),
    .B1(net153));
 sg13g2_xor2_1 _759_ (.B(_087_),
    .A(net178),
    .X(_323_));
 sg13g2_nor2_1 _760_ (.A(net153),
    .B(_323_),
    .Y(_030_));
 sg13g2_o21ai_1 _761_ (.B1(net93),
    .Y(_324_),
    .A1(\ticks[8] ),
    .A2(_087_));
 sg13g2_or3_1 _762_ (.A(net93),
    .B(\ticks[8] ),
    .C(_087_),
    .X(_325_));
 sg13g2_a21oi_1 _763_ (.A1(net94),
    .A2(_325_),
    .Y(_031_),
    .B1(net153));
 sg13g2_xor2_1 _764_ (.B(_325_),
    .A(net175),
    .X(_326_));
 sg13g2_nor2_1 _765_ (.A(net153),
    .B(_326_),
    .Y(_032_));
 sg13g2_o21ai_1 _766_ (.B1(net79),
    .Y(_327_),
    .A1(\ticks[10] ),
    .A2(_325_));
 sg13g2_a21oi_1 _767_ (.A1(_089_),
    .A2(net80),
    .Y(_033_),
    .B1(net153));
 sg13g2_a21oi_1 _768_ (.A1(_075_),
    .A2(net161),
    .Y(_034_),
    .B1(_125_));
 sg13g2_nand2_1 _769_ (.Y(_328_),
    .A(net113),
    .B(net158));
 sg13g2_o21ai_1 _770_ (.B1(_328_),
    .Y(_035_),
    .A1(_076_),
    .A2(_137_));
 sg13g2_o21ai_1 _771_ (.B1(_131_),
    .Y(_036_),
    .A1(_074_),
    .A2(net155));
 sg13g2_o21ai_1 _772_ (.B1(_118_),
    .Y(_037_),
    .A1(_073_),
    .A2(net155));
 sg13g2_a21o_1 _773_ (.A2(net158),
    .A1(net112),
    .B1(_113_),
    .X(_038_));
 sg13g2_o21ai_1 _774_ (.B1(_157_),
    .Y(_039_),
    .A1(_071_),
    .A2(net154));
 sg13g2_o21ai_1 _775_ (.B1(_106_),
    .Y(_040_),
    .A1(_070_),
    .A2(net155));
 sg13g2_nand3_1 _776_ (.B(net168),
    .C(net164),
    .A(\db_entry[4] ),
    .Y(_329_));
 sg13g2_o21ai_1 _777_ (.B1(_329_),
    .Y(_041_),
    .A1(_069_),
    .A2(net156));
 sg13g2_nand3_1 _778_ (.B(net1),
    .C(net164),
    .A(net104),
    .Y(_330_));
 sg13g2_o21ai_1 _779_ (.B1(_330_),
    .Y(_042_),
    .A1(_068_),
    .A2(net157));
 sg13g2_nand3_1 _780_ (.B(net168),
    .C(net164),
    .A(net88),
    .Y(_331_));
 sg13g2_o21ai_1 _781_ (.B1(_331_),
    .Y(_043_),
    .A1(_067_),
    .A2(net157));
 sg13g2_nand3_1 _782_ (.B(net168),
    .C(net164),
    .A(net74),
    .Y(_332_));
 sg13g2_o21ai_1 _783_ (.B1(_332_),
    .Y(_044_),
    .A1(_066_),
    .A2(net157));
 sg13g2_nand3_1 _784_ (.B(net168),
    .C(net165),
    .A(net169),
    .Y(_333_));
 sg13g2_o21ai_1 _785_ (.B1(_333_),
    .Y(_045_),
    .A1(_065_),
    .A2(net157));
 sg13g2_nand3_1 _786_ (.B(net167),
    .C(net164),
    .A(net98),
    .Y(_334_));
 sg13g2_o21ai_1 _787_ (.B1(_334_),
    .Y(_046_),
    .A1(_064_),
    .A2(net156));
 sg13g2_nand3_1 _788_ (.B(net167),
    .C(net164),
    .A(net72),
    .Y(_335_));
 sg13g2_o21ai_1 _789_ (.B1(_335_),
    .Y(_047_),
    .A1(_063_),
    .A2(net156));
 sg13g2_nand3_1 _790_ (.B(net167),
    .C(net164),
    .A(net70),
    .Y(_336_));
 sg13g2_o21ai_1 _791_ (.B1(_336_),
    .Y(_048_),
    .A1(_062_),
    .A2(net156));
 sg13g2_xnor2_1 _792_ (.Y(_337_),
    .A(\ticks[12] ),
    .B(_089_));
 sg13g2_o21ai_1 _793_ (.B1(net166),
    .Y(_338_),
    .A1(net108),
    .A2(net160));
 sg13g2_nor2b_1 _794_ (.A(_338_),
    .B_N(_337_),
    .Y(_049_));
 sg13g2_o21ai_1 _795_ (.B1(net117),
    .Y(_339_),
    .A1(\ticks[12] ),
    .A2(_089_));
 sg13g2_o21ai_1 _796_ (.B1(_090_),
    .Y(_340_),
    .A1(\db_entry[1] ),
    .A2(_091_));
 sg13g2_a21oi_1 _797_ (.A1(net118),
    .A2(_340_),
    .Y(_050_),
    .B1(_076_));
 sg13g2_and2_1 _798_ (.A(net180),
    .B(_090_),
    .X(_341_));
 sg13g2_nor2_1 _799_ (.A(net180),
    .B(_090_),
    .Y(_342_));
 sg13g2_a221oi_1 _800_ (.B2(_091_),
    .C1(_342_),
    .B1(_341_),
    .A1(\db_entry[2] ),
    .Y(_343_),
    .A2(net162));
 sg13g2_nor2_1 _801_ (.A(_076_),
    .B(net181),
    .Y(_051_));
 sg13g2_xnor2_1 _802_ (.Y(_344_),
    .A(\ticks[15] ),
    .B(_341_));
 sg13g2_o21ai_1 _803_ (.B1(net166),
    .Y(_345_),
    .A1(net102),
    .A2(net160));
 sg13g2_a21oi_1 _804_ (.A1(net160),
    .A2(_344_),
    .Y(_052_),
    .B1(_345_));
 sg13g2_nand2_1 _805_ (.Y(_346_),
    .A(_067_),
    .B(\counter[1] ));
 sg13g2_nor2_1 _806_ (.A(_068_),
    .B(\counter[0] ),
    .Y(_347_));
 sg13g2_nand2b_1 _807_ (.Y(_348_),
    .B(\freq[3] ),
    .A_N(\counter[2] ));
 sg13g2_o21ai_1 _808_ (.B1(_348_),
    .Y(_349_),
    .A1(_067_),
    .A2(\counter[1] ));
 sg13g2_a21oi_1 _809_ (.A1(_346_),
    .A2(_347_),
    .Y(_350_),
    .B1(_349_));
 sg13g2_a221oi_1 _810_ (.B2(_066_),
    .C1(_350_),
    .B1(\counter[2] ),
    .A1(_065_),
    .Y(_351_),
    .A2(\counter[3] ));
 sg13g2_nor2_1 _811_ (.A(_063_),
    .B(\counter[5] ),
    .Y(_352_));
 sg13g2_nor3_2 _812_ (.A(\counter[0] ),
    .B(\counter[2] ),
    .C(\counter[1] ),
    .Y(_353_));
 sg13g2_and2_1 _813_ (.A(_080_),
    .B(_353_),
    .X(_354_));
 sg13g2_and2_1 _814_ (.A(_079_),
    .B(_354_),
    .X(_355_));
 sg13g2_nor2b_1 _815_ (.A(\counter[5] ),
    .B_N(_355_),
    .Y(_356_));
 sg13g2_nor2b_2 _816_ (.A(\counter[6] ),
    .B_N(_356_),
    .Y(_357_));
 sg13g2_a221oi_1 _817_ (.B2(\freq[4] ),
    .C1(_351_),
    .B1(_080_),
    .A1(\freq[5] ),
    .Y(_358_),
    .A2(_079_));
 sg13g2_a221oi_1 _818_ (.B2(_064_),
    .C1(_358_),
    .B1(\counter[4] ),
    .A1(_063_),
    .Y(_359_),
    .A2(\counter[5] ));
 sg13g2_nor2_1 _819_ (.A(_062_),
    .B(\counter[6] ),
    .Y(_360_));
 sg13g2_nor4_1 _820_ (.A(_352_),
    .B(_357_),
    .C(_359_),
    .D(_360_),
    .Y(_361_));
 sg13g2_nor2b_1 _821_ (.A(\freq[7] ),
    .B_N(\counter[6] ),
    .Y(_362_));
 sg13g2_nor4_1 _822_ (.A(\counter[7] ),
    .B(net164),
    .C(_361_),
    .D(_362_),
    .Y(_363_));
 sg13g2_o21ai_1 _823_ (.B1(net167),
    .Y(_364_),
    .A1(net173),
    .A2(net161));
 sg13g2_nor2_1 _824_ (.A(_363_),
    .B(_364_),
    .Y(_053_));
 sg13g2_nand2b_2 _825_ (.Y(_365_),
    .B(_357_),
    .A_N(\counter[7] ));
 sg13g2_a21oi_1 _826_ (.A1(_107_),
    .A2(_365_),
    .Y(_366_),
    .B1(_041_));
 sg13g2_nor2b_1 _827_ (.A(net68),
    .B_N(_365_),
    .Y(_367_));
 sg13g2_a21oi_1 _828_ (.A1(_329_),
    .A2(_367_),
    .Y(_054_),
    .B1(_366_));
 sg13g2_xnor2_1 _829_ (.Y(_368_),
    .A(\counter[0] ),
    .B(\counter[1] ));
 sg13g2_o21ai_1 _830_ (.B1(_368_),
    .Y(_369_),
    .A1(net100),
    .A2(_365_));
 sg13g2_o21ai_1 _831_ (.B1(_330_),
    .Y(_055_),
    .A1(net157),
    .A2(_369_));
 sg13g2_o21ai_1 _832_ (.B1(\counter[2] ),
    .Y(_370_),
    .A1(\counter[0] ),
    .A2(\counter[1] ));
 sg13g2_nand2b_1 _833_ (.Y(_371_),
    .B(_370_),
    .A_N(_353_));
 sg13g2_o21ai_1 _834_ (.B1(_371_),
    .Y(_372_),
    .A1(net96),
    .A2(_365_));
 sg13g2_o21ai_1 _835_ (.B1(_331_),
    .Y(_056_),
    .A1(net157),
    .A2(net97));
 sg13g2_xnor2_1 _836_ (.Y(_373_),
    .A(_080_),
    .B(_353_));
 sg13g2_o21ai_1 _837_ (.B1(_373_),
    .Y(_374_),
    .A1(\freq[3] ),
    .A2(_365_));
 sg13g2_o21ai_1 _838_ (.B1(_332_),
    .Y(_057_),
    .A1(net156),
    .A2(_374_));
 sg13g2_a21oi_1 _839_ (.A1(net158),
    .A2(_365_),
    .Y(_375_),
    .B1(net123));
 sg13g2_xnor2_1 _840_ (.Y(_376_),
    .A(\counter[4] ),
    .B(_354_));
 sg13g2_a21oi_1 _841_ (.A1(_333_),
    .A2(_376_),
    .Y(_058_),
    .B1(_375_));
 sg13g2_a21oi_1 _842_ (.A1(net158),
    .A2(_365_),
    .Y(_377_),
    .B1(_046_));
 sg13g2_xnor2_1 _843_ (.Y(_378_),
    .A(\counter[5] ),
    .B(_355_));
 sg13g2_a21oi_1 _844_ (.A1(_334_),
    .A2(_378_),
    .Y(_059_),
    .B1(_377_));
 sg13g2_nor2b_1 _845_ (.A(_356_),
    .B_N(\counter[6] ),
    .Y(_379_));
 sg13g2_or2_1 _846_ (.X(_380_),
    .B(\counter[7] ),
    .A(\freq[6] ));
 sg13g2_a21oi_1 _847_ (.A1(_357_),
    .A2(_380_),
    .Y(_381_),
    .B1(_379_));
 sg13g2_o21ai_1 _848_ (.B1(_335_),
    .Y(_060_),
    .A1(net156),
    .A2(_381_));
 sg13g2_nand2b_1 _849_ (.Y(_382_),
    .B(net185),
    .A_N(_357_));
 sg13g2_nor3_1 _850_ (.A(_062_),
    .B(net156),
    .C(_365_),
    .Y(_383_));
 sg13g2_o21ai_1 _851_ (.B1(_336_),
    .Y(_384_),
    .A1(net156),
    .A2(_382_));
 sg13g2_or2_1 _852_ (.X(_061_),
    .B(_384_),
    .A(_383_));
 sg13g2_dfrbp_1 _853_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net9),
    .D(_020_),
    .Q_N(_416_),
    .Q(\db_entry[3] ));
 sg13g2_dfrbp_1 _854_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net10),
    .D(_000_),
    .Q_N(_417_),
    .Q(\db_entry[0] ));
 sg13g2_dfrbp_1 _855_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net11),
    .D(_002_),
    .Q_N(_418_),
    .Q(\db_entry[1] ));
 sg13g2_dfrbp_1 _856_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net12),
    .D(_003_),
    .Q_N(_419_),
    .Q(\db_entry[2] ));
 sg13g2_dfrbp_1 _857_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net13),
    .D(_004_),
    .Q_N(_420_),
    .Q(\db_entry[4] ));
 sg13g2_dfrbp_1 _858_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net14),
    .D(_005_),
    .Q_N(_421_),
    .Q(\db_entry[5] ));
 sg13g2_dfrbp_1 _859_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net15),
    .D(_006_),
    .Q_N(_422_),
    .Q(\db_entry[6] ));
 sg13g2_dfrbp_1 _860_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net16),
    .D(_007_),
    .Q_N(_423_),
    .Q(\db_entry[7] ));
 sg13g2_dfrbp_1 _861_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net17),
    .D(_008_),
    .Q_N(_424_),
    .Q(\db_entry[8] ));
 sg13g2_dfrbp_1 _862_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net36),
    .D(_009_),
    .Q_N(_425_),
    .Q(\db_entry[9] ));
 sg13g2_dfrbp_1 _863_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net8),
    .D(_001_),
    .Q_N(_415_),
    .Q(\db_entry[10] ));
 sg13g2_dfrbp_1 _864_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net20),
    .D(_021_),
    .Q_N(_414_),
    .Q(\db_entry[11] ));
 sg13g2_dfrbp_1 _865_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net19),
    .D(_022_),
    .Q_N(_019_),
    .Q(\ticks[0] ));
 sg13g2_dfrbp_1 _866_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net18),
    .D(_023_),
    .Q_N(_413_),
    .Q(\ticks[1] ));
 sg13g2_dfrbp_1 _867_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net7),
    .D(_024_),
    .Q_N(_412_),
    .Q(\ticks[2] ));
 sg13g2_dfrbp_1 _868_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net58),
    .D(net107),
    .Q_N(_411_),
    .Q(\ticks[3] ));
 sg13g2_dfrbp_1 _869_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net57),
    .D(_026_),
    .Q_N(_410_),
    .Q(\ticks[4] ));
 sg13g2_dfrbp_1 _870_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net56),
    .D(net92),
    .Q_N(_409_),
    .Q(\ticks[5] ));
 sg13g2_dfrbp_1 _871_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net55),
    .D(_028_),
    .Q_N(_408_),
    .Q(\ticks[6] ));
 sg13g2_dfrbp_1 _872_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net54),
    .D(net87),
    .Q_N(_407_),
    .Q(\ticks[7] ));
 sg13g2_dfrbp_1 _873_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net53),
    .D(_030_),
    .Q_N(_406_),
    .Q(\ticks[8] ));
 sg13g2_dfrbp_1 _874_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net52),
    .D(net95),
    .Q_N(_405_),
    .Q(\ticks[9] ));
 sg13g2_dfrbp_1 _875_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net51),
    .D(_032_),
    .Q_N(_404_),
    .Q(\ticks[10] ));
 sg13g2_dfrbp_1 _876_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net50),
    .D(net81),
    .Q_N(_403_),
    .Q(\ticks[11] ));
 sg13g2_dfrbp_1 _877_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net49),
    .D(_034_),
    .Q_N(_013_),
    .Q(\meriac_tune_db.address[0] ));
 sg13g2_dfrbp_1 _878_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net47),
    .D(net114),
    .Q_N(_014_),
    .Q(\meriac_tune_db.address[1] ));
 sg13g2_dfrbp_1 _879_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net45),
    .D(_036_),
    .Q_N(_015_),
    .Q(\meriac_tune_db.address[2] ));
 sg13g2_dfrbp_1 _880_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net43),
    .D(net121),
    .Q_N(_016_),
    .Q(\meriac_tune_db.address[3] ));
 sg13g2_dfrbp_1 _881_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net41),
    .D(_038_),
    .Q_N(_017_),
    .Q(\meriac_tune_db.address[4] ));
 sg13g2_dfrbp_1 _882_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net39),
    .D(net125),
    .Q_N(_011_),
    .Q(\meriac_tune_db.address[5] ));
 sg13g2_dfrbp_1 _883_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net37),
    .D(net78),
    .Q_N(_010_),
    .Q(\meriac_tune_db.address[6] ));
 sg13g2_dfrbp_1 _884_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net35),
    .D(net84),
    .Q_N(_402_),
    .Q(\freq[0] ));
 sg13g2_dfrbp_1 _885_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net33),
    .D(net101),
    .Q_N(_401_),
    .Q(\freq[1] ));
 sg13g2_dfrbp_1 _886_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net31),
    .D(net89),
    .Q_N(_400_),
    .Q(\freq[2] ));
 sg13g2_dfrbp_1 _887_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net29),
    .D(_044_),
    .Q_N(_399_),
    .Q(\freq[3] ));
 sg13g2_dfrbp_1 _888_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net27),
    .D(net123),
    .Q_N(_398_),
    .Q(\freq[4] ));
 sg13g2_dfrbp_1 _889_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net25),
    .D(_046_),
    .Q_N(_397_),
    .Q(\freq[5] ));
 sg13g2_dfrbp_1 _890_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net23),
    .D(_047_),
    .Q_N(_396_),
    .Q(\freq[6] ));
 sg13g2_dfrbp_1 _891_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net21),
    .D(net71),
    .Q_N(_395_),
    .Q(\freq[7] ));
 sg13g2_dfrbp_1 _892_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net46),
    .D(net109),
    .Q_N(_394_),
    .Q(\ticks[12] ));
 sg13g2_dfrbp_1 _893_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net44),
    .D(net119),
    .Q_N(_393_),
    .Q(\ticks[13] ));
 sg13g2_dfrbp_1 _894_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net42),
    .D(_051_),
    .Q_N(_012_),
    .Q(\ticks[14] ));
 sg13g2_dfrbp_1 _895_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net40),
    .D(net103),
    .Q_N(_392_),
    .Q(\ticks[15] ));
 sg13g2_dfrbp_1 _896_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net38),
    .D(net174),
    .Q_N(uio_out[1]),
    .Q(speaker));
 sg13g2_dfrbp_1 _897_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net34),
    .D(net69),
    .Q_N(_018_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 _898_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net32),
    .D(net105),
    .Q_N(_391_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 _899_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net30),
    .D(_056_),
    .Q_N(_390_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 _900_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net28),
    .D(net75),
    .Q_N(_389_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 _901_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net26),
    .D(net170),
    .Q_N(_388_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 _902_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net24),
    .D(net99),
    .Q_N(_387_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 _903_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net22),
    .D(net73),
    .Q_N(_386_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 _904_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net48),
    .D(net186),
    .Q_N(_385_),
    .Q(\counter[7] ));
 sg13g2_tiehi _863__8 (.L_HI(net8));
 sg13g2_tiehi _853__9 (.L_HI(net9));
 sg13g2_tiehi _854__10 (.L_HI(net10));
 sg13g2_tiehi _855__11 (.L_HI(net11));
 sg13g2_tiehi _856__12 (.L_HI(net12));
 sg13g2_tiehi _857__13 (.L_HI(net13));
 sg13g2_tiehi _858__14 (.L_HI(net14));
 sg13g2_tiehi _859__15 (.L_HI(net15));
 sg13g2_tiehi _860__16 (.L_HI(net16));
 sg13g2_tiehi _861__17 (.L_HI(net17));
 sg13g2_tiehi _866__18 (.L_HI(net18));
 sg13g2_tiehi _865__19 (.L_HI(net19));
 sg13g2_tiehi _864__20 (.L_HI(net20));
 sg13g2_tiehi _891__21 (.L_HI(net21));
 sg13g2_tiehi _903__22 (.L_HI(net22));
 sg13g2_tiehi _890__23 (.L_HI(net23));
 sg13g2_tiehi _902__24 (.L_HI(net24));
 sg13g2_tiehi _889__25 (.L_HI(net25));
 sg13g2_tiehi _901__26 (.L_HI(net26));
 sg13g2_tiehi _888__27 (.L_HI(net27));
 sg13g2_tiehi _900__28 (.L_HI(net28));
 sg13g2_tiehi _887__29 (.L_HI(net29));
 sg13g2_tiehi _899__30 (.L_HI(net30));
 sg13g2_tiehi _886__31 (.L_HI(net31));
 sg13g2_tiehi _898__32 (.L_HI(net32));
 sg13g2_tiehi _885__33 (.L_HI(net33));
 sg13g2_tiehi _897__34 (.L_HI(net34));
 sg13g2_tiehi _884__35 (.L_HI(net35));
 sg13g2_tiehi _862__36 (.L_HI(net36));
 sg13g2_tiehi _883__37 (.L_HI(net37));
 sg13g2_tiehi _896__38 (.L_HI(net38));
 sg13g2_tiehi _882__39 (.L_HI(net39));
 sg13g2_tiehi _895__40 (.L_HI(net40));
 sg13g2_tiehi _881__41 (.L_HI(net41));
 sg13g2_tiehi _894__42 (.L_HI(net42));
 sg13g2_tiehi _880__43 (.L_HI(net43));
 sg13g2_tiehi _893__44 (.L_HI(net44));
 sg13g2_tiehi _879__45 (.L_HI(net45));
 sg13g2_tiehi _892__46 (.L_HI(net46));
 sg13g2_tiehi _878__47 (.L_HI(net47));
 sg13g2_tiehi _904__48 (.L_HI(net48));
 sg13g2_tiehi _877__49 (.L_HI(net49));
 sg13g2_tiehi _876__50 (.L_HI(net50));
 sg13g2_tiehi _875__51 (.L_HI(net51));
 sg13g2_tiehi _874__52 (.L_HI(net52));
 sg13g2_tiehi _873__53 (.L_HI(net53));
 sg13g2_tiehi _872__54 (.L_HI(net54));
 sg13g2_tiehi _871__55 (.L_HI(net55));
 sg13g2_tiehi _870__56 (.L_HI(net56));
 sg13g2_tiehi _869__57 (.L_HI(net57));
 sg13g2_tiehi _868__58 (.L_HI(net58));
 sg13g2_tiehi tt_um_meriac_play_tune_59 (.L_HI(net59));
 sg13g2_tiehi tt_um_meriac_play_tune_60 (.L_HI(net60));
 sg13g2_tiehi tt_um_meriac_play_tune_61 (.L_HI(net61));
 sg13g2_tiehi tt_um_meriac_play_tune_62 (.L_HI(net62));
 sg13g2_tiehi tt_um_meriac_play_tune_63 (.L_HI(net63));
 sg13g2_tiehi tt_um_meriac_play_tune_64 (.L_HI(net64));
 sg13g2_tiehi tt_um_meriac_play_tune_65 (.L_HI(net65));
 sg13g2_tiehi tt_um_meriac_play_tune_66 (.L_HI(net66));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_meriac_play_tune_3 (.L_LO(net3));
 sg13g2_tielo tt_um_meriac_play_tune_4 (.L_LO(net4));
 sg13g2_tielo tt_um_meriac_play_tune_5 (.L_LO(net5));
 sg13g2_tielo tt_um_meriac_play_tune_6 (.L_LO(net6));
 sg13g2_tiehi _867__7 (.L_HI(net7));
 sg13g2_buf_1 _970_ (.A(speaker),
    .X(uio_out[0]));
 sg13g2_buf_1 _971_ (.A(speaker),
    .X(uio_out[7]));
 sg13g2_buf_1 _972_ (.A(ui_in[0]),
    .X(uo_out[0]));
 sg13g2_buf_1 _973_ (.A(ui_in[1]),
    .X(uo_out[1]));
 sg13g2_buf_1 _974_ (.A(ui_in[2]),
    .X(uo_out[2]));
 sg13g2_buf_1 _975_ (.A(ui_in[3]),
    .X(uo_out[3]));
 sg13g2_buf_1 _976_ (.A(ui_in[4]),
    .X(uo_out[4]));
 sg13g2_buf_1 _977_ (.A(ui_in[5]),
    .X(uo_out[5]));
 sg13g2_buf_1 _978_ (.A(ui_in[6]),
    .X(uo_out[6]));
 sg13g2_buf_1 _979_ (.A(ui_in[7]),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout126 (.A(_122_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(net128),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_109_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(net130),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_158_),
    .X(net130));
 sg13g2_buf_4 fanout131 (.X(net131),
    .A(_141_));
 sg13g2_buf_1 fanout132 (.A(_141_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(net134),
    .X(net133));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(_140_));
 sg13g2_buf_2 fanout135 (.A(_135_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_135_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(net138),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_128_),
    .X(net138));
 sg13g2_buf_4 fanout139 (.X(net139),
    .A(_127_));
 sg13g2_buf_2 fanout140 (.A(_127_),
    .X(net140));
 sg13g2_buf_4 fanout141 (.X(net141),
    .A(net142));
 sg13g2_buf_2 fanout142 (.A(_121_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(net146),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(net146),
    .X(net145));
 sg13g2_buf_1 fanout146 (.A(_120_),
    .X(net146));
 sg13g2_buf_4 fanout147 (.X(net147),
    .A(_115_));
 sg13g2_buf_2 fanout148 (.A(_115_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(net150),
    .X(net149));
 sg13g2_buf_1 fanout150 (.A(net152),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(net152),
    .X(net151));
 sg13g2_buf_1 fanout152 (.A(_114_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(net155),
    .X(net153));
 sg13g2_buf_1 fanout154 (.A(net155),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_108_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_108_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_108_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_107_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_100_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(net161),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_093_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(net165),
    .X(net162));
 sg13g2_buf_1 fanout163 (.A(net165),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(net165),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_092_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(net167),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(net1),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(net1),
    .X(net168));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_tielo tt_um_meriac_play_tune_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_3_5__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_019_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold2 (.A(_018_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold3 (.A(_054_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold4 (.A(\db_entry[11] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold5 (.A(_048_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold6 (.A(\db_entry[10] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold7 (.A(_060_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold8 (.A(\db_entry[7] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold9 (.A(_057_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold10 (.A(\freq[3] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold11 (.A(\meriac_tune_db.address[6] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold12 (.A(_040_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold13 (.A(\ticks[11] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold14 (.A(_327_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold15 (.A(_033_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold16 (.A(\freq[6] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold17 (.A(\freq[0] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold18 (.A(_041_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold19 (.A(\ticks[7] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold20 (.A(_322_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold21 (.A(_029_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold22 (.A(\db_entry[6] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold23 (.A(_043_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold24 (.A(\ticks[5] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold25 (.A(_320_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold26 (.A(_027_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold27 (.A(\ticks[9] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold28 (.A(_324_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold29 (.A(_031_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold30 (.A(\freq[2] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold31 (.A(_372_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold32 (.A(\db_entry[9] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold33 (.A(_059_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold34 (.A(\freq[1] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold35 (.A(_042_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold36 (.A(\db_entry[3] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold37 (.A(_052_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold38 (.A(\db_entry[5] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold39 (.A(_055_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold40 (.A(\ticks[3] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold41 (.A(_025_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold42 (.A(\db_entry[0] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold43 (.A(_049_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold44 (.A(\freq[5] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold45 (.A(\meriac_tune_db.address[2] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold46 (.A(\meriac_tune_db.address[4] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold47 (.A(\meriac_tune_db.address[1] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold48 (.A(_035_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold49 (.A(\ticks[4] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold50 (.A(_319_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold51 (.A(\ticks[13] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold52 (.A(_339_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold53 (.A(_050_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold54 (.A(\meriac_tune_db.address[3] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold55 (.A(_037_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold56 (.A(\freq[4] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold57 (.A(_045_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold58 (.A(\meriac_tune_db.address[5] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold59 (.A(_039_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold60 (.A(\db_entry[8] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold61 (.A(_058_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold62 (.A(\ticks[1] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold63 (.A(_315_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold64 (.A(speaker),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold65 (.A(_053_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold66 (.A(\ticks[10] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold67 (.A(\ticks[6] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold68 (.A(_321_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold69 (.A(\ticks[8] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold70 (.A(\meriac_tune_db.address[0] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold71 (.A(_012_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold72 (.A(_343_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold73 (.A(\ticks[2] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold74 (.A(_081_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold75 (.A(_317_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold76 (.A(\counter[7] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold77 (.A(_061_),
    .X(net186));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_4 FILLER_15_240 ();
 sg13g2_fill_2 FILLER_15_254 ();
 sg13g2_decap_8 FILLER_15_260 ();
 sg13g2_decap_8 FILLER_15_267 ();
 sg13g2_decap_8 FILLER_15_274 ();
 sg13g2_decap_8 FILLER_15_281 ();
 sg13g2_decap_8 FILLER_15_288 ();
 sg13g2_decap_8 FILLER_15_295 ();
 sg13g2_decap_8 FILLER_15_302 ();
 sg13g2_decap_8 FILLER_15_309 ();
 sg13g2_decap_8 FILLER_15_316 ();
 sg13g2_decap_4 FILLER_15_323 ();
 sg13g2_fill_2 FILLER_15_327 ();
 sg13g2_fill_1 FILLER_15_345 ();
 sg13g2_decap_4 FILLER_15_355 ();
 sg13g2_fill_1 FILLER_15_359 ();
 sg13g2_decap_8 FILLER_15_373 ();
 sg13g2_decap_8 FILLER_15_380 ();
 sg13g2_decap_8 FILLER_15_387 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_fill_1 FILLER_16_210 ();
 sg13g2_decap_4 FILLER_16_215 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_4 FILLER_16_294 ();
 sg13g2_fill_1 FILLER_16_298 ();
 sg13g2_fill_2 FILLER_16_325 ();
 sg13g2_fill_1 FILLER_16_327 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_4 FILLER_17_140 ();
 sg13g2_fill_2 FILLER_17_144 ();
 sg13g2_decap_8 FILLER_17_150 ();
 sg13g2_decap_8 FILLER_17_157 ();
 sg13g2_decap_4 FILLER_17_164 ();
 sg13g2_fill_2 FILLER_17_172 ();
 sg13g2_decap_8 FILLER_17_283 ();
 sg13g2_decap_8 FILLER_17_290 ();
 sg13g2_decap_8 FILLER_17_297 ();
 sg13g2_decap_4 FILLER_17_304 ();
 sg13g2_fill_2 FILLER_17_308 ();
 sg13g2_fill_2 FILLER_17_374 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_4 FILLER_18_126 ();
 sg13g2_fill_1 FILLER_18_130 ();
 sg13g2_decap_8 FILLER_18_183 ();
 sg13g2_fill_2 FILLER_18_216 ();
 sg13g2_fill_1 FILLER_18_218 ();
 sg13g2_fill_2 FILLER_18_271 ();
 sg13g2_fill_1 FILLER_18_299 ();
 sg13g2_fill_2 FILLER_18_326 ();
 sg13g2_fill_1 FILLER_18_328 ();
 sg13g2_fill_1 FILLER_18_362 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_fill_2 FILLER_19_185 ();
 sg13g2_decap_4 FILLER_19_192 ();
 sg13g2_fill_1 FILLER_19_196 ();
 sg13g2_fill_2 FILLER_19_202 ();
 sg13g2_fill_2 FILLER_19_214 ();
 sg13g2_fill_2 FILLER_19_227 ();
 sg13g2_fill_2 FILLER_19_248 ();
 sg13g2_fill_1 FILLER_19_274 ();
 sg13g2_decap_4 FILLER_19_306 ();
 sg13g2_fill_1 FILLER_19_314 ();
 sg13g2_fill_1 FILLER_19_324 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_fill_1 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_157 ();
 sg13g2_decap_4 FILLER_20_164 ();
 sg13g2_fill_1 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_173 ();
 sg13g2_fill_2 FILLER_20_189 ();
 sg13g2_fill_1 FILLER_20_208 ();
 sg13g2_decap_4 FILLER_20_226 ();
 sg13g2_fill_2 FILLER_20_255 ();
 sg13g2_fill_1 FILLER_20_257 ();
 sg13g2_fill_1 FILLER_20_350 ();
 sg13g2_fill_1 FILLER_20_360 ();
 sg13g2_fill_2 FILLER_20_378 ();
 sg13g2_fill_1 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_4 FILLER_21_119 ();
 sg13g2_fill_2 FILLER_21_129 ();
 sg13g2_fill_2 FILLER_21_142 ();
 sg13g2_decap_8 FILLER_21_162 ();
 sg13g2_fill_2 FILLER_21_200 ();
 sg13g2_fill_1 FILLER_21_202 ();
 sg13g2_decap_8 FILLER_21_212 ();
 sg13g2_fill_1 FILLER_21_219 ();
 sg13g2_decap_8 FILLER_21_228 ();
 sg13g2_decap_8 FILLER_21_256 ();
 sg13g2_fill_1 FILLER_21_263 ();
 sg13g2_fill_2 FILLER_21_292 ();
 sg13g2_fill_2 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_fill_1 FILLER_22_132 ();
 sg13g2_decap_8 FILLER_22_139 ();
 sg13g2_fill_2 FILLER_22_146 ();
 sg13g2_decap_4 FILLER_22_153 ();
 sg13g2_fill_1 FILLER_22_157 ();
 sg13g2_fill_2 FILLER_22_188 ();
 sg13g2_fill_2 FILLER_22_198 ();
 sg13g2_fill_1 FILLER_22_200 ();
 sg13g2_decap_4 FILLER_22_207 ();
 sg13g2_fill_2 FILLER_22_221 ();
 sg13g2_fill_1 FILLER_22_223 ();
 sg13g2_decap_8 FILLER_22_232 ();
 sg13g2_fill_2 FILLER_22_239 ();
 sg13g2_fill_1 FILLER_22_241 ();
 sg13g2_decap_8 FILLER_22_260 ();
 sg13g2_decap_8 FILLER_22_267 ();
 sg13g2_decap_8 FILLER_22_296 ();
 sg13g2_fill_2 FILLER_22_323 ();
 sg13g2_fill_1 FILLER_22_325 ();
 sg13g2_fill_1 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_fill_1 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_fill_2 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_158 ();
 sg13g2_decap_4 FILLER_23_165 ();
 sg13g2_decap_4 FILLER_23_192 ();
 sg13g2_decap_4 FILLER_23_217 ();
 sg13g2_fill_1 FILLER_23_221 ();
 sg13g2_fill_2 FILLER_23_255 ();
 sg13g2_fill_1 FILLER_23_257 ();
 sg13g2_fill_2 FILLER_23_278 ();
 sg13g2_fill_1 FILLER_23_280 ();
 sg13g2_fill_1 FILLER_23_307 ();
 sg13g2_fill_1 FILLER_23_360 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_fill_1 FILLER_24_112 ();
 sg13g2_fill_2 FILLER_24_158 ();
 sg13g2_fill_2 FILLER_24_177 ();
 sg13g2_fill_2 FILLER_24_186 ();
 sg13g2_fill_2 FILLER_24_204 ();
 sg13g2_fill_1 FILLER_24_206 ();
 sg13g2_fill_2 FILLER_24_211 ();
 sg13g2_fill_1 FILLER_24_213 ();
 sg13g2_decap_8 FILLER_24_218 ();
 sg13g2_fill_1 FILLER_24_225 ();
 sg13g2_fill_2 FILLER_24_241 ();
 sg13g2_fill_1 FILLER_24_243 ();
 sg13g2_fill_1 FILLER_24_257 ();
 sg13g2_decap_4 FILLER_24_271 ();
 sg13g2_fill_1 FILLER_24_275 ();
 sg13g2_decap_8 FILLER_24_282 ();
 sg13g2_fill_2 FILLER_24_289 ();
 sg13g2_fill_1 FILLER_24_291 ();
 sg13g2_decap_4 FILLER_24_304 ();
 sg13g2_fill_1 FILLER_24_323 ();
 sg13g2_fill_1 FILLER_24_372 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_4 FILLER_25_105 ();
 sg13g2_fill_2 FILLER_25_109 ();
 sg13g2_fill_2 FILLER_25_130 ();
 sg13g2_decap_4 FILLER_25_136 ();
 sg13g2_decap_4 FILLER_25_151 ();
 sg13g2_fill_2 FILLER_25_167 ();
 sg13g2_fill_1 FILLER_25_169 ();
 sg13g2_fill_2 FILLER_25_188 ();
 sg13g2_fill_1 FILLER_25_190 ();
 sg13g2_fill_2 FILLER_25_216 ();
 sg13g2_fill_1 FILLER_25_218 ();
 sg13g2_decap_8 FILLER_25_248 ();
 sg13g2_decap_4 FILLER_25_265 ();
 sg13g2_fill_1 FILLER_25_278 ();
 sg13g2_decap_4 FILLER_25_307 ();
 sg13g2_fill_2 FILLER_25_311 ();
 sg13g2_fill_2 FILLER_25_347 ();
 sg13g2_fill_1 FILLER_25_366 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_4 FILLER_26_98 ();
 sg13g2_fill_2 FILLER_26_102 ();
 sg13g2_decap_4 FILLER_26_130 ();
 sg13g2_decap_8 FILLER_26_158 ();
 sg13g2_decap_8 FILLER_26_165 ();
 sg13g2_decap_4 FILLER_26_172 ();
 sg13g2_fill_1 FILLER_26_176 ();
 sg13g2_fill_2 FILLER_26_186 ();
 sg13g2_fill_1 FILLER_26_188 ();
 sg13g2_fill_1 FILLER_26_199 ();
 sg13g2_fill_2 FILLER_26_205 ();
 sg13g2_fill_1 FILLER_26_207 ();
 sg13g2_fill_2 FILLER_26_214 ();
 sg13g2_decap_8 FILLER_26_221 ();
 sg13g2_fill_1 FILLER_26_234 ();
 sg13g2_decap_4 FILLER_26_262 ();
 sg13g2_decap_4 FILLER_26_286 ();
 sg13g2_fill_2 FILLER_26_290 ();
 sg13g2_fill_2 FILLER_26_315 ();
 sg13g2_fill_1 FILLER_26_317 ();
 sg13g2_fill_1 FILLER_26_332 ();
 sg13g2_fill_2 FILLER_26_345 ();
 sg13g2_fill_1 FILLER_26_347 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_fill_2 FILLER_27_105 ();
 sg13g2_fill_1 FILLER_27_107 ();
 sg13g2_fill_2 FILLER_27_131 ();
 sg13g2_fill_1 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_157 ();
 sg13g2_fill_2 FILLER_27_175 ();
 sg13g2_fill_2 FILLER_27_193 ();
 sg13g2_decap_8 FILLER_27_202 ();
 sg13g2_decap_4 FILLER_27_209 ();
 sg13g2_decap_8 FILLER_27_278 ();
 sg13g2_decap_8 FILLER_27_289 ();
 sg13g2_decap_4 FILLER_27_296 ();
 sg13g2_fill_2 FILLER_27_326 ();
 sg13g2_fill_1 FILLER_27_328 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_fill_1 FILLER_28_112 ();
 sg13g2_decap_4 FILLER_28_131 ();
 sg13g2_fill_1 FILLER_28_139 ();
 sg13g2_fill_1 FILLER_28_155 ();
 sg13g2_fill_2 FILLER_28_176 ();
 sg13g2_fill_1 FILLER_28_178 ();
 sg13g2_decap_4 FILLER_28_185 ();
 sg13g2_decap_4 FILLER_28_208 ();
 sg13g2_fill_1 FILLER_28_212 ();
 sg13g2_fill_2 FILLER_28_223 ();
 sg13g2_fill_1 FILLER_28_225 ();
 sg13g2_decap_8 FILLER_28_236 ();
 sg13g2_decap_4 FILLER_28_243 ();
 sg13g2_decap_8 FILLER_28_264 ();
 sg13g2_fill_2 FILLER_28_271 ();
 sg13g2_fill_1 FILLER_28_273 ();
 sg13g2_fill_2 FILLER_28_300 ();
 sg13g2_fill_1 FILLER_28_309 ();
 sg13g2_fill_2 FILLER_28_314 ();
 sg13g2_decap_8 FILLER_28_325 ();
 sg13g2_decap_4 FILLER_28_332 ();
 sg13g2_fill_2 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_359 ();
 sg13g2_decap_8 FILLER_28_366 ();
 sg13g2_decap_8 FILLER_28_373 ();
 sg13g2_decap_8 FILLER_28_380 ();
 sg13g2_decap_8 FILLER_28_387 ();
 sg13g2_decap_8 FILLER_28_394 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_fill_2 FILLER_29_105 ();
 sg13g2_fill_1 FILLER_29_107 ();
 sg13g2_fill_2 FILLER_29_130 ();
 sg13g2_fill_2 FILLER_29_148 ();
 sg13g2_fill_1 FILLER_29_150 ();
 sg13g2_fill_2 FILLER_29_157 ();
 sg13g2_fill_1 FILLER_29_159 ();
 sg13g2_fill_2 FILLER_29_178 ();
 sg13g2_fill_1 FILLER_29_180 ();
 sg13g2_fill_1 FILLER_29_206 ();
 sg13g2_decap_8 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_252 ();
 sg13g2_fill_2 FILLER_29_290 ();
 sg13g2_decap_4 FILLER_29_297 ();
 sg13g2_decap_4 FILLER_29_334 ();
 sg13g2_fill_2 FILLER_29_338 ();
 sg13g2_decap_8 FILLER_29_344 ();
 sg13g2_decap_8 FILLER_29_351 ();
 sg13g2_decap_8 FILLER_29_358 ();
 sg13g2_decap_8 FILLER_29_365 ();
 sg13g2_decap_8 FILLER_29_372 ();
 sg13g2_decap_8 FILLER_29_379 ();
 sg13g2_decap_8 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_4 FILLER_30_112 ();
 sg13g2_fill_2 FILLER_30_121 ();
 sg13g2_decap_8 FILLER_30_132 ();
 sg13g2_decap_8 FILLER_30_139 ();
 sg13g2_fill_2 FILLER_30_146 ();
 sg13g2_fill_1 FILLER_30_148 ();
 sg13g2_decap_4 FILLER_30_168 ();
 sg13g2_fill_2 FILLER_30_172 ();
 sg13g2_decap_8 FILLER_30_183 ();
 sg13g2_fill_2 FILLER_30_190 ();
 sg13g2_fill_1 FILLER_30_192 ();
 sg13g2_decap_8 FILLER_30_206 ();
 sg13g2_fill_2 FILLER_30_213 ();
 sg13g2_fill_1 FILLER_30_215 ();
 sg13g2_decap_8 FILLER_30_220 ();
 sg13g2_decap_8 FILLER_30_227 ();
 sg13g2_fill_2 FILLER_30_263 ();
 sg13g2_fill_1 FILLER_30_265 ();
 sg13g2_fill_1 FILLER_30_274 ();
 sg13g2_fill_2 FILLER_30_288 ();
 sg13g2_fill_2 FILLER_30_295 ();
 sg13g2_decap_8 FILLER_30_358 ();
 sg13g2_decap_8 FILLER_30_365 ();
 sg13g2_decap_8 FILLER_30_372 ();
 sg13g2_decap_8 FILLER_30_379 ();
 sg13g2_decap_8 FILLER_30_386 ();
 sg13g2_decap_8 FILLER_30_393 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_151 ();
 sg13g2_decap_8 FILLER_31_158 ();
 sg13g2_decap_8 FILLER_31_165 ();
 sg13g2_decap_8 FILLER_31_176 ();
 sg13g2_decap_8 FILLER_31_183 ();
 sg13g2_fill_2 FILLER_31_190 ();
 sg13g2_decap_4 FILLER_31_205 ();
 sg13g2_decap_8 FILLER_31_235 ();
 sg13g2_fill_2 FILLER_31_242 ();
 sg13g2_decap_4 FILLER_31_253 ();
 sg13g2_fill_2 FILLER_31_257 ();
 sg13g2_fill_2 FILLER_31_263 ();
 sg13g2_fill_1 FILLER_31_270 ();
 sg13g2_fill_2 FILLER_31_323 ();
 sg13g2_fill_1 FILLER_31_344 ();
 sg13g2_decap_8 FILLER_31_367 ();
 sg13g2_decap_8 FILLER_31_374 ();
 sg13g2_decap_8 FILLER_31_381 ();
 sg13g2_decap_8 FILLER_31_388 ();
 sg13g2_decap_8 FILLER_31_395 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_fill_2 FILLER_32_234 ();
 sg13g2_fill_1 FILLER_32_236 ();
 sg13g2_fill_1 FILLER_32_296 ();
 sg13g2_decap_8 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_decap_8 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_4 FILLER_33_189 ();
 sg13g2_fill_1 FILLER_33_219 ();
 sg13g2_decap_4 FILLER_33_261 ();
 sg13g2_fill_2 FILLER_33_265 ();
 sg13g2_fill_1 FILLER_33_293 ();
 sg13g2_decap_8 FILLER_33_374 ();
 sg13g2_decap_8 FILLER_33_381 ();
 sg13g2_decap_8 FILLER_33_388 ();
 sg13g2_decap_8 FILLER_33_395 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_fill_2 FILLER_34_182 ();
 sg13g2_fill_1 FILLER_34_215 ();
 sg13g2_decap_4 FILLER_34_250 ();
 sg13g2_fill_1 FILLER_34_254 ();
 sg13g2_fill_2 FILLER_34_260 ();
 sg13g2_fill_2 FILLER_34_266 ();
 sg13g2_fill_1 FILLER_34_268 ();
 sg13g2_fill_1 FILLER_34_272 ();
 sg13g2_decap_8 FILLER_34_378 ();
 sg13g2_decap_8 FILLER_34_385 ();
 sg13g2_decap_8 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_4 FILLER_35_189 ();
 sg13g2_fill_2 FILLER_35_193 ();
 sg13g2_fill_2 FILLER_35_199 ();
 sg13g2_fill_1 FILLER_35_201 ();
 sg13g2_fill_2 FILLER_35_215 ();
 sg13g2_fill_1 FILLER_35_230 ();
 sg13g2_fill_1 FILLER_35_245 ();
 sg13g2_fill_1 FILLER_35_313 ();
 sg13g2_fill_1 FILLER_35_341 ();
 sg13g2_decap_8 FILLER_35_368 ();
 sg13g2_decap_8 FILLER_35_375 ();
 sg13g2_decap_8 FILLER_35_382 ();
 sg13g2_decap_8 FILLER_35_389 ();
 sg13g2_decap_8 FILLER_35_396 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_4 FILLER_36_189 ();
 sg13g2_fill_2 FILLER_36_193 ();
 sg13g2_fill_2 FILLER_36_226 ();
 sg13g2_fill_2 FILLER_36_245 ();
 sg13g2_fill_2 FILLER_36_260 ();
 sg13g2_fill_1 FILLER_36_262 ();
 sg13g2_decap_4 FILLER_36_271 ();
 sg13g2_fill_1 FILLER_36_275 ();
 sg13g2_decap_4 FILLER_36_355 ();
 sg13g2_decap_8 FILLER_36_363 ();
 sg13g2_decap_8 FILLER_36_370 ();
 sg13g2_decap_8 FILLER_36_377 ();
 sg13g2_decap_8 FILLER_36_384 ();
 sg13g2_decap_8 FILLER_36_391 ();
 sg13g2_decap_8 FILLER_36_398 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_fill_2 FILLER_37_203 ();
 sg13g2_fill_1 FILLER_37_205 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_4 FILLER_37_217 ();
 sg13g2_fill_1 FILLER_37_239 ();
 sg13g2_decap_8 FILLER_37_271 ();
 sg13g2_decap_4 FILLER_37_278 ();
 sg13g2_decap_8 FILLER_37_326 ();
 sg13g2_fill_2 FILLER_37_333 ();
 sg13g2_fill_2 FILLER_37_347 ();
 sg13g2_fill_2 FILLER_37_353 ();
 sg13g2_decap_8 FILLER_37_359 ();
 sg13g2_decap_8 FILLER_37_366 ();
 sg13g2_fill_1 FILLER_37_373 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_123 ();
 sg13g2_fill_1 FILLER_38_127 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_8 FILLER_38_164 ();
 sg13g2_decap_8 FILLER_38_171 ();
 sg13g2_decap_8 FILLER_38_178 ();
 sg13g2_decap_8 FILLER_38_185 ();
 sg13g2_decap_8 FILLER_38_192 ();
 sg13g2_decap_8 FILLER_38_199 ();
 sg13g2_decap_8 FILLER_38_206 ();
 sg13g2_decap_8 FILLER_38_213 ();
 sg13g2_decap_8 FILLER_38_304 ();
 sg13g2_fill_1 FILLER_38_315 ();
 sg13g2_decap_8 FILLER_38_319 ();
 sg13g2_decap_4 FILLER_38_326 ();
 sg13g2_fill_1 FILLER_38_330 ();
 sg13g2_decap_8 FILLER_38_335 ();
 sg13g2_decap_8 FILLER_38_342 ();
 sg13g2_decap_8 FILLER_38_349 ();
 sg13g2_decap_8 FILLER_38_356 ();
 sg13g2_fill_2 FILLER_38_363 ();
 sg13g2_fill_1 FILLER_38_365 ();
 sg13g2_decap_4 FILLER_38_370 ();
 sg13g2_fill_2 FILLER_38_374 ();
 sg13g2_decap_8 FILLER_38_380 ();
 sg13g2_decap_8 FILLER_38_387 ();
 sg13g2_decap_8 FILLER_38_394 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net59;
 assign uio_oe[1] = net60;
 assign uio_oe[2] = net61;
 assign uio_oe[3] = net62;
 assign uio_oe[4] = net63;
 assign uio_oe[5] = net64;
 assign uio_oe[6] = net65;
 assign uio_oe[7] = net66;
 assign uio_out[2] = net2;
 assign uio_out[3] = net3;
 assign uio_out[4] = net4;
 assign uio_out[5] = net5;
 assign uio_out[6] = net6;
endmodule

module tt_um_rejunity_ay8913 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net41;
 wire net33;
 wire net25;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire active;
 wire \amplitude_A[0] ;
 wire \amplitude_A[1] ;
 wire \amplitude_A[2] ;
 wire \amplitude_A[3] ;
 wire \amplitude_B[0] ;
 wire \amplitude_B[1] ;
 wire \amplitude_B[2] ;
 wire \amplitude_B[3] ;
 wire \amplitude_C[0] ;
 wire \amplitude_C[1] ;
 wire \amplitude_C[2] ;
 wire \amplitude_C[3] ;
 wire \attenuation_A.out[0] ;
 wire \attenuation_A.out[1] ;
 wire \attenuation_A.out[2] ;
 wire \attenuation_A.out[3] ;
 wire \attenuation_A.out[4] ;
 wire \attenuation_A.out[5] ;
 wire \attenuation_A.out[6] ;
 wire \attenuation_A.out[7] ;
 wire \attenuation_B.out[0] ;
 wire \attenuation_B.out[1] ;
 wire \attenuation_B.out[2] ;
 wire \attenuation_B.out[3] ;
 wire \attenuation_B.out[4] ;
 wire \attenuation_B.out[5] ;
 wire \attenuation_B.out[6] ;
 wire \attenuation_B.out[7] ;
 wire \attenuation_C.out[0] ;
 wire \attenuation_C.out[1] ;
 wire \attenuation_C.out[2] ;
 wire \attenuation_C.out[3] ;
 wire \attenuation_C.out[4] ;
 wire \attenuation_C.out[5] ;
 wire \attenuation_C.out[6] ;
 wire \attenuation_C.out[7] ;
 wire \clk_counter[0] ;
 wire \clk_counter[1] ;
 wire \clk_counter[2] ;
 wire \clk_counter[3] ;
 wire \clk_counter[4] ;
 wire \clk_counter[5] ;
 wire \clk_counter[6] ;
 wire envelope_A;
 wire envelope_B;
 wire envelope_C;
 wire envelope_alternate;
 wire envelope_attack;
 wire envelope_continue;
 wire \envelope_generator.envelope_counter[0] ;
 wire \envelope_generator.envelope_counter[1] ;
 wire \envelope_generator.envelope_counter[2] ;
 wire \envelope_generator.envelope_counter[3] ;
 wire \envelope_generator.hold ;
 wire \envelope_generator.invert_output ;
 wire \envelope_generator.period[0] ;
 wire \envelope_generator.period[10] ;
 wire \envelope_generator.period[11] ;
 wire \envelope_generator.period[12] ;
 wire \envelope_generator.period[13] ;
 wire \envelope_generator.period[14] ;
 wire \envelope_generator.period[15] ;
 wire \envelope_generator.period[1] ;
 wire \envelope_generator.period[2] ;
 wire \envelope_generator.period[3] ;
 wire \envelope_generator.period[4] ;
 wire \envelope_generator.period[5] ;
 wire \envelope_generator.period[6] ;
 wire \envelope_generator.period[7] ;
 wire \envelope_generator.period[8] ;
 wire \envelope_generator.period[9] ;
 wire \envelope_generator.signal_edge.previous_signal_state_0 ;
 wire \envelope_generator.signal_edge.signal ;
 wire \envelope_generator.stop ;
 wire \envelope_generator.tone.counter[0] ;
 wire \envelope_generator.tone.counter[10] ;
 wire \envelope_generator.tone.counter[11] ;
 wire \envelope_generator.tone.counter[12] ;
 wire \envelope_generator.tone.counter[13] ;
 wire \envelope_generator.tone.counter[14] ;
 wire \envelope_generator.tone.counter[15] ;
 wire \envelope_generator.tone.counter[1] ;
 wire \envelope_generator.tone.counter[2] ;
 wire \envelope_generator.tone.counter[3] ;
 wire \envelope_generator.tone.counter[4] ;
 wire \envelope_generator.tone.counter[5] ;
 wire \envelope_generator.tone.counter[6] ;
 wire \envelope_generator.tone.counter[7] ;
 wire \envelope_generator.tone.counter[8] ;
 wire \envelope_generator.tone.counter[9] ;
 wire \latched_register[0] ;
 wire \latched_register[1] ;
 wire \latched_register[2] ;
 wire \latched_register[3] ;
 wire noise_disable_A;
 wire noise_disable_B;
 wire noise_disable_C;
 wire \noise_generator.lfsr[0] ;
 wire \noise_generator.lfsr[10] ;
 wire \noise_generator.lfsr[11] ;
 wire \noise_generator.lfsr[12] ;
 wire \noise_generator.lfsr[13] ;
 wire \noise_generator.lfsr[14] ;
 wire \noise_generator.lfsr[15] ;
 wire \noise_generator.lfsr[16] ;
 wire \noise_generator.lfsr[1] ;
 wire \noise_generator.lfsr[2] ;
 wire \noise_generator.lfsr[3] ;
 wire \noise_generator.lfsr[4] ;
 wire \noise_generator.lfsr[5] ;
 wire \noise_generator.lfsr[6] ;
 wire \noise_generator.lfsr[7] ;
 wire \noise_generator.lfsr[8] ;
 wire \noise_generator.lfsr[9] ;
 wire \noise_generator.period[0] ;
 wire \noise_generator.period[1] ;
 wire \noise_generator.period[2] ;
 wire \noise_generator.period[3] ;
 wire \noise_generator.period[4] ;
 wire \noise_generator.signal_edge.previous_signal_state_0 ;
 wire \noise_generator.signal_edge.signal ;
 wire \noise_generator.tone.counter[0] ;
 wire \noise_generator.tone.counter[1] ;
 wire \noise_generator.tone.counter[2] ;
 wire \noise_generator.tone.counter[3] ;
 wire \noise_generator.tone.counter[4] ;
 wire \pwm_A.accumulator[0] ;
 wire \pwm_A.accumulator[1] ;
 wire \pwm_A.accumulator[2] ;
 wire \pwm_A.accumulator[3] ;
 wire \pwm_A.accumulator[4] ;
 wire \pwm_A.accumulator[5] ;
 wire \pwm_A.accumulator[6] ;
 wire \pwm_A.accumulator[7] ;
 wire \pwm_A.accumulator[8] ;
 wire \pwm_B.accumulator[0] ;
 wire \pwm_B.accumulator[1] ;
 wire \pwm_B.accumulator[2] ;
 wire \pwm_B.accumulator[3] ;
 wire \pwm_B.accumulator[4] ;
 wire \pwm_B.accumulator[5] ;
 wire \pwm_B.accumulator[6] ;
 wire \pwm_B.accumulator[7] ;
 wire \pwm_B.accumulator[8] ;
 wire \pwm_C.accumulator[0] ;
 wire \pwm_C.accumulator[1] ;
 wire \pwm_C.accumulator[2] ;
 wire \pwm_C.accumulator[3] ;
 wire \pwm_C.accumulator[4] ;
 wire \pwm_C.accumulator[5] ;
 wire \pwm_C.accumulator[6] ;
 wire \pwm_C.accumulator[7] ;
 wire \pwm_C.accumulator[8] ;
 wire \pwm_master.accumulator[0] ;
 wire \pwm_master.accumulator[1] ;
 wire \pwm_master.accumulator[2] ;
 wire \pwm_master.accumulator[3] ;
 wire \pwm_master.accumulator[4] ;
 wire \pwm_master.accumulator[5] ;
 wire \pwm_master.accumulator[6] ;
 wire \pwm_master.accumulator[7] ;
 wire \pwm_master.accumulator[8] ;
 wire \pwm_master.accumulator[9] ;
 wire \register[0][0] ;
 wire \register[0][1] ;
 wire \register[0][2] ;
 wire \register[0][3] ;
 wire \register[0][4] ;
 wire \register[0][5] ;
 wire \register[0][6] ;
 wire \register[0][7] ;
 wire \register[1][0] ;
 wire \register[1][1] ;
 wire \register[1][2] ;
 wire \register[1][3] ;
 wire \register[2][0] ;
 wire \register[2][1] ;
 wire \register[2][2] ;
 wire \register[2][3] ;
 wire \register[2][4] ;
 wire \register[2][5] ;
 wire \register[2][6] ;
 wire \register[2][7] ;
 wire \register[3][0] ;
 wire \register[3][1] ;
 wire \register[3][2] ;
 wire \register[3][3] ;
 wire \register[4][0] ;
 wire \register[4][1] ;
 wire \register[4][2] ;
 wire \register[4][3] ;
 wire \register[4][4] ;
 wire \register[4][5] ;
 wire \register[4][6] ;
 wire \register[4][7] ;
 wire \register[5][0] ;
 wire \register[5][1] ;
 wire \register[5][2] ;
 wire \register[5][3] ;
 wire restart_envelope;
 wire tone_A;
 wire \tone_A_generator.counter[0] ;
 wire \tone_A_generator.counter[10] ;
 wire \tone_A_generator.counter[11] ;
 wire \tone_A_generator.counter[1] ;
 wire \tone_A_generator.counter[2] ;
 wire \tone_A_generator.counter[3] ;
 wire \tone_A_generator.counter[4] ;
 wire \tone_A_generator.counter[5] ;
 wire \tone_A_generator.counter[6] ;
 wire \tone_A_generator.counter[7] ;
 wire \tone_A_generator.counter[8] ;
 wire \tone_A_generator.counter[9] ;
 wire tone_B;
 wire \tone_B_generator.counter[0] ;
 wire \tone_B_generator.counter[10] ;
 wire \tone_B_generator.counter[11] ;
 wire \tone_B_generator.counter[1] ;
 wire \tone_B_generator.counter[2] ;
 wire \tone_B_generator.counter[3] ;
 wire \tone_B_generator.counter[4] ;
 wire \tone_B_generator.counter[5] ;
 wire \tone_B_generator.counter[6] ;
 wire \tone_B_generator.counter[7] ;
 wire \tone_B_generator.counter[8] ;
 wire \tone_B_generator.counter[9] ;
 wire tone_C;
 wire \tone_C_generator.counter[0] ;
 wire \tone_C_generator.counter[10] ;
 wire \tone_C_generator.counter[11] ;
 wire \tone_C_generator.counter[1] ;
 wire \tone_C_generator.counter[2] ;
 wire \tone_C_generator.counter[3] ;
 wire \tone_C_generator.counter[4] ;
 wire \tone_C_generator.counter[5] ;
 wire \tone_C_generator.counter[6] ;
 wire \tone_C_generator.counter[7] ;
 wire \tone_C_generator.counter[8] ;
 wire \tone_C_generator.counter[9] ;
 wire tone_disable_A;
 wire tone_disable_B;
 wire tone_disable_C;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net330;
 wire net331;
 wire net332;
 wire clknet_leaf_0_clk;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;

 sg13g2_inv_1 _1545_ (.Y(_0723_),
    .A(net334));
 sg13g2_inv_1 _1546_ (.Y(_0724_),
    .A(net387));
 sg13g2_inv_1 _1547_ (.Y(_0725_),
    .A(\envelope_generator.tone.counter[15] ));
 sg13g2_inv_1 _1548_ (.Y(_0726_),
    .A(\envelope_generator.tone.counter[13] ));
 sg13g2_inv_1 _1549_ (.Y(_0727_),
    .A(\envelope_generator.tone.counter[10] ));
 sg13g2_inv_1 _1550_ (.Y(_0728_),
    .A(\envelope_generator.tone.counter[8] ));
 sg13g2_inv_1 _1551_ (.Y(_0729_),
    .A(\envelope_generator.tone.counter[7] ));
 sg13g2_inv_1 _1552_ (.Y(_0730_),
    .A(net544));
 sg13g2_inv_1 _1553_ (.Y(_0731_),
    .A(net619));
 sg13g2_inv_1 _1554_ (.Y(_0732_),
    .A(\envelope_generator.tone.counter[2] ));
 sg13g2_inv_1 _1555_ (.Y(_0733_),
    .A(net429));
 sg13g2_inv_1 _1556_ (.Y(_0734_),
    .A(\envelope_generator.tone.counter[0] ));
 sg13g2_inv_1 _1557_ (.Y(_0735_),
    .A(net469));
 sg13g2_inv_1 _1558_ (.Y(_0736_),
    .A(net432));
 sg13g2_inv_1 _1559_ (.Y(_0737_),
    .A(net495));
 sg13g2_inv_1 _1560_ (.Y(_0738_),
    .A(net453));
 sg13g2_inv_1 _1561_ (.Y(_0739_),
    .A(net465));
 sg13g2_inv_1 _1562_ (.Y(_0740_),
    .A(net449));
 sg13g2_inv_1 _1563_ (.Y(_0741_),
    .A(net480));
 sg13g2_inv_1 _1564_ (.Y(_0742_),
    .A(net416));
 sg13g2_inv_1 _1565_ (.Y(_0743_),
    .A(net456));
 sg13g2_inv_1 _1566_ (.Y(_0744_),
    .A(net459));
 sg13g2_inv_1 _1567_ (.Y(_0745_),
    .A(net473));
 sg13g2_inv_1 _1568_ (.Y(_0746_),
    .A(net503));
 sg13g2_inv_1 _1569_ (.Y(_0747_),
    .A(net462));
 sg13g2_inv_1 _1570_ (.Y(_0748_),
    .A(net471));
 sg13g2_inv_1 _1571_ (.Y(_0749_),
    .A(net434));
 sg13g2_inv_1 _1572_ (.Y(_0750_),
    .A(net472));
 sg13g2_inv_1 _1573_ (.Y(_0751_),
    .A(\noise_generator.tone.counter[4] ));
 sg13g2_inv_1 _1574_ (.Y(_0752_),
    .A(\noise_generator.tone.counter[3] ));
 sg13g2_inv_1 _1575_ (.Y(_0753_),
    .A(net375));
 sg13g2_inv_1 _1576_ (.Y(_0754_),
    .A(\noise_generator.tone.counter[0] ));
 sg13g2_inv_1 _1577_ (.Y(_0755_),
    .A(\tone_C_generator.counter[11] ));
 sg13g2_inv_1 _1578_ (.Y(_0756_),
    .A(\tone_C_generator.counter[10] ));
 sg13g2_inv_1 _1579_ (.Y(_0757_),
    .A(\tone_C_generator.counter[9] ));
 sg13g2_inv_1 _1580_ (.Y(_0758_),
    .A(net610));
 sg13g2_inv_1 _1581_ (.Y(_0759_),
    .A(\tone_C_generator.counter[6] ));
 sg13g2_inv_1 _1582_ (.Y(_0760_),
    .A(\tone_C_generator.counter[5] ));
 sg13g2_inv_1 _1583_ (.Y(_0761_),
    .A(\tone_C_generator.counter[4] ));
 sg13g2_inv_1 _1584_ (.Y(_0762_),
    .A(\tone_B_generator.counter[11] ));
 sg13g2_inv_1 _1585_ (.Y(_0763_),
    .A(\tone_B_generator.counter[10] ));
 sg13g2_inv_1 _1586_ (.Y(_0764_),
    .A(\tone_B_generator.counter[8] ));
 sg13g2_inv_1 _1587_ (.Y(_0765_),
    .A(\tone_B_generator.counter[3] ));
 sg13g2_inv_1 _1588_ (.Y(_0766_),
    .A(\tone_B_generator.counter[2] ));
 sg13g2_inv_1 _1589_ (.Y(_0767_),
    .A(\tone_B_generator.counter[1] ));
 sg13g2_inv_1 _1590_ (.Y(_0768_),
    .A(tone_B));
 sg13g2_inv_1 _1591_ (.Y(_0769_),
    .A(\tone_A_generator.counter[11] ));
 sg13g2_inv_1 _1592_ (.Y(_0770_),
    .A(\tone_A_generator.counter[10] ));
 sg13g2_inv_1 _1593_ (.Y(_0771_),
    .A(\tone_A_generator.counter[8] ));
 sg13g2_inv_1 _1594_ (.Y(_0772_),
    .A(net611));
 sg13g2_inv_1 _1595_ (.Y(_0773_),
    .A(\tone_A_generator.counter[5] ));
 sg13g2_inv_1 _1596_ (.Y(_0774_),
    .A(\tone_A_generator.counter[4] ));
 sg13g2_inv_1 _1597_ (.Y(_0775_),
    .A(\tone_A_generator.counter[2] ));
 sg13g2_inv_1 _1598_ (.Y(_0776_),
    .A(net384));
 sg13g2_inv_1 _1599_ (.Y(_0777_),
    .A(\tone_A_generator.counter[0] ));
 sg13g2_inv_1 _1600_ (.Y(_0778_),
    .A(net598));
 sg13g2_inv_1 _1601_ (.Y(_0779_),
    .A(net595));
 sg13g2_inv_1 _1602_ (.Y(_0780_),
    .A(net599));
 sg13g2_inv_1 _1603_ (.Y(_0781_),
    .A(net596));
 sg13g2_inv_1 _1604_ (.Y(_0782_),
    .A(net593));
 sg13g2_inv_1 _1605_ (.Y(_0783_),
    .A(net451));
 sg13g2_inv_1 _1606_ (.Y(_0784_),
    .A(\noise_generator.period[4] ));
 sg13g2_inv_1 _1607_ (.Y(_0785_),
    .A(\envelope_generator.period[11] ));
 sg13g2_inv_1 _1608_ (.Y(_0786_),
    .A(\envelope_generator.period[10] ));
 sg13g2_inv_1 _1609_ (.Y(_0787_),
    .A(\envelope_generator.period[9] ));
 sg13g2_inv_1 _1610_ (.Y(_0788_),
    .A(\envelope_generator.period[7] ));
 sg13g2_inv_1 _1611_ (.Y(_0789_),
    .A(\envelope_generator.period[6] ));
 sg13g2_inv_1 _1612_ (.Y(_0790_),
    .A(\envelope_generator.period[5] ));
 sg13g2_inv_1 _1613_ (.Y(_0791_),
    .A(\envelope_generator.period[4] ));
 sg13g2_inv_1 _1614_ (.Y(_0792_),
    .A(\envelope_generator.period[3] ));
 sg13g2_inv_1 _1615_ (.Y(_0793_),
    .A(\register[4][0] ));
 sg13g2_inv_1 _1616_ (.Y(_0794_),
    .A(\register[4][1] ));
 sg13g2_inv_1 _1617_ (.Y(_0795_),
    .A(\register[4][4] ));
 sg13g2_inv_1 _1618_ (.Y(_0796_),
    .A(\register[5][2] ));
 sg13g2_inv_1 _1619_ (.Y(_0797_),
    .A(\register[5][1] ));
 sg13g2_inv_1 _1620_ (.Y(_0798_),
    .A(\register[3][2] ));
 sg13g2_inv_1 _1621_ (.Y(_0799_),
    .A(\register[3][1] ));
 sg13g2_inv_1 _1622_ (.Y(_0800_),
    .A(\register[3][0] ));
 sg13g2_inv_1 _1623_ (.Y(_0801_),
    .A(\register[2][7] ));
 sg13g2_inv_1 _1624_ (.Y(_0802_),
    .A(\register[2][6] ));
 sg13g2_inv_1 _1625_ (.Y(_0803_),
    .A(\register[2][5] ));
 sg13g2_inv_1 _1626_ (.Y(_0804_),
    .A(\register[2][4] ));
 sg13g2_inv_1 _1627_ (.Y(_0805_),
    .A(\register[2][3] ));
 sg13g2_inv_1 _1628_ (.Y(_0806_),
    .A(\register[1][3] ));
 sg13g2_inv_1 _1629_ (.Y(_0807_),
    .A(\register[1][2] ));
 sg13g2_inv_1 _1630_ (.Y(_0808_),
    .A(\register[1][1] ));
 sg13g2_inv_1 _1631_ (.Y(_0809_),
    .A(\register[1][0] ));
 sg13g2_inv_1 _1632_ (.Y(_0810_),
    .A(\register[0][6] ));
 sg13g2_inv_1 _1633_ (.Y(_0811_),
    .A(\register[0][4] ));
 sg13g2_inv_1 _1634_ (.Y(_0812_),
    .A(\register[0][3] ));
 sg13g2_inv_1 _1635_ (.Y(_0813_),
    .A(\register[0][2] ));
 sg13g2_inv_2 _1636_ (.Y(_0814_),
    .A(net186));
 sg13g2_inv_1 _1637_ (.Y(_0815_),
    .A(net5));
 sg13g2_inv_1 _1638_ (.Y(_0816_),
    .A(net6));
 sg13g2_inv_1 _1639_ (.Y(_0817_),
    .A(net336));
 sg13g2_inv_1 _1640_ (.Y(_0818_),
    .A(noise_disable_A));
 sg13g2_inv_1 _1641_ (.Y(_0819_),
    .A(_0018_));
 sg13g2_inv_1 _1642_ (.Y(_0820_),
    .A(_0021_));
 sg13g2_inv_1 _1643_ (.Y(_0821_),
    .A(\pwm_master.accumulator[1] ));
 sg13g2_inv_1 _1644_ (.Y(_0822_),
    .A(net620));
 sg13g2_inv_1 _1645_ (.Y(_0823_),
    .A(net634));
 sg13g2_inv_1 _1646_ (.Y(_0824_),
    .A(net622));
 sg13g2_and2_1 _1647_ (.A(\attenuation_B.out[7] ),
    .B(\attenuation_A.out[7] ),
    .X(_0825_));
 sg13g2_xor2_1 _1648_ (.B(\attenuation_A.out[7] ),
    .A(\attenuation_B.out[7] ),
    .X(_0826_));
 sg13g2_a21oi_1 _1649_ (.A1(\attenuation_C.out[7] ),
    .A2(_0826_),
    .Y(_0827_),
    .B1(_0825_));
 sg13g2_and2_1 _1650_ (.A(\attenuation_B.out[6] ),
    .B(\attenuation_A.out[6] ),
    .X(_0828_));
 sg13g2_xor2_1 _1651_ (.B(\attenuation_A.out[6] ),
    .A(\attenuation_B.out[6] ),
    .X(_0829_));
 sg13g2_a21oi_1 _1652_ (.A1(\attenuation_C.out[6] ),
    .A2(_0829_),
    .Y(_0830_),
    .B1(_0828_));
 sg13g2_xnor2_1 _1653_ (.Y(_0831_),
    .A(\attenuation_C.out[7] ),
    .B(_0826_));
 sg13g2_or2_1 _1654_ (.X(_0832_),
    .B(_0831_),
    .A(_0830_));
 sg13g2_and2_1 _1655_ (.A(\attenuation_B.out[5] ),
    .B(\attenuation_A.out[5] ),
    .X(_0833_));
 sg13g2_xor2_1 _1656_ (.B(\attenuation_A.out[5] ),
    .A(\attenuation_B.out[5] ),
    .X(_0834_));
 sg13g2_a21oi_2 _1657_ (.B1(_0833_),
    .Y(_0835_),
    .A2(_0834_),
    .A1(\attenuation_C.out[5] ));
 sg13g2_xnor2_1 _1658_ (.Y(_0836_),
    .A(\attenuation_C.out[6] ),
    .B(_0829_));
 sg13g2_nor2_1 _1659_ (.A(_0835_),
    .B(_0836_),
    .Y(_0837_));
 sg13g2_xor2_1 _1660_ (.B(_0836_),
    .A(_0835_),
    .X(_0838_));
 sg13g2_inv_1 _1661_ (.Y(_0839_),
    .A(_0838_));
 sg13g2_and2_1 _1662_ (.A(\attenuation_B.out[4] ),
    .B(\attenuation_A.out[4] ),
    .X(_0840_));
 sg13g2_xor2_1 _1663_ (.B(\attenuation_A.out[4] ),
    .A(\attenuation_B.out[4] ),
    .X(_0841_));
 sg13g2_a21oi_2 _1664_ (.B1(_0840_),
    .Y(_0842_),
    .A2(_0841_),
    .A1(\attenuation_C.out[4] ));
 sg13g2_xnor2_1 _1665_ (.Y(_0843_),
    .A(\attenuation_C.out[5] ),
    .B(_0834_));
 sg13g2_nor2_1 _1666_ (.A(_0842_),
    .B(_0843_),
    .Y(_0844_));
 sg13g2_nand2_1 _1667_ (.Y(_0845_),
    .A(_0842_),
    .B(_0843_));
 sg13g2_xnor2_1 _1668_ (.Y(_0846_),
    .A(\attenuation_C.out[4] ),
    .B(_0841_));
 sg13g2_and2_1 _1669_ (.A(\attenuation_B.out[3] ),
    .B(\attenuation_A.out[3] ),
    .X(_0847_));
 sg13g2_xor2_1 _1670_ (.B(\attenuation_A.out[3] ),
    .A(\attenuation_B.out[3] ),
    .X(_0848_));
 sg13g2_a21oi_2 _1671_ (.B1(_0847_),
    .Y(_0849_),
    .A2(_0848_),
    .A1(\attenuation_C.out[3] ));
 sg13g2_nor2_1 _1672_ (.A(_0846_),
    .B(_0849_),
    .Y(_0850_));
 sg13g2_and2_1 _1673_ (.A(\attenuation_B.out[2] ),
    .B(\attenuation_A.out[2] ),
    .X(_0851_));
 sg13g2_xor2_1 _1674_ (.B(\attenuation_A.out[2] ),
    .A(\attenuation_B.out[2] ),
    .X(_0852_));
 sg13g2_xnor2_1 _1675_ (.Y(_0853_),
    .A(\attenuation_C.out[2] ),
    .B(_0852_));
 sg13g2_and2_1 _1676_ (.A(\attenuation_B.out[1] ),
    .B(\attenuation_A.out[1] ),
    .X(_0854_));
 sg13g2_xor2_1 _1677_ (.B(\attenuation_A.out[1] ),
    .A(\attenuation_B.out[1] ),
    .X(_0855_));
 sg13g2_a21oi_2 _1678_ (.B1(_0854_),
    .Y(_0856_),
    .A2(_0855_),
    .A1(\attenuation_C.out[1] ));
 sg13g2_nor2_1 _1679_ (.A(_0853_),
    .B(_0856_),
    .Y(_0857_));
 sg13g2_nand2_1 _1680_ (.Y(_0858_),
    .A(_0853_),
    .B(_0856_));
 sg13g2_xnor2_1 _1681_ (.Y(_0859_),
    .A(_0853_),
    .B(_0856_));
 sg13g2_xnor2_1 _1682_ (.Y(_0860_),
    .A(\attenuation_C.out[1] ),
    .B(_0855_));
 sg13g2_and2_1 _1683_ (.A(\attenuation_B.out[0] ),
    .B(\attenuation_A.out[0] ),
    .X(_0861_));
 sg13g2_xor2_1 _1684_ (.B(\attenuation_A.out[0] ),
    .A(\attenuation_B.out[0] ),
    .X(_0862_));
 sg13g2_a21oi_2 _1685_ (.B1(_0861_),
    .Y(_0863_),
    .A2(_0862_),
    .A1(\attenuation_C.out[0] ));
 sg13g2_nor2_1 _1686_ (.A(_0860_),
    .B(_0863_),
    .Y(_0864_));
 sg13g2_a21oi_2 _1687_ (.B1(_0851_),
    .Y(_0865_),
    .A2(_0852_),
    .A1(\attenuation_C.out[2] ));
 sg13g2_xnor2_1 _1688_ (.Y(_0866_),
    .A(\attenuation_C.out[3] ),
    .B(_0848_));
 sg13g2_nand2_1 _1689_ (.Y(_0867_),
    .A(_0865_),
    .B(_0866_));
 sg13g2_nor2_1 _1690_ (.A(_0865_),
    .B(_0866_),
    .Y(_0868_));
 sg13g2_xor2_1 _1691_ (.B(_0866_),
    .A(_0865_),
    .X(_0869_));
 sg13g2_nand3b_1 _1692_ (.B(_0864_),
    .C(_0869_),
    .Y(_0870_),
    .A_N(_0859_));
 sg13g2_a21oi_1 _1693_ (.A1(_0857_),
    .A2(_0867_),
    .Y(_0871_),
    .B1(_0868_));
 sg13g2_nand2_1 _1694_ (.Y(_0872_),
    .A(_0870_),
    .B(_0871_));
 sg13g2_xnor2_1 _1695_ (.Y(_0873_),
    .A(_0846_),
    .B(_0849_));
 sg13g2_inv_1 _1696_ (.Y(_0874_),
    .A(_0873_));
 sg13g2_a21oi_1 _1697_ (.A1(_0872_),
    .A2(_0874_),
    .Y(_0875_),
    .B1(_0850_));
 sg13g2_a21oi_1 _1698_ (.A1(_0845_),
    .A2(_0850_),
    .Y(_0876_),
    .B1(_0844_));
 sg13g2_xor2_1 _1699_ (.B(_0843_),
    .A(_0842_),
    .X(_0877_));
 sg13g2_nand2b_1 _1700_ (.Y(_0878_),
    .B(_0877_),
    .A_N(_0873_));
 sg13g2_a21o_1 _1701_ (.A2(_0871_),
    .A1(_0870_),
    .B1(_0878_),
    .X(_0879_));
 sg13g2_a21oi_2 _1702_ (.B1(_0839_),
    .Y(_0880_),
    .A2(_0879_),
    .A1(_0876_));
 sg13g2_xor2_1 _1703_ (.B(_0831_),
    .A(_0830_),
    .X(_0881_));
 sg13g2_o21ai_1 _1704_ (.B1(_0881_),
    .Y(_0882_),
    .A1(_0837_),
    .A2(_0880_));
 sg13g2_a21o_2 _1705_ (.A2(_0882_),
    .A1(_0832_),
    .B1(_0827_),
    .X(_0883_));
 sg13g2_inv_1 _1706_ (.Y(_0884_),
    .A(_0883_));
 sg13g2_xnor2_1 _1707_ (.Y(_0885_),
    .A(_0860_),
    .B(_0863_));
 sg13g2_nand2_1 _1708_ (.Y(uo_out[0]),
    .A(_0883_),
    .B(_0885_));
 sg13g2_xnor2_1 _1709_ (.Y(_0886_),
    .A(_0859_),
    .B(_0864_));
 sg13g2_or2_1 _1710_ (.X(uo_out[1]),
    .B(_0886_),
    .A(_0884_));
 sg13g2_a21oi_1 _1711_ (.A1(_0858_),
    .A2(_0864_),
    .Y(_0887_),
    .B1(_0857_));
 sg13g2_xnor2_1 _1712_ (.Y(_0888_),
    .A(_0869_),
    .B(_0887_));
 sg13g2_or2_1 _1713_ (.X(uo_out[2]),
    .B(_0888_),
    .A(_0884_));
 sg13g2_xnor2_1 _1714_ (.Y(_0889_),
    .A(_0872_),
    .B(_0874_));
 sg13g2_nand2_1 _1715_ (.Y(uo_out[3]),
    .A(_0883_),
    .B(_0889_));
 sg13g2_xor2_1 _1716_ (.B(_0877_),
    .A(_0875_),
    .X(_0890_));
 sg13g2_nand2_1 _1717_ (.Y(uo_out[4]),
    .A(_0883_),
    .B(_0890_));
 sg13g2_nand3_1 _1718_ (.B(_0876_),
    .C(_0879_),
    .A(_0839_),
    .Y(_0891_));
 sg13g2_nor2b_2 _1719_ (.A(_0880_),
    .B_N(_0891_),
    .Y(_0892_));
 sg13g2_or2_1 _1720_ (.X(uo_out[5]),
    .B(_0892_),
    .A(_0884_));
 sg13g2_or3_1 _1721_ (.A(_0837_),
    .B(_0880_),
    .C(_0881_),
    .X(_0893_));
 sg13g2_nand2_1 _1722_ (.Y(_0894_),
    .A(_0882_),
    .B(_0893_));
 sg13g2_nand2_1 _1723_ (.Y(uo_out[6]),
    .A(_0883_),
    .B(_0894_));
 sg13g2_nand3_1 _1724_ (.B(_0832_),
    .C(_0882_),
    .A(_0827_),
    .Y(uo_out[7]));
 sg13g2_xnor2_1 _1725_ (.Y(_0895_),
    .A(\envelope_generator.envelope_counter[2] ),
    .B(\envelope_generator.invert_output ));
 sg13g2_nor2_1 _1726_ (.A(tone_A),
    .B(tone_disable_A),
    .Y(_0896_));
 sg13g2_a21oi_2 _1727_ (.B1(_0896_),
    .Y(_0897_),
    .A2(_0818_),
    .A1(\noise_generator.lfsr[0] ));
 sg13g2_nor2b_1 _1728_ (.A(net161),
    .B_N(_0010_),
    .Y(_0898_));
 sg13g2_a21oi_2 _1729_ (.B1(_0898_),
    .Y(_0899_),
    .A2(_0895_),
    .A1(envelope_A));
 sg13g2_nand2_2 _1730_ (.Y(_0900_),
    .A(_0897_),
    .B(_0899_));
 sg13g2_xnor2_1 _1731_ (.Y(_0901_),
    .A(\envelope_generator.envelope_counter[0] ),
    .B(\envelope_generator.invert_output ));
 sg13g2_nand2_1 _1732_ (.Y(_0902_),
    .A(net161),
    .B(_0901_));
 sg13g2_nand2b_1 _1733_ (.Y(_0903_),
    .B(_0012_),
    .A_N(net161));
 sg13g2_and3_1 _1734_ (.X(_0904_),
    .A(_0897_),
    .B(_0902_),
    .C(_0903_));
 sg13g2_nand3_1 _1735_ (.B(_0902_),
    .C(_0903_),
    .A(_0897_),
    .Y(_0905_));
 sg13g2_xnor2_1 _1736_ (.Y(_0906_),
    .A(\envelope_generator.envelope_counter[1] ),
    .B(\envelope_generator.invert_output ));
 sg13g2_nor2b_1 _1737_ (.A(net161),
    .B_N(_0013_),
    .Y(_0907_));
 sg13g2_a21oi_2 _1738_ (.B1(_0907_),
    .Y(_0908_),
    .A2(_0906_),
    .A1(net161));
 sg13g2_nand2_1 _1739_ (.Y(_0909_),
    .A(_0897_),
    .B(_0908_));
 sg13g2_nand4_1 _1740_ (.B(_0900_),
    .C(_0905_),
    .A(_0897_),
    .Y(_0910_),
    .D(_0908_));
 sg13g2_xnor2_1 _1741_ (.Y(_0911_),
    .A(\envelope_generator.envelope_counter[3] ),
    .B(\envelope_generator.invert_output ));
 sg13g2_nand2_1 _1742_ (.Y(_0912_),
    .A(net161),
    .B(_0911_));
 sg13g2_nand2b_1 _1743_ (.Y(_0913_),
    .B(_0011_),
    .A_N(net161));
 sg13g2_and3_2 _1744_ (.X(_0914_),
    .A(_0897_),
    .B(_0912_),
    .C(_0913_));
 sg13g2_nand3_1 _1745_ (.B(_0912_),
    .C(_0913_),
    .A(_0897_),
    .Y(_0915_));
 sg13g2_nor2_1 _1746_ (.A(_0904_),
    .B(_0914_),
    .Y(_0916_));
 sg13g2_nor3_1 _1747_ (.A(_0900_),
    .B(_0904_),
    .C(_0914_),
    .Y(_0917_));
 sg13g2_o21ai_1 _1748_ (.B1(_0910_),
    .Y(_0918_),
    .A1(_0905_),
    .A2(_0915_));
 sg13g2_or2_1 _1749_ (.X(_0243_),
    .B(_0918_),
    .A(_0917_));
 sg13g2_o21ai_1 _1750_ (.B1(_0914_),
    .Y(_0919_),
    .A1(_0904_),
    .A2(_0909_));
 sg13g2_nor2_1 _1751_ (.A(_0900_),
    .B(_0905_),
    .Y(_0920_));
 sg13g2_nor2_1 _1752_ (.A(_0905_),
    .B(_0909_),
    .Y(_0921_));
 sg13g2_nor2_1 _1753_ (.A(_0914_),
    .B(_0921_),
    .Y(_0922_));
 sg13g2_nand2_1 _1754_ (.Y(_0923_),
    .A(_0905_),
    .B(_0909_));
 sg13g2_nand2_1 _1755_ (.Y(_0924_),
    .A(_0922_),
    .B(_0923_));
 sg13g2_o21ai_1 _1756_ (.B1(_0919_),
    .Y(_0244_),
    .A1(_0920_),
    .A2(_0924_));
 sg13g2_nand3_1 _1757_ (.B(_0899_),
    .C(_0908_),
    .A(_0897_),
    .Y(_0925_));
 sg13g2_o21ai_1 _1758_ (.B1(_0925_),
    .Y(_0926_),
    .A1(_0917_),
    .A2(_0921_));
 sg13g2_o21ai_1 _1759_ (.B1(_0914_),
    .Y(_0927_),
    .A1(_0900_),
    .A2(_0923_));
 sg13g2_nand2_1 _1760_ (.Y(_0245_),
    .A(_0926_),
    .B(_0927_));
 sg13g2_or2_1 _1761_ (.X(_0928_),
    .B(_0919_),
    .A(_0900_));
 sg13g2_inv_1 _1762_ (.Y(_0249_),
    .A(_0928_));
 sg13g2_o21ai_1 _1763_ (.B1(_0923_),
    .Y(_0929_),
    .A1(_0900_),
    .A2(_0922_));
 sg13g2_a22oi_1 _1764_ (.Y(_0246_),
    .B1(_0928_),
    .B2(_0929_),
    .A2(_0915_),
    .A1(_0900_));
 sg13g2_a21oi_1 _1765_ (.A1(_0919_),
    .A2(_0925_),
    .Y(_0247_),
    .B1(_0916_));
 sg13g2_o21ai_1 _1766_ (.B1(_0909_),
    .Y(_0930_),
    .A1(_0900_),
    .A2(_0905_));
 sg13g2_and2_1 _1767_ (.A(_0914_),
    .B(_0930_),
    .X(_0248_));
 sg13g2_nor2_2 _1768_ (.A(_0915_),
    .B(_0925_),
    .Y(_0250_));
 sg13g2_nand2b_1 _1769_ (.Y(_0931_),
    .B(\noise_generator.lfsr[0] ),
    .A_N(noise_disable_B));
 sg13g2_o21ai_1 _1770_ (.B1(_0931_),
    .Y(_0932_),
    .A1(tone_B),
    .A2(tone_disable_B));
 sg13g2_nand2b_1 _1771_ (.Y(_0933_),
    .B(_0014_),
    .A_N(envelope_B));
 sg13g2_a21oi_1 _1772_ (.A1(envelope_B),
    .A2(_0895_),
    .Y(_0934_),
    .B1(_0932_));
 sg13g2_and2_1 _1773_ (.A(_0933_),
    .B(_0934_),
    .X(_0935_));
 sg13g2_nand2_2 _1774_ (.Y(_0936_),
    .A(_0933_),
    .B(_0934_));
 sg13g2_mux2_2 _1775_ (.A0(_0016_),
    .A1(_0901_),
    .S(envelope_B),
    .X(_0937_));
 sg13g2_nor2_2 _1776_ (.A(_0932_),
    .B(_0937_),
    .Y(_0938_));
 sg13g2_mux2_2 _1777_ (.A0(_0017_),
    .A1(_0906_),
    .S(envelope_B),
    .X(_0939_));
 sg13g2_nor2_1 _1778_ (.A(_0932_),
    .B(_0939_),
    .Y(_0940_));
 sg13g2_nor2b_1 _1779_ (.A(_0938_),
    .B_N(_0940_),
    .Y(_0941_));
 sg13g2_nand2b_1 _1780_ (.Y(_0942_),
    .B(_0015_),
    .A_N(envelope_B));
 sg13g2_a21oi_1 _1781_ (.A1(envelope_B),
    .A2(_0911_),
    .Y(_0943_),
    .B1(_0932_));
 sg13g2_and2_2 _1782_ (.A(_0942_),
    .B(_0943_),
    .X(_0944_));
 sg13g2_nand2_1 _1783_ (.Y(_0945_),
    .A(_0942_),
    .B(_0943_));
 sg13g2_nor2_1 _1784_ (.A(_0938_),
    .B(_0944_),
    .Y(_0946_));
 sg13g2_nand2_1 _1785_ (.Y(_0947_),
    .A(_0935_),
    .B(_0946_));
 sg13g2_a22oi_1 _1786_ (.Y(_0948_),
    .B1(_0944_),
    .B2(_0938_),
    .A2(_0941_),
    .A1(_0936_));
 sg13g2_nand2_1 _1787_ (.Y(_0251_),
    .A(_0947_),
    .B(_0948_));
 sg13g2_nand2b_1 _1788_ (.Y(_0949_),
    .B(_0944_),
    .A_N(_0941_));
 sg13g2_nor3_2 _1789_ (.A(_0932_),
    .B(_0937_),
    .C(_0939_),
    .Y(_0950_));
 sg13g2_a21oi_2 _1790_ (.B1(_0932_),
    .Y(_0951_),
    .A2(_0939_),
    .A1(_0937_));
 sg13g2_a21oi_1 _1791_ (.A1(_0935_),
    .A2(_0938_),
    .Y(_0952_),
    .B1(_0944_));
 sg13g2_nand2_1 _1792_ (.Y(_0953_),
    .A(_0951_),
    .B(_0952_));
 sg13g2_o21ai_1 _1793_ (.B1(_0949_),
    .Y(_0252_),
    .A1(_0950_),
    .A2(_0953_));
 sg13g2_nand2_1 _1794_ (.Y(_0954_),
    .A(_0935_),
    .B(_0940_));
 sg13g2_nor3_1 _1795_ (.A(_0936_),
    .B(_0944_),
    .C(_0951_),
    .Y(_0955_));
 sg13g2_a21oi_1 _1796_ (.A1(_0936_),
    .A2(_0950_),
    .Y(_0956_),
    .B1(_0955_));
 sg13g2_o21ai_1 _1797_ (.B1(_0944_),
    .Y(_0957_),
    .A1(_0936_),
    .A2(_0951_));
 sg13g2_nand2_1 _1798_ (.Y(_0253_),
    .A(_0956_),
    .B(_0957_));
 sg13g2_nor2_2 _1799_ (.A(_0936_),
    .B(_0949_),
    .Y(_0257_));
 sg13g2_nor2_1 _1800_ (.A(_0935_),
    .B(_0945_),
    .Y(_0958_));
 sg13g2_nor3_1 _1801_ (.A(_0936_),
    .B(_0944_),
    .C(_0950_),
    .Y(_0959_));
 sg13g2_o21ai_1 _1802_ (.B1(_0951_),
    .Y(_0960_),
    .A1(_0958_),
    .A2(_0959_));
 sg13g2_nand2b_1 _1803_ (.Y(_0254_),
    .B(_0960_),
    .A_N(_0257_));
 sg13g2_o21ai_1 _1804_ (.B1(_0949_),
    .Y(_0255_),
    .A1(_0946_),
    .A2(_0954_));
 sg13g2_a21oi_1 _1805_ (.A1(_0935_),
    .A2(_0938_),
    .Y(_0961_),
    .B1(_0940_));
 sg13g2_nor2_1 _1806_ (.A(_0945_),
    .B(_0961_),
    .Y(_0256_));
 sg13g2_nor2_1 _1807_ (.A(_0945_),
    .B(_0954_),
    .Y(_0258_));
 sg13g2_nand2b_1 _1808_ (.Y(_0962_),
    .B(\noise_generator.lfsr[0] ),
    .A_N(noise_disable_C));
 sg13g2_o21ai_1 _1809_ (.B1(_0962_),
    .Y(_0963_),
    .A1(tone_C),
    .A2(tone_disable_C));
 sg13g2_a21oi_1 _1810_ (.A1(envelope_C),
    .A2(_0895_),
    .Y(_0964_),
    .B1(_0963_));
 sg13g2_o21ai_1 _1811_ (.B1(_0964_),
    .Y(_0965_),
    .A1(_0819_),
    .A2(envelope_C));
 sg13g2_mux2_1 _1812_ (.A0(_0020_),
    .A1(_0901_),
    .S(envelope_C),
    .X(_0966_));
 sg13g2_nor2_2 _1813_ (.A(_0963_),
    .B(_0966_),
    .Y(_0967_));
 sg13g2_a21oi_1 _1814_ (.A1(envelope_C),
    .A2(_0906_),
    .Y(_0968_),
    .B1(_0963_));
 sg13g2_o21ai_1 _1815_ (.B1(_0968_),
    .Y(_0969_),
    .A1(envelope_C),
    .A2(_0820_));
 sg13g2_inv_1 _1816_ (.Y(_0970_),
    .A(_0969_));
 sg13g2_nor2_1 _1817_ (.A(_0967_),
    .B(_0969_),
    .Y(_0971_));
 sg13g2_nand2b_1 _1818_ (.Y(_0972_),
    .B(_0019_),
    .A_N(envelope_C));
 sg13g2_a21oi_1 _1819_ (.A1(envelope_C),
    .A2(_0911_),
    .Y(_0973_),
    .B1(_0963_));
 sg13g2_and2_1 _1820_ (.A(_0972_),
    .B(_0973_),
    .X(_0974_));
 sg13g2_nand2_2 _1821_ (.Y(_0975_),
    .A(_0972_),
    .B(_0973_));
 sg13g2_nor2_1 _1822_ (.A(_0967_),
    .B(_0974_),
    .Y(_0976_));
 sg13g2_nand2b_1 _1823_ (.Y(_0977_),
    .B(_0975_),
    .A_N(_0965_));
 sg13g2_a22oi_1 _1824_ (.Y(_0978_),
    .B1(_0974_),
    .B2(_0967_),
    .A2(_0971_),
    .A1(_0965_));
 sg13g2_o21ai_1 _1825_ (.B1(_0978_),
    .Y(_0259_),
    .A1(_0967_),
    .A2(_0977_));
 sg13g2_o21ai_1 _1826_ (.B1(_0974_),
    .Y(_0979_),
    .A1(_0967_),
    .A2(_0969_));
 sg13g2_nor2b_1 _1827_ (.A(_0965_),
    .B_N(_0967_),
    .Y(_0980_));
 sg13g2_nand2b_1 _1828_ (.Y(_0981_),
    .B(_0969_),
    .A_N(_0967_));
 sg13g2_a21oi_1 _1829_ (.A1(_0967_),
    .A2(_0970_),
    .Y(_0982_),
    .B1(_0974_));
 sg13g2_inv_1 _1830_ (.Y(_0983_),
    .A(_0982_));
 sg13g2_nand2_1 _1831_ (.Y(_0984_),
    .A(_0981_),
    .B(_0982_));
 sg13g2_o21ai_1 _1832_ (.B1(_0979_),
    .Y(_0260_),
    .A1(_0980_),
    .A2(_0984_));
 sg13g2_a22oi_1 _1833_ (.Y(_0985_),
    .B1(_0983_),
    .B2(_0965_),
    .A2(_0981_),
    .A1(_0974_));
 sg13g2_o21ai_1 _1834_ (.B1(_0985_),
    .Y(_0261_),
    .A1(_0977_),
    .A2(_0981_));
 sg13g2_nor2_1 _1835_ (.A(_0965_),
    .B(_0979_),
    .Y(_0265_));
 sg13g2_a21oi_1 _1836_ (.A1(_0965_),
    .A2(_0981_),
    .Y(_0986_),
    .B1(_0265_));
 sg13g2_a22oi_1 _1837_ (.Y(_0262_),
    .B1(_0984_),
    .B2(_0986_),
    .A2(_0975_),
    .A1(_0965_));
 sg13g2_or2_1 _1838_ (.X(_0987_),
    .B(_0969_),
    .A(_0965_));
 sg13g2_o21ai_1 _1839_ (.B1(_0979_),
    .Y(_0263_),
    .A1(_0976_),
    .A2(_0987_));
 sg13g2_nor2_1 _1840_ (.A(_0970_),
    .B(_0980_),
    .Y(_0988_));
 sg13g2_nor2_1 _1841_ (.A(_0975_),
    .B(_0988_),
    .Y(_0264_));
 sg13g2_nor2_1 _1842_ (.A(_0975_),
    .B(_0987_),
    .Y(_0266_));
 sg13g2_nand4_1 _1843_ (.B(net185),
    .C(_0815_),
    .A(active),
    .Y(_0989_),
    .D(net6));
 sg13g2_nor3_2 _1844_ (.A(\latched_register[1] ),
    .B(_0781_),
    .C(_0989_),
    .Y(_0990_));
 sg13g2_and3_2 _1845_ (.X(_0024_),
    .A(net598),
    .B(net595),
    .C(_0990_));
 sg13g2_nor2_2 _1846_ (.A(\latched_register[3] ),
    .B(\latched_register[2] ),
    .Y(_0991_));
 sg13g2_and2_2 _1847_ (.A(_0990_),
    .B(_0991_),
    .X(_0992_));
 sg13g2_nor2_2 _1848_ (.A(net162),
    .B(_0992_),
    .Y(_0993_));
 sg13g2_a22oi_1 _1849_ (.Y(_0994_),
    .B1(_0993_),
    .B2(net468),
    .A2(_0992_),
    .A1(net175));
 sg13g2_inv_1 _1850_ (.Y(_0025_),
    .A(_0994_));
 sg13g2_a22oi_1 _1851_ (.Y(_0995_),
    .B1(_0993_),
    .B2(net351),
    .A2(_0992_),
    .A1(net173));
 sg13g2_inv_1 _1852_ (.Y(_0026_),
    .A(_0995_));
 sg13g2_a22oi_1 _1853_ (.Y(_0996_),
    .B1(_0993_),
    .B2(net386),
    .A2(_0992_),
    .A1(net171));
 sg13g2_inv_1 _1854_ (.Y(_0027_),
    .A(_0996_));
 sg13g2_a22oi_1 _1855_ (.Y(_0997_),
    .B1(_0993_),
    .B2(net425),
    .A2(_0992_),
    .A1(net169));
 sg13g2_inv_1 _1856_ (.Y(_0028_),
    .A(_0997_));
 sg13g2_nor3_2 _1857_ (.A(_0780_),
    .B(\latched_register[0] ),
    .C(_0989_),
    .Y(_0998_));
 sg13g2_and2_1 _1858_ (.A(_0991_),
    .B(_0998_),
    .X(_0999_));
 sg13g2_nor2_2 _1859_ (.A(net164),
    .B(net152),
    .Y(_1000_));
 sg13g2_a22oi_1 _1860_ (.Y(_1001_),
    .B1(_1000_),
    .B2(net411),
    .A2(net152),
    .A1(net176));
 sg13g2_inv_1 _1861_ (.Y(_0029_),
    .A(_1001_));
 sg13g2_a22oi_1 _1862_ (.Y(_1002_),
    .B1(_1000_),
    .B2(net424),
    .A2(net152),
    .A1(net174));
 sg13g2_inv_1 _1863_ (.Y(_0030_),
    .A(_1002_));
 sg13g2_a22oi_1 _1864_ (.Y(_1003_),
    .B1(_1000_),
    .B2(net400),
    .A2(net152),
    .A1(net172));
 sg13g2_inv_1 _1865_ (.Y(_0031_),
    .A(_1003_));
 sg13g2_a22oi_1 _1866_ (.Y(_1004_),
    .B1(_1000_),
    .B2(net404),
    .A2(net152),
    .A1(net170));
 sg13g2_inv_1 _1867_ (.Y(_0032_),
    .A(_1004_));
 sg13g2_a22oi_1 _1868_ (.Y(_1005_),
    .B1(_1000_),
    .B2(net379),
    .A2(_0999_),
    .A1(net168));
 sg13g2_inv_1 _1869_ (.Y(_0033_),
    .A(_1005_));
 sg13g2_a22oi_1 _1870_ (.Y(_1006_),
    .B1(_1000_),
    .B2(net438),
    .A2(net152),
    .A1(net2));
 sg13g2_inv_1 _1871_ (.Y(_0034_),
    .A(_1006_));
 sg13g2_a22oi_1 _1872_ (.Y(_1007_),
    .B1(_1000_),
    .B2(net370),
    .A2(net152),
    .A1(net3));
 sg13g2_inv_1 _1873_ (.Y(_0035_),
    .A(_1007_));
 sg13g2_a22oi_1 _1874_ (.Y(_1008_),
    .B1(_1000_),
    .B2(net410),
    .A2(net152),
    .A1(net4));
 sg13g2_inv_1 _1875_ (.Y(_0036_),
    .A(_1008_));
 sg13g2_nor2_2 _1876_ (.A(\latched_register[3] ),
    .B(_0779_),
    .Y(_1009_));
 sg13g2_and2_2 _1877_ (.A(_0998_),
    .B(_1009_),
    .X(_1010_));
 sg13g2_nor2_2 _1878_ (.A(net162),
    .B(_1010_),
    .Y(_1011_));
 sg13g2_a22oi_1 _1879_ (.Y(_1012_),
    .B1(_1011_),
    .B2(net361),
    .A2(_1010_),
    .A1(net175));
 sg13g2_inv_1 _1880_ (.Y(_0037_),
    .A(_1012_));
 sg13g2_a22oi_1 _1881_ (.Y(_1013_),
    .B1(_1011_),
    .B2(net423),
    .A2(_1010_),
    .A1(net173));
 sg13g2_inv_1 _1882_ (.Y(_0038_),
    .A(_1013_));
 sg13g2_a22oi_1 _1883_ (.Y(_1014_),
    .B1(_1011_),
    .B2(net415),
    .A2(_1010_),
    .A1(net171));
 sg13g2_inv_1 _1884_ (.Y(_0039_),
    .A(_1014_));
 sg13g2_a22oi_1 _1885_ (.Y(_1015_),
    .B1(_1011_),
    .B2(net437),
    .A2(_1010_),
    .A1(net169));
 sg13g2_inv_1 _1886_ (.Y(_0040_),
    .A(_1015_));
 sg13g2_a22oi_1 _1887_ (.Y(_1016_),
    .B1(_1011_),
    .B2(net401),
    .A2(_1010_),
    .A1(net168));
 sg13g2_inv_1 _1888_ (.Y(_0041_),
    .A(_1016_));
 sg13g2_and2_2 _1889_ (.A(_0990_),
    .B(_1009_),
    .X(_1017_));
 sg13g2_nor2_2 _1890_ (.A(net162),
    .B(_1017_),
    .Y(_1018_));
 sg13g2_a22oi_1 _1891_ (.Y(_1019_),
    .B1(_1018_),
    .B2(net441),
    .A2(_1017_),
    .A1(net175));
 sg13g2_inv_1 _1892_ (.Y(_0042_),
    .A(_1019_));
 sg13g2_a22oi_1 _1893_ (.Y(_1020_),
    .B1(_1018_),
    .B2(net461),
    .A2(_1017_),
    .A1(net173));
 sg13g2_inv_1 _1894_ (.Y(_0043_),
    .A(_1020_));
 sg13g2_a22oi_1 _1895_ (.Y(_1021_),
    .B1(_1018_),
    .B2(net440),
    .A2(_1017_),
    .A1(net171));
 sg13g2_inv_1 _1896_ (.Y(_0044_),
    .A(_1021_));
 sg13g2_a22oi_1 _1897_ (.Y(_1022_),
    .B1(_1018_),
    .B2(net494),
    .A2(_1017_),
    .A1(net169));
 sg13g2_inv_1 _1898_ (.Y(_0045_),
    .A(_1022_));
 sg13g2_xor2_1 _1899_ (.B(_0862_),
    .A(\attenuation_C.out[0] ),
    .X(_1023_));
 sg13g2_or2_1 _1900_ (.X(_1024_),
    .B(_1023_),
    .A(net572));
 sg13g2_nand2_1 _1901_ (.Y(_1025_),
    .A(net572),
    .B(_1023_));
 sg13g2_and3_1 _1902_ (.X(_0046_),
    .A(net183),
    .B(_1024_),
    .C(_1025_));
 sg13g2_or2_1 _1903_ (.X(_1026_),
    .B(_0885_),
    .A(_0821_));
 sg13g2_xnor2_1 _1904_ (.Y(_1027_),
    .A(_0821_),
    .B(_0885_));
 sg13g2_o21ai_1 _1905_ (.B1(net183),
    .Y(_1028_),
    .A1(_1025_),
    .A2(_1027_));
 sg13g2_a21oi_1 _1906_ (.A1(_1025_),
    .A2(_1027_),
    .Y(_0047_),
    .B1(_1028_));
 sg13g2_o21ai_1 _1907_ (.B1(_1026_),
    .Y(_1029_),
    .A1(_1025_),
    .A2(_1027_));
 sg13g2_and2_1 _1908_ (.A(net628),
    .B(_0886_),
    .X(_1030_));
 sg13g2_or2_1 _1909_ (.X(_1031_),
    .B(_0886_),
    .A(net628));
 sg13g2_nor2b_1 _1910_ (.A(_1030_),
    .B_N(_1031_),
    .Y(_1032_));
 sg13g2_o21ai_1 _1911_ (.B1(net183),
    .Y(_1033_),
    .A1(_1029_),
    .A2(_1032_));
 sg13g2_a21oi_1 _1912_ (.A1(_1029_),
    .A2(_1032_),
    .Y(_0048_),
    .B1(_1033_));
 sg13g2_a21oi_1 _1913_ (.A1(_1029_),
    .A2(_1031_),
    .Y(_1034_),
    .B1(_1030_));
 sg13g2_nand2_1 _1914_ (.Y(_1035_),
    .A(net605),
    .B(_0888_));
 sg13g2_xnor2_1 _1915_ (.Y(_1036_),
    .A(net605),
    .B(_0888_));
 sg13g2_o21ai_1 _1916_ (.B1(net183),
    .Y(_1037_),
    .A1(_1034_),
    .A2(_1036_));
 sg13g2_a21oi_1 _1917_ (.A1(_1034_),
    .A2(_1036_),
    .Y(_0049_),
    .B1(_1037_));
 sg13g2_o21ai_1 _1918_ (.B1(_1035_),
    .Y(_1038_),
    .A1(_1034_),
    .A2(_1036_));
 sg13g2_nor2_1 _1919_ (.A(_0822_),
    .B(_0889_),
    .Y(_1039_));
 sg13g2_nand2_1 _1920_ (.Y(_1040_),
    .A(_0822_),
    .B(_0889_));
 sg13g2_nor2b_1 _1921_ (.A(_1039_),
    .B_N(_1040_),
    .Y(_1041_));
 sg13g2_o21ai_1 _1922_ (.B1(net182),
    .Y(_1042_),
    .A1(_1038_),
    .A2(_1041_));
 sg13g2_a21oi_1 _1923_ (.A1(_1038_),
    .A2(_1041_),
    .Y(_0050_),
    .B1(_1042_));
 sg13g2_a21oi_1 _1924_ (.A1(_1038_),
    .A2(_1040_),
    .Y(_1043_),
    .B1(_1039_));
 sg13g2_or2_1 _1925_ (.X(_1044_),
    .B(_0890_),
    .A(_0823_));
 sg13g2_xnor2_1 _1926_ (.Y(_1045_),
    .A(_0823_),
    .B(_0890_));
 sg13g2_o21ai_1 _1927_ (.B1(net182),
    .Y(_1046_),
    .A1(_1043_),
    .A2(_1045_));
 sg13g2_a21oi_1 _1928_ (.A1(_1043_),
    .A2(_1045_),
    .Y(_0051_),
    .B1(_1046_));
 sg13g2_o21ai_1 _1929_ (.B1(_1044_),
    .Y(_1047_),
    .A1(_1043_),
    .A2(_1045_));
 sg13g2_and2_1 _1930_ (.A(\pwm_master.accumulator[6] ),
    .B(_0892_),
    .X(_1048_));
 sg13g2_nand2_1 _1931_ (.Y(_1049_),
    .A(\pwm_master.accumulator[6] ),
    .B(_0892_));
 sg13g2_xnor2_1 _1932_ (.Y(_1050_),
    .A(net635),
    .B(_0892_));
 sg13g2_inv_1 _1933_ (.Y(_1051_),
    .A(_1050_));
 sg13g2_xnor2_1 _1934_ (.Y(_1052_),
    .A(_1047_),
    .B(_1051_));
 sg13g2_nor2_1 _1935_ (.A(net165),
    .B(_1052_),
    .Y(_0052_));
 sg13g2_a21oi_1 _1936_ (.A1(_0882_),
    .A2(_0893_),
    .Y(_1053_),
    .B1(net622));
 sg13g2_xnor2_1 _1937_ (.Y(_1054_),
    .A(_0824_),
    .B(_0894_));
 sg13g2_a21oi_1 _1938_ (.A1(_1047_),
    .A2(_1051_),
    .Y(_1055_),
    .B1(_1048_));
 sg13g2_o21ai_1 _1939_ (.B1(net183),
    .Y(_1056_),
    .A1(_1054_),
    .A2(_1055_));
 sg13g2_a21oi_1 _1940_ (.A1(_1054_),
    .A2(_1055_),
    .Y(_0053_),
    .B1(_1056_));
 sg13g2_nand3_1 _1941_ (.B(_0883_),
    .C(uo_out[7]),
    .A(net568),
    .Y(_1057_));
 sg13g2_a21o_1 _1942_ (.A2(uo_out[7]),
    .A1(_0883_),
    .B1(net629),
    .X(_1058_));
 sg13g2_nand2_1 _1943_ (.Y(_1059_),
    .A(_1057_),
    .B(_1058_));
 sg13g2_o21ai_1 _1944_ (.B1(_1049_),
    .Y(_1060_),
    .A1(_0824_),
    .A2(_0894_));
 sg13g2_a21oi_1 _1945_ (.A1(_1047_),
    .A2(_1051_),
    .Y(_1061_),
    .B1(_1060_));
 sg13g2_o21ai_1 _1946_ (.B1(_1059_),
    .Y(_1062_),
    .A1(_1053_),
    .A2(_1061_));
 sg13g2_or3_1 _1947_ (.A(_1053_),
    .B(_1059_),
    .C(_1061_),
    .X(_1063_));
 sg13g2_and3_1 _1948_ (.X(_0054_),
    .A(net182),
    .B(_1062_),
    .C(_1063_));
 sg13g2_a21oi_1 _1949_ (.A1(_1057_),
    .A2(_1063_),
    .Y(_0055_),
    .B1(net165));
 sg13g2_nor4_1 _1950_ (.A(net4),
    .B(net3),
    .C(net2),
    .D(net1),
    .Y(_1064_));
 sg13g2_nand3_1 _1951_ (.B(net6),
    .C(_1064_),
    .A(net5),
    .Y(_1065_));
 sg13g2_o21ai_1 _1952_ (.B1(net181),
    .Y(_1066_),
    .A1(net175),
    .A2(net160));
 sg13g2_a21oi_1 _1953_ (.A1(_0781_),
    .A2(net160),
    .Y(_0056_),
    .B1(_1066_));
 sg13g2_o21ai_1 _1954_ (.B1(net181),
    .Y(_1067_),
    .A1(net173),
    .A2(net160));
 sg13g2_a21oi_1 _1955_ (.A1(_0780_),
    .A2(net160),
    .Y(_0057_),
    .B1(_1067_));
 sg13g2_o21ai_1 _1956_ (.B1(net181),
    .Y(_1068_),
    .A1(net171),
    .A2(net160));
 sg13g2_a21oi_1 _1957_ (.A1(_0779_),
    .A2(net160),
    .Y(_0058_),
    .B1(_1068_));
 sg13g2_o21ai_1 _1958_ (.B1(net180),
    .Y(_1069_),
    .A1(net169),
    .A2(net160));
 sg13g2_a21oi_1 _1959_ (.A1(_0778_),
    .A2(net160),
    .Y(_0059_),
    .B1(_1069_));
 sg13g2_o21ai_1 _1960_ (.B1(net448),
    .Y(_1070_),
    .A1(_0815_),
    .A2(_0816_));
 sg13g2_a21oi_1 _1961_ (.A1(_1065_),
    .A2(_1070_),
    .Y(_0060_),
    .B1(net167));
 sg13g2_and2_1 _1962_ (.A(net185),
    .B(net333),
    .X(_0061_));
 sg13g2_xnor2_1 _1963_ (.Y(_1071_),
    .A(\clk_counter[1] ),
    .B(net549));
 sg13g2_nor2_1 _1964_ (.A(net166),
    .B(net550),
    .Y(_0062_));
 sg13g2_a21oi_1 _1965_ (.A1(\clk_counter[1] ),
    .A2(\clk_counter[0] ),
    .Y(_1072_),
    .B1(net418));
 sg13g2_nand3_1 _1966_ (.B(net549),
    .C(net418),
    .A(\clk_counter[1] ),
    .Y(_1073_));
 sg13g2_nand2_1 _1967_ (.Y(_1074_),
    .A(net185),
    .B(_1073_));
 sg13g2_nor2_1 _1968_ (.A(net419),
    .B(_1074_),
    .Y(_0063_));
 sg13g2_nor2_1 _1969_ (.A(_0782_),
    .B(_1073_),
    .Y(_1075_));
 sg13g2_a21oi_1 _1970_ (.A1(_0782_),
    .A2(_1073_),
    .Y(_1076_),
    .B1(net166));
 sg13g2_nor2b_1 _1971_ (.A(_1075_),
    .B_N(net594),
    .Y(_0064_));
 sg13g2_nor2_1 _1972_ (.A(net527),
    .B(_1075_),
    .Y(_1077_));
 sg13g2_and2_1 _1973_ (.A(net527),
    .B(_1075_),
    .X(_1078_));
 sg13g2_nor3_1 _1974_ (.A(net166),
    .B(net528),
    .C(_1078_),
    .Y(_0065_));
 sg13g2_nand2_1 _1975_ (.Y(_1079_),
    .A(net567),
    .B(_1078_));
 sg13g2_o21ai_1 _1976_ (.B1(net185),
    .Y(_1080_),
    .A1(net567),
    .A2(_1078_));
 sg13g2_nor2b_1 _1977_ (.A(_1080_),
    .B_N(_1079_),
    .Y(_0066_));
 sg13g2_o21ai_1 _1978_ (.B1(net185),
    .Y(_1081_),
    .A1(_0783_),
    .A2(_1079_));
 sg13g2_a21oi_1 _1979_ (.A1(_0783_),
    .A2(_1079_),
    .Y(_0067_),
    .B1(_1081_));
 sg13g2_nor2_2 _1980_ (.A(net166),
    .B(_0024_),
    .Y(_1082_));
 sg13g2_a22oi_1 _1981_ (.Y(_1083_),
    .B1(_1082_),
    .B2(net506),
    .A2(_0024_),
    .A1(net176));
 sg13g2_inv_1 _1982_ (.Y(_0068_),
    .A(_1083_));
 sg13g2_a22oi_1 _1983_ (.Y(_1084_),
    .B1(_1082_),
    .B2(net394),
    .A2(_0024_),
    .A1(net174));
 sg13g2_inv_1 _1984_ (.Y(_0069_),
    .A(_1084_));
 sg13g2_a22oi_1 _1985_ (.Y(_1085_),
    .B1(_1082_),
    .B2(net354),
    .A2(_0024_),
    .A1(net172));
 sg13g2_inv_1 _1986_ (.Y(_0070_),
    .A(_1085_));
 sg13g2_a22oi_1 _1987_ (.Y(_1086_),
    .B1(_1082_),
    .B2(net476),
    .A2(_0024_),
    .A1(net170));
 sg13g2_inv_1 _1988_ (.Y(_0071_),
    .A(_1086_));
 sg13g2_nor3_2 _1989_ (.A(\latched_register[1] ),
    .B(\latched_register[0] ),
    .C(_0989_),
    .Y(_1087_));
 sg13g2_and3_2 _1990_ (.X(_1088_),
    .A(\latched_register[3] ),
    .B(net638),
    .C(_1087_));
 sg13g2_nor2_2 _1991_ (.A(net167),
    .B(net151),
    .Y(_1089_));
 sg13g2_a22oi_1 _1992_ (.Y(_1090_),
    .B1(_1089_),
    .B2(net439),
    .A2(net151),
    .A1(net176));
 sg13g2_inv_1 _1993_ (.Y(_0072_),
    .A(_1090_));
 sg13g2_a22oi_1 _1994_ (.Y(_1091_),
    .B1(_1089_),
    .B2(net381),
    .A2(net151),
    .A1(net174));
 sg13g2_inv_1 _1995_ (.Y(_0073_),
    .A(_1091_));
 sg13g2_a22oi_1 _1996_ (.Y(_1092_),
    .B1(_1089_),
    .B2(net466),
    .A2(net151),
    .A1(net172));
 sg13g2_inv_1 _1997_ (.Y(_0074_),
    .A(_1092_));
 sg13g2_a22oi_1 _1998_ (.Y(_1093_),
    .B1(_1089_),
    .B2(net371),
    .A2(net639),
    .A1(net170));
 sg13g2_inv_1 _1999_ (.Y(_0075_),
    .A(_1093_));
 sg13g2_a22oi_1 _2000_ (.Y(_1094_),
    .B1(_1089_),
    .B2(net392),
    .A2(net151),
    .A1(net1));
 sg13g2_inv_1 _2001_ (.Y(_0076_),
    .A(_1094_));
 sg13g2_a22oi_1 _2002_ (.Y(_1095_),
    .B1(_1089_),
    .B2(net407),
    .A2(net151),
    .A1(net2));
 sg13g2_inv_1 _2003_ (.Y(_0077_),
    .A(_1095_));
 sg13g2_a22oi_1 _2004_ (.Y(_1096_),
    .B1(_1089_),
    .B2(net477),
    .A2(net151),
    .A1(net3));
 sg13g2_inv_1 _2005_ (.Y(_0078_),
    .A(_1096_));
 sg13g2_a22oi_1 _2006_ (.Y(_1097_),
    .B1(_1089_),
    .B2(net412),
    .A2(net151),
    .A1(net4));
 sg13g2_inv_1 _2007_ (.Y(_0079_),
    .A(_1097_));
 sg13g2_nor2_2 _2008_ (.A(_0778_),
    .B(\latched_register[2] ),
    .Y(_1098_));
 sg13g2_and2_2 _2009_ (.A(_0998_),
    .B(_1098_),
    .X(_1099_));
 sg13g2_nor2_2 _2010_ (.A(net166),
    .B(_1099_),
    .Y(_1100_));
 sg13g2_a22oi_1 _2011_ (.Y(_1101_),
    .B1(_1100_),
    .B2(net345),
    .A2(_1099_),
    .A1(net176));
 sg13g2_inv_1 _2012_ (.Y(_0080_),
    .A(_1101_));
 sg13g2_a22oi_1 _2013_ (.Y(_1102_),
    .B1(_1100_),
    .B2(net358),
    .A2(_1099_),
    .A1(net174));
 sg13g2_inv_1 _2014_ (.Y(_0081_),
    .A(_1102_));
 sg13g2_a22oi_1 _2015_ (.Y(_1103_),
    .B1(_1100_),
    .B2(net352),
    .A2(_1099_),
    .A1(net172));
 sg13g2_inv_1 _2016_ (.Y(_0082_),
    .A(_1103_));
 sg13g2_a22oi_1 _2017_ (.Y(_0267_),
    .B1(_1100_),
    .B2(net346),
    .A2(_1099_),
    .A1(net170));
 sg13g2_inv_1 _2018_ (.Y(_0083_),
    .A(_0267_));
 sg13g2_a22oi_1 _2019_ (.Y(_0268_),
    .B1(_1100_),
    .B2(net589),
    .A2(_1099_),
    .A1(net1));
 sg13g2_inv_1 _2020_ (.Y(_0084_),
    .A(_0268_));
 sg13g2_nor3_2 _2021_ (.A(_0780_),
    .B(_0781_),
    .C(_0989_),
    .Y(_0269_));
 sg13g2_and2_1 _2022_ (.A(_1098_),
    .B(_0269_),
    .X(_0270_));
 sg13g2_nor2_2 _2023_ (.A(net166),
    .B(net150),
    .Y(_0271_));
 sg13g2_a22oi_1 _2024_ (.Y(_0272_),
    .B1(_0271_),
    .B2(net378),
    .A2(net150),
    .A1(net176));
 sg13g2_inv_1 _2025_ (.Y(_0085_),
    .A(_0272_));
 sg13g2_a22oi_1 _2026_ (.Y(_0273_),
    .B1(_0271_),
    .B2(net403),
    .A2(net150),
    .A1(net174));
 sg13g2_inv_1 _2027_ (.Y(_0086_),
    .A(_0273_));
 sg13g2_a22oi_1 _2028_ (.Y(_0274_),
    .B1(_0271_),
    .B2(net402),
    .A2(net150),
    .A1(net172));
 sg13g2_inv_1 _2029_ (.Y(_0087_),
    .A(_0274_));
 sg13g2_a22oi_1 _2030_ (.Y(_0275_),
    .B1(_0271_),
    .B2(net426),
    .A2(net150),
    .A1(net170));
 sg13g2_inv_1 _2031_ (.Y(_0088_),
    .A(_0275_));
 sg13g2_a22oi_1 _2032_ (.Y(_0276_),
    .B1(_0271_),
    .B2(net422),
    .A2(net150),
    .A1(net168));
 sg13g2_inv_1 _2033_ (.Y(_0089_),
    .A(_0276_));
 sg13g2_a22oi_1 _2034_ (.Y(_0277_),
    .B1(_0271_),
    .B2(net364),
    .A2(_0270_),
    .A1(net2));
 sg13g2_inv_1 _2035_ (.Y(_0090_),
    .A(_0277_));
 sg13g2_a22oi_1 _2036_ (.Y(_0278_),
    .B1(_0271_),
    .B2(net479),
    .A2(net150),
    .A1(net3));
 sg13g2_inv_1 _2037_ (.Y(_0091_),
    .A(_0278_));
 sg13g2_a22oi_1 _2038_ (.Y(_0279_),
    .B1(_0271_),
    .B2(net393),
    .A2(net150),
    .A1(net4));
 sg13g2_inv_1 _2039_ (.Y(_0092_),
    .A(_0279_));
 sg13g2_or3_1 _2040_ (.A(\clk_counter[1] ),
    .B(\clk_counter[0] ),
    .C(\clk_counter[2] ),
    .X(_0280_));
 sg13g2_nand2b_1 _2041_ (.Y(_0281_),
    .B(net7),
    .A_N(net8));
 sg13g2_or4_1 _2042_ (.A(\clk_counter[3] ),
    .B(\clk_counter[5] ),
    .C(\clk_counter[4] ),
    .D(\clk_counter[6] ),
    .X(_0282_));
 sg13g2_nor2b_1 _2043_ (.A(net7),
    .B_N(net8),
    .Y(_0283_));
 sg13g2_a22oi_1 _2044_ (.Y(_0284_),
    .B1(_0282_),
    .B2(_0283_),
    .A2(_0281_),
    .A1(_0280_));
 sg13g2_inv_4 _2045_ (.A(_0284_),
    .Y(_0285_));
 sg13g2_a22oi_1 _2046_ (.Y(_0286_),
    .B1(\register[0][7] ),
    .B2(_0772_),
    .A2(\register[1][0] ),
    .A1(_0771_));
 sg13g2_nor2_1 _2047_ (.A(_0773_),
    .B(\register[0][5] ),
    .Y(_0287_));
 sg13g2_a21oi_1 _2048_ (.A1(\tone_A_generator.counter[6] ),
    .A2(_0810_),
    .Y(_0288_),
    .B1(_0287_));
 sg13g2_a22oi_1 _2049_ (.Y(_0289_),
    .B1(\register[0][4] ),
    .B2(_0774_),
    .A2(\register[0][5] ),
    .A1(_0773_));
 sg13g2_a22oi_1 _2050_ (.Y(_0290_),
    .B1(_0812_),
    .B2(\tone_A_generator.counter[3] ),
    .A2(_0811_),
    .A1(\tone_A_generator.counter[4] ));
 sg13g2_nand2b_1 _2051_ (.Y(_0291_),
    .B(\tone_A_generator.counter[0] ),
    .A_N(\register[0][0] ));
 sg13g2_o21ai_1 _2052_ (.B1(_0291_),
    .Y(_0292_),
    .A1(_0776_),
    .A2(\register[0][1] ));
 sg13g2_a22oi_1 _2053_ (.Y(_0293_),
    .B1(\register[0][1] ),
    .B2(_0776_),
    .A2(\register[0][2] ),
    .A1(_0775_));
 sg13g2_a22oi_1 _2054_ (.Y(_0294_),
    .B1(_0292_),
    .B2(_0293_),
    .A2(_0813_),
    .A1(\tone_A_generator.counter[2] ));
 sg13g2_nor2_1 _2055_ (.A(\tone_A_generator.counter[3] ),
    .B(_0812_),
    .Y(_0295_));
 sg13g2_o21ai_1 _2056_ (.B1(_0290_),
    .Y(_0296_),
    .A1(_0294_),
    .A2(_0295_));
 sg13g2_a221oi_1 _2057_ (.B2(_0296_),
    .C1(_0287_),
    .B1(_0289_),
    .A1(\tone_A_generator.counter[6] ),
    .Y(_0297_),
    .A2(_0810_));
 sg13g2_nor2_1 _2058_ (.A(\tone_A_generator.counter[6] ),
    .B(_0810_),
    .Y(_0298_));
 sg13g2_nand2b_1 _2059_ (.Y(_0299_),
    .B(\register[0][6] ),
    .A_N(\tone_A_generator.counter[6] ));
 sg13g2_nand2b_1 _2060_ (.Y(_0300_),
    .B(\tone_A_generator.counter[7] ),
    .A_N(\register[0][7] ));
 sg13g2_o21ai_1 _2061_ (.B1(_0300_),
    .Y(_0301_),
    .A1(_0297_),
    .A2(_0298_));
 sg13g2_a22oi_1 _2062_ (.Y(_0302_),
    .B1(_0286_),
    .B2(_0301_),
    .A2(_0809_),
    .A1(\tone_A_generator.counter[8] ));
 sg13g2_nor2_1 _2063_ (.A(\tone_A_generator.counter[9] ),
    .B(_0808_),
    .Y(_0303_));
 sg13g2_a22oi_1 _2064_ (.Y(_0304_),
    .B1(_0808_),
    .B2(\tone_A_generator.counter[9] ),
    .A2(_0807_),
    .A1(\tone_A_generator.counter[10] ));
 sg13g2_o21ai_1 _2065_ (.B1(_0304_),
    .Y(_0305_),
    .A1(_0302_),
    .A2(_0303_));
 sg13g2_a22oi_1 _2066_ (.Y(_0306_),
    .B1(\register[1][2] ),
    .B2(_0770_),
    .A2(\register[1][3] ),
    .A1(_0769_));
 sg13g2_nor2b_1 _2067_ (.A(_0292_),
    .B_N(_0306_),
    .Y(_0307_));
 sg13g2_nand3_1 _2068_ (.B(_0304_),
    .C(_0307_),
    .A(_0293_),
    .Y(_0308_));
 sg13g2_nand4_1 _2069_ (.B(_0288_),
    .C(_0289_),
    .A(_0286_),
    .Y(_0309_),
    .D(_0290_));
 sg13g2_a221oi_1 _2070_ (.B2(_0777_),
    .C1(_0303_),
    .B1(\register[0][0] ),
    .A1(\tone_A_generator.counter[8] ),
    .Y(_0310_),
    .A2(_0809_));
 sg13g2_a21oi_1 _2071_ (.A1(\tone_A_generator.counter[2] ),
    .A2(_0813_),
    .Y(_0311_),
    .B1(_0295_));
 sg13g2_nand4_1 _2072_ (.B(_0300_),
    .C(_0310_),
    .A(_0299_),
    .Y(_0312_),
    .D(_0311_));
 sg13g2_nor3_1 _2073_ (.A(_0308_),
    .B(_0309_),
    .C(_0312_),
    .Y(_0313_));
 sg13g2_a221oi_1 _2074_ (.B2(_0306_),
    .C1(_0313_),
    .B1(_0305_),
    .A1(\tone_A_generator.counter[11] ),
    .Y(_0314_),
    .A2(_0806_));
 sg13g2_nand2b_2 _2075_ (.Y(_0315_),
    .B(net158),
    .A_N(_0314_));
 sg13g2_nor2b_1 _2076_ (.A(tone_A),
    .B_N(_0315_),
    .Y(_0316_));
 sg13g2_nor2_1 _2077_ (.A(net382),
    .B(_0315_),
    .Y(_0317_));
 sg13g2_o21ai_1 _2078_ (.B1(net181),
    .Y(_0093_),
    .A1(_0316_),
    .A2(_0317_));
 sg13g2_nand2_1 _2079_ (.Y(_0318_),
    .A(net180),
    .B(_0315_));
 sg13g2_xnor2_1 _2080_ (.Y(_0319_),
    .A(net602),
    .B(net158));
 sg13g2_nand3_1 _2081_ (.B(_0315_),
    .C(_0319_),
    .A(net180),
    .Y(_0094_));
 sg13g2_nor3_2 _2082_ (.A(_0776_),
    .B(_0777_),
    .C(_0285_),
    .Y(_0320_));
 sg13g2_a21oi_1 _2083_ (.A1(\tone_A_generator.counter[0] ),
    .A2(net158),
    .Y(_0321_),
    .B1(net384));
 sg13g2_nor3_1 _2084_ (.A(net145),
    .B(_0320_),
    .C(net385),
    .Y(_0095_));
 sg13g2_and2_1 _2085_ (.A(net565),
    .B(_0320_),
    .X(_0322_));
 sg13g2_nor2_1 _2086_ (.A(net565),
    .B(_0320_),
    .Y(_0323_));
 sg13g2_nor3_1 _2087_ (.A(_0318_),
    .B(_0322_),
    .C(net566),
    .Y(_0096_));
 sg13g2_and2_1 _2088_ (.A(net558),
    .B(_0322_),
    .X(_0324_));
 sg13g2_nor2_1 _2089_ (.A(net558),
    .B(_0322_),
    .Y(_0325_));
 sg13g2_nor3_1 _2090_ (.A(net145),
    .B(_0324_),
    .C(net559),
    .Y(_0097_));
 sg13g2_and2_1 _2091_ (.A(net538),
    .B(_0324_),
    .X(_0326_));
 sg13g2_nor2_1 _2092_ (.A(net538),
    .B(_0324_),
    .Y(_0327_));
 sg13g2_nor3_1 _2093_ (.A(net145),
    .B(_0326_),
    .C(net539),
    .Y(_0098_));
 sg13g2_xnor2_1 _2094_ (.Y(_0328_),
    .A(net557),
    .B(_0326_));
 sg13g2_nor2_1 _2095_ (.A(net145),
    .B(_0328_),
    .Y(_0099_));
 sg13g2_nand3_1 _2096_ (.B(net557),
    .C(_0326_),
    .A(\tone_A_generator.counter[6] ),
    .Y(_0329_));
 sg13g2_a21o_1 _2097_ (.A2(_0326_),
    .A1(net557),
    .B1(net621),
    .X(_0330_));
 sg13g2_and4_1 _2098_ (.A(net180),
    .B(_0315_),
    .C(_0329_),
    .D(_0330_),
    .X(_0100_));
 sg13g2_nor2_2 _2099_ (.A(_0772_),
    .B(_0329_),
    .Y(_0331_));
 sg13g2_and2_1 _2100_ (.A(_0772_),
    .B(_0329_),
    .X(_0332_));
 sg13g2_nor3_1 _2101_ (.A(_0318_),
    .B(_0331_),
    .C(net612),
    .Y(_0101_));
 sg13g2_xnor2_1 _2102_ (.Y(_0333_),
    .A(net591),
    .B(_0331_));
 sg13g2_nor2_1 _2103_ (.A(net145),
    .B(net592),
    .Y(_0102_));
 sg13g2_and3_1 _2104_ (.X(_0334_),
    .A(net501),
    .B(net637),
    .C(_0331_));
 sg13g2_a21oi_1 _2105_ (.A1(\tone_A_generator.counter[8] ),
    .A2(_0331_),
    .Y(_0335_),
    .B1(net501));
 sg13g2_nor3_1 _2106_ (.A(net145),
    .B(_0334_),
    .C(net502),
    .Y(_0103_));
 sg13g2_xnor2_1 _2107_ (.Y(_0336_),
    .A(net548),
    .B(_0334_));
 sg13g2_nor2_1 _2108_ (.A(net145),
    .B(_0336_),
    .Y(_0104_));
 sg13g2_a21oi_1 _2109_ (.A1(\tone_A_generator.counter[10] ),
    .A2(_0334_),
    .Y(_0337_),
    .B1(net413));
 sg13g2_nor2_1 _2110_ (.A(net145),
    .B(net414),
    .Y(_0105_));
 sg13g2_nor2_1 _2111_ (.A(_0762_),
    .B(\register[3][3] ),
    .Y(_0338_));
 sg13g2_a22oi_1 _2112_ (.Y(_0339_),
    .B1(\register[3][2] ),
    .B2(_0763_),
    .A2(\register[3][3] ),
    .A1(_0762_));
 sg13g2_o21ai_1 _2113_ (.B1(net159),
    .Y(_0340_),
    .A1(_0338_),
    .A2(_0339_));
 sg13g2_a221oi_1 _2114_ (.B2(\tone_B_generator.counter[9] ),
    .C1(_0338_),
    .B1(_0799_),
    .A1(\tone_B_generator.counter[10] ),
    .Y(_0341_),
    .A2(_0798_));
 sg13g2_and2_1 _2115_ (.A(_0339_),
    .B(_0341_),
    .X(_0342_));
 sg13g2_nor2b_1 _2116_ (.A(\tone_B_generator.counter[9] ),
    .B_N(\register[3][1] ),
    .Y(_0343_));
 sg13g2_nor2_1 _2117_ (.A(\tone_B_generator.counter[8] ),
    .B(_0800_),
    .Y(_0344_));
 sg13g2_nand2b_1 _2118_ (.Y(_0345_),
    .B(\register[2][7] ),
    .A_N(\tone_B_generator.counter[7] ));
 sg13g2_o21ai_1 _2119_ (.B1(_0345_),
    .Y(_0346_),
    .A1(\tone_B_generator.counter[6] ),
    .A2(_0802_));
 sg13g2_a22oi_1 _2120_ (.Y(_0347_),
    .B1(_0801_),
    .B2(\tone_B_generator.counter[7] ),
    .A2(_0800_),
    .A1(\tone_B_generator.counter[8] ));
 sg13g2_a221oi_1 _2121_ (.B2(_0347_),
    .C1(_0343_),
    .B1(_0346_),
    .A1(_0764_),
    .Y(_0348_),
    .A2(\register[3][0] ));
 sg13g2_nor2b_1 _2122_ (.A(\tone_B_generator.counter[0] ),
    .B_N(\register[2][0] ),
    .Y(_0349_));
 sg13g2_or4_1 _2123_ (.A(_0343_),
    .B(_0344_),
    .C(_0346_),
    .D(_0349_),
    .X(_0350_));
 sg13g2_nand2b_1 _2124_ (.Y(_0351_),
    .B(\tone_B_generator.counter[0] ),
    .A_N(\register[2][0] ));
 sg13g2_a22oi_1 _2125_ (.Y(_0352_),
    .B1(_0350_),
    .B2(_0351_),
    .A2(\register[2][1] ),
    .A1(_0767_));
 sg13g2_nand2b_1 _2126_ (.Y(_0353_),
    .B(\tone_B_generator.counter[2] ),
    .A_N(\register[2][2] ));
 sg13g2_o21ai_1 _2127_ (.B1(_0353_),
    .Y(_0354_),
    .A1(_0767_),
    .A2(\register[2][1] ));
 sg13g2_a22oi_1 _2128_ (.Y(_0355_),
    .B1(\register[2][2] ),
    .B2(_0766_),
    .A2(\register[2][3] ),
    .A1(_0765_));
 sg13g2_o21ai_1 _2129_ (.B1(_0355_),
    .Y(_0356_),
    .A1(_0352_),
    .A2(_0354_));
 sg13g2_a22oi_1 _2130_ (.Y(_0357_),
    .B1(_0805_),
    .B2(\tone_B_generator.counter[3] ),
    .A2(_0804_),
    .A1(\tone_B_generator.counter[4] ));
 sg13g2_nand2b_1 _2131_ (.Y(_0358_),
    .B(\register[2][5] ),
    .A_N(\tone_B_generator.counter[5] ));
 sg13g2_o21ai_1 _2132_ (.B1(_0358_),
    .Y(_0359_),
    .A1(\tone_B_generator.counter[4] ),
    .A2(_0804_));
 sg13g2_a21oi_1 _2133_ (.A1(_0356_),
    .A2(_0357_),
    .Y(_0360_),
    .B1(_0359_));
 sg13g2_a22oi_1 _2134_ (.Y(_0361_),
    .B1(_0803_),
    .B2(\tone_B_generator.counter[5] ),
    .A2(_0802_),
    .A1(\tone_B_generator.counter[6] ));
 sg13g2_nand2_1 _2135_ (.Y(_0362_),
    .A(_0347_),
    .B(_0361_));
 sg13g2_o21ai_1 _2136_ (.B1(_0348_),
    .Y(_0363_),
    .A1(_0360_),
    .A2(_0362_));
 sg13g2_a21oi_2 _2137_ (.B1(_0340_),
    .Y(_0364_),
    .A2(_0363_),
    .A1(_0342_));
 sg13g2_a21oi_1 _2138_ (.A1(net343),
    .A2(_0364_),
    .Y(_0365_),
    .B1(net164));
 sg13g2_o21ai_1 _2139_ (.B1(_0365_),
    .Y(_0106_),
    .A1(_0768_),
    .A2(_0364_));
 sg13g2_nand2b_1 _2140_ (.Y(_0366_),
    .B(net181),
    .A_N(_0364_));
 sg13g2_xnor2_1 _2141_ (.Y(_0367_),
    .A(net597),
    .B(net159));
 sg13g2_nand2b_1 _2142_ (.Y(_0107_),
    .B(_0367_),
    .A_N(net146));
 sg13g2_and3_1 _2143_ (.X(_0368_),
    .A(net442),
    .B(\tone_B_generator.counter[0] ),
    .C(net159));
 sg13g2_a21oi_1 _2144_ (.A1(\tone_B_generator.counter[0] ),
    .A2(net159),
    .Y(_0369_),
    .B1(net442));
 sg13g2_nor3_1 _2145_ (.A(net146),
    .B(_0368_),
    .C(net443),
    .Y(_0108_));
 sg13g2_and2_1 _2146_ (.A(net518),
    .B(_0368_),
    .X(_0370_));
 sg13g2_nor2_1 _2147_ (.A(net518),
    .B(_0368_),
    .Y(_0371_));
 sg13g2_nor3_1 _2148_ (.A(net147),
    .B(_0370_),
    .C(net519),
    .Y(_0109_));
 sg13g2_and2_1 _2149_ (.A(net526),
    .B(_0370_),
    .X(_0372_));
 sg13g2_nor2_1 _2150_ (.A(net526),
    .B(_0370_),
    .Y(_0373_));
 sg13g2_nor3_1 _2151_ (.A(net147),
    .B(_0372_),
    .C(_0373_),
    .Y(_0110_));
 sg13g2_and2_1 _2152_ (.A(net511),
    .B(_0372_),
    .X(_0374_));
 sg13g2_nor2_1 _2153_ (.A(net511),
    .B(_0372_),
    .Y(_0375_));
 sg13g2_nor3_1 _2154_ (.A(net147),
    .B(_0374_),
    .C(net512),
    .Y(_0111_));
 sg13g2_and2_1 _2155_ (.A(net533),
    .B(_0374_),
    .X(_0376_));
 sg13g2_nor2_1 _2156_ (.A(net533),
    .B(_0374_),
    .Y(_0377_));
 sg13g2_nor3_1 _2157_ (.A(net147),
    .B(_0376_),
    .C(_0377_),
    .Y(_0112_));
 sg13g2_and2_1 _2158_ (.A(net509),
    .B(_0376_),
    .X(_0378_));
 sg13g2_nor2_1 _2159_ (.A(net509),
    .B(_0376_),
    .Y(_0379_));
 sg13g2_nor3_1 _2160_ (.A(net146),
    .B(_0378_),
    .C(net510),
    .Y(_0113_));
 sg13g2_and2_1 _2161_ (.A(net547),
    .B(_0378_),
    .X(_0380_));
 sg13g2_nor2_1 _2162_ (.A(net547),
    .B(_0378_),
    .Y(_0381_));
 sg13g2_nor3_1 _2163_ (.A(net146),
    .B(_0380_),
    .C(_0381_),
    .Y(_0114_));
 sg13g2_xnor2_1 _2164_ (.Y(_0382_),
    .A(net582),
    .B(_0380_));
 sg13g2_nor2_1 _2165_ (.A(net146),
    .B(_0382_),
    .Y(_0115_));
 sg13g2_and3_1 _2166_ (.X(_0383_),
    .A(net445),
    .B(net636),
    .C(_0380_));
 sg13g2_a21oi_1 _2167_ (.A1(\tone_B_generator.counter[8] ),
    .A2(_0380_),
    .Y(_0384_),
    .B1(net445));
 sg13g2_nor3_1 _2168_ (.A(net146),
    .B(_0383_),
    .C(net446),
    .Y(_0116_));
 sg13g2_xnor2_1 _2169_ (.Y(_0385_),
    .A(net570),
    .B(_0383_));
 sg13g2_nor2_1 _2170_ (.A(net146),
    .B(net571),
    .Y(_0117_));
 sg13g2_a21oi_1 _2171_ (.A1(\tone_B_generator.counter[10] ),
    .A2(_0383_),
    .Y(_0386_),
    .B1(net365));
 sg13g2_nor2_1 _2172_ (.A(net146),
    .B(net366),
    .Y(_0118_));
 sg13g2_and2_2 _2173_ (.A(_1087_),
    .B(_1098_),
    .X(_0387_));
 sg13g2_nor2_2 _2174_ (.A(net162),
    .B(_0387_),
    .Y(_0388_));
 sg13g2_a22oi_1 _2175_ (.Y(_0389_),
    .B1(_0388_),
    .B2(net339),
    .A2(_0387_),
    .A1(net176));
 sg13g2_inv_1 _2176_ (.Y(_0119_),
    .A(_0389_));
 sg13g2_a22oi_1 _2177_ (.Y(_0390_),
    .B1(_0388_),
    .B2(net348),
    .A2(_0387_),
    .A1(net174));
 sg13g2_inv_1 _2178_ (.Y(_0120_),
    .A(_0390_));
 sg13g2_a22oi_1 _2179_ (.Y(_0391_),
    .B1(_0388_),
    .B2(net342),
    .A2(_0387_),
    .A1(net172));
 sg13g2_inv_1 _2180_ (.Y(_0121_),
    .A(_0391_));
 sg13g2_a22oi_1 _2181_ (.Y(_0392_),
    .B1(_0388_),
    .B2(net341),
    .A2(_0387_),
    .A1(net170));
 sg13g2_inv_1 _2182_ (.Y(_0122_),
    .A(_0392_));
 sg13g2_a22oi_1 _2183_ (.Y(_0393_),
    .B1(_0388_),
    .B2(net161),
    .A2(_0387_),
    .A1(net168));
 sg13g2_inv_1 _2184_ (.Y(_0123_),
    .A(_0393_));
 sg13g2_a22oi_1 _2185_ (.Y(_0394_),
    .B1(\register[5][2] ),
    .B2(_0756_),
    .A2(\register[5][3] ),
    .A1(_0755_));
 sg13g2_a22oi_1 _2186_ (.Y(_0395_),
    .B1(_0797_),
    .B2(\tone_C_generator.counter[9] ),
    .A2(_0796_),
    .A1(\tone_C_generator.counter[10] ));
 sg13g2_nor2b_1 _2187_ (.A(\tone_C_generator.counter[8] ),
    .B_N(\register[5][0] ),
    .Y(_0396_));
 sg13g2_nand2_1 _2188_ (.Y(_0397_),
    .A(_0757_),
    .B(\register[5][1] ));
 sg13g2_nand2b_1 _2189_ (.Y(_0398_),
    .B(\tone_C_generator.counter[8] ),
    .A_N(\register[5][0] ));
 sg13g2_a22oi_1 _2190_ (.Y(_0399_),
    .B1(\register[4][6] ),
    .B2(_0759_),
    .A2(\register[4][7] ),
    .A1(_0758_));
 sg13g2_nor2_1 _2191_ (.A(_0758_),
    .B(\register[4][7] ),
    .Y(_0400_));
 sg13g2_nand2b_1 _2192_ (.Y(_0401_),
    .B(\tone_C_generator.counter[6] ),
    .A_N(\register[4][6] ));
 sg13g2_o21ai_1 _2193_ (.B1(_0401_),
    .Y(_0402_),
    .A1(_0760_),
    .A2(\register[4][5] ));
 sg13g2_nor2_1 _2194_ (.A(_0400_),
    .B(_0402_),
    .Y(_0403_));
 sg13g2_and2_1 _2195_ (.A(_0399_),
    .B(_0403_),
    .X(_0404_));
 sg13g2_a22oi_1 _2196_ (.Y(_0405_),
    .B1(\register[4][4] ),
    .B2(_0761_),
    .A2(\register[4][5] ),
    .A1(_0760_));
 sg13g2_nor2b_1 _2197_ (.A(\tone_C_generator.counter[2] ),
    .B_N(\register[4][2] ),
    .Y(_0406_));
 sg13g2_nor2b_1 _2198_ (.A(\tone_C_generator.counter[3] ),
    .B_N(\register[4][3] ),
    .Y(_0407_));
 sg13g2_nor2b_1 _2199_ (.A(\register[4][3] ),
    .B_N(\tone_C_generator.counter[3] ),
    .Y(_0408_));
 sg13g2_nand2b_1 _2200_ (.Y(_0409_),
    .B(\tone_C_generator.counter[3] ),
    .A_N(\register[4][3] ));
 sg13g2_o21ai_1 _2201_ (.B1(_0409_),
    .Y(_0410_),
    .A1(_0406_),
    .A2(_0407_));
 sg13g2_nor2b_1 _2202_ (.A(\register[4][2] ),
    .B_N(\tone_C_generator.counter[2] ),
    .Y(_0411_));
 sg13g2_nor4_2 _2203_ (.A(_0406_),
    .B(_0407_),
    .C(_0408_),
    .Y(_0412_),
    .D(_0411_));
 sg13g2_nor2_1 _2204_ (.A(\tone_C_generator.counter[1] ),
    .B(_0794_),
    .Y(_0413_));
 sg13g2_a22oi_1 _2205_ (.Y(_0414_),
    .B1(_0794_),
    .B2(\tone_C_generator.counter[1] ),
    .A2(_0793_),
    .A1(\tone_C_generator.counter[0] ));
 sg13g2_o21ai_1 _2206_ (.B1(_0412_),
    .Y(_0415_),
    .A1(_0413_),
    .A2(_0414_));
 sg13g2_a22oi_1 _2207_ (.Y(_0416_),
    .B1(_0410_),
    .B2(_0415_),
    .A2(_0795_),
    .A1(\tone_C_generator.counter[4] ));
 sg13g2_nand2b_1 _2208_ (.Y(_0417_),
    .B(_0405_),
    .A_N(_0416_));
 sg13g2_nor2_1 _2209_ (.A(_0399_),
    .B(_0400_),
    .Y(_0418_));
 sg13g2_a21o_1 _2210_ (.A2(_0417_),
    .A1(_0404_),
    .B1(_0418_),
    .X(_0419_));
 sg13g2_a221oi_1 _2211_ (.B2(_0419_),
    .C1(_0396_),
    .B1(_0398_),
    .A1(_0757_),
    .Y(_0420_),
    .A2(\register[5][1] ));
 sg13g2_nand2b_1 _2212_ (.Y(_0421_),
    .B(_0395_),
    .A_N(_0420_));
 sg13g2_and2_1 _2213_ (.A(_0394_),
    .B(_0421_),
    .X(_0422_));
 sg13g2_o21ai_1 _2214_ (.B1(_0398_),
    .Y(_0423_),
    .A1(_0761_),
    .A2(\register[4][4] ));
 sg13g2_nor2_1 _2215_ (.A(\tone_C_generator.counter[0] ),
    .B(_0793_),
    .Y(_0424_));
 sg13g2_nand3b_1 _2216_ (.B(_0397_),
    .C(_0394_),
    .Y(_0425_),
    .A_N(_0396_));
 sg13g2_nor4_1 _2217_ (.A(_0413_),
    .B(_0423_),
    .C(_0424_),
    .D(_0425_),
    .Y(_0426_));
 sg13g2_and4_1 _2218_ (.A(_0395_),
    .B(_0404_),
    .C(_0405_),
    .D(_0414_),
    .X(_0427_));
 sg13g2_nand3_1 _2219_ (.B(_0426_),
    .C(_0427_),
    .A(_0412_),
    .Y(_0428_));
 sg13g2_o21ai_1 _2220_ (.B1(_0428_),
    .Y(_0429_),
    .A1(_0755_),
    .A2(\register[5][3] ));
 sg13g2_o21ai_1 _2221_ (.B1(net158),
    .Y(_0430_),
    .A1(_0422_),
    .A2(_0429_));
 sg13g2_nor2b_1 _2222_ (.A(tone_C),
    .B_N(_0430_),
    .Y(_0431_));
 sg13g2_nor2_1 _2223_ (.A(net355),
    .B(_0430_),
    .Y(_0432_));
 sg13g2_o21ai_1 _2224_ (.B1(net180),
    .Y(_0124_),
    .A1(_0431_),
    .A2(_0432_));
 sg13g2_nand2_1 _2225_ (.Y(_0433_),
    .A(net180),
    .B(_0430_));
 sg13g2_xnor2_1 _2226_ (.Y(_0434_),
    .A(net600),
    .B(net158));
 sg13g2_nand3_1 _2227_ (.B(_0430_),
    .C(_0434_),
    .A(net180),
    .Y(_0125_));
 sg13g2_and3_1 _2228_ (.X(_0435_),
    .A(net482),
    .B(\tone_C_generator.counter[0] ),
    .C(net159));
 sg13g2_a21oi_1 _2229_ (.A1(\tone_C_generator.counter[0] ),
    .A2(net158),
    .Y(_0436_),
    .B1(net482));
 sg13g2_nor3_1 _2230_ (.A(_0433_),
    .B(_0435_),
    .C(net483),
    .Y(_0126_));
 sg13g2_and2_1 _2231_ (.A(net540),
    .B(_0435_),
    .X(_0437_));
 sg13g2_nor2_1 _2232_ (.A(net540),
    .B(_0435_),
    .Y(_0438_));
 sg13g2_nor3_1 _2233_ (.A(_0433_),
    .B(_0437_),
    .C(net541),
    .Y(_0127_));
 sg13g2_and2_1 _2234_ (.A(net579),
    .B(_0437_),
    .X(_0439_));
 sg13g2_nor2_1 _2235_ (.A(net579),
    .B(_0437_),
    .Y(_0440_));
 sg13g2_nor3_1 _2236_ (.A(net144),
    .B(_0439_),
    .C(_0440_),
    .Y(_0128_));
 sg13g2_and2_1 _2237_ (.A(net529),
    .B(_0439_),
    .X(_0441_));
 sg13g2_nor2_1 _2238_ (.A(net529),
    .B(_0439_),
    .Y(_0442_));
 sg13g2_nor3_1 _2239_ (.A(net144),
    .B(_0441_),
    .C(net530),
    .Y(_0129_));
 sg13g2_xnor2_1 _2240_ (.Y(_0443_),
    .A(net560),
    .B(_0441_));
 sg13g2_nor2_1 _2241_ (.A(net144),
    .B(_0443_),
    .Y(_0130_));
 sg13g2_nand3_1 _2242_ (.B(net560),
    .C(_0441_),
    .A(net601),
    .Y(_0444_));
 sg13g2_a21o_1 _2243_ (.A2(_0441_),
    .A1(net560),
    .B1(net601),
    .X(_0445_));
 sg13g2_and4_1 _2244_ (.A(net180),
    .B(_0430_),
    .C(_0444_),
    .D(_0445_),
    .X(_0131_));
 sg13g2_nor2_1 _2245_ (.A(_0758_),
    .B(_0444_),
    .Y(_0446_));
 sg13g2_and2_1 _2246_ (.A(_0758_),
    .B(_0444_),
    .X(_0447_));
 sg13g2_nor3_1 _2247_ (.A(net144),
    .B(_0446_),
    .C(_0447_),
    .Y(_0132_));
 sg13g2_and2_1 _2248_ (.A(net561),
    .B(_0446_),
    .X(_0448_));
 sg13g2_nor2_1 _2249_ (.A(net561),
    .B(_0446_),
    .Y(_0449_));
 sg13g2_nor3_1 _2250_ (.A(net144),
    .B(_0448_),
    .C(net562),
    .Y(_0133_));
 sg13g2_and2_1 _2251_ (.A(net536),
    .B(_0448_),
    .X(_0450_));
 sg13g2_nor2_1 _2252_ (.A(net536),
    .B(_0448_),
    .Y(_0451_));
 sg13g2_nor3_1 _2253_ (.A(net144),
    .B(_0450_),
    .C(net537),
    .Y(_0134_));
 sg13g2_xnor2_1 _2254_ (.Y(_0452_),
    .A(net574),
    .B(_0450_));
 sg13g2_nor2_1 _2255_ (.A(net144),
    .B(_0452_),
    .Y(_0135_));
 sg13g2_a21oi_1 _2256_ (.A1(\tone_C_generator.counter[10] ),
    .A2(_0450_),
    .Y(_0453_),
    .B1(net362));
 sg13g2_nor2_1 _2257_ (.A(net144),
    .B(net363),
    .Y(_0136_));
 sg13g2_and2_2 _2258_ (.A(_1009_),
    .B(_0269_),
    .X(_0454_));
 sg13g2_nor2_2 _2259_ (.A(net162),
    .B(_0454_),
    .Y(_0455_));
 sg13g2_a22oi_1 _2260_ (.Y(_0456_),
    .B1(_0455_),
    .B2(net357),
    .A2(_0454_),
    .A1(net176));
 sg13g2_inv_1 _2261_ (.Y(_0137_),
    .A(_0456_));
 sg13g2_a22oi_1 _2262_ (.Y(_0457_),
    .B1(_0455_),
    .B2(net396),
    .A2(_0454_),
    .A1(net174));
 sg13g2_inv_1 _2263_ (.Y(_0138_),
    .A(_0457_));
 sg13g2_a22oi_1 _2264_ (.Y(_0458_),
    .B1(_0455_),
    .B2(net372),
    .A2(_0454_),
    .A1(net172));
 sg13g2_inv_1 _2265_ (.Y(_0139_),
    .A(_0458_));
 sg13g2_a22oi_1 _2266_ (.Y(_0459_),
    .B1(_0455_),
    .B2(net353),
    .A2(_0454_),
    .A1(net170));
 sg13g2_inv_1 _2267_ (.Y(_0140_),
    .A(_0459_));
 sg13g2_a22oi_1 _2268_ (.Y(_0460_),
    .B1(_0455_),
    .B2(net349),
    .A2(_0454_),
    .A1(net168));
 sg13g2_inv_1 _2269_ (.Y(_0141_),
    .A(_0460_));
 sg13g2_a22oi_1 _2270_ (.Y(_0461_),
    .B1(_0455_),
    .B2(net391),
    .A2(_0454_),
    .A1(net2));
 sg13g2_inv_1 _2271_ (.Y(_0142_),
    .A(_0461_));
 sg13g2_and2_2 _2272_ (.A(_0990_),
    .B(_1098_),
    .X(_0462_));
 sg13g2_nor2_2 _2273_ (.A(net164),
    .B(_0462_),
    .Y(_0463_));
 sg13g2_a22oi_1 _2274_ (.Y(_0464_),
    .B1(_0463_),
    .B2(net338),
    .A2(_0462_),
    .A1(net175));
 sg13g2_inv_1 _2275_ (.Y(_0143_),
    .A(_0464_));
 sg13g2_a22oi_1 _2276_ (.Y(_0465_),
    .B1(_0463_),
    .B2(net347),
    .A2(_0462_),
    .A1(net173));
 sg13g2_inv_1 _2277_ (.Y(_0144_),
    .A(_0465_));
 sg13g2_a22oi_1 _2278_ (.Y(_0466_),
    .B1(_0463_),
    .B2(net350),
    .A2(_0462_),
    .A1(net171));
 sg13g2_inv_1 _2279_ (.Y(_0145_),
    .A(_0466_));
 sg13g2_a22oi_1 _2280_ (.Y(_0467_),
    .B1(_0463_),
    .B2(net340),
    .A2(_0462_),
    .A1(net169));
 sg13g2_inv_1 _2281_ (.Y(_0146_),
    .A(_0467_));
 sg13g2_a22oi_1 _2282_ (.Y(_0468_),
    .B1(_0463_),
    .B2(net581),
    .A2(_0462_),
    .A1(net168));
 sg13g2_inv_1 _2283_ (.Y(_0147_),
    .A(_0468_));
 sg13g2_nor2_2 _2284_ (.A(net563),
    .B(net166),
    .Y(_0469_));
 sg13g2_nand2b_2 _2285_ (.Y(_0470_),
    .B(net185),
    .A_N(restart_envelope));
 sg13g2_nor2_1 _2286_ (.A(_0724_),
    .B(_0470_),
    .Y(_0148_));
 sg13g2_xnor2_1 _2287_ (.Y(_0471_),
    .A(net578),
    .B(net158));
 sg13g2_nand2b_1 _2288_ (.Y(_0472_),
    .B(\noise_generator.period[2] ),
    .A_N(\noise_generator.tone.counter[2] ));
 sg13g2_a22oi_1 _2289_ (.Y(_0473_),
    .B1(\noise_generator.period[1] ),
    .B2(_0753_),
    .A2(\noise_generator.period[0] ),
    .A1(_0754_));
 sg13g2_nand2b_1 _2290_ (.Y(_0474_),
    .B(\noise_generator.tone.counter[2] ),
    .A_N(\noise_generator.period[2] ));
 sg13g2_o21ai_1 _2291_ (.B1(_0474_),
    .Y(_0475_),
    .A1(_0753_),
    .A2(\noise_generator.period[1] ));
 sg13g2_o21ai_1 _2292_ (.B1(_0472_),
    .Y(_0476_),
    .A1(_0473_),
    .A2(_0475_));
 sg13g2_o21ai_1 _2293_ (.B1(_0476_),
    .Y(_0477_),
    .A1(_0752_),
    .A2(\noise_generator.period[3] ));
 sg13g2_a22oi_1 _2294_ (.Y(_0478_),
    .B1(\noise_generator.period[4] ),
    .B2(_0751_),
    .A2(\noise_generator.period[3] ),
    .A1(_0752_));
 sg13g2_a22oi_1 _2295_ (.Y(_0479_),
    .B1(_0477_),
    .B2(_0478_),
    .A2(_0784_),
    .A1(\noise_generator.tone.counter[4] ));
 sg13g2_nor2_1 _2296_ (.A(_0285_),
    .B(_0479_),
    .Y(_0480_));
 sg13g2_o21ai_1 _2297_ (.B1(net179),
    .Y(_0481_),
    .A1(_0285_),
    .A2(_0479_));
 sg13g2_nand2b_1 _2298_ (.Y(_0149_),
    .B(_0471_),
    .A_N(_0481_));
 sg13g2_nor3_2 _2299_ (.A(_0753_),
    .B(_0754_),
    .C(_0285_),
    .Y(_0482_));
 sg13g2_a21oi_1 _2300_ (.A1(\noise_generator.tone.counter[0] ),
    .A2(net158),
    .Y(_0483_),
    .B1(net375));
 sg13g2_nor3_1 _2301_ (.A(_0481_),
    .B(_0482_),
    .C(net376),
    .Y(_0150_));
 sg13g2_and2_1 _2302_ (.A(net504),
    .B(_0482_),
    .X(_0484_));
 sg13g2_nor2_1 _2303_ (.A(net504),
    .B(_0482_),
    .Y(_0485_));
 sg13g2_nor3_1 _2304_ (.A(_0481_),
    .B(_0484_),
    .C(net505),
    .Y(_0151_));
 sg13g2_xnor2_1 _2305_ (.Y(_0486_),
    .A(net516),
    .B(_0484_));
 sg13g2_nor2_1 _2306_ (.A(_0481_),
    .B(_0486_),
    .Y(_0152_));
 sg13g2_a21oi_1 _2307_ (.A1(\noise_generator.tone.counter[3] ),
    .A2(_0484_),
    .Y(_0487_),
    .B1(net405));
 sg13g2_nor2_1 _2308_ (.A(_0481_),
    .B(net406),
    .Y(_0153_));
 sg13g2_a21oi_1 _2309_ (.A1(net373),
    .A2(_0480_),
    .Y(_0488_),
    .B1(net163));
 sg13g2_o21ai_1 _2310_ (.B1(_0488_),
    .Y(_0154_),
    .A1(_0750_),
    .A2(_0480_));
 sg13g2_nor2_1 _2311_ (.A(_0750_),
    .B(\noise_generator.signal_edge.previous_signal_state_0 ),
    .Y(_0489_));
 sg13g2_nand2b_2 _2312_ (.Y(_0490_),
    .B(net472),
    .A_N(net531));
 sg13g2_o21ai_1 _2313_ (.B1(net179),
    .Y(_0491_),
    .A1(\noise_generator.lfsr[0] ),
    .A2(net157));
 sg13g2_a21oi_1 _2314_ (.A1(_0749_),
    .A2(net157),
    .Y(_0155_),
    .B1(_0491_));
 sg13g2_o21ai_1 _2315_ (.B1(net179),
    .Y(_0492_),
    .A1(net434),
    .A2(net156));
 sg13g2_a21oi_1 _2316_ (.A1(_0748_),
    .A2(net156),
    .Y(_0156_),
    .B1(_0492_));
 sg13g2_o21ai_1 _2317_ (.B1(net177),
    .Y(_0493_),
    .A1(net498),
    .A2(_0490_));
 sg13g2_a21oi_1 _2318_ (.A1(_0748_),
    .A2(_0490_),
    .Y(_0157_),
    .B1(net499));
 sg13g2_o21ai_1 _2319_ (.B1(net177),
    .Y(_0494_),
    .A1(\noise_generator.lfsr[3] ),
    .A2(net156));
 sg13g2_a21oi_1 _2320_ (.A1(_0747_),
    .A2(net156),
    .Y(_0158_),
    .B1(_0494_));
 sg13g2_o21ai_1 _2321_ (.B1(net177),
    .Y(_0495_),
    .A1(net462),
    .A2(net156));
 sg13g2_a21oi_1 _2322_ (.A1(_0746_),
    .A2(net156),
    .Y(_0159_),
    .B1(_0495_));
 sg13g2_o21ai_1 _2323_ (.B1(net177),
    .Y(_0496_),
    .A1(\noise_generator.lfsr[5] ),
    .A2(net156));
 sg13g2_a21oi_1 _2324_ (.A1(_0745_),
    .A2(net156),
    .Y(_0160_),
    .B1(_0496_));
 sg13g2_o21ai_1 _2325_ (.B1(net177),
    .Y(_0497_),
    .A1(\noise_generator.lfsr[6] ),
    .A2(net157));
 sg13g2_a21oi_1 _2326_ (.A1(_0744_),
    .A2(net157),
    .Y(_0161_),
    .B1(_0497_));
 sg13g2_o21ai_1 _2327_ (.B1(net177),
    .Y(_0498_),
    .A1(\noise_generator.lfsr[7] ),
    .A2(net157));
 sg13g2_a21oi_1 _2328_ (.A1(_0743_),
    .A2(net157),
    .Y(_0162_),
    .B1(_0498_));
 sg13g2_o21ai_1 _2329_ (.B1(net177),
    .Y(_0499_),
    .A1(\noise_generator.lfsr[8] ),
    .A2(net155));
 sg13g2_a21oi_1 _2330_ (.A1(_0742_),
    .A2(net155),
    .Y(_0163_),
    .B1(_0499_));
 sg13g2_o21ai_1 _2331_ (.B1(net178),
    .Y(_0500_),
    .A1(net416),
    .A2(net153));
 sg13g2_a21oi_1 _2332_ (.A1(_0741_),
    .A2(net153),
    .Y(_0164_),
    .B1(_0500_));
 sg13g2_o21ai_1 _2333_ (.B1(net178),
    .Y(_0501_),
    .A1(\noise_generator.lfsr[10] ),
    .A2(net153));
 sg13g2_a21oi_1 _2334_ (.A1(_0740_),
    .A2(net153),
    .Y(_0165_),
    .B1(_0501_));
 sg13g2_o21ai_1 _2335_ (.B1(net178),
    .Y(_0502_),
    .A1(net449),
    .A2(net153));
 sg13g2_a21oi_1 _2336_ (.A1(_0739_),
    .A2(net153),
    .Y(_0166_),
    .B1(_0502_));
 sg13g2_o21ai_1 _2337_ (.B1(net178),
    .Y(_0503_),
    .A1(\noise_generator.lfsr[12] ),
    .A2(net154));
 sg13g2_a21oi_1 _2338_ (.A1(_0738_),
    .A2(net154),
    .Y(_0167_),
    .B1(_0503_));
 sg13g2_o21ai_1 _2339_ (.B1(net178),
    .Y(_0504_),
    .A1(net453),
    .A2(net154));
 sg13g2_a21oi_1 _2340_ (.A1(_0737_),
    .A2(net154),
    .Y(_0168_),
    .B1(_0504_));
 sg13g2_o21ai_1 _2341_ (.B1(net178),
    .Y(_0505_),
    .A1(\noise_generator.lfsr[14] ),
    .A2(net153));
 sg13g2_a21oi_1 _2342_ (.A1(_0736_),
    .A2(net153),
    .Y(_0169_),
    .B1(_0505_));
 sg13g2_o21ai_1 _2343_ (.B1(net178),
    .Y(_0506_),
    .A1(net432),
    .A2(net155));
 sg13g2_a21oi_1 _2344_ (.A1(_0735_),
    .A2(net155),
    .Y(_0170_),
    .B1(_0506_));
 sg13g2_nor4_1 _2345_ (.A(net465),
    .B(net449),
    .C(net480),
    .D(net416),
    .Y(_0507_));
 sg13g2_nor4_1 _2346_ (.A(net469),
    .B(net432),
    .C(net495),
    .D(net453),
    .Y(_0508_));
 sg13g2_nand4_1 _2347_ (.B(_0744_),
    .C(_0745_),
    .A(_0743_),
    .Y(_0509_),
    .D(_0746_));
 sg13g2_nor4_1 _2348_ (.A(net462),
    .B(net471),
    .C(net434),
    .D(_0509_),
    .Y(_0510_));
 sg13g2_nand3_1 _2349_ (.B(_0508_),
    .C(_0510_),
    .A(_0507_),
    .Y(_0511_));
 sg13g2_nor3_1 _2350_ (.A(net498),
    .B(\noise_generator.lfsr[0] ),
    .C(_0490_),
    .Y(_0512_));
 sg13g2_nand2_1 _2351_ (.Y(_0513_),
    .A(net498),
    .B(\noise_generator.lfsr[0] ));
 sg13g2_o21ai_1 _2352_ (.B1(net177),
    .Y(_0514_),
    .A1(_0490_),
    .A2(_0513_));
 sg13g2_a221oi_1 _2353_ (.B2(_0512_),
    .C1(_0514_),
    .B1(_0511_),
    .A1(_0735_),
    .Y(_0171_),
    .A2(_0490_));
 sg13g2_and2_1 _2354_ (.A(_1009_),
    .B(_1087_),
    .X(_0515_));
 sg13g2_nor2_2 _2355_ (.A(net162),
    .B(net149),
    .Y(_0516_));
 sg13g2_a22oi_1 _2356_ (.Y(_0517_),
    .B1(_0516_),
    .B2(net408),
    .A2(net149),
    .A1(net175));
 sg13g2_inv_1 _2357_ (.Y(_0172_),
    .A(_0517_));
 sg13g2_a22oi_1 _2358_ (.Y(_0518_),
    .B1(_0516_),
    .B2(net390),
    .A2(net149),
    .A1(net173));
 sg13g2_inv_1 _2359_ (.Y(_0173_),
    .A(_0518_));
 sg13g2_a22oi_1 _2360_ (.Y(_0519_),
    .B1(_0516_),
    .B2(net427),
    .A2(_0515_),
    .A1(net171));
 sg13g2_inv_1 _2361_ (.Y(_0174_),
    .A(_0519_));
 sg13g2_a22oi_1 _2362_ (.Y(_0520_),
    .B1(_0516_),
    .B2(net436),
    .A2(net149),
    .A1(net169));
 sg13g2_inv_1 _2363_ (.Y(_0175_),
    .A(_0520_));
 sg13g2_a22oi_1 _2364_ (.Y(_0521_),
    .B1(_0516_),
    .B2(net522),
    .A2(net149),
    .A1(net168));
 sg13g2_inv_1 _2365_ (.Y(_0176_),
    .A(_0521_));
 sg13g2_a22oi_1 _2366_ (.Y(_0522_),
    .B1(_0516_),
    .B2(net507),
    .A2(net149),
    .A1(net2));
 sg13g2_inv_1 _2367_ (.Y(_0177_),
    .A(_0522_));
 sg13g2_a22oi_1 _2368_ (.Y(_0523_),
    .B1(_0516_),
    .B2(net475),
    .A2(net149),
    .A1(net3));
 sg13g2_inv_1 _2369_ (.Y(_0178_),
    .A(_0523_));
 sg13g2_a22oi_1 _2370_ (.Y(_0524_),
    .B1(_0516_),
    .B2(net520),
    .A2(net149),
    .A1(net4));
 sg13g2_inv_1 _2371_ (.Y(_0179_),
    .A(_0524_));
 sg13g2_xnor2_1 _2372_ (.Y(_0525_),
    .A(\envelope_generator.hold ),
    .B(envelope_alternate));
 sg13g2_nand2_1 _2373_ (.Y(_0526_),
    .A(envelope_continue),
    .B(_0525_));
 sg13g2_nand2b_1 _2374_ (.Y(_0527_),
    .B(net387),
    .A_N(\envelope_generator.signal_edge.previous_signal_state_0 ));
 sg13g2_and3_1 _2375_ (.X(_0528_),
    .A(\envelope_generator.envelope_counter[2] ),
    .B(\envelope_generator.envelope_counter[1] ),
    .C(\envelope_generator.envelope_counter[0] ));
 sg13g2_nand2_1 _2376_ (.Y(_0529_),
    .A(\envelope_generator.envelope_counter[3] ),
    .B(_0528_));
 sg13g2_nor2_1 _2377_ (.A(_0527_),
    .B(_0529_),
    .Y(_0530_));
 sg13g2_inv_1 _2378_ (.Y(_0531_),
    .A(_0530_));
 sg13g2_nand2b_1 _2379_ (.Y(_0532_),
    .B(envelope_attack),
    .A_N(envelope_continue));
 sg13g2_nand3_1 _2380_ (.B(_0530_),
    .C(_0532_),
    .A(_0526_),
    .Y(_0533_));
 sg13g2_nor2_1 _2381_ (.A(\envelope_generator.invert_output ),
    .B(_0470_),
    .Y(_0534_));
 sg13g2_nor3_1 _2382_ (.A(_0009_),
    .B(_0470_),
    .C(_0533_),
    .Y(_0535_));
 sg13g2_a221oi_1 _2383_ (.B2(_0534_),
    .C1(_0535_),
    .B1(_0533_),
    .A1(_0817_),
    .Y(_0180_),
    .A2(_0470_));
 sg13g2_a22oi_1 _2384_ (.Y(_0536_),
    .B1(\envelope_generator.period[0] ),
    .B2(_0734_),
    .A2(\envelope_generator.period[1] ),
    .A1(_0733_));
 sg13g2_nand2b_1 _2385_ (.Y(_0537_),
    .B(\envelope_generator.tone.counter[2] ),
    .A_N(\envelope_generator.period[2] ));
 sg13g2_o21ai_1 _2386_ (.B1(_0537_),
    .Y(_0538_),
    .A1(_0733_),
    .A2(\envelope_generator.period[1] ));
 sg13g2_a22oi_1 _2387_ (.Y(_0539_),
    .B1(\envelope_generator.period[2] ),
    .B2(_0732_),
    .A2(\envelope_generator.period[3] ),
    .A1(_0731_));
 sg13g2_o21ai_1 _2388_ (.B1(_0539_),
    .Y(_0540_),
    .A1(_0536_),
    .A2(_0538_));
 sg13g2_a22oi_1 _2389_ (.Y(_0541_),
    .B1(_0792_),
    .B2(\envelope_generator.tone.counter[3] ),
    .A2(_0791_),
    .A1(\envelope_generator.tone.counter[4] ));
 sg13g2_a22oi_1 _2390_ (.Y(_0542_),
    .B1(_0540_),
    .B2(_0541_),
    .A2(\envelope_generator.period[4] ),
    .A1(_0730_));
 sg13g2_a21oi_1 _2391_ (.A1(\envelope_generator.tone.counter[5] ),
    .A2(_0790_),
    .Y(_0543_),
    .B1(_0542_));
 sg13g2_nand2b_1 _2392_ (.Y(_0544_),
    .B(\envelope_generator.period[6] ),
    .A_N(\envelope_generator.tone.counter[6] ));
 sg13g2_o21ai_1 _2393_ (.B1(_0544_),
    .Y(_0545_),
    .A1(\envelope_generator.tone.counter[5] ),
    .A2(_0790_));
 sg13g2_a22oi_1 _2394_ (.Y(_0546_),
    .B1(_0789_),
    .B2(\envelope_generator.tone.counter[6] ),
    .A2(_0788_),
    .A1(\envelope_generator.tone.counter[7] ));
 sg13g2_o21ai_1 _2395_ (.B1(_0546_),
    .Y(_0547_),
    .A1(_0543_),
    .A2(_0545_));
 sg13g2_nor2_1 _2396_ (.A(\envelope_generator.tone.counter[9] ),
    .B(_0787_),
    .Y(_0548_));
 sg13g2_a221oi_1 _2397_ (.B2(_0729_),
    .C1(_0548_),
    .B1(\envelope_generator.period[7] ),
    .A1(_0728_),
    .Y(_0549_),
    .A2(\envelope_generator.period[8] ));
 sg13g2_nor2_1 _2398_ (.A(_0728_),
    .B(\envelope_generator.period[8] ),
    .Y(_0550_));
 sg13g2_a221oi_1 _2399_ (.B2(_0549_),
    .C1(_0550_),
    .B1(_0547_),
    .A1(\envelope_generator.tone.counter[9] ),
    .Y(_0551_),
    .A2(_0787_));
 sg13g2_a22oi_1 _2400_ (.Y(_0552_),
    .B1(_0548_),
    .B2(_0550_),
    .A2(\envelope_generator.period[10] ),
    .A1(_0727_));
 sg13g2_o21ai_1 _2401_ (.B1(_0552_),
    .Y(_0553_),
    .A1(\envelope_generator.tone.counter[11] ),
    .A2(_0785_));
 sg13g2_a22oi_1 _2402_ (.Y(_0554_),
    .B1(_0786_),
    .B2(\envelope_generator.tone.counter[10] ),
    .A2(_0785_),
    .A1(\envelope_generator.tone.counter[11] ));
 sg13g2_o21ai_1 _2403_ (.B1(_0554_),
    .Y(_0555_),
    .A1(_0551_),
    .A2(_0553_));
 sg13g2_nand2b_1 _2404_ (.Y(_0556_),
    .B(\envelope_generator.tone.counter[12] ),
    .A_N(\envelope_generator.period[12] ));
 sg13g2_o21ai_1 _2405_ (.B1(_0556_),
    .Y(_0557_),
    .A1(_0726_),
    .A2(\envelope_generator.period[13] ));
 sg13g2_nand2_1 _2406_ (.Y(_0558_),
    .A(_0725_),
    .B(\envelope_generator.period[15] ));
 sg13g2_nor2b_1 _2407_ (.A(\envelope_generator.tone.counter[12] ),
    .B_N(\envelope_generator.period[12] ),
    .Y(_0559_));
 sg13g2_nand2b_1 _2408_ (.Y(_0560_),
    .B(\envelope_generator.tone.counter[14] ),
    .A_N(\envelope_generator.period[14] ));
 sg13g2_o21ai_1 _2409_ (.B1(_0560_),
    .Y(_0561_),
    .A1(_0725_),
    .A2(\envelope_generator.period[15] ));
 sg13g2_nor4_1 _2410_ (.A(\envelope_generator.tone.counter[11] ),
    .B(_0727_),
    .C(_0785_),
    .D(\envelope_generator.period[10] ),
    .Y(_0562_));
 sg13g2_nand2_1 _2411_ (.Y(_0563_),
    .A(_0726_),
    .B(\envelope_generator.period[13] ));
 sg13g2_nand2b_1 _2412_ (.Y(_0564_),
    .B(\envelope_generator.period[14] ),
    .A_N(\envelope_generator.tone.counter[14] ));
 sg13g2_nand3_1 _2413_ (.B(_0563_),
    .C(_0564_),
    .A(_0558_),
    .Y(_0565_));
 sg13g2_nor2_1 _2414_ (.A(_0561_),
    .B(_0565_),
    .Y(_0566_));
 sg13g2_nor3_1 _2415_ (.A(_0557_),
    .B(_0559_),
    .C(_0562_),
    .Y(_0567_));
 sg13g2_nand3_1 _2416_ (.B(_0566_),
    .C(_0567_),
    .A(_0555_),
    .Y(_0568_));
 sg13g2_a22oi_1 _2417_ (.Y(_0569_),
    .B1(_0566_),
    .B2(_0557_),
    .A2(_0561_),
    .A1(_0558_));
 sg13g2_a21oi_2 _2418_ (.B1(_0285_),
    .Y(_0570_),
    .A2(_0569_),
    .A1(_0568_));
 sg13g2_nand2b_1 _2419_ (.Y(_0571_),
    .B(_0469_),
    .A_N(_0570_));
 sg13g2_xnor2_1 _2420_ (.Y(_0572_),
    .A(net590),
    .B(_0284_));
 sg13g2_nand2b_1 _2421_ (.Y(_0181_),
    .B(_0572_),
    .A_N(net142));
 sg13g2_a21oi_1 _2422_ (.A1(\envelope_generator.tone.counter[0] ),
    .A2(net159),
    .Y(_0573_),
    .B1(net429));
 sg13g2_nor3_1 _2423_ (.A(_0733_),
    .B(_0734_),
    .C(_0285_),
    .Y(_0574_));
 sg13g2_nor3_1 _2424_ (.A(net142),
    .B(net430),
    .C(_0574_),
    .Y(_0182_));
 sg13g2_nand4_1 _2425_ (.B(net429),
    .C(net590),
    .A(net553),
    .Y(_0575_),
    .D(net159));
 sg13g2_xnor2_1 _2426_ (.Y(_0576_),
    .A(net553),
    .B(_0574_));
 sg13g2_nor2_1 _2427_ (.A(net142),
    .B(net554),
    .Y(_0183_));
 sg13g2_and2_1 _2428_ (.A(_0731_),
    .B(_0575_),
    .X(_0577_));
 sg13g2_nor2_1 _2429_ (.A(_0731_),
    .B(_0575_),
    .Y(_0578_));
 sg13g2_nor3_1 _2430_ (.A(net142),
    .B(_0577_),
    .C(_0578_),
    .Y(_0184_));
 sg13g2_nor2_1 _2431_ (.A(net544),
    .B(_0578_),
    .Y(_0579_));
 sg13g2_nor3_2 _2432_ (.A(_0730_),
    .B(_0731_),
    .C(_0575_),
    .Y(_0580_));
 sg13g2_nor3_1 _2433_ (.A(net142),
    .B(net545),
    .C(_0580_),
    .Y(_0185_));
 sg13g2_xnor2_1 _2434_ (.Y(_0581_),
    .A(net575),
    .B(_0580_));
 sg13g2_nor2_1 _2435_ (.A(net142),
    .B(net576),
    .Y(_0186_));
 sg13g2_and3_1 _2436_ (.X(_0582_),
    .A(net491),
    .B(\envelope_generator.tone.counter[5] ),
    .C(_0580_));
 sg13g2_a21oi_1 _2437_ (.A1(\envelope_generator.tone.counter[5] ),
    .A2(_0580_),
    .Y(_0583_),
    .B1(net491));
 sg13g2_nor3_1 _2438_ (.A(net142),
    .B(_0582_),
    .C(net492),
    .Y(_0187_));
 sg13g2_and2_1 _2439_ (.A(net542),
    .B(_0582_),
    .X(_0584_));
 sg13g2_nor2_1 _2440_ (.A(net542),
    .B(_0582_),
    .Y(_0585_));
 sg13g2_nor3_1 _2441_ (.A(net142),
    .B(_0584_),
    .C(net543),
    .Y(_0188_));
 sg13g2_nor2_1 _2442_ (.A(net534),
    .B(_0584_),
    .Y(_0586_));
 sg13g2_and2_1 _2443_ (.A(net534),
    .B(_0584_),
    .X(_0587_));
 sg13g2_nor3_1 _2444_ (.A(net143),
    .B(net535),
    .C(_0587_),
    .Y(_0189_));
 sg13g2_xnor2_1 _2445_ (.Y(_0588_),
    .A(net580),
    .B(_0587_));
 sg13g2_nor2_1 _2446_ (.A(net143),
    .B(_0588_),
    .Y(_0190_));
 sg13g2_a21oi_1 _2447_ (.A1(\envelope_generator.tone.counter[9] ),
    .A2(_0587_),
    .Y(_0589_),
    .B1(net523));
 sg13g2_and3_1 _2448_ (.X(_0590_),
    .A(net523),
    .B(\envelope_generator.tone.counter[9] ),
    .C(_0587_));
 sg13g2_nor3_1 _2449_ (.A(net143),
    .B(net524),
    .C(_0590_),
    .Y(_0191_));
 sg13g2_nor2_1 _2450_ (.A(net555),
    .B(_0590_),
    .Y(_0591_));
 sg13g2_and2_1 _2451_ (.A(net555),
    .B(_0590_),
    .X(_0592_));
 sg13g2_nor3_1 _2452_ (.A(net143),
    .B(net556),
    .C(_0592_),
    .Y(_0192_));
 sg13g2_xnor2_1 _2453_ (.Y(_0593_),
    .A(net577),
    .B(_0592_));
 sg13g2_nor2_1 _2454_ (.A(net143),
    .B(_0593_),
    .Y(_0193_));
 sg13g2_and3_1 _2455_ (.X(_0594_),
    .A(net397),
    .B(\envelope_generator.tone.counter[12] ),
    .C(_0592_));
 sg13g2_a21oi_1 _2456_ (.A1(\envelope_generator.tone.counter[12] ),
    .A2(_0592_),
    .Y(_0595_),
    .B1(net397));
 sg13g2_nor3_1 _2457_ (.A(net143),
    .B(_0594_),
    .C(net398),
    .Y(_0194_));
 sg13g2_xnor2_1 _2458_ (.Y(_0596_),
    .A(net551),
    .B(_0594_));
 sg13g2_nor2_1 _2459_ (.A(net143),
    .B(net552),
    .Y(_0195_));
 sg13g2_a21oi_1 _2460_ (.A1(\envelope_generator.tone.counter[14] ),
    .A2(_0594_),
    .Y(_0597_),
    .B1(net359));
 sg13g2_nor2_1 _2461_ (.A(net143),
    .B(net360),
    .Y(_0196_));
 sg13g2_a21oi_1 _2462_ (.A1(net367),
    .A2(_0570_),
    .Y(_0598_),
    .B1(_0470_));
 sg13g2_o21ai_1 _2463_ (.B1(net368),
    .Y(_0197_),
    .A1(_0724_),
    .A2(_0570_));
 sg13g2_nand2b_1 _2464_ (.Y(_0599_),
    .B(net476),
    .A_N(\envelope_generator.hold ));
 sg13g2_o21ai_1 _2465_ (.B1(net485),
    .Y(_0600_),
    .A1(_0527_),
    .A2(_0599_));
 sg13g2_a21oi_1 _2466_ (.A1(_0531_),
    .A2(net486),
    .Y(_0198_),
    .B1(_0470_));
 sg13g2_a21oi_2 _2467_ (.B1(_0527_),
    .Y(_0601_),
    .A2(_0599_),
    .A1(net485));
 sg13g2_o21ai_1 _2468_ (.B1(_0469_),
    .Y(_0602_),
    .A1(\envelope_generator.envelope_counter[0] ),
    .A2(_0601_));
 sg13g2_a21oi_1 _2469_ (.A1(_0723_),
    .A2(_0601_),
    .Y(_0199_),
    .B1(_0602_));
 sg13g2_a21oi_1 _2470_ (.A1(\envelope_generator.envelope_counter[0] ),
    .A2(_0601_),
    .Y(_0603_),
    .B1(net513));
 sg13g2_and3_1 _2471_ (.X(_0604_),
    .A(net513),
    .B(\envelope_generator.envelope_counter[0] ),
    .C(_0601_));
 sg13g2_nor3_1 _2472_ (.A(_0470_),
    .B(net514),
    .C(_0604_),
    .Y(_0200_));
 sg13g2_and2_1 _2473_ (.A(_0528_),
    .B(_0601_),
    .X(_0605_));
 sg13g2_o21ai_1 _2474_ (.B1(_0469_),
    .Y(_0606_),
    .A1(\envelope_generator.envelope_counter[2] ),
    .A2(_0604_));
 sg13g2_nor2_1 _2475_ (.A(_0605_),
    .B(net564),
    .Y(_0201_));
 sg13g2_o21ai_1 _2476_ (.B1(_0469_),
    .Y(_0607_),
    .A1(net496),
    .A2(_0605_));
 sg13g2_a21oi_1 _2477_ (.A1(net496),
    .A2(_0605_),
    .Y(_0202_),
    .B1(_0607_));
 sg13g2_and2_2 _2478_ (.A(_0991_),
    .B(_0269_),
    .X(_0608_));
 sg13g2_nor2_2 _2479_ (.A(net162),
    .B(_0608_),
    .Y(_0609_));
 sg13g2_a22oi_1 _2480_ (.Y(_0610_),
    .B1(_0609_),
    .B2(net409),
    .A2(_0608_),
    .A1(net175));
 sg13g2_inv_1 _2481_ (.Y(_0203_),
    .A(_0610_));
 sg13g2_a22oi_1 _2482_ (.Y(_0611_),
    .B1(_0609_),
    .B2(net395),
    .A2(_0608_),
    .A1(net173));
 sg13g2_inv_1 _2483_ (.Y(_0204_),
    .A(_0611_));
 sg13g2_a22oi_1 _2484_ (.Y(_0612_),
    .B1(_0609_),
    .B2(net389),
    .A2(_0608_),
    .A1(net171));
 sg13g2_inv_1 _2485_ (.Y(_0205_),
    .A(_0612_));
 sg13g2_a22oi_1 _2486_ (.Y(_0613_),
    .B1(_0609_),
    .B2(net447),
    .A2(_0608_),
    .A1(net169));
 sg13g2_inv_1 _2487_ (.Y(_0206_),
    .A(_0613_));
 sg13g2_nor2_1 _2488_ (.A(_0750_),
    .B(net163),
    .Y(_0207_));
 sg13g2_and2_1 _2489_ (.A(_0991_),
    .B(_1087_),
    .X(_0614_));
 sg13g2_nor2_2 _2490_ (.A(net162),
    .B(_0614_),
    .Y(_0615_));
 sg13g2_a22oi_1 _2491_ (.Y(_0616_),
    .B1(_0615_),
    .B2(net478),
    .A2(net148),
    .A1(net175));
 sg13g2_inv_1 _2492_ (.Y(_0208_),
    .A(_0616_));
 sg13g2_a22oi_1 _2493_ (.Y(_0617_),
    .B1(_0615_),
    .B2(net464),
    .A2(net148),
    .A1(net173));
 sg13g2_inv_1 _2494_ (.Y(_0209_),
    .A(_0617_));
 sg13g2_a22oi_1 _2495_ (.Y(_0618_),
    .B1(_0615_),
    .B2(net455),
    .A2(net148),
    .A1(net171));
 sg13g2_inv_1 _2496_ (.Y(_0210_),
    .A(_0618_));
 sg13g2_a22oi_1 _2497_ (.Y(_0619_),
    .B1(_0615_),
    .B2(net380),
    .A2(net148),
    .A1(net169));
 sg13g2_inv_1 _2498_ (.Y(_0211_),
    .A(_0619_));
 sg13g2_a22oi_1 _2499_ (.Y(_0620_),
    .B1(_0615_),
    .B2(net467),
    .A2(net148),
    .A1(net168));
 sg13g2_inv_1 _2500_ (.Y(_0212_),
    .A(_0620_));
 sg13g2_a22oi_1 _2501_ (.Y(_0621_),
    .B1(_0615_),
    .B2(net508),
    .A2(net148),
    .A1(net2));
 sg13g2_inv_1 _2502_ (.Y(_0213_),
    .A(_0621_));
 sg13g2_a22oi_1 _2503_ (.Y(_0622_),
    .B1(_0615_),
    .B2(net458),
    .A2(net148),
    .A1(net3));
 sg13g2_inv_1 _2504_ (.Y(_0214_),
    .A(_0622_));
 sg13g2_a22oi_1 _2505_ (.Y(_0623_),
    .B1(_0615_),
    .B2(net521),
    .A2(net148),
    .A1(net4));
 sg13g2_inv_1 _2506_ (.Y(_0215_),
    .A(_0623_));
 sg13g2_nor2_1 _2507_ (.A(\attenuation_A.out[0] ),
    .B(net428),
    .Y(_0624_));
 sg13g2_and2_1 _2508_ (.A(\attenuation_A.out[0] ),
    .B(net428),
    .X(_0625_));
 sg13g2_nor3_1 _2509_ (.A(net163),
    .B(_0624_),
    .C(_0625_),
    .Y(_0216_));
 sg13g2_and2_1 _2510_ (.A(\attenuation_A.out[1] ),
    .B(net609),
    .X(_0626_));
 sg13g2_xor2_1 _2511_ (.B(net609),
    .A(\attenuation_A.out[1] ),
    .X(_0627_));
 sg13g2_nor2_1 _2512_ (.A(_0625_),
    .B(_0627_),
    .Y(_0628_));
 sg13g2_a21oi_1 _2513_ (.A1(_0625_),
    .A2(_0627_),
    .Y(_0629_),
    .B1(net163));
 sg13g2_nor2b_1 _2514_ (.A(_0628_),
    .B_N(_0629_),
    .Y(_0217_));
 sg13g2_xnor2_1 _2515_ (.Y(_0630_),
    .A(\attenuation_A.out[2] ),
    .B(net627));
 sg13g2_a21oi_1 _2516_ (.A1(_0625_),
    .A2(_0627_),
    .Y(_0631_),
    .B1(_0626_));
 sg13g2_and2_1 _2517_ (.A(_0630_),
    .B(_0631_),
    .X(_0632_));
 sg13g2_nor2_1 _2518_ (.A(_0630_),
    .B(_0631_),
    .Y(_0633_));
 sg13g2_nor3_1 _2519_ (.A(net163),
    .B(_0632_),
    .C(_0633_),
    .Y(_0218_));
 sg13g2_nand2_1 _2520_ (.Y(_0634_),
    .A(\attenuation_A.out[3] ),
    .B(net587));
 sg13g2_xnor2_1 _2521_ (.Y(_0635_),
    .A(\attenuation_A.out[3] ),
    .B(net587));
 sg13g2_a21oi_1 _2522_ (.A1(\attenuation_A.out[2] ),
    .A2(\pwm_A.accumulator[2] ),
    .Y(_0636_),
    .B1(_0633_));
 sg13g2_or2_1 _2523_ (.X(_0637_),
    .B(_0636_),
    .A(_0635_));
 sg13g2_nand2_1 _2524_ (.Y(_0638_),
    .A(net184),
    .B(_0637_));
 sg13g2_a21oi_1 _2525_ (.A1(_0635_),
    .A2(_0636_),
    .Y(_0219_),
    .B1(_0638_));
 sg13g2_nand2_1 _2526_ (.Y(_0639_),
    .A(\attenuation_A.out[4] ),
    .B(\pwm_A.accumulator[4] ));
 sg13g2_xnor2_1 _2527_ (.Y(_0640_),
    .A(\attenuation_A.out[4] ),
    .B(net625));
 sg13g2_nand3_1 _2528_ (.B(_0637_),
    .C(_0640_),
    .A(_0634_),
    .Y(_0641_));
 sg13g2_a21o_1 _2529_ (.A2(_0637_),
    .A1(_0634_),
    .B1(_0640_),
    .X(_0642_));
 sg13g2_and3_1 _2530_ (.X(_0220_),
    .A(net184),
    .B(_0641_),
    .C(_0642_));
 sg13g2_and2_1 _2531_ (.A(_0639_),
    .B(_0642_),
    .X(_0643_));
 sg13g2_nor2_1 _2532_ (.A(\attenuation_A.out[5] ),
    .B(net614),
    .Y(_0644_));
 sg13g2_nand2_1 _2533_ (.Y(_0645_),
    .A(\attenuation_A.out[5] ),
    .B(net614));
 sg13g2_nand2b_1 _2534_ (.Y(_0646_),
    .B(_0645_),
    .A_N(_0644_));
 sg13g2_o21ai_1 _2535_ (.B1(net184),
    .Y(_0647_),
    .A1(_0643_),
    .A2(_0646_));
 sg13g2_a21oi_1 _2536_ (.A1(_0643_),
    .A2(_0646_),
    .Y(_0221_),
    .B1(_0647_));
 sg13g2_xor2_1 _2537_ (.B(net626),
    .A(\attenuation_A.out[6] ),
    .X(_0648_));
 sg13g2_o21ai_1 _2538_ (.B1(_0645_),
    .Y(_0649_),
    .A1(_0643_),
    .A2(_0644_));
 sg13g2_and2_1 _2539_ (.A(_0648_),
    .B(_0649_),
    .X(_0650_));
 sg13g2_o21ai_1 _2540_ (.B1(net182),
    .Y(_0651_),
    .A1(_0648_),
    .A2(_0649_));
 sg13g2_nor2_1 _2541_ (.A(_0650_),
    .B(_0651_),
    .Y(_0222_));
 sg13g2_nand2_1 _2542_ (.Y(_0652_),
    .A(\attenuation_A.out[7] ),
    .B(net490));
 sg13g2_xnor2_1 _2543_ (.Y(_0653_),
    .A(\attenuation_A.out[7] ),
    .B(net490));
 sg13g2_a21oi_1 _2544_ (.A1(\attenuation_A.out[6] ),
    .A2(net626),
    .Y(_0654_),
    .B1(_0650_));
 sg13g2_or2_1 _2545_ (.X(_0655_),
    .B(_0654_),
    .A(_0653_));
 sg13g2_a21oi_1 _2546_ (.A1(_0653_),
    .A2(_0654_),
    .Y(_0656_),
    .B1(net165));
 sg13g2_and2_1 _2547_ (.A(_0655_),
    .B(_0656_),
    .X(_0223_));
 sg13g2_a21oi_1 _2548_ (.A1(_0652_),
    .A2(_0655_),
    .Y(_0224_),
    .B1(net167));
 sg13g2_nor2_1 _2549_ (.A(\attenuation_B.out[0] ),
    .B(net481),
    .Y(_0657_));
 sg13g2_and2_1 _2550_ (.A(\attenuation_B.out[0] ),
    .B(net481),
    .X(_0658_));
 sg13g2_nor3_1 _2551_ (.A(net163),
    .B(_0657_),
    .C(_0658_),
    .Y(_0225_));
 sg13g2_and2_1 _2552_ (.A(\attenuation_B.out[1] ),
    .B(\pwm_B.accumulator[1] ),
    .X(_0659_));
 sg13g2_xor2_1 _2553_ (.B(net617),
    .A(\attenuation_B.out[1] ),
    .X(_0660_));
 sg13g2_nor2_1 _2554_ (.A(_0658_),
    .B(_0660_),
    .Y(_0661_));
 sg13g2_a21oi_1 _2555_ (.A1(_0658_),
    .A2(_0660_),
    .Y(_0662_),
    .B1(net163));
 sg13g2_nor2b_1 _2556_ (.A(_0661_),
    .B_N(_0662_),
    .Y(_0226_));
 sg13g2_xnor2_1 _2557_ (.Y(_0663_),
    .A(\attenuation_B.out[2] ),
    .B(net630));
 sg13g2_a21oi_1 _2558_ (.A1(_0658_),
    .A2(_0660_),
    .Y(_0664_),
    .B1(_0659_));
 sg13g2_and2_1 _2559_ (.A(_0663_),
    .B(_0664_),
    .X(_0665_));
 sg13g2_nor2_1 _2560_ (.A(_0663_),
    .B(_0664_),
    .Y(_0666_));
 sg13g2_nor3_1 _2561_ (.A(net163),
    .B(net631),
    .C(_0666_),
    .Y(_0227_));
 sg13g2_nand2_1 _2562_ (.Y(_0667_),
    .A(\attenuation_B.out[3] ),
    .B(net585));
 sg13g2_xnor2_1 _2563_ (.Y(_0668_),
    .A(\attenuation_B.out[3] ),
    .B(net585));
 sg13g2_a21oi_1 _2564_ (.A1(\attenuation_B.out[2] ),
    .A2(\pwm_B.accumulator[2] ),
    .Y(_0669_),
    .B1(_0666_));
 sg13g2_or2_1 _2565_ (.X(_0670_),
    .B(_0669_),
    .A(_0668_));
 sg13g2_nand2_1 _2566_ (.Y(_0671_),
    .A(net184),
    .B(_0670_));
 sg13g2_a21oi_1 _2567_ (.A1(_0668_),
    .A2(_0669_),
    .Y(_0228_),
    .B1(_0671_));
 sg13g2_nand2_1 _2568_ (.Y(_0672_),
    .A(\attenuation_B.out[4] ),
    .B(\pwm_B.accumulator[4] ));
 sg13g2_xnor2_1 _2569_ (.Y(_0673_),
    .A(\attenuation_B.out[4] ),
    .B(\pwm_B.accumulator[4] ));
 sg13g2_nand3_1 _2570_ (.B(_0670_),
    .C(_0673_),
    .A(_0667_),
    .Y(_0674_));
 sg13g2_a21o_1 _2571_ (.A2(_0670_),
    .A1(_0667_),
    .B1(_0673_),
    .X(_0675_));
 sg13g2_and3_1 _2572_ (.X(_0229_),
    .A(net184),
    .B(_0674_),
    .C(_0675_));
 sg13g2_and2_1 _2573_ (.A(_0672_),
    .B(_0675_),
    .X(_0676_));
 sg13g2_nor2_1 _2574_ (.A(\attenuation_B.out[5] ),
    .B(net603),
    .Y(_0677_));
 sg13g2_nand2_1 _2575_ (.Y(_0678_),
    .A(\attenuation_B.out[5] ),
    .B(net603));
 sg13g2_nand2b_1 _2576_ (.Y(_0679_),
    .B(_0678_),
    .A_N(_0677_));
 sg13g2_o21ai_1 _2577_ (.B1(net184),
    .Y(_0680_),
    .A1(_0676_),
    .A2(_0679_));
 sg13g2_a21oi_1 _2578_ (.A1(_0676_),
    .A2(_0679_),
    .Y(_0230_),
    .B1(_0680_));
 sg13g2_xor2_1 _2579_ (.B(net633),
    .A(\attenuation_B.out[6] ),
    .X(_0681_));
 sg13g2_o21ai_1 _2580_ (.B1(_0678_),
    .Y(_0682_),
    .A1(_0676_),
    .A2(_0677_));
 sg13g2_and2_1 _2581_ (.A(_0681_),
    .B(_0682_),
    .X(_0683_));
 sg13g2_o21ai_1 _2582_ (.B1(net182),
    .Y(_0684_),
    .A1(_0681_),
    .A2(_0682_));
 sg13g2_nor2_1 _2583_ (.A(_0683_),
    .B(_0684_),
    .Y(_0231_));
 sg13g2_nand2_1 _2584_ (.Y(_0685_),
    .A(\attenuation_B.out[7] ),
    .B(net517));
 sg13g2_xnor2_1 _2585_ (.Y(_0686_),
    .A(\attenuation_B.out[7] ),
    .B(net517));
 sg13g2_a21oi_1 _2586_ (.A1(\attenuation_B.out[6] ),
    .A2(net633),
    .Y(_0687_),
    .B1(_0683_));
 sg13g2_or2_1 _2587_ (.X(_0688_),
    .B(_0687_),
    .A(_0686_));
 sg13g2_a21oi_1 _2588_ (.A1(_0686_),
    .A2(_0687_),
    .Y(_0689_),
    .B1(net165));
 sg13g2_and2_1 _2589_ (.A(_0688_),
    .B(_0689_),
    .X(_0232_));
 sg13g2_a21oi_1 _2590_ (.A1(_0685_),
    .A2(_0688_),
    .Y(_0233_),
    .B1(net167));
 sg13g2_nor2_1 _2591_ (.A(\attenuation_C.out[0] ),
    .B(net421),
    .Y(_0690_));
 sg13g2_and2_1 _2592_ (.A(\attenuation_C.out[0] ),
    .B(net421),
    .X(_0691_));
 sg13g2_nor3_1 _2593_ (.A(net166),
    .B(_0690_),
    .C(_0691_),
    .Y(_0234_));
 sg13g2_and2_1 _2594_ (.A(\attenuation_C.out[1] ),
    .B(net613),
    .X(_0692_));
 sg13g2_xor2_1 _2595_ (.B(net613),
    .A(\attenuation_C.out[1] ),
    .X(_0693_));
 sg13g2_nor2_1 _2596_ (.A(_0691_),
    .B(_0693_),
    .Y(_0694_));
 sg13g2_a21oi_1 _2597_ (.A1(_0691_),
    .A2(_0693_),
    .Y(_0695_),
    .B1(net165));
 sg13g2_nor2b_1 _2598_ (.A(_0694_),
    .B_N(_0695_),
    .Y(_0235_));
 sg13g2_xnor2_1 _2599_ (.Y(_0696_),
    .A(\attenuation_C.out[2] ),
    .B(net624));
 sg13g2_a21oi_1 _2600_ (.A1(_0691_),
    .A2(_0693_),
    .Y(_0697_),
    .B1(_0692_));
 sg13g2_and2_1 _2601_ (.A(_0696_),
    .B(_0697_),
    .X(_0698_));
 sg13g2_nor2_1 _2602_ (.A(_0696_),
    .B(_0697_),
    .Y(_0699_));
 sg13g2_nor3_1 _2603_ (.A(net165),
    .B(_0698_),
    .C(_0699_),
    .Y(_0236_));
 sg13g2_nand2_1 _2604_ (.Y(_0700_),
    .A(\attenuation_C.out[3] ),
    .B(net583));
 sg13g2_xnor2_1 _2605_ (.Y(_0701_),
    .A(\attenuation_C.out[3] ),
    .B(net583));
 sg13g2_a21oi_1 _2606_ (.A1(\attenuation_C.out[2] ),
    .A2(\pwm_C.accumulator[2] ),
    .Y(_0702_),
    .B1(_0699_));
 sg13g2_or2_1 _2607_ (.X(_0703_),
    .B(_0702_),
    .A(_0701_));
 sg13g2_nand2_1 _2608_ (.Y(_0704_),
    .A(net184),
    .B(_0703_));
 sg13g2_a21oi_1 _2609_ (.A1(_0701_),
    .A2(_0702_),
    .Y(_0237_),
    .B1(_0704_));
 sg13g2_nand2_1 _2610_ (.Y(_0705_),
    .A(\attenuation_C.out[4] ),
    .B(\pwm_C.accumulator[4] ));
 sg13g2_xnor2_1 _2611_ (.Y(_0706_),
    .A(\attenuation_C.out[4] ),
    .B(\pwm_C.accumulator[4] ));
 sg13g2_nand3_1 _2612_ (.B(_0703_),
    .C(_0706_),
    .A(_0700_),
    .Y(_0707_));
 sg13g2_a21o_1 _2613_ (.A2(_0703_),
    .A1(_0700_),
    .B1(_0706_),
    .X(_0708_));
 sg13g2_and3_1 _2614_ (.X(_0238_),
    .A(net182),
    .B(_0707_),
    .C(_0708_));
 sg13g2_and2_1 _2615_ (.A(_0705_),
    .B(_0708_),
    .X(_0709_));
 sg13g2_nor2_1 _2616_ (.A(\attenuation_C.out[5] ),
    .B(net607),
    .Y(_0710_));
 sg13g2_nand2_1 _2617_ (.Y(_0711_),
    .A(\attenuation_C.out[5] ),
    .B(net607));
 sg13g2_nand2b_1 _2618_ (.Y(_0712_),
    .B(_0711_),
    .A_N(_0710_));
 sg13g2_o21ai_1 _2619_ (.B1(net182),
    .Y(_0713_),
    .A1(_0709_),
    .A2(_0712_));
 sg13g2_a21oi_1 _2620_ (.A1(_0709_),
    .A2(_0712_),
    .Y(_0239_),
    .B1(_0713_));
 sg13g2_xor2_1 _2621_ (.B(net618),
    .A(\attenuation_C.out[6] ),
    .X(_0714_));
 sg13g2_o21ai_1 _2622_ (.B1(_0711_),
    .Y(_0715_),
    .A1(_0709_),
    .A2(_0710_));
 sg13g2_and2_1 _2623_ (.A(_0714_),
    .B(_0715_),
    .X(_0716_));
 sg13g2_o21ai_1 _2624_ (.B1(net182),
    .Y(_0717_),
    .A1(_0714_),
    .A2(_0715_));
 sg13g2_nor2_1 _2625_ (.A(_0716_),
    .B(_0717_),
    .Y(_0240_));
 sg13g2_nand2_1 _2626_ (.Y(_0718_),
    .A(\attenuation_C.out[7] ),
    .B(net488));
 sg13g2_xnor2_1 _2627_ (.Y(_0719_),
    .A(\attenuation_C.out[7] ),
    .B(net488));
 sg13g2_a21oi_1 _2628_ (.A1(\attenuation_C.out[6] ),
    .A2(net618),
    .Y(_0720_),
    .B1(_0716_));
 sg13g2_or2_1 _2629_ (.X(_0721_),
    .B(_0720_),
    .A(_0719_));
 sg13g2_a21oi_1 _2630_ (.A1(_0719_),
    .A2(_0720_),
    .Y(_0722_),
    .B1(net165));
 sg13g2_and2_1 _2631_ (.A(_0721_),
    .B(_0722_),
    .X(_0241_));
 sg13g2_a21oi_1 _2632_ (.A1(_0718_),
    .A2(_0721_),
    .Y(_0242_),
    .B1(net165));
 sg13g2_dfrbp_1 _2633_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net318),
    .D(_0024_),
    .Q_N(_1301_),
    .Q(restart_envelope));
 sg13g2_dfrbp_1 _2634_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net263),
    .D(_0025_),
    .Q_N(_1300_),
    .Q(\register[1][0] ));
 sg13g2_dfrbp_1 _2635_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net261),
    .D(_0026_),
    .Q_N(_1299_),
    .Q(\register[1][1] ));
 sg13g2_dfrbp_1 _2636_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net259),
    .D(_0027_),
    .Q_N(_1298_),
    .Q(\register[1][2] ));
 sg13g2_dfrbp_1 _2637_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net257),
    .D(_0028_),
    .Q_N(_1297_),
    .Q(\register[1][3] ));
 sg13g2_dfrbp_1 _2638_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net255),
    .D(_0029_),
    .Q_N(_1296_),
    .Q(\register[2][0] ));
 sg13g2_dfrbp_1 _2639_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net253),
    .D(_0030_),
    .Q_N(_1295_),
    .Q(\register[2][1] ));
 sg13g2_dfrbp_1 _2640_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net251),
    .D(_0031_),
    .Q_N(_1294_),
    .Q(\register[2][2] ));
 sg13g2_dfrbp_1 _2641_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net249),
    .D(_0032_),
    .Q_N(_1293_),
    .Q(\register[2][3] ));
 sg13g2_dfrbp_1 _2642_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net247),
    .D(_0033_),
    .Q_N(_1292_),
    .Q(\register[2][4] ));
 sg13g2_dfrbp_1 _2643_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net245),
    .D(_0034_),
    .Q_N(_1291_),
    .Q(\register[2][5] ));
 sg13g2_dfrbp_1 _2644_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net243),
    .D(_0035_),
    .Q_N(_1290_),
    .Q(\register[2][6] ));
 sg13g2_dfrbp_1 _2645_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net241),
    .D(_0036_),
    .Q_N(_1289_),
    .Q(\register[2][7] ));
 sg13g2_dfrbp_1 _2646_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net239),
    .D(_0037_),
    .Q_N(_1288_),
    .Q(\noise_generator.period[0] ));
 sg13g2_dfrbp_1 _2647_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net237),
    .D(_0038_),
    .Q_N(_1287_),
    .Q(\noise_generator.period[1] ));
 sg13g2_dfrbp_1 _2648_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net235),
    .D(_0039_),
    .Q_N(_1286_),
    .Q(\noise_generator.period[2] ));
 sg13g2_dfrbp_1 _2649_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net233),
    .D(_0040_),
    .Q_N(_1285_),
    .Q(\noise_generator.period[3] ));
 sg13g2_dfrbp_1 _2650_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net231),
    .D(_0041_),
    .Q_N(_1284_),
    .Q(\noise_generator.period[4] ));
 sg13g2_dfrbp_1 _2651_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net229),
    .D(_0042_),
    .Q_N(_1283_),
    .Q(\register[5][0] ));
 sg13g2_dfrbp_1 _2652_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net227),
    .D(_0043_),
    .Q_N(_1282_),
    .Q(\register[5][1] ));
 sg13g2_dfrbp_1 _2653_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net225),
    .D(_0044_),
    .Q_N(_1281_),
    .Q(\register[5][2] ));
 sg13g2_dfrbp_1 _2654_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net223),
    .D(_0045_),
    .Q_N(_1280_),
    .Q(\register[5][3] ));
 sg13g2_dfrbp_1 _2655_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net221),
    .D(_0046_),
    .Q_N(_1279_),
    .Q(\pwm_master.accumulator[0] ));
 sg13g2_dfrbp_1 _2656_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net220),
    .D(net573),
    .Q_N(_1278_),
    .Q(\pwm_master.accumulator[1] ));
 sg13g2_dfrbp_1 _2657_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net219),
    .D(_0048_),
    .Q_N(_1277_),
    .Q(\pwm_master.accumulator[2] ));
 sg13g2_dfrbp_1 _2658_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net218),
    .D(net606),
    .Q_N(_1276_),
    .Q(\pwm_master.accumulator[3] ));
 sg13g2_dfrbp_1 _2659_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net217),
    .D(_0050_),
    .Q_N(_1275_),
    .Q(\pwm_master.accumulator[4] ));
 sg13g2_dfrbp_1 _2660_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net216),
    .D(_0051_),
    .Q_N(_1274_),
    .Q(\pwm_master.accumulator[5] ));
 sg13g2_dfrbp_1 _2661_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net215),
    .D(_0052_),
    .Q_N(_1273_),
    .Q(\pwm_master.accumulator[6] ));
 sg13g2_dfrbp_1 _2662_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net214),
    .D(net623),
    .Q_N(_1272_),
    .Q(\pwm_master.accumulator[7] ));
 sg13g2_dfrbp_1 _2663_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net213),
    .D(_0054_),
    .Q_N(_1271_),
    .Q(\pwm_master.accumulator[8] ));
 sg13g2_dfrbp_1 _2664_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net212),
    .D(net569),
    .Q_N(_1270_),
    .Q(\pwm_master.accumulator[9] ));
 sg13g2_dfrbp_1 _2665_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net211),
    .D(_0056_),
    .Q_N(_1269_),
    .Q(\latched_register[0] ));
 sg13g2_dfrbp_1 _2666_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net209),
    .D(_0057_),
    .Q_N(_1268_),
    .Q(\latched_register[1] ));
 sg13g2_dfrbp_1 _2667_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net207),
    .D(_0058_),
    .Q_N(_1267_),
    .Q(\latched_register[2] ));
 sg13g2_dfrbp_1 _2668_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net205),
    .D(_0059_),
    .Q_N(_1266_),
    .Q(\latched_register[3] ));
 sg13g2_dfrbp_1 _2669_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net203),
    .D(_0060_),
    .Q_N(_1265_),
    .Q(active));
 sg13g2_dfrbp_1 _2670_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net201),
    .D(_0061_),
    .Q_N(_0023_),
    .Q(\clk_counter[0] ));
 sg13g2_dfrbp_1 _2671_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net200),
    .D(_0062_),
    .Q_N(_1264_),
    .Q(\clk_counter[1] ));
 sg13g2_dfrbp_1 _2672_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net199),
    .D(net420),
    .Q_N(_1263_),
    .Q(\clk_counter[2] ));
 sg13g2_dfrbp_1 _2673_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net198),
    .D(_0064_),
    .Q_N(_1262_),
    .Q(\clk_counter[3] ));
 sg13g2_dfrbp_1 _2674_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net197),
    .D(_0065_),
    .Q_N(_1261_),
    .Q(\clk_counter[4] ));
 sg13g2_dfrbp_1 _2675_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net196),
    .D(_0066_),
    .Q_N(_1260_),
    .Q(\clk_counter[5] ));
 sg13g2_dfrbp_1 _2676_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net195),
    .D(net452),
    .Q_N(_1259_),
    .Q(\clk_counter[6] ));
 sg13g2_dfrbp_1 _2677_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net194),
    .D(_0068_),
    .Q_N(_1258_),
    .Q(\envelope_generator.hold ));
 sg13g2_dfrbp_1 _2678_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net192),
    .D(_0069_),
    .Q_N(_1257_),
    .Q(envelope_alternate));
 sg13g2_dfrbp_1 _2679_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net190),
    .D(_0070_),
    .Q_N(_0008_),
    .Q(envelope_attack));
 sg13g2_dfrbp_1 _2680_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net188),
    .D(_0071_),
    .Q_N(_1256_),
    .Q(envelope_continue));
 sg13g2_dfrbp_1 _2681_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net141),
    .D(_0072_),
    .Q_N(_1255_),
    .Q(\envelope_generator.period[8] ));
 sg13g2_dfrbp_1 _2682_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net139),
    .D(_0073_),
    .Q_N(_1254_),
    .Q(\envelope_generator.period[9] ));
 sg13g2_dfrbp_1 _2683_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net137),
    .D(_0074_),
    .Q_N(_1253_),
    .Q(\envelope_generator.period[10] ));
 sg13g2_dfrbp_1 _2684_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net135),
    .D(_0075_),
    .Q_N(_1252_),
    .Q(\envelope_generator.period[11] ));
 sg13g2_dfrbp_1 _2685_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net133),
    .D(_0076_),
    .Q_N(_1251_),
    .Q(\envelope_generator.period[12] ));
 sg13g2_dfrbp_1 _2686_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net131),
    .D(_0077_),
    .Q_N(_1250_),
    .Q(\envelope_generator.period[13] ));
 sg13g2_dfrbp_1 _2687_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net129),
    .D(_0078_),
    .Q_N(_1249_),
    .Q(\envelope_generator.period[14] ));
 sg13g2_dfrbp_1 _2688_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net127),
    .D(_0079_),
    .Q_N(_1248_),
    .Q(\envelope_generator.period[15] ));
 sg13g2_dfrbp_1 _2689_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net125),
    .D(_0080_),
    .Q_N(_0020_),
    .Q(\amplitude_C[0] ));
 sg13g2_dfrbp_1 _2690_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net123),
    .D(_0081_),
    .Q_N(_0021_),
    .Q(\amplitude_C[1] ));
 sg13g2_dfrbp_1 _2691_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net121),
    .D(_0082_),
    .Q_N(_0018_),
    .Q(\amplitude_C[2] ));
 sg13g2_dfrbp_1 _2692_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net119),
    .D(_0083_),
    .Q_N(_0019_),
    .Q(\amplitude_C[3] ));
 sg13g2_dfrbp_1 _2693_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net117),
    .D(_0084_),
    .Q_N(_1247_),
    .Q(envelope_C));
 sg13g2_dfrbp_1 _2694_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net115),
    .D(_0085_),
    .Q_N(_1246_),
    .Q(\envelope_generator.period[0] ));
 sg13g2_dfrbp_1 _2695_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net113),
    .D(_0086_),
    .Q_N(_1245_),
    .Q(\envelope_generator.period[1] ));
 sg13g2_dfrbp_1 _2696_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net111),
    .D(_0087_),
    .Q_N(_1244_),
    .Q(\envelope_generator.period[2] ));
 sg13g2_dfrbp_1 _2697_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net109),
    .D(_0088_),
    .Q_N(_1243_),
    .Q(\envelope_generator.period[3] ));
 sg13g2_dfrbp_1 _2698_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net107),
    .D(_0089_),
    .Q_N(_1242_),
    .Q(\envelope_generator.period[4] ));
 sg13g2_dfrbp_1 _2699_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net105),
    .D(_0090_),
    .Q_N(_1241_),
    .Q(\envelope_generator.period[5] ));
 sg13g2_dfrbp_1 _2700_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net103),
    .D(_0091_),
    .Q_N(_1240_),
    .Q(\envelope_generator.period[6] ));
 sg13g2_dfrbp_1 _2701_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net101),
    .D(_0092_),
    .Q_N(_1239_),
    .Q(\envelope_generator.period[7] ));
 sg13g2_dfrbp_1 _2702_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net99),
    .D(net383),
    .Q_N(_0005_),
    .Q(tone_A));
 sg13g2_dfrbp_1 _2703_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net97),
    .D(_0094_),
    .Q_N(_1238_),
    .Q(\tone_A_generator.counter[0] ));
 sg13g2_dfrbp_1 _2704_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net95),
    .D(_0095_),
    .Q_N(_1237_),
    .Q(\tone_A_generator.counter[1] ));
 sg13g2_dfrbp_1 _2705_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net93),
    .D(_0096_),
    .Q_N(_1236_),
    .Q(\tone_A_generator.counter[2] ));
 sg13g2_dfrbp_1 _2706_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net91),
    .D(_0097_),
    .Q_N(_1235_),
    .Q(\tone_A_generator.counter[3] ));
 sg13g2_dfrbp_1 _2707_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net89),
    .D(_0098_),
    .Q_N(_1234_),
    .Q(\tone_A_generator.counter[4] ));
 sg13g2_dfrbp_1 _2708_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net87),
    .D(_0099_),
    .Q_N(_1233_),
    .Q(\tone_A_generator.counter[5] ));
 sg13g2_dfrbp_1 _2709_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net85),
    .D(_0100_),
    .Q_N(_1232_),
    .Q(\tone_A_generator.counter[6] ));
 sg13g2_dfrbp_1 _2710_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net83),
    .D(_0101_),
    .Q_N(_1231_),
    .Q(\tone_A_generator.counter[7] ));
 sg13g2_dfrbp_1 _2711_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net81),
    .D(_0102_),
    .Q_N(_1230_),
    .Q(\tone_A_generator.counter[8] ));
 sg13g2_dfrbp_1 _2712_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net79),
    .D(_0103_),
    .Q_N(_1229_),
    .Q(\tone_A_generator.counter[9] ));
 sg13g2_dfrbp_1 _2713_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net77),
    .D(_0104_),
    .Q_N(_1228_),
    .Q(\tone_A_generator.counter[10] ));
 sg13g2_dfrbp_1 _2714_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net75),
    .D(_0105_),
    .Q_N(_1227_),
    .Q(\tone_A_generator.counter[11] ));
 sg13g2_dfrbp_1 _2715_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net73),
    .D(net344),
    .Q_N(_0006_),
    .Q(tone_B));
 sg13g2_dfrbp_1 _2716_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net71),
    .D(_0107_),
    .Q_N(_1226_),
    .Q(\tone_B_generator.counter[0] ));
 sg13g2_dfrbp_1 _2717_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net69),
    .D(net444),
    .Q_N(_1225_),
    .Q(\tone_B_generator.counter[1] ));
 sg13g2_dfrbp_1 _2718_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net67),
    .D(_0109_),
    .Q_N(_1224_),
    .Q(\tone_B_generator.counter[2] ));
 sg13g2_dfrbp_1 _2719_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net65),
    .D(_0110_),
    .Q_N(_1223_),
    .Q(\tone_B_generator.counter[3] ));
 sg13g2_dfrbp_1 _2720_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net63),
    .D(_0111_),
    .Q_N(_1222_),
    .Q(\tone_B_generator.counter[4] ));
 sg13g2_dfrbp_1 _2721_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net61),
    .D(_0112_),
    .Q_N(_1221_),
    .Q(\tone_B_generator.counter[5] ));
 sg13g2_dfrbp_1 _2722_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net59),
    .D(_0113_),
    .Q_N(_1220_),
    .Q(\tone_B_generator.counter[6] ));
 sg13g2_dfrbp_1 _2723_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net57),
    .D(_0114_),
    .Q_N(_1219_),
    .Q(\tone_B_generator.counter[7] ));
 sg13g2_dfrbp_1 _2724_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net55),
    .D(_0115_),
    .Q_N(_1218_),
    .Q(\tone_B_generator.counter[8] ));
 sg13g2_dfrbp_1 _2725_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net53),
    .D(_0116_),
    .Q_N(_1217_),
    .Q(\tone_B_generator.counter[9] ));
 sg13g2_dfrbp_1 _2726_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net51),
    .D(_0117_),
    .Q_N(_1216_),
    .Q(\tone_B_generator.counter[10] ));
 sg13g2_dfrbp_1 _2727_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net49),
    .D(_0118_),
    .Q_N(_1215_),
    .Q(\tone_B_generator.counter[11] ));
 sg13g2_dfrbp_1 _2728_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net47),
    .D(_0119_),
    .Q_N(_0012_),
    .Q(\amplitude_A[0] ));
 sg13g2_dfrbp_1 _2729_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net45),
    .D(_0120_),
    .Q_N(_0013_),
    .Q(\amplitude_A[1] ));
 sg13g2_dfrbp_1 _2730_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net43),
    .D(_0121_),
    .Q_N(_0010_),
    .Q(\amplitude_A[2] ));
 sg13g2_dfrbp_1 _2731_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net41),
    .D(_0122_),
    .Q_N(_0011_),
    .Q(\amplitude_A[3] ));
 sg13g2_dfrbp_1 _2732_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net327),
    .D(_0123_),
    .Q_N(_1214_),
    .Q(envelope_A));
 sg13g2_dfrbp_1 _2733_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net325),
    .D(net356),
    .Q_N(_0007_),
    .Q(tone_C));
 sg13g2_dfrbp_1 _2734_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net323),
    .D(_0125_),
    .Q_N(_1213_),
    .Q(\tone_C_generator.counter[0] ));
 sg13g2_dfrbp_1 _2735_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net321),
    .D(net484),
    .Q_N(_1212_),
    .Q(\tone_C_generator.counter[1] ));
 sg13g2_dfrbp_1 _2736_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net319),
    .D(_0127_),
    .Q_N(_1211_),
    .Q(\tone_C_generator.counter[2] ));
 sg13g2_dfrbp_1 _2737_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net317),
    .D(_0128_),
    .Q_N(_1210_),
    .Q(\tone_C_generator.counter[3] ));
 sg13g2_dfrbp_1 _2738_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net315),
    .D(_0129_),
    .Q_N(_1209_),
    .Q(\tone_C_generator.counter[4] ));
 sg13g2_dfrbp_1 _2739_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net313),
    .D(_0130_),
    .Q_N(_1208_),
    .Q(\tone_C_generator.counter[5] ));
 sg13g2_dfrbp_1 _2740_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net311),
    .D(_0131_),
    .Q_N(_1207_),
    .Q(\tone_C_generator.counter[6] ));
 sg13g2_dfrbp_1 _2741_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net309),
    .D(_0132_),
    .Q_N(_1206_),
    .Q(\tone_C_generator.counter[7] ));
 sg13g2_dfrbp_1 _2742_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net307),
    .D(_0133_),
    .Q_N(_1205_),
    .Q(\tone_C_generator.counter[8] ));
 sg13g2_dfrbp_1 _2743_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net305),
    .D(_0134_),
    .Q_N(_1204_),
    .Q(\tone_C_generator.counter[9] ));
 sg13g2_dfrbp_1 _2744_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net303),
    .D(_0135_),
    .Q_N(_1203_),
    .Q(\tone_C_generator.counter[10] ));
 sg13g2_dfrbp_1 _2745_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net301),
    .D(_0136_),
    .Q_N(_1202_),
    .Q(\tone_C_generator.counter[11] ));
 sg13g2_dfrbp_1 _2746_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net299),
    .D(_0137_),
    .Q_N(_1201_),
    .Q(tone_disable_A));
 sg13g2_dfrbp_1 _2747_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net297),
    .D(_0138_),
    .Q_N(_1200_),
    .Q(tone_disable_B));
 sg13g2_dfrbp_1 _2748_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net295),
    .D(_0139_),
    .Q_N(_1199_),
    .Q(tone_disable_C));
 sg13g2_dfrbp_1 _2749_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net293),
    .D(_0140_),
    .Q_N(_1198_),
    .Q(noise_disable_A));
 sg13g2_dfrbp_1 _2750_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net267),
    .D(_0141_),
    .Q_N(_1197_),
    .Q(noise_disable_B));
 sg13g2_dfrbp_1 _2751_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net265),
    .D(_0142_),
    .Q_N(_1196_),
    .Q(noise_disable_C));
 sg13g2_dfrbp_1 _2752_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net262),
    .D(_0143_),
    .Q_N(_0016_),
    .Q(\amplitude_B[0] ));
 sg13g2_dfrbp_1 _2753_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net258),
    .D(_0144_),
    .Q_N(_0017_),
    .Q(\amplitude_B[1] ));
 sg13g2_dfrbp_1 _2754_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net254),
    .D(_0145_),
    .Q_N(_0014_),
    .Q(\amplitude_B[2] ));
 sg13g2_dfrbp_1 _2755_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net250),
    .D(_0146_),
    .Q_N(_0015_),
    .Q(\amplitude_B[3] ));
 sg13g2_dfrbp_1 _2756_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net246),
    .D(_0147_),
    .Q_N(_1195_),
    .Q(envelope_B));
 sg13g2_dfrbp_1 _2757_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net242),
    .D(net388),
    .Q_N(_1194_),
    .Q(\envelope_generator.signal_edge.previous_signal_state_0 ));
 sg13g2_dfrbp_1 _2758_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net240),
    .D(_0149_),
    .Q_N(_1193_),
    .Q(\noise_generator.tone.counter[0] ));
 sg13g2_dfrbp_1 _2759_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net236),
    .D(net377),
    .Q_N(_1192_),
    .Q(\noise_generator.tone.counter[1] ));
 sg13g2_dfrbp_1 _2760_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net232),
    .D(_0151_),
    .Q_N(_1191_),
    .Q(\noise_generator.tone.counter[2] ));
 sg13g2_dfrbp_1 _2761_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net228),
    .D(_0152_),
    .Q_N(_1190_),
    .Q(\noise_generator.tone.counter[3] ));
 sg13g2_dfrbp_1 _2762_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net224),
    .D(_0153_),
    .Q_N(_1189_),
    .Q(\noise_generator.tone.counter[4] ));
 sg13g2_dfrbp_1 _2763_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net210),
    .D(net374),
    .Q_N(_0004_),
    .Q(\noise_generator.signal_edge.signal ));
 sg13g2_dfrbp_1 _2764_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net206),
    .D(net435),
    .Q_N(_1188_),
    .Q(\noise_generator.lfsr[0] ));
 sg13g2_dfrbp_1 _2765_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net202),
    .D(_0156_),
    .Q_N(_1187_),
    .Q(\noise_generator.lfsr[1] ));
 sg13g2_dfrbp_1 _2766_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net191),
    .D(net500),
    .Q_N(_1186_),
    .Q(\noise_generator.lfsr[2] ));
 sg13g2_dfrbp_1 _2767_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net187),
    .D(net463),
    .Q_N(_1185_),
    .Q(\noise_generator.lfsr[3] ));
 sg13g2_dfrbp_1 _2768_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net138),
    .D(_0159_),
    .Q_N(_1184_),
    .Q(\noise_generator.lfsr[4] ));
 sg13g2_dfrbp_1 _2769_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net134),
    .D(net474),
    .Q_N(_1183_),
    .Q(\noise_generator.lfsr[5] ));
 sg13g2_dfrbp_1 _2770_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net130),
    .D(net460),
    .Q_N(_1182_),
    .Q(\noise_generator.lfsr[6] ));
 sg13g2_dfrbp_1 _2771_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net126),
    .D(net457),
    .Q_N(_1181_),
    .Q(\noise_generator.lfsr[7] ));
 sg13g2_dfrbp_1 _2772_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net122),
    .D(net417),
    .Q_N(_1180_),
    .Q(\noise_generator.lfsr[8] ));
 sg13g2_dfrbp_1 _2773_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net118),
    .D(_0164_),
    .Q_N(_1179_),
    .Q(\noise_generator.lfsr[9] ));
 sg13g2_dfrbp_1 _2774_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net114),
    .D(net450),
    .Q_N(_1178_),
    .Q(\noise_generator.lfsr[10] ));
 sg13g2_dfrbp_1 _2775_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net110),
    .D(_0166_),
    .Q_N(_1177_),
    .Q(\noise_generator.lfsr[11] ));
 sg13g2_dfrbp_1 _2776_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net106),
    .D(net454),
    .Q_N(_1176_),
    .Q(\noise_generator.lfsr[12] ));
 sg13g2_dfrbp_1 _2777_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net102),
    .D(_0168_),
    .Q_N(_1175_),
    .Q(\noise_generator.lfsr[13] ));
 sg13g2_dfrbp_1 _2778_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net98),
    .D(net433),
    .Q_N(_1174_),
    .Q(\noise_generator.lfsr[14] ));
 sg13g2_dfrbp_1 _2779_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net94),
    .D(net470),
    .Q_N(_1173_),
    .Q(\noise_generator.lfsr[15] ));
 sg13g2_dfrbp_1 _2780_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net90),
    .D(net532),
    .Q_N(_1172_),
    .Q(\noise_generator.lfsr[16] ));
 sg13g2_dfrbp_1 _2781_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net86),
    .D(_0172_),
    .Q_N(_1171_),
    .Q(\register[4][0] ));
 sg13g2_dfrbp_1 _2782_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net82),
    .D(_0173_),
    .Q_N(_1170_),
    .Q(\register[4][1] ));
 sg13g2_dfrbp_1 _2783_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net78),
    .D(_0174_),
    .Q_N(_1169_),
    .Q(\register[4][2] ));
 sg13g2_dfrbp_1 _2784_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net74),
    .D(_0175_),
    .Q_N(_1168_),
    .Q(\register[4][3] ));
 sg13g2_dfrbp_1 _2785_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net70),
    .D(_0176_),
    .Q_N(_1167_),
    .Q(\register[4][4] ));
 sg13g2_dfrbp_1 _2786_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net66),
    .D(_0177_),
    .Q_N(_1166_),
    .Q(\register[4][5] ));
 sg13g2_dfrbp_1 _2787_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net62),
    .D(_0178_),
    .Q_N(_1165_),
    .Q(\register[4][6] ));
 sg13g2_dfrbp_1 _2788_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net58),
    .D(_0179_),
    .Q_N(_1164_),
    .Q(\register[4][7] ));
 sg13g2_dfrbp_1 _2789_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net54),
    .D(net337),
    .Q_N(_0009_),
    .Q(\envelope_generator.invert_output ));
 sg13g2_dfrbp_1 _2790_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net52),
    .D(_0181_),
    .Q_N(_1163_),
    .Q(\envelope_generator.tone.counter[0] ));
 sg13g2_dfrbp_1 _2791_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net48),
    .D(net431),
    .Q_N(_1162_),
    .Q(\envelope_generator.tone.counter[1] ));
 sg13g2_dfrbp_1 _2792_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net44),
    .D(_0183_),
    .Q_N(_1161_),
    .Q(\envelope_generator.tone.counter[2] ));
 sg13g2_dfrbp_1 _2793_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net328),
    .D(_0184_),
    .Q_N(_1160_),
    .Q(\envelope_generator.tone.counter[3] ));
 sg13g2_dfrbp_1 _2794_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net324),
    .D(net546),
    .Q_N(_1159_),
    .Q(\envelope_generator.tone.counter[4] ));
 sg13g2_dfrbp_1 _2795_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net320),
    .D(_0186_),
    .Q_N(_1158_),
    .Q(\envelope_generator.tone.counter[5] ));
 sg13g2_dfrbp_1 _2796_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net316),
    .D(net493),
    .Q_N(_1157_),
    .Q(\envelope_generator.tone.counter[6] ));
 sg13g2_dfrbp_1 _2797_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net312),
    .D(_0188_),
    .Q_N(_1156_),
    .Q(\envelope_generator.tone.counter[7] ));
 sg13g2_dfrbp_1 _2798_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net308),
    .D(_0189_),
    .Q_N(_1155_),
    .Q(\envelope_generator.tone.counter[8] ));
 sg13g2_dfrbp_1 _2799_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net304),
    .D(_0190_),
    .Q_N(_1154_),
    .Q(\envelope_generator.tone.counter[9] ));
 sg13g2_dfrbp_1 _2800_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net300),
    .D(net525),
    .Q_N(_1153_),
    .Q(\envelope_generator.tone.counter[10] ));
 sg13g2_dfrbp_1 _2801_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net296),
    .D(_0192_),
    .Q_N(_1152_),
    .Q(\envelope_generator.tone.counter[11] ));
 sg13g2_dfrbp_1 _2802_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net268),
    .D(_0193_),
    .Q_N(_1151_),
    .Q(\envelope_generator.tone.counter[12] ));
 sg13g2_dfrbp_1 _2803_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net264),
    .D(net399),
    .Q_N(_1150_),
    .Q(\envelope_generator.tone.counter[13] ));
 sg13g2_dfrbp_1 _2804_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net256),
    .D(_0195_),
    .Q_N(_1149_),
    .Q(\envelope_generator.tone.counter[14] ));
 sg13g2_dfrbp_1 _2805_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net248),
    .D(_0196_),
    .Q_N(_1148_),
    .Q(\envelope_generator.tone.counter[15] ));
 sg13g2_dfrbp_1 _2806_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net238),
    .D(net369),
    .Q_N(_0003_),
    .Q(\envelope_generator.signal_edge.signal ));
 sg13g2_dfrbp_1 _2807_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net230),
    .D(net487),
    .Q_N(_1147_),
    .Q(\envelope_generator.stop ));
 sg13g2_dfrbp_1 _2808_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net222),
    .D(net335),
    .Q_N(_0022_),
    .Q(\envelope_generator.envelope_counter[0] ));
 sg13g2_dfrbp_1 _2809_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net204),
    .D(net515),
    .Q_N(_1146_),
    .Q(\envelope_generator.envelope_counter[1] ));
 sg13g2_dfrbp_1 _2810_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net189),
    .D(_0201_),
    .Q_N(_1145_),
    .Q(\envelope_generator.envelope_counter[2] ));
 sg13g2_dfrbp_1 _2811_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net136),
    .D(net497),
    .Q_N(_1144_),
    .Q(\envelope_generator.envelope_counter[3] ));
 sg13g2_dfrbp_1 _2812_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net128),
    .D(_0203_),
    .Q_N(_1143_),
    .Q(\register[3][0] ));
 sg13g2_dfrbp_1 _2813_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net120),
    .D(_0204_),
    .Q_N(_1142_),
    .Q(\register[3][1] ));
 sg13g2_dfrbp_1 _2814_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net112),
    .D(_0205_),
    .Q_N(_1141_),
    .Q(\register[3][2] ));
 sg13g2_dfrbp_1 _2815_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net104),
    .D(_0206_),
    .Q_N(_1140_),
    .Q(\register[3][3] ));
 sg13g2_dllrq_1 _2816_ (.D(_0243_),
    .GATE_N(net33),
    .RESET_B(net269),
    .Q(\attenuation_A.out[0] ));
 sg13g2_dllrq_1 _2817_ (.D(_0244_),
    .GATE_N(net34),
    .RESET_B(net270),
    .Q(\attenuation_A.out[1] ));
 sg13g2_dllrq_1 _2818_ (.D(_0245_),
    .GATE_N(net35),
    .RESET_B(net271),
    .Q(\attenuation_A.out[2] ));
 sg13g2_dllrq_1 _2819_ (.D(_0246_),
    .GATE_N(net36),
    .RESET_B(net272),
    .Q(\attenuation_A.out[3] ));
 sg13g2_dllrq_1 _2820_ (.D(_0247_),
    .GATE_N(net37),
    .RESET_B(net273),
    .Q(\attenuation_A.out[4] ));
 sg13g2_dllrq_1 _2821_ (.D(_0248_),
    .GATE_N(net38),
    .RESET_B(net274),
    .Q(\attenuation_A.out[5] ));
 sg13g2_dllrq_1 _2822_ (.D(_0249_),
    .GATE_N(net39),
    .RESET_B(net275),
    .Q(\attenuation_A.out[6] ));
 sg13g2_dllrq_1 _2823_ (.D(_0250_),
    .GATE_N(net40),
    .RESET_B(net276),
    .Q(\attenuation_A.out[7] ));
 sg13g2_dllrq_1 _2824_ (.D(_0251_),
    .GATE_N(net25),
    .RESET_B(net277),
    .Q(\attenuation_B.out[0] ));
 sg13g2_dllrq_1 _2825_ (.D(_0252_),
    .GATE_N(net26),
    .RESET_B(net278),
    .Q(\attenuation_B.out[1] ));
 sg13g2_dllrq_1 _2826_ (.D(_0253_),
    .GATE_N(net27),
    .RESET_B(net279),
    .Q(\attenuation_B.out[2] ));
 sg13g2_dllrq_1 _2827_ (.D(_0254_),
    .GATE_N(net28),
    .RESET_B(net280),
    .Q(\attenuation_B.out[3] ));
 sg13g2_dllrq_1 _2828_ (.D(_0255_),
    .GATE_N(net29),
    .RESET_B(net281),
    .Q(\attenuation_B.out[4] ));
 sg13g2_dllrq_1 _2829_ (.D(_0256_),
    .GATE_N(net30),
    .RESET_B(net282),
    .Q(\attenuation_B.out[5] ));
 sg13g2_dllrq_1 _2830_ (.D(_0257_),
    .GATE_N(net31),
    .RESET_B(net283),
    .Q(\attenuation_B.out[6] ));
 sg13g2_dllrq_1 _2831_ (.D(_0258_),
    .GATE_N(net32),
    .RESET_B(net284),
    .Q(\attenuation_B.out[7] ));
 sg13g2_dllrq_1 _2832_ (.D(_0259_),
    .GATE_N(net17),
    .RESET_B(net285),
    .Q(\attenuation_C.out[0] ));
 sg13g2_dllrq_1 _2833_ (.D(_0260_),
    .GATE_N(net18),
    .RESET_B(net286),
    .Q(\attenuation_C.out[1] ));
 sg13g2_dllrq_1 _2834_ (.D(_0261_),
    .GATE_N(net19),
    .RESET_B(net287),
    .Q(\attenuation_C.out[2] ));
 sg13g2_dllrq_1 _2835_ (.D(_0262_),
    .GATE_N(net20),
    .RESET_B(net288),
    .Q(\attenuation_C.out[3] ));
 sg13g2_dllrq_1 _2836_ (.D(_0263_),
    .GATE_N(net21),
    .RESET_B(net289),
    .Q(\attenuation_C.out[4] ));
 sg13g2_dllrq_1 _2837_ (.D(_0264_),
    .GATE_N(net22),
    .RESET_B(net290),
    .Q(\attenuation_C.out[5] ));
 sg13g2_dllrq_1 _2838_ (.D(_0265_),
    .GATE_N(net23),
    .RESET_B(net291),
    .Q(\attenuation_C.out[6] ));
 sg13g2_dllrq_1 _2839_ (.D(_0266_),
    .GATE_N(net24),
    .RESET_B(net292),
    .Q(\attenuation_C.out[7] ));
 sg13g2_dfrbp_1 _2840_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net96),
    .D(_0207_),
    .Q_N(_1139_),
    .Q(\noise_generator.signal_edge.previous_signal_state_0 ));
 sg13g2_dfrbp_1 _2841_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net92),
    .D(_0208_),
    .Q_N(_1138_),
    .Q(\register[0][0] ));
 sg13g2_dfrbp_1 _2842_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net84),
    .D(_0209_),
    .Q_N(_1137_),
    .Q(\register[0][1] ));
 sg13g2_dfrbp_1 _2843_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net76),
    .D(_0210_),
    .Q_N(_1136_),
    .Q(\register[0][2] ));
 sg13g2_dfrbp_1 _2844_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net68),
    .D(_0211_),
    .Q_N(_1135_),
    .Q(\register[0][3] ));
 sg13g2_dfrbp_1 _2845_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net60),
    .D(_0212_),
    .Q_N(_1134_),
    .Q(\register[0][4] ));
 sg13g2_dfrbp_1 _2846_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net50),
    .D(_0213_),
    .Q_N(_1133_),
    .Q(\register[0][5] ));
 sg13g2_dfrbp_1 _2847_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net42),
    .D(_0214_),
    .Q_N(_1132_),
    .Q(\register[0][6] ));
 sg13g2_dfrbp_1 _2848_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net322),
    .D(_0215_),
    .Q_N(_1131_),
    .Q(\register[0][7] ));
 sg13g2_dfrbp_1 _2849_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net314),
    .D(_0216_),
    .Q_N(_1130_),
    .Q(\pwm_A.accumulator[0] ));
 sg13g2_dfrbp_1 _2850_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net310),
    .D(_0217_),
    .Q_N(_1129_),
    .Q(\pwm_A.accumulator[1] ));
 sg13g2_dfrbp_1 _2851_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net306),
    .D(_0218_),
    .Q_N(_1128_),
    .Q(\pwm_A.accumulator[2] ));
 sg13g2_dfrbp_1 _2852_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net302),
    .D(net588),
    .Q_N(_1127_),
    .Q(\pwm_A.accumulator[3] ));
 sg13g2_dfrbp_1 _2853_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net298),
    .D(_0220_),
    .Q_N(_1126_),
    .Q(\pwm_A.accumulator[4] ));
 sg13g2_dfrbp_1 _2854_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net294),
    .D(net615),
    .Q_N(_1125_),
    .Q(\pwm_A.accumulator[5] ));
 sg13g2_dfrbp_1 _2855_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net266),
    .D(_0222_),
    .Q_N(_1124_),
    .Q(\pwm_A.accumulator[6] ));
 sg13g2_dfrbp_1 _2856_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net260),
    .D(_0223_),
    .Q_N(_1123_),
    .Q(\pwm_A.accumulator[7] ));
 sg13g2_dfrbp_1 _2857_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net252),
    .D(_0224_),
    .Q_N(_1122_),
    .Q(\pwm_A.accumulator[8] ));
 sg13g2_dfrbp_1 _2858_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net244),
    .D(_0225_),
    .Q_N(_1121_),
    .Q(\pwm_B.accumulator[0] ));
 sg13g2_dfrbp_1 _2859_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net234),
    .D(_0226_),
    .Q_N(_1120_),
    .Q(\pwm_B.accumulator[1] ));
 sg13g2_dfrbp_1 _2860_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net226),
    .D(net632),
    .Q_N(_1119_),
    .Q(\pwm_B.accumulator[2] ));
 sg13g2_dfrbp_1 _2861_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net208),
    .D(net586),
    .Q_N(_1118_),
    .Q(\pwm_B.accumulator[3] ));
 sg13g2_dfrbp_1 _2862_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net193),
    .D(_0229_),
    .Q_N(_1117_),
    .Q(\pwm_B.accumulator[4] ));
 sg13g2_dfrbp_1 _2863_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net140),
    .D(net604),
    .Q_N(_1116_),
    .Q(\pwm_B.accumulator[5] ));
 sg13g2_dfrbp_1 _2864_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net132),
    .D(_0231_),
    .Q_N(_1115_),
    .Q(\pwm_B.accumulator[6] ));
 sg13g2_dfrbp_1 _2865_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net124),
    .D(_0232_),
    .Q_N(_1114_),
    .Q(\pwm_B.accumulator[7] ));
 sg13g2_dfrbp_1 _2866_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net116),
    .D(_0233_),
    .Q_N(_1113_),
    .Q(\pwm_B.accumulator[8] ));
 sg13g2_dfrbp_1 _2867_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net108),
    .D(_0234_),
    .Q_N(_1112_),
    .Q(\pwm_C.accumulator[0] ));
 sg13g2_dfrbp_1 _2868_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net100),
    .D(_0235_),
    .Q_N(_1111_),
    .Q(\pwm_C.accumulator[1] ));
 sg13g2_dfrbp_1 _2869_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net88),
    .D(_0236_),
    .Q_N(_1110_),
    .Q(\pwm_C.accumulator[2] ));
 sg13g2_dfrbp_1 _2870_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net80),
    .D(net584),
    .Q_N(_1109_),
    .Q(\pwm_C.accumulator[3] ));
 sg13g2_dfrbp_1 _2871_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net72),
    .D(_0238_),
    .Q_N(_1108_),
    .Q(\pwm_C.accumulator[4] ));
 sg13g2_dfrbp_1 _2872_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net64),
    .D(net608),
    .Q_N(_1107_),
    .Q(\pwm_C.accumulator[5] ));
 sg13g2_dfrbp_1 _2873_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net56),
    .D(_0240_),
    .Q_N(_1106_),
    .Q(\pwm_C.accumulator[6] ));
 sg13g2_dfrbp_1 _2874_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net46),
    .D(_0241_),
    .Q_N(_1105_),
    .Q(\pwm_C.accumulator[7] ));
 sg13g2_dfrbp_1 _2875_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net326),
    .D(net489),
    .Q_N(_1104_),
    .Q(\pwm_C.accumulator[8] ));
 sg13g2_tiehi _2847__42 (.L_HI(net42));
 sg13g2_tiehi _2730__43 (.L_HI(net43));
 sg13g2_tiehi _2792__44 (.L_HI(net44));
 sg13g2_tiehi _2729__45 (.L_HI(net45));
 sg13g2_tiehi _2874__46 (.L_HI(net46));
 sg13g2_tiehi _2728__47 (.L_HI(net47));
 sg13g2_tiehi _2791__48 (.L_HI(net48));
 sg13g2_tiehi _2727__49 (.L_HI(net49));
 sg13g2_tiehi _2846__50 (.L_HI(net50));
 sg13g2_tiehi _2726__51 (.L_HI(net51));
 sg13g2_tiehi _2790__52 (.L_HI(net52));
 sg13g2_tiehi _2725__53 (.L_HI(net53));
 sg13g2_tiehi _2789__54 (.L_HI(net54));
 sg13g2_tiehi _2724__55 (.L_HI(net55));
 sg13g2_tiehi _2873__56 (.L_HI(net56));
 sg13g2_tiehi _2723__57 (.L_HI(net57));
 sg13g2_tiehi _2788__58 (.L_HI(net58));
 sg13g2_tiehi _2722__59 (.L_HI(net59));
 sg13g2_tiehi _2845__60 (.L_HI(net60));
 sg13g2_tiehi _2721__61 (.L_HI(net61));
 sg13g2_tiehi _2787__62 (.L_HI(net62));
 sg13g2_tiehi _2720__63 (.L_HI(net63));
 sg13g2_tiehi _2872__64 (.L_HI(net64));
 sg13g2_tiehi _2719__65 (.L_HI(net65));
 sg13g2_tiehi _2786__66 (.L_HI(net66));
 sg13g2_tiehi _2718__67 (.L_HI(net67));
 sg13g2_tiehi _2844__68 (.L_HI(net68));
 sg13g2_tiehi _2717__69 (.L_HI(net69));
 sg13g2_tiehi _2785__70 (.L_HI(net70));
 sg13g2_tiehi _2716__71 (.L_HI(net71));
 sg13g2_tiehi _2871__72 (.L_HI(net72));
 sg13g2_tiehi _2715__73 (.L_HI(net73));
 sg13g2_tiehi _2784__74 (.L_HI(net74));
 sg13g2_tiehi _2714__75 (.L_HI(net75));
 sg13g2_tiehi _2843__76 (.L_HI(net76));
 sg13g2_tiehi _2713__77 (.L_HI(net77));
 sg13g2_tiehi _2783__78 (.L_HI(net78));
 sg13g2_tiehi _2712__79 (.L_HI(net79));
 sg13g2_tiehi _2870__80 (.L_HI(net80));
 sg13g2_tiehi _2711__81 (.L_HI(net81));
 sg13g2_tiehi _2782__82 (.L_HI(net82));
 sg13g2_tiehi _2710__83 (.L_HI(net83));
 sg13g2_tiehi _2842__84 (.L_HI(net84));
 sg13g2_tiehi _2709__85 (.L_HI(net85));
 sg13g2_tiehi _2781__86 (.L_HI(net86));
 sg13g2_tiehi _2708__87 (.L_HI(net87));
 sg13g2_tiehi _2869__88 (.L_HI(net88));
 sg13g2_tiehi _2707__89 (.L_HI(net89));
 sg13g2_tiehi _2780__90 (.L_HI(net90));
 sg13g2_tiehi _2706__91 (.L_HI(net91));
 sg13g2_tiehi _2841__92 (.L_HI(net92));
 sg13g2_tiehi _2705__93 (.L_HI(net93));
 sg13g2_tiehi _2779__94 (.L_HI(net94));
 sg13g2_tiehi _2704__95 (.L_HI(net95));
 sg13g2_tiehi _2840__96 (.L_HI(net96));
 sg13g2_tiehi _2703__97 (.L_HI(net97));
 sg13g2_tiehi _2778__98 (.L_HI(net98));
 sg13g2_tiehi _2702__99 (.L_HI(net99));
 sg13g2_tiehi _2868__100 (.L_HI(net100));
 sg13g2_tiehi _2701__101 (.L_HI(net101));
 sg13g2_tiehi _2777__102 (.L_HI(net102));
 sg13g2_tiehi _2700__103 (.L_HI(net103));
 sg13g2_tiehi _2815__104 (.L_HI(net104));
 sg13g2_tiehi _2699__105 (.L_HI(net105));
 sg13g2_tiehi _2776__106 (.L_HI(net106));
 sg13g2_tiehi _2698__107 (.L_HI(net107));
 sg13g2_tiehi _2867__108 (.L_HI(net108));
 sg13g2_tiehi _2697__109 (.L_HI(net109));
 sg13g2_tiehi _2775__110 (.L_HI(net110));
 sg13g2_tiehi _2696__111 (.L_HI(net111));
 sg13g2_tiehi _2814__112 (.L_HI(net112));
 sg13g2_tiehi _2695__113 (.L_HI(net113));
 sg13g2_tiehi _2774__114 (.L_HI(net114));
 sg13g2_tiehi _2694__115 (.L_HI(net115));
 sg13g2_tiehi _2866__116 (.L_HI(net116));
 sg13g2_tiehi _2693__117 (.L_HI(net117));
 sg13g2_tiehi _2773__118 (.L_HI(net118));
 sg13g2_tiehi _2692__119 (.L_HI(net119));
 sg13g2_tiehi _2813__120 (.L_HI(net120));
 sg13g2_tiehi _2691__121 (.L_HI(net121));
 sg13g2_tiehi _2772__122 (.L_HI(net122));
 sg13g2_tiehi _2690__123 (.L_HI(net123));
 sg13g2_tiehi _2865__124 (.L_HI(net124));
 sg13g2_tiehi _2689__125 (.L_HI(net125));
 sg13g2_tiehi _2771__126 (.L_HI(net126));
 sg13g2_tiehi _2688__127 (.L_HI(net127));
 sg13g2_tiehi _2812__128 (.L_HI(net128));
 sg13g2_tiehi _2687__129 (.L_HI(net129));
 sg13g2_tiehi _2770__130 (.L_HI(net130));
 sg13g2_tiehi _2686__131 (.L_HI(net131));
 sg13g2_tiehi _2864__132 (.L_HI(net132));
 sg13g2_tiehi _2685__133 (.L_HI(net133));
 sg13g2_tiehi _2769__134 (.L_HI(net134));
 sg13g2_tiehi _2684__135 (.L_HI(net135));
 sg13g2_tiehi _2811__136 (.L_HI(net136));
 sg13g2_tiehi _2683__137 (.L_HI(net137));
 sg13g2_tiehi _2768__138 (.L_HI(net138));
 sg13g2_tiehi _2682__139 (.L_HI(net139));
 sg13g2_tiehi _2863__140 (.L_HI(net140));
 sg13g2_tiehi _2681__141 (.L_HI(net141));
 sg13g2_tiehi _2767__142 (.L_HI(net187));
 sg13g2_tiehi _2680__143 (.L_HI(net188));
 sg13g2_tiehi _2810__144 (.L_HI(net189));
 sg13g2_tiehi _2679__145 (.L_HI(net190));
 sg13g2_tiehi _2766__146 (.L_HI(net191));
 sg13g2_tiehi _2678__147 (.L_HI(net192));
 sg13g2_tiehi _2862__148 (.L_HI(net193));
 sg13g2_tiehi _2677__149 (.L_HI(net194));
 sg13g2_tiehi _2676__150 (.L_HI(net195));
 sg13g2_tiehi _2675__151 (.L_HI(net196));
 sg13g2_tiehi _2674__152 (.L_HI(net197));
 sg13g2_tiehi _2673__153 (.L_HI(net198));
 sg13g2_tiehi _2672__154 (.L_HI(net199));
 sg13g2_tiehi _2671__155 (.L_HI(net200));
 sg13g2_tiehi _2670__156 (.L_HI(net201));
 sg13g2_tiehi _2765__157 (.L_HI(net202));
 sg13g2_tiehi _2669__158 (.L_HI(net203));
 sg13g2_tiehi _2809__159 (.L_HI(net204));
 sg13g2_tiehi _2668__160 (.L_HI(net205));
 sg13g2_tiehi _2764__161 (.L_HI(net206));
 sg13g2_tiehi _2667__162 (.L_HI(net207));
 sg13g2_tiehi _2861__163 (.L_HI(net208));
 sg13g2_tiehi _2666__164 (.L_HI(net209));
 sg13g2_tiehi _2763__165 (.L_HI(net210));
 sg13g2_tiehi _2665__166 (.L_HI(net211));
 sg13g2_tiehi _2664__167 (.L_HI(net212));
 sg13g2_tiehi _2663__168 (.L_HI(net213));
 sg13g2_tiehi _2662__169 (.L_HI(net214));
 sg13g2_tiehi _2661__170 (.L_HI(net215));
 sg13g2_tiehi _2660__171 (.L_HI(net216));
 sg13g2_tiehi _2659__172 (.L_HI(net217));
 sg13g2_tiehi _2658__173 (.L_HI(net218));
 sg13g2_tiehi _2657__174 (.L_HI(net219));
 sg13g2_tiehi _2656__175 (.L_HI(net220));
 sg13g2_tiehi _2655__176 (.L_HI(net221));
 sg13g2_tiehi _2808__177 (.L_HI(net222));
 sg13g2_tiehi _2654__178 (.L_HI(net223));
 sg13g2_tiehi _2762__179 (.L_HI(net224));
 sg13g2_tiehi _2653__180 (.L_HI(net225));
 sg13g2_tiehi _2860__181 (.L_HI(net226));
 sg13g2_tiehi _2652__182 (.L_HI(net227));
 sg13g2_tiehi _2761__183 (.L_HI(net228));
 sg13g2_tiehi _2651__184 (.L_HI(net229));
 sg13g2_tiehi _2807__185 (.L_HI(net230));
 sg13g2_tiehi _2650__186 (.L_HI(net231));
 sg13g2_tiehi _2760__187 (.L_HI(net232));
 sg13g2_tiehi _2649__188 (.L_HI(net233));
 sg13g2_tiehi _2859__189 (.L_HI(net234));
 sg13g2_tiehi _2648__190 (.L_HI(net235));
 sg13g2_tiehi _2759__191 (.L_HI(net236));
 sg13g2_tiehi _2647__192 (.L_HI(net237));
 sg13g2_tiehi _2806__193 (.L_HI(net238));
 sg13g2_tiehi _2646__194 (.L_HI(net239));
 sg13g2_tiehi _2758__195 (.L_HI(net240));
 sg13g2_tiehi _2645__196 (.L_HI(net241));
 sg13g2_tiehi _2757__197 (.L_HI(net242));
 sg13g2_tiehi _2644__198 (.L_HI(net243));
 sg13g2_tiehi _2858__199 (.L_HI(net244));
 sg13g2_tiehi _2643__200 (.L_HI(net245));
 sg13g2_tiehi _2756__201 (.L_HI(net246));
 sg13g2_tiehi _2642__202 (.L_HI(net247));
 sg13g2_tiehi _2805__203 (.L_HI(net248));
 sg13g2_tiehi _2641__204 (.L_HI(net249));
 sg13g2_tiehi _2755__205 (.L_HI(net250));
 sg13g2_tiehi _2640__206 (.L_HI(net251));
 sg13g2_tiehi _2857__207 (.L_HI(net252));
 sg13g2_tiehi _2639__208 (.L_HI(net253));
 sg13g2_tiehi _2754__209 (.L_HI(net254));
 sg13g2_tiehi _2638__210 (.L_HI(net255));
 sg13g2_tiehi _2804__211 (.L_HI(net256));
 sg13g2_tiehi _2637__212 (.L_HI(net257));
 sg13g2_tiehi _2753__213 (.L_HI(net258));
 sg13g2_tiehi _2636__214 (.L_HI(net259));
 sg13g2_tiehi _2856__215 (.L_HI(net260));
 sg13g2_tiehi _2635__216 (.L_HI(net261));
 sg13g2_tiehi _2752__217 (.L_HI(net262));
 sg13g2_tiehi _2634__218 (.L_HI(net263));
 sg13g2_tiehi _2803__219 (.L_HI(net264));
 sg13g2_tiehi _2751__220 (.L_HI(net265));
 sg13g2_tiehi _2855__221 (.L_HI(net266));
 sg13g2_tiehi _2750__222 (.L_HI(net267));
 sg13g2_tiehi _2802__223 (.L_HI(net268));
 sg13g2_tiehi _2816__224 (.L_HI(net269));
 sg13g2_tiehi _2817__225 (.L_HI(net270));
 sg13g2_tiehi _2818__226 (.L_HI(net271));
 sg13g2_tiehi _2819__227 (.L_HI(net272));
 sg13g2_tiehi _2820__228 (.L_HI(net273));
 sg13g2_tiehi _2821__229 (.L_HI(net274));
 sg13g2_tiehi _2822__230 (.L_HI(net275));
 sg13g2_tiehi _2823__231 (.L_HI(net276));
 sg13g2_tiehi _2824__232 (.L_HI(net277));
 sg13g2_tiehi _2825__233 (.L_HI(net278));
 sg13g2_tiehi _2826__234 (.L_HI(net279));
 sg13g2_tiehi _2827__235 (.L_HI(net280));
 sg13g2_tiehi _2828__236 (.L_HI(net281));
 sg13g2_tiehi _2829__237 (.L_HI(net282));
 sg13g2_tiehi _2830__238 (.L_HI(net283));
 sg13g2_tiehi _2831__239 (.L_HI(net284));
 sg13g2_tiehi _2832__240 (.L_HI(net285));
 sg13g2_tiehi _2833__241 (.L_HI(net286));
 sg13g2_tiehi _2834__242 (.L_HI(net287));
 sg13g2_tiehi _2835__243 (.L_HI(net288));
 sg13g2_tiehi _2836__244 (.L_HI(net289));
 sg13g2_tiehi _2837__245 (.L_HI(net290));
 sg13g2_tiehi _2838__246 (.L_HI(net291));
 sg13g2_tiehi _2839__247 (.L_HI(net292));
 sg13g2_tiehi _2749__248 (.L_HI(net293));
 sg13g2_tiehi _2854__249 (.L_HI(net294));
 sg13g2_tiehi _2748__250 (.L_HI(net295));
 sg13g2_tiehi _2801__251 (.L_HI(net296));
 sg13g2_tiehi _2747__252 (.L_HI(net297));
 sg13g2_tiehi _2853__253 (.L_HI(net298));
 sg13g2_tiehi _2746__254 (.L_HI(net299));
 sg13g2_tiehi _2800__255 (.L_HI(net300));
 sg13g2_tiehi _2745__256 (.L_HI(net301));
 sg13g2_tiehi _2852__257 (.L_HI(net302));
 sg13g2_tiehi _2744__258 (.L_HI(net303));
 sg13g2_tiehi _2799__259 (.L_HI(net304));
 sg13g2_tiehi _2743__260 (.L_HI(net305));
 sg13g2_tiehi _2851__261 (.L_HI(net306));
 sg13g2_tiehi _2742__262 (.L_HI(net307));
 sg13g2_tiehi _2798__263 (.L_HI(net308));
 sg13g2_tiehi _2741__264 (.L_HI(net309));
 sg13g2_tiehi _2850__265 (.L_HI(net310));
 sg13g2_tiehi _2740__266 (.L_HI(net311));
 sg13g2_tiehi _2797__267 (.L_HI(net312));
 sg13g2_tiehi _2739__268 (.L_HI(net313));
 sg13g2_tiehi _2849__269 (.L_HI(net314));
 sg13g2_tiehi _2738__270 (.L_HI(net315));
 sg13g2_tiehi _2796__271 (.L_HI(net316));
 sg13g2_tiehi _2737__272 (.L_HI(net317));
 sg13g2_tiehi _2633__273 (.L_HI(net318));
 sg13g2_tiehi _2736__274 (.L_HI(net319));
 sg13g2_tiehi _2795__275 (.L_HI(net320));
 sg13g2_tiehi _2735__276 (.L_HI(net321));
 sg13g2_tiehi _2848__277 (.L_HI(net322));
 sg13g2_tiehi _2734__278 (.L_HI(net323));
 sg13g2_tiehi _2794__279 (.L_HI(net324));
 sg13g2_tiehi _2733__280 (.L_HI(net325));
 sg13g2_tiehi _2875__281 (.L_HI(net326));
 sg13g2_tiehi _2732__282 (.L_HI(net327));
 sg13g2_tiehi _2793__283 (.L_HI(net328));
 sg13g2_tiehi tt_um_rejunity_ay8913_284 (.L_HI(net329));
 sg13g2_tiehi tt_um_rejunity_ay8913_285 (.L_HI(net330));
 sg13g2_tiehi tt_um_rejunity_ay8913_286 (.L_HI(net331));
 sg13g2_tiehi tt_um_rejunity_ay8913_287 (.L_HI(net332));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_rejunity_ay8913_10 (.L_LO(net10));
 sg13g2_tielo tt_um_rejunity_ay8913_11 (.L_LO(net11));
 sg13g2_tielo tt_um_rejunity_ay8913_12 (.L_LO(net12));
 sg13g2_tielo tt_um_rejunity_ay8913_13 (.L_LO(net13));
 sg13g2_tielo tt_um_rejunity_ay8913_14 (.L_LO(net14));
 sg13g2_tielo tt_um_rejunity_ay8913_15 (.L_LO(net15));
 sg13g2_tielo tt_um_rejunity_ay8913_16 (.L_LO(net16));
 sg13g2_tielo _2832__17 (.L_LO(net17));
 sg13g2_tielo _2824__25 (.L_LO(net25));
 sg13g2_tielo _2816__33 (.L_LO(net33));
 sg13g2_tiehi _2731__41 (.L_HI(net41));
 sg13g2_buf_1 _3134_ (.A(\pwm_A.accumulator[8] ),
    .X(uio_out[4]));
 sg13g2_buf_1 _3135_ (.A(\pwm_B.accumulator[8] ),
    .X(uio_out[5]));
 sg13g2_buf_1 _3136_ (.A(\pwm_C.accumulator[8] ),
    .X(uio_out[6]));
 sg13g2_buf_1 _3137_ (.A(\pwm_master.accumulator[9] ),
    .X(uio_out[7]));
 sg13g2_buf_2 fanout142 (.A(_0571_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_0571_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_0433_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_0318_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_0366_),
    .X(net146));
 sg13g2_buf_1 fanout147 (.A(_0366_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_0614_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_0515_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_0270_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_1088_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_0999_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(net155),
    .X(net153));
 sg13g2_buf_1 fanout154 (.A(net155),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_0489_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(net157),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_0489_),
    .X(net157));
 sg13g2_buf_4 fanout158 (.X(net158),
    .A(net159));
 sg13g2_buf_4 fanout159 (.X(net159),
    .A(_0284_));
 sg13g2_buf_2 fanout160 (.A(_1065_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(net616),
    .X(net161));
 sg13g2_buf_4 fanout162 (.X(net162),
    .A(net164));
 sg13g2_buf_4 fanout163 (.X(net163),
    .A(_0814_));
 sg13g2_buf_2 fanout164 (.A(_0814_),
    .X(net164));
 sg13g2_buf_4 fanout165 (.X(net165),
    .A(net167));
 sg13g2_buf_4 fanout166 (.X(net166),
    .A(net167));
 sg13g2_buf_4 fanout167 (.X(net167),
    .A(_0814_));
 sg13g2_buf_4 fanout168 (.X(net168),
    .A(net1));
 sg13g2_buf_4 fanout169 (.X(net169),
    .A(net170));
 sg13g2_buf_4 fanout170 (.X(net170),
    .A(ui_in[3]));
 sg13g2_buf_4 fanout171 (.X(net171),
    .A(net172));
 sg13g2_buf_4 fanout172 (.X(net172),
    .A(ui_in[2]));
 sg13g2_buf_4 fanout173 (.X(net173),
    .A(net174));
 sg13g2_buf_4 fanout174 (.X(net174),
    .A(ui_in[1]));
 sg13g2_buf_4 fanout175 (.X(net175),
    .A(net176));
 sg13g2_buf_4 fanout176 (.X(net176),
    .A(ui_in[0]));
 sg13g2_buf_2 fanout177 (.A(net178),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(net179),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(net186),
    .X(net179));
 sg13g2_buf_4 fanout180 (.X(net180),
    .A(net186));
 sg13g2_buf_2 fanout181 (.A(net186),
    .X(net181));
 sg13g2_buf_4 fanout182 (.X(net182),
    .A(net185));
 sg13g2_buf_2 fanout183 (.A(net184),
    .X(net183));
 sg13g2_buf_4 fanout184 (.X(net184),
    .A(net185));
 sg13g2_buf_4 fanout185 (.X(net185),
    .A(net186));
 sg13g2_buf_2 fanout186 (.A(rst_n),
    .X(net186));
 sg13g2_buf_2 input1 (.A(ui_in[4]),
    .X(net1));
 sg13g2_buf_4 input2 (.X(net2),
    .A(ui_in[5]));
 sg13g2_buf_4 input3 (.X(net3),
    .A(ui_in[6]));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[7]));
 sg13g2_buf_2 input5 (.A(uio_in[0]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(uio_in[1]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[2]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[3]),
    .X(net8));
 sg13g2_tielo tt_um_rejunity_ay8913_9 (.L_LO(net9));
 sg13g2_tielo _2833__18 (.L_LO(net18));
 sg13g2_tielo _2834__19 (.L_LO(net19));
 sg13g2_tielo _2835__20 (.L_LO(net20));
 sg13g2_tielo _2836__21 (.L_LO(net21));
 sg13g2_tielo _2837__22 (.L_LO(net22));
 sg13g2_tielo _2838__23 (.L_LO(net23));
 sg13g2_tielo _2839__24 (.L_LO(net24));
 sg13g2_tielo _2825__26 (.L_LO(net26));
 sg13g2_tielo _2826__27 (.L_LO(net27));
 sg13g2_tielo _2827__28 (.L_LO(net28));
 sg13g2_tielo _2828__29 (.L_LO(net29));
 sg13g2_tielo _2829__30 (.L_LO(net30));
 sg13g2_tielo _2830__31 (.L_LO(net31));
 sg13g2_tielo _2831__32 (.L_LO(net32));
 sg13g2_tielo _2817__34 (.L_LO(net34));
 sg13g2_tielo _2818__35 (.L_LO(net35));
 sg13g2_tielo _2819__36 (.L_LO(net36));
 sg13g2_tielo _2820__37 (.L_LO(net37));
 sg13g2_tielo _2821__38 (.L_LO(net38));
 sg13g2_tielo _2822__39 (.L_LO(net39));
 sg13g2_tielo _2823__40 (.L_LO(net40));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_leaf_25_clk));
 sg13g2_inv_2 clkload4 (.A(clknet_leaf_26_clk));
 sg13g2_inv_4 clkload5 (.A(clknet_leaf_27_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_2_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_28_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_19_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_7_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_8_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_15_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0023_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0022_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0199_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0008_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0180_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold6 (.A(\amplitude_B[0] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold7 (.A(\amplitude_A[0] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold8 (.A(\amplitude_B[3] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold9 (.A(\amplitude_A[3] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold10 (.A(\amplitude_A[2] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0006_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0106_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold13 (.A(\amplitude_C[0] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold14 (.A(\amplitude_C[3] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold15 (.A(\amplitude_B[1] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold16 (.A(\amplitude_A[1] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold17 (.A(noise_disable_B),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold18 (.A(\amplitude_B[2] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold19 (.A(\register[1][1] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold20 (.A(\amplitude_C[2] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold21 (.A(noise_disable_A),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold22 (.A(envelope_attack),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0007_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0124_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold25 (.A(tone_disable_A),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold26 (.A(\amplitude_C[1] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold27 (.A(\envelope_generator.tone.counter[15] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0597_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold29 (.A(\noise_generator.period[0] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold30 (.A(\tone_C_generator.counter[11] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0453_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold32 (.A(\envelope_generator.period[5] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold33 (.A(\tone_B_generator.counter[11] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0386_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0003_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0598_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0197_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold38 (.A(\register[2][6] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold39 (.A(\envelope_generator.period[11] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold40 (.A(tone_disable_C),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0004_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0154_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold43 (.A(\noise_generator.tone.counter[1] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0483_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0150_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold46 (.A(\envelope_generator.period[0] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold47 (.A(\register[2][4] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold48 (.A(\register[0][3] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold49 (.A(\envelope_generator.period[9] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0005_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0093_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold52 (.A(\tone_A_generator.counter[1] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0321_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold54 (.A(\register[1][2] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold55 (.A(\envelope_generator.signal_edge.signal ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0148_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold57 (.A(\register[3][2] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold58 (.A(\register[4][1] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold59 (.A(noise_disable_C),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold60 (.A(\envelope_generator.period[12] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold61 (.A(\envelope_generator.period[7] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold62 (.A(envelope_alternate),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold63 (.A(\register[3][1] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold64 (.A(tone_disable_B),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold65 (.A(\envelope_generator.tone.counter[13] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0595_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0194_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold68 (.A(\register[2][2] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold69 (.A(\noise_generator.period[4] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold70 (.A(\envelope_generator.period[2] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold71 (.A(\envelope_generator.period[1] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold72 (.A(\register[2][3] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold73 (.A(\noise_generator.tone.counter[4] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0487_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold75 (.A(\envelope_generator.period[13] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold76 (.A(\register[4][0] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold77 (.A(\register[3][0] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold78 (.A(\register[2][7] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold79 (.A(\register[2][0] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold80 (.A(\envelope_generator.period[15] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold81 (.A(\tone_A_generator.counter[11] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0337_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold83 (.A(\noise_generator.period[2] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold84 (.A(\noise_generator.lfsr[9] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0163_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold86 (.A(\clk_counter[2] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold87 (.A(_1072_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0063_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold89 (.A(\pwm_C.accumulator[0] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold90 (.A(\envelope_generator.period[4] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold91 (.A(\noise_generator.period[1] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold92 (.A(\register[2][1] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold93 (.A(\register[1][3] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold94 (.A(\envelope_generator.period[3] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold95 (.A(\register[4][2] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold96 (.A(\pwm_A.accumulator[0] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold97 (.A(\envelope_generator.tone.counter[1] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0573_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0182_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold100 (.A(\noise_generator.lfsr[15] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0169_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold102 (.A(\noise_generator.lfsr[1] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0155_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold104 (.A(\register[4][3] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold105 (.A(\noise_generator.period[3] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold106 (.A(\register[2][5] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold107 (.A(\envelope_generator.period[8] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold108 (.A(\register[5][2] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold109 (.A(\register[5][0] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold110 (.A(\tone_B_generator.counter[1] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0369_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0108_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold113 (.A(\tone_B_generator.counter[9] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0384_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold115 (.A(\register[3][3] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold116 (.A(active),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold117 (.A(\noise_generator.lfsr[11] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0165_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold119 (.A(\clk_counter[6] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0067_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold121 (.A(\noise_generator.lfsr[13] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0167_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold123 (.A(\register[0][2] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold124 (.A(\noise_generator.lfsr[8] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0162_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold126 (.A(\register[0][6] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold127 (.A(\noise_generator.lfsr[7] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0161_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold129 (.A(\register[5][1] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold130 (.A(\noise_generator.lfsr[4] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0158_),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold132 (.A(\register[0][1] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold133 (.A(\noise_generator.lfsr[12] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold134 (.A(\envelope_generator.period[10] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold135 (.A(\register[0][4] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold136 (.A(\register[1][0] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold137 (.A(\noise_generator.lfsr[16] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0170_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold139 (.A(\noise_generator.lfsr[2] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold140 (.A(\noise_generator.signal_edge.signal ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold141 (.A(\noise_generator.lfsr[6] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0160_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold143 (.A(\register[4][6] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold144 (.A(envelope_continue),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold145 (.A(\envelope_generator.period[14] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold146 (.A(\register[0][0] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold147 (.A(\envelope_generator.period[6] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold148 (.A(\noise_generator.lfsr[10] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold149 (.A(\pwm_B.accumulator[0] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold150 (.A(\tone_C_generator.counter[1] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0436_),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0126_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold153 (.A(\envelope_generator.stop ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0600_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0198_),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold156 (.A(\pwm_C.accumulator[7] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0242_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold158 (.A(\pwm_A.accumulator[7] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold159 (.A(\envelope_generator.tone.counter[6] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0583_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0187_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold162 (.A(\register[5][3] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold163 (.A(\noise_generator.lfsr[14] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold164 (.A(\envelope_generator.envelope_counter[3] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0202_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold166 (.A(\noise_generator.lfsr[3] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0493_),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0157_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold169 (.A(\tone_A_generator.counter[9] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0335_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold171 (.A(\noise_generator.lfsr[5] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold172 (.A(\noise_generator.tone.counter[2] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0485_),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold174 (.A(\envelope_generator.hold ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold175 (.A(\register[4][5] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold176 (.A(\register[0][5] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold177 (.A(\tone_B_generator.counter[6] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0379_),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold179 (.A(\tone_B_generator.counter[4] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0375_),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold181 (.A(\envelope_generator.envelope_counter[1] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0603_),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0200_),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold184 (.A(\noise_generator.tone.counter[3] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold185 (.A(\pwm_B.accumulator[7] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold186 (.A(\tone_B_generator.counter[2] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0371_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold188 (.A(\register[4][7] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold189 (.A(\register[0][7] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold190 (.A(\register[4][4] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold191 (.A(\envelope_generator.tone.counter[10] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0589_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0191_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold194 (.A(\tone_B_generator.counter[3] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold195 (.A(\clk_counter[4] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold196 (.A(_1077_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold197 (.A(\tone_C_generator.counter[4] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0442_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold199 (.A(\noise_generator.signal_edge.previous_signal_state_0 ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0171_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold201 (.A(\tone_B_generator.counter[5] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold202 (.A(\envelope_generator.tone.counter[8] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0586_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold204 (.A(\tone_C_generator.counter[9] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0451_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold206 (.A(\tone_A_generator.counter[4] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0327_),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold208 (.A(\tone_C_generator.counter[2] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0438_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold210 (.A(\envelope_generator.tone.counter[7] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0585_),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold212 (.A(\envelope_generator.tone.counter[4] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0579_),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0185_),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold215 (.A(\tone_B_generator.counter[7] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold216 (.A(\tone_A_generator.counter[10] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold217 (.A(\clk_counter[0] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold218 (.A(_1071_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold219 (.A(\envelope_generator.tone.counter[14] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0596_),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold221 (.A(\envelope_generator.tone.counter[2] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0576_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold223 (.A(\envelope_generator.tone.counter[11] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0591_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold225 (.A(\tone_A_generator.counter[5] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold226 (.A(\tone_A_generator.counter[3] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0325_),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold228 (.A(\tone_C_generator.counter[5] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold229 (.A(\tone_C_generator.counter[8] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0449_),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold231 (.A(restart_envelope),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0606_),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold233 (.A(\tone_A_generator.counter[2] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0323_),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold235 (.A(\clk_counter[5] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold236 (.A(\pwm_master.accumulator[8] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0055_),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold238 (.A(\tone_B_generator.counter[10] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0385_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold240 (.A(\pwm_master.accumulator[0] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0047_),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold242 (.A(\tone_C_generator.counter[10] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold243 (.A(\envelope_generator.tone.counter[5] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0581_),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold245 (.A(\envelope_generator.tone.counter[12] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold246 (.A(\noise_generator.tone.counter[0] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold247 (.A(\tone_C_generator.counter[3] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold248 (.A(\envelope_generator.tone.counter[9] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold249 (.A(envelope_B),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold250 (.A(\tone_B_generator.counter[8] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold251 (.A(\pwm_C.accumulator[3] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0237_),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold253 (.A(\pwm_B.accumulator[3] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0228_),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold255 (.A(\pwm_A.accumulator[3] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0219_),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold257 (.A(envelope_C),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold258 (.A(\envelope_generator.tone.counter[0] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold259 (.A(\tone_A_generator.counter[8] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0333_),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold261 (.A(\clk_counter[3] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold262 (.A(_1076_),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold263 (.A(\latched_register[2] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold264 (.A(\latched_register[0] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold265 (.A(\tone_B_generator.counter[0] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold266 (.A(\latched_register[3] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold267 (.A(\latched_register[1] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold268 (.A(\tone_C_generator.counter[0] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold269 (.A(\tone_C_generator.counter[6] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold270 (.A(\tone_A_generator.counter[0] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold271 (.A(\pwm_B.accumulator[5] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold272 (.A(_0230_),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold273 (.A(\pwm_master.accumulator[3] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0049_),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold275 (.A(\pwm_C.accumulator[5] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0239_),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold277 (.A(\pwm_A.accumulator[1] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold278 (.A(\tone_C_generator.counter[7] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold279 (.A(\tone_A_generator.counter[7] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0332_),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold281 (.A(\pwm_C.accumulator[1] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold282 (.A(\pwm_A.accumulator[5] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0221_),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold284 (.A(envelope_A),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold285 (.A(\pwm_B.accumulator[1] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold286 (.A(\pwm_C.accumulator[6] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold287 (.A(\envelope_generator.tone.counter[3] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold288 (.A(\pwm_master.accumulator[4] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold289 (.A(\tone_A_generator.counter[6] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold290 (.A(\pwm_master.accumulator[7] ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0053_),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold292 (.A(\pwm_C.accumulator[2] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold293 (.A(\pwm_A.accumulator[4] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold294 (.A(\pwm_A.accumulator[6] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold295 (.A(\pwm_A.accumulator[2] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold296 (.A(\pwm_master.accumulator[2] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold297 (.A(\pwm_master.accumulator[8] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold298 (.A(\pwm_B.accumulator[2] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold299 (.A(_0665_),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0227_),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold301 (.A(\pwm_B.accumulator[6] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold302 (.A(\pwm_master.accumulator[5] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold303 (.A(\pwm_master.accumulator[6] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold304 (.A(\tone_B_generator.counter[8] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold305 (.A(\tone_A_generator.counter[8] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold306 (.A(\latched_register[2] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold307 (.A(_1088_),
    .X(net639));
 sg13g2_antennanp ANTENNA_1 (.A(rst_n));
 sg13g2_antennanp ANTENNA_2 (.A(rst_n));
 sg13g2_antennanp ANTENNA_3 (.A(rst_n));
 sg13g2_antennanp ANTENNA_4 (.A(rst_n));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_4 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_274 ();
 sg13g2_fill_1 FILLER_3_281 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_fill_2 FILLER_4_264 ();
 sg13g2_decap_8 FILLER_4_311 ();
 sg13g2_decap_8 FILLER_4_318 ();
 sg13g2_decap_8 FILLER_4_325 ();
 sg13g2_decap_8 FILLER_4_332 ();
 sg13g2_decap_8 FILLER_4_339 ();
 sg13g2_decap_8 FILLER_4_346 ();
 sg13g2_decap_8 FILLER_4_353 ();
 sg13g2_decap_8 FILLER_4_360 ();
 sg13g2_decap_8 FILLER_4_367 ();
 sg13g2_decap_8 FILLER_4_374 ();
 sg13g2_decap_8 FILLER_4_381 ();
 sg13g2_decap_8 FILLER_4_388 ();
 sg13g2_decap_8 FILLER_4_395 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_fill_2 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_318 ();
 sg13g2_decap_8 FILLER_5_325 ();
 sg13g2_decap_8 FILLER_5_332 ();
 sg13g2_decap_8 FILLER_5_339 ();
 sg13g2_decap_8 FILLER_5_346 ();
 sg13g2_decap_8 FILLER_5_353 ();
 sg13g2_decap_8 FILLER_5_360 ();
 sg13g2_decap_8 FILLER_5_367 ();
 sg13g2_decap_8 FILLER_5_374 ();
 sg13g2_decap_8 FILLER_5_381 ();
 sg13g2_decap_8 FILLER_5_388 ();
 sg13g2_decap_8 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_fill_2 FILLER_6_224 ();
 sg13g2_fill_2 FILLER_6_275 ();
 sg13g2_fill_1 FILLER_6_277 ();
 sg13g2_decap_8 FILLER_6_326 ();
 sg13g2_decap_8 FILLER_6_333 ();
 sg13g2_decap_8 FILLER_6_340 ();
 sg13g2_decap_8 FILLER_6_347 ();
 sg13g2_decap_8 FILLER_6_354 ();
 sg13g2_decap_8 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_decap_8 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_396 ();
 sg13g2_decap_4 FILLER_6_403 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_fill_1 FILLER_7_231 ();
 sg13g2_fill_2 FILLER_7_276 ();
 sg13g2_fill_1 FILLER_7_278 ();
 sg13g2_decap_8 FILLER_7_320 ();
 sg13g2_decap_8 FILLER_7_327 ();
 sg13g2_decap_8 FILLER_7_334 ();
 sg13g2_decap_8 FILLER_7_341 ();
 sg13g2_decap_8 FILLER_7_348 ();
 sg13g2_decap_8 FILLER_7_355 ();
 sg13g2_decap_8 FILLER_7_362 ();
 sg13g2_decap_8 FILLER_7_369 ();
 sg13g2_decap_8 FILLER_7_376 ();
 sg13g2_decap_8 FILLER_7_383 ();
 sg13g2_decap_8 FILLER_7_390 ();
 sg13g2_decap_8 FILLER_7_397 ();
 sg13g2_decap_4 FILLER_7_404 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_fill_2 FILLER_8_231 ();
 sg13g2_fill_1 FILLER_8_233 ();
 sg13g2_fill_1 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_316 ();
 sg13g2_decap_8 FILLER_8_323 ();
 sg13g2_fill_1 FILLER_8_330 ();
 sg13g2_decap_8 FILLER_8_335 ();
 sg13g2_decap_8 FILLER_8_342 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_356 ();
 sg13g2_decap_8 FILLER_8_363 ();
 sg13g2_decap_8 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_fill_2 FILLER_9_231 ();
 sg13g2_decap_4 FILLER_9_314 ();
 sg13g2_decap_8 FILLER_9_374 ();
 sg13g2_decap_8 FILLER_9_381 ();
 sg13g2_decap_8 FILLER_9_388 ();
 sg13g2_decap_8 FILLER_9_395 ();
 sg13g2_decap_8 FILLER_9_402 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_fill_2 FILLER_10_300 ();
 sg13g2_decap_8 FILLER_10_380 ();
 sg13g2_decap_8 FILLER_10_387 ();
 sg13g2_decap_8 FILLER_10_394 ();
 sg13g2_decap_8 FILLER_10_401 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_fill_2 FILLER_11_224 ();
 sg13g2_fill_2 FILLER_11_257 ();
 sg13g2_fill_2 FILLER_11_268 ();
 sg13g2_decap_8 FILLER_11_288 ();
 sg13g2_decap_4 FILLER_11_295 ();
 sg13g2_fill_1 FILLER_11_299 ();
 sg13g2_decap_8 FILLER_11_307 ();
 sg13g2_fill_2 FILLER_11_314 ();
 sg13g2_fill_1 FILLER_11_316 ();
 sg13g2_fill_2 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_fill_2 FILLER_12_231 ();
 sg13g2_fill_1 FILLER_12_245 ();
 sg13g2_fill_2 FILLER_12_264 ();
 sg13g2_decap_4 FILLER_12_316 ();
 sg13g2_fill_2 FILLER_12_320 ();
 sg13g2_fill_1 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_384 ();
 sg13g2_decap_8 FILLER_12_391 ();
 sg13g2_decap_8 FILLER_12_398 ();
 sg13g2_decap_4 FILLER_12_405 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_4 FILLER_13_245 ();
 sg13g2_fill_2 FILLER_13_249 ();
 sg13g2_fill_2 FILLER_13_254 ();
 sg13g2_fill_1 FILLER_13_256 ();
 sg13g2_fill_1 FILLER_13_283 ();
 sg13g2_fill_2 FILLER_13_310 ();
 sg13g2_fill_2 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_321 ();
 sg13g2_fill_2 FILLER_13_328 ();
 sg13g2_fill_1 FILLER_13_334 ();
 sg13g2_fill_2 FILLER_13_347 ();
 sg13g2_fill_1 FILLER_13_354 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_4 FILLER_14_238 ();
 sg13g2_fill_2 FILLER_14_242 ();
 sg13g2_fill_1 FILLER_14_257 ();
 sg13g2_fill_2 FILLER_14_266 ();
 sg13g2_fill_1 FILLER_14_291 ();
 sg13g2_fill_1 FILLER_14_305 ();
 sg13g2_fill_2 FILLER_14_335 ();
 sg13g2_fill_2 FILLER_14_352 ();
 sg13g2_fill_1 FILLER_14_361 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_4 FILLER_15_224 ();
 sg13g2_fill_1 FILLER_15_273 ();
 sg13g2_fill_1 FILLER_15_279 ();
 sg13g2_fill_2 FILLER_15_286 ();
 sg13g2_fill_2 FILLER_15_334 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_4 FILLER_16_217 ();
 sg13g2_fill_2 FILLER_16_221 ();
 sg13g2_fill_1 FILLER_16_287 ();
 sg13g2_fill_2 FILLER_16_291 ();
 sg13g2_decap_4 FILLER_16_300 ();
 sg13g2_fill_1 FILLER_16_304 ();
 sg13g2_decap_4 FILLER_16_361 ();
 sg13g2_fill_2 FILLER_16_365 ();
 sg13g2_decap_8 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_4 FILLER_17_224 ();
 sg13g2_fill_2 FILLER_17_228 ();
 sg13g2_fill_2 FILLER_17_266 ();
 sg13g2_fill_1 FILLER_17_268 ();
 sg13g2_decap_8 FILLER_17_275 ();
 sg13g2_decap_8 FILLER_17_282 ();
 sg13g2_decap_8 FILLER_17_289 ();
 sg13g2_fill_1 FILLER_17_296 ();
 sg13g2_decap_8 FILLER_17_300 ();
 sg13g2_fill_1 FILLER_17_307 ();
 sg13g2_decap_4 FILLER_17_356 ();
 sg13g2_decap_8 FILLER_17_377 ();
 sg13g2_decap_8 FILLER_17_384 ();
 sg13g2_decap_8 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_17_398 ();
 sg13g2_decap_4 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_fill_1 FILLER_18_224 ();
 sg13g2_fill_2 FILLER_18_263 ();
 sg13g2_fill_1 FILLER_18_265 ();
 sg13g2_fill_2 FILLER_18_320 ();
 sg13g2_fill_1 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_fill_2 FILLER_18_343 ();
 sg13g2_fill_1 FILLER_18_368 ();
 sg13g2_decap_8 FILLER_18_384 ();
 sg13g2_decap_8 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_4 FILLER_19_238 ();
 sg13g2_fill_1 FILLER_19_242 ();
 sg13g2_decap_4 FILLER_19_248 ();
 sg13g2_fill_1 FILLER_19_284 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_fill_2 FILLER_20_224 ();
 sg13g2_fill_2 FILLER_20_286 ();
 sg13g2_fill_2 FILLER_20_365 ();
 sg13g2_fill_2 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_395 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_4 FILLER_21_147 ();
 sg13g2_fill_2 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_159 ();
 sg13g2_decap_8 FILLER_21_166 ();
 sg13g2_decap_8 FILLER_21_173 ();
 sg13g2_decap_8 FILLER_21_180 ();
 sg13g2_decap_8 FILLER_21_187 ();
 sg13g2_decap_8 FILLER_21_194 ();
 sg13g2_decap_8 FILLER_21_201 ();
 sg13g2_decap_8 FILLER_21_208 ();
 sg13g2_decap_4 FILLER_21_215 ();
 sg13g2_fill_2 FILLER_21_245 ();
 sg13g2_fill_1 FILLER_21_247 ();
 sg13g2_decap_4 FILLER_21_274 ();
 sg13g2_fill_2 FILLER_21_278 ();
 sg13g2_fill_2 FILLER_21_284 ();
 sg13g2_fill_1 FILLER_21_286 ();
 sg13g2_fill_2 FILLER_21_293 ();
 sg13g2_fill_1 FILLER_21_295 ();
 sg13g2_fill_1 FILLER_21_345 ();
 sg13g2_fill_2 FILLER_21_354 ();
 sg13g2_fill_1 FILLER_21_365 ();
 sg13g2_fill_1 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_fill_2 FILLER_22_140 ();
 sg13g2_fill_1 FILLER_22_142 ();
 sg13g2_fill_2 FILLER_22_157 ();
 sg13g2_decap_8 FILLER_22_172 ();
 sg13g2_decap_8 FILLER_22_179 ();
 sg13g2_decap_8 FILLER_22_186 ();
 sg13g2_decap_8 FILLER_22_193 ();
 sg13g2_decap_8 FILLER_22_200 ();
 sg13g2_decap_8 FILLER_22_207 ();
 sg13g2_fill_2 FILLER_22_214 ();
 sg13g2_fill_1 FILLER_22_268 ();
 sg13g2_fill_2 FILLER_22_273 ();
 sg13g2_decap_4 FILLER_22_300 ();
 sg13g2_fill_2 FILLER_22_304 ();
 sg13g2_decap_8 FILLER_22_309 ();
 sg13g2_decap_8 FILLER_22_316 ();
 sg13g2_fill_2 FILLER_22_323 ();
 sg13g2_fill_2 FILLER_22_333 ();
 sg13g2_fill_1 FILLER_22_335 ();
 sg13g2_fill_2 FILLER_22_351 ();
 sg13g2_decap_8 FILLER_22_387 ();
 sg13g2_decap_8 FILLER_22_394 ();
 sg13g2_decap_8 FILLER_22_401 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_fill_1 FILLER_23_137 ();
 sg13g2_decap_8 FILLER_23_183 ();
 sg13g2_decap_8 FILLER_23_190 ();
 sg13g2_decap_8 FILLER_23_197 ();
 sg13g2_decap_4 FILLER_23_204 ();
 sg13g2_fill_1 FILLER_23_208 ();
 sg13g2_fill_1 FILLER_23_330 ();
 sg13g2_decap_8 FILLER_23_397 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_4 FILLER_24_119 ();
 sg13g2_fill_1 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_181 ();
 sg13g2_decap_8 FILLER_24_188 ();
 sg13g2_decap_8 FILLER_24_195 ();
 sg13g2_decap_8 FILLER_24_202 ();
 sg13g2_decap_8 FILLER_24_209 ();
 sg13g2_fill_1 FILLER_24_225 ();
 sg13g2_fill_1 FILLER_24_250 ();
 sg13g2_decap_8 FILLER_24_278 ();
 sg13g2_fill_2 FILLER_24_285 ();
 sg13g2_fill_2 FILLER_24_290 ();
 sg13g2_fill_1 FILLER_24_292 ();
 sg13g2_fill_2 FILLER_24_299 ();
 sg13g2_fill_1 FILLER_24_301 ();
 sg13g2_fill_2 FILLER_24_337 ();
 sg13g2_fill_2 FILLER_24_365 ();
 sg13g2_decap_8 FILLER_24_393 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_fill_2 FILLER_25_119 ();
 sg13g2_fill_1 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_181 ();
 sg13g2_decap_8 FILLER_25_188 ();
 sg13g2_decap_8 FILLER_25_195 ();
 sg13g2_decap_8 FILLER_25_202 ();
 sg13g2_fill_1 FILLER_25_209 ();
 sg13g2_decap_4 FILLER_25_276 ();
 sg13g2_decap_8 FILLER_25_389 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_decap_4 FILLER_25_403 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_4 FILLER_26_112 ();
 sg13g2_fill_1 FILLER_26_145 ();
 sg13g2_fill_2 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_190 ();
 sg13g2_decap_8 FILLER_26_197 ();
 sg13g2_decap_8 FILLER_26_204 ();
 sg13g2_decap_8 FILLER_26_211 ();
 sg13g2_fill_2 FILLER_26_278 ();
 sg13g2_fill_2 FILLER_26_289 ();
 sg13g2_fill_2 FILLER_26_295 ();
 sg13g2_fill_2 FILLER_26_314 ();
 sg13g2_fill_2 FILLER_26_362 ();
 sg13g2_fill_2 FILLER_26_373 ();
 sg13g2_fill_1 FILLER_26_375 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_fill_2 FILLER_27_119 ();
 sg13g2_fill_1 FILLER_27_187 ();
 sg13g2_decap_8 FILLER_27_197 ();
 sg13g2_decap_8 FILLER_27_204 ();
 sg13g2_decap_4 FILLER_27_211 ();
 sg13g2_decap_4 FILLER_27_219 ();
 sg13g2_fill_1 FILLER_27_223 ();
 sg13g2_fill_1 FILLER_27_264 ();
 sg13g2_fill_1 FILLER_27_311 ();
 sg13g2_fill_1 FILLER_27_322 ();
 sg13g2_fill_2 FILLER_27_339 ();
 sg13g2_fill_2 FILLER_27_347 ();
 sg13g2_decap_8 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_27_396 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_fill_1 FILLER_28_119 ();
 sg13g2_fill_1 FILLER_28_155 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_4 FILLER_28_203 ();
 sg13g2_fill_2 FILLER_28_207 ();
 sg13g2_fill_1 FILLER_28_230 ();
 sg13g2_fill_2 FILLER_28_236 ();
 sg13g2_fill_1 FILLER_28_262 ();
 sg13g2_fill_2 FILLER_28_334 ();
 sg13g2_fill_2 FILLER_28_345 ();
 sg13g2_decap_8 FILLER_28_373 ();
 sg13g2_decap_8 FILLER_28_380 ();
 sg13g2_decap_8 FILLER_28_387 ();
 sg13g2_decap_8 FILLER_28_394 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_fill_2 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_188 ();
 sg13g2_decap_8 FILLER_29_195 ();
 sg13g2_fill_2 FILLER_29_202 ();
 sg13g2_fill_1 FILLER_29_204 ();
 sg13g2_fill_2 FILLER_29_275 ();
 sg13g2_decap_8 FILLER_29_384 ();
 sg13g2_decap_8 FILLER_29_391 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_fill_2 FILLER_30_133 ();
 sg13g2_fill_1 FILLER_30_135 ();
 sg13g2_fill_1 FILLER_30_174 ();
 sg13g2_fill_1 FILLER_30_193 ();
 sg13g2_fill_2 FILLER_30_206 ();
 sg13g2_fill_1 FILLER_30_356 ();
 sg13g2_decap_8 FILLER_30_383 ();
 sg13g2_decap_8 FILLER_30_390 ();
 sg13g2_decap_8 FILLER_30_397 ();
 sg13g2_decap_4 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_fill_2 FILLER_31_177 ();
 sg13g2_fill_1 FILLER_31_179 ();
 sg13g2_fill_1 FILLER_31_185 ();
 sg13g2_fill_2 FILLER_31_225 ();
 sg13g2_fill_1 FILLER_31_227 ();
 sg13g2_fill_2 FILLER_31_260 ();
 sg13g2_fill_2 FILLER_31_266 ();
 sg13g2_decap_8 FILLER_31_282 ();
 sg13g2_fill_2 FILLER_31_289 ();
 sg13g2_fill_1 FILLER_31_291 ();
 sg13g2_decap_8 FILLER_31_297 ();
 sg13g2_fill_2 FILLER_31_317 ();
 sg13g2_fill_2 FILLER_31_330 ();
 sg13g2_fill_1 FILLER_31_332 ();
 sg13g2_fill_1 FILLER_31_347 ();
 sg13g2_decap_8 FILLER_31_374 ();
 sg13g2_decap_8 FILLER_31_381 ();
 sg13g2_decap_8 FILLER_31_388 ();
 sg13g2_decap_8 FILLER_31_395 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_fill_2 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_142 ();
 sg13g2_fill_1 FILLER_32_171 ();
 sg13g2_decap_4 FILLER_32_233 ();
 sg13g2_fill_1 FILLER_32_237 ();
 sg13g2_fill_2 FILLER_32_289 ();
 sg13g2_fill_2 FILLER_32_299 ();
 sg13g2_decap_8 FILLER_32_307 ();
 sg13g2_decap_8 FILLER_32_314 ();
 sg13g2_decap_8 FILLER_32_321 ();
 sg13g2_fill_2 FILLER_32_328 ();
 sg13g2_decap_8 FILLER_32_338 ();
 sg13g2_decap_8 FILLER_32_345 ();
 sg13g2_decap_4 FILLER_32_352 ();
 sg13g2_decap_4 FILLER_32_362 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_4 FILLER_33_133 ();
 sg13g2_fill_1 FILLER_33_194 ();
 sg13g2_fill_2 FILLER_33_203 ();
 sg13g2_fill_1 FILLER_33_205 ();
 sg13g2_decap_8 FILLER_33_225 ();
 sg13g2_fill_1 FILLER_33_232 ();
 sg13g2_decap_8 FILLER_33_237 ();
 sg13g2_fill_1 FILLER_33_249 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_decap_4 FILLER_33_266 ();
 sg13g2_fill_1 FILLER_33_274 ();
 sg13g2_decap_4 FILLER_33_280 ();
 sg13g2_fill_2 FILLER_33_293 ();
 sg13g2_fill_1 FILLER_33_295 ();
 sg13g2_decap_4 FILLER_33_322 ();
 sg13g2_fill_1 FILLER_33_326 ();
 sg13g2_decap_8 FILLER_33_395 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_fill_2 FILLER_34_126 ();
 sg13g2_fill_1 FILLER_34_154 ();
 sg13g2_fill_2 FILLER_34_233 ();
 sg13g2_fill_2 FILLER_34_244 ();
 sg13g2_fill_1 FILLER_34_246 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_4 FILLER_34_266 ();
 sg13g2_fill_1 FILLER_34_270 ();
 sg13g2_fill_1 FILLER_34_279 ();
 sg13g2_fill_2 FILLER_34_322 ();
 sg13g2_fill_1 FILLER_34_363 ();
 sg13g2_fill_2 FILLER_34_381 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_fill_2 FILLER_35_126 ();
 sg13g2_fill_1 FILLER_35_163 ();
 sg13g2_fill_1 FILLER_35_209 ();
 sg13g2_fill_1 FILLER_35_241 ();
 sg13g2_decap_4 FILLER_35_294 ();
 sg13g2_fill_1 FILLER_35_298 ();
 sg13g2_fill_2 FILLER_35_369 ();
 sg13g2_decap_8 FILLER_35_396 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_fill_2 FILLER_36_126 ();
 sg13g2_fill_1 FILLER_36_128 ();
 sg13g2_fill_1 FILLER_36_162 ();
 sg13g2_fill_1 FILLER_36_201 ();
 sg13g2_fill_2 FILLER_36_216 ();
 sg13g2_fill_1 FILLER_36_240 ();
 sg13g2_fill_1 FILLER_36_275 ();
 sg13g2_fill_2 FILLER_36_314 ();
 sg13g2_fill_2 FILLER_36_325 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_4 FILLER_37_126 ();
 sg13g2_fill_1 FILLER_37_130 ();
 sg13g2_fill_1 FILLER_37_163 ();
 sg13g2_fill_2 FILLER_37_177 ();
 sg13g2_fill_2 FILLER_37_192 ();
 sg13g2_decap_8 FILLER_37_198 ();
 sg13g2_decap_8 FILLER_37_205 ();
 sg13g2_fill_2 FILLER_37_212 ();
 sg13g2_fill_1 FILLER_37_214 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_fill_2 FILLER_37_231 ();
 sg13g2_fill_1 FILLER_37_233 ();
 sg13g2_fill_1 FILLER_37_246 ();
 sg13g2_fill_2 FILLER_37_284 ();
 sg13g2_decap_4 FILLER_37_290 ();
 sg13g2_fill_1 FILLER_37_300 ();
 sg13g2_fill_2 FILLER_37_311 ();
 sg13g2_fill_1 FILLER_37_313 ();
 sg13g2_decap_4 FILLER_37_320 ();
 sg13g2_fill_2 FILLER_37_324 ();
 sg13g2_fill_2 FILLER_37_332 ();
 sg13g2_fill_1 FILLER_37_334 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_4 FILLER_38_126 ();
 sg13g2_fill_1 FILLER_38_130 ();
 sg13g2_fill_1 FILLER_38_184 ();
 sg13g2_fill_2 FILLER_38_197 ();
 sg13g2_fill_1 FILLER_38_199 ();
 sg13g2_decap_8 FILLER_38_204 ();
 sg13g2_decap_8 FILLER_38_211 ();
 sg13g2_decap_8 FILLER_38_218 ();
 sg13g2_fill_2 FILLER_38_225 ();
 sg13g2_fill_2 FILLER_38_272 ();
 sg13g2_fill_1 FILLER_38_274 ();
 sg13g2_decap_8 FILLER_38_354 ();
 sg13g2_decap_8 FILLER_38_361 ();
 sg13g2_decap_8 FILLER_38_368 ();
 sg13g2_fill_2 FILLER_38_375 ();
 sg13g2_fill_2 FILLER_38_385 ();
 sg13g2_fill_1 FILLER_38_387 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_fill_2 FILLER_39_150 ();
 sg13g2_decap_8 FILLER_39_245 ();
 sg13g2_fill_2 FILLER_39_252 ();
 sg13g2_fill_1 FILLER_39_254 ();
 sg13g2_decap_4 FILLER_39_264 ();
 sg13g2_fill_2 FILLER_39_338 ();
 sg13g2_decap_8 FILLER_39_353 ();
 sg13g2_decap_4 FILLER_39_360 ();
 sg13g2_fill_1 FILLER_39_364 ();
 sg13g2_fill_1 FILLER_39_375 ();
 sg13g2_decap_8 FILLER_39_401 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_fill_2 FILLER_40_147 ();
 sg13g2_fill_1 FILLER_40_149 ();
 sg13g2_fill_1 FILLER_40_207 ();
 sg13g2_fill_2 FILLER_40_224 ();
 sg13g2_fill_2 FILLER_40_252 ();
 sg13g2_fill_2 FILLER_40_287 ();
 sg13g2_fill_1 FILLER_40_298 ();
 sg13g2_fill_1 FILLER_40_325 ();
 sg13g2_fill_2 FILLER_40_335 ();
 sg13g2_fill_1 FILLER_40_377 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_165 ();
 sg13g2_decap_4 FILLER_41_172 ();
 sg13g2_fill_1 FILLER_41_216 ();
 sg13g2_fill_1 FILLER_41_245 ();
 sg13g2_fill_2 FILLER_41_295 ();
 sg13g2_fill_1 FILLER_41_318 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_8 FILLER_42_154 ();
 sg13g2_fill_2 FILLER_42_161 ();
 sg13g2_fill_1 FILLER_42_163 ();
 sg13g2_decap_8 FILLER_42_167 ();
 sg13g2_decap_8 FILLER_42_174 ();
 sg13g2_decap_4 FILLER_42_181 ();
 sg13g2_fill_2 FILLER_42_190 ();
 sg13g2_fill_2 FILLER_42_204 ();
 sg13g2_fill_1 FILLER_42_206 ();
 sg13g2_decap_4 FILLER_42_211 ();
 sg13g2_fill_2 FILLER_42_215 ();
 sg13g2_decap_8 FILLER_42_221 ();
 sg13g2_decap_4 FILLER_42_228 ();
 sg13g2_fill_2 FILLER_42_232 ();
 sg13g2_decap_8 FILLER_42_239 ();
 sg13g2_decap_4 FILLER_42_246 ();
 sg13g2_fill_1 FILLER_42_250 ();
 sg13g2_fill_1 FILLER_42_271 ();
 sg13g2_fill_1 FILLER_42_313 ();
 sg13g2_fill_1 FILLER_42_337 ();
 sg13g2_fill_1 FILLER_42_344 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_decap_4 FILLER_43_154 ();
 sg13g2_fill_2 FILLER_43_158 ();
 sg13g2_decap_8 FILLER_43_184 ();
 sg13g2_decap_8 FILLER_43_191 ();
 sg13g2_decap_8 FILLER_43_198 ();
 sg13g2_decap_8 FILLER_43_205 ();
 sg13g2_decap_8 FILLER_43_216 ();
 sg13g2_fill_2 FILLER_43_223 ();
 sg13g2_decap_8 FILLER_43_260 ();
 sg13g2_fill_2 FILLER_43_267 ();
 sg13g2_fill_1 FILLER_43_305 ();
 sg13g2_fill_2 FILLER_43_366 ();
 sg13g2_fill_1 FILLER_43_368 ();
 sg13g2_fill_2 FILLER_43_373 ();
 sg13g2_fill_1 FILLER_43_379 ();
 sg13g2_fill_1 FILLER_43_393 ();
 sg13g2_fill_2 FILLER_43_398 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_decap_8 FILLER_44_140 ();
 sg13g2_decap_8 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_decap_8 FILLER_44_161 ();
 sg13g2_decap_8 FILLER_44_168 ();
 sg13g2_decap_4 FILLER_44_175 ();
 sg13g2_decap_8 FILLER_44_188 ();
 sg13g2_fill_1 FILLER_44_211 ();
 sg13g2_fill_2 FILLER_44_222 ();
 sg13g2_fill_1 FILLER_44_224 ();
 sg13g2_decap_4 FILLER_44_251 ();
 sg13g2_fill_1 FILLER_44_255 ();
 sg13g2_decap_8 FILLER_44_291 ();
 sg13g2_fill_1 FILLER_44_309 ();
 sg13g2_fill_1 FILLER_44_338 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_fill_2 FILLER_45_140 ();
 sg13g2_fill_1 FILLER_45_142 ();
 sg13g2_fill_2 FILLER_45_230 ();
 sg13g2_fill_1 FILLER_45_232 ();
 sg13g2_fill_1 FILLER_45_247 ();
 sg13g2_fill_1 FILLER_45_260 ();
 sg13g2_decap_8 FILLER_45_286 ();
 sg13g2_fill_1 FILLER_45_293 ();
 sg13g2_decap_4 FILLER_45_304 ();
 sg13g2_fill_2 FILLER_45_308 ();
 sg13g2_fill_2 FILLER_45_317 ();
 sg13g2_fill_2 FILLER_45_330 ();
 sg13g2_fill_2 FILLER_45_364 ();
 sg13g2_fill_1 FILLER_45_374 ();
 sg13g2_fill_2 FILLER_45_393 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_8 FILLER_46_133 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_fill_2 FILLER_46_199 ();
 sg13g2_fill_1 FILLER_46_201 ();
 sg13g2_decap_8 FILLER_46_231 ();
 sg13g2_decap_8 FILLER_46_238 ();
 sg13g2_fill_2 FILLER_46_245 ();
 sg13g2_fill_1 FILLER_46_247 ();
 sg13g2_fill_1 FILLER_46_270 ();
 sg13g2_decap_4 FILLER_46_294 ();
 sg13g2_decap_4 FILLER_46_323 ();
 sg13g2_fill_1 FILLER_46_327 ();
 sg13g2_fill_2 FILLER_46_359 ();
 sg13g2_fill_1 FILLER_46_377 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_4 FILLER_47_154 ();
 sg13g2_fill_1 FILLER_47_158 ();
 sg13g2_fill_1 FILLER_47_177 ();
 sg13g2_fill_1 FILLER_47_183 ();
 sg13g2_decap_8 FILLER_47_205 ();
 sg13g2_decap_8 FILLER_47_212 ();
 sg13g2_fill_2 FILLER_47_224 ();
 sg13g2_fill_1 FILLER_47_226 ();
 sg13g2_fill_2 FILLER_47_289 ();
 sg13g2_fill_2 FILLER_47_346 ();
 sg13g2_fill_1 FILLER_47_364 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_4 FILLER_48_161 ();
 sg13g2_fill_2 FILLER_48_165 ();
 sg13g2_decap_8 FILLER_48_171 ();
 sg13g2_fill_1 FILLER_48_178 ();
 sg13g2_decap_8 FILLER_48_187 ();
 sg13g2_fill_1 FILLER_48_194 ();
 sg13g2_decap_8 FILLER_48_199 ();
 sg13g2_fill_2 FILLER_48_225 ();
 sg13g2_fill_1 FILLER_48_227 ();
 sg13g2_fill_1 FILLER_48_234 ();
 sg13g2_fill_2 FILLER_48_241 ();
 sg13g2_fill_1 FILLER_48_306 ();
 sg13g2_decap_4 FILLER_48_328 ();
 sg13g2_fill_2 FILLER_48_332 ();
 sg13g2_fill_2 FILLER_48_406 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_decap_4 FILLER_49_140 ();
 sg13g2_fill_1 FILLER_49_144 ();
 sg13g2_decap_4 FILLER_49_172 ();
 sg13g2_fill_1 FILLER_49_176 ();
 sg13g2_fill_2 FILLER_49_181 ();
 sg13g2_fill_1 FILLER_49_183 ();
 sg13g2_fill_2 FILLER_49_188 ();
 sg13g2_fill_1 FILLER_49_190 ();
 sg13g2_fill_2 FILLER_49_195 ();
 sg13g2_fill_1 FILLER_49_197 ();
 sg13g2_decap_4 FILLER_49_259 ();
 sg13g2_fill_2 FILLER_49_263 ();
 sg13g2_fill_2 FILLER_49_269 ();
 sg13g2_fill_1 FILLER_49_271 ();
 sg13g2_decap_4 FILLER_49_283 ();
 sg13g2_fill_2 FILLER_49_287 ();
 sg13g2_fill_2 FILLER_49_293 ();
 sg13g2_fill_1 FILLER_49_295 ();
 sg13g2_decap_8 FILLER_49_318 ();
 sg13g2_fill_1 FILLER_49_325 ();
 sg13g2_fill_2 FILLER_49_329 ();
 sg13g2_fill_2 FILLER_49_386 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_decap_8 FILLER_50_119 ();
 sg13g2_decap_8 FILLER_50_126 ();
 sg13g2_decap_8 FILLER_50_133 ();
 sg13g2_decap_8 FILLER_50_140 ();
 sg13g2_fill_1 FILLER_50_147 ();
 sg13g2_fill_1 FILLER_50_206 ();
 sg13g2_fill_2 FILLER_50_213 ();
 sg13g2_fill_1 FILLER_50_234 ();
 sg13g2_decap_8 FILLER_50_240 ();
 sg13g2_decap_8 FILLER_50_255 ();
 sg13g2_decap_8 FILLER_50_262 ();
 sg13g2_fill_1 FILLER_50_269 ();
 sg13g2_decap_8 FILLER_50_274 ();
 sg13g2_decap_8 FILLER_50_281 ();
 sg13g2_fill_2 FILLER_50_288 ();
 sg13g2_decap_4 FILLER_50_295 ();
 sg13g2_decap_4 FILLER_50_312 ();
 sg13g2_fill_2 FILLER_50_316 ();
 sg13g2_fill_1 FILLER_50_365 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_8 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_decap_8 FILLER_51_119 ();
 sg13g2_decap_8 FILLER_51_126 ();
 sg13g2_decap_8 FILLER_51_133 ();
 sg13g2_fill_1 FILLER_51_140 ();
 sg13g2_fill_1 FILLER_51_159 ();
 sg13g2_fill_2 FILLER_51_207 ();
 sg13g2_fill_1 FILLER_51_209 ();
 sg13g2_fill_1 FILLER_51_215 ();
 sg13g2_decap_8 FILLER_51_233 ();
 sg13g2_decap_8 FILLER_51_240 ();
 sg13g2_decap_8 FILLER_51_247 ();
 sg13g2_fill_1 FILLER_51_254 ();
 sg13g2_decap_4 FILLER_51_259 ();
 sg13g2_fill_2 FILLER_51_271 ();
 sg13g2_fill_1 FILLER_51_273 ();
 sg13g2_fill_2 FILLER_51_277 ();
 sg13g2_fill_1 FILLER_51_279 ();
 sg13g2_fill_1 FILLER_51_382 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_8 FILLER_52_112 ();
 sg13g2_decap_8 FILLER_52_119 ();
 sg13g2_decap_4 FILLER_52_126 ();
 sg13g2_fill_1 FILLER_52_130 ();
 sg13g2_fill_2 FILLER_52_179 ();
 sg13g2_fill_2 FILLER_52_195 ();
 sg13g2_decap_4 FILLER_52_214 ();
 sg13g2_decap_4 FILLER_52_222 ();
 sg13g2_fill_2 FILLER_52_226 ();
 sg13g2_fill_1 FILLER_52_232 ();
 sg13g2_fill_2 FILLER_52_237 ();
 sg13g2_fill_1 FILLER_52_239 ();
 sg13g2_decap_8 FILLER_52_245 ();
 sg13g2_fill_2 FILLER_52_252 ();
 sg13g2_decap_4 FILLER_52_262 ();
 sg13g2_fill_1 FILLER_52_266 ();
 sg13g2_fill_2 FILLER_52_308 ();
 sg13g2_decap_8 FILLER_52_342 ();
 sg13g2_fill_1 FILLER_52_363 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_112 ();
 sg13g2_decap_8 FILLER_53_119 ();
 sg13g2_decap_8 FILLER_53_126 ();
 sg13g2_fill_2 FILLER_53_133 ();
 sg13g2_fill_1 FILLER_53_148 ();
 sg13g2_fill_1 FILLER_53_154 ();
 sg13g2_fill_2 FILLER_53_169 ();
 sg13g2_fill_1 FILLER_53_175 ();
 sg13g2_fill_2 FILLER_53_197 ();
 sg13g2_fill_1 FILLER_53_203 ();
 sg13g2_fill_2 FILLER_53_208 ();
 sg13g2_fill_1 FILLER_53_210 ();
 sg13g2_fill_1 FILLER_53_215 ();
 sg13g2_fill_2 FILLER_53_236 ();
 sg13g2_fill_1 FILLER_53_296 ();
 sg13g2_decap_8 FILLER_53_327 ();
 sg13g2_fill_1 FILLER_53_334 ();
 sg13g2_decap_8 FILLER_53_341 ();
 sg13g2_fill_1 FILLER_53_348 ();
 sg13g2_fill_1 FILLER_53_373 ();
 sg13g2_fill_2 FILLER_53_392 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_decap_8 FILLER_54_112 ();
 sg13g2_decap_8 FILLER_54_119 ();
 sg13g2_decap_8 FILLER_54_126 ();
 sg13g2_decap_8 FILLER_54_133 ();
 sg13g2_decap_4 FILLER_54_140 ();
 sg13g2_fill_1 FILLER_54_144 ();
 sg13g2_fill_1 FILLER_54_149 ();
 sg13g2_fill_2 FILLER_54_172 ();
 sg13g2_decap_4 FILLER_54_183 ();
 sg13g2_fill_2 FILLER_54_191 ();
 sg13g2_fill_1 FILLER_54_193 ();
 sg13g2_fill_1 FILLER_54_214 ();
 sg13g2_fill_1 FILLER_54_231 ();
 sg13g2_fill_1 FILLER_54_269 ();
 sg13g2_fill_1 FILLER_54_279 ();
 sg13g2_decap_4 FILLER_54_306 ();
 sg13g2_fill_1 FILLER_54_310 ();
 sg13g2_fill_2 FILLER_54_319 ();
 sg13g2_decap_4 FILLER_54_324 ();
 sg13g2_fill_2 FILLER_54_334 ();
 sg13g2_fill_2 FILLER_54_375 ();
 sg13g2_fill_2 FILLER_54_407 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_decap_8 FILLER_55_112 ();
 sg13g2_decap_8 FILLER_55_119 ();
 sg13g2_decap_8 FILLER_55_126 ();
 sg13g2_fill_2 FILLER_55_179 ();
 sg13g2_fill_1 FILLER_55_225 ();
 sg13g2_fill_2 FILLER_55_234 ();
 sg13g2_fill_1 FILLER_55_266 ();
 sg13g2_decap_8 FILLER_55_270 ();
 sg13g2_fill_1 FILLER_55_281 ();
 sg13g2_decap_8 FILLER_55_304 ();
 sg13g2_decap_4 FILLER_55_311 ();
 sg13g2_fill_1 FILLER_55_367 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_8 FILLER_56_105 ();
 sg13g2_decap_8 FILLER_56_112 ();
 sg13g2_decap_8 FILLER_56_119 ();
 sg13g2_decap_8 FILLER_56_126 ();
 sg13g2_decap_4 FILLER_56_133 ();
 sg13g2_fill_2 FILLER_56_150 ();
 sg13g2_decap_8 FILLER_56_174 ();
 sg13g2_decap_4 FILLER_56_181 ();
 sg13g2_fill_2 FILLER_56_185 ();
 sg13g2_decap_4 FILLER_56_258 ();
 sg13g2_fill_2 FILLER_56_262 ();
 sg13g2_decap_4 FILLER_56_270 ();
 sg13g2_fill_1 FILLER_56_274 ();
 sg13g2_decap_8 FILLER_56_286 ();
 sg13g2_decap_8 FILLER_56_293 ();
 sg13g2_decap_8 FILLER_56_300 ();
 sg13g2_decap_8 FILLER_56_307 ();
 sg13g2_decap_8 FILLER_56_314 ();
 sg13g2_fill_1 FILLER_56_321 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_decap_8 FILLER_57_105 ();
 sg13g2_decap_8 FILLER_57_112 ();
 sg13g2_decap_8 FILLER_57_119 ();
 sg13g2_decap_8 FILLER_57_126 ();
 sg13g2_decap_8 FILLER_57_133 ();
 sg13g2_decap_8 FILLER_57_140 ();
 sg13g2_fill_2 FILLER_57_152 ();
 sg13g2_fill_2 FILLER_57_171 ();
 sg13g2_fill_1 FILLER_57_173 ();
 sg13g2_fill_2 FILLER_57_186 ();
 sg13g2_fill_1 FILLER_57_188 ();
 sg13g2_fill_2 FILLER_57_207 ();
 sg13g2_fill_1 FILLER_57_209 ();
 sg13g2_decap_4 FILLER_57_218 ();
 sg13g2_fill_2 FILLER_57_222 ();
 sg13g2_decap_4 FILLER_57_230 ();
 sg13g2_fill_1 FILLER_57_234 ();
 sg13g2_decap_4 FILLER_57_244 ();
 sg13g2_fill_1 FILLER_57_248 ();
 sg13g2_fill_1 FILLER_57_282 ();
 sg13g2_decap_4 FILLER_57_297 ();
 sg13g2_fill_2 FILLER_57_388 ();
 sg13g2_fill_1 FILLER_57_399 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_8 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_decap_8 FILLER_58_126 ();
 sg13g2_decap_4 FILLER_58_133 ();
 sg13g2_fill_1 FILLER_58_137 ();
 sg13g2_fill_2 FILLER_58_164 ();
 sg13g2_fill_2 FILLER_58_186 ();
 sg13g2_decap_8 FILLER_58_192 ();
 sg13g2_decap_8 FILLER_58_199 ();
 sg13g2_decap_8 FILLER_58_206 ();
 sg13g2_fill_1 FILLER_58_213 ();
 sg13g2_fill_2 FILLER_58_293 ();
 sg13g2_fill_1 FILLER_58_335 ();
 sg13g2_fill_1 FILLER_58_355 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_decap_8 FILLER_59_119 ();
 sg13g2_decap_8 FILLER_59_126 ();
 sg13g2_decap_8 FILLER_59_133 ();
 sg13g2_decap_4 FILLER_59_140 ();
 sg13g2_fill_1 FILLER_59_144 ();
 sg13g2_fill_2 FILLER_59_158 ();
 sg13g2_fill_2 FILLER_59_174 ();
 sg13g2_fill_1 FILLER_59_176 ();
 sg13g2_decap_4 FILLER_59_205 ();
 sg13g2_fill_1 FILLER_59_256 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_decap_8 FILLER_60_105 ();
 sg13g2_decap_8 FILLER_60_112 ();
 sg13g2_decap_8 FILLER_60_119 ();
 sg13g2_decap_8 FILLER_60_126 ();
 sg13g2_decap_8 FILLER_60_133 ();
 sg13g2_fill_2 FILLER_60_140 ();
 sg13g2_fill_2 FILLER_60_173 ();
 sg13g2_fill_2 FILLER_60_191 ();
 sg13g2_decap_8 FILLER_60_261 ();
 sg13g2_fill_1 FILLER_60_272 ();
 sg13g2_fill_2 FILLER_60_310 ();
 sg13g2_fill_2 FILLER_60_348 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_8 FILLER_61_91 ();
 sg13g2_decap_8 FILLER_61_98 ();
 sg13g2_decap_8 FILLER_61_105 ();
 sg13g2_decap_8 FILLER_61_112 ();
 sg13g2_decap_8 FILLER_61_119 ();
 sg13g2_decap_8 FILLER_61_126 ();
 sg13g2_fill_2 FILLER_61_133 ();
 sg13g2_fill_1 FILLER_61_135 ();
 sg13g2_fill_1 FILLER_61_161 ();
 sg13g2_fill_1 FILLER_61_218 ();
 sg13g2_fill_1 FILLER_61_229 ();
 sg13g2_decap_4 FILLER_61_235 ();
 sg13g2_fill_1 FILLER_61_239 ();
 sg13g2_fill_2 FILLER_61_244 ();
 sg13g2_fill_1 FILLER_61_246 ();
 sg13g2_decap_8 FILLER_61_265 ();
 sg13g2_decap_8 FILLER_61_272 ();
 sg13g2_fill_2 FILLER_61_279 ();
 sg13g2_fill_1 FILLER_61_346 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_112 ();
 sg13g2_fill_2 FILLER_62_119 ();
 sg13g2_fill_1 FILLER_62_121 ();
 sg13g2_fill_1 FILLER_62_148 ();
 sg13g2_fill_2 FILLER_62_158 ();
 sg13g2_fill_2 FILLER_62_170 ();
 sg13g2_fill_1 FILLER_62_172 ();
 sg13g2_decap_8 FILLER_62_225 ();
 sg13g2_decap_8 FILLER_62_232 ();
 sg13g2_decap_8 FILLER_62_239 ();
 sg13g2_decap_4 FILLER_62_246 ();
 sg13g2_fill_2 FILLER_62_290 ();
 sg13g2_fill_2 FILLER_62_328 ();
 sg13g2_fill_1 FILLER_62_336 ();
 sg13g2_fill_1 FILLER_62_343 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_8 FILLER_63_105 ();
 sg13g2_decap_8 FILLER_63_112 ();
 sg13g2_decap_8 FILLER_63_119 ();
 sg13g2_decap_4 FILLER_63_126 ();
 sg13g2_fill_1 FILLER_63_130 ();
 sg13g2_fill_2 FILLER_63_156 ();
 sg13g2_fill_2 FILLER_63_178 ();
 sg13g2_fill_1 FILLER_63_180 ();
 sg13g2_decap_8 FILLER_63_185 ();
 sg13g2_fill_1 FILLER_63_192 ();
 sg13g2_fill_2 FILLER_63_207 ();
 sg13g2_decap_4 FILLER_63_259 ();
 sg13g2_fill_1 FILLER_63_263 ();
 sg13g2_fill_2 FILLER_63_321 ();
 sg13g2_fill_1 FILLER_63_362 ();
 sg13g2_fill_1 FILLER_63_367 ();
 sg13g2_fill_1 FILLER_63_382 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_8 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_decap_8 FILLER_64_133 ();
 sg13g2_fill_2 FILLER_64_140 ();
 sg13g2_decap_8 FILLER_64_176 ();
 sg13g2_decap_8 FILLER_64_183 ();
 sg13g2_decap_8 FILLER_64_190 ();
 sg13g2_decap_8 FILLER_64_197 ();
 sg13g2_decap_8 FILLER_64_204 ();
 sg13g2_fill_2 FILLER_64_227 ();
 sg13g2_fill_1 FILLER_64_229 ();
 sg13g2_fill_2 FILLER_64_281 ();
 sg13g2_fill_1 FILLER_64_300 ();
 sg13g2_fill_2 FILLER_64_372 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_decap_4 FILLER_65_119 ();
 sg13g2_fill_2 FILLER_65_123 ();
 sg13g2_fill_1 FILLER_65_179 ();
 sg13g2_fill_2 FILLER_65_188 ();
 sg13g2_fill_1 FILLER_65_194 ();
 sg13g2_fill_2 FILLER_65_203 ();
 sg13g2_fill_1 FILLER_65_210 ();
 sg13g2_fill_2 FILLER_65_223 ();
 sg13g2_fill_2 FILLER_65_304 ();
 sg13g2_fill_1 FILLER_65_324 ();
 sg13g2_fill_1 FILLER_65_388 ();
 sg13g2_fill_2 FILLER_65_398 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_decap_8 FILLER_66_119 ();
 sg13g2_decap_4 FILLER_66_126 ();
 sg13g2_fill_2 FILLER_66_130 ();
 sg13g2_decap_4 FILLER_66_183 ();
 sg13g2_fill_1 FILLER_66_187 ();
 sg13g2_fill_2 FILLER_66_206 ();
 sg13g2_fill_2 FILLER_66_211 ();
 sg13g2_fill_2 FILLER_66_232 ();
 sg13g2_fill_2 FILLER_66_259 ();
 sg13g2_fill_1 FILLER_66_261 ();
 sg13g2_fill_2 FILLER_66_307 ();
 sg13g2_fill_2 FILLER_66_350 ();
 sg13g2_fill_1 FILLER_66_361 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_decap_8 FILLER_67_119 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_fill_2 FILLER_67_149 ();
 sg13g2_fill_1 FILLER_67_151 ();
 sg13g2_decap_8 FILLER_67_156 ();
 sg13g2_decap_4 FILLER_67_163 ();
 sg13g2_fill_1 FILLER_67_167 ();
 sg13g2_decap_4 FILLER_67_177 ();
 sg13g2_fill_1 FILLER_67_274 ();
 sg13g2_fill_2 FILLER_67_380 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_119 ();
 sg13g2_fill_2 FILLER_68_126 ();
 sg13g2_fill_1 FILLER_68_128 ();
 sg13g2_fill_1 FILLER_68_155 ();
 sg13g2_decap_8 FILLER_68_185 ();
 sg13g2_fill_1 FILLER_68_192 ();
 sg13g2_decap_8 FILLER_68_201 ();
 sg13g2_decap_8 FILLER_68_219 ();
 sg13g2_decap_8 FILLER_68_226 ();
 sg13g2_decap_8 FILLER_68_233 ();
 sg13g2_decap_8 FILLER_68_240 ();
 sg13g2_decap_8 FILLER_68_247 ();
 sg13g2_decap_4 FILLER_68_254 ();
 sg13g2_fill_1 FILLER_68_258 ();
 sg13g2_fill_1 FILLER_68_263 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_fill_2 FILLER_69_119 ();
 sg13g2_fill_2 FILLER_69_147 ();
 sg13g2_fill_1 FILLER_69_149 ();
 sg13g2_fill_1 FILLER_69_174 ();
 sg13g2_fill_2 FILLER_69_194 ();
 sg13g2_fill_1 FILLER_69_196 ();
 sg13g2_decap_8 FILLER_69_204 ();
 sg13g2_decap_8 FILLER_69_211 ();
 sg13g2_decap_8 FILLER_69_218 ();
 sg13g2_decap_8 FILLER_69_225 ();
 sg13g2_fill_2 FILLER_69_232 ();
 sg13g2_fill_1 FILLER_69_234 ();
 sg13g2_decap_8 FILLER_69_261 ();
 sg13g2_decap_4 FILLER_69_268 ();
 sg13g2_fill_2 FILLER_69_272 ();
 sg13g2_fill_1 FILLER_69_309 ();
 sg13g2_fill_1 FILLER_69_328 ();
 sg13g2_fill_2 FILLER_69_338 ();
 sg13g2_fill_2 FILLER_69_371 ();
 sg13g2_fill_2 FILLER_69_381 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_fill_2 FILLER_70_126 ();
 sg13g2_fill_1 FILLER_70_128 ();
 sg13g2_fill_2 FILLER_70_144 ();
 sg13g2_fill_1 FILLER_70_146 ();
 sg13g2_fill_2 FILLER_70_155 ();
 sg13g2_fill_1 FILLER_70_157 ();
 sg13g2_fill_2 FILLER_70_181 ();
 sg13g2_decap_8 FILLER_70_191 ();
 sg13g2_fill_2 FILLER_70_198 ();
 sg13g2_fill_1 FILLER_70_200 ();
 sg13g2_decap_4 FILLER_70_206 ();
 sg13g2_fill_2 FILLER_70_218 ();
 sg13g2_fill_1 FILLER_70_220 ();
 sg13g2_fill_2 FILLER_70_236 ();
 sg13g2_fill_2 FILLER_70_262 ();
 sg13g2_fill_2 FILLER_70_272 ();
 sg13g2_fill_1 FILLER_70_377 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_fill_1 FILLER_71_126 ();
 sg13g2_fill_2 FILLER_71_176 ();
 sg13g2_fill_1 FILLER_71_178 ();
 sg13g2_fill_1 FILLER_71_191 ();
 sg13g2_decap_4 FILLER_71_205 ();
 sg13g2_fill_1 FILLER_71_213 ();
 sg13g2_decap_4 FILLER_71_218 ();
 sg13g2_fill_1 FILLER_71_236 ();
 sg13g2_fill_1 FILLER_71_257 ();
 sg13g2_fill_2 FILLER_71_351 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_fill_1 FILLER_72_133 ();
 sg13g2_fill_2 FILLER_72_148 ();
 sg13g2_fill_1 FILLER_72_150 ();
 sg13g2_fill_1 FILLER_72_190 ();
 sg13g2_fill_2 FILLER_72_213 ();
 sg13g2_fill_1 FILLER_72_215 ();
 sg13g2_decap_4 FILLER_72_228 ();
 sg13g2_fill_1 FILLER_72_267 ();
 sg13g2_fill_2 FILLER_72_320 ();
 sg13g2_fill_1 FILLER_72_356 ();
 sg13g2_fill_1 FILLER_72_378 ();
 sg13g2_fill_2 FILLER_72_397 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_4 FILLER_73_147 ();
 sg13g2_fill_1 FILLER_73_151 ();
 sg13g2_fill_2 FILLER_73_213 ();
 sg13g2_fill_1 FILLER_73_246 ();
 sg13g2_fill_2 FILLER_73_273 ();
 sg13g2_fill_1 FILLER_73_278 ();
 sg13g2_fill_2 FILLER_73_283 ();
 sg13g2_fill_1 FILLER_73_315 ();
 sg13g2_fill_1 FILLER_73_339 ();
 sg13g2_fill_2 FILLER_73_352 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_fill_2 FILLER_74_159 ();
 sg13g2_fill_1 FILLER_74_174 ();
 sg13g2_fill_2 FILLER_74_216 ();
 sg13g2_fill_1 FILLER_74_218 ();
 sg13g2_fill_2 FILLER_74_275 ();
 sg13g2_fill_1 FILLER_74_295 ();
 sg13g2_fill_1 FILLER_74_337 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_4 FILLER_75_126 ();
 sg13g2_fill_2 FILLER_75_130 ();
 sg13g2_decap_8 FILLER_75_166 ();
 sg13g2_decap_4 FILLER_75_173 ();
 sg13g2_fill_1 FILLER_75_225 ();
 sg13g2_fill_2 FILLER_75_230 ();
 sg13g2_fill_1 FILLER_75_232 ();
 sg13g2_fill_2 FILLER_75_238 ();
 sg13g2_fill_1 FILLER_75_240 ();
 sg13g2_fill_1 FILLER_75_307 ();
 sg13g2_fill_1 FILLER_75_359 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_fill_2 FILLER_76_140 ();
 sg13g2_fill_1 FILLER_76_142 ();
 sg13g2_decap_4 FILLER_76_151 ();
 sg13g2_decap_4 FILLER_76_159 ();
 sg13g2_fill_1 FILLER_76_163 ();
 sg13g2_fill_2 FILLER_76_176 ();
 sg13g2_fill_1 FILLER_76_239 ();
 sg13g2_fill_1 FILLER_76_249 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_fill_2 FILLER_77_199 ();
 sg13g2_fill_1 FILLER_77_201 ();
 sg13g2_fill_2 FILLER_77_217 ();
 sg13g2_fill_1 FILLER_77_250 ();
 sg13g2_fill_1 FILLER_77_291 ();
 sg13g2_fill_1 FILLER_77_301 ();
 sg13g2_fill_2 FILLER_77_348 ();
 sg13g2_fill_2 FILLER_77_368 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_fill_1 FILLER_78_147 ();
 sg13g2_fill_2 FILLER_78_179 ();
 sg13g2_fill_1 FILLER_78_181 ();
 sg13g2_fill_2 FILLER_78_208 ();
 sg13g2_fill_1 FILLER_78_224 ();
 sg13g2_fill_1 FILLER_78_238 ();
 sg13g2_fill_1 FILLER_78_265 ();
 sg13g2_fill_1 FILLER_78_330 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_fill_2 FILLER_79_185 ();
 sg13g2_fill_1 FILLER_79_187 ();
 sg13g2_fill_2 FILLER_79_197 ();
 sg13g2_fill_1 FILLER_79_199 ();
 sg13g2_fill_2 FILLER_79_252 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_8 FILLER_80_116 ();
 sg13g2_decap_8 FILLER_80_123 ();
 sg13g2_decap_8 FILLER_80_130 ();
 sg13g2_decap_8 FILLER_80_137 ();
 sg13g2_decap_4 FILLER_80_144 ();
 sg13g2_fill_1 FILLER_80_148 ();
 sg13g2_fill_1 FILLER_80_182 ();
 sg13g2_fill_1 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_192 ();
 sg13g2_decap_8 FILLER_80_199 ();
 sg13g2_decap_4 FILLER_80_206 ();
 sg13g2_fill_1 FILLER_80_210 ();
 sg13g2_decap_8 FILLER_80_215 ();
 sg13g2_decap_8 FILLER_80_225 ();
 sg13g2_decap_4 FILLER_80_236 ();
 sg13g2_fill_1 FILLER_80_290 ();
 sg13g2_fill_1 FILLER_80_301 ();
 sg13g2_fill_1 FILLER_80_387 ();
 sg13g2_fill_2 FILLER_80_392 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net329;
 assign uio_oe[5] = net330;
 assign uio_oe[6] = net331;
 assign uio_oe[7] = net332;
 assign uio_out[0] = net13;
 assign uio_out[1] = net14;
 assign uio_out[2] = net15;
 assign uio_out[3] = net16;
endmodule

module tt_um_spacewar (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire clknet_0_clk;
 wire \counter[0] ;
 wire \counter[10] ;
 wire \counter[11] ;
 wire \counter[12] ;
 wire \counter[13] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire \driver.decoder.data_reg[0] ;
 wire \driver.decoder.data_reg[10] ;
 wire \driver.decoder.data_reg[11] ;
 wire \driver.decoder.data_reg[1] ;
 wire \driver.decoder.data_reg[2] ;
 wire \driver.decoder.data_reg[3] ;
 wire \driver.decoder.data_reg[4] ;
 wire \driver.decoder.data_reg[5] ;
 wire \driver.decoder.data_reg[6] ;
 wire \driver.decoder.data_reg[7] ;
 wire \driver.decoder.data_reg[8] ;
 wire \driver.decoder.data_reg[9] ;
 wire \driver.driver.pmod_clk_prev ;
 wire \driver.driver.pmod_clk_sync[0] ;
 wire \driver.driver.pmod_clk_sync[1] ;
 wire \driver.driver.pmod_data_sync[0] ;
 wire \driver.driver.pmod_data_sync[1] ;
 wire \driver.driver.pmod_latch_prev ;
 wire \driver.driver.pmod_latch_sync[0] ;
 wire \driver.driver.pmod_latch_sync[1] ;
 wire \driver.driver.shift_reg[0] ;
 wire \driver.driver.shift_reg[10] ;
 wire \driver.driver.shift_reg[11] ;
 wire \driver.driver.shift_reg[1] ;
 wire \driver.driver.shift_reg[2] ;
 wire \driver.driver.shift_reg[3] ;
 wire \driver.driver.shift_reg[4] ;
 wire \driver.driver.shift_reg[5] ;
 wire \driver.driver.shift_reg[6] ;
 wire \driver.driver.shift_reg[7] ;
 wire \driver.driver.shift_reg[8] ;
 wire \driver.driver.shift_reg[9] ;
 wire hsync;
 wire \pix_x[0] ;
 wire \pix_x[1] ;
 wire \pix_x[2] ;
 wire \pix_x[3] ;
 wire \pix_x[4] ;
 wire \pix_x[5] ;
 wire \pix_x[6] ;
 wire \pix_x[7] ;
 wire \pix_x[8] ;
 wire \pix_x[9] ;
 wire \pix_y[0] ;
 wire \pix_y[1] ;
 wire \pix_y[2] ;
 wire \pix_y[3] ;
 wire \pix_y[4] ;
 wire \pix_y[5] ;
 wire \pix_y[6] ;
 wire \pix_y[7] ;
 wire \pix_y[8] ;
 wire \pix_y[9] ;
 wire \square_x[0] ;
 wire \square_x[1] ;
 wire \square_x[2] ;
 wire \square_x[3] ;
 wire \square_x[4] ;
 wire \square_x[5] ;
 wire \square_x[6] ;
 wire \square_x[7] ;
 wire \square_x[8] ;
 wire \square_x[9] ;
 wire \square_y[0] ;
 wire \square_y[1] ;
 wire \square_y[2] ;
 wire \square_y[3] ;
 wire \square_y[4] ;
 wire \square_y[5] ;
 wire \square_y[6] ;
 wire \square_y[7] ;
 wire \square_y[8] ;
 wire \square_y[9] ;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire \vga_sync_gen.vsync ;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;

 sg13g2_inv_1 _0968_ (.Y(_0120_),
    .A(net163));
 sg13g2_inv_1 _0969_ (.Y(_0121_),
    .A(net170));
 sg13g2_inv_1 _0970_ (.Y(_0122_),
    .A(net168));
 sg13g2_inv_1 _0971_ (.Y(_0123_),
    .A(net171));
 sg13g2_inv_1 _0972_ (.Y(_0124_),
    .A(net174));
 sg13g2_inv_1 _0973_ (.Y(_0125_),
    .A(net159));
 sg13g2_inv_1 _0974_ (.Y(_0126_),
    .A(net165));
 sg13g2_inv_1 _0975_ (.Y(_0127_),
    .A(net153));
 sg13g2_inv_1 _0976_ (.Y(_0128_),
    .A(net173));
 sg13g2_inv_1 _0977_ (.Y(_0129_),
    .A(net157));
 sg13g2_inv_1 _0978_ (.Y(_0130_),
    .A(\driver.driver.shift_reg[0] ));
 sg13g2_inv_1 _0979_ (.Y(_0131_),
    .A(net130));
 sg13g2_inv_1 _0980_ (.Y(_0132_),
    .A(\square_y[9] ));
 sg13g2_inv_1 _0981_ (.Y(_0133_),
    .A(\square_y[8] ));
 sg13g2_inv_1 _0982_ (.Y(_0134_),
    .A(\square_y[7] ));
 sg13g2_inv_1 _0983_ (.Y(_0135_),
    .A(\square_y[6] ));
 sg13g2_inv_1 _0984_ (.Y(_0136_),
    .A(\square_y[5] ));
 sg13g2_inv_1 _0985_ (.Y(_0137_),
    .A(\square_y[4] ));
 sg13g2_inv_1 _0986_ (.Y(_0138_),
    .A(\square_y[0] ));
 sg13g2_inv_1 _0987_ (.Y(_0139_),
    .A(net119));
 sg13g2_inv_1 _0988_ (.Y(_0140_),
    .A(\square_x[9] ));
 sg13g2_inv_1 _0989_ (.Y(_0141_),
    .A(\square_x[8] ));
 sg13g2_inv_1 _0990_ (.Y(_0142_),
    .A(\square_x[7] ));
 sg13g2_inv_1 _0991_ (.Y(_0143_),
    .A(\square_x[2] ));
 sg13g2_inv_1 _0992_ (.Y(_0144_),
    .A(\square_x[1] ));
 sg13g2_inv_1 _0993_ (.Y(_0145_),
    .A(net141));
 sg13g2_inv_1 _0994_ (.Y(_0146_),
    .A(net274));
 sg13g2_inv_1 _0995_ (.Y(_0147_),
    .A(net276));
 sg13g2_inv_2 _0996_ (.Y(_0148_),
    .A(\pix_x[8] ));
 sg13g2_inv_2 _0997_ (.Y(_0149_),
    .A(net260));
 sg13g2_inv_2 _0998_ (.Y(_0150_),
    .A(net311));
 sg13g2_inv_2 _0999_ (.Y(_0151_),
    .A(\pix_y[8] ));
 sg13g2_inv_2 _1000_ (.Y(_0152_),
    .A(\pix_y[6] ));
 sg13g2_inv_1 _1001_ (.Y(_0153_),
    .A(net243));
 sg13g2_inv_1 _1002_ (.Y(_0154_),
    .A(net245));
 sg13g2_inv_1 _1003_ (.Y(_0155_),
    .A(net246));
 sg13g2_inv_2 _1004_ (.Y(_0156_),
    .A(net249));
 sg13g2_inv_2 _1005_ (.Y(_0157_),
    .A(net305));
 sg13g2_inv_1 _1006_ (.Y(_0158_),
    .A(net255));
 sg13g2_inv_1 _1007_ (.Y(_0159_),
    .A(net147));
 sg13g2_inv_1 _1008_ (.Y(_0160_),
    .A(net139));
 sg13g2_inv_1 _1009_ (.Y(_0161_),
    .A(net135));
 sg13g2_inv_1 _1010_ (.Y(_0162_),
    .A(net155));
 sg13g2_inv_1 _1011_ (.Y(_0163_),
    .A(net195));
 sg13g2_inv_1 _1012_ (.Y(_0164_),
    .A(net175));
 sg13g2_inv_1 _1013_ (.Y(_0165_),
    .A(net194));
 sg13g2_inv_2 _1014_ (.Y(_0166_),
    .A(net178));
 sg13g2_inv_1 _1015_ (.Y(_0167_),
    .A(net143));
 sg13g2_inv_1 _1016_ (.Y(_0168_),
    .A(net149));
 sg13g2_inv_1 _1017_ (.Y(_0169_),
    .A(net137));
 sg13g2_inv_1 _1018_ (.Y(_0170_),
    .A(net145));
 sg13g2_inv_1 _1019_ (.Y(_0171_),
    .A(net269));
 sg13g2_inv_1 _1020_ (.Y(_0172_),
    .A(net261));
 sg13g2_inv_1 _1021_ (.Y(_0173_),
    .A(net262));
 sg13g2_inv_2 _1022_ (.Y(_0174_),
    .A(\pix_x[3] ));
 sg13g2_inv_2 _1023_ (.Y(_0175_),
    .A(\pix_x[2] ));
 sg13g2_inv_1 _1024_ (.Y(_0176_),
    .A(net283));
 sg13g2_inv_2 _1025_ (.Y(_0177_),
    .A(\pix_x[1] ));
 sg13g2_inv_1 _1026_ (.Y(_0178_),
    .A(_0020_));
 sg13g2_inv_1 _1027_ (.Y(_0179_),
    .A(_0022_));
 sg13g2_inv_1 _1028_ (.Y(_0180_),
    .A(_0025_));
 sg13g2_inv_1 _1029_ (.Y(_0181_),
    .A(_0019_));
 sg13g2_inv_1 _1030_ (.Y(_0182_),
    .A(_0013_));
 sg13g2_nand3_1 _1031_ (.B(_0155_),
    .C(net255),
    .A(net245),
    .Y(_0183_));
 sg13g2_and2_2 _1032_ (.A(\pix_y[6] ),
    .B(net243),
    .X(_0184_));
 sg13g2_nand2_2 _1033_ (.Y(_0185_),
    .A(\pix_y[6] ),
    .B(net243));
 sg13g2_nor2b_1 _1034_ (.A(\pix_y[2] ),
    .B_N(net249),
    .Y(_0186_));
 sg13g2_nand2b_1 _1035_ (.Y(_0187_),
    .B(net248),
    .A_N(net250));
 sg13g2_nand2b_1 _1036_ (.Y(_0188_),
    .B(net242),
    .A_N(net292));
 sg13g2_nor4_1 _1037_ (.A(_0183_),
    .B(_0185_),
    .C(_0187_),
    .D(net293),
    .Y(_0001_));
 sg13g2_nor2_2 _1038_ (.A(\pix_x[5] ),
    .B(net263),
    .Y(_0189_));
 sg13g2_nor3_2 _1039_ (.A(\pix_x[6] ),
    .B(net262),
    .C(net263),
    .Y(_0190_));
 sg13g2_nor2_2 _1040_ (.A(net258),
    .B(_0150_),
    .Y(_0191_));
 sg13g2_nand3_1 _1041_ (.B(net262),
    .C(net263),
    .A(net318),
    .Y(_0192_));
 sg13g2_nand3_1 _1042_ (.B(_0191_),
    .C(_0192_),
    .A(net259),
    .Y(_0193_));
 sg13g2_nor2_1 _1043_ (.A(_0190_),
    .B(_0193_),
    .Y(_0000_));
 sg13g2_nand4_1 _1044_ (.B(\driver.decoder.data_reg[8] ),
    .C(\driver.decoder.data_reg[11] ),
    .A(\driver.decoder.data_reg[9] ),
    .Y(_0194_),
    .D(\driver.decoder.data_reg[10] ));
 sg13g2_nand4_1 _1045_ (.B(\driver.decoder.data_reg[0] ),
    .C(\driver.decoder.data_reg[3] ),
    .A(\driver.decoder.data_reg[1] ),
    .Y(_0195_),
    .D(\driver.decoder.data_reg[2] ));
 sg13g2_nor2_2 _1046_ (.A(_0165_),
    .B(_0166_),
    .Y(_0196_));
 sg13g2_nand4_1 _1047_ (.B(\driver.decoder.data_reg[4] ),
    .C(\driver.decoder.data_reg[7] ),
    .A(\driver.decoder.data_reg[5] ),
    .Y(_0197_),
    .D(\driver.decoder.data_reg[6] ));
 sg13g2_or3_1 _1048_ (.A(_0194_),
    .B(_0195_),
    .C(_0197_),
    .X(_0198_));
 sg13g2_and2_1 _1049_ (.A(net245),
    .B(net246),
    .X(_0199_));
 sg13g2_nand2_2 _1050_ (.Y(_0200_),
    .A(net244),
    .B(net247));
 sg13g2_nor2_1 _1051_ (.A(net241),
    .B(net242),
    .Y(_0201_));
 sg13g2_nand2_2 _1052_ (.Y(_0202_),
    .A(_0184_),
    .B(_0201_));
 sg13g2_nor2_1 _1053_ (.A(_0152_),
    .B(_0200_),
    .Y(_0203_));
 sg13g2_nor2_1 _1054_ (.A(_0200_),
    .B(_0202_),
    .Y(_0204_));
 sg13g2_nor4_2 _1055_ (.A(_0148_),
    .B(net257),
    .C(_0200_),
    .Y(_0205_),
    .D(_0202_));
 sg13g2_nand3_1 _1056_ (.B(_0150_),
    .C(_0204_),
    .A(net258),
    .Y(_0206_));
 sg13g2_nor2b_1 _1057_ (.A(net264),
    .B_N(\pix_x[5] ),
    .Y(_0207_));
 sg13g2_and4_1 _1058_ (.A(net259),
    .B(net261),
    .C(_0205_),
    .D(net236),
    .X(_0208_));
 sg13g2_nand4_1 _1059_ (.B(net261),
    .C(_0205_),
    .A(net259),
    .Y(_0209_),
    .D(net236));
 sg13g2_nor2_2 _1060_ (.A(net255),
    .B(\pix_y[0] ),
    .Y(_0210_));
 sg13g2_or2_2 _1061_ (.X(_0211_),
    .B(\pix_y[0] ),
    .A(net255));
 sg13g2_nand2b_1 _1062_ (.Y(_0212_),
    .B(net250),
    .A_N(net248));
 sg13g2_nand3b_1 _1063_ (.B(net245),
    .C(\pix_y[6] ),
    .Y(_0213_),
    .A_N(\pix_y[7] ));
 sg13g2_nor2_1 _1064_ (.A(net246),
    .B(_0213_),
    .Y(_0214_));
 sg13g2_nor4_1 _1065_ (.A(net246),
    .B(_0211_),
    .C(_0212_),
    .D(_0213_),
    .Y(_0215_));
 sg13g2_nand4_1 _1066_ (.B(net250),
    .C(_0210_),
    .A(_0156_),
    .Y(_0216_),
    .D(_0214_));
 sg13g2_nor2_1 _1067_ (.A(net248),
    .B(net250),
    .Y(_0217_));
 sg13g2_o21ai_1 _1068_ (.B1(_0156_),
    .Y(_0218_),
    .A1(_0157_),
    .A2(_0210_));
 sg13g2_a21oi_1 _1069_ (.A1(net250),
    .A2(_0211_),
    .Y(_0219_),
    .B1(net248));
 sg13g2_a21oi_1 _1070_ (.A1(\pix_y[6] ),
    .A2(_0178_),
    .Y(_0220_),
    .B1(\pix_y[7] ));
 sg13g2_a21oi_1 _1071_ (.A1(_0214_),
    .A2(_0219_),
    .Y(_0221_),
    .B1(_0220_));
 sg13g2_a21o_1 _1072_ (.A2(_0219_),
    .A1(_0214_),
    .B1(_0220_),
    .X(_0222_));
 sg13g2_nand2_1 _1073_ (.Y(_0223_),
    .A(_0153_),
    .B(_0201_));
 sg13g2_a21o_1 _1074_ (.A2(_0218_),
    .A1(_0203_),
    .B1(_0223_),
    .X(_0224_));
 sg13g2_nor4_1 _1075_ (.A(_0152_),
    .B(net243),
    .C(_0211_),
    .D(_0212_),
    .Y(_0225_));
 sg13g2_a221oi_1 _1076_ (.B2(_0199_),
    .C1(_0223_),
    .B1(_0225_),
    .A1(_0203_),
    .Y(_0226_),
    .A2(_0218_));
 sg13g2_a221oi_1 _1077_ (.B2(_0199_),
    .C1(_0224_),
    .B1(_0225_),
    .A1(_0216_),
    .Y(_0227_),
    .A2(_0222_));
 sg13g2_o21ai_1 _1078_ (.B1(_0226_),
    .Y(_0228_),
    .A1(_0215_),
    .A2(_0221_));
 sg13g2_nor2b_1 _1079_ (.A(net259),
    .B_N(net261),
    .Y(_0229_));
 sg13g2_nand2b_1 _1080_ (.Y(_0230_),
    .B(net263),
    .A_N(\pix_x[5] ));
 sg13g2_nor3_2 _1081_ (.A(net260),
    .B(_0172_),
    .C(_0230_),
    .Y(_0231_));
 sg13g2_and2_1 _1082_ (.A(_0191_),
    .B(_0231_),
    .X(_0232_));
 sg13g2_nand2_1 _1083_ (.Y(_0233_),
    .A(_0191_),
    .B(_0231_));
 sg13g2_nor2_1 _1084_ (.A(_0228_),
    .B(_0233_),
    .Y(_0234_));
 sg13g2_nand2_2 _1085_ (.Y(_0235_),
    .A(_0227_),
    .B(_0232_));
 sg13g2_nor2_1 _1086_ (.A(net259),
    .B(net261),
    .Y(_0236_));
 sg13g2_nand2_1 _1087_ (.Y(_0237_),
    .A(_0149_),
    .B(_0172_));
 sg13g2_nor2_2 _1088_ (.A(net283),
    .B(\pix_x[1] ),
    .Y(_0238_));
 sg13g2_nor2_1 _1089_ (.A(\pix_x[3] ),
    .B(\pix_x[2] ),
    .Y(_0239_));
 sg13g2_nand4_1 _1090_ (.B(_0236_),
    .C(_0238_),
    .A(net236),
    .Y(_0240_),
    .D(_0239_));
 sg13g2_nand2_1 _1091_ (.Y(_0241_),
    .A(_0021_),
    .B(_0240_));
 sg13g2_nor2_2 _1092_ (.A(net258),
    .B(net257),
    .Y(_0242_));
 sg13g2_a21oi_1 _1093_ (.A1(net262),
    .A2(net263),
    .Y(_0243_),
    .B1(_0237_));
 sg13g2_and3_1 _1094_ (.X(_0244_),
    .A(_0241_),
    .B(_0242_),
    .C(_0243_));
 sg13g2_nand3_1 _1095_ (.B(_0242_),
    .C(_0243_),
    .A(_0241_),
    .Y(_0245_));
 sg13g2_nand2_2 _1096_ (.Y(_0246_),
    .A(_0227_),
    .B(_0244_));
 sg13g2_o21ai_1 _1097_ (.B1(_0227_),
    .Y(_0247_),
    .A1(_0232_),
    .A2(_0244_));
 sg13g2_a21oi_2 _1098_ (.B1(_0228_),
    .Y(_0248_),
    .A2(_0245_),
    .A1(_0233_));
 sg13g2_xnor2_1 _1099_ (.Y(_0249_),
    .A(_0027_),
    .B(net217));
 sg13g2_xnor2_1 _1100_ (.Y(_0250_),
    .A(_0027_),
    .B(_0248_));
 sg13g2_a21oi_2 _1101_ (.B1(_0179_),
    .Y(_0251_),
    .A2(_0210_),
    .A1(_0186_));
 sg13g2_o21ai_1 _1102_ (.B1(_0022_),
    .Y(_0252_),
    .A1(_0187_),
    .A2(_0211_));
 sg13g2_nor2_2 _1103_ (.A(net245),
    .B(_0252_),
    .Y(_0253_));
 sg13g2_nor2_2 _1104_ (.A(net244),
    .B(net247),
    .Y(_0254_));
 sg13g2_o21ai_1 _1105_ (.B1(_0154_),
    .Y(_0255_),
    .A1(_0155_),
    .A2(_0251_));
 sg13g2_a21oi_1 _1106_ (.A1(net247),
    .A2(_0252_),
    .Y(_0256_),
    .B1(net245));
 sg13g2_a21oi_1 _1107_ (.A1(_0251_),
    .A2(_0254_),
    .Y(_0257_),
    .B1(_0202_));
 sg13g2_a21o_1 _1108_ (.A2(_0254_),
    .A1(_0251_),
    .B1(_0202_),
    .X(_0258_));
 sg13g2_and2_1 _1109_ (.A(_0149_),
    .B(_0190_),
    .X(_0259_));
 sg13g2_nand2_1 _1110_ (.Y(_0260_),
    .A(_0191_),
    .B(_0259_));
 sg13g2_nor3_1 _1111_ (.A(_0255_),
    .B(_0258_),
    .C(_0260_),
    .Y(_0261_));
 sg13g2_nand4_1 _1112_ (.B(_0256_),
    .C(_0257_),
    .A(_0191_),
    .Y(_0262_),
    .D(_0259_));
 sg13g2_nor2_1 _1113_ (.A(_0208_),
    .B(net221),
    .Y(_0263_));
 sg13g2_nand2_1 _1114_ (.Y(_0264_),
    .A(_0209_),
    .B(_0262_));
 sg13g2_nand3_1 _1115_ (.B(_0229_),
    .C(_0242_),
    .A(net236),
    .Y(_0265_));
 sg13g2_nor4_1 _1116_ (.A(\pix_y[6] ),
    .B(net243),
    .C(_0188_),
    .D(_0199_),
    .Y(_0266_));
 sg13g2_o21ai_1 _1117_ (.B1(_0266_),
    .Y(_0267_),
    .A1(net246),
    .A2(_0251_));
 sg13g2_nor3_2 _1118_ (.A(_0253_),
    .B(_0265_),
    .C(_0267_),
    .Y(_0268_));
 sg13g2_inv_2 _1119_ (.Y(_0269_),
    .A(_0268_));
 sg13g2_nor3_2 _1120_ (.A(_0253_),
    .B(_0260_),
    .C(_0267_),
    .Y(_0270_));
 sg13g2_inv_1 _1121_ (.Y(_0271_),
    .A(_0270_));
 sg13g2_and4_2 _1122_ (.A(_0191_),
    .B(_0204_),
    .C(net236),
    .D(_0236_),
    .X(_0272_));
 sg13g2_nor2_2 _1123_ (.A(_0270_),
    .B(_0272_),
    .Y(_0273_));
 sg13g2_or2_1 _1124_ (.X(_0274_),
    .B(_0272_),
    .A(_0270_));
 sg13g2_nor2_1 _1125_ (.A(net220),
    .B(_0270_),
    .Y(_0275_));
 sg13g2_or2_1 _1126_ (.X(_0276_),
    .B(_0270_),
    .A(net220));
 sg13g2_nor3_2 _1127_ (.A(_0268_),
    .B(_0270_),
    .C(_0272_),
    .Y(_0277_));
 sg13g2_nor3_1 _1128_ (.A(_0255_),
    .B(_0258_),
    .C(_0265_),
    .Y(_0278_));
 sg13g2_nand3b_1 _1129_ (.B(_0256_),
    .C(_0257_),
    .Y(_0279_),
    .A_N(_0265_));
 sg13g2_and2_1 _1130_ (.A(_0189_),
    .B(_0229_),
    .X(_0280_));
 sg13g2_and4_2 _1131_ (.A(_0184_),
    .B(_0199_),
    .C(_0201_),
    .D(_0242_),
    .X(_0281_));
 sg13g2_and2_2 _1132_ (.A(_0280_),
    .B(_0281_),
    .X(_0282_));
 sg13g2_nand2_2 _1133_ (.Y(_0283_),
    .A(_0280_),
    .B(_0281_));
 sg13g2_and3_1 _1134_ (.X(_0284_),
    .A(net259),
    .B(_0190_),
    .C(_0281_));
 sg13g2_and3_2 _1135_ (.X(_0285_),
    .A(net259),
    .B(_0190_),
    .C(_0281_));
 sg13g2_nand3_1 _1136_ (.B(_0190_),
    .C(_0281_),
    .A(net259),
    .Y(_0286_));
 sg13g2_and2_1 _1137_ (.A(_0283_),
    .B(_0286_),
    .X(_0287_));
 sg13g2_nand2_2 _1138_ (.Y(_0288_),
    .A(_0279_),
    .B(_0287_));
 sg13g2_nor4_2 _1139_ (.A(net216),
    .B(net220),
    .C(_0274_),
    .Y(_0289_),
    .D(_0288_));
 sg13g2_mux2_1 _1140_ (.A0(\pix_y[2] ),
    .A1(_0250_),
    .S(_0289_),
    .X(_0290_));
 sg13g2_mux2_1 _1141_ (.A0(_0157_),
    .A1(_0249_),
    .S(_0289_),
    .X(_0291_));
 sg13g2_xnor2_1 _1142_ (.Y(_0292_),
    .A(net246),
    .B(_0217_));
 sg13g2_nor2_1 _1143_ (.A(_0180_),
    .B(_0213_),
    .Y(_0293_));
 sg13g2_nand2_1 _1144_ (.Y(_0294_),
    .A(_0292_),
    .B(_0293_));
 sg13g2_nand2_1 _1145_ (.Y(_0295_),
    .A(net242),
    .B(_0024_));
 sg13g2_o21ai_1 _1146_ (.B1(_0151_),
    .Y(_0296_),
    .A1(_0185_),
    .A2(_0200_));
 sg13g2_nor2_1 _1147_ (.A(_0151_),
    .B(_0154_),
    .Y(_0297_));
 sg13g2_nand3_1 _1148_ (.B(_0184_),
    .C(_0199_),
    .A(net242),
    .Y(_0298_));
 sg13g2_xor2_1 _1149_ (.B(_0023_),
    .A(net243),
    .X(_0299_));
 sg13g2_xor2_1 _1150_ (.B(_0295_),
    .A(net241),
    .X(_0300_));
 sg13g2_and4_1 _1151_ (.A(_0203_),
    .B(_0298_),
    .C(_0299_),
    .D(_0300_),
    .X(_0301_));
 sg13g2_a21oi_1 _1152_ (.A1(_0296_),
    .A2(_0301_),
    .Y(_0302_),
    .B1(net222));
 sg13g2_o21ai_1 _1153_ (.B1(_0302_),
    .Y(_0303_),
    .A1(net217),
    .A2(_0294_));
 sg13g2_nor3_1 _1154_ (.A(net244),
    .B(net247),
    .C(net248),
    .Y(_0304_));
 sg13g2_xnor2_1 _1155_ (.Y(_0305_),
    .A(net242),
    .B(_0304_));
 sg13g2_nor2_1 _1156_ (.A(_0178_),
    .B(_0185_),
    .Y(_0306_));
 sg13g2_xor2_1 _1157_ (.B(net248),
    .A(net247),
    .X(_0307_));
 sg13g2_xnor2_1 _1158_ (.Y(_0308_),
    .A(_0025_),
    .B(_0295_));
 sg13g2_nand4_1 _1159_ (.B(_0306_),
    .C(_0307_),
    .A(_0305_),
    .Y(_0309_),
    .D(_0308_));
 sg13g2_a21oi_1 _1160_ (.A1(net222),
    .A2(_0309_),
    .Y(_0310_),
    .B1(_0276_));
 sg13g2_nor2b_1 _1161_ (.A(_0254_),
    .B_N(_0026_),
    .Y(_0311_));
 sg13g2_nand4_1 _1162_ (.B(_0025_),
    .C(_0200_),
    .A(net242),
    .Y(_0312_),
    .D(_0311_));
 sg13g2_a21oi_1 _1163_ (.A1(net244),
    .A2(_0020_),
    .Y(_0313_),
    .B1(_0023_));
 sg13g2_and3_1 _1164_ (.X(_0314_),
    .A(net244),
    .B(_0020_),
    .C(_0023_));
 sg13g2_nor4_2 _1165_ (.A(_0307_),
    .B(_0312_),
    .C(_0313_),
    .Y(_0315_),
    .D(_0314_));
 sg13g2_a21o_1 _1166_ (.A2(_0315_),
    .A1(_0276_),
    .B1(net218),
    .X(_0316_));
 sg13g2_a221oi_1 _1167_ (.B2(_0276_),
    .C1(net218),
    .B1(_0315_),
    .A1(_0303_),
    .Y(_0317_),
    .A2(_0310_));
 sg13g2_a21o_2 _1168_ (.A2(_0310_),
    .A1(_0303_),
    .B1(_0316_),
    .X(_0318_));
 sg13g2_and2_1 _1169_ (.A(net219),
    .B(_0309_),
    .X(_0319_));
 sg13g2_nand2_2 _1170_ (.Y(_0320_),
    .A(net219),
    .B(_0309_));
 sg13g2_nor2_2 _1171_ (.A(_0317_),
    .B(_0319_),
    .Y(_0321_));
 sg13g2_nand2_2 _1172_ (.Y(_0322_),
    .A(_0318_),
    .B(_0320_));
 sg13g2_nand2_1 _1173_ (.Y(_0323_),
    .A(net222),
    .B(net207));
 sg13g2_nor2_1 _1174_ (.A(_0322_),
    .B(_0323_),
    .Y(_0324_));
 sg13g2_nand2_1 _1175_ (.Y(_0325_),
    .A(net239),
    .B(net207));
 sg13g2_o21ai_1 _1176_ (.B1(_0325_),
    .Y(_0326_),
    .A1(_0322_),
    .A2(_0323_));
 sg13g2_o21ai_1 _1177_ (.B1(net240),
    .Y(_0327_),
    .A1(net217),
    .A2(_0294_));
 sg13g2_or4_1 _1178_ (.A(net222),
    .B(net220),
    .C(_0270_),
    .D(net218),
    .X(_0328_));
 sg13g2_o21ai_1 _1179_ (.B1(_0156_),
    .Y(_0329_),
    .A1(net250),
    .A2(net217));
 sg13g2_a21oi_1 _1180_ (.A1(_0186_),
    .A2(_0248_),
    .Y(_0330_),
    .B1(_0328_));
 sg13g2_and2_1 _1181_ (.A(_0022_),
    .B(_0328_),
    .X(_0331_));
 sg13g2_a22oi_1 _1182_ (.Y(_0332_),
    .B1(_0329_),
    .B2(_0330_),
    .A2(_0328_),
    .A1(_0022_));
 sg13g2_a21o_1 _1183_ (.A2(_0330_),
    .A1(_0329_),
    .B1(_0331_),
    .X(_0333_));
 sg13g2_nor2_1 _1184_ (.A(net251),
    .B(_0285_),
    .Y(_0334_));
 sg13g2_nand2_1 _1185_ (.Y(_0335_),
    .A(_0279_),
    .B(_0334_));
 sg13g2_nor4_1 _1186_ (.A(net216),
    .B(_0274_),
    .C(_0282_),
    .D(_0335_),
    .Y(_0336_));
 sg13g2_nor2b_1 _1187_ (.A(\pix_x[2] ),
    .B_N(\pix_x[3] ),
    .Y(_0337_));
 sg13g2_and2_1 _1188_ (.A(_0238_),
    .B(_0337_),
    .X(_0338_));
 sg13g2_a21o_1 _1189_ (.A2(_0337_),
    .A1(_0238_),
    .B1(_0017_),
    .X(_0339_));
 sg13g2_a21o_1 _1190_ (.A2(_0339_),
    .A1(_0231_),
    .B1(_0280_),
    .X(_0340_));
 sg13g2_nand3_1 _1191_ (.B(_0189_),
    .C(_0229_),
    .A(_0017_),
    .Y(_0341_));
 sg13g2_a21o_1 _1192_ (.A2(_0341_),
    .A1(_0237_),
    .B1(_0338_),
    .X(_0342_));
 sg13g2_nand2_1 _1193_ (.Y(_0343_),
    .A(_0231_),
    .B(_0338_));
 sg13g2_and4_1 _1194_ (.A(_0205_),
    .B(_0340_),
    .C(_0342_),
    .D(_0343_),
    .X(_0344_));
 sg13g2_and4_2 _1195_ (.A(_0205_),
    .B(_0340_),
    .C(_0342_),
    .D(_0343_),
    .X(_0345_));
 sg13g2_nand2b_2 _1196_ (.Y(_0346_),
    .B(_0247_),
    .A_N(_0345_));
 sg13g2_a21oi_1 _1197_ (.A1(net252),
    .A2(_0346_),
    .Y(_0347_),
    .B1(_0336_));
 sg13g2_nor2_1 _1198_ (.A(net206),
    .B(_0347_),
    .Y(_0348_));
 sg13g2_a221oi_1 _1199_ (.B2(_0321_),
    .C1(_0332_),
    .B1(_0348_),
    .A1(_0326_),
    .Y(_0349_),
    .A2(_0327_));
 sg13g2_nand2_1 _1200_ (.Y(_0350_),
    .A(_0246_),
    .B(_0263_));
 sg13g2_nor3_1 _1201_ (.A(net251),
    .B(_0248_),
    .C(net216),
    .Y(_0351_));
 sg13g2_a21oi_1 _1202_ (.A1(net251),
    .A2(_0224_),
    .Y(_0352_),
    .B1(_0351_));
 sg13g2_or2_1 _1203_ (.X(_0353_),
    .B(_0352_),
    .A(net206));
 sg13g2_a21o_1 _1204_ (.A2(_0277_),
    .A1(_0263_),
    .B1(net239),
    .X(_0354_));
 sg13g2_o21ai_1 _1205_ (.B1(_0354_),
    .Y(_0355_),
    .A1(net253),
    .A2(_0346_));
 sg13g2_a21oi_1 _1206_ (.A1(net206),
    .A2(_0355_),
    .Y(_0356_),
    .B1(_0322_));
 sg13g2_a21oi_1 _1207_ (.A1(_0353_),
    .A2(_0356_),
    .Y(_0357_),
    .B1(_0333_));
 sg13g2_or3_1 _1208_ (.A(\pix_x[1] ),
    .B(_0349_),
    .C(_0357_),
    .X(_0358_));
 sg13g2_nor2_1 _1209_ (.A(net237),
    .B(_0332_),
    .Y(_0359_));
 sg13g2_nor3_1 _1210_ (.A(net219),
    .B(_0285_),
    .C(_0345_),
    .Y(_0360_));
 sg13g2_nor3_1 _1211_ (.A(_0208_),
    .B(_0288_),
    .C(_0345_),
    .Y(_0361_));
 sg13g2_nand3_1 _1212_ (.B(_0320_),
    .C(_0361_),
    .A(_0318_),
    .Y(_0362_));
 sg13g2_o21ai_1 _1213_ (.B1(net253),
    .Y(_0363_),
    .A1(net222),
    .A2(_0362_));
 sg13g2_nand3_1 _1214_ (.B(_0277_),
    .C(_0283_),
    .A(_0247_),
    .Y(_0364_));
 sg13g2_nand3_1 _1215_ (.B(_0320_),
    .C(_0364_),
    .A(_0318_),
    .Y(_0365_));
 sg13g2_a21oi_1 _1216_ (.A1(net239),
    .A2(_0365_),
    .Y(_0366_),
    .B1(net207));
 sg13g2_nor2_1 _1217_ (.A(net221),
    .B(_0346_),
    .Y(_0367_));
 sg13g2_nor3_1 _1218_ (.A(net221),
    .B(_0274_),
    .C(_0346_),
    .Y(_0368_));
 sg13g2_a221oi_1 _1219_ (.B2(_0273_),
    .C1(_0322_),
    .B1(_0367_),
    .A1(_0323_),
    .Y(_0369_),
    .A2(_0325_));
 sg13g2_a21o_1 _1220_ (.A2(_0366_),
    .A1(_0363_),
    .B1(_0369_),
    .X(_0370_));
 sg13g2_nand2_1 _1221_ (.Y(_0371_),
    .A(_0235_),
    .B(_0273_));
 sg13g2_nand2_1 _1222_ (.Y(_0372_),
    .A(_0247_),
    .B(_0273_));
 sg13g2_nor2_1 _1223_ (.A(_0288_),
    .B(_0372_),
    .Y(_0373_));
 sg13g2_nor3_1 _1224_ (.A(_0317_),
    .B(_0319_),
    .C(_0373_),
    .Y(_0374_));
 sg13g2_nor2_1 _1225_ (.A(net239),
    .B(_0374_),
    .Y(_0375_));
 sg13g2_or2_1 _1226_ (.X(_0376_),
    .B(_0345_),
    .A(net220));
 sg13g2_inv_1 _1227_ (.Y(_0377_),
    .A(_0376_));
 sg13g2_nor3_1 _1228_ (.A(net216),
    .B(_0285_),
    .C(_0376_),
    .Y(_0378_));
 sg13g2_nor3_2 _1229_ (.A(_0208_),
    .B(net221),
    .C(_0345_),
    .Y(_0379_));
 sg13g2_a21oi_1 _1230_ (.A1(_0321_),
    .A2(_0378_),
    .Y(_0380_),
    .B1(net252));
 sg13g2_o21ai_1 _1231_ (.B1(net207),
    .Y(_0381_),
    .A1(_0375_),
    .A2(_0380_));
 sg13g2_nor2_1 _1232_ (.A(net237),
    .B(net205),
    .Y(_0382_));
 sg13g2_a22oi_1 _1233_ (.Y(_0383_),
    .B1(_0368_),
    .B2(_0209_),
    .A2(_0351_),
    .A1(_0271_));
 sg13g2_a21oi_1 _1234_ (.A1(_0321_),
    .A2(_0383_),
    .Y(_0384_),
    .B1(net206));
 sg13g2_nor2b_1 _1235_ (.A(_0384_),
    .B_N(_0382_),
    .Y(_0385_));
 sg13g2_a221oi_1 _1236_ (.B2(_0385_),
    .C1(\pix_x[2] ),
    .B1(_0381_),
    .A1(_0359_),
    .Y(_0386_),
    .A2(_0370_));
 sg13g2_a21oi_1 _1237_ (.A1(_0028_),
    .A2(net217),
    .Y(_0387_),
    .B1(net222));
 sg13g2_o21ai_1 _1238_ (.B1(_0387_),
    .Y(_0388_),
    .A1(net217),
    .A2(_0292_));
 sg13g2_nand2_1 _1239_ (.Y(_0389_),
    .A(net222),
    .B(_0307_));
 sg13g2_nand3_1 _1240_ (.B(_0388_),
    .C(_0389_),
    .A(_0275_),
    .Y(_0390_));
 sg13g2_a21oi_1 _1241_ (.A1(_0276_),
    .A2(_0307_),
    .Y(_0391_),
    .B1(net218));
 sg13g2_a22oi_1 _1242_ (.Y(_0392_),
    .B1(_0390_),
    .B2(_0391_),
    .A2(_0307_),
    .A1(net218));
 sg13g2_nor2_1 _1243_ (.A(net218),
    .B(_0282_),
    .Y(_0393_));
 sg13g2_nor3_1 _1244_ (.A(net238),
    .B(net218),
    .C(_0282_),
    .Y(_0394_));
 sg13g2_nor2b_1 _1245_ (.A(_0376_),
    .B_N(_0394_),
    .Y(_0395_));
 sg13g2_nor4_1 _1246_ (.A(_0285_),
    .B(net205),
    .C(_0350_),
    .D(_0395_),
    .Y(_0396_));
 sg13g2_nor3_2 _1247_ (.A(net254),
    .B(net218),
    .C(_0282_),
    .Y(_0397_));
 sg13g2_nor3_1 _1248_ (.A(_0234_),
    .B(net216),
    .C(_0376_),
    .Y(_0398_));
 sg13g2_nand3_1 _1249_ (.B(_0269_),
    .C(_0379_),
    .A(_0235_),
    .Y(_0399_));
 sg13g2_nor3_1 _1250_ (.A(_0248_),
    .B(net216),
    .C(net220),
    .Y(_0400_));
 sg13g2_a221oi_1 _1251_ (.B2(_0394_),
    .C1(_0332_),
    .B1(_0400_),
    .A1(_0397_),
    .Y(_0401_),
    .A2(_0398_));
 sg13g2_o21ai_1 _1252_ (.B1(_0291_),
    .Y(_0402_),
    .A1(_0396_),
    .A2(_0401_));
 sg13g2_nand3_1 _1253_ (.B(_0279_),
    .C(_0283_),
    .A(_0269_),
    .Y(_0403_));
 sg13g2_nand2_1 _1254_ (.Y(_0404_),
    .A(net251),
    .B(_0286_));
 sg13g2_nand2_1 _1255_ (.Y(_0405_),
    .A(net238),
    .B(_0379_));
 sg13g2_nand2_1 _1256_ (.Y(_0406_),
    .A(_0404_),
    .B(_0405_));
 sg13g2_nand3_1 _1257_ (.B(_0273_),
    .C(_0379_),
    .A(_0235_),
    .Y(_0407_));
 sg13g2_and2_1 _1258_ (.A(net251),
    .B(_0407_),
    .X(_0408_));
 sg13g2_a21oi_1 _1259_ (.A1(net254),
    .A2(_0407_),
    .Y(_0409_),
    .B1(_0403_));
 sg13g2_nand3_1 _1260_ (.B(_0406_),
    .C(_0409_),
    .A(_0332_),
    .Y(_0410_));
 sg13g2_nor3_1 _1261_ (.A(net221),
    .B(_0282_),
    .C(_0284_),
    .Y(_0411_));
 sg13g2_nand3_1 _1262_ (.B(_0262_),
    .C(_0287_),
    .A(net251),
    .Y(_0412_));
 sg13g2_nor2_1 _1263_ (.A(_0372_),
    .B(_0412_),
    .Y(_0413_));
 sg13g2_nand4_1 _1264_ (.B(_0246_),
    .C(_0275_),
    .A(_0209_),
    .Y(_0414_),
    .D(_0393_));
 sg13g2_and2_1 _1265_ (.A(net240),
    .B(_0414_),
    .X(_0415_));
 sg13g2_or3_1 _1266_ (.A(_0332_),
    .B(_0413_),
    .C(_0415_),
    .X(_0416_));
 sg13g2_nand3_1 _1267_ (.B(_0410_),
    .C(_0416_),
    .A(net208),
    .Y(_0417_));
 sg13g2_a21o_1 _1268_ (.A2(_0417_),
    .A1(_0402_),
    .B1(net237),
    .X(_0418_));
 sg13g2_nor2_1 _1269_ (.A(\pix_x[1] ),
    .B(net206),
    .Y(_0419_));
 sg13g2_o21ai_1 _1270_ (.B1(_0377_),
    .Y(_0420_),
    .A1(net251),
    .A2(_0372_));
 sg13g2_nor3_1 _1271_ (.A(_0285_),
    .B(net205),
    .C(_0420_),
    .Y(_0421_));
 sg13g2_o21ai_1 _1272_ (.B1(net205),
    .Y(_0422_),
    .A1(net221),
    .A2(_0364_));
 sg13g2_a21oi_1 _1273_ (.A1(net238),
    .A2(_0365_),
    .Y(_0423_),
    .B1(_0422_));
 sg13g2_o21ai_1 _1274_ (.B1(_0419_),
    .Y(_0424_),
    .A1(_0421_),
    .A2(_0423_));
 sg13g2_a21o_1 _1275_ (.A2(_0424_),
    .A1(_0418_),
    .B1(_0322_),
    .X(_0425_));
 sg13g2_nor2_1 _1276_ (.A(_0350_),
    .B(_0371_),
    .Y(_0426_));
 sg13g2_a221oi_1 _1277_ (.B2(_0426_),
    .C1(_0322_),
    .B1(_0397_),
    .A1(net252),
    .Y(_0427_),
    .A2(_0373_));
 sg13g2_nand2b_1 _1278_ (.Y(_0428_),
    .B(_0332_),
    .A_N(_0427_));
 sg13g2_nand2_1 _1279_ (.Y(_0429_),
    .A(net237),
    .B(net207));
 sg13g2_nand3_1 _1280_ (.B(_0320_),
    .C(_0345_),
    .A(_0318_),
    .Y(_0430_));
 sg13g2_nand2_1 _1281_ (.Y(_0431_),
    .A(net253),
    .B(_0430_));
 sg13g2_mux2_1 _1282_ (.A0(_0362_),
    .A1(_0430_),
    .S(net252),
    .X(_0432_));
 sg13g2_a21oi_1 _1283_ (.A1(net205),
    .A2(_0432_),
    .Y(_0433_),
    .B1(_0429_));
 sg13g2_a21oi_1 _1284_ (.A1(_0428_),
    .A2(_0433_),
    .Y(_0434_),
    .B1(_0175_));
 sg13g2_a221oi_1 _1285_ (.B2(_0434_),
    .C1(_0392_),
    .B1(_0425_),
    .A1(_0358_),
    .Y(_0435_),
    .A2(_0386_));
 sg13g2_o21ai_1 _1286_ (.B1(net207),
    .Y(_0436_),
    .A1(net252),
    .A2(_0269_));
 sg13g2_and2_1 _1287_ (.A(_0277_),
    .B(_0334_),
    .X(_0437_));
 sg13g2_nor4_2 _1288_ (.A(net208),
    .B(_0317_),
    .C(_0319_),
    .Y(_0438_),
    .D(_0437_));
 sg13g2_and4_1 _1289_ (.A(net217),
    .B(_0262_),
    .C(_0277_),
    .D(_0286_),
    .X(_0439_));
 sg13g2_nand2b_1 _1290_ (.Y(_0440_),
    .B(_0438_),
    .A_N(_0439_));
 sg13g2_o21ai_1 _1291_ (.B1(_0440_),
    .Y(_0441_),
    .A1(_0432_),
    .A2(_0436_));
 sg13g2_nand4_1 _1292_ (.B(_0279_),
    .C(_0283_),
    .A(net251),
    .Y(_0442_),
    .D(_0286_));
 sg13g2_o21ai_1 _1293_ (.B1(_0442_),
    .Y(_0443_),
    .A1(_0264_),
    .A2(_0335_));
 sg13g2_nand2b_1 _1294_ (.Y(_0444_),
    .B(_0443_),
    .A_N(_0371_));
 sg13g2_nand3_1 _1295_ (.B(_0235_),
    .C(_0273_),
    .A(net238),
    .Y(_0445_));
 sg13g2_and4_1 _1296_ (.A(_0246_),
    .B(_0377_),
    .C(_0393_),
    .D(_0445_),
    .X(_0446_));
 sg13g2_mux2_1 _1297_ (.A0(_0444_),
    .A1(_0446_),
    .S(_0291_),
    .X(_0447_));
 sg13g2_o21ai_1 _1298_ (.B1(_0335_),
    .Y(_0448_),
    .A1(_0371_),
    .A2(_0442_));
 sg13g2_nand3_1 _1299_ (.B(_0379_),
    .C(_0448_),
    .A(_0332_),
    .Y(_0449_));
 sg13g2_nand4_1 _1300_ (.B(net217),
    .C(_0275_),
    .A(_0209_),
    .Y(_0450_),
    .D(_0286_));
 sg13g2_a22oi_1 _1301_ (.Y(_0451_),
    .B1(_0450_),
    .B2(net238),
    .A2(_0439_),
    .A1(_0394_));
 sg13g2_nand2_1 _1302_ (.Y(_0452_),
    .A(net205),
    .B(_0451_));
 sg13g2_nand4_1 _1303_ (.B(net208),
    .C(_0449_),
    .A(net237),
    .Y(_0453_),
    .D(_0452_));
 sg13g2_nor4_1 _1304_ (.A(_0248_),
    .B(net216),
    .C(net220),
    .D(_0404_),
    .Y(_0454_));
 sg13g2_a21oi_1 _1305_ (.A1(_0334_),
    .A2(_0398_),
    .Y(_0455_),
    .B1(_0454_));
 sg13g2_nand4_1 _1306_ (.B(_0263_),
    .C(_0269_),
    .A(_0246_),
    .Y(_0456_),
    .D(_0397_));
 sg13g2_o21ai_1 _1307_ (.B1(_0456_),
    .Y(_0457_),
    .A1(net238),
    .A2(_0360_));
 sg13g2_mux2_1 _1308_ (.A0(_0455_),
    .A1(_0457_),
    .S(_0332_),
    .X(_0458_));
 sg13g2_a22oi_1 _1309_ (.Y(_0459_),
    .B1(_0458_),
    .B2(_0419_),
    .A2(_0447_),
    .A1(_0382_));
 sg13g2_a21oi_1 _1310_ (.A1(_0453_),
    .A2(_0459_),
    .Y(_0460_),
    .B1(_0322_));
 sg13g2_a21o_1 _1311_ (.A2(_0441_),
    .A1(_0359_),
    .B1(_0460_),
    .X(_0461_));
 sg13g2_o21ai_1 _1312_ (.B1(net252),
    .Y(_0462_),
    .A1(_0288_),
    .A2(_0399_));
 sg13g2_nor3_1 _1313_ (.A(net221),
    .B(_0272_),
    .C(_0346_),
    .Y(_0463_));
 sg13g2_nor2_1 _1314_ (.A(_0322_),
    .B(_0463_),
    .Y(_0464_));
 sg13g2_a221oi_1 _1315_ (.B2(_0326_),
    .C1(\pix_x[1] ),
    .B1(_0464_),
    .A1(_0438_),
    .Y(_0465_),
    .A2(_0462_));
 sg13g2_nand4_1 _1316_ (.B(_0279_),
    .C(_0318_),
    .A(_0269_),
    .Y(_0466_),
    .D(_0426_));
 sg13g2_nor4_1 _1317_ (.A(_0282_),
    .B(_0285_),
    .C(net206),
    .D(_0466_),
    .Y(_0467_));
 sg13g2_a221oi_1 _1318_ (.B2(_0467_),
    .C1(net237),
    .B1(_0431_),
    .A1(_0181_),
    .Y(_0468_),
    .A2(_0324_));
 sg13g2_o21ai_1 _1319_ (.B1(net205),
    .Y(_0469_),
    .A1(_0465_),
    .A2(_0468_));
 sg13g2_nand2_1 _1320_ (.Y(_0470_),
    .A(net238),
    .B(_0430_));
 sg13g2_nand2_1 _1321_ (.Y(_0471_),
    .A(\pix_x[1] ),
    .B(net207));
 sg13g2_a21oi_1 _1322_ (.A1(net252),
    .A2(_0466_),
    .Y(_0472_),
    .B1(_0471_));
 sg13g2_o21ai_1 _1323_ (.B1(net252),
    .Y(_0473_),
    .A1(_0272_),
    .A2(_0288_));
 sg13g2_o21ai_1 _1324_ (.B1(_0473_),
    .Y(_0474_),
    .A1(_0345_),
    .A2(_0456_));
 sg13g2_nand3_1 _1325_ (.B(net206),
    .C(_0474_),
    .A(net237),
    .Y(_0475_));
 sg13g2_a22oi_1 _1326_ (.Y(_0476_),
    .B1(_0408_),
    .B2(net237),
    .A2(net216),
    .A1(net238));
 sg13g2_o21ai_1 _1327_ (.B1(_0475_),
    .Y(_0477_),
    .A1(net206),
    .A2(_0476_));
 sg13g2_a221oi_1 _1328_ (.B2(_0321_),
    .C1(net205),
    .B1(_0477_),
    .A1(_0470_),
    .Y(_0478_),
    .A2(_0472_));
 sg13g2_nor2_1 _1329_ (.A(_0175_),
    .B(_0478_),
    .Y(_0479_));
 sg13g2_a22oi_1 _1330_ (.Y(_0480_),
    .B1(_0469_),
    .B2(_0479_),
    .A2(_0461_),
    .A1(_0175_));
 sg13g2_o21ai_1 _1331_ (.B1(\pix_x[3] ),
    .Y(_0481_),
    .A1(_0392_),
    .A2(_0480_));
 sg13g2_or2_2 _1332_ (.X(_0482_),
    .B(_0435_),
    .A(\pix_x[3] ));
 sg13g2_nand3_1 _1333_ (.B(_0481_),
    .C(_0482_),
    .A(_0207_),
    .Y(_0483_));
 sg13g2_or3_1 _1334_ (.A(_0170_),
    .B(_0209_),
    .C(_0483_),
    .X(_0484_));
 sg13g2_and4_1 _1335_ (.A(net236),
    .B(net220),
    .C(_0481_),
    .D(_0482_),
    .X(_0485_));
 sg13g2_nand3_1 _1336_ (.B(_0481_),
    .C(_0482_),
    .A(_0189_),
    .Y(_0486_));
 sg13g2_and4_1 _1337_ (.A(_0189_),
    .B(_0270_),
    .C(_0481_),
    .D(_0482_),
    .X(_0487_));
 sg13g2_a22oi_1 _1338_ (.Y(_0488_),
    .B1(_0487_),
    .B2(net137),
    .A2(_0485_),
    .A1(net178));
 sg13g2_and4_1 _1339_ (.A(net236),
    .B(_0272_),
    .C(_0481_),
    .D(_0482_),
    .X(_0489_));
 sg13g2_nor3_1 _1340_ (.A(net262),
    .B(_0002_),
    .C(_0235_),
    .Y(_0490_));
 sg13g2_and3_1 _1341_ (.X(_0491_),
    .A(_0481_),
    .B(_0482_),
    .C(_0490_));
 sg13g2_a22oi_1 _1342_ (.Y(_0492_),
    .B1(_0491_),
    .B2(net139),
    .A2(_0489_),
    .A1(net135));
 sg13g2_nor2_1 _1343_ (.A(net263),
    .B(_0174_),
    .Y(_0493_));
 sg13g2_nor2b_1 _1344_ (.A(\pix_x[3] ),
    .B_N(net264),
    .Y(_0494_));
 sg13g2_a21o_1 _1345_ (.A2(_0493_),
    .A1(_0435_),
    .B1(_0494_),
    .X(_0495_));
 sg13g2_o21ai_1 _1346_ (.B1(_0174_),
    .Y(_0496_),
    .A1(_0392_),
    .A2(_0480_));
 sg13g2_and4_1 _1347_ (.A(_0021_),
    .B(_0344_),
    .C(_0495_),
    .D(_0496_),
    .X(_0497_));
 sg13g2_a21oi_1 _1348_ (.A1(_0017_),
    .A2(_0259_),
    .Y(_0498_),
    .B1(_0242_));
 sg13g2_nor2_1 _1349_ (.A(_0338_),
    .B(_0498_),
    .Y(_0499_));
 sg13g2_nor2_1 _1350_ (.A(_0230_),
    .B(_0237_),
    .Y(_0500_));
 sg13g2_a21oi_1 _1351_ (.A1(_0339_),
    .A2(_0500_),
    .Y(_0501_),
    .B1(_0259_));
 sg13g2_and2_1 _1352_ (.A(_0338_),
    .B(_0500_),
    .X(_0502_));
 sg13g2_nor4_1 _1353_ (.A(_0206_),
    .B(_0499_),
    .C(_0501_),
    .D(_0502_),
    .Y(_0503_));
 sg13g2_and4_1 _1354_ (.A(_0021_),
    .B(_0495_),
    .C(_0496_),
    .D(_0503_),
    .X(_0504_));
 sg13g2_a22oi_1 _1355_ (.Y(_0505_),
    .B1(_0504_),
    .B2(net143),
    .A2(_0497_),
    .A1(net149));
 sg13g2_nand4_1 _1356_ (.B(_0488_),
    .C(_0492_),
    .A(_0484_),
    .Y(_0506_),
    .D(_0505_));
 sg13g2_a21oi_1 _1357_ (.A1(_0209_),
    .A2(_0246_),
    .Y(_0507_),
    .B1(_0483_));
 sg13g2_nand4_1 _1358_ (.B(net219),
    .C(_0481_),
    .A(net236),
    .Y(_0508_),
    .D(_0482_));
 sg13g2_o21ai_1 _1359_ (.B1(_0508_),
    .Y(_0509_),
    .A1(_0411_),
    .A2(_0486_));
 sg13g2_nor2_1 _1360_ (.A(_0507_),
    .B(_0509_),
    .Y(_0510_));
 sg13g2_or2_1 _1361_ (.X(_0511_),
    .B(_0491_),
    .A(_0489_));
 sg13g2_or4_1 _1362_ (.A(_0485_),
    .B(_0487_),
    .C(_0497_),
    .D(_0504_),
    .X(_0512_));
 sg13g2_nor2_1 _1363_ (.A(_0511_),
    .B(_0512_),
    .Y(_0513_));
 sg13g2_nor4_1 _1364_ (.A(_0507_),
    .B(_0509_),
    .C(_0511_),
    .D(_0512_),
    .Y(_0514_));
 sg13g2_nand2_1 _1365_ (.Y(_0515_),
    .A(\driver.decoder.data_reg[1] ),
    .B(_0198_));
 sg13g2_nor3_1 _1366_ (.A(_0246_),
    .B(_0483_),
    .C(_0515_),
    .Y(_0516_));
 sg13g2_nand2_2 _1367_ (.Y(_0517_),
    .A(\driver.decoder.data_reg[7] ),
    .B(net231));
 sg13g2_nor2_1 _1368_ (.A(_0508_),
    .B(_0517_),
    .Y(_0518_));
 sg13g2_nand2_1 _1369_ (.Y(_0519_),
    .A(_0148_),
    .B(_0149_));
 sg13g2_a221oi_1 _1370_ (.B2(net257),
    .C1(net241),
    .B1(_0519_),
    .A1(_0184_),
    .Y(_0520_),
    .A2(_0297_));
 sg13g2_nand2_1 _1371_ (.Y(_0521_),
    .A(net271),
    .B(_0520_));
 sg13g2_nand3_1 _1372_ (.B(net231),
    .C(net221),
    .A(\driver.decoder.data_reg[2] ),
    .Y(_0522_));
 sg13g2_and2_1 _1373_ (.A(\driver.decoder.data_reg[5] ),
    .B(net231),
    .X(_0523_));
 sg13g2_and2_1 _1374_ (.A(\driver.decoder.data_reg[4] ),
    .B(net231),
    .X(_0524_));
 sg13g2_a22oi_1 _1375_ (.Y(_0525_),
    .B1(_0524_),
    .B2(_0284_),
    .A2(_0523_),
    .A1(_0282_));
 sg13g2_a21oi_1 _1376_ (.A1(_0522_),
    .A2(_0525_),
    .Y(_0526_),
    .B1(_0486_));
 sg13g2_or4_1 _1377_ (.A(_0516_),
    .B(_0518_),
    .C(_0521_),
    .D(_0526_),
    .X(_0527_));
 sg13g2_a221oi_1 _1378_ (.B2(_0513_),
    .C1(_0527_),
    .B1(_0510_),
    .A1(net231),
    .Y(_0034_),
    .A2(_0506_));
 sg13g2_nor2b_1 _1379_ (.A(\driver.driver.pmod_latch_prev ),
    .B_N(net110),
    .Y(_0528_));
 sg13g2_nor2_1 _1380_ (.A(_0171_),
    .B(net234),
    .Y(_0529_));
 sg13g2_a22oi_1 _1381_ (.Y(_0035_),
    .B1(net230),
    .B2(_0160_),
    .A2(net235),
    .A1(_0130_));
 sg13g2_a22oi_1 _1382_ (.Y(_0036_),
    .B1(net230),
    .B2(_0159_),
    .A2(net235),
    .A1(_0129_));
 sg13g2_a22oi_1 _1383_ (.Y(_0037_),
    .B1(net230),
    .B2(_0162_),
    .A2(net235),
    .A1(_0128_));
 sg13g2_a22oi_1 _1384_ (.Y(_0038_),
    .B1(net230),
    .B2(_0161_),
    .A2(net235),
    .A1(_0127_));
 sg13g2_a22oi_1 _1385_ (.Y(_0039_),
    .B1(net229),
    .B2(_0164_),
    .A2(net234),
    .A1(_0126_));
 sg13g2_a22oi_1 _1386_ (.Y(_0040_),
    .B1(net229),
    .B2(_0163_),
    .A2(net234),
    .A1(_0125_));
 sg13g2_a22oi_1 _1387_ (.Y(_0041_),
    .B1(net229),
    .B2(_0166_),
    .A2(net234),
    .A1(_0124_));
 sg13g2_a22oi_1 _1388_ (.Y(_0042_),
    .B1(net229),
    .B2(_0165_),
    .A2(net234),
    .A1(_0123_));
 sg13g2_a22oi_1 _1389_ (.Y(_0043_),
    .B1(net229),
    .B2(_0168_),
    .A2(net235),
    .A1(_0122_));
 sg13g2_a22oi_1 _1390_ (.Y(_0044_),
    .B1(net229),
    .B2(_0167_),
    .A2(net234),
    .A1(_0121_));
 sg13g2_a22oi_1 _1391_ (.Y(_0045_),
    .B1(net229),
    .B2(_0170_),
    .A2(net234),
    .A1(_0120_));
 sg13g2_a22oi_1 _1392_ (.Y(_0046_),
    .B1(net229),
    .B2(_0169_),
    .A2(net234),
    .A1(_0145_));
 sg13g2_and2_1 _1393_ (.A(net269),
    .B(net113),
    .X(_0047_));
 sg13g2_and2_1 _1394_ (.A(net183),
    .B(\counter[0] ),
    .X(_0530_));
 sg13g2_nor2_1 _1395_ (.A(net183),
    .B(\counter[0] ),
    .Y(_0531_));
 sg13g2_nor3_1 _1396_ (.A(net265),
    .B(_0530_),
    .C(net184),
    .Y(_0048_));
 sg13g2_nor2_1 _1397_ (.A(net166),
    .B(_0530_),
    .Y(_0532_));
 sg13g2_nand2_1 _1398_ (.Y(_0533_),
    .A(net166),
    .B(_0530_));
 sg13g2_nand2_1 _1399_ (.Y(_0534_),
    .A(net269),
    .B(_0533_));
 sg13g2_nor2_1 _1400_ (.A(net167),
    .B(_0534_),
    .Y(_0049_));
 sg13g2_and2_1 _1401_ (.A(_0146_),
    .B(_0533_),
    .X(_0535_));
 sg13g2_nor2_1 _1402_ (.A(_0146_),
    .B(_0533_),
    .Y(_0536_));
 sg13g2_nor3_1 _1403_ (.A(net265),
    .B(_0535_),
    .C(_0536_),
    .Y(_0050_));
 sg13g2_and2_1 _1404_ (.A(net196),
    .B(_0536_),
    .X(_0537_));
 sg13g2_o21ai_1 _1405_ (.B1(net270),
    .Y(_0538_),
    .A1(net196),
    .A2(_0536_));
 sg13g2_nor2_1 _1406_ (.A(_0537_),
    .B(net197),
    .Y(_0051_));
 sg13g2_xnor2_1 _1407_ (.Y(_0539_),
    .A(net186),
    .B(_0537_));
 sg13g2_nor2_1 _1408_ (.A(net265),
    .B(net187),
    .Y(_0052_));
 sg13g2_a21oi_1 _1409_ (.A1(\counter[5] ),
    .A2(_0537_),
    .Y(_0540_),
    .B1(net126));
 sg13g2_nand3_1 _1410_ (.B(net126),
    .C(_0537_),
    .A(net186),
    .Y(_0541_));
 sg13g2_nand2_1 _1411_ (.Y(_0542_),
    .A(net270),
    .B(_0541_));
 sg13g2_nor2_1 _1412_ (.A(net127),
    .B(_0542_),
    .Y(_0053_));
 sg13g2_and2_1 _1413_ (.A(_0147_),
    .B(_0541_),
    .X(_0543_));
 sg13g2_nor2_1 _1414_ (.A(_0147_),
    .B(_0541_),
    .Y(_0544_));
 sg13g2_nor3_1 _1415_ (.A(net265),
    .B(_0543_),
    .C(_0544_),
    .Y(_0054_));
 sg13g2_and2_1 _1416_ (.A(net192),
    .B(_0544_),
    .X(_0545_));
 sg13g2_o21ai_1 _1417_ (.B1(net269),
    .Y(_0546_),
    .A1(net192),
    .A2(_0544_));
 sg13g2_nor2_1 _1418_ (.A(_0545_),
    .B(net193),
    .Y(_0055_));
 sg13g2_xnor2_1 _1419_ (.Y(_0547_),
    .A(net188),
    .B(_0545_));
 sg13g2_nor2_1 _1420_ (.A(net265),
    .B(net189),
    .Y(_0056_));
 sg13g2_a21oi_1 _1421_ (.A1(\counter[9] ),
    .A2(_0545_),
    .Y(_0548_),
    .B1(net132));
 sg13g2_and3_1 _1422_ (.X(_0549_),
    .A(\counter[9] ),
    .B(net132),
    .C(_0545_));
 sg13g2_nor3_1 _1423_ (.A(net266),
    .B(net133),
    .C(_0549_),
    .Y(_0057_));
 sg13g2_xnor2_1 _1424_ (.Y(_0550_),
    .A(net179),
    .B(_0549_));
 sg13g2_nor2_1 _1425_ (.A(net266),
    .B(net180),
    .Y(_0058_));
 sg13g2_a21oi_1 _1426_ (.A1(\counter[11] ),
    .A2(_0549_),
    .Y(_0551_),
    .B1(net123));
 sg13g2_nand3_1 _1427_ (.B(net123),
    .C(_0549_),
    .A(\counter[11] ),
    .Y(_0552_));
 sg13g2_nand2_1 _1428_ (.Y(_0553_),
    .A(net268),
    .B(_0552_));
 sg13g2_nor2_1 _1429_ (.A(net124),
    .B(_0553_),
    .Y(_0059_));
 sg13g2_xor2_1 _1430_ (.B(_0552_),
    .A(net176),
    .X(_0554_));
 sg13g2_nor2_1 _1431_ (.A(net266),
    .B(net177),
    .Y(_0060_));
 sg13g2_nor2_2 _1432_ (.A(_0176_),
    .B(_0177_),
    .Y(_0555_));
 sg13g2_nor4_2 _1433_ (.A(_0174_),
    .B(_0175_),
    .C(_0176_),
    .Y(_0556_),
    .D(_0177_));
 sg13g2_nand3_1 _1434_ (.B(\pix_x[2] ),
    .C(_0555_),
    .A(\pix_x[3] ),
    .Y(_0557_));
 sg13g2_nand4_1 _1435_ (.B(net257),
    .C(_0500_),
    .A(net258),
    .Y(_0558_),
    .D(_0556_));
 sg13g2_and2_1 _1436_ (.A(net268),
    .B(_0558_),
    .X(_0559_));
 sg13g2_nand2_1 _1437_ (.Y(_0560_),
    .A(net268),
    .B(_0558_));
 sg13g2_and2_1 _1438_ (.A(net112),
    .B(_0559_),
    .X(_0061_));
 sg13g2_nor3_1 _1439_ (.A(_0171_),
    .B(net284),
    .C(_0555_),
    .Y(_0062_));
 sg13g2_o21ai_1 _1440_ (.B1(net271),
    .Y(_0561_),
    .A1(net285),
    .A2(_0555_));
 sg13g2_a21oi_1 _1441_ (.A1(net285),
    .A2(_0555_),
    .Y(_0063_),
    .B1(_0561_));
 sg13g2_nor2b_1 _1442_ (.A(net161),
    .B_N(_0555_),
    .Y(_0562_));
 sg13g2_xnor2_1 _1443_ (.Y(_0563_),
    .A(\pix_x[3] ),
    .B(_0562_));
 sg13g2_nor2_1 _1444_ (.A(_0560_),
    .B(net162),
    .Y(_0064_));
 sg13g2_xnor2_1 _1445_ (.Y(_0564_),
    .A(net129),
    .B(_0557_));
 sg13g2_nor2_1 _1446_ (.A(net214),
    .B(_0564_),
    .Y(_0065_));
 sg13g2_and3_1 _1447_ (.X(_0565_),
    .A(net262),
    .B(net263),
    .C(_0556_));
 sg13g2_a21oi_1 _1448_ (.A1(net263),
    .A2(_0556_),
    .Y(_0566_),
    .B1(net262));
 sg13g2_nor3_1 _1449_ (.A(net214),
    .B(_0565_),
    .C(net301),
    .Y(_0066_));
 sg13g2_nor2_1 _1450_ (.A(net261),
    .B(_0565_),
    .Y(_0567_));
 sg13g2_nor2_1 _1451_ (.A(_0192_),
    .B(_0557_),
    .Y(_0568_));
 sg13g2_nor3_1 _1452_ (.A(net214),
    .B(_0567_),
    .C(_0568_),
    .Y(_0067_));
 sg13g2_nor2_1 _1453_ (.A(net260),
    .B(_0568_),
    .Y(_0569_));
 sg13g2_nor3_2 _1454_ (.A(_0149_),
    .B(_0192_),
    .C(_0557_),
    .Y(_0570_));
 sg13g2_nor3_1 _1455_ (.A(net214),
    .B(net303),
    .C(_0570_),
    .Y(_0068_));
 sg13g2_and2_1 _1456_ (.A(net258),
    .B(_0570_),
    .X(_0571_));
 sg13g2_o21ai_1 _1457_ (.B1(net215),
    .Y(_0572_),
    .A1(net258),
    .A2(_0570_));
 sg13g2_nor2_1 _1458_ (.A(_0571_),
    .B(_0572_),
    .Y(_0069_));
 sg13g2_a21oi_1 _1459_ (.A1(net257),
    .A2(_0571_),
    .Y(_0573_),
    .B1(net214));
 sg13g2_o21ai_1 _1460_ (.B1(_0573_),
    .Y(_0574_),
    .A1(net257),
    .A2(_0571_));
 sg13g2_inv_1 _1461_ (.Y(_0070_),
    .A(_0574_));
 sg13g2_nor2_1 _1462_ (.A(\square_x[3] ),
    .B(_0174_),
    .Y(_0575_));
 sg13g2_a22oi_1 _1463_ (.Y(_0576_),
    .B1(_0177_),
    .B2(\square_x[1] ),
    .A2(_0176_),
    .A1(\square_x[0] ));
 sg13g2_a221oi_1 _1464_ (.B2(_0144_),
    .C1(_0576_),
    .B1(\pix_x[1] ),
    .A1(_0143_),
    .Y(_0577_),
    .A2(\pix_x[2] ));
 sg13g2_a221oi_1 _1465_ (.B2(\square_x[2] ),
    .C1(_0577_),
    .B1(_0175_),
    .A1(\square_x[3] ),
    .Y(_0578_),
    .A2(_0174_));
 sg13g2_or2_1 _1466_ (.X(_0579_),
    .B(_0578_),
    .A(_0575_));
 sg13g2_a21oi_1 _1467_ (.A1(net256),
    .A2(net264),
    .Y(_0580_),
    .B1(_0579_));
 sg13g2_nand2_1 _1468_ (.Y(_0581_),
    .A(\square_x[5] ),
    .B(net256));
 sg13g2_xnor2_1 _1469_ (.Y(_0582_),
    .A(\square_x[5] ),
    .B(net256));
 sg13g2_nor2_1 _1470_ (.A(net256),
    .B(net264),
    .Y(_0583_));
 sg13g2_xor2_1 _1471_ (.B(_0582_),
    .A(_0021_),
    .X(_0584_));
 sg13g2_nor3_1 _1472_ (.A(_0580_),
    .B(_0583_),
    .C(_0584_),
    .Y(_0585_));
 sg13g2_a21o_1 _1473_ (.A2(_0582_),
    .A1(net262),
    .B1(_0585_),
    .X(_0586_));
 sg13g2_nor2_1 _1474_ (.A(_0005_),
    .B(_0581_),
    .Y(_0587_));
 sg13g2_xnor2_1 _1475_ (.Y(_0588_),
    .A(_0005_),
    .B(_0581_));
 sg13g2_o21ai_1 _1476_ (.B1(_0586_),
    .Y(_0589_),
    .A1(net261),
    .A2(_0588_));
 sg13g2_xor2_1 _1477_ (.B(_0587_),
    .A(_0016_),
    .X(_0590_));
 sg13g2_a22oi_1 _1478_ (.Y(_0591_),
    .B1(_0590_),
    .B2(net260),
    .A2(_0588_),
    .A1(net261));
 sg13g2_nand4_1 _1479_ (.B(\square_x[6] ),
    .C(\square_x[5] ),
    .A(\square_x[7] ),
    .Y(_0592_),
    .D(net256));
 sg13g2_nor2_1 _1480_ (.A(_0004_),
    .B(_0592_),
    .Y(_0593_));
 sg13g2_xor2_1 _1481_ (.B(_0592_),
    .A(_0004_),
    .X(_0594_));
 sg13g2_a22oi_1 _1482_ (.Y(_0595_),
    .B1(_0594_),
    .B2(_0148_),
    .A2(_0591_),
    .A1(_0589_));
 sg13g2_o21ai_1 _1483_ (.B1(_0595_),
    .Y(_0596_),
    .A1(net260),
    .A2(_0590_));
 sg13g2_nand2b_1 _1484_ (.Y(_0597_),
    .B(net258),
    .A_N(_0594_));
 sg13g2_xnor2_1 _1485_ (.Y(_0598_),
    .A(_0003_),
    .B(_0593_));
 sg13g2_o21ai_1 _1486_ (.B1(_0597_),
    .Y(_0599_),
    .A1(_0150_),
    .A2(_0598_));
 sg13g2_nand2b_1 _1487_ (.Y(_0600_),
    .B(_0596_),
    .A_N(_0599_));
 sg13g2_nor2_1 _1488_ (.A(_0141_),
    .B(_0592_),
    .Y(_0601_));
 sg13g2_a22oi_1 _1489_ (.Y(_0602_),
    .B1(_0601_),
    .B2(\square_x[9] ),
    .A2(_0598_),
    .A1(_0150_));
 sg13g2_nand2_1 _1490_ (.Y(_0603_),
    .A(\square_y[5] ),
    .B(\square_y[4] ));
 sg13g2_nor2_1 _1491_ (.A(\square_y[5] ),
    .B(\square_y[4] ),
    .Y(_0604_));
 sg13g2_xnor2_1 _1492_ (.Y(_0605_),
    .A(\square_y[5] ),
    .B(\square_y[4] ));
 sg13g2_nand2_1 _1493_ (.Y(_0606_),
    .A(\square_y[3] ),
    .B(_0156_));
 sg13g2_nor2_1 _1494_ (.A(\square_y[1] ),
    .B(net240),
    .Y(_0607_));
 sg13g2_nor3_1 _1495_ (.A(_0138_),
    .B(\pix_y[0] ),
    .C(_0607_),
    .Y(_0608_));
 sg13g2_a221oi_1 _1496_ (.B2(\square_y[1] ),
    .C1(_0608_),
    .B1(net240),
    .A1(\square_y[2] ),
    .Y(_0609_),
    .A2(_0157_));
 sg13g2_nand2b_1 _1497_ (.Y(_0610_),
    .B(net249),
    .A_N(\square_y[3] ));
 sg13g2_o21ai_1 _1498_ (.B1(_0610_),
    .Y(_0611_),
    .A1(\square_y[2] ),
    .A2(_0157_));
 sg13g2_o21ai_1 _1499_ (.B1(_0606_),
    .Y(_0612_),
    .A1(_0609_),
    .A2(_0611_));
 sg13g2_nand2_1 _1500_ (.Y(_0613_),
    .A(\square_y[4] ),
    .B(net246));
 sg13g2_nand2_1 _1501_ (.Y(_0614_),
    .A(_0137_),
    .B(_0155_));
 sg13g2_o21ai_1 _1502_ (.B1(_0614_),
    .Y(_0615_),
    .A1(_0178_),
    .A2(_0605_));
 sg13g2_a221oi_1 _1503_ (.B2(_0613_),
    .C1(_0615_),
    .B1(_0612_),
    .A1(_0178_),
    .Y(_0616_),
    .A2(_0605_));
 sg13g2_a21oi_1 _1504_ (.A1(net244),
    .A2(_0605_),
    .Y(_0617_),
    .B1(_0616_));
 sg13g2_nor2_1 _1505_ (.A(_0009_),
    .B(_0603_),
    .Y(_0618_));
 sg13g2_xor2_1 _1506_ (.B(_0603_),
    .A(_0009_),
    .X(_0619_));
 sg13g2_xnor2_1 _1507_ (.Y(_0620_),
    .A(_0023_),
    .B(_0619_));
 sg13g2_xor2_1 _1508_ (.B(_0618_),
    .A(_0008_),
    .X(_0621_));
 sg13g2_nor2_1 _1509_ (.A(_0152_),
    .B(_0619_),
    .Y(_0622_));
 sg13g2_a21oi_1 _1510_ (.A1(net243),
    .A2(_0621_),
    .Y(_0623_),
    .B1(_0622_));
 sg13g2_o21ai_1 _1511_ (.B1(_0623_),
    .Y(_0624_),
    .A1(_0617_),
    .A2(_0620_));
 sg13g2_nand4_1 _1512_ (.B(\square_y[6] ),
    .C(\square_y[5] ),
    .A(\square_y[7] ),
    .Y(_0625_),
    .D(\square_y[4] ));
 sg13g2_nor2_1 _1513_ (.A(_0007_),
    .B(_0625_),
    .Y(_0626_));
 sg13g2_xor2_1 _1514_ (.B(_0625_),
    .A(_0007_),
    .X(_0627_));
 sg13g2_xnor2_1 _1515_ (.Y(_0628_),
    .A(_0024_),
    .B(_0627_));
 sg13g2_o21ai_1 _1516_ (.B1(_0624_),
    .Y(_0629_),
    .A1(net243),
    .A2(_0621_));
 sg13g2_nor2_1 _1517_ (.A(_0151_),
    .B(_0627_),
    .Y(_0630_));
 sg13g2_xor2_1 _1518_ (.B(_0626_),
    .A(_0006_),
    .X(_0631_));
 sg13g2_a21oi_1 _1519_ (.A1(\pix_y[9] ),
    .A2(_0631_),
    .Y(_0632_),
    .B1(_0630_));
 sg13g2_o21ai_1 _1520_ (.B1(_0632_),
    .Y(_0633_),
    .A1(_0628_),
    .A2(_0629_));
 sg13g2_nor2_1 _1521_ (.A(net241),
    .B(_0631_),
    .Y(_0634_));
 sg13g2_nand2_1 _1522_ (.Y(_0635_),
    .A(\square_y[9] ),
    .B(\square_y[8] ));
 sg13g2_o21ai_1 _1523_ (.B1(_0633_),
    .Y(_0636_),
    .A1(_0625_),
    .A2(_0635_));
 sg13g2_nand2b_1 _1524_ (.Y(_0637_),
    .B(net256),
    .A_N(net264));
 sg13g2_nor2b_1 _1525_ (.A(net256),
    .B_N(net264),
    .Y(_0638_));
 sg13g2_o21ai_1 _1526_ (.B1(_0637_),
    .Y(_0639_),
    .A1(_0579_),
    .A2(_0638_));
 sg13g2_o21ai_1 _1527_ (.B1(_0639_),
    .Y(_0640_),
    .A1(\square_x[5] ),
    .A2(_0173_));
 sg13g2_a22oi_1 _1528_ (.Y(_0641_),
    .B1(_0173_),
    .B2(\square_x[5] ),
    .A2(_0172_),
    .A1(\square_x[6] ));
 sg13g2_nor2_1 _1529_ (.A(\square_x[6] ),
    .B(_0172_),
    .Y(_0642_));
 sg13g2_a221oi_1 _1530_ (.B2(_0641_),
    .C1(_0642_),
    .B1(_0640_),
    .A1(_0142_),
    .Y(_0643_),
    .A2(net260));
 sg13g2_a221oi_1 _1531_ (.B2(\square_x[7] ),
    .C1(_0643_),
    .B1(_0149_),
    .A1(\square_x[8] ),
    .Y(_0644_),
    .A2(_0148_));
 sg13g2_a221oi_1 _1532_ (.B2(_0140_),
    .C1(_0644_),
    .B1(net257),
    .A1(_0141_),
    .Y(_0645_),
    .A2(net258));
 sg13g2_a21oi_1 _1533_ (.A1(_0613_),
    .A2(_0614_),
    .Y(_0646_),
    .B1(_0612_));
 sg13g2_a221oi_1 _1534_ (.B2(_0137_),
    .C1(_0646_),
    .B1(net246),
    .A1(_0136_),
    .Y(_0647_),
    .A2(net245));
 sg13g2_a221oi_1 _1535_ (.B2(\square_y[5] ),
    .C1(_0647_),
    .B1(_0154_),
    .A1(\square_y[6] ),
    .Y(_0648_),
    .A2(_0152_));
 sg13g2_a221oi_1 _1536_ (.B2(_0134_),
    .C1(_0648_),
    .B1(\pix_y[7] ),
    .A1(_0135_),
    .Y(_0649_),
    .A2(\pix_y[6] ));
 sg13g2_a221oi_1 _1537_ (.B2(\square_y[7] ),
    .C1(_0649_),
    .B1(_0153_),
    .A1(\square_y[8] ),
    .Y(_0650_),
    .A2(_0151_));
 sg13g2_a221oi_1 _1538_ (.B2(_0133_),
    .C1(_0650_),
    .B1(net242),
    .A1(_0132_),
    .Y(_0651_),
    .A2(net241));
 sg13g2_nor2_1 _1539_ (.A(_0140_),
    .B(net257),
    .Y(_0652_));
 sg13g2_nor2_1 _1540_ (.A(_0132_),
    .B(net241),
    .Y(_0653_));
 sg13g2_nor4_1 _1541_ (.A(_0645_),
    .B(_0651_),
    .C(_0652_),
    .D(_0653_),
    .Y(_0654_));
 sg13g2_o21ai_1 _1542_ (.B1(_0654_),
    .Y(_0655_),
    .A1(_0634_),
    .A2(_0636_));
 sg13g2_a21o_1 _1543_ (.A2(_0602_),
    .A1(_0600_),
    .B1(_0655_),
    .X(_0656_));
 sg13g2_a21oi_1 _1544_ (.A1(_0514_),
    .A2(_0656_),
    .Y(_0071_),
    .B1(_0521_));
 sg13g2_nor4_1 _1545_ (.A(\square_x[3] ),
    .B(\square_x[2] ),
    .C(\square_x[1] ),
    .D(\square_x[0] ),
    .Y(_0657_));
 sg13g2_nor4_1 _1546_ (.A(\square_x[9] ),
    .B(\square_x[6] ),
    .C(\square_x[5] ),
    .D(net256),
    .Y(_0658_));
 sg13g2_nand4_1 _1547_ (.B(_0142_),
    .C(_0657_),
    .A(_0141_),
    .Y(_0659_),
    .D(_0658_));
 sg13g2_and3_1 _1548_ (.X(_0660_),
    .A(\driver.decoder.data_reg[5] ),
    .B(net231),
    .C(_0659_));
 sg13g2_nand2_2 _1549_ (.Y(_0661_),
    .A(_0523_),
    .B(_0659_));
 sg13g2_nand2_1 _1550_ (.Y(_0662_),
    .A(_0142_),
    .B(\square_x[6] ));
 sg13g2_o21ai_1 _1551_ (.B1(_0016_),
    .Y(_0663_),
    .A1(_0581_),
    .A2(_0662_));
 sg13g2_o21ai_1 _1552_ (.B1(\square_x[9] ),
    .Y(_0664_),
    .A1(\square_x[8] ),
    .A2(_0663_));
 sg13g2_nand2_1 _1553_ (.Y(_0665_),
    .A(_0524_),
    .B(_0664_));
 sg13g2_nor4_1 _1554_ (.A(\counter[3] ),
    .B(\counter[2] ),
    .C(\counter[5] ),
    .D(\counter[4] ),
    .Y(_0666_));
 sg13g2_nor4_1 _1555_ (.A(\counter[11] ),
    .B(\counter[10] ),
    .C(\counter[13] ),
    .D(\counter[12] ),
    .Y(_0667_));
 sg13g2_nor4_1 _1556_ (.A(\counter[7] ),
    .B(\counter[6] ),
    .C(\counter[9] ),
    .D(\counter[8] ),
    .Y(_0668_));
 sg13g2_nand4_1 _1557_ (.B(_0666_),
    .C(_0667_),
    .A(_0531_),
    .Y(_0669_),
    .D(_0668_));
 sg13g2_or2_1 _1558_ (.X(_0670_),
    .B(_0669_),
    .A(_0520_));
 sg13g2_a221oi_1 _1559_ (.B2(_0665_),
    .C1(_0670_),
    .B1(_0661_),
    .A1(\driver.decoder.data_reg[5] ),
    .Y(_0671_),
    .A2(net175));
 sg13g2_nor2_1 _1560_ (.A(\square_x[0] ),
    .B(net212),
    .Y(_0672_));
 sg13g2_nor2b_1 _1561_ (.A(net121),
    .B_N(net212),
    .Y(_0673_));
 sg13g2_nor3_1 _1562_ (.A(net266),
    .B(_0672_),
    .C(_0673_),
    .Y(_0072_));
 sg13g2_o21ai_1 _1563_ (.B1(net269),
    .Y(_0674_),
    .A1(net272),
    .A2(net212));
 sg13g2_nor2_1 _1564_ (.A(_0182_),
    .B(net226),
    .Y(_0675_));
 sg13g2_xnor2_1 _1565_ (.Y(_0676_),
    .A(_0013_),
    .B(net226));
 sg13g2_or2_1 _1566_ (.X(_0677_),
    .B(_0676_),
    .A(net121));
 sg13g2_nand2_1 _1567_ (.Y(_0678_),
    .A(net121),
    .B(_0676_));
 sg13g2_and3_1 _1568_ (.X(_0679_),
    .A(net212),
    .B(_0677_),
    .C(_0678_));
 sg13g2_nor2_1 _1569_ (.A(_0674_),
    .B(_0679_),
    .Y(_0073_));
 sg13g2_xnor2_1 _1570_ (.Y(_0680_),
    .A(\square_x[2] ),
    .B(net226));
 sg13g2_a21oi_1 _1571_ (.A1(_0182_),
    .A2(net226),
    .Y(_0681_),
    .B1(\square_x[0] ));
 sg13g2_or3_1 _1572_ (.A(_0675_),
    .B(_0680_),
    .C(_0681_),
    .X(_0682_));
 sg13g2_o21ai_1 _1573_ (.B1(_0680_),
    .Y(_0683_),
    .A1(_0675_),
    .A2(_0681_));
 sg13g2_and2_1 _1574_ (.A(_0682_),
    .B(_0683_),
    .X(_0684_));
 sg13g2_mux2_1 _1575_ (.A0(net310),
    .A1(_0684_),
    .S(net212),
    .X(_0685_));
 sg13g2_and2_1 _1576_ (.A(net269),
    .B(_0685_),
    .X(_0074_));
 sg13g2_o21ai_1 _1577_ (.B1(_0682_),
    .Y(_0686_),
    .A1(_0143_),
    .A2(_0661_));
 sg13g2_nor2_1 _1578_ (.A(_0014_),
    .B(_0661_),
    .Y(_0687_));
 sg13g2_nand2_1 _1579_ (.Y(_0688_),
    .A(_0014_),
    .B(_0661_));
 sg13g2_nand2b_1 _1580_ (.Y(_0689_),
    .B(_0688_),
    .A_N(_0687_));
 sg13g2_xnor2_1 _1581_ (.Y(_0690_),
    .A(_0686_),
    .B(_0689_));
 sg13g2_mux2_1 _1582_ (.A0(net288),
    .A1(_0690_),
    .S(net212),
    .X(_0691_));
 sg13g2_and2_1 _1583_ (.A(net269),
    .B(_0691_),
    .X(_0075_));
 sg13g2_nand2_1 _1584_ (.Y(_0692_),
    .A(\square_x[4] ),
    .B(net226));
 sg13g2_xnor2_1 _1585_ (.Y(_0693_),
    .A(\square_x[4] ),
    .B(net225));
 sg13g2_a21oi_1 _1586_ (.A1(_0686_),
    .A2(_0688_),
    .Y(_0694_),
    .B1(_0687_));
 sg13g2_xnor2_1 _1587_ (.Y(_0695_),
    .A(_0693_),
    .B(_0694_));
 sg13g2_nand2_1 _1588_ (.Y(_0696_),
    .A(net213),
    .B(_0695_));
 sg13g2_o21ai_1 _1589_ (.B1(_0696_),
    .Y(_0697_),
    .A1(net200),
    .A2(_0671_));
 sg13g2_nor2_1 _1590_ (.A(net265),
    .B(net201),
    .Y(_0076_));
 sg13g2_o21ai_1 _1591_ (.B1(_0692_),
    .Y(_0698_),
    .A1(_0693_),
    .A2(_0694_));
 sg13g2_nand2_1 _1592_ (.Y(_0699_),
    .A(_0015_),
    .B(_0661_));
 sg13g2_nor2_1 _1593_ (.A(_0015_),
    .B(_0661_),
    .Y(_0700_));
 sg13g2_xnor2_1 _1594_ (.Y(_0701_),
    .A(_0015_),
    .B(net225));
 sg13g2_xnor2_1 _1595_ (.Y(_0702_),
    .A(_0698_),
    .B(_0701_));
 sg13g2_nand2_1 _1596_ (.Y(_0703_),
    .A(net212),
    .B(_0702_));
 sg13g2_o21ai_1 _1597_ (.B1(_0703_),
    .Y(_0704_),
    .A1(net291),
    .A2(net212));
 sg13g2_nor2_1 _1598_ (.A(net265),
    .B(_0704_),
    .Y(_0077_));
 sg13g2_a21o_1 _1599_ (.A2(_0699_),
    .A1(_0698_),
    .B1(_0700_),
    .X(_0705_));
 sg13g2_xnor2_1 _1600_ (.Y(_0706_),
    .A(_0005_),
    .B(net225));
 sg13g2_xor2_1 _1601_ (.B(_0706_),
    .A(_0705_),
    .X(_0707_));
 sg13g2_mux2_1 _1602_ (.A0(net313),
    .A1(_0707_),
    .S(net213),
    .X(_0708_));
 sg13g2_and2_1 _1603_ (.A(net269),
    .B(_0708_),
    .X(_0078_));
 sg13g2_and2_1 _1604_ (.A(\square_x[6] ),
    .B(net225),
    .X(_0709_));
 sg13g2_a21o_1 _1605_ (.A2(_0706_),
    .A1(_0705_),
    .B1(_0709_),
    .X(_0710_));
 sg13g2_xnor2_1 _1606_ (.Y(_0711_),
    .A(_0016_),
    .B(net225));
 sg13g2_and2_1 _1607_ (.A(_0710_),
    .B(_0711_),
    .X(_0712_));
 sg13g2_nor2_1 _1608_ (.A(_0710_),
    .B(_0711_),
    .Y(_0713_));
 sg13g2_o21ai_1 _1609_ (.B1(net213),
    .Y(_0714_),
    .A1(_0712_),
    .A2(_0713_));
 sg13g2_o21ai_1 _1610_ (.B1(_0714_),
    .Y(_0715_),
    .A1(net275),
    .A2(net213));
 sg13g2_nor2_1 _1611_ (.A(net266),
    .B(_0715_),
    .Y(_0079_));
 sg13g2_a21oi_1 _1612_ (.A1(\square_x[7] ),
    .A2(net225),
    .Y(_0716_),
    .B1(_0712_));
 sg13g2_nor2_1 _1613_ (.A(_0004_),
    .B(net225),
    .Y(_0717_));
 sg13g2_xnor2_1 _1614_ (.Y(_0718_),
    .A(_0004_),
    .B(net225));
 sg13g2_nand2b_1 _1615_ (.Y(_0719_),
    .B(_0718_),
    .A_N(_0716_));
 sg13g2_xnor2_1 _1616_ (.Y(_0720_),
    .A(_0716_),
    .B(_0718_));
 sg13g2_mux2_1 _1617_ (.A0(net308),
    .A1(_0720_),
    .S(net213),
    .X(_0721_));
 sg13g2_and2_1 _1618_ (.A(net268),
    .B(_0721_),
    .X(_0080_));
 sg13g2_nor2_1 _1619_ (.A(net198),
    .B(net213),
    .Y(_0722_));
 sg13g2_nor2_1 _1620_ (.A(\square_x[8] ),
    .B(_0661_),
    .Y(_0723_));
 sg13g2_a22oi_1 _1621_ (.Y(_0724_),
    .B1(_0719_),
    .B2(_0723_),
    .A2(_0717_),
    .A1(_0712_));
 sg13g2_nand2b_1 _1622_ (.Y(_0725_),
    .B(_0003_),
    .A_N(_0724_));
 sg13g2_nand2b_1 _1623_ (.Y(_0726_),
    .B(_0724_),
    .A_N(_0003_));
 sg13g2_and3_1 _1624_ (.X(_0727_),
    .A(net213),
    .B(_0725_),
    .C(_0726_));
 sg13g2_nor3_1 _1625_ (.A(net266),
    .B(_0722_),
    .C(_0727_),
    .Y(_0081_));
 sg13g2_nor4_1 _1626_ (.A(\square_y[3] ),
    .B(\square_y[2] ),
    .C(\square_y[1] ),
    .D(\square_y[0] ),
    .Y(_0728_));
 sg13g2_nor4_1 _1627_ (.A(\square_y[9] ),
    .B(\square_y[8] ),
    .C(\square_y[7] ),
    .D(\square_y[6] ),
    .Y(_0729_));
 sg13g2_nand3_1 _1628_ (.B(_0728_),
    .C(_0729_),
    .A(_0604_),
    .Y(_0730_));
 sg13g2_nand3_1 _1629_ (.B(net231),
    .C(_0730_),
    .A(\driver.decoder.data_reg[7] ),
    .Y(_0731_));
 sg13g2_inv_1 _1630_ (.Y(_0732_),
    .A(net224));
 sg13g2_nor4_1 _1631_ (.A(_0133_),
    .B(_0134_),
    .C(_0135_),
    .D(_0604_),
    .Y(_0733_));
 sg13g2_nor3_1 _1632_ (.A(\square_y[9] ),
    .B(_0166_),
    .C(_0733_),
    .Y(_0734_));
 sg13g2_a21oi_1 _1633_ (.A1(net231),
    .A2(_0734_),
    .Y(_0735_),
    .B1(_0732_));
 sg13g2_nor3_1 _1634_ (.A(_0196_),
    .B(_0670_),
    .C(_0735_),
    .Y(_0736_));
 sg13g2_nor3_1 _1635_ (.A(_0196_),
    .B(_0670_),
    .C(_0735_),
    .Y(_0737_));
 sg13g2_inv_1 _1636_ (.Y(_0738_),
    .A(_0737_));
 sg13g2_o21ai_1 _1637_ (.B1(net267),
    .Y(_0739_),
    .A1(\square_y[0] ),
    .A2(net211));
 sg13g2_a21oi_1 _1638_ (.A1(_0139_),
    .A2(net211),
    .Y(_0082_),
    .B1(_0739_));
 sg13g2_o21ai_1 _1639_ (.B1(net267),
    .Y(_0740_),
    .A1(net151),
    .A2(net211));
 sg13g2_nor2_1 _1640_ (.A(_0010_),
    .B(net224),
    .Y(_0741_));
 sg13g2_nand2_1 _1641_ (.Y(_0742_),
    .A(_0010_),
    .B(net224));
 sg13g2_nor2b_1 _1642_ (.A(_0741_),
    .B_N(_0742_),
    .Y(_0743_));
 sg13g2_or2_1 _1643_ (.X(_0744_),
    .B(_0743_),
    .A(net119));
 sg13g2_a21oi_1 _1644_ (.A1(net119),
    .A2(_0743_),
    .Y(_0745_),
    .B1(_0738_));
 sg13g2_a21oi_1 _1645_ (.A1(_0744_),
    .A2(_0745_),
    .Y(_0083_),
    .B1(_0740_));
 sg13g2_nand2_1 _1646_ (.Y(_0746_),
    .A(\square_y[2] ),
    .B(_0732_));
 sg13g2_xor2_1 _1647_ (.B(net224),
    .A(\square_y[2] ),
    .X(_0747_));
 sg13g2_o21ai_1 _1648_ (.B1(_0742_),
    .Y(_0748_),
    .A1(\square_y[0] ),
    .A2(_0741_));
 sg13g2_xnor2_1 _1649_ (.Y(_0749_),
    .A(_0747_),
    .B(_0748_));
 sg13g2_o21ai_1 _1650_ (.B1(net267),
    .Y(_0750_),
    .A1(net286),
    .A2(net209));
 sg13g2_a21oi_1 _1651_ (.A1(net209),
    .A2(_0749_),
    .Y(_0084_),
    .B1(_0750_));
 sg13g2_nor2_1 _1652_ (.A(net190),
    .B(net211),
    .Y(_0751_));
 sg13g2_o21ai_1 _1653_ (.B1(_0746_),
    .Y(_0752_),
    .A1(_0747_),
    .A2(_0748_));
 sg13g2_nor2_1 _1654_ (.A(_0011_),
    .B(net224),
    .Y(_0753_));
 sg13g2_nand2_1 _1655_ (.Y(_0754_),
    .A(_0011_),
    .B(net224));
 sg13g2_nand2b_1 _1656_ (.Y(_0755_),
    .B(_0754_),
    .A_N(_0753_));
 sg13g2_xnor2_1 _1657_ (.Y(_0756_),
    .A(_0752_),
    .B(_0755_));
 sg13g2_nor2_1 _1658_ (.A(_0738_),
    .B(_0756_),
    .Y(_0757_));
 sg13g2_nor3_1 _1659_ (.A(net266),
    .B(_0751_),
    .C(_0757_),
    .Y(_0085_));
 sg13g2_nand2_1 _1660_ (.Y(_0758_),
    .A(\square_y[4] ),
    .B(_0732_));
 sg13g2_xnor2_1 _1661_ (.Y(_0759_),
    .A(_0137_),
    .B(net223));
 sg13g2_a21oi_2 _1662_ (.B1(_0753_),
    .Y(_0760_),
    .A2(_0754_),
    .A1(_0752_));
 sg13g2_xnor2_1 _1663_ (.Y(_0761_),
    .A(_0759_),
    .B(_0760_));
 sg13g2_o21ai_1 _1664_ (.B1(net267),
    .Y(_0762_),
    .A1(net297),
    .A2(net209));
 sg13g2_a21oi_1 _1665_ (.A1(net209),
    .A2(_0761_),
    .Y(_0086_),
    .B1(_0762_));
 sg13g2_o21ai_1 _1666_ (.B1(net267),
    .Y(_0763_),
    .A1(\square_y[5] ),
    .A2(net209));
 sg13g2_o21ai_1 _1667_ (.B1(_0758_),
    .Y(_0764_),
    .A1(_0759_),
    .A2(_0760_));
 sg13g2_nand2_1 _1668_ (.Y(_0765_),
    .A(_0012_),
    .B(net223));
 sg13g2_nor2_1 _1669_ (.A(_0012_),
    .B(net223),
    .Y(_0766_));
 sg13g2_xor2_1 _1670_ (.B(net223),
    .A(net295),
    .X(_0767_));
 sg13g2_xnor2_1 _1671_ (.Y(_0768_),
    .A(_0764_),
    .B(_0767_));
 sg13g2_a21oi_1 _1672_ (.A1(net209),
    .A2(_0768_),
    .Y(_0087_),
    .B1(_0763_));
 sg13g2_o21ai_1 _1673_ (.B1(_0765_),
    .Y(_0769_),
    .A1(_0764_),
    .A2(_0766_));
 sg13g2_xor2_1 _1674_ (.B(net223),
    .A(_0009_),
    .X(_0770_));
 sg13g2_nand2b_1 _1675_ (.Y(_0771_),
    .B(_0770_),
    .A_N(_0769_));
 sg13g2_xor2_1 _1676_ (.B(_0770_),
    .A(_0769_),
    .X(_0772_));
 sg13g2_o21ai_1 _1677_ (.B1(net267),
    .Y(_0773_),
    .A1(net277),
    .A2(net210));
 sg13g2_a21oi_1 _1678_ (.A1(net209),
    .A2(_0772_),
    .Y(_0088_),
    .B1(_0773_));
 sg13g2_o21ai_1 _1679_ (.B1(_0771_),
    .Y(_0774_),
    .A1(_0135_),
    .A2(net223));
 sg13g2_xor2_1 _1680_ (.B(net223),
    .A(_0008_),
    .X(_0775_));
 sg13g2_xnor2_1 _1681_ (.Y(_0776_),
    .A(_0774_),
    .B(_0775_));
 sg13g2_o21ai_1 _1682_ (.B1(net268),
    .Y(_0777_),
    .A1(net279),
    .A2(net210));
 sg13g2_a21oi_1 _1683_ (.A1(net210),
    .A2(_0776_),
    .Y(_0089_),
    .B1(_0777_));
 sg13g2_nor2_1 _1684_ (.A(_0134_),
    .B(_0517_),
    .Y(_0778_));
 sg13g2_a21o_1 _1685_ (.A2(_0775_),
    .A1(_0774_),
    .B1(_0778_),
    .X(_0779_));
 sg13g2_nor2_1 _1686_ (.A(_0007_),
    .B(_0732_),
    .Y(_0780_));
 sg13g2_xor2_1 _1687_ (.B(net223),
    .A(_0007_),
    .X(_0781_));
 sg13g2_nand2_1 _1688_ (.Y(_0782_),
    .A(_0779_),
    .B(_0781_));
 sg13g2_xnor2_1 _1689_ (.Y(_0783_),
    .A(_0779_),
    .B(_0781_));
 sg13g2_o21ai_1 _1690_ (.B1(net267),
    .Y(_0784_),
    .A1(net281),
    .A2(net210));
 sg13g2_a21oi_1 _1691_ (.A1(net209),
    .A2(_0783_),
    .Y(_0090_),
    .B1(_0784_));
 sg13g2_o21ai_1 _1692_ (.B1(net267),
    .Y(_0785_),
    .A1(\square_y[9] ),
    .A2(net211));
 sg13g2_nor2_1 _1693_ (.A(\square_y[8] ),
    .B(net224),
    .Y(_0786_));
 sg13g2_a22oi_1 _1694_ (.Y(_0787_),
    .B1(_0782_),
    .B2(_0786_),
    .A2(_0780_),
    .A1(_0779_));
 sg13g2_xnor2_1 _1695_ (.Y(_0788_),
    .A(net181),
    .B(_0787_));
 sg13g2_a21oi_1 _1696_ (.A1(net211),
    .A2(_0788_),
    .Y(_0091_),
    .B1(_0785_));
 sg13g2_and2_1 _1697_ (.A(net271),
    .B(net1),
    .X(_0092_));
 sg13g2_and2_1 _1698_ (.A(net270),
    .B(net118),
    .X(_0093_));
 sg13g2_nand4_1 _1699_ (.B(_0153_),
    .C(net249),
    .A(_0152_),
    .Y(_0789_),
    .D(net250));
 sg13g2_nand4_1 _1700_ (.B(_0151_),
    .C(_0210_),
    .A(\pix_y[9] ),
    .Y(_0790_),
    .D(_0254_));
 sg13g2_o21ai_1 _1701_ (.B1(net271),
    .Y(_0791_),
    .A1(_0789_),
    .A2(_0790_));
 sg13g2_or2_2 _1702_ (.X(_0792_),
    .B(_0791_),
    .A(_0558_));
 sg13g2_inv_1 _1703_ (.Y(_0793_),
    .A(_0792_));
 sg13g2_a22oi_1 _1704_ (.Y(_0794_),
    .B1(_0793_),
    .B2(net114),
    .A2(net215),
    .A1(\pix_y[0] ));
 sg13g2_inv_1 _1705_ (.Y(_0094_),
    .A(net115));
 sg13g2_nand2_1 _1706_ (.Y(_0795_),
    .A(net255),
    .B(net319));
 sg13g2_nand3_1 _1707_ (.B(_0793_),
    .C(_0795_),
    .A(_0211_),
    .Y(_0796_));
 sg13g2_o21ai_1 _1708_ (.B1(_0796_),
    .Y(_0095_),
    .A1(net240),
    .A2(net214));
 sg13g2_nand3_1 _1709_ (.B(\pix_y[0] ),
    .C(net214),
    .A(net255),
    .Y(_0797_));
 sg13g2_and2_2 _1710_ (.A(net214),
    .B(_0791_),
    .X(_0798_));
 sg13g2_xnor2_1 _1711_ (.Y(_0799_),
    .A(_0157_),
    .B(_0797_));
 sg13g2_nor2_1 _1712_ (.A(_0798_),
    .B(net306),
    .Y(_0096_));
 sg13g2_nand2_1 _1713_ (.Y(_0800_),
    .A(net248),
    .B(net215));
 sg13g2_nand3b_1 _1714_ (.B(net320),
    .C(net255),
    .Y(_0801_),
    .A_N(net316));
 sg13g2_xnor2_1 _1715_ (.Y(_0802_),
    .A(_0156_),
    .B(_0801_));
 sg13g2_o21ai_1 _1716_ (.B1(_0800_),
    .Y(_0097_),
    .A1(_0792_),
    .A2(_0802_));
 sg13g2_nand4_1 _1717_ (.B(net250),
    .C(net255),
    .A(net248),
    .Y(_0803_),
    .D(\pix_y[0] ));
 sg13g2_nor2_1 _1718_ (.A(net215),
    .B(_0803_),
    .Y(_0804_));
 sg13g2_xnor2_1 _1719_ (.Y(_0805_),
    .A(net247),
    .B(_0804_));
 sg13g2_nor2_1 _1720_ (.A(_0798_),
    .B(_0805_),
    .Y(_0098_));
 sg13g2_nand2_1 _1721_ (.Y(_0806_),
    .A(net244),
    .B(net215));
 sg13g2_nor2_1 _1722_ (.A(net202),
    .B(_0803_),
    .Y(_0807_));
 sg13g2_xnor2_1 _1723_ (.Y(_0808_),
    .A(net244),
    .B(_0807_));
 sg13g2_o21ai_1 _1724_ (.B1(_0806_),
    .Y(_0099_),
    .A1(_0792_),
    .A2(net203));
 sg13g2_nor3_2 _1725_ (.A(_0200_),
    .B(net215),
    .C(_0803_),
    .Y(_0809_));
 sg13g2_xnor2_1 _1726_ (.Y(_0810_),
    .A(net299),
    .B(_0809_));
 sg13g2_nor2_1 _1727_ (.A(_0798_),
    .B(_0810_),
    .Y(_0100_));
 sg13g2_nor3_1 _1728_ (.A(_0153_),
    .B(_0798_),
    .C(_0809_),
    .Y(_0811_));
 sg13g2_nor4_1 _1729_ (.A(_0200_),
    .B(_0299_),
    .C(_0792_),
    .D(_0803_),
    .Y(_0812_));
 sg13g2_or2_1 _1730_ (.X(_0101_),
    .B(_0812_),
    .A(_0811_));
 sg13g2_nor3_1 _1731_ (.A(_0298_),
    .B(net215),
    .C(_0803_),
    .Y(_0813_));
 sg13g2_a21oi_1 _1732_ (.A1(_0184_),
    .A2(_0809_),
    .Y(_0814_),
    .B1(net242));
 sg13g2_nor3_1 _1733_ (.A(_0798_),
    .B(_0813_),
    .C(_0814_),
    .Y(_0102_));
 sg13g2_nand2_1 _1734_ (.Y(_0815_),
    .A(net241),
    .B(net215));
 sg13g2_nor4_1 _1735_ (.A(net289),
    .B(_0185_),
    .C(_0200_),
    .D(_0803_),
    .Y(_0816_));
 sg13g2_xnor2_1 _1736_ (.Y(_0817_),
    .A(net241),
    .B(_0816_));
 sg13g2_o21ai_1 _1737_ (.B1(_0815_),
    .Y(_0103_),
    .A1(_0792_),
    .A2(_0817_));
 sg13g2_nor2b_1 _1738_ (.A(\driver.driver.pmod_clk_prev ),
    .B_N(\driver.driver.pmod_clk_sync[1] ),
    .Y(_0818_));
 sg13g2_nor2_1 _1739_ (.A(net265),
    .B(net232),
    .Y(_0819_));
 sg13g2_a22oi_1 _1740_ (.Y(_0104_),
    .B1(net228),
    .B2(_0130_),
    .A2(net233),
    .A1(_0131_));
 sg13g2_a22oi_1 _1741_ (.Y(_0105_),
    .B1(net228),
    .B2(_0129_),
    .A2(net233),
    .A1(_0130_));
 sg13g2_a22oi_1 _1742_ (.Y(_0106_),
    .B1(net227),
    .B2(_0128_),
    .A2(net233),
    .A1(_0129_));
 sg13g2_a22oi_1 _1743_ (.Y(_0107_),
    .B1(net227),
    .B2(_0127_),
    .A2(net232),
    .A1(_0128_));
 sg13g2_a22oi_1 _1744_ (.Y(_0108_),
    .B1(net227),
    .B2(_0126_),
    .A2(net232),
    .A1(_0127_));
 sg13g2_a22oi_1 _1745_ (.Y(_0109_),
    .B1(net227),
    .B2(_0125_),
    .A2(net232),
    .A1(_0126_));
 sg13g2_a22oi_1 _1746_ (.Y(_0110_),
    .B1(net227),
    .B2(_0124_),
    .A2(net232),
    .A1(_0125_));
 sg13g2_a22oi_1 _1747_ (.Y(_0111_),
    .B1(net227),
    .B2(_0123_),
    .A2(net232),
    .A1(_0124_));
 sg13g2_a22oi_1 _1748_ (.Y(_0112_),
    .B1(net227),
    .B2(_0122_),
    .A2(net232),
    .A1(_0123_));
 sg13g2_a22oi_1 _1749_ (.Y(_0113_),
    .B1(net227),
    .B2(_0121_),
    .A2(net232),
    .A1(_0122_));
 sg13g2_a22oi_1 _1750_ (.Y(_0114_),
    .B1(net228),
    .B2(_0120_),
    .A2(net233),
    .A1(_0121_));
 sg13g2_a22oi_1 _1751_ (.Y(_0115_),
    .B1(net228),
    .B2(_0145_),
    .A2(net233),
    .A1(_0120_));
 sg13g2_and2_1 _1752_ (.A(net270),
    .B(net3),
    .X(_0116_));
 sg13g2_and2_1 _1753_ (.A(net270),
    .B(net116),
    .X(_0117_));
 sg13g2_and2_1 _1754_ (.A(net270),
    .B(net2),
    .X(_0118_));
 sg13g2_and2_1 _1755_ (.A(net270),
    .B(net117),
    .X(_0119_));
 sg13g2_dfrbp_1 _1756_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net80),
    .D(_0034_),
    .Q_N(_0874_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _1757_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net102),
    .D(net140),
    .Q_N(_0873_),
    .Q(\driver.decoder.data_reg[0] ));
 sg13g2_dfrbp_1 _1758_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net100),
    .D(net148),
    .Q_N(_0872_),
    .Q(\driver.decoder.data_reg[1] ));
 sg13g2_dfrbp_1 _1759_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net98),
    .D(net156),
    .Q_N(_0871_),
    .Q(\driver.decoder.data_reg[2] ));
 sg13g2_dfrbp_1 _1760_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net96),
    .D(net136),
    .Q_N(_0870_),
    .Q(\driver.decoder.data_reg[3] ));
 sg13g2_dfrbp_1 _1761_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net94),
    .D(_0039_),
    .Q_N(_0869_),
    .Q(\driver.decoder.data_reg[4] ));
 sg13g2_dfrbp_1 _1762_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net89),
    .D(_0040_),
    .Q_N(_0868_),
    .Q(\driver.decoder.data_reg[5] ));
 sg13g2_dfrbp_1 _1763_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net87),
    .D(_0041_),
    .Q_N(_0867_),
    .Q(\driver.decoder.data_reg[6] ));
 sg13g2_dfrbp_1 _1764_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net85),
    .D(_0042_),
    .Q_N(_0866_),
    .Q(\driver.decoder.data_reg[7] ));
 sg13g2_dfrbp_1 _1765_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net83),
    .D(net150),
    .Q_N(_0865_),
    .Q(\driver.decoder.data_reg[8] ));
 sg13g2_dfrbp_1 _1766_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net81),
    .D(net144),
    .Q_N(_0864_),
    .Q(\driver.decoder.data_reg[9] ));
 sg13g2_dfrbp_1 _1767_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net78),
    .D(net146),
    .Q_N(_0863_),
    .Q(\driver.decoder.data_reg[10] ));
 sg13g2_dfrbp_1 _1768_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net76),
    .D(net138),
    .Q_N(_0862_),
    .Q(\driver.decoder.data_reg[11] ));
 sg13g2_dfrbp_1 _1769_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net74),
    .D(_0047_),
    .Q_N(_0033_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 _1770_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net73),
    .D(net185),
    .Q_N(_0861_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 _1771_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net72),
    .D(_0049_),
    .Q_N(_0860_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 _1772_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net71),
    .D(_0050_),
    .Q_N(_0859_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 _1773_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net70),
    .D(_0051_),
    .Q_N(_0858_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 _1774_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net69),
    .D(_0052_),
    .Q_N(_0857_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 _1775_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net68),
    .D(net128),
    .Q_N(_0856_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 _1776_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net67),
    .D(_0054_),
    .Q_N(_0855_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 _1777_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net66),
    .D(_0055_),
    .Q_N(_0854_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 _1778_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net65),
    .D(_0056_),
    .Q_N(_0853_),
    .Q(\counter[9] ));
 sg13g2_dfrbp_1 _1779_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net64),
    .D(net134),
    .Q_N(_0852_),
    .Q(\counter[10] ));
 sg13g2_dfrbp_1 _1780_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net63),
    .D(_0058_),
    .Q_N(_0851_),
    .Q(\counter[11] ));
 sg13g2_dfrbp_1 _1781_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net62),
    .D(net125),
    .Q_N(_0850_),
    .Q(\counter[12] ));
 sg13g2_dfrbp_1 _1782_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net61),
    .D(_0060_),
    .Q_N(_0849_),
    .Q(\counter[13] ));
 sg13g2_dfrbp_1 _1783_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net60),
    .D(_0061_),
    .Q_N(_0032_),
    .Q(\pix_x[0] ));
 sg13g2_dfrbp_1 _1784_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net59),
    .D(_0062_),
    .Q_N(_0848_),
    .Q(\pix_x[1] ));
 sg13g2_dfrbp_1 _1785_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net58),
    .D(_0063_),
    .Q_N(_0018_),
    .Q(\pix_x[2] ));
 sg13g2_dfrbp_1 _1786_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net57),
    .D(_0064_),
    .Q_N(_0017_),
    .Q(\pix_x[3] ));
 sg13g2_dfrbp_1 _1787_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net56),
    .D(_0065_),
    .Q_N(_0002_),
    .Q(\pix_x[4] ));
 sg13g2_dfrbp_1 _1788_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net55),
    .D(_0066_),
    .Q_N(_0021_),
    .Q(\pix_x[5] ));
 sg13g2_dfrbp_1 _1789_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net54),
    .D(net315),
    .Q_N(_0847_),
    .Q(\pix_x[6] ));
 sg13g2_dfrbp_1 _1790_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net53),
    .D(net304),
    .Q_N(_0846_),
    .Q(\pix_x[7] ));
 sg13g2_dfrbp_1 _1791_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net52),
    .D(_0069_),
    .Q_N(_0845_),
    .Q(\pix_x[8] ));
 sg13g2_dfrbp_1 _1792_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net51),
    .D(_0070_),
    .Q_N(_0844_),
    .Q(\pix_x[9] ));
 sg13g2_dfrbp_1 _1793_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net50),
    .D(_0071_),
    .Q_N(_0843_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _1794_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net49),
    .D(net122),
    .Q_N(_0031_),
    .Q(\square_x[0] ));
 sg13g2_dfrbp_1 _1795_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net47),
    .D(net273),
    .Q_N(_0013_),
    .Q(\square_x[1] ));
 sg13g2_dfrbp_1 _1796_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net45),
    .D(_0074_),
    .Q_N(_0842_),
    .Q(\square_x[2] ));
 sg13g2_dfrbp_1 _1797_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net43),
    .D(_0075_),
    .Q_N(_0014_),
    .Q(\square_x[3] ));
 sg13g2_dfrbp_1 _1798_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net41),
    .D(_0076_),
    .Q_N(_0841_),
    .Q(\square_x[4] ));
 sg13g2_dfrbp_1 _1799_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net39),
    .D(_0077_),
    .Q_N(_0015_),
    .Q(\square_x[5] ));
 sg13g2_dfrbp_1 _1800_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net37),
    .D(_0078_),
    .Q_N(_0005_),
    .Q(\square_x[6] ));
 sg13g2_dfrbp_1 _1801_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net35),
    .D(_0079_),
    .Q_N(_0016_),
    .Q(\square_x[7] ));
 sg13g2_dfrbp_1 _1802_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net33),
    .D(_0080_),
    .Q_N(_0004_),
    .Q(\square_x[8] ));
 sg13g2_dfrbp_1 _1803_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net31),
    .D(net199),
    .Q_N(_0003_),
    .Q(\square_x[9] ));
 sg13g2_dfrbp_1 _1804_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net29),
    .D(net120),
    .Q_N(_0030_),
    .Q(\square_y[0] ));
 sg13g2_dfrbp_1 _1805_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net27),
    .D(net152),
    .Q_N(_0010_),
    .Q(\square_y[1] ));
 sg13g2_dfrbp_1 _1806_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net25),
    .D(net287),
    .Q_N(_0840_),
    .Q(\square_y[2] ));
 sg13g2_dfrbp_1 _1807_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net23),
    .D(net191),
    .Q_N(_0011_),
    .Q(\square_y[3] ));
 sg13g2_dfrbp_1 _1808_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net21),
    .D(net298),
    .Q_N(_0839_),
    .Q(\square_y[4] ));
 sg13g2_dfrbp_1 _1809_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net109),
    .D(net296),
    .Q_N(_0012_),
    .Q(\square_y[5] ));
 sg13g2_dfrbp_1 _1810_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net107),
    .D(net278),
    .Q_N(_0009_),
    .Q(\square_y[6] ));
 sg13g2_dfrbp_1 _1811_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net105),
    .D(net280),
    .Q_N(_0008_),
    .Q(\square_y[7] ));
 sg13g2_dfrbp_1 _1812_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net103),
    .D(net282),
    .Q_N(_0007_),
    .Q(\square_y[8] ));
 sg13g2_dfrbp_1 _1813_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net99),
    .D(net182),
    .Q_N(_0006_),
    .Q(\square_y[9] ));
 sg13g2_dfrbp_1 _1814_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net95),
    .D(_0092_),
    .Q_N(_0838_),
    .Q(\driver.driver.pmod_latch_sync[0] ));
 sg13g2_dfrbp_1 _1815_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net91),
    .D(_0093_),
    .Q_N(_0875_),
    .Q(\driver.driver.pmod_latch_sync[1] ));
 sg13g2_dfrbp_1 _1816_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net90),
    .D(net312),
    .Q_N(_0837_),
    .Q(hsync));
 sg13g2_dfrbp_1 _1817_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net88),
    .D(_0094_),
    .Q_N(_0029_),
    .Q(\pix_y[0] ));
 sg13g2_dfrbp_1 _1818_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net84),
    .D(_0095_),
    .Q_N(_0019_),
    .Q(\pix_y[1] ));
 sg13g2_dfrbp_1 _1819_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net79),
    .D(_0096_),
    .Q_N(_0027_),
    .Q(\pix_y[2] ));
 sg13g2_dfrbp_1 _1820_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net75),
    .D(_0097_),
    .Q_N(_0022_),
    .Q(\pix_y[3] ));
 sg13g2_dfrbp_1 _1821_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net46),
    .D(_0098_),
    .Q_N(_0028_),
    .Q(\pix_y[4] ));
 sg13g2_dfrbp_1 _1822_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net42),
    .D(net204),
    .Q_N(_0020_),
    .Q(\pix_y[5] ));
 sg13g2_dfrbp_1 _1823_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net38),
    .D(_0100_),
    .Q_N(_0023_),
    .Q(\pix_y[6] ));
 sg13g2_dfrbp_1 _1824_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net34),
    .D(_0101_),
    .Q_N(_0026_),
    .Q(\pix_y[7] ));
 sg13g2_dfrbp_1 _1825_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net30),
    .D(_0102_),
    .Q_N(_0024_),
    .Q(\pix_y[8] ));
 sg13g2_dfrbp_1 _1826_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net92),
    .D(net290),
    .Q_N(_0025_),
    .Q(\pix_y[9] ));
 sg13g2_dfrbp_1 _1827_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net93),
    .D(net294),
    .Q_N(_0876_),
    .Q(\vga_sync_gen.vsync ));
 sg13g2_dfrbp_1 _1828_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net36),
    .D(net111),
    .Q_N(_0877_),
    .Q(\driver.driver.pmod_clk_prev ));
 sg13g2_dfrbp_1 _1829_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net26),
    .D(net110),
    .Q_N(_0836_),
    .Q(\driver.driver.pmod_latch_prev ));
 sg13g2_dfrbp_1 _1830_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net22),
    .D(net131),
    .Q_N(_0835_),
    .Q(\driver.driver.shift_reg[0] ));
 sg13g2_dfrbp_1 _1831_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net108),
    .D(net158),
    .Q_N(_0834_),
    .Q(\driver.driver.shift_reg[1] ));
 sg13g2_dfrbp_1 _1832_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net104),
    .D(_0106_),
    .Q_N(_0833_),
    .Q(\driver.driver.shift_reg[2] ));
 sg13g2_dfrbp_1 _1833_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net97),
    .D(net154),
    .Q_N(_0832_),
    .Q(\driver.driver.shift_reg[3] ));
 sg13g2_dfrbp_1 _1834_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net82),
    .D(_0108_),
    .Q_N(_0831_),
    .Q(\driver.driver.shift_reg[4] ));
 sg13g2_dfrbp_1 _1835_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net48),
    .D(net160),
    .Q_N(_0830_),
    .Q(\driver.driver.shift_reg[5] ));
 sg13g2_dfrbp_1 _1836_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net40),
    .D(_0110_),
    .Q_N(_0829_),
    .Q(\driver.driver.shift_reg[6] ));
 sg13g2_dfrbp_1 _1837_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net32),
    .D(net172),
    .Q_N(_0828_),
    .Q(\driver.driver.shift_reg[7] ));
 sg13g2_dfrbp_1 _1838_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net24),
    .D(net169),
    .Q_N(_0827_),
    .Q(\driver.driver.shift_reg[8] ));
 sg13g2_dfrbp_1 _1839_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net106),
    .D(_0113_),
    .Q_N(_0826_),
    .Q(\driver.driver.shift_reg[9] ));
 sg13g2_dfrbp_1 _1840_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net86),
    .D(net164),
    .Q_N(_0825_),
    .Q(\driver.driver.shift_reg[10] ));
 sg13g2_dfrbp_1 _1841_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net44),
    .D(net142),
    .Q_N(_0824_),
    .Q(\driver.driver.shift_reg[11] ));
 sg13g2_dfrbp_1 _1842_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net28),
    .D(_0116_),
    .Q_N(_0823_),
    .Q(\driver.driver.pmod_data_sync[0] ));
 sg13g2_dfrbp_1 _1843_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net20),
    .D(_0117_),
    .Q_N(_0822_),
    .Q(\driver.driver.pmod_data_sync[1] ));
 sg13g2_dfrbp_1 _1844_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net101),
    .D(_0118_),
    .Q_N(_0821_),
    .Q(\driver.driver.pmod_clk_sync[0] ));
 sg13g2_dfrbp_1 _1845_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net77),
    .D(_0119_),
    .Q_N(_0820_),
    .Q(\driver.driver.pmod_clk_sync[1] ));
 sg13g2_tiehi _1808__21 (.L_HI(net21));
 sg13g2_tiehi _1830__22 (.L_HI(net22));
 sg13g2_tiehi _1807__23 (.L_HI(net23));
 sg13g2_tiehi _1838__24 (.L_HI(net24));
 sg13g2_tiehi _1806__25 (.L_HI(net25));
 sg13g2_tiehi _1829__26 (.L_HI(net26));
 sg13g2_tiehi _1805__27 (.L_HI(net27));
 sg13g2_tiehi _1842__28 (.L_HI(net28));
 sg13g2_tiehi _1804__29 (.L_HI(net29));
 sg13g2_tiehi _1825__30 (.L_HI(net30));
 sg13g2_tiehi _1803__31 (.L_HI(net31));
 sg13g2_tiehi _1837__32 (.L_HI(net32));
 sg13g2_tiehi _1802__33 (.L_HI(net33));
 sg13g2_tiehi _1824__34 (.L_HI(net34));
 sg13g2_tiehi _1801__35 (.L_HI(net35));
 sg13g2_tiehi _1828__36 (.L_HI(net36));
 sg13g2_tiehi _1800__37 (.L_HI(net37));
 sg13g2_tiehi _1823__38 (.L_HI(net38));
 sg13g2_tiehi _1799__39 (.L_HI(net39));
 sg13g2_tiehi _1836__40 (.L_HI(net40));
 sg13g2_tiehi _1798__41 (.L_HI(net41));
 sg13g2_tiehi _1822__42 (.L_HI(net42));
 sg13g2_tiehi _1797__43 (.L_HI(net43));
 sg13g2_tiehi _1841__44 (.L_HI(net44));
 sg13g2_tiehi _1796__45 (.L_HI(net45));
 sg13g2_tiehi _1821__46 (.L_HI(net46));
 sg13g2_tiehi _1795__47 (.L_HI(net47));
 sg13g2_tiehi _1835__48 (.L_HI(net48));
 sg13g2_tiehi _1794__49 (.L_HI(net49));
 sg13g2_tiehi _1793__50 (.L_HI(net50));
 sg13g2_tiehi _1792__51 (.L_HI(net51));
 sg13g2_tiehi _1791__52 (.L_HI(net52));
 sg13g2_tiehi _1790__53 (.L_HI(net53));
 sg13g2_tiehi _1789__54 (.L_HI(net54));
 sg13g2_tiehi _1788__55 (.L_HI(net55));
 sg13g2_tiehi _1787__56 (.L_HI(net56));
 sg13g2_tiehi _1786__57 (.L_HI(net57));
 sg13g2_tiehi _1785__58 (.L_HI(net58));
 sg13g2_tiehi _1784__59 (.L_HI(net59));
 sg13g2_tiehi _1783__60 (.L_HI(net60));
 sg13g2_tiehi _1782__61 (.L_HI(net61));
 sg13g2_tiehi _1781__62 (.L_HI(net62));
 sg13g2_tiehi _1780__63 (.L_HI(net63));
 sg13g2_tiehi _1779__64 (.L_HI(net64));
 sg13g2_tiehi _1778__65 (.L_HI(net65));
 sg13g2_tiehi _1777__66 (.L_HI(net66));
 sg13g2_tiehi _1776__67 (.L_HI(net67));
 sg13g2_tiehi _1775__68 (.L_HI(net68));
 sg13g2_tiehi _1774__69 (.L_HI(net69));
 sg13g2_tiehi _1773__70 (.L_HI(net70));
 sg13g2_tiehi _1772__71 (.L_HI(net71));
 sg13g2_tiehi _1771__72 (.L_HI(net72));
 sg13g2_tiehi _1770__73 (.L_HI(net73));
 sg13g2_tiehi _1769__74 (.L_HI(net74));
 sg13g2_tiehi _1820__75 (.L_HI(net75));
 sg13g2_tiehi _1768__76 (.L_HI(net76));
 sg13g2_tiehi _1845__77 (.L_HI(net77));
 sg13g2_tiehi _1767__78 (.L_HI(net78));
 sg13g2_tiehi _1819__79 (.L_HI(net79));
 sg13g2_tiehi _1756__80 (.L_HI(net80));
 sg13g2_tiehi _1766__81 (.L_HI(net81));
 sg13g2_tiehi _1834__82 (.L_HI(net82));
 sg13g2_tiehi _1765__83 (.L_HI(net83));
 sg13g2_tiehi _1818__84 (.L_HI(net84));
 sg13g2_tiehi _1764__85 (.L_HI(net85));
 sg13g2_tiehi _1840__86 (.L_HI(net86));
 sg13g2_tiehi _1763__87 (.L_HI(net87));
 sg13g2_tiehi _1817__88 (.L_HI(net88));
 sg13g2_tiehi _1762__89 (.L_HI(net89));
 sg13g2_tiehi _1816__90 (.L_HI(net90));
 sg13g2_tiehi _1815__91 (.L_HI(net91));
 sg13g2_tiehi _1826__92 (.L_HI(net92));
 sg13g2_tiehi _1827__93 (.L_HI(net93));
 sg13g2_tiehi _1761__94 (.L_HI(net94));
 sg13g2_tiehi _1814__95 (.L_HI(net95));
 sg13g2_tiehi _1760__96 (.L_HI(net96));
 sg13g2_tiehi _1833__97 (.L_HI(net97));
 sg13g2_tiehi _1759__98 (.L_HI(net98));
 sg13g2_tiehi _1813__99 (.L_HI(net99));
 sg13g2_tiehi _1758__100 (.L_HI(net100));
 sg13g2_tiehi _1844__101 (.L_HI(net101));
 sg13g2_tiehi _1757__102 (.L_HI(net102));
 sg13g2_tiehi _1812__103 (.L_HI(net103));
 sg13g2_tiehi _1832__104 (.L_HI(net104));
 sg13g2_tiehi _1811__105 (.L_HI(net105));
 sg13g2_tiehi _1839__106 (.L_HI(net106));
 sg13g2_tiehi _1810__107 (.L_HI(net107));
 sg13g2_tiehi _1831__108 (.L_HI(net108));
 sg13g2_tiehi _1809__109 (.L_HI(net109));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_spacewar_5 (.L_LO(net5));
 sg13g2_tielo tt_um_spacewar_6 (.L_LO(net6));
 sg13g2_tielo tt_um_spacewar_7 (.L_LO(net7));
 sg13g2_tielo tt_um_spacewar_8 (.L_LO(net8));
 sg13g2_tielo tt_um_spacewar_9 (.L_LO(net9));
 sg13g2_tielo tt_um_spacewar_10 (.L_LO(net10));
 sg13g2_tielo tt_um_spacewar_11 (.L_LO(net11));
 sg13g2_tielo tt_um_spacewar_12 (.L_LO(net12));
 sg13g2_tielo tt_um_spacewar_13 (.L_LO(net13));
 sg13g2_tielo tt_um_spacewar_14 (.L_LO(net14));
 sg13g2_tielo tt_um_spacewar_15 (.L_LO(net15));
 sg13g2_tielo tt_um_spacewar_16 (.L_LO(net16));
 sg13g2_tielo tt_um_spacewar_17 (.L_LO(net17));
 sg13g2_tielo tt_um_spacewar_18 (.L_LO(net18));
 sg13g2_tielo tt_um_spacewar_19 (.L_LO(net19));
 sg13g2_tiehi _1843__20 (.L_HI(net20));
 sg13g2_buf_1 _1952_ (.A(uo_out[6]),
    .X(uo_out[0]));
 sg13g2_buf_1 _1953_ (.A(uo_out[5]),
    .X(uo_out[1]));
 sg13g2_buf_1 _1954_ (.A(uo_out[6]),
    .X(uo_out[2]));
 sg13g2_buf_1 _1955_ (.A(\vga_sync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _1956_ (.A(uo_out[6]),
    .X(uo_out[4]));
 sg13g2_buf_1 _1957_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout205 (.A(_0333_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(net208),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(net208),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_0290_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(net211),
    .X(net209));
 sg13g2_buf_1 fanout210 (.A(net211),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_0736_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(net213),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_0671_),
    .X(net213));
 sg13g2_buf_4 fanout214 (.X(net214),
    .A(_0560_));
 sg13g2_buf_4 fanout215 (.X(net215),
    .A(_0559_));
 sg13g2_buf_2 fanout216 (.A(_0264_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_0247_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(net219),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_0278_),
    .X(net219));
 sg13g2_buf_4 fanout220 (.X(net220),
    .A(_0268_));
 sg13g2_buf_2 fanout221 (.A(net222),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_0261_),
    .X(net222));
 sg13g2_buf_4 fanout223 (.X(net223),
    .A(_0731_));
 sg13g2_buf_2 fanout224 (.A(_0731_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_0660_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_0660_),
    .X(net226));
 sg13g2_buf_4 fanout227 (.X(net227),
    .A(_0819_));
 sg13g2_buf_2 fanout228 (.A(_0819_),
    .X(net228));
 sg13g2_buf_4 fanout229 (.X(net229),
    .A(_0529_));
 sg13g2_buf_2 fanout230 (.A(_0529_),
    .X(net230));
 sg13g2_buf_4 fanout231 (.X(net231),
    .A(_0198_));
 sg13g2_buf_2 fanout232 (.A(_0818_),
    .X(net232));
 sg13g2_buf_1 fanout233 (.A(_0818_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_0528_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_0528_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_0207_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_0177_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(net240),
    .X(net238));
 sg13g2_buf_1 fanout239 (.A(net240),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_0158_),
    .X(net240));
 sg13g2_buf_4 fanout241 (.X(net241),
    .A(\pix_y[9] ));
 sg13g2_buf_2 fanout242 (.A(net307),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(\pix_y[7] ),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(\pix_y[5] ),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(\pix_y[5] ),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(net247),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(net309),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(net249),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(\pix_y[3] ),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(\pix_y[2] ),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(net254),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(net253),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(net254),
    .X(net253));
 sg13g2_buf_1 fanout254 (.A(\pix_y[1] ),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(\pix_y[1] ),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(\square_x[4] ),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(net311),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(net317),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(net260),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(net302),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(net314),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(\pix_x[5] ),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(net300),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(\pix_x[4] ),
    .X(net264));
 sg13g2_buf_4 fanout265 (.X(net265),
    .A(net266));
 sg13g2_buf_4 fanout266 (.X(net266),
    .A(_0171_));
 sg13g2_buf_2 fanout267 (.A(net268),
    .X(net267));
 sg13g2_buf_4 fanout268 (.X(net268),
    .A(net271));
 sg13g2_buf_2 fanout269 (.A(net270),
    .X(net269));
 sg13g2_buf_4 fanout270 (.X(net270),
    .A(net271));
 sg13g2_buf_2 fanout271 (.A(rst_n),
    .X(net271));
 sg13g2_buf_1 input1 (.A(ui_in[4]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[5]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[6]),
    .X(net3));
 sg13g2_tielo tt_um_spacewar_4 (.L_LO(net4));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\driver.driver.pmod_latch_sync[1] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold2 (.A(\driver.driver.pmod_clk_sync[1] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0032_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0033_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0029_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0794_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold7 (.A(\driver.driver.pmod_data_sync[0] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold8 (.A(\driver.driver.pmod_clk_sync[0] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold9 (.A(\driver.driver.pmod_latch_sync[0] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0030_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0082_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0031_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0072_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold14 (.A(\counter[12] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0551_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0059_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold17 (.A(\counter[6] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0540_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0053_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0002_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold21 (.A(\driver.driver.pmod_data_sync[1] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0104_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold23 (.A(\counter[10] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0548_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0057_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold26 (.A(\driver.decoder.data_reg[3] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0038_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold28 (.A(\driver.decoder.data_reg[11] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0046_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold30 (.A(\driver.decoder.data_reg[0] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0035_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold32 (.A(\driver.driver.shift_reg[11] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0115_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold34 (.A(\driver.decoder.data_reg[9] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0044_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold36 (.A(\driver.decoder.data_reg[10] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0045_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold38 (.A(\driver.decoder.data_reg[1] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0036_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold40 (.A(\driver.decoder.data_reg[8] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0043_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold42 (.A(\square_y[1] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0083_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold44 (.A(\driver.driver.shift_reg[3] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0107_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold46 (.A(\driver.decoder.data_reg[2] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0037_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold48 (.A(\driver.driver.shift_reg[1] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0105_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold50 (.A(\driver.driver.shift_reg[5] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0109_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0018_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0563_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold54 (.A(\driver.driver.shift_reg[10] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0114_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold56 (.A(\driver.driver.shift_reg[4] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold57 (.A(\counter[2] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0532_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold59 (.A(\driver.driver.shift_reg[8] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0112_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold61 (.A(\driver.driver.shift_reg[9] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold62 (.A(\driver.driver.shift_reg[7] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0111_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold64 (.A(\driver.driver.shift_reg[2] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold65 (.A(\driver.driver.shift_reg[6] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold66 (.A(\driver.decoder.data_reg[4] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold67 (.A(\counter[13] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0554_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold69 (.A(\driver.decoder.data_reg[6] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold70 (.A(\counter[11] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0550_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0006_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0091_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold74 (.A(\counter[1] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0531_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0048_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold77 (.A(\counter[5] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0539_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold79 (.A(\counter[9] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0547_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold81 (.A(\square_y[3] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0085_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold83 (.A(\counter[8] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0546_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold85 (.A(\driver.decoder.data_reg[7] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold86 (.A(\driver.decoder.data_reg[5] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold87 (.A(\counter[4] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0538_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold89 (.A(\square_x[9] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0081_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold91 (.A(\square_x[4] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0697_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0028_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0808_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0099_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold96 (.A(\square_x[1] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0073_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold98 (.A(\counter[3] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold99 (.A(\square_x[7] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold100 (.A(\counter[7] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold101 (.A(\square_y[6] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0088_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold103 (.A(\square_y[7] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0089_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold105 (.A(\square_y[8] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0090_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold107 (.A(\pix_x[0] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0238_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold109 (.A(\pix_x[2] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold110 (.A(\square_y[2] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0084_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold112 (.A(\square_x[3] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0024_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0103_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold115 (.A(\square_x[5] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold116 (.A(\pix_y[9] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0188_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0001_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0012_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0087_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold121 (.A(\square_y[4] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0086_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold123 (.A(\pix_y[6] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold124 (.A(\pix_x[4] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0566_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold126 (.A(\pix_x[7] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0569_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0068_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold129 (.A(\pix_y[2] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0799_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold131 (.A(\pix_y[8] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold132 (.A(\square_x[8] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold133 (.A(\pix_y[4] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold134 (.A(\square_x[2] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold135 (.A(\pix_x[9] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0000_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold137 (.A(\square_x[6] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold138 (.A(\pix_x[6] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0067_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0027_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold141 (.A(\pix_x[8] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold142 (.A(\pix_x[6] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold143 (.A(\pix_y[0] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold144 (.A(\pix_y[0] ),
    .X(net320));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_221 ();
 sg13g2_decap_8 FILLER_8_233 ();
 sg13g2_decap_8 FILLER_8_240 ();
 sg13g2_decap_8 FILLER_8_247 ();
 sg13g2_decap_8 FILLER_8_254 ();
 sg13g2_decap_8 FILLER_8_261 ();
 sg13g2_decap_8 FILLER_8_268 ();
 sg13g2_fill_2 FILLER_8_275 ();
 sg13g2_fill_1 FILLER_8_277 ();
 sg13g2_decap_8 FILLER_8_282 ();
 sg13g2_decap_8 FILLER_8_289 ();
 sg13g2_decap_8 FILLER_8_296 ();
 sg13g2_decap_8 FILLER_8_303 ();
 sg13g2_decap_8 FILLER_8_310 ();
 sg13g2_decap_4 FILLER_8_317 ();
 sg13g2_fill_2 FILLER_8_321 ();
 sg13g2_decap_8 FILLER_8_327 ();
 sg13g2_decap_8 FILLER_8_334 ();
 sg13g2_decap_8 FILLER_8_341 ();
 sg13g2_decap_8 FILLER_8_348 ();
 sg13g2_decap_8 FILLER_8_355 ();
 sg13g2_decap_8 FILLER_8_362 ();
 sg13g2_decap_8 FILLER_8_369 ();
 sg13g2_decap_8 FILLER_8_376 ();
 sg13g2_decap_8 FILLER_8_383 ();
 sg13g2_decap_8 FILLER_8_390 ();
 sg13g2_decap_8 FILLER_8_397 ();
 sg13g2_decap_4 FILLER_8_404 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_fill_2 FILLER_9_189 ();
 sg13g2_fill_2 FILLER_9_242 ();
 sg13g2_fill_1 FILLER_9_244 ();
 sg13g2_decap_8 FILLER_9_250 ();
 sg13g2_fill_2 FILLER_9_257 ();
 sg13g2_decap_8 FILLER_9_296 ();
 sg13g2_fill_1 FILLER_9_303 ();
 sg13g2_decap_4 FILLER_9_308 ();
 sg13g2_fill_2 FILLER_9_312 ();
 sg13g2_fill_2 FILLER_9_332 ();
 sg13g2_decap_4 FILLER_9_341 ();
 sg13g2_fill_2 FILLER_9_345 ();
 sg13g2_fill_2 FILLER_9_351 ();
 sg13g2_decap_8 FILLER_9_370 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_384 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_fill_2 FILLER_10_175 ();
 sg13g2_fill_1 FILLER_10_177 ();
 sg13g2_fill_2 FILLER_10_191 ();
 sg13g2_fill_1 FILLER_10_193 ();
 sg13g2_fill_2 FILLER_10_207 ();
 sg13g2_fill_2 FILLER_10_231 ();
 sg13g2_fill_2 FILLER_10_268 ();
 sg13g2_fill_1 FILLER_10_292 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_fill_2 FILLER_11_198 ();
 sg13g2_fill_2 FILLER_11_237 ();
 sg13g2_fill_1 FILLER_11_277 ();
 sg13g2_fill_2 FILLER_11_359 ();
 sg13g2_fill_1 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_397 ();
 sg13g2_decap_4 FILLER_11_404 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_4 FILLER_12_189 ();
 sg13g2_fill_2 FILLER_12_193 ();
 sg13g2_fill_2 FILLER_12_235 ();
 sg13g2_fill_1 FILLER_12_237 ();
 sg13g2_decap_4 FILLER_12_251 ();
 sg13g2_fill_1 FILLER_12_320 ();
 sg13g2_fill_2 FILLER_12_329 ();
 sg13g2_fill_1 FILLER_12_331 ();
 sg13g2_fill_1 FILLER_12_351 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_4 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_4 FILLER_13_77 ();
 sg13g2_fill_2 FILLER_13_81 ();
 sg13g2_decap_8 FILLER_13_86 ();
 sg13g2_decap_8 FILLER_13_93 ();
 sg13g2_decap_4 FILLER_13_100 ();
 sg13g2_fill_2 FILLER_13_104 ();
 sg13g2_fill_2 FILLER_13_110 ();
 sg13g2_fill_1 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_121 ();
 sg13g2_decap_8 FILLER_13_128 ();
 sg13g2_decap_8 FILLER_13_143 ();
 sg13g2_decap_8 FILLER_13_150 ();
 sg13g2_decap_8 FILLER_13_157 ();
 sg13g2_decap_8 FILLER_13_164 ();
 sg13g2_decap_8 FILLER_13_171 ();
 sg13g2_fill_1 FILLER_13_178 ();
 sg13g2_decap_4 FILLER_13_205 ();
 sg13g2_fill_1 FILLER_13_265 ();
 sg13g2_fill_2 FILLER_13_275 ();
 sg13g2_fill_1 FILLER_13_277 ();
 sg13g2_decap_4 FILLER_13_292 ();
 sg13g2_fill_2 FILLER_13_315 ();
 sg13g2_fill_2 FILLER_13_362 ();
 sg13g2_decap_8 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_397 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_fill_2 FILLER_14_49 ();
 sg13g2_fill_2 FILLER_14_55 ();
 sg13g2_decap_8 FILLER_14_62 ();
 sg13g2_fill_1 FILLER_14_69 ();
 sg13g2_fill_2 FILLER_14_78 ();
 sg13g2_fill_1 FILLER_14_94 ();
 sg13g2_fill_1 FILLER_14_121 ();
 sg13g2_decap_8 FILLER_14_152 ();
 sg13g2_decap_4 FILLER_14_159 ();
 sg13g2_decap_8 FILLER_14_167 ();
 sg13g2_decap_4 FILLER_14_174 ();
 sg13g2_fill_1 FILLER_14_178 ();
 sg13g2_fill_1 FILLER_14_196 ();
 sg13g2_fill_2 FILLER_14_220 ();
 sg13g2_decap_4 FILLER_14_249 ();
 sg13g2_fill_1 FILLER_14_253 ();
 sg13g2_fill_2 FILLER_14_332 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_fill_2 FILLER_15_42 ();
 sg13g2_fill_1 FILLER_15_44 ();
 sg13g2_fill_1 FILLER_15_50 ();
 sg13g2_fill_1 FILLER_15_61 ();
 sg13g2_fill_2 FILLER_15_116 ();
 sg13g2_fill_1 FILLER_15_118 ();
 sg13g2_fill_2 FILLER_15_124 ();
 sg13g2_fill_1 FILLER_15_126 ();
 sg13g2_fill_2 FILLER_15_150 ();
 sg13g2_fill_2 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_215 ();
 sg13g2_decap_4 FILLER_15_222 ();
 sg13g2_decap_4 FILLER_15_238 ();
 sg13g2_fill_2 FILLER_15_300 ();
 sg13g2_fill_1 FILLER_15_310 ();
 sg13g2_fill_2 FILLER_15_316 ();
 sg13g2_fill_2 FILLER_15_356 ();
 sg13g2_fill_1 FILLER_15_358 ();
 sg13g2_decap_8 FILLER_15_372 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_4 FILLER_16_28 ();
 sg13g2_fill_1 FILLER_16_98 ();
 sg13g2_fill_1 FILLER_16_113 ();
 sg13g2_fill_2 FILLER_16_119 ();
 sg13g2_fill_2 FILLER_16_126 ();
 sg13g2_fill_2 FILLER_16_145 ();
 sg13g2_fill_1 FILLER_16_208 ();
 sg13g2_decap_4 FILLER_16_235 ();
 sg13g2_decap_8 FILLER_16_244 ();
 sg13g2_fill_2 FILLER_16_251 ();
 sg13g2_fill_1 FILLER_16_262 ();
 sg13g2_fill_2 FILLER_16_285 ();
 sg13g2_fill_1 FILLER_16_287 ();
 sg13g2_fill_1 FILLER_16_298 ();
 sg13g2_fill_1 FILLER_16_329 ();
 sg13g2_decap_4 FILLER_16_363 ();
 sg13g2_fill_1 FILLER_16_367 ();
 sg13g2_decap_8 FILLER_16_372 ();
 sg13g2_decap_8 FILLER_16_379 ();
 sg13g2_decap_8 FILLER_16_386 ();
 sg13g2_decap_8 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_4 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_25 ();
 sg13g2_fill_2 FILLER_17_39 ();
 sg13g2_fill_1 FILLER_17_55 ();
 sg13g2_fill_1 FILLER_17_70 ();
 sg13g2_fill_1 FILLER_17_131 ();
 sg13g2_fill_1 FILLER_17_189 ();
 sg13g2_fill_2 FILLER_17_200 ();
 sg13g2_fill_1 FILLER_17_202 ();
 sg13g2_decap_8 FILLER_17_235 ();
 sg13g2_decap_4 FILLER_17_242 ();
 sg13g2_fill_2 FILLER_17_271 ();
 sg13g2_fill_1 FILLER_17_273 ();
 sg13g2_decap_4 FILLER_17_288 ();
 sg13g2_fill_1 FILLER_17_300 ();
 sg13g2_fill_1 FILLER_17_324 ();
 sg13g2_fill_2 FILLER_17_351 ();
 sg13g2_fill_1 FILLER_17_353 ();
 sg13g2_fill_2 FILLER_17_380 ();
 sg13g2_fill_1 FILLER_17_382 ();
 sg13g2_decap_4 FILLER_17_389 ();
 sg13g2_fill_1 FILLER_17_393 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_fill_2 FILLER_18_14 ();
 sg13g2_fill_1 FILLER_18_16 ();
 sg13g2_fill_1 FILLER_18_43 ();
 sg13g2_fill_1 FILLER_18_66 ();
 sg13g2_fill_1 FILLER_18_84 ();
 sg13g2_fill_2 FILLER_18_119 ();
 sg13g2_fill_2 FILLER_18_128 ();
 sg13g2_decap_8 FILLER_18_145 ();
 sg13g2_decap_4 FILLER_18_152 ();
 sg13g2_fill_2 FILLER_18_156 ();
 sg13g2_decap_8 FILLER_18_162 ();
 sg13g2_decap_4 FILLER_18_169 ();
 sg13g2_fill_1 FILLER_18_173 ();
 sg13g2_fill_2 FILLER_18_194 ();
 sg13g2_fill_1 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_236 ();
 sg13g2_fill_1 FILLER_18_262 ();
 sg13g2_fill_1 FILLER_18_306 ();
 sg13g2_fill_1 FILLER_18_318 ();
 sg13g2_fill_2 FILLER_18_323 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_4 FILLER_19_21 ();
 sg13g2_fill_1 FILLER_19_25 ();
 sg13g2_fill_2 FILLER_19_52 ();
 sg13g2_fill_1 FILLER_19_54 ();
 sg13g2_fill_2 FILLER_19_86 ();
 sg13g2_fill_1 FILLER_19_88 ();
 sg13g2_decap_4 FILLER_19_123 ();
 sg13g2_decap_4 FILLER_19_137 ();
 sg13g2_fill_1 FILLER_19_141 ();
 sg13g2_fill_2 FILLER_19_168 ();
 sg13g2_fill_1 FILLER_19_170 ();
 sg13g2_fill_1 FILLER_19_175 ();
 sg13g2_fill_1 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_207 ();
 sg13g2_decap_4 FILLER_19_214 ();
 sg13g2_fill_1 FILLER_19_241 ();
 sg13g2_fill_2 FILLER_19_265 ();
 sg13g2_decap_8 FILLER_19_272 ();
 sg13g2_decap_8 FILLER_19_279 ();
 sg13g2_fill_2 FILLER_19_292 ();
 sg13g2_fill_2 FILLER_19_300 ();
 sg13g2_fill_1 FILLER_19_331 ();
 sg13g2_fill_1 FILLER_19_338 ();
 sg13g2_fill_2 FILLER_19_361 ();
 sg13g2_fill_1 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_4 FILLER_20_14 ();
 sg13g2_fill_1 FILLER_20_44 ();
 sg13g2_fill_1 FILLER_20_59 ();
 sg13g2_fill_2 FILLER_20_85 ();
 sg13g2_fill_1 FILLER_20_107 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_4 FILLER_20_119 ();
 sg13g2_fill_1 FILLER_20_141 ();
 sg13g2_decap_8 FILLER_20_145 ();
 sg13g2_fill_1 FILLER_20_178 ();
 sg13g2_fill_1 FILLER_20_185 ();
 sg13g2_fill_1 FILLER_20_191 ();
 sg13g2_fill_2 FILLER_20_200 ();
 sg13g2_fill_2 FILLER_20_216 ();
 sg13g2_decap_8 FILLER_20_236 ();
 sg13g2_fill_2 FILLER_20_243 ();
 sg13g2_fill_1 FILLER_20_245 ();
 sg13g2_fill_1 FILLER_20_281 ();
 sg13g2_fill_2 FILLER_20_303 ();
 sg13g2_fill_1 FILLER_20_315 ();
 sg13g2_fill_2 FILLER_20_398 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_fill_1 FILLER_21_28 ();
 sg13g2_fill_2 FILLER_21_69 ();
 sg13g2_fill_1 FILLER_21_71 ();
 sg13g2_fill_2 FILLER_21_90 ();
 sg13g2_fill_1 FILLER_21_92 ();
 sg13g2_fill_2 FILLER_21_105 ();
 sg13g2_fill_1 FILLER_21_127 ();
 sg13g2_fill_2 FILLER_21_132 ();
 sg13g2_fill_1 FILLER_21_145 ();
 sg13g2_fill_1 FILLER_21_159 ();
 sg13g2_fill_2 FILLER_21_163 ();
 sg13g2_fill_1 FILLER_21_165 ();
 sg13g2_decap_8 FILLER_21_170 ();
 sg13g2_fill_2 FILLER_21_177 ();
 sg13g2_fill_1 FILLER_21_179 ();
 sg13g2_fill_1 FILLER_21_196 ();
 sg13g2_decap_4 FILLER_21_246 ();
 sg13g2_fill_1 FILLER_21_250 ();
 sg13g2_decap_4 FILLER_21_256 ();
 sg13g2_fill_1 FILLER_21_260 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_fill_1 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_300 ();
 sg13g2_fill_2 FILLER_21_307 ();
 sg13g2_fill_1 FILLER_21_309 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_fill_1 FILLER_22_82 ();
 sg13g2_fill_1 FILLER_22_106 ();
 sg13g2_fill_2 FILLER_22_141 ();
 sg13g2_fill_1 FILLER_22_143 ();
 sg13g2_fill_1 FILLER_22_154 ();
 sg13g2_fill_2 FILLER_22_181 ();
 sg13g2_fill_2 FILLER_22_261 ();
 sg13g2_fill_1 FILLER_22_263 ();
 sg13g2_decap_8 FILLER_22_334 ();
 sg13g2_fill_2 FILLER_22_341 ();
 sg13g2_fill_1 FILLER_22_381 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_fill_1 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_58 ();
 sg13g2_decap_8 FILLER_23_75 ();
 sg13g2_fill_1 FILLER_23_82 ();
 sg13g2_fill_2 FILLER_23_91 ();
 sg13g2_fill_1 FILLER_23_93 ();
 sg13g2_decap_8 FILLER_23_104 ();
 sg13g2_fill_1 FILLER_23_111 ();
 sg13g2_decap_8 FILLER_23_123 ();
 sg13g2_decap_8 FILLER_23_130 ();
 sg13g2_decap_4 FILLER_23_137 ();
 sg13g2_fill_1 FILLER_23_154 ();
 sg13g2_fill_2 FILLER_23_186 ();
 sg13g2_fill_2 FILLER_23_246 ();
 sg13g2_fill_1 FILLER_23_248 ();
 sg13g2_fill_1 FILLER_23_294 ();
 sg13g2_fill_2 FILLER_23_309 ();
 sg13g2_decap_8 FILLER_23_319 ();
 sg13g2_fill_1 FILLER_23_326 ();
 sg13g2_fill_1 FILLER_23_340 ();
 sg13g2_fill_2 FILLER_23_398 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_fill_1 FILLER_24_42 ();
 sg13g2_fill_2 FILLER_24_47 ();
 sg13g2_fill_1 FILLER_24_49 ();
 sg13g2_fill_2 FILLER_24_86 ();
 sg13g2_fill_2 FILLER_24_96 ();
 sg13g2_fill_2 FILLER_24_114 ();
 sg13g2_fill_2 FILLER_24_133 ();
 sg13g2_fill_2 FILLER_24_213 ();
 sg13g2_fill_2 FILLER_24_270 ();
 sg13g2_fill_2 FILLER_24_289 ();
 sg13g2_fill_2 FILLER_24_322 ();
 sg13g2_fill_1 FILLER_24_324 ();
 sg13g2_fill_2 FILLER_24_362 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_4 FILLER_25_35 ();
 sg13g2_fill_1 FILLER_25_39 ();
 sg13g2_fill_1 FILLER_25_48 ();
 sg13g2_fill_2 FILLER_25_65 ();
 sg13g2_fill_1 FILLER_25_72 ();
 sg13g2_fill_2 FILLER_25_83 ();
 sg13g2_fill_1 FILLER_25_85 ();
 sg13g2_decap_8 FILLER_25_113 ();
 sg13g2_decap_4 FILLER_25_142 ();
 sg13g2_fill_2 FILLER_25_151 ();
 sg13g2_decap_8 FILLER_25_159 ();
 sg13g2_fill_2 FILLER_25_166 ();
 sg13g2_fill_1 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_173 ();
 sg13g2_fill_1 FILLER_25_180 ();
 sg13g2_fill_1 FILLER_25_187 ();
 sg13g2_fill_2 FILLER_25_197 ();
 sg13g2_fill_1 FILLER_25_199 ();
 sg13g2_fill_1 FILLER_25_209 ();
 sg13g2_fill_2 FILLER_25_215 ();
 sg13g2_decap_4 FILLER_25_244 ();
 sg13g2_fill_2 FILLER_25_248 ();
 sg13g2_fill_1 FILLER_25_260 ();
 sg13g2_fill_2 FILLER_25_272 ();
 sg13g2_fill_2 FILLER_25_290 ();
 sg13g2_fill_1 FILLER_25_292 ();
 sg13g2_fill_2 FILLER_25_349 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_4 FILLER_26_21 ();
 sg13g2_fill_1 FILLER_26_25 ();
 sg13g2_fill_1 FILLER_26_52 ();
 sg13g2_fill_1 FILLER_26_62 ();
 sg13g2_fill_2 FILLER_26_95 ();
 sg13g2_fill_2 FILLER_26_113 ();
 sg13g2_fill_1 FILLER_26_115 ();
 sg13g2_decap_8 FILLER_26_132 ();
 sg13g2_fill_2 FILLER_26_139 ();
 sg13g2_decap_4 FILLER_26_153 ();
 sg13g2_fill_1 FILLER_26_157 ();
 sg13g2_fill_2 FILLER_26_164 ();
 sg13g2_fill_1 FILLER_26_166 ();
 sg13g2_fill_1 FILLER_26_190 ();
 sg13g2_decap_8 FILLER_26_267 ();
 sg13g2_fill_2 FILLER_26_274 ();
 sg13g2_fill_1 FILLER_26_276 ();
 sg13g2_fill_2 FILLER_26_300 ();
 sg13g2_fill_1 FILLER_26_302 ();
 sg13g2_fill_1 FILLER_26_308 ();
 sg13g2_fill_1 FILLER_26_321 ();
 sg13g2_fill_1 FILLER_26_335 ();
 sg13g2_fill_1 FILLER_26_342 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_fill_2 FILLER_27_35 ();
 sg13g2_fill_2 FILLER_27_45 ();
 sg13g2_fill_1 FILLER_27_47 ();
 sg13g2_fill_1 FILLER_27_69 ();
 sg13g2_fill_1 FILLER_27_75 ();
 sg13g2_decap_4 FILLER_27_105 ();
 sg13g2_fill_1 FILLER_27_109 ();
 sg13g2_fill_2 FILLER_27_127 ();
 sg13g2_decap_8 FILLER_27_145 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_fill_2 FILLER_27_172 ();
 sg13g2_fill_1 FILLER_27_174 ();
 sg13g2_fill_2 FILLER_27_192 ();
 sg13g2_fill_1 FILLER_27_194 ();
 sg13g2_fill_2 FILLER_27_222 ();
 sg13g2_fill_1 FILLER_27_224 ();
 sg13g2_decap_4 FILLER_27_244 ();
 sg13g2_fill_1 FILLER_27_248 ();
 sg13g2_fill_1 FILLER_27_253 ();
 sg13g2_fill_2 FILLER_27_258 ();
 sg13g2_fill_1 FILLER_27_260 ();
 sg13g2_decap_8 FILLER_27_286 ();
 sg13g2_fill_1 FILLER_27_293 ();
 sg13g2_fill_1 FILLER_27_352 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_4 FILLER_28_21 ();
 sg13g2_fill_1 FILLER_28_25 ();
 sg13g2_fill_1 FILLER_28_52 ();
 sg13g2_fill_1 FILLER_28_64 ();
 sg13g2_decap_4 FILLER_28_70 ();
 sg13g2_fill_1 FILLER_28_119 ();
 sg13g2_fill_1 FILLER_28_125 ();
 sg13g2_decap_4 FILLER_28_153 ();
 sg13g2_decap_8 FILLER_28_169 ();
 sg13g2_fill_2 FILLER_28_176 ();
 sg13g2_fill_1 FILLER_28_178 ();
 sg13g2_decap_4 FILLER_28_200 ();
 sg13g2_fill_2 FILLER_28_204 ();
 sg13g2_fill_2 FILLER_28_212 ();
 sg13g2_fill_1 FILLER_28_214 ();
 sg13g2_fill_2 FILLER_28_223 ();
 sg13g2_fill_1 FILLER_28_225 ();
 sg13g2_fill_2 FILLER_28_247 ();
 sg13g2_fill_1 FILLER_28_249 ();
 sg13g2_decap_4 FILLER_28_256 ();
 sg13g2_fill_2 FILLER_28_286 ();
 sg13g2_fill_1 FILLER_28_288 ();
 sg13g2_fill_2 FILLER_28_307 ();
 sg13g2_fill_1 FILLER_28_320 ();
 sg13g2_fill_2 FILLER_28_375 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_fill_2 FILLER_29_28 ();
 sg13g2_decap_4 FILLER_29_47 ();
 sg13g2_decap_4 FILLER_29_70 ();
 sg13g2_fill_2 FILLER_29_74 ();
 sg13g2_decap_8 FILLER_29_94 ();
 sg13g2_fill_2 FILLER_29_112 ();
 sg13g2_fill_2 FILLER_29_120 ();
 sg13g2_decap_4 FILLER_29_144 ();
 sg13g2_fill_2 FILLER_29_148 ();
 sg13g2_fill_1 FILLER_29_201 ();
 sg13g2_fill_2 FILLER_29_212 ();
 sg13g2_fill_1 FILLER_29_214 ();
 sg13g2_decap_8 FILLER_29_241 ();
 sg13g2_decap_4 FILLER_29_248 ();
 sg13g2_decap_8 FILLER_29_257 ();
 sg13g2_fill_2 FILLER_29_264 ();
 sg13g2_fill_1 FILLER_29_266 ();
 sg13g2_decap_4 FILLER_29_282 ();
 sg13g2_decap_4 FILLER_29_291 ();
 sg13g2_fill_1 FILLER_29_295 ();
 sg13g2_fill_2 FILLER_29_315 ();
 sg13g2_fill_2 FILLER_29_350 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_fill_1 FILLER_30_56 ();
 sg13g2_fill_2 FILLER_30_78 ();
 sg13g2_fill_1 FILLER_30_80 ();
 sg13g2_fill_2 FILLER_30_101 ();
 sg13g2_fill_1 FILLER_30_103 ();
 sg13g2_fill_2 FILLER_30_109 ();
 sg13g2_fill_1 FILLER_30_111 ();
 sg13g2_fill_2 FILLER_30_123 ();
 sg13g2_decap_8 FILLER_30_141 ();
 sg13g2_decap_8 FILLER_30_148 ();
 sg13g2_decap_4 FILLER_30_155 ();
 sg13g2_fill_2 FILLER_30_159 ();
 sg13g2_fill_2 FILLER_30_175 ();
 sg13g2_fill_1 FILLER_30_177 ();
 sg13g2_decap_4 FILLER_30_193 ();
 sg13g2_fill_2 FILLER_30_197 ();
 sg13g2_fill_2 FILLER_30_204 ();
 sg13g2_fill_1 FILLER_30_206 ();
 sg13g2_decap_8 FILLER_30_215 ();
 sg13g2_decap_8 FILLER_30_222 ();
 sg13g2_fill_2 FILLER_30_229 ();
 sg13g2_fill_1 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_274 ();
 sg13g2_decap_4 FILLER_30_281 ();
 sg13g2_fill_2 FILLER_30_285 ();
 sg13g2_fill_1 FILLER_30_291 ();
 sg13g2_decap_4 FILLER_30_297 ();
 sg13g2_decap_4 FILLER_30_310 ();
 sg13g2_fill_2 FILLER_30_314 ();
 sg13g2_fill_1 FILLER_30_378 ();
 sg13g2_fill_1 FILLER_30_388 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_4 FILLER_31_21 ();
 sg13g2_fill_2 FILLER_31_25 ();
 sg13g2_fill_2 FILLER_31_52 ();
 sg13g2_fill_2 FILLER_31_95 ();
 sg13g2_fill_1 FILLER_31_117 ();
 sg13g2_fill_2 FILLER_31_124 ();
 sg13g2_fill_1 FILLER_31_126 ();
 sg13g2_fill_1 FILLER_31_152 ();
 sg13g2_fill_2 FILLER_31_174 ();
 sg13g2_decap_8 FILLER_31_181 ();
 sg13g2_decap_8 FILLER_31_188 ();
 sg13g2_fill_1 FILLER_31_195 ();
 sg13g2_decap_4 FILLER_31_211 ();
 sg13g2_fill_1 FILLER_31_220 ();
 sg13g2_fill_1 FILLER_31_226 ();
 sg13g2_decap_8 FILLER_31_241 ();
 sg13g2_fill_1 FILLER_31_268 ();
 sg13g2_fill_2 FILLER_31_275 ();
 sg13g2_decap_4 FILLER_31_283 ();
 sg13g2_decap_4 FILLER_31_300 ();
 sg13g2_fill_1 FILLER_31_304 ();
 sg13g2_fill_2 FILLER_31_352 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_fill_1 FILLER_32_28 ();
 sg13g2_decap_4 FILLER_32_65 ();
 sg13g2_decap_8 FILLER_32_74 ();
 sg13g2_decap_4 FILLER_32_93 ();
 sg13g2_fill_1 FILLER_32_101 ();
 sg13g2_fill_1 FILLER_32_107 ();
 sg13g2_decap_8 FILLER_32_118 ();
 sg13g2_decap_8 FILLER_32_129 ();
 sg13g2_fill_1 FILLER_32_136 ();
 sg13g2_fill_1 FILLER_32_142 ();
 sg13g2_decap_8 FILLER_32_148 ();
 sg13g2_decap_4 FILLER_32_155 ();
 sg13g2_decap_4 FILLER_32_177 ();
 sg13g2_fill_2 FILLER_32_199 ();
 sg13g2_fill_1 FILLER_32_201 ();
 sg13g2_decap_4 FILLER_32_219 ();
 sg13g2_fill_2 FILLER_32_229 ();
 sg13g2_fill_1 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_244 ();
 sg13g2_fill_2 FILLER_32_274 ();
 sg13g2_fill_1 FILLER_32_276 ();
 sg13g2_decap_4 FILLER_32_311 ();
 sg13g2_fill_2 FILLER_32_315 ();
 sg13g2_fill_2 FILLER_32_343 ();
 sg13g2_fill_2 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_4 FILLER_33_28 ();
 sg13g2_fill_1 FILLER_33_32 ();
 sg13g2_decap_8 FILLER_33_46 ();
 sg13g2_fill_2 FILLER_33_53 ();
 sg13g2_fill_1 FILLER_33_68 ();
 sg13g2_fill_2 FILLER_33_83 ();
 sg13g2_fill_1 FILLER_33_85 ();
 sg13g2_fill_2 FILLER_33_123 ();
 sg13g2_fill_2 FILLER_33_129 ();
 sg13g2_fill_2 FILLER_33_146 ();
 sg13g2_fill_2 FILLER_33_159 ();
 sg13g2_fill_1 FILLER_33_161 ();
 sg13g2_fill_2 FILLER_33_175 ();
 sg13g2_fill_2 FILLER_33_186 ();
 sg13g2_fill_1 FILLER_33_188 ();
 sg13g2_fill_2 FILLER_33_198 ();
 sg13g2_fill_2 FILLER_33_204 ();
 sg13g2_fill_2 FILLER_33_215 ();
 sg13g2_fill_1 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_222 ();
 sg13g2_fill_2 FILLER_33_234 ();
 sg13g2_fill_1 FILLER_33_236 ();
 sg13g2_decap_4 FILLER_33_252 ();
 sg13g2_fill_2 FILLER_33_256 ();
 sg13g2_decap_4 FILLER_33_262 ();
 sg13g2_fill_2 FILLER_33_266 ();
 sg13g2_fill_2 FILLER_33_296 ();
 sg13g2_decap_4 FILLER_33_317 ();
 sg13g2_fill_2 FILLER_33_342 ();
 sg13g2_fill_1 FILLER_33_357 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_4 FILLER_34_42 ();
 sg13g2_fill_1 FILLER_34_46 ();
 sg13g2_fill_1 FILLER_34_90 ();
 sg13g2_fill_1 FILLER_34_119 ();
 sg13g2_fill_2 FILLER_34_144 ();
 sg13g2_fill_1 FILLER_34_146 ();
 sg13g2_fill_2 FILLER_34_167 ();
 sg13g2_fill_2 FILLER_34_173 ();
 sg13g2_fill_1 FILLER_34_175 ();
 sg13g2_fill_1 FILLER_34_188 ();
 sg13g2_fill_2 FILLER_34_200 ();
 sg13g2_fill_1 FILLER_34_207 ();
 sg13g2_fill_2 FILLER_34_214 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_fill_1 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_237 ();
 sg13g2_decap_4 FILLER_34_244 ();
 sg13g2_fill_1 FILLER_34_248 ();
 sg13g2_decap_4 FILLER_34_288 ();
 sg13g2_fill_1 FILLER_34_292 ();
 sg13g2_fill_2 FILLER_34_298 ();
 sg13g2_decap_8 FILLER_34_310 ();
 sg13g2_fill_2 FILLER_34_317 ();
 sg13g2_fill_2 FILLER_34_332 ();
 sg13g2_fill_1 FILLER_34_334 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_4 FILLER_35_49 ();
 sg13g2_fill_1 FILLER_35_53 ();
 sg13g2_fill_2 FILLER_35_58 ();
 sg13g2_fill_1 FILLER_35_60 ();
 sg13g2_fill_1 FILLER_35_65 ();
 sg13g2_fill_2 FILLER_35_115 ();
 sg13g2_fill_2 FILLER_35_139 ();
 sg13g2_fill_1 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_169 ();
 sg13g2_fill_2 FILLER_35_176 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_fill_2 FILLER_35_205 ();
 sg13g2_decap_4 FILLER_35_217 ();
 sg13g2_fill_2 FILLER_35_226 ();
 sg13g2_decap_4 FILLER_35_262 ();
 sg13g2_fill_2 FILLER_35_266 ();
 sg13g2_decap_4 FILLER_35_278 ();
 sg13g2_fill_2 FILLER_35_292 ();
 sg13g2_fill_1 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_319 ();
 sg13g2_decap_8 FILLER_35_326 ();
 sg13g2_decap_4 FILLER_35_333 ();
 sg13g2_fill_2 FILLER_35_337 ();
 sg13g2_fill_1 FILLER_35_373 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_fill_1 FILLER_36_49 ();
 sg13g2_fill_2 FILLER_36_76 ();
 sg13g2_fill_2 FILLER_36_147 ();
 sg13g2_fill_2 FILLER_36_152 ();
 sg13g2_fill_2 FILLER_36_164 ();
 sg13g2_fill_1 FILLER_36_166 ();
 sg13g2_fill_2 FILLER_36_172 ();
 sg13g2_fill_1 FILLER_36_174 ();
 sg13g2_fill_1 FILLER_36_201 ();
 sg13g2_fill_1 FILLER_36_208 ();
 sg13g2_fill_1 FILLER_36_214 ();
 sg13g2_fill_1 FILLER_36_219 ();
 sg13g2_decap_8 FILLER_36_240 ();
 sg13g2_fill_1 FILLER_36_247 ();
 sg13g2_decap_4 FILLER_36_258 ();
 sg13g2_fill_2 FILLER_36_268 ();
 sg13g2_decap_4 FILLER_36_283 ();
 sg13g2_fill_1 FILLER_36_287 ();
 sg13g2_fill_1 FILLER_36_294 ();
 sg13g2_decap_8 FILLER_36_309 ();
 sg13g2_fill_2 FILLER_36_316 ();
 sg13g2_fill_2 FILLER_36_349 ();
 sg13g2_fill_1 FILLER_36_377 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_fill_1 FILLER_37_98 ();
 sg13g2_fill_2 FILLER_37_108 ();
 sg13g2_fill_1 FILLER_37_110 ();
 sg13g2_fill_1 FILLER_37_119 ();
 sg13g2_fill_1 FILLER_37_133 ();
 sg13g2_fill_1 FILLER_37_151 ();
 sg13g2_decap_8 FILLER_37_160 ();
 sg13g2_decap_4 FILLER_37_167 ();
 sg13g2_fill_2 FILLER_37_193 ();
 sg13g2_fill_1 FILLER_37_246 ();
 sg13g2_fill_1 FILLER_37_263 ();
 sg13g2_fill_2 FILLER_37_284 ();
 sg13g2_decap_8 FILLER_37_311 ();
 sg13g2_fill_1 FILLER_37_318 ();
 sg13g2_fill_2 FILLER_37_327 ();
 sg13g2_fill_1 FILLER_37_346 ();
 sg13g2_fill_1 FILLER_37_355 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_fill_1 FILLER_38_108 ();
 sg13g2_fill_1 FILLER_38_143 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_fill_2 FILLER_38_199 ();
 sg13g2_fill_1 FILLER_38_201 ();
 sg13g2_fill_2 FILLER_38_207 ();
 sg13g2_decap_8 FILLER_38_214 ();
 sg13g2_decap_8 FILLER_38_221 ();
 sg13g2_decap_8 FILLER_38_237 ();
 sg13g2_fill_1 FILLER_38_244 ();
 sg13g2_fill_1 FILLER_38_250 ();
 sg13g2_fill_1 FILLER_38_271 ();
 sg13g2_fill_1 FILLER_38_276 ();
 sg13g2_decap_4 FILLER_38_281 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_decap_4 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_307 ();
 sg13g2_fill_2 FILLER_38_338 ();
 sg13g2_decap_4 FILLER_38_390 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net4;
 assign uio_oe[1] = net5;
 assign uio_oe[2] = net6;
 assign uio_oe[3] = net7;
 assign uio_oe[4] = net8;
 assign uio_oe[5] = net9;
 assign uio_oe[6] = net10;
 assign uio_oe[7] = net11;
 assign uio_out[0] = net12;
 assign uio_out[1] = net13;
 assign uio_out[2] = net14;
 assign uio_out[3] = net15;
 assign uio_out[4] = net16;
 assign uio_out[5] = net17;
 assign uio_out[6] = net18;
 assign uio_out[7] = net19;
endmodule

module tt_um_shuangyu_top (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire \inst_calculator.bcd[0] ;
 wire \inst_calculator.denominator[0] ;
 wire \inst_calculator.denominator[1] ;
 wire \inst_calculator.denominator[2] ;
 wire \inst_calculator.denominator[3] ;
 wire \inst_calculator.denominator[4] ;
 wire \inst_calculator.denominator[5] ;
 wire \inst_calculator.denominator[6] ;
 wire \inst_calculator.denominator[7] ;
 wire \inst_calculator.denominator[8] ;
 wire \inst_calculator.denominator[9] ;
 wire \inst_calculator.divider_done ;
 wire \inst_calculator.divider_start ;
 wire \inst_calculator.inst_bin2bcd.bin_in[1] ;
 wire \inst_calculator.inst_bin2bcd.bin_in[2] ;
 wire \inst_calculator.inst_bin2bcd.bin_in[3] ;
 wire \inst_calculator.inst_bin2bcd.bin_in[4] ;
 wire \inst_calculator.inst_bin2bcd.bin_in[5] ;
 wire \inst_calculator.inst_bin2bcd.bin_in[6] ;
 wire \inst_calculator.inst_bin2bcd.bin_in[7] ;
 wire \inst_calculator.inst_bin2bcd.bin_in[8] ;
 wire \inst_calculator.inst_bin2bcd.bin_in[9] ;
 wire \inst_calculator.inst_divider.busy ;
 wire \inst_calculator.inst_divider.d[0] ;
 wire \inst_calculator.inst_divider.d[1] ;
 wire \inst_calculator.inst_divider.d[2] ;
 wire \inst_calculator.inst_divider.d[3] ;
 wire \inst_calculator.inst_divider.d[4] ;
 wire \inst_calculator.inst_divider.d[5] ;
 wire \inst_calculator.inst_divider.d[6] ;
 wire \inst_calculator.inst_divider.d[7] ;
 wire \inst_calculator.inst_divider.d[8] ;
 wire \inst_calculator.inst_divider.d[9] ;
 wire \inst_calculator.inst_divider.n[0] ;
 wire \inst_calculator.inst_divider.n[1] ;
 wire \inst_calculator.inst_divider.n[2] ;
 wire \inst_calculator.inst_divider.n[3] ;
 wire \inst_calculator.inst_divider.n[4] ;
 wire \inst_calculator.inst_divider.n[5] ;
 wire \inst_calculator.inst_divider.n[6] ;
 wire \inst_calculator.inst_divider.n[7] ;
 wire \inst_calculator.inst_divider.n[8] ;
 wire \inst_calculator.inst_divider.n[9] ;
 wire \inst_calculator.inst_divider.numerator[0] ;
 wire \inst_calculator.inst_divider.numerator[1] ;
 wire \inst_calculator.inst_divider.numerator[2] ;
 wire \inst_calculator.inst_divider.numerator[3] ;
 wire \inst_calculator.inst_divider.numerator[4] ;
 wire \inst_calculator.inst_divider.numerator[5] ;
 wire \inst_calculator.inst_divider.numerator[6] ;
 wire \inst_calculator.inst_divider.numerator[7] ;
 wire \inst_calculator.inst_divider.numerator[8] ;
 wire \inst_calculator.inst_divider.numerator[9] ;
 wire \inst_calculator.inst_divider.q[0] ;
 wire \inst_calculator.inst_divider.q[1] ;
 wire \inst_calculator.inst_divider.q[2] ;
 wire \inst_calculator.inst_divider.q[3] ;
 wire \inst_calculator.inst_divider.q[4] ;
 wire \inst_calculator.inst_divider.q[5] ;
 wire \inst_calculator.inst_divider.q[6] ;
 wire \inst_calculator.inst_divider.q[7] ;
 wire \inst_calculator.inst_divider.q[8] ;
 wire \inst_calculator.inst_divider.q[9] ;
 wire \inst_calculator.inst_drive.cnt0[0] ;
 wire \inst_calculator.inst_drive.cnt0[10] ;
 wire \inst_calculator.inst_drive.cnt0[11] ;
 wire \inst_calculator.inst_drive.cnt0[12] ;
 wire \inst_calculator.inst_drive.cnt0[13] ;
 wire \inst_calculator.inst_drive.cnt0[1] ;
 wire \inst_calculator.inst_drive.cnt0[2] ;
 wire \inst_calculator.inst_drive.cnt0[3] ;
 wire \inst_calculator.inst_drive.cnt0[4] ;
 wire \inst_calculator.inst_drive.cnt0[5] ;
 wire \inst_calculator.inst_drive.cnt0[6] ;
 wire \inst_calculator.inst_drive.cnt0[7] ;
 wire \inst_calculator.inst_drive.cnt0[8] ;
 wire \inst_calculator.inst_drive.cnt0[9] ;
 wire \inst_calculator.inst_drive.cnt_sel[0] ;
 wire \inst_calculator.inst_drive.cnt_sel[1] ;
 wire \inst_calculator.inst_drive.flag ;
 wire \inst_calculator.inst_drive.num_disp[0] ;
 wire \inst_calculator.inst_drive.num_disp[1] ;
 wire \inst_calculator.inst_drive.num_disp[2] ;
 wire \inst_calculator.inst_drive.num_disp[3] ;
 wire \inst_calculator.inst_keypad_encoder.key[0] ;
 wire \inst_calculator.inst_keypad_encoder.key[1] ;
 wire \inst_calculator.inst_keypad_encoder.key[2] ;
 wire \inst_calculator.inst_keypad_encoder.key[3] ;
 wire \inst_calculator.inst_keypad_encoder.rows[0] ;
 wire \inst_calculator.inst_keypad_encoder.rows[1] ;
 wire \inst_calculator.inst_keypad_encoder.rows[2] ;
 wire \inst_calculator.inst_keypad_encoder.rows[3] ;
 wire \inst_calculator.inst_keypad_poller.clk_counter[0] ;
 wire \inst_calculator.inst_keypad_poller.clk_counter[10] ;
 wire \inst_calculator.inst_keypad_poller.clk_counter[11] ;
 wire \inst_calculator.inst_keypad_poller.clk_counter[12] ;
 wire \inst_calculator.inst_keypad_poller.clk_counter[13] ;
 wire \inst_calculator.inst_keypad_poller.clk_counter[14] ;
 wire \inst_calculator.inst_keypad_poller.clk_counter[15] ;
 wire \inst_calculator.inst_keypad_poller.clk_counter[16] ;
 wire \inst_calculator.inst_keypad_poller.clk_counter[1] ;
 wire \inst_calculator.inst_keypad_poller.clk_counter[2] ;
 wire \inst_calculator.inst_keypad_poller.clk_counter[3] ;
 wire \inst_calculator.inst_keypad_poller.clk_counter[4] ;
 wire \inst_calculator.inst_keypad_poller.clk_counter[5] ;
 wire \inst_calculator.inst_keypad_poller.clk_counter[6] ;
 wire \inst_calculator.inst_keypad_poller.clk_counter[7] ;
 wire \inst_calculator.inst_keypad_poller.clk_counter[8] ;
 wire \inst_calculator.inst_keypad_poller.clk_counter[9] ;
 wire \inst_calculator.inst_keypad_poller.key_pressed ;
 wire \inst_calculator.inst_keypad_poller.state[0] ;
 wire \inst_calculator.inst_keypad_poller.state[1] ;
 wire \inst_calculator.inst_keypad_poller.state[2] ;
 wire \inst_calculator.inst_keypad_poller.state[3] ;
 wire \inst_calculator.inst_keypad_poller.state[4] ;
 wire \inst_calculator.inst_keypad_poller.state[5] ;
 wire \inst_calculator.key_pressed_prev ;
 wire \inst_calculator.reg_arg[0] ;
 wire \inst_calculator.reg_arg[1] ;
 wire \inst_calculator.reg_arg[2] ;
 wire \inst_calculator.reg_arg[3] ;
 wire \inst_calculator.reg_arg[4] ;
 wire \inst_calculator.reg_arg[5] ;
 wire \inst_calculator.reg_arg[6] ;
 wire \inst_calculator.reg_arg[7] ;
 wire \inst_calculator.reg_arg[8] ;
 wire \inst_calculator.reg_arg[9] ;
 wire \inst_calculator.reg_operator[0] ;
 wire \inst_calculator.reg_operator[1] ;
 wire \inst_calculator.reg_operator_next[0] ;
 wire \inst_calculator.reg_operator_next[1] ;
 wire \inst_calculator.reg_result[0] ;
 wire \inst_calculator.reg_result[1] ;
 wire \inst_calculator.reg_result[2] ;
 wire \inst_calculator.reg_result[3] ;
 wire \inst_calculator.reg_result[4] ;
 wire \inst_calculator.reg_result[5] ;
 wire \inst_calculator.reg_result[6] ;
 wire \inst_calculator.reg_result[7] ;
 wire \inst_calculator.reg_result[8] ;
 wire \inst_calculator.reg_result[9] ;
 wire \inst_calculator.state[0] ;
 wire \inst_calculator.state[10] ;
 wire \inst_calculator.state[1] ;
 wire \inst_calculator.state[2] ;
 wire \inst_calculator.state[3] ;
 wire \inst_calculator.state[4] ;
 wire \inst_calculator.state[5] ;
 wire \inst_calculator.state[6] ;
 wire \inst_calculator.state[7] ;
 wire \inst_calculator.state[8] ;
 wire \inst_calculator.state[9] ;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net6;
 wire clknet_0_clk;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;

 sg13g2_inv_1 _1297_ (.Y(_0559_),
    .A(net134));
 sg13g2_inv_1 _1298_ (.Y(_0560_),
    .A(net151));
 sg13g2_inv_1 _1299_ (.Y(_0561_),
    .A(uio_out[7]));
 sg13g2_inv_1 _1300_ (.Y(_0562_),
    .A(net308));
 sg13g2_inv_1 _1301_ (.Y(_0563_),
    .A(net190));
 sg13g2_inv_1 _1302_ (.Y(_0564_),
    .A(\inst_calculator.reg_operator[0] ));
 sg13g2_inv_1 _1303_ (.Y(_0565_),
    .A(net110));
 sg13g2_inv_1 _1304_ (.Y(_0566_),
    .A(net357));
 sg13g2_inv_1 _1305_ (.Y(_0567_),
    .A(net145));
 sg13g2_inv_1 _1306_ (.Y(_0568_),
    .A(net314));
 sg13g2_inv_2 _1307_ (.Y(_0569_),
    .A(net316));
 sg13g2_inv_1 _1308_ (.Y(_0570_),
    .A(net319));
 sg13g2_inv_2 _1309_ (.Y(_0571_),
    .A(net320));
 sg13g2_inv_1 _1310_ (.Y(_0572_),
    .A(net324));
 sg13g2_inv_1 _1311_ (.Y(_0573_),
    .A(net102));
 sg13g2_inv_1 _1312_ (.Y(_0574_),
    .A(\inst_calculator.inst_keypad_poller.clk_counter[5] ));
 sg13g2_inv_1 _1313_ (.Y(_0575_),
    .A(\inst_calculator.inst_keypad_poller.clk_counter[9] ));
 sg13g2_inv_1 _1314_ (.Y(_0576_),
    .A(net165));
 sg13g2_inv_1 _1315_ (.Y(_0577_),
    .A(net162));
 sg13g2_inv_1 _1316_ (.Y(_0578_),
    .A(\inst_calculator.inst_divider.busy ));
 sg13g2_inv_1 _1317_ (.Y(_0579_),
    .A(net425));
 sg13g2_inv_1 _1318_ (.Y(_0580_),
    .A(net416));
 sg13g2_inv_2 _1319_ (.Y(_0581_),
    .A(net438));
 sg13g2_inv_2 _1320_ (.Y(_0582_),
    .A(net291));
 sg13g2_inv_1 _1321_ (.Y(_0583_),
    .A(net289));
 sg13g2_inv_1 _1322_ (.Y(_0584_),
    .A(\inst_calculator.inst_divider.q[3] ));
 sg13g2_inv_1 _1323_ (.Y(_0585_),
    .A(\inst_calculator.inst_drive.num_disp[0] ));
 sg13g2_inv_1 _1324_ (.Y(_0586_),
    .A(\inst_calculator.inst_drive.cnt0[11] ));
 sg13g2_inv_1 _1325_ (.Y(_0587_),
    .A(net355));
 sg13g2_inv_1 _1326_ (.Y(_0588_),
    .A(net136));
 sg13g2_inv_1 _1327_ (.Y(_0589_),
    .A(_0037_));
 sg13g2_inv_1 _1328_ (.Y(_0590_),
    .A(_0036_));
 sg13g2_inv_1 _1329_ (.Y(_0591_),
    .A(_0038_));
 sg13g2_inv_1 _1330_ (.Y(_0592_),
    .A(_0040_));
 sg13g2_inv_1 _1331_ (.Y(_0593_),
    .A(_0041_));
 sg13g2_inv_1 _1332_ (.Y(_0594_),
    .A(_0042_));
 sg13g2_inv_1 _1333_ (.Y(_0595_),
    .A(_0043_));
 sg13g2_inv_1 _1334_ (.Y(_0596_),
    .A(_0044_));
 sg13g2_o21ai_1 _1335_ (.B1(_0566_),
    .Y(_0597_),
    .A1(net312),
    .A2(\inst_calculator.inst_keypad_encoder.key[2] ));
 sg13g2_nor2_1 _1336_ (.A(_0567_),
    .B(net119),
    .Y(_0598_));
 sg13g2_nand2_1 _1337_ (.Y(_0599_),
    .A(net171),
    .B(_0598_));
 sg13g2_nor2_1 _1338_ (.A(_0597_),
    .B(_0599_),
    .Y(_0600_));
 sg13g2_or2_1 _1339_ (.X(_0601_),
    .B(_0599_),
    .A(_0597_));
 sg13g2_nand2_1 _1340_ (.Y(_0602_),
    .A(net364),
    .B(\inst_calculator.inst_keypad_encoder.key[2] ));
 sg13g2_nand4_1 _1341_ (.B(net364),
    .C(net381),
    .A(net312),
    .Y(_0068_),
    .D(_0600_));
 sg13g2_or2_1 _1342_ (.X(_0603_),
    .B(\inst_calculator.inst_drive.num_disp[1] ),
    .A(\inst_calculator.inst_drive.num_disp[2] ));
 sg13g2_nand2b_1 _1343_ (.Y(_0604_),
    .B(net426),
    .A_N(net418));
 sg13g2_nand3_1 _1344_ (.B(net441),
    .C(net108),
    .A(net426),
    .Y(_0605_));
 sg13g2_nor2_1 _1345_ (.A(net418),
    .B(_0605_),
    .Y(_0606_));
 sg13g2_nor2_1 _1346_ (.A(\inst_calculator.inst_drive.num_disp[2] ),
    .B(\inst_calculator.inst_drive.num_disp[3] ),
    .Y(_0607_));
 sg13g2_a221oi_1 _1347_ (.B2(net90),
    .C1(_0606_),
    .B1(_0607_),
    .A1(\inst_calculator.inst_drive.num_disp[3] ),
    .Y(_0067_),
    .A2(_0603_));
 sg13g2_nor2b_2 _1348_ (.A(net311),
    .B_N(net405),
    .Y(_0066_));
 sg13g2_nand2b_2 _1349_ (.Y(_0608_),
    .B(net311),
    .A_N(net405));
 sg13g2_inv_1 _1350_ (.Y(_0065_),
    .A(_0608_));
 sg13g2_nor2_2 _1351_ (.A(net405),
    .B(net311),
    .Y(_0064_));
 sg13g2_nor4_2 _1352_ (.A(net2),
    .B(net1),
    .C(net4),
    .Y(_0609_),
    .D(net3));
 sg13g2_nand2_1 _1353_ (.Y(_0063_),
    .A(net107),
    .B(_0609_));
 sg13g2_nand2b_1 _1354_ (.Y(_0610_),
    .B(net298),
    .A_N(net305));
 sg13g2_nand2_1 _1355_ (.Y(_0611_),
    .A(net298),
    .B(_0564_));
 sg13g2_nand2_1 _1356_ (.Y(_0612_),
    .A(net303),
    .B(net409));
 sg13g2_nand3_1 _1357_ (.B(_0611_),
    .C(_0612_),
    .A(_0610_),
    .Y(_0018_));
 sg13g2_nor3_1 _1358_ (.A(\inst_calculator.state[4] ),
    .B(\inst_calculator.state[0] ),
    .C(\inst_calculator.state[7] ),
    .Y(_0613_));
 sg13g2_o21ai_1 _1359_ (.B1(_0598_),
    .Y(_0614_),
    .A1(\inst_calculator.inst_keypad_encoder.key[3] ),
    .A2(_0597_));
 sg13g2_nand2_1 _1360_ (.Y(_0615_),
    .A(net171),
    .B(_0614_));
 sg13g2_nand2_1 _1361_ (.Y(_0019_),
    .A(_0613_),
    .B(net172));
 sg13g2_nand2_1 _1362_ (.Y(_0616_),
    .A(\inst_calculator.inst_keypad_poller.state[5] ),
    .B(_0609_));
 sg13g2_nand2_1 _1363_ (.Y(_0015_),
    .A(_0573_),
    .B(_0616_));
 sg13g2_nand2_1 _1364_ (.Y(_0617_),
    .A(\inst_calculator.inst_keypad_poller.clk_counter[15] ),
    .B(\inst_calculator.inst_keypad_poller.clk_counter[16] ));
 sg13g2_nand2_1 _1365_ (.Y(_0618_),
    .A(\inst_calculator.inst_keypad_poller.clk_counter[7] ),
    .B(\inst_calculator.inst_keypad_poller.clk_counter[10] ));
 sg13g2_nor4_1 _1366_ (.A(\inst_calculator.inst_keypad_poller.clk_counter[11] ),
    .B(\inst_calculator.inst_keypad_poller.clk_counter[14] ),
    .C(_0617_),
    .D(_0618_),
    .Y(_0619_));
 sg13g2_nor4_1 _1367_ (.A(\inst_calculator.inst_keypad_poller.clk_counter[4] ),
    .B(_0574_),
    .C(\inst_calculator.inst_keypad_poller.clk_counter[6] ),
    .D(\inst_calculator.inst_keypad_poller.clk_counter[8] ),
    .Y(_0620_));
 sg13g2_nor2_1 _1368_ (.A(\inst_calculator.inst_keypad_poller.clk_counter[0] ),
    .B(net200),
    .Y(_0621_));
 sg13g2_nor2_1 _1369_ (.A(\inst_calculator.inst_keypad_poller.clk_counter[3] ),
    .B(\inst_calculator.inst_keypad_poller.clk_counter[2] ),
    .Y(_0622_));
 sg13g2_nand3_1 _1370_ (.B(_0621_),
    .C(_0622_),
    .A(_0620_),
    .Y(_0623_));
 sg13g2_nor4_2 _1371_ (.A(_0575_),
    .B(\inst_calculator.inst_keypad_poller.clk_counter[13] ),
    .C(\inst_calculator.inst_keypad_poller.clk_counter[12] ),
    .Y(_0624_),
    .D(_0623_));
 sg13g2_nand2_1 _1372_ (.Y(_0625_),
    .A(_0619_),
    .B(_0624_));
 sg13g2_a21o_1 _1373_ (.A2(_0625_),
    .A1(net160),
    .B1(net263),
    .X(_0014_));
 sg13g2_or4_1 _1374_ (.A(net187),
    .B(\inst_calculator.state[5] ),
    .C(net390),
    .D(net174),
    .X(_0016_));
 sg13g2_nand2b_1 _1375_ (.Y(_0626_),
    .B(\inst_calculator.inst_keypad_poller.clk_counter[11] ),
    .A_N(\inst_calculator.inst_keypad_poller.clk_counter[7] ));
 sg13g2_nand2_1 _1376_ (.Y(_0627_),
    .A(\inst_calculator.inst_keypad_poller.clk_counter[10] ),
    .B(\inst_calculator.inst_keypad_poller.clk_counter[14] ));
 sg13g2_nor4_1 _1377_ (.A(\inst_calculator.inst_keypad_poller.clk_counter[15] ),
    .B(\inst_calculator.inst_keypad_poller.clk_counter[16] ),
    .C(_0626_),
    .D(_0627_),
    .Y(_0628_));
 sg13g2_nand2_1 _1378_ (.Y(_0629_),
    .A(_0624_),
    .B(_0628_));
 sg13g2_a21oi_1 _1379_ (.A1(net178),
    .A2(_0048_),
    .Y(_0630_),
    .B1(_0609_));
 sg13g2_a21o_1 _1380_ (.A2(_0629_),
    .A1(net156),
    .B1(net179),
    .X(_0013_));
 sg13g2_nand2b_1 _1381_ (.Y(_0631_),
    .B(net303),
    .A_N(net409));
 sg13g2_nand2_1 _1382_ (.Y(_0632_),
    .A(net298),
    .B(net305));
 sg13g2_o21ai_1 _1383_ (.B1(net410),
    .Y(_0017_),
    .A1(_0564_),
    .A2(_0632_));
 sg13g2_and3_1 _1384_ (.X(_0002_),
    .A(_0585_),
    .B(net108),
    .C(net104));
 sg13g2_nand2_1 _1385_ (.Y(_0633_),
    .A(net104),
    .B(\inst_calculator.inst_drive.num_disp[3] ));
 sg13g2_nand2_1 _1386_ (.Y(_0634_),
    .A(net418),
    .B(_0002_));
 sg13g2_and2_1 _1387_ (.A(net441),
    .B(_0603_),
    .X(_0635_));
 sg13g2_nand2b_1 _1388_ (.Y(_0636_),
    .B(\inst_calculator.inst_drive.num_disp[2] ),
    .A_N(\inst_calculator.inst_drive.num_disp[1] ));
 sg13g2_a21oi_1 _1389_ (.A1(_0585_),
    .A2(_0636_),
    .Y(_0637_),
    .B1(net418));
 sg13g2_inv_1 _1390_ (.Y(_0638_),
    .A(_0637_));
 sg13g2_o21ai_1 _1391_ (.B1(_0634_),
    .Y(_0000_),
    .A1(net442),
    .A2(_0638_));
 sg13g2_xnor2_1 _1392_ (.Y(_0639_),
    .A(\inst_calculator.inst_drive.num_disp[0] ),
    .B(net108));
 sg13g2_o21ai_1 _1393_ (.B1(_0634_),
    .Y(_0001_),
    .A1(_0604_),
    .A2(_0639_));
 sg13g2_or2_1 _1394_ (.X(_0003_),
    .B(_0000_),
    .A(_0606_));
 sg13g2_o21ai_1 _1395_ (.B1(_0638_),
    .Y(_0004_),
    .A1(net105),
    .A2(_0639_));
 sg13g2_nor2_1 _1396_ (.A(\inst_calculator.inst_drive.num_disp[0] ),
    .B(net108),
    .Y(_0640_));
 sg13g2_o21ai_1 _1397_ (.B1(_0605_),
    .Y(_0641_),
    .A1(\inst_calculator.inst_drive.num_disp[2] ),
    .A2(_0640_));
 sg13g2_inv_1 _1398_ (.Y(_0642_),
    .A(_0641_));
 sg13g2_o21ai_1 _1399_ (.B1(_0634_),
    .Y(_0005_),
    .A1(net418),
    .A2(_0642_));
 sg13g2_and3_1 _1400_ (.X(_0643_),
    .A(net129),
    .B(net183),
    .C(net114));
 sg13g2_and2_1 _1401_ (.A(net186),
    .B(_0643_),
    .X(_0644_));
 sg13g2_nor2_1 _1402_ (.A(net406),
    .B(_0644_),
    .Y(_0645_));
 sg13g2_nor3_1 _1403_ (.A(\inst_calculator.inst_drive.cnt0[7] ),
    .B(\inst_calculator.inst_drive.cnt0[6] ),
    .C(\inst_calculator.inst_drive.cnt0[5] ),
    .Y(_0646_));
 sg13g2_nand4_1 _1404_ (.B(\inst_calculator.inst_drive.cnt0[10] ),
    .C(net401),
    .A(_0586_),
    .Y(_0647_),
    .D(\inst_calculator.inst_drive.cnt0[8] ));
 sg13g2_a21oi_1 _1405_ (.A1(_0645_),
    .A2(_0646_),
    .Y(_0648_),
    .B1(_0647_));
 sg13g2_nor3_2 _1406_ (.A(net197),
    .B(_0587_),
    .C(_0648_),
    .Y(_0649_));
 sg13g2_nor2b_2 _1407_ (.A(_0649_),
    .B_N(net386),
    .Y(_0052_));
 sg13g2_nor2_1 _1408_ (.A(net114),
    .B(net267),
    .Y(_0022_));
 sg13g2_xnor2_1 _1409_ (.Y(_0650_),
    .A(net183),
    .B(net114));
 sg13g2_nor2_1 _1410_ (.A(net267),
    .B(_0650_),
    .Y(_0027_));
 sg13g2_a21oi_1 _1411_ (.A1(\inst_calculator.inst_drive.cnt0[1] ),
    .A2(net114),
    .Y(_0651_),
    .B1(net129));
 sg13g2_nor3_1 _1412_ (.A(_0643_),
    .B(net267),
    .C(net130),
    .Y(_0028_));
 sg13g2_nor2_1 _1413_ (.A(net186),
    .B(_0643_),
    .Y(_0652_));
 sg13g2_nor3_1 _1414_ (.A(_0644_),
    .B(net266),
    .C(_0652_),
    .Y(_0029_));
 sg13g2_and2_1 _1415_ (.A(net406),
    .B(_0644_),
    .X(_0653_));
 sg13g2_nor3_1 _1416_ (.A(_0645_),
    .B(net266),
    .C(_0653_),
    .Y(_0030_));
 sg13g2_xnor2_1 _1417_ (.Y(_0654_),
    .A(net413),
    .B(_0653_));
 sg13g2_nor2_1 _1418_ (.A(net267),
    .B(_0654_),
    .Y(_0031_));
 sg13g2_a21oi_1 _1419_ (.A1(\inst_calculator.inst_drive.cnt0[5] ),
    .A2(_0653_),
    .Y(_0655_),
    .B1(net168));
 sg13g2_and3_1 _1420_ (.X(_0656_),
    .A(net168),
    .B(\inst_calculator.inst_drive.cnt0[5] ),
    .C(_0653_));
 sg13g2_nor3_1 _1421_ (.A(net267),
    .B(net169),
    .C(_0656_),
    .Y(_0032_));
 sg13g2_nor2_1 _1422_ (.A(net362),
    .B(_0656_),
    .Y(_0657_));
 sg13g2_and2_1 _1423_ (.A(net362),
    .B(_0656_),
    .X(_0658_));
 sg13g2_nor3_1 _1424_ (.A(net266),
    .B(net363),
    .C(_0658_),
    .Y(_0033_));
 sg13g2_and2_1 _1425_ (.A(net220),
    .B(_0658_),
    .X(_0659_));
 sg13g2_nor2_1 _1426_ (.A(net220),
    .B(_0658_),
    .Y(_0660_));
 sg13g2_nor3_1 _1427_ (.A(net266),
    .B(_0659_),
    .C(net221),
    .Y(_0034_));
 sg13g2_nor2_1 _1428_ (.A(net372),
    .B(_0659_),
    .Y(_0661_));
 sg13g2_and2_1 _1429_ (.A(net372),
    .B(_0659_),
    .X(_0662_));
 sg13g2_nor3_1 _1430_ (.A(net266),
    .B(_0661_),
    .C(_0662_),
    .Y(_0035_));
 sg13g2_nor2_1 _1431_ (.A(net367),
    .B(_0662_),
    .Y(_0663_));
 sg13g2_and2_1 _1432_ (.A(net367),
    .B(_0662_),
    .X(_0664_));
 sg13g2_nor3_1 _1433_ (.A(net266),
    .B(net368),
    .C(_0664_),
    .Y(_0023_));
 sg13g2_nor2_1 _1434_ (.A(_0587_),
    .B(_0664_),
    .Y(_0665_));
 sg13g2_a21oi_1 _1435_ (.A1(_0587_),
    .A2(_0664_),
    .Y(_0666_),
    .B1(net266));
 sg13g2_nor2b_1 _1436_ (.A(net356),
    .B_N(_0666_),
    .Y(_0024_));
 sg13g2_a21oi_1 _1437_ (.A1(\inst_calculator.inst_drive.cnt0[11] ),
    .A2(_0664_),
    .Y(_0667_),
    .B1(net197));
 sg13g2_and3_1 _1438_ (.X(_0668_),
    .A(net197),
    .B(\inst_calculator.inst_drive.cnt0[11] ),
    .C(_0664_));
 sg13g2_nor3_1 _1439_ (.A(net266),
    .B(net198),
    .C(_0668_),
    .Y(_0025_));
 sg13g2_mux2_1 _1440_ (.A0(_0668_),
    .A1(_0649_),
    .S(net386),
    .X(_0026_));
 sg13g2_nor2b_1 _1441_ (.A(\inst_calculator.inst_bin2bcd.bin_in[8] ),
    .B_N(\inst_calculator.inst_bin2bcd.bin_in[9] ),
    .Y(_0669_));
 sg13g2_mux2_2 _1442_ (.A0(_0037_),
    .A1(_0036_),
    .S(_0669_),
    .X(_0670_));
 sg13g2_nor2_1 _1443_ (.A(\inst_calculator.inst_bin2bcd.bin_in[7] ),
    .B(\inst_calculator.inst_bin2bcd.bin_in[8] ),
    .Y(_0671_));
 sg13g2_xnor2_1 _1444_ (.Y(_0672_),
    .A(_0589_),
    .B(_0671_));
 sg13g2_mux2_1 _1445_ (.A0(_0672_),
    .A1(\inst_calculator.inst_bin2bcd.bin_in[9] ),
    .S(_0670_),
    .X(_0673_));
 sg13g2_o21ai_1 _1446_ (.B1(_0590_),
    .Y(_0674_),
    .A1(_0589_),
    .A2(_0669_));
 sg13g2_o21ai_1 _1447_ (.B1(_0036_),
    .Y(_0675_),
    .A1(_0037_),
    .A2(_0669_));
 sg13g2_nand2_1 _1448_ (.Y(_0676_),
    .A(_0674_),
    .B(_0675_));
 sg13g2_xnor2_1 _1449_ (.Y(_0677_),
    .A(\inst_calculator.inst_bin2bcd.bin_in[7] ),
    .B(\inst_calculator.inst_bin2bcd.bin_in[8] ));
 sg13g2_mux2_2 _1450_ (.A0(_0677_),
    .A1(_0591_),
    .S(_0670_),
    .X(_0678_));
 sg13g2_a21oi_1 _1451_ (.A1(_0674_),
    .A2(_0675_),
    .Y(_0679_),
    .B1(_0039_));
 sg13g2_a21oi_2 _1452_ (.B1(_0673_),
    .Y(_0680_),
    .A2(_0679_),
    .A1(_0678_));
 sg13g2_a21o_2 _1453_ (.A2(_0679_),
    .A1(_0678_),
    .B1(_0673_),
    .X(_0681_));
 sg13g2_xor2_1 _1454_ (.B(_0670_),
    .A(\inst_calculator.inst_bin2bcd.bin_in[7] ),
    .X(_0682_));
 sg13g2_xnor2_1 _1455_ (.Y(_0683_),
    .A(\inst_calculator.inst_bin2bcd.bin_in[7] ),
    .B(_0670_));
 sg13g2_or3_1 _1456_ (.A(\inst_calculator.inst_bin2bcd.bin_in[7] ),
    .B(\inst_calculator.inst_bin2bcd.bin_in[8] ),
    .C(_0670_),
    .X(_0684_));
 sg13g2_o21ai_1 _1457_ (.B1(\inst_calculator.inst_bin2bcd.bin_in[8] ),
    .Y(_0685_),
    .A1(\inst_calculator.inst_bin2bcd.bin_in[7] ),
    .A2(_0037_));
 sg13g2_nand2_1 _1458_ (.Y(_0686_),
    .A(_0684_),
    .B(_0685_));
 sg13g2_a21oi_2 _1459_ (.B1(_0682_),
    .Y(_0687_),
    .A2(_0685_),
    .A1(_0684_));
 sg13g2_a21o_1 _1460_ (.A2(_0685_),
    .A1(_0684_),
    .B1(_0682_),
    .X(_0688_));
 sg13g2_nor2_1 _1461_ (.A(_0681_),
    .B(_0687_),
    .Y(_0689_));
 sg13g2_nand2_1 _1462_ (.Y(_0690_),
    .A(_0680_),
    .B(_0688_));
 sg13g2_xnor2_1 _1463_ (.Y(_0691_),
    .A(_0039_),
    .B(_0683_));
 sg13g2_o21ai_1 _1464_ (.B1(_0691_),
    .Y(_0692_),
    .A1(_0681_),
    .A2(_0687_));
 sg13g2_nand3_1 _1465_ (.B(_0680_),
    .C(_0688_),
    .A(_0676_),
    .Y(_0693_));
 sg13g2_and2_1 _1466_ (.A(_0692_),
    .B(_0693_),
    .X(_0694_));
 sg13g2_nor2_1 _1467_ (.A(_0681_),
    .B(_0683_),
    .Y(_0695_));
 sg13g2_nand2_1 _1468_ (.Y(_0696_),
    .A(_0680_),
    .B(_0682_));
 sg13g2_and3_1 _1469_ (.X(_0697_),
    .A(_0680_),
    .B(_0682_),
    .C(_0686_));
 sg13g2_nand2_1 _1470_ (.Y(_0698_),
    .A(_0039_),
    .B(_0676_));
 sg13g2_xor2_1 _1471_ (.B(_0698_),
    .A(_0678_),
    .X(_0699_));
 sg13g2_a22oi_1 _1472_ (.Y(_0700_),
    .B1(_0699_),
    .B2(_0690_),
    .A2(_0695_),
    .A1(_0686_));
 sg13g2_a21o_1 _1473_ (.A2(_0699_),
    .A1(_0690_),
    .B1(_0697_),
    .X(_0701_));
 sg13g2_o21ai_1 _1474_ (.B1(\inst_calculator.inst_bin2bcd.bin_in[6] ),
    .Y(_0702_),
    .A1(_0681_),
    .A2(_0687_));
 sg13g2_nand3b_1 _1475_ (.B(_0680_),
    .C(_0688_),
    .Y(_0703_),
    .A_N(\inst_calculator.inst_bin2bcd.bin_in[6] ));
 sg13g2_and2_1 _1476_ (.A(_0702_),
    .B(_0703_),
    .X(_0704_));
 sg13g2_nand2_1 _1477_ (.Y(_0705_),
    .A(_0702_),
    .B(_0703_));
 sg13g2_nand4_1 _1478_ (.B(_0693_),
    .C(_0702_),
    .A(_0692_),
    .Y(_0706_),
    .D(_0703_));
 sg13g2_and2_1 _1479_ (.A(_0692_),
    .B(_0696_),
    .X(_0707_));
 sg13g2_nand3b_1 _1480_ (.B(_0680_),
    .C(_0688_),
    .Y(_0708_),
    .A_N(_0039_));
 sg13g2_o21ai_1 _1481_ (.B1(_0039_),
    .Y(_0709_),
    .A1(_0681_),
    .A2(_0687_));
 sg13g2_nand2_1 _1482_ (.Y(_0710_),
    .A(_0708_),
    .B(_0709_));
 sg13g2_and3_1 _1483_ (.X(_0711_),
    .A(_0592_),
    .B(_0708_),
    .C(_0709_));
 sg13g2_nand4_1 _1484_ (.B(_0696_),
    .C(_0708_),
    .A(_0692_),
    .Y(_0712_),
    .D(_0709_));
 sg13g2_a221oi_1 _1485_ (.B2(_0711_),
    .C1(_0701_),
    .B1(_0707_),
    .A1(_0694_),
    .Y(_0713_),
    .A2(_0704_));
 sg13g2_nand3_1 _1486_ (.B(_0708_),
    .C(_0709_),
    .A(_0040_),
    .Y(_0714_));
 sg13g2_xor2_1 _1487_ (.B(_0714_),
    .A(_0707_),
    .X(_0715_));
 sg13g2_mux2_2 _1488_ (.A0(_0715_),
    .A1(_0694_),
    .S(_0713_),
    .X(_0716_));
 sg13g2_xnor2_1 _1489_ (.Y(_0717_),
    .A(_0040_),
    .B(_0704_));
 sg13g2_nand3_1 _1490_ (.B(_0706_),
    .C(_0710_),
    .A(_0700_),
    .Y(_0718_));
 sg13g2_o21ai_1 _1491_ (.B1(_0718_),
    .Y(_0719_),
    .A1(_0713_),
    .A2(_0717_));
 sg13g2_xnor2_1 _1492_ (.Y(_0720_),
    .A(\inst_calculator.inst_bin2bcd.bin_in[5] ),
    .B(_0713_));
 sg13g2_a21oi_2 _1493_ (.B1(_0716_),
    .Y(_0721_),
    .A2(_0720_),
    .A1(_0719_));
 sg13g2_a21o_1 _1494_ (.A2(_0720_),
    .A1(_0719_),
    .B1(_0716_),
    .X(_0722_));
 sg13g2_nand4_1 _1495_ (.B(_0700_),
    .C(_0706_),
    .A(_0592_),
    .Y(_0723_),
    .D(_0712_));
 sg13g2_a21oi_1 _1496_ (.A1(_0700_),
    .A2(_0706_),
    .Y(_0724_),
    .B1(_0592_));
 sg13g2_a21o_1 _1497_ (.A2(_0713_),
    .A1(_0592_),
    .B1(_0724_),
    .X(_0725_));
 sg13g2_mux2_1 _1498_ (.A0(_0717_),
    .A1(_0705_),
    .S(_0713_),
    .X(_0726_));
 sg13g2_nor3_2 _1499_ (.A(_0041_),
    .B(_0725_),
    .C(_0726_),
    .Y(_0727_));
 sg13g2_or3_2 _1500_ (.A(_0041_),
    .B(_0725_),
    .C(_0726_),
    .X(_0728_));
 sg13g2_nor2_1 _1501_ (.A(_0722_),
    .B(_0727_),
    .Y(_0729_));
 sg13g2_xnor2_1 _1502_ (.Y(_0730_),
    .A(_0593_),
    .B(_0720_));
 sg13g2_o21ai_1 _1503_ (.B1(_0730_),
    .Y(_0731_),
    .A1(_0722_),
    .A2(_0727_));
 sg13g2_nand2_1 _1504_ (.Y(_0732_),
    .A(_0721_),
    .B(_0725_));
 sg13g2_nand2_1 _1505_ (.Y(_0733_),
    .A(_0731_),
    .B(_0732_));
 sg13g2_nand3_1 _1506_ (.B(_0721_),
    .C(_0728_),
    .A(\inst_calculator.inst_bin2bcd.bin_in[4] ),
    .Y(_0734_));
 sg13g2_a21o_1 _1507_ (.A2(_0728_),
    .A1(_0721_),
    .B1(\inst_calculator.inst_bin2bcd.bin_in[4] ),
    .X(_0735_));
 sg13g2_nand2_2 _1508_ (.Y(_0736_),
    .A(_0734_),
    .B(_0735_));
 sg13g2_inv_1 _1509_ (.Y(_0737_),
    .A(_0736_));
 sg13g2_a22oi_1 _1510_ (.Y(_0738_),
    .B1(_0734_),
    .B2(_0735_),
    .A2(_0732_),
    .A1(_0731_));
 sg13g2_nand3b_1 _1511_ (.B(_0041_),
    .C(_0723_),
    .Y(_0739_),
    .A_N(_0724_));
 sg13g2_xnor2_1 _1512_ (.Y(_0740_),
    .A(_0726_),
    .B(_0739_));
 sg13g2_nand3b_1 _1513_ (.B(_0721_),
    .C(_0728_),
    .Y(_0741_),
    .A_N(_0719_));
 sg13g2_o21ai_1 _1514_ (.B1(_0741_),
    .Y(_0742_),
    .A1(_0729_),
    .A2(_0740_));
 sg13g2_mux2_1 _1515_ (.A0(_0740_),
    .A1(_0719_),
    .S(_0729_),
    .X(_0743_));
 sg13g2_nand2_1 _1516_ (.Y(_0744_),
    .A(_0041_),
    .B(_0721_));
 sg13g2_o21ai_1 _1517_ (.B1(_0593_),
    .Y(_0745_),
    .A1(_0722_),
    .A2(_0727_));
 sg13g2_and2_1 _1518_ (.A(_0744_),
    .B(_0745_),
    .X(_0746_));
 sg13g2_nand3_1 _1519_ (.B(_0721_),
    .C(_0728_),
    .A(_0720_),
    .Y(_0747_));
 sg13g2_nand2_1 _1520_ (.Y(_0748_),
    .A(_0731_),
    .B(_0747_));
 sg13g2_a221oi_1 _1521_ (.B2(_0731_),
    .C1(_0042_),
    .B1(_0747_),
    .A1(_0744_),
    .Y(_0749_),
    .A2(_0745_));
 sg13g2_or3_2 _1522_ (.A(_0738_),
    .B(_0743_),
    .C(_0749_),
    .X(_0750_));
 sg13g2_a21o_1 _1523_ (.A2(_0745_),
    .A1(_0744_),
    .B1(_0594_),
    .X(_0751_));
 sg13g2_xor2_1 _1524_ (.B(_0751_),
    .A(_0748_),
    .X(_0752_));
 sg13g2_mux2_1 _1525_ (.A0(_0733_),
    .A1(_0752_),
    .S(_0750_),
    .X(_0753_));
 sg13g2_xnor2_1 _1526_ (.Y(_0754_),
    .A(_0042_),
    .B(_0736_));
 sg13g2_xnor2_1 _1527_ (.Y(_0755_),
    .A(_0594_),
    .B(_0736_));
 sg13g2_mux2_1 _1528_ (.A0(_0746_),
    .A1(_0755_),
    .S(_0750_),
    .X(_0756_));
 sg13g2_xor2_1 _1529_ (.B(_0750_),
    .A(\inst_calculator.inst_bin2bcd.bin_in[3] ),
    .X(_0757_));
 sg13g2_a21oi_2 _1530_ (.B1(_0753_),
    .Y(_0758_),
    .A2(_0757_),
    .A1(_0756_));
 sg13g2_a21o_1 _1531_ (.A2(_0757_),
    .A1(_0756_),
    .B1(_0753_),
    .X(_0759_));
 sg13g2_or4_1 _1532_ (.A(_0042_),
    .B(_0738_),
    .C(_0743_),
    .D(_0749_),
    .X(_0760_));
 sg13g2_o21ai_1 _1533_ (.B1(_0042_),
    .Y(_0761_),
    .A1(_0738_),
    .A2(_0743_));
 sg13g2_nand2_1 _1534_ (.Y(_0762_),
    .A(_0760_),
    .B(_0761_));
 sg13g2_mux2_1 _1535_ (.A0(_0737_),
    .A1(_0754_),
    .S(_0750_),
    .X(_0763_));
 sg13g2_nor3_1 _1536_ (.A(_0043_),
    .B(_0762_),
    .C(_0763_),
    .Y(_0764_));
 sg13g2_or3_2 _1537_ (.A(_0043_),
    .B(_0762_),
    .C(_0763_),
    .X(_0765_));
 sg13g2_nand2_1 _1538_ (.Y(_0766_),
    .A(_0758_),
    .B(_0765_));
 sg13g2_xnor2_1 _1539_ (.Y(_0767_),
    .A(_0595_),
    .B(_0757_));
 sg13g2_o21ai_1 _1540_ (.B1(_0767_),
    .Y(_0768_),
    .A1(_0759_),
    .A2(_0764_));
 sg13g2_nand2_1 _1541_ (.Y(_0769_),
    .A(_0758_),
    .B(_0762_));
 sg13g2_nand2_1 _1542_ (.Y(_0770_),
    .A(_0768_),
    .B(_0769_));
 sg13g2_nand3_1 _1543_ (.B(_0758_),
    .C(_0765_),
    .A(\inst_calculator.inst_bin2bcd.bin_in[2] ),
    .Y(_0771_));
 sg13g2_a21o_1 _1544_ (.A2(_0765_),
    .A1(_0758_),
    .B1(\inst_calculator.inst_bin2bcd.bin_in[2] ),
    .X(_0772_));
 sg13g2_nand2_1 _1545_ (.Y(_0773_),
    .A(_0771_),
    .B(_0772_));
 sg13g2_a22oi_1 _1546_ (.Y(_0774_),
    .B1(_0771_),
    .B2(_0772_),
    .A2(_0769_),
    .A1(_0768_));
 sg13g2_nand3_1 _1547_ (.B(_0760_),
    .C(_0761_),
    .A(_0043_),
    .Y(_0775_));
 sg13g2_xnor2_1 _1548_ (.Y(_0776_),
    .A(_0763_),
    .B(_0775_));
 sg13g2_mux2_1 _1549_ (.A0(_0756_),
    .A1(_0776_),
    .S(_0766_),
    .X(_0777_));
 sg13g2_nand2_1 _1550_ (.Y(_0778_),
    .A(_0043_),
    .B(_0758_));
 sg13g2_o21ai_1 _1551_ (.B1(_0595_),
    .Y(_0779_),
    .A1(_0759_),
    .A2(_0764_));
 sg13g2_nand3_1 _1552_ (.B(_0758_),
    .C(_0765_),
    .A(_0757_),
    .Y(_0780_));
 sg13g2_nand2_1 _1553_ (.Y(_0781_),
    .A(_0768_),
    .B(_0780_));
 sg13g2_a21oi_1 _1554_ (.A1(_0778_),
    .A2(_0779_),
    .Y(_0782_),
    .B1(_0044_));
 sg13g2_a221oi_1 _1555_ (.B2(_0782_),
    .C1(_0777_),
    .B1(_0781_),
    .A1(_0770_),
    .Y(_0783_),
    .A2(_0773_));
 sg13g2_a21oi_1 _1556_ (.A1(_0778_),
    .A2(_0779_),
    .Y(_0784_),
    .B1(_0596_));
 sg13g2_a21o_1 _1557_ (.A2(_0769_),
    .A1(_0768_),
    .B1(_0784_),
    .X(_0785_));
 sg13g2_xor2_1 _1558_ (.B(_0785_),
    .A(_0777_),
    .X(_0786_));
 sg13g2_nor3_1 _1559_ (.A(_0608_),
    .B(_0783_),
    .C(_0786_),
    .Y(_0787_));
 sg13g2_and2_1 _1560_ (.A(_0756_),
    .B(_0775_),
    .X(_0788_));
 sg13g2_or2_1 _1561_ (.X(_0789_),
    .B(_0788_),
    .A(_0753_));
 sg13g2_a22oi_1 _1562_ (.Y(_0790_),
    .B1(_0788_),
    .B2(_0753_),
    .A2(_0765_),
    .A1(_0758_));
 sg13g2_and2_1 _1563_ (.A(_0789_),
    .B(_0790_),
    .X(_0791_));
 sg13g2_and2_1 _1564_ (.A(_0719_),
    .B(_0739_),
    .X(_0792_));
 sg13g2_a21oi_1 _1565_ (.A1(_0719_),
    .A2(_0739_),
    .Y(_0793_),
    .B1(_0716_));
 sg13g2_nand2_1 _1566_ (.Y(_0794_),
    .A(_0716_),
    .B(_0792_));
 sg13g2_a21oi_1 _1567_ (.A1(_0721_),
    .A2(_0728_),
    .Y(_0795_),
    .B1(_0793_));
 sg13g2_a221oi_1 _1568_ (.B2(_0716_),
    .C1(_0793_),
    .B1(_0792_),
    .A1(_0721_),
    .Y(_0796_),
    .A2(_0728_));
 sg13g2_nand2_2 _1569_ (.Y(_0797_),
    .A(_0794_),
    .B(_0795_));
 sg13g2_nor3_2 _1570_ (.A(_0037_),
    .B(_0670_),
    .C(_0671_),
    .Y(_0798_));
 sg13g2_nand2_1 _1571_ (.Y(_0799_),
    .A(_0686_),
    .B(_0698_));
 sg13g2_xor2_1 _1572_ (.B(_0799_),
    .A(_0673_),
    .X(_0800_));
 sg13g2_nor2_1 _1573_ (.A(_0689_),
    .B(_0800_),
    .Y(_0801_));
 sg13g2_nor3_1 _1574_ (.A(_0689_),
    .B(_0798_),
    .C(_0800_),
    .Y(_0802_));
 sg13g2_a21o_1 _1575_ (.A2(_0714_),
    .A1(_0694_),
    .B1(_0700_),
    .X(_0803_));
 sg13g2_nand3_1 _1576_ (.B(_0700_),
    .C(_0714_),
    .A(_0694_),
    .Y(_0804_));
 sg13g2_o21ai_1 _1577_ (.B1(_0803_),
    .Y(_0805_),
    .A1(_0713_),
    .A2(_0804_));
 sg13g2_nor2_1 _1578_ (.A(_0801_),
    .B(_0805_),
    .Y(_0806_));
 sg13g2_nor2b_1 _1579_ (.A(_0806_),
    .B_N(_0798_),
    .Y(_0807_));
 sg13g2_a21oi_1 _1580_ (.A1(_0798_),
    .A2(_0801_),
    .Y(_0808_),
    .B1(_0805_));
 sg13g2_a21oi_1 _1581_ (.A1(_0798_),
    .A2(_0805_),
    .Y(_0809_),
    .B1(_0808_));
 sg13g2_a21o_1 _1582_ (.A2(_0805_),
    .A1(_0798_),
    .B1(_0808_),
    .X(_0810_));
 sg13g2_o21ai_1 _1583_ (.B1(_0802_),
    .Y(_0811_),
    .A1(_0796_),
    .A2(_0809_));
 sg13g2_and2_1 _1584_ (.A(_0798_),
    .B(_0806_),
    .X(_0812_));
 sg13g2_inv_1 _1585_ (.Y(_0813_),
    .A(_0812_));
 sg13g2_nand2_2 _1586_ (.Y(_0814_),
    .A(_0811_),
    .B(_0813_));
 sg13g2_a21oi_1 _1587_ (.A1(_0811_),
    .A2(_0813_),
    .Y(_0815_),
    .B1(_0796_));
 sg13g2_xnor2_1 _1588_ (.Y(_0816_),
    .A(_0796_),
    .B(_0814_));
 sg13g2_xnor2_1 _1589_ (.Y(_0817_),
    .A(_0797_),
    .B(_0814_));
 sg13g2_a21oi_1 _1590_ (.A1(_0733_),
    .A2(_0751_),
    .Y(_0818_),
    .B1(_0742_));
 sg13g2_and3_1 _1591_ (.X(_0819_),
    .A(_0733_),
    .B(_0742_),
    .C(_0751_));
 sg13g2_a21oi_1 _1592_ (.A1(_0750_),
    .A2(_0819_),
    .Y(_0820_),
    .B1(_0818_));
 sg13g2_a21o_1 _1593_ (.A2(_0819_),
    .A1(_0750_),
    .B1(_0818_),
    .X(_0821_));
 sg13g2_nand3_1 _1594_ (.B(_0802_),
    .C(_0810_),
    .A(_0797_),
    .Y(_0822_));
 sg13g2_o21ai_1 _1595_ (.B1(_0822_),
    .Y(_0823_),
    .A1(_0797_),
    .A2(_0813_));
 sg13g2_inv_1 _1596_ (.Y(_0824_),
    .A(_0823_));
 sg13g2_nand3_1 _1597_ (.B(_0810_),
    .C(_0812_),
    .A(_0797_),
    .Y(_0825_));
 sg13g2_o21ai_1 _1598_ (.B1(_0825_),
    .Y(_0826_),
    .A1(_0810_),
    .A2(_0815_));
 sg13g2_nand2_1 _1599_ (.Y(_0827_),
    .A(_0816_),
    .B(_0820_));
 sg13g2_o21ai_1 _1600_ (.B1(_0826_),
    .Y(_0828_),
    .A1(_0817_),
    .A2(_0821_));
 sg13g2_and2_1 _1601_ (.A(_0824_),
    .B(_0828_),
    .X(_0829_));
 sg13g2_nor3_1 _1602_ (.A(_0820_),
    .B(_0823_),
    .C(_0826_),
    .Y(_0830_));
 sg13g2_or2_1 _1603_ (.X(_0831_),
    .B(_0830_),
    .A(_0816_));
 sg13g2_a21o_1 _1604_ (.A2(_0790_),
    .A1(_0789_),
    .B1(_0831_),
    .X(_0832_));
 sg13g2_a21oi_1 _1605_ (.A1(_0824_),
    .A2(_0828_),
    .Y(_0833_),
    .B1(_0821_));
 sg13g2_xnor2_1 _1606_ (.Y(_0834_),
    .A(_0816_),
    .B(_0833_));
 sg13g2_a21oi_1 _1607_ (.A1(_0823_),
    .A2(_0827_),
    .Y(_0835_),
    .B1(_0826_));
 sg13g2_a21oi_1 _1608_ (.A1(_0826_),
    .A2(_0827_),
    .Y(_0836_),
    .B1(_0835_));
 sg13g2_a21oi_2 _1609_ (.B1(_0836_),
    .Y(_0837_),
    .A2(_0834_),
    .A1(_0832_));
 sg13g2_nor2b_1 _1610_ (.A(_0837_),
    .B_N(_0066_),
    .Y(_0838_));
 sg13g2_a21oi_1 _1611_ (.A1(net177),
    .A2(_0064_),
    .Y(_0839_),
    .B1(_0838_));
 sg13g2_nand2b_1 _1612_ (.Y(_0185_),
    .B(_0839_),
    .A_N(_0787_));
 sg13g2_xnor2_1 _1613_ (.Y(_0840_),
    .A(_0791_),
    .B(_0837_));
 sg13g2_xnor2_1 _1614_ (.Y(_0841_),
    .A(\inst_calculator.inst_bin2bcd.bin_in[1] ),
    .B(_0783_));
 sg13g2_nand2_1 _1615_ (.Y(_0842_),
    .A(_0064_),
    .B(_0841_));
 sg13g2_nor2_1 _1616_ (.A(_0807_),
    .B(_0829_),
    .Y(_0843_));
 sg13g2_a22oi_1 _1617_ (.Y(_0844_),
    .B1(_0843_),
    .B2(_0066_),
    .A2(_0840_),
    .A1(net311));
 sg13g2_a22oi_1 _1618_ (.Y(_0186_),
    .B1(_0842_),
    .B2(_0844_),
    .A2(net166),
    .A1(\inst_calculator.inst_drive.cnt_sel[1] ));
 sg13g2_nor2_1 _1619_ (.A(_0830_),
    .B(_0833_),
    .Y(_0845_));
 sg13g2_o21ai_1 _1620_ (.B1(_0845_),
    .Y(_0846_),
    .A1(_0791_),
    .A2(_0837_));
 sg13g2_or3_1 _1621_ (.A(_0791_),
    .B(_0837_),
    .C(_0845_),
    .X(_0847_));
 sg13g2_nand3_1 _1622_ (.B(_0846_),
    .C(_0847_),
    .A(net311),
    .Y(_0848_));
 sg13g2_o21ai_1 _1623_ (.B1(net420),
    .Y(_0849_),
    .A1(_0774_),
    .A2(_0777_));
 sg13g2_xnor2_1 _1624_ (.Y(_0850_),
    .A(_0773_),
    .B(_0849_));
 sg13g2_a22oi_1 _1625_ (.Y(_0851_),
    .B1(_0850_),
    .B2(_0064_),
    .A2(_0814_),
    .A1(_0066_));
 sg13g2_a22oi_1 _1626_ (.Y(_0187_),
    .B1(_0848_),
    .B2(_0851_),
    .A2(net311),
    .A1(net405));
 sg13g2_xnor2_1 _1627_ (.Y(_0852_),
    .A(_0770_),
    .B(_0784_));
 sg13g2_nor2_1 _1628_ (.A(_0783_),
    .B(_0852_),
    .Y(_0853_));
 sg13g2_nor3_1 _1629_ (.A(_0774_),
    .B(_0777_),
    .C(_0781_),
    .Y(_0854_));
 sg13g2_nor4_1 _1630_ (.A(net405),
    .B(net311),
    .C(_0853_),
    .D(_0854_),
    .Y(_0855_));
 sg13g2_nand2b_1 _1631_ (.Y(_0856_),
    .B(_0845_),
    .A_N(_0791_));
 sg13g2_a21oi_1 _1632_ (.A1(_0836_),
    .A2(_0856_),
    .Y(_0857_),
    .B1(_0834_));
 sg13g2_a21o_1 _1633_ (.A2(_0834_),
    .A1(_0832_),
    .B1(_0608_),
    .X(_0858_));
 sg13g2_nand3_1 _1634_ (.B(_0807_),
    .C(_0829_),
    .A(_0066_),
    .Y(_0859_));
 sg13g2_o21ai_1 _1635_ (.B1(_0859_),
    .Y(_0860_),
    .A1(_0857_),
    .A2(_0858_));
 sg13g2_or2_1 _1636_ (.X(_0188_),
    .B(_0860_),
    .A(_0855_));
 sg13g2_nor2_1 _1637_ (.A(\inst_calculator.inst_keypad_encoder.rows[2] ),
    .B(\inst_calculator.inst_keypad_encoder.rows[3] ),
    .Y(_0861_));
 sg13g2_nand3b_1 _1638_ (.B(_0861_),
    .C(\inst_calculator.inst_keypad_encoder.rows[1] ),
    .Y(_0862_),
    .A_N(\inst_calculator.inst_keypad_encoder.rows[0] ));
 sg13g2_nor2_1 _1639_ (.A(\inst_calculator.inst_keypad_encoder.rows[1] ),
    .B(\inst_calculator.inst_keypad_encoder.rows[0] ),
    .Y(_0863_));
 sg13g2_nand3b_1 _1640_ (.B(\inst_calculator.inst_keypad_encoder.rows[3] ),
    .C(_0863_),
    .Y(_0864_),
    .A_N(\inst_calculator.inst_keypad_encoder.rows[2] ));
 sg13g2_nand2_1 _1641_ (.Y(_0865_),
    .A(_0862_),
    .B(_0864_));
 sg13g2_nand3b_1 _1642_ (.B(_0863_),
    .C(net402),
    .Y(_0866_),
    .A_N(\inst_calculator.inst_keypad_encoder.rows[3] ));
 sg13g2_nand2_1 _1643_ (.Y(_0867_),
    .A(_0864_),
    .B(_0866_));
 sg13g2_nor2b_1 _1644_ (.A(_0867_),
    .B_N(_0862_),
    .Y(_0868_));
 sg13g2_nand3b_1 _1645_ (.B(net195),
    .C(_0861_),
    .Y(_0869_),
    .A_N(\inst_calculator.inst_keypad_encoder.rows[1] ));
 sg13g2_and2_1 _1646_ (.A(_0868_),
    .B(_0869_),
    .X(_0870_));
 sg13g2_nor2_1 _1647_ (.A(uio_out[7]),
    .B(uio_out[6]),
    .Y(_0871_));
 sg13g2_nand3b_1 _1648_ (.B(net451),
    .C(_0871_),
    .Y(_0872_),
    .A_N(uio_out[5]));
 sg13g2_nor2_1 _1649_ (.A(_0865_),
    .B(_0872_),
    .Y(_0873_));
 sg13g2_nor2_1 _1650_ (.A(uio_out[5]),
    .B(net433),
    .Y(_0874_));
 sg13g2_nand3_1 _1651_ (.B(uio_out[6]),
    .C(_0874_),
    .A(_0561_),
    .Y(_0875_));
 sg13g2_nor2_1 _1652_ (.A(net379),
    .B(_0875_),
    .Y(_0876_));
 sg13g2_nor2_1 _1653_ (.A(_0873_),
    .B(_0876_),
    .Y(_0877_));
 sg13g2_nand3b_1 _1654_ (.B(_0874_),
    .C(net444),
    .Y(_0878_),
    .A_N(uio_out[6]));
 sg13g2_nand3b_1 _1655_ (.B(_0871_),
    .C(uio_out[5]),
    .Y(_0879_),
    .A_N(uio_out[4]));
 sg13g2_o21ai_1 _1656_ (.B1(_0878_),
    .Y(_0880_),
    .A1(_0862_),
    .A2(_0879_));
 sg13g2_nand2_1 _1657_ (.Y(_0881_),
    .A(_0865_),
    .B(net446));
 sg13g2_o21ai_1 _1658_ (.B1(net447),
    .Y(_0189_),
    .A1(_0870_),
    .A2(_0877_));
 sg13g2_nor3_1 _1659_ (.A(net402),
    .B(_0870_),
    .C(_0875_),
    .Y(_0882_));
 sg13g2_a21oi_1 _1660_ (.A1(_0862_),
    .A2(_0869_),
    .Y(_0883_),
    .B1(_0878_));
 sg13g2_nand2b_1 _1661_ (.Y(_0884_),
    .B(_0867_),
    .A_N(_0872_));
 sg13g2_o21ai_1 _1662_ (.B1(_0884_),
    .Y(_0885_),
    .A1(_0869_),
    .A2(_0879_));
 sg13g2_or3_1 _1663_ (.A(_0882_),
    .B(_0883_),
    .C(_0885_),
    .X(_0190_));
 sg13g2_nand2b_1 _1664_ (.Y(_0886_),
    .B(_0867_),
    .A_N(_0878_));
 sg13g2_o21ai_1 _1665_ (.B1(_0886_),
    .Y(_0887_),
    .A1(_0868_),
    .A2(_0872_));
 sg13g2_o21ai_1 _1666_ (.B1(_0875_),
    .Y(_0888_),
    .A1(_0862_),
    .A2(_0879_));
 sg13g2_a21o_1 _1667_ (.A2(_0888_),
    .A1(_0865_),
    .B1(_0887_),
    .X(_0191_));
 sg13g2_nor2_1 _1668_ (.A(_0866_),
    .B(_0879_),
    .Y(_0889_));
 sg13g2_o21ai_1 _1669_ (.B1(_0875_),
    .Y(_0890_),
    .A1(_0864_),
    .A2(_0872_));
 sg13g2_a21oi_1 _1670_ (.A1(_0867_),
    .A2(_0890_),
    .Y(_0891_),
    .B1(_0889_));
 sg13g2_o21ai_1 _1671_ (.B1(_0891_),
    .Y(_0192_),
    .A1(_0870_),
    .A2(net445));
 sg13g2_nor4_1 _1672_ (.A(_0563_),
    .B(net312),
    .C(_0601_),
    .D(net365),
    .Y(_0010_));
 sg13g2_and3_1 _1673_ (.X(_0006_),
    .A(net156),
    .B(_0624_),
    .C(_0628_));
 sg13g2_nand3b_1 _1674_ (.B(_0600_),
    .C(net364),
    .Y(_0892_),
    .A_N(net381));
 sg13g2_nor3_1 _1675_ (.A(\inst_calculator.inst_keypad_encoder.key[0] ),
    .B(_0565_),
    .C(_0892_),
    .Y(_0012_));
 sg13g2_nor4_1 _1676_ (.A(net190),
    .B(net312),
    .C(_0601_),
    .D(_0602_),
    .Y(_0011_));
 sg13g2_nor2b_1 _1677_ (.A(_0599_),
    .B_N(net358),
    .Y(_0009_));
 sg13g2_a21oi_1 _1678_ (.A1(_0563_),
    .A2(net312),
    .Y(_0008_),
    .B1(_0892_));
 sg13g2_and3_1 _1679_ (.X(_0007_),
    .A(net160),
    .B(_0619_),
    .C(_0624_));
 sg13g2_nor3_1 _1680_ (.A(net321),
    .B(net324),
    .C(net326),
    .Y(_0893_));
 sg13g2_nand2_1 _1681_ (.Y(_0894_),
    .A(net316),
    .B(net319));
 sg13g2_nor3_1 _1682_ (.A(\inst_calculator.reg_arg[9] ),
    .B(net313),
    .C(\inst_calculator.reg_arg[7] ),
    .Y(_0895_));
 sg13g2_o21ai_1 _1683_ (.B1(_0895_),
    .Y(_0896_),
    .A1(_0893_),
    .A2(_0894_));
 sg13g2_nor3_1 _1684_ (.A(net298),
    .B(\inst_calculator.state[0] ),
    .C(net89),
    .Y(_0897_));
 sg13g2_a21oi_1 _1685_ (.A1(net89),
    .A2(_0896_),
    .Y(_0898_),
    .B1(_0897_));
 sg13g2_nand2_2 _1686_ (.Y(_0899_),
    .A(net339),
    .B(_0898_));
 sg13g2_nor3_2 _1687_ (.A(net298),
    .B(net206),
    .C(_0899_),
    .Y(_0900_));
 sg13g2_a22oi_1 _1688_ (.Y(_0901_),
    .B1(_0900_),
    .B2(net190),
    .A2(net271),
    .A1(net332));
 sg13g2_inv_1 _1689_ (.Y(_0069_),
    .A(net207));
 sg13g2_xor2_1 _1690_ (.B(net332),
    .A(net312),
    .X(_0902_));
 sg13g2_a22oi_1 _1691_ (.Y(_0903_),
    .B1(_0900_),
    .B2(_0902_),
    .A2(net271),
    .A1(net330));
 sg13g2_inv_1 _1692_ (.Y(_0070_),
    .A(_0903_));
 sg13g2_nand2_1 _1693_ (.Y(_0904_),
    .A(net326),
    .B(net271));
 sg13g2_nand2_1 _1694_ (.Y(_0905_),
    .A(\inst_calculator.inst_keypad_encoder.key[2] ),
    .B(net330));
 sg13g2_xor2_1 _1695_ (.B(net330),
    .A(net408),
    .X(_0906_));
 sg13g2_a21oi_1 _1696_ (.A1(net312),
    .A2(net332),
    .Y(_0907_),
    .B1(_0906_));
 sg13g2_nand3_1 _1697_ (.B(net332),
    .C(_0906_),
    .A(net312),
    .Y(_0908_));
 sg13g2_nand2_1 _1698_ (.Y(_0909_),
    .A(net268),
    .B(_0908_));
 sg13g2_o21ai_1 _1699_ (.B1(_0904_),
    .Y(_0071_),
    .A1(_0907_),
    .A2(_0909_));
 sg13g2_nand2_1 _1700_ (.Y(_0910_),
    .A(net325),
    .B(net331));
 sg13g2_xor2_1 _1701_ (.B(net331),
    .A(net326),
    .X(_0911_));
 sg13g2_xnor2_1 _1702_ (.Y(_0912_),
    .A(\inst_calculator.inst_keypad_encoder.key[3] ),
    .B(_0911_));
 sg13g2_a21oi_1 _1703_ (.A1(_0905_),
    .A2(_0908_),
    .Y(_0913_),
    .B1(_0912_));
 sg13g2_nand3_1 _1704_ (.B(_0908_),
    .C(_0912_),
    .A(_0905_),
    .Y(_0914_));
 sg13g2_nor2b_1 _1705_ (.A(_0913_),
    .B_N(_0914_),
    .Y(_0915_));
 sg13g2_a22oi_1 _1706_ (.Y(_0916_),
    .B1(net268),
    .B2(_0915_),
    .A2(_0899_),
    .A1(net323));
 sg13g2_inv_1 _1707_ (.Y(_0072_),
    .A(_0916_));
 sg13g2_xnor2_1 _1708_ (.Y(_0917_),
    .A(net323),
    .B(net329));
 sg13g2_nor2_1 _1709_ (.A(_0910_),
    .B(_0917_),
    .Y(_0918_));
 sg13g2_inv_1 _1710_ (.Y(_0919_),
    .A(_0918_));
 sg13g2_xnor2_1 _1711_ (.Y(_0920_),
    .A(_0910_),
    .B(_0917_));
 sg13g2_a21oi_1 _1712_ (.A1(_0566_),
    .A2(_0911_),
    .Y(_0921_),
    .B1(_0913_));
 sg13g2_nor2_1 _1713_ (.A(_0920_),
    .B(_0921_),
    .Y(_0922_));
 sg13g2_nand2b_1 _1714_ (.Y(_0923_),
    .B(net268),
    .A_N(_0922_));
 sg13g2_a21oi_1 _1715_ (.A1(_0920_),
    .A2(_0921_),
    .Y(_0924_),
    .B1(_0923_));
 sg13g2_a21o_1 _1716_ (.A2(net271),
    .A1(net321),
    .B1(_0924_),
    .X(_0073_));
 sg13g2_nand2_1 _1717_ (.Y(_0925_),
    .A(net321),
    .B(net326));
 sg13g2_xor2_1 _1718_ (.B(net326),
    .A(net321),
    .X(_0926_));
 sg13g2_nand3_1 _1719_ (.B(net329),
    .C(_0926_),
    .A(net323),
    .Y(_0927_));
 sg13g2_a21o_1 _1720_ (.A2(net329),
    .A1(net323),
    .B1(_0926_),
    .X(_0928_));
 sg13g2_a21oi_1 _1721_ (.A1(_0927_),
    .A2(_0928_),
    .Y(_0929_),
    .B1(_0918_));
 sg13g2_a21oi_1 _1722_ (.A1(_0571_),
    .A2(_0918_),
    .Y(_0930_),
    .B1(_0929_));
 sg13g2_nand2_1 _1723_ (.Y(_0931_),
    .A(_0922_),
    .B(_0930_));
 sg13g2_o21ai_1 _1724_ (.B1(net268),
    .Y(_0932_),
    .A1(_0922_),
    .A2(_0930_));
 sg13g2_nor2b_1 _1725_ (.A(_0932_),
    .B_N(_0931_),
    .Y(_0933_));
 sg13g2_a21o_1 _1726_ (.A2(net271),
    .A1(net317),
    .B1(_0933_),
    .X(_0074_));
 sg13g2_o21ai_1 _1727_ (.B1(_0927_),
    .Y(_0934_),
    .A1(net320),
    .A2(_0919_));
 sg13g2_xor2_1 _1728_ (.B(net323),
    .A(net317),
    .X(_0935_));
 sg13g2_nand2b_1 _1729_ (.Y(_0936_),
    .B(_0935_),
    .A_N(_0925_));
 sg13g2_xnor2_1 _1730_ (.Y(_0937_),
    .A(_0925_),
    .B(_0935_));
 sg13g2_xnor2_1 _1731_ (.Y(_0938_),
    .A(_0934_),
    .B(_0937_));
 sg13g2_nor2_1 _1732_ (.A(_0931_),
    .B(_0938_),
    .Y(_0939_));
 sg13g2_o21ai_1 _1733_ (.B1(net268),
    .Y(_0940_),
    .A1(_0931_),
    .A2(_0938_));
 sg13g2_a21oi_1 _1734_ (.A1(_0931_),
    .A2(_0938_),
    .Y(_0941_),
    .B1(_0940_));
 sg13g2_a21o_1 _1735_ (.A2(net271),
    .A1(net315),
    .B1(_0941_),
    .X(_0075_));
 sg13g2_nand2_2 _1736_ (.Y(_0942_),
    .A(net315),
    .B(net321));
 sg13g2_nand2_1 _1737_ (.Y(_0943_),
    .A(_0569_),
    .B(_0571_));
 sg13g2_a22oi_1 _1738_ (.Y(_0944_),
    .B1(_0942_),
    .B2(_0943_),
    .A2(net323),
    .A1(net318));
 sg13g2_nand4_1 _1739_ (.B(net323),
    .C(_0942_),
    .A(net317),
    .Y(_0945_),
    .D(_0943_));
 sg13g2_nor2b_1 _1740_ (.A(_0944_),
    .B_N(_0945_),
    .Y(_0946_));
 sg13g2_nand3_1 _1741_ (.B(_0926_),
    .C(_0935_),
    .A(_0918_),
    .Y(_0947_));
 sg13g2_o21ai_1 _1742_ (.B1(_0936_),
    .Y(_0948_),
    .A1(net317),
    .A2(_0927_));
 sg13g2_nor2b_1 _1743_ (.A(_0948_),
    .B_N(_0947_),
    .Y(_0949_));
 sg13g2_xnor2_1 _1744_ (.Y(_0950_),
    .A(_0946_),
    .B(_0949_));
 sg13g2_nand2_1 _1745_ (.Y(_0951_),
    .A(_0939_),
    .B(_0950_));
 sg13g2_o21ai_1 _1746_ (.B1(net268),
    .Y(_0952_),
    .A1(_0939_),
    .A2(_0950_));
 sg13g2_nor2b_1 _1747_ (.A(_0952_),
    .B_N(_0951_),
    .Y(_0953_));
 sg13g2_a21o_1 _1748_ (.A2(net271),
    .A1(net314),
    .B1(_0953_),
    .X(_0076_));
 sg13g2_o21ai_1 _1749_ (.B1(_0945_),
    .Y(_0954_),
    .A1(_0944_),
    .A2(_0949_));
 sg13g2_nand2_1 _1750_ (.Y(_0955_),
    .A(net314),
    .B(net317));
 sg13g2_xnor2_1 _1751_ (.Y(_0956_),
    .A(net314),
    .B(net317));
 sg13g2_xor2_1 _1752_ (.B(_0956_),
    .A(_0942_),
    .X(_0957_));
 sg13g2_nand2_1 _1753_ (.Y(_0958_),
    .A(_0954_),
    .B(_0957_));
 sg13g2_xnor2_1 _1754_ (.Y(_0959_),
    .A(_0954_),
    .B(_0957_));
 sg13g2_nor2_1 _1755_ (.A(_0951_),
    .B(_0959_),
    .Y(_0960_));
 sg13g2_xor2_1 _1756_ (.B(_0959_),
    .A(_0951_),
    .X(_0961_));
 sg13g2_a22oi_1 _1757_ (.Y(_0962_),
    .B1(net268),
    .B2(_0961_),
    .A2(net271),
    .A1(net313));
 sg13g2_inv_1 _1758_ (.Y(_0077_),
    .A(_0962_));
 sg13g2_nand2_1 _1759_ (.Y(_0963_),
    .A(net423),
    .B(_0899_));
 sg13g2_xnor2_1 _1760_ (.Y(_0964_),
    .A(net313),
    .B(net315));
 sg13g2_xnor2_1 _1761_ (.Y(_0965_),
    .A(_0955_),
    .B(_0964_));
 sg13g2_o21ai_1 _1762_ (.B1(_0958_),
    .Y(_0966_),
    .A1(_0942_),
    .A2(_0956_));
 sg13g2_xnor2_1 _1763_ (.Y(_0967_),
    .A(_0960_),
    .B(_0965_));
 sg13g2_o21ai_1 _1764_ (.B1(net268),
    .Y(_0968_),
    .A1(_0966_),
    .A2(_0967_));
 sg13g2_nand2_1 _1765_ (.Y(_0078_),
    .A(_0963_),
    .B(_0968_));
 sg13g2_nor2_1 _1766_ (.A(net160),
    .B(net156),
    .Y(_0969_));
 sg13g2_or2_1 _1767_ (.X(_0970_),
    .B(\inst_calculator.inst_keypad_poller.state[1] ),
    .A(\inst_calculator.inst_keypad_poller.state[2] ));
 sg13g2_o21ai_1 _1768_ (.B1(_0609_),
    .Y(_0971_),
    .A1(\inst_calculator.inst_keypad_poller.state[5] ),
    .A2(\inst_calculator.inst_keypad_poller.state[4] ));
 sg13g2_or4_1 _1769_ (.A(\inst_calculator.inst_keypad_poller.state[5] ),
    .B(\inst_calculator.inst_keypad_poller.state[3] ),
    .C(\inst_calculator.inst_keypad_poller.state[4] ),
    .D(_0970_),
    .X(_0972_));
 sg13g2_nand3_1 _1770_ (.B(_0971_),
    .C(_0972_),
    .A(net353),
    .Y(_0973_));
 sg13g2_inv_1 _1771_ (.Y(_0974_),
    .A(_0973_));
 sg13g2_nor2_1 _1772_ (.A(_0969_),
    .B(_0973_),
    .Y(_0975_));
 sg13g2_a22oi_1 _1773_ (.Y(_0976_),
    .B1(_0975_),
    .B2(net94),
    .A2(_0973_),
    .A1(\inst_calculator.inst_keypad_poller.clk_counter[0] ));
 sg13g2_inv_1 _1774_ (.Y(_0079_),
    .A(net95));
 sg13g2_and2_1 _1775_ (.A(\inst_calculator.inst_keypad_poller.clk_counter[0] ),
    .B(net200),
    .X(_0977_));
 sg13g2_nor4_1 _1776_ (.A(_0621_),
    .B(_0969_),
    .C(_0973_),
    .D(_0977_),
    .Y(_0978_));
 sg13g2_a21o_1 _1777_ (.A2(_0973_),
    .A1(net200),
    .B1(_0978_),
    .X(_0080_));
 sg13g2_a21oi_1 _1778_ (.A1(_0974_),
    .A2(_0977_),
    .Y(_0979_),
    .B1(net163));
 sg13g2_nor2_1 _1779_ (.A(_0970_),
    .B(_0973_),
    .Y(_0980_));
 sg13g2_nand2_1 _1780_ (.Y(_0981_),
    .A(net163),
    .B(_0977_));
 sg13g2_nor2_1 _1781_ (.A(_0973_),
    .B(_0981_),
    .Y(_0982_));
 sg13g2_nor3_1 _1782_ (.A(net164),
    .B(net270),
    .C(_0982_),
    .Y(_0081_));
 sg13g2_nor2_1 _1783_ (.A(net247),
    .B(_0982_),
    .Y(_0983_));
 sg13g2_and2_1 _1784_ (.A(net247),
    .B(_0982_),
    .X(_0984_));
 sg13g2_nor3_1 _1785_ (.A(net270),
    .B(net248),
    .C(_0984_),
    .Y(_0082_));
 sg13g2_nor2_1 _1786_ (.A(net239),
    .B(_0984_),
    .Y(_0985_));
 sg13g2_and2_1 _1787_ (.A(net239),
    .B(_0984_),
    .X(_0986_));
 sg13g2_nor3_1 _1788_ (.A(net270),
    .B(net240),
    .C(_0986_),
    .Y(_0083_));
 sg13g2_nor2_1 _1789_ (.A(net243),
    .B(_0986_),
    .Y(_0987_));
 sg13g2_and2_1 _1790_ (.A(net243),
    .B(_0986_),
    .X(_0988_));
 sg13g2_nor3_1 _1791_ (.A(net270),
    .B(_0987_),
    .C(_0988_),
    .Y(_0084_));
 sg13g2_nor2_1 _1792_ (.A(net211),
    .B(_0988_),
    .Y(_0989_));
 sg13g2_and2_1 _1793_ (.A(net211),
    .B(_0988_),
    .X(_0990_));
 sg13g2_nor3_1 _1794_ (.A(net270),
    .B(net212),
    .C(_0990_),
    .Y(_0085_));
 sg13g2_nor2_1 _1795_ (.A(net407),
    .B(_0990_),
    .Y(_0991_));
 sg13g2_and2_1 _1796_ (.A(net407),
    .B(_0990_),
    .X(_0992_));
 sg13g2_nor3_1 _1797_ (.A(net269),
    .B(_0991_),
    .C(_0992_),
    .Y(_0086_));
 sg13g2_nor2_1 _1798_ (.A(net232),
    .B(_0992_),
    .Y(_0993_));
 sg13g2_and2_1 _1799_ (.A(net232),
    .B(_0992_),
    .X(_0994_));
 sg13g2_nor3_1 _1800_ (.A(net269),
    .B(net233),
    .C(_0994_),
    .Y(_0087_));
 sg13g2_nor2_1 _1801_ (.A(net382),
    .B(_0994_),
    .Y(_0995_));
 sg13g2_and2_1 _1802_ (.A(net382),
    .B(_0994_),
    .X(_0996_));
 sg13g2_nor3_1 _1803_ (.A(net270),
    .B(_0995_),
    .C(_0996_),
    .Y(_0088_));
 sg13g2_nor2_1 _1804_ (.A(net369),
    .B(_0996_),
    .Y(_0997_));
 sg13g2_and2_1 _1805_ (.A(net369),
    .B(_0996_),
    .X(_0998_));
 sg13g2_nor3_1 _1806_ (.A(net269),
    .B(net370),
    .C(_0998_),
    .Y(_0089_));
 sg13g2_nor2_1 _1807_ (.A(net398),
    .B(_0998_),
    .Y(_0999_));
 sg13g2_and2_1 _1808_ (.A(net398),
    .B(_0998_),
    .X(_1000_));
 sg13g2_nor3_1 _1809_ (.A(net269),
    .B(_0999_),
    .C(_1000_),
    .Y(_0090_));
 sg13g2_nor2_1 _1810_ (.A(net395),
    .B(_1000_),
    .Y(_1001_));
 sg13g2_and2_1 _1811_ (.A(net395),
    .B(_1000_),
    .X(_1002_));
 sg13g2_nor3_1 _1812_ (.A(net270),
    .B(net396),
    .C(_1002_),
    .Y(_0091_));
 sg13g2_nor2_1 _1813_ (.A(net392),
    .B(_1002_),
    .Y(_1003_));
 sg13g2_and2_1 _1814_ (.A(net392),
    .B(_1002_),
    .X(_1004_));
 sg13g2_nor3_1 _1815_ (.A(net269),
    .B(net393),
    .C(_1004_),
    .Y(_0092_));
 sg13g2_nor2_1 _1816_ (.A(net388),
    .B(_1004_),
    .Y(_1005_));
 sg13g2_and2_1 _1817_ (.A(net388),
    .B(_1004_),
    .X(_1006_));
 sg13g2_nor3_1 _1818_ (.A(net269),
    .B(net389),
    .C(_1006_),
    .Y(_0093_));
 sg13g2_nor2_1 _1819_ (.A(net397),
    .B(_1006_),
    .Y(_1007_));
 sg13g2_and2_1 _1820_ (.A(net397),
    .B(_1006_),
    .X(_1008_));
 sg13g2_nor3_1 _1821_ (.A(net269),
    .B(_1007_),
    .C(_1008_),
    .Y(_0094_));
 sg13g2_a21oi_1 _1822_ (.A1(net412),
    .A2(_1008_),
    .Y(_1009_),
    .B1(net269));
 sg13g2_o21ai_1 _1823_ (.B1(_1009_),
    .Y(_1010_),
    .A1(net412),
    .A2(_1008_));
 sg13g2_inv_1 _1824_ (.Y(_0095_),
    .A(_1010_));
 sg13g2_nor2b_1 _1825_ (.A(net218),
    .B_N(net225),
    .Y(_1011_));
 sg13g2_nand2b_1 _1826_ (.Y(_1012_),
    .B(\inst_calculator.inst_divider.n[8] ),
    .A_N(\inst_calculator.inst_divider.d[8] ));
 sg13g2_nor2b_1 _1827_ (.A(\inst_calculator.inst_divider.n[8] ),
    .B_N(\inst_calculator.inst_divider.d[8] ),
    .Y(_1013_));
 sg13g2_xnor2_1 _1828_ (.Y(_1014_),
    .A(net165),
    .B(\inst_calculator.inst_divider.n[7] ));
 sg13g2_xor2_1 _1829_ (.B(net261),
    .A(net162),
    .X(_1015_));
 sg13g2_nor2b_1 _1830_ (.A(net208),
    .B_N(\inst_calculator.inst_divider.n[5] ),
    .Y(_1016_));
 sg13g2_xnor2_1 _1831_ (.Y(_1017_),
    .A(net208),
    .B(net244));
 sg13g2_nand2b_1 _1832_ (.Y(_1018_),
    .B(net450),
    .A_N(\inst_calculator.inst_divider.d[4] ));
 sg13g2_xor2_1 _1833_ (.B(net249),
    .A(\inst_calculator.inst_divider.d[4] ),
    .X(_1019_));
 sg13g2_nor2b_1 _1834_ (.A(net204),
    .B_N(\inst_calculator.inst_divider.n[3] ),
    .Y(_1020_));
 sg13g2_xnor2_1 _1835_ (.Y(_1021_),
    .A(\inst_calculator.inst_divider.d[3] ),
    .B(net257));
 sg13g2_nand2b_1 _1836_ (.Y(_1022_),
    .B(\inst_calculator.inst_divider.n[2] ),
    .A_N(\inst_calculator.inst_divider.d[2] ));
 sg13g2_xor2_1 _1837_ (.B(net377),
    .A(\inst_calculator.inst_divider.d[2] ),
    .X(_1023_));
 sg13g2_nor2b_1 _1838_ (.A(\inst_calculator.inst_divider.d[1] ),
    .B_N(\inst_calculator.inst_divider.n[1] ),
    .Y(_1024_));
 sg13g2_xnor2_1 _1839_ (.Y(_1025_),
    .A(\inst_calculator.inst_divider.d[1] ),
    .B(net214));
 sg13g2_nor2b_1 _1840_ (.A(net142),
    .B_N(\inst_calculator.inst_divider.d[0] ),
    .Y(_1026_));
 sg13g2_nand2b_1 _1841_ (.Y(_1027_),
    .B(\inst_calculator.inst_divider.d[0] ),
    .A_N(net142));
 sg13g2_a21oi_1 _1842_ (.A1(_1025_),
    .A2(_1027_),
    .Y(_1028_),
    .B1(_1024_));
 sg13g2_o21ai_1 _1843_ (.B1(_1022_),
    .Y(_1029_),
    .A1(_1023_),
    .A2(_1028_));
 sg13g2_a21oi_1 _1844_ (.A1(_1021_),
    .A2(_1029_),
    .Y(_1030_),
    .B1(_1020_));
 sg13g2_o21ai_1 _1845_ (.B1(_1018_),
    .Y(_1031_),
    .A1(_1019_),
    .A2(_1030_));
 sg13g2_a21oi_1 _1846_ (.A1(_1017_),
    .A2(_1031_),
    .Y(_1032_),
    .B1(_1016_));
 sg13g2_nor2_1 _1847_ (.A(_1015_),
    .B(_1032_),
    .Y(_1033_));
 sg13g2_a21oi_1 _1848_ (.A1(_0577_),
    .A2(net261),
    .Y(_1034_),
    .B1(_1033_));
 sg13g2_nor2b_1 _1849_ (.A(_1034_),
    .B_N(_1014_),
    .Y(_1035_));
 sg13g2_a21oi_1 _1850_ (.A1(_0576_),
    .A2(net373),
    .Y(_1036_),
    .B1(_1035_));
 sg13g2_o21ai_1 _1851_ (.B1(_1012_),
    .Y(_1037_),
    .A1(_1013_),
    .A2(_1036_));
 sg13g2_nand2b_1 _1852_ (.Y(_1038_),
    .B(\inst_calculator.inst_divider.d[9] ),
    .A_N(\inst_calculator.inst_divider.n[9] ));
 sg13g2_a21oi_1 _1853_ (.A1(_1037_),
    .A2(_1038_),
    .Y(_1039_),
    .B1(_1011_));
 sg13g2_nor3_2 _1854_ (.A(net309),
    .B(_0578_),
    .C(_1039_),
    .Y(_1040_));
 sg13g2_inv_2 _1855_ (.Y(_1041_),
    .A(_1040_));
 sg13g2_mux2_1 _1856_ (.A0(\inst_calculator.inst_divider.q[0] ),
    .A1(net100),
    .S(_1040_),
    .X(_0096_));
 sg13g2_nand3_1 _1857_ (.B(net436),
    .C(_1040_),
    .A(net430),
    .Y(_1042_));
 sg13g2_a21o_1 _1858_ (.A2(_1040_),
    .A1(net436),
    .B1(net430),
    .X(_1043_));
 sg13g2_and2_1 _1859_ (.A(_1042_),
    .B(_1043_),
    .X(_0097_));
 sg13g2_nand4_1 _1860_ (.B(\inst_calculator.inst_divider.q[1] ),
    .C(\inst_calculator.inst_divider.q[0] ),
    .A(\inst_calculator.inst_divider.q[2] ),
    .Y(_1044_),
    .D(_1040_));
 sg13g2_xnor2_1 _1861_ (.Y(_0098_),
    .A(net209),
    .B(_1042_));
 sg13g2_nor2_1 _1862_ (.A(_0584_),
    .B(_1044_),
    .Y(_1045_));
 sg13g2_xnor2_1 _1863_ (.Y(_0099_),
    .A(net184),
    .B(_1044_));
 sg13g2_and2_1 _1864_ (.A(net158),
    .B(_1045_),
    .X(_1046_));
 sg13g2_xor2_1 _1865_ (.B(_1045_),
    .A(net158),
    .X(_0100_));
 sg13g2_xor2_1 _1866_ (.B(_1046_),
    .A(net182),
    .X(_0101_));
 sg13g2_and3_1 _1867_ (.X(_1047_),
    .A(net153),
    .B(net182),
    .C(_1046_));
 sg13g2_a21oi_1 _1868_ (.A1(\inst_calculator.inst_divider.q[5] ),
    .A2(_1046_),
    .Y(_1048_),
    .B1(net153));
 sg13g2_nor2_1 _1869_ (.A(_1047_),
    .B(net154),
    .Y(_0102_));
 sg13g2_xor2_1 _1870_ (.B(_1047_),
    .A(net234),
    .X(_0103_));
 sg13g2_nand3_1 _1871_ (.B(net234),
    .C(_1047_),
    .A(net383),
    .Y(_1049_));
 sg13g2_a21o_1 _1872_ (.A2(_1047_),
    .A1(net234),
    .B1(net383),
    .X(_1050_));
 sg13g2_and2_1 _1873_ (.A(_1049_),
    .B(_1050_),
    .X(_0104_));
 sg13g2_xnor2_1 _1874_ (.Y(_0105_),
    .A(net148),
    .B(_1049_));
 sg13g2_nor2_2 _1875_ (.A(net308),
    .B(_1040_),
    .Y(_1051_));
 sg13g2_nor2_1 _1876_ (.A(net352),
    .B(net359),
    .Y(_1052_));
 sg13g2_a21oi_1 _1877_ (.A1(net352),
    .A2(_1051_),
    .Y(_0106_),
    .B1(_1052_));
 sg13g2_nand4_1 _1878_ (.B(net305),
    .C(\inst_calculator.reg_operator[0] ),
    .A(net298),
    .Y(_1053_),
    .D(net348));
 sg13g2_mux2_1 _1879_ (.A0(net333),
    .A1(net245),
    .S(net280),
    .X(_0107_));
 sg13g2_mux2_1 _1880_ (.A0(net330),
    .A1(net228),
    .S(net280),
    .X(_0108_));
 sg13g2_mux2_1 _1881_ (.A0(net327),
    .A1(net237),
    .S(net281),
    .X(_0109_));
 sg13g2_nand2_1 _1882_ (.Y(_1054_),
    .A(net124),
    .B(net280));
 sg13g2_o21ai_1 _1883_ (.B1(_1054_),
    .Y(_0110_),
    .A1(_0572_),
    .A2(net282));
 sg13g2_nand2_1 _1884_ (.Y(_1055_),
    .A(net128),
    .B(net281));
 sg13g2_o21ai_1 _1885_ (.B1(_1055_),
    .Y(_0111_),
    .A1(_0571_),
    .A2(net282));
 sg13g2_nand2_1 _1886_ (.Y(_1056_),
    .A(net112),
    .B(net283));
 sg13g2_o21ai_1 _1887_ (.B1(_1056_),
    .Y(_0112_),
    .A1(_0570_),
    .A2(net283));
 sg13g2_nand2_1 _1888_ (.Y(_1057_),
    .A(net115),
    .B(net283));
 sg13g2_o21ai_1 _1889_ (.B1(_1057_),
    .Y(_0113_),
    .A1(_0569_),
    .A2(net283));
 sg13g2_nand2_1 _1890_ (.Y(_1058_),
    .A(net140),
    .B(net283));
 sg13g2_o21ai_1 _1891_ (.B1(_1058_),
    .Y(_0114_),
    .A1(_0568_),
    .A2(net283));
 sg13g2_mux2_1 _1892_ (.A0(net313),
    .A1(net235),
    .S(net284),
    .X(_0115_));
 sg13g2_mux2_1 _1893_ (.A0(\inst_calculator.reg_arg[9] ),
    .A1(net259),
    .S(net284),
    .X(_0116_));
 sg13g2_a21oi_1 _1894_ (.A1(\inst_calculator.inst_divider.busy ),
    .A2(_1039_),
    .Y(_1059_),
    .B1(net309));
 sg13g2_mux2_1 _1895_ (.A0(net96),
    .A1(\inst_calculator.divider_done ),
    .S(_1059_),
    .X(_0117_));
 sg13g2_mux2_1 _1896_ (.A0(\inst_calculator.inst_divider.d[0] ),
    .A1(net245),
    .S(net307),
    .X(_0118_));
 sg13g2_mux2_1 _1897_ (.A0(\inst_calculator.inst_divider.d[1] ),
    .A1(net228),
    .S(net306),
    .X(_0119_));
 sg13g2_mux2_1 _1898_ (.A0(\inst_calculator.inst_divider.d[2] ),
    .A1(net237),
    .S(net307),
    .X(_0120_));
 sg13g2_mux2_1 _1899_ (.A0(net204),
    .A1(net124),
    .S(net306),
    .X(_0121_));
 sg13g2_mux2_1 _1900_ (.A0(net150),
    .A1(net128),
    .S(net306),
    .X(_0122_));
 sg13g2_mux2_1 _1901_ (.A0(net208),
    .A1(net112),
    .S(net308),
    .X(_0123_));
 sg13g2_nand2_1 _1902_ (.Y(_1060_),
    .A(net308),
    .B(net115));
 sg13g2_o21ai_1 _1903_ (.B1(_1060_),
    .Y(_0124_),
    .A1(net308),
    .A2(_0577_));
 sg13g2_nand2_1 _1904_ (.Y(_1061_),
    .A(net308),
    .B(net140));
 sg13g2_o21ai_1 _1905_ (.B1(_1061_),
    .Y(_0125_),
    .A1(net309),
    .A2(_0576_));
 sg13g2_mux2_1 _1906_ (.A0(\inst_calculator.inst_divider.d[8] ),
    .A1(net235),
    .S(net309),
    .X(_0126_));
 sg13g2_mux2_1 _1907_ (.A0(net218),
    .A1(\inst_calculator.denominator[9] ),
    .S(net310),
    .X(_0127_));
 sg13g2_nand2_1 _1908_ (.Y(_1062_),
    .A(\inst_calculator.inst_divider.d[0] ),
    .B(_1040_));
 sg13g2_a221oi_1 _1909_ (.B2(net142),
    .C1(net307),
    .B1(_1062_),
    .A1(_1026_),
    .Y(_1063_),
    .A2(_1040_));
 sg13g2_a21oi_1 _1910_ (.A1(net307),
    .A2(_0588_),
    .Y(_0128_),
    .B1(net143));
 sg13g2_xnor2_1 _1911_ (.Y(_1064_),
    .A(_1025_),
    .B(_1027_));
 sg13g2_a22oi_1 _1912_ (.Y(_1065_),
    .B1(net265),
    .B2(net214),
    .A2(net138),
    .A1(net306));
 sg13g2_o21ai_1 _1913_ (.B1(_1065_),
    .Y(_0129_),
    .A1(_1041_),
    .A2(_1064_));
 sg13g2_xnor2_1 _1914_ (.Y(_1066_),
    .A(_1023_),
    .B(_1028_));
 sg13g2_a22oi_1 _1915_ (.Y(_1067_),
    .B1(net265),
    .B2(net377),
    .A2(net122),
    .A1(net306));
 sg13g2_o21ai_1 _1916_ (.B1(_1067_),
    .Y(_0130_),
    .A1(_1041_),
    .A2(_1066_));
 sg13g2_xnor2_1 _1917_ (.Y(_1068_),
    .A(_1021_),
    .B(_1029_));
 sg13g2_a22oi_1 _1918_ (.Y(_1069_),
    .B1(net265),
    .B2(net257),
    .A2(net132),
    .A1(net306));
 sg13g2_o21ai_1 _1919_ (.B1(_1069_),
    .Y(_0131_),
    .A1(_1041_),
    .A2(_1068_));
 sg13g2_xnor2_1 _1920_ (.Y(_1070_),
    .A(_1019_),
    .B(_1030_));
 sg13g2_a22oi_1 _1921_ (.Y(_1071_),
    .B1(net265),
    .B2(net249),
    .A2(net146),
    .A1(net306));
 sg13g2_o21ai_1 _1922_ (.B1(_1071_),
    .Y(_0132_),
    .A1(_1041_),
    .A2(_1070_));
 sg13g2_xnor2_1 _1923_ (.Y(_1072_),
    .A(_1017_),
    .B(_1031_));
 sg13g2_a22oi_1 _1924_ (.Y(_1073_),
    .B1(net265),
    .B2(net244),
    .A2(net126),
    .A1(net306));
 sg13g2_o21ai_1 _1925_ (.B1(_1073_),
    .Y(_0133_),
    .A1(_1041_),
    .A2(_1072_));
 sg13g2_xnor2_1 _1926_ (.Y(_1074_),
    .A(_1015_),
    .B(_1032_));
 sg13g2_a22oi_1 _1927_ (.Y(_1075_),
    .B1(_1051_),
    .B2(net261),
    .A2(net216),
    .A1(net308));
 sg13g2_o21ai_1 _1928_ (.B1(_1075_),
    .Y(_0134_),
    .A1(_1041_),
    .A2(_1074_));
 sg13g2_xor2_1 _1929_ (.B(_1034_),
    .A(_1014_),
    .X(_1076_));
 sg13g2_a22oi_1 _1930_ (.Y(_1077_),
    .B1(net265),
    .B2(net373),
    .A2(net223),
    .A1(net309));
 sg13g2_o21ai_1 _1931_ (.B1(_1077_),
    .Y(_0135_),
    .A1(_1041_),
    .A2(_1076_));
 sg13g2_xor2_1 _1932_ (.B(net399),
    .A(\inst_calculator.inst_divider.d[8] ),
    .X(_1078_));
 sg13g2_xnor2_1 _1933_ (.Y(_1079_),
    .A(_1036_),
    .B(_1078_));
 sg13g2_a22oi_1 _1934_ (.Y(_1080_),
    .B1(net265),
    .B2(net399),
    .A2(net360),
    .A1(net309));
 sg13g2_o21ai_1 _1935_ (.B1(_1080_),
    .Y(_0136_),
    .A1(_1041_),
    .A2(_1079_));
 sg13g2_nand4_1 _1936_ (.B(\inst_calculator.inst_divider.busy ),
    .C(_1011_),
    .A(_0562_),
    .Y(_1081_),
    .D(_1037_));
 sg13g2_a22oi_1 _1937_ (.Y(_1082_),
    .B1(net265),
    .B2(net225),
    .A2(\inst_calculator.inst_divider.numerator[9] ),
    .A1(net308));
 sg13g2_nand2_1 _1938_ (.Y(_0137_),
    .A(_1081_),
    .B(net226));
 sg13g2_o21ai_1 _1939_ (.B1(_0616_),
    .Y(_1083_),
    .A1(\inst_calculator.inst_keypad_poller.state[5] ),
    .A2(net102));
 sg13g2_a22oi_1 _1940_ (.Y(_1084_),
    .B1(net195),
    .B2(_1083_),
    .A2(\inst_calculator.inst_keypad_poller.state[5] ),
    .A1(net1));
 sg13g2_inv_1 _1941_ (.Y(_0138_),
    .A(net196));
 sg13g2_a22oi_1 _1942_ (.Y(_0193_),
    .B1(net379),
    .B2(_1083_),
    .A2(\inst_calculator.inst_keypad_poller.state[5] ),
    .A1(net2));
 sg13g2_inv_1 _1943_ (.Y(_0139_),
    .A(net380));
 sg13g2_a22oi_1 _1944_ (.Y(_0194_),
    .B1(net402),
    .B2(_1083_),
    .A2(\inst_calculator.inst_keypad_poller.state[5] ),
    .A1(net3));
 sg13g2_inv_1 _1945_ (.Y(_0140_),
    .A(net403));
 sg13g2_a22oi_1 _1946_ (.Y(_0195_),
    .B1(net202),
    .B2(_1083_),
    .A2(\inst_calculator.inst_keypad_poller.state[5] ),
    .A1(net4));
 sg13g2_inv_1 _1947_ (.Y(_0141_),
    .A(net203));
 sg13g2_mux2_1 _1948_ (.A0(net311),
    .A1(_0064_),
    .S(net117),
    .X(_0142_));
 sg13g2_nor2_1 _1949_ (.A(\inst_calculator.inst_drive.cnt_sel[1] ),
    .B(net117),
    .Y(_0196_));
 sg13g2_a21oi_1 _1950_ (.A1(net117),
    .A2(_0608_),
    .Y(_0143_),
    .B1(_0196_));
 sg13g2_mux2_1 _1951_ (.A0(_0061_),
    .A1(net98),
    .S(\inst_calculator.inst_keypad_poller.state[3] ),
    .X(_0144_));
 sg13g2_mux2_1 _1952_ (.A0(net424),
    .A1(net433),
    .S(net263),
    .X(_0145_));
 sg13g2_mux2_1 _1953_ (.A0(net421),
    .A1(net424),
    .S(net263),
    .X(_0146_));
 sg13g2_nand2_1 _1954_ (.Y(_0197_),
    .A(net263),
    .B(net421));
 sg13g2_o21ai_1 _1955_ (.B1(_0197_),
    .Y(_0147_),
    .A1(_0561_),
    .A2(net263));
 sg13g2_a21oi_1 _1956_ (.A1(net145),
    .A2(_0573_),
    .Y(_0198_),
    .B1(net107));
 sg13g2_a21oi_1 _1957_ (.A1(_0567_),
    .A2(_0609_),
    .Y(_0148_),
    .B1(_0198_));
 sg13g2_nand2_1 _1958_ (.Y(_0199_),
    .A(\inst_calculator.state[6] ),
    .B(net349));
 sg13g2_nand2_1 _1959_ (.Y(_0200_),
    .A(net119),
    .B(_0199_));
 sg13g2_o21ai_1 _1960_ (.B1(net120),
    .Y(_0149_),
    .A1(_0567_),
    .A2(_0199_));
 sg13g2_nor2b_2 _1961_ (.A(net305),
    .B_N(\inst_calculator.reg_operator[0] ),
    .Y(_0201_));
 sg13g2_nand2b_1 _1962_ (.Y(_0202_),
    .B(net279),
    .A_N(_0046_));
 sg13g2_or2_1 _1963_ (.X(_0203_),
    .B(net303),
    .A(net299));
 sg13g2_nand4_1 _1964_ (.B(_0611_),
    .C(_0202_),
    .A(net343),
    .Y(_0204_),
    .D(_0203_));
 sg13g2_mux2_1 _1965_ (.A0(net92),
    .A1(net310),
    .S(_0204_),
    .X(_0150_));
 sg13g2_o21ai_1 _1966_ (.B1(net347),
    .Y(_0205_),
    .A1(net298),
    .A2(\inst_calculator.state[0] ));
 sg13g2_and2_1 _1967_ (.A(net298),
    .B(net348),
    .X(_0206_));
 sg13g2_a22oi_1 _1968_ (.Y(_0207_),
    .B1(_0206_),
    .B2(net151),
    .A2(_0205_),
    .A1(\inst_calculator.reg_operator[0] ));
 sg13g2_inv_1 _1969_ (.Y(_0151_),
    .A(net152));
 sg13g2_a22oi_1 _1970_ (.Y(_0208_),
    .B1(_0206_),
    .B2(net134),
    .A2(_0205_),
    .A1(net305));
 sg13g2_inv_1 _1971_ (.Y(_0152_),
    .A(net135));
 sg13g2_nor2_1 _1972_ (.A(net287),
    .B(net280),
    .Y(_0209_));
 sg13g2_a21oi_1 _1973_ (.A1(_0588_),
    .A2(net280),
    .Y(_0153_),
    .B1(_0209_));
 sg13g2_nand2_1 _1974_ (.Y(_0210_),
    .A(net138),
    .B(net281));
 sg13g2_o21ai_1 _1975_ (.B1(_0210_),
    .Y(_0154_),
    .A1(_0583_),
    .A2(net281));
 sg13g2_nand2_1 _1976_ (.Y(_0211_),
    .A(net122),
    .B(net281));
 sg13g2_o21ai_1 _1977_ (.B1(_0211_),
    .Y(_0155_),
    .A1(_0582_),
    .A2(net282));
 sg13g2_nand2_1 _1978_ (.Y(_0212_),
    .A(net132),
    .B(net280));
 sg13g2_o21ai_1 _1979_ (.B1(_0212_),
    .Y(_0156_),
    .A1(_0581_),
    .A2(net281));
 sg13g2_nand2_1 _1980_ (.Y(_0213_),
    .A(net146),
    .B(net280));
 sg13g2_o21ai_1 _1981_ (.B1(_0213_),
    .Y(_0157_),
    .A1(_0580_),
    .A2(net280));
 sg13g2_nand2_1 _1982_ (.Y(_0214_),
    .A(net126),
    .B(net281));
 sg13g2_o21ai_1 _1983_ (.B1(_0214_),
    .Y(_0158_),
    .A1(_0579_),
    .A2(net282));
 sg13g2_mux2_1 _1984_ (.A0(net295),
    .A1(net216),
    .S(net283),
    .X(_0159_));
 sg13g2_mux2_1 _1985_ (.A0(net296),
    .A1(net223),
    .S(net283),
    .X(_0160_));
 sg13g2_mux2_1 _1986_ (.A0(\inst_calculator.reg_result[8] ),
    .A1(net360),
    .S(net284),
    .X(_0161_));
 sg13g2_mux2_1 _1987_ (.A0(\inst_calculator.reg_result[9] ),
    .A1(net255),
    .S(net284),
    .X(_0162_));
 sg13g2_nand2_2 _1988_ (.Y(_0215_),
    .A(net322),
    .B(net292));
 sg13g2_inv_1 _1989_ (.Y(_0216_),
    .A(_0215_));
 sg13g2_and2_2 _1990_ (.A(net325),
    .B(net290),
    .X(_0217_));
 sg13g2_and2_1 _1991_ (.A(net322),
    .B(net290),
    .X(_0218_));
 sg13g2_and2_1 _1992_ (.A(net328),
    .B(net293),
    .X(_0219_));
 sg13g2_a21oi_1 _1993_ (.A1(net325),
    .A2(net292),
    .Y(_0220_),
    .B1(_0218_));
 sg13g2_a21oi_1 _1994_ (.A1(_0216_),
    .A2(_0217_),
    .Y(_0221_),
    .B1(_0220_));
 sg13g2_a22oi_1 _1995_ (.Y(_0222_),
    .B1(_0219_),
    .B2(_0221_),
    .A2(_0217_),
    .A1(_0216_));
 sg13g2_nand2_2 _1996_ (.Y(_0223_),
    .A(net318),
    .B(net288));
 sg13g2_nand2_2 _1997_ (.Y(_0224_),
    .A(net320),
    .B(net286));
 sg13g2_nor2_2 _1998_ (.A(_0223_),
    .B(_0224_),
    .Y(_0225_));
 sg13g2_nand2_1 _1999_ (.Y(_0226_),
    .A(net328),
    .B(net294));
 sg13g2_nand2_1 _2000_ (.Y(_0227_),
    .A(net322),
    .B(net293));
 sg13g2_nand2_1 _2001_ (.Y(_0228_),
    .A(net325),
    .B(net293));
 sg13g2_xor2_1 _2002_ (.B(_0228_),
    .A(_0215_),
    .X(_0229_));
 sg13g2_nand2b_1 _2003_ (.Y(_0230_),
    .B(_0229_),
    .A_N(_0226_));
 sg13g2_xnor2_1 _2004_ (.Y(_0231_),
    .A(_0226_),
    .B(_0229_));
 sg13g2_nand2_1 _2005_ (.Y(_0232_),
    .A(_0225_),
    .B(_0231_));
 sg13g2_nor2_1 _2006_ (.A(_0225_),
    .B(_0231_),
    .Y(_0233_));
 sg13g2_xor2_1 _2007_ (.B(_0231_),
    .A(_0225_),
    .X(_0234_));
 sg13g2_xnor2_1 _2008_ (.Y(_0235_),
    .A(_0222_),
    .B(_0234_));
 sg13g2_nand2_1 _2009_ (.Y(_0236_),
    .A(net320),
    .B(net290));
 sg13g2_nand2_1 _2010_ (.Y(_0237_),
    .A(net315),
    .B(net286));
 sg13g2_or2_1 _2011_ (.X(_0238_),
    .B(_0237_),
    .A(_0223_));
 sg13g2_xor2_1 _2012_ (.B(_0237_),
    .A(_0223_),
    .X(_0239_));
 sg13g2_nand2b_1 _2013_ (.Y(_0240_),
    .B(_0239_),
    .A_N(_0236_));
 sg13g2_xnor2_1 _2014_ (.Y(_0241_),
    .A(_0236_),
    .B(_0239_));
 sg13g2_nand2_1 _2015_ (.Y(_0242_),
    .A(_0235_),
    .B(_0241_));
 sg13g2_xor2_1 _2016_ (.B(_0241_),
    .A(_0235_),
    .X(_0243_));
 sg13g2_xor2_1 _2017_ (.B(_0221_),
    .A(_0219_),
    .X(_0244_));
 sg13g2_and2_1 _2018_ (.A(net325),
    .B(net288),
    .X(_0245_));
 sg13g2_nand2_1 _2019_ (.Y(_0246_),
    .A(net322),
    .B(net288));
 sg13g2_and2_1 _2020_ (.A(net328),
    .B(net292),
    .X(_0247_));
 sg13g2_xnor2_1 _2021_ (.Y(_0248_),
    .A(_0217_),
    .B(_0246_));
 sg13g2_a22oi_1 _2022_ (.Y(_0249_),
    .B1(_0247_),
    .B2(_0248_),
    .A2(_0245_),
    .A1(_0218_));
 sg13g2_nor2b_1 _2023_ (.A(_0249_),
    .B_N(_0244_),
    .Y(_0250_));
 sg13g2_xnor2_1 _2024_ (.Y(_0251_),
    .A(_0244_),
    .B(_0249_));
 sg13g2_a22oi_1 _2025_ (.Y(_0252_),
    .B1(net286),
    .B2(net318),
    .A2(net288),
    .A1(net320));
 sg13g2_nor2_1 _2026_ (.A(_0225_),
    .B(_0252_),
    .Y(_0253_));
 sg13g2_a21o_1 _2027_ (.A2(_0253_),
    .A1(_0251_),
    .B1(_0250_),
    .X(_0254_));
 sg13g2_nand2_1 _2028_ (.Y(_0255_),
    .A(_0243_),
    .B(_0254_));
 sg13g2_o21ai_1 _2029_ (.B1(_0232_),
    .Y(_0256_),
    .A1(_0222_),
    .A2(_0233_));
 sg13g2_o21ai_1 _2030_ (.B1(_0230_),
    .Y(_0257_),
    .A1(_0215_),
    .A2(_0228_));
 sg13g2_and2_1 _2031_ (.A(_0238_),
    .B(_0240_),
    .X(_0258_));
 sg13g2_nand2_1 _2032_ (.Y(_0259_),
    .A(net328),
    .B(net295));
 sg13g2_nand2_1 _2033_ (.Y(_0260_),
    .A(net322),
    .B(net294));
 sg13g2_nand2_1 _2034_ (.Y(_0261_),
    .A(net325),
    .B(net294));
 sg13g2_xor2_1 _2035_ (.B(_0261_),
    .A(_0227_),
    .X(_0262_));
 sg13g2_nand2b_1 _2036_ (.Y(_0263_),
    .B(_0262_),
    .A_N(_0259_));
 sg13g2_xnor2_1 _2037_ (.Y(_0264_),
    .A(_0259_),
    .B(_0262_));
 sg13g2_nor2b_1 _2038_ (.A(_0258_),
    .B_N(_0264_),
    .Y(_0265_));
 sg13g2_xnor2_1 _2039_ (.Y(_0266_),
    .A(_0258_),
    .B(_0264_));
 sg13g2_xnor2_1 _2040_ (.Y(_0267_),
    .A(_0257_),
    .B(_0266_));
 sg13g2_nand2_2 _2041_ (.Y(_0268_),
    .A(net314),
    .B(net287));
 sg13g2_nor2_1 _2042_ (.A(_0571_),
    .B(_0581_),
    .Y(_0269_));
 sg13g2_nor3_1 _2043_ (.A(_0569_),
    .B(_0582_),
    .C(_0223_),
    .Y(_0270_));
 sg13g2_a22oi_1 _2044_ (.Y(_0271_),
    .B1(net288),
    .B2(net315),
    .A2(net291),
    .A1(net318));
 sg13g2_nor2_1 _2045_ (.A(_0270_),
    .B(_0271_),
    .Y(_0272_));
 sg13g2_xor2_1 _2046_ (.B(_0272_),
    .A(_0269_),
    .X(_0273_));
 sg13g2_nand2b_1 _2047_ (.Y(_0274_),
    .B(_0273_),
    .A_N(_0268_));
 sg13g2_xnor2_1 _2048_ (.Y(_0275_),
    .A(_0268_),
    .B(_0273_));
 sg13g2_nand2b_1 _2049_ (.Y(_0276_),
    .B(_0275_),
    .A_N(_0267_));
 sg13g2_xor2_1 _2050_ (.B(_0275_),
    .A(_0267_),
    .X(_0277_));
 sg13g2_nor2_1 _2051_ (.A(_0242_),
    .B(_0277_),
    .Y(_0278_));
 sg13g2_xor2_1 _2052_ (.B(_0277_),
    .A(_0242_),
    .X(_0279_));
 sg13g2_xnor2_1 _2053_ (.Y(_0280_),
    .A(_0256_),
    .B(_0279_));
 sg13g2_nor2_1 _2054_ (.A(_0255_),
    .B(_0280_),
    .Y(_0281_));
 sg13g2_and2_1 _2055_ (.A(net333),
    .B(net296),
    .X(_0282_));
 sg13g2_xor2_1 _2056_ (.B(_0280_),
    .A(_0255_),
    .X(_0283_));
 sg13g2_a21oi_1 _2057_ (.A1(_0282_),
    .A2(_0283_),
    .Y(_0284_),
    .B1(_0281_));
 sg13g2_nand2_1 _2058_ (.Y(_0285_),
    .A(net333),
    .B(\inst_calculator.reg_result[8] ));
 sg13g2_a21oi_1 _2059_ (.A1(_0256_),
    .A2(_0279_),
    .Y(_0286_),
    .B1(_0278_));
 sg13g2_a21o_1 _2060_ (.A2(_0266_),
    .A1(_0257_),
    .B1(_0265_),
    .X(_0287_));
 sg13g2_nand2_1 _2061_ (.Y(_0288_),
    .A(net313),
    .B(net289));
 sg13g2_nor2_1 _2062_ (.A(_0268_),
    .B(_0288_),
    .Y(_0289_));
 sg13g2_a22oi_1 _2063_ (.Y(_0290_),
    .B1(net287),
    .B2(net313),
    .A2(net288),
    .A1(net314));
 sg13g2_nor2_1 _2064_ (.A(_0289_),
    .B(_0290_),
    .Y(_0291_));
 sg13g2_nand2_1 _2065_ (.Y(_0292_),
    .A(net320),
    .B(net293));
 sg13g2_inv_1 _2066_ (.Y(_0293_),
    .A(_0292_));
 sg13g2_a22oi_1 _2067_ (.Y(_0294_),
    .B1(net290),
    .B2(net315),
    .A2(net292),
    .A1(net318));
 sg13g2_nand2_1 _2068_ (.Y(_0295_),
    .A(net315),
    .B(net292));
 sg13g2_nand4_1 _2069_ (.B(net318),
    .C(net292),
    .A(net315),
    .Y(_0296_),
    .D(net290));
 sg13g2_nand2b_1 _2070_ (.Y(_0297_),
    .B(_0296_),
    .A_N(_0294_));
 sg13g2_xnor2_1 _2071_ (.Y(_0298_),
    .A(_0293_),
    .B(_0297_));
 sg13g2_nand2_1 _2072_ (.Y(_0299_),
    .A(_0291_),
    .B(_0298_));
 sg13g2_xnor2_1 _2073_ (.Y(_0300_),
    .A(_0291_),
    .B(_0298_));
 sg13g2_nor2_1 _2074_ (.A(_0274_),
    .B(_0300_),
    .Y(_0301_));
 sg13g2_xor2_1 _2075_ (.B(_0300_),
    .A(_0274_),
    .X(_0302_));
 sg13g2_o21ai_1 _2076_ (.B1(_0263_),
    .Y(_0303_),
    .A1(_0227_),
    .A2(_0261_));
 sg13g2_a21oi_2 _2077_ (.B1(_0270_),
    .Y(_0304_),
    .A2(_0272_),
    .A1(_0269_));
 sg13g2_nand2_1 _2078_ (.Y(_0305_),
    .A(net328),
    .B(net296));
 sg13g2_nand2_1 _2079_ (.Y(_0306_),
    .A(net322),
    .B(net295));
 sg13g2_nand2_1 _2080_ (.Y(_0307_),
    .A(net325),
    .B(net295));
 sg13g2_xor2_1 _2081_ (.B(_0307_),
    .A(_0260_),
    .X(_0308_));
 sg13g2_nand2b_1 _2082_ (.Y(_0309_),
    .B(_0308_),
    .A_N(_0305_));
 sg13g2_xnor2_1 _2083_ (.Y(_0310_),
    .A(_0305_),
    .B(_0308_));
 sg13g2_nor2b_1 _2084_ (.A(_0304_),
    .B_N(_0310_),
    .Y(_0311_));
 sg13g2_xnor2_1 _2085_ (.Y(_0312_),
    .A(_0304_),
    .B(_0310_));
 sg13g2_xor2_1 _2086_ (.B(_0312_),
    .A(_0303_),
    .X(_0313_));
 sg13g2_xnor2_1 _2087_ (.Y(_0314_),
    .A(_0302_),
    .B(_0313_));
 sg13g2_nor2_1 _2088_ (.A(_0276_),
    .B(_0314_),
    .Y(_0315_));
 sg13g2_xor2_1 _2089_ (.B(_0314_),
    .A(_0276_),
    .X(_0316_));
 sg13g2_xnor2_1 _2090_ (.Y(_0317_),
    .A(_0287_),
    .B(_0316_));
 sg13g2_xor2_1 _2091_ (.B(_0317_),
    .A(_0286_),
    .X(_0318_));
 sg13g2_nand2b_1 _2092_ (.Y(_0319_),
    .B(_0318_),
    .A_N(_0285_));
 sg13g2_xnor2_1 _2093_ (.Y(_0320_),
    .A(_0285_),
    .B(_0318_));
 sg13g2_inv_1 _2094_ (.Y(_0321_),
    .A(_0320_));
 sg13g2_xor2_1 _2095_ (.B(_0254_),
    .A(_0243_),
    .X(_0322_));
 sg13g2_xor2_1 _2096_ (.B(_0253_),
    .A(_0251_),
    .X(_0323_));
 sg13g2_xor2_1 _2097_ (.B(_0248_),
    .A(_0247_),
    .X(_0324_));
 sg13g2_nand2_1 _2098_ (.Y(_0325_),
    .A(net325),
    .B(net286));
 sg13g2_nand2_1 _2099_ (.Y(_0326_),
    .A(net322),
    .B(net286));
 sg13g2_nor2_1 _2100_ (.A(_0246_),
    .B(_0325_),
    .Y(_0327_));
 sg13g2_and2_1 _2101_ (.A(net328),
    .B(net290),
    .X(_0328_));
 sg13g2_xnor2_1 _2102_ (.Y(_0329_),
    .A(_0245_),
    .B(_0326_));
 sg13g2_a21oi_1 _2103_ (.A1(_0328_),
    .A2(_0329_),
    .Y(_0330_),
    .B1(_0327_));
 sg13g2_nand2b_1 _2104_ (.Y(_0331_),
    .B(_0324_),
    .A_N(_0330_));
 sg13g2_xnor2_1 _2105_ (.Y(_0332_),
    .A(_0324_),
    .B(_0330_));
 sg13g2_nand2b_1 _2106_ (.Y(_0333_),
    .B(_0332_),
    .A_N(_0224_));
 sg13g2_nand2_1 _2107_ (.Y(_0334_),
    .A(_0331_),
    .B(_0333_));
 sg13g2_nand2_1 _2108_ (.Y(_0335_),
    .A(_0323_),
    .B(_0334_));
 sg13g2_inv_1 _2109_ (.Y(_0336_),
    .A(_0335_));
 sg13g2_nand2_1 _2110_ (.Y(_0337_),
    .A(net333),
    .B(net295));
 sg13g2_xor2_1 _2111_ (.B(_0335_),
    .A(_0322_),
    .X(_0338_));
 sg13g2_nor2_1 _2112_ (.A(_0337_),
    .B(_0338_),
    .Y(_0339_));
 sg13g2_a21oi_1 _2113_ (.A1(_0322_),
    .A2(_0336_),
    .Y(_0340_),
    .B1(_0339_));
 sg13g2_xor2_1 _2114_ (.B(_0283_),
    .A(_0282_),
    .X(_0341_));
 sg13g2_nor2b_1 _2115_ (.A(_0340_),
    .B_N(_0341_),
    .Y(_0342_));
 sg13g2_and2_1 _2116_ (.A(net328),
    .B(net286),
    .X(_0343_));
 sg13g2_nand2_1 _2117_ (.Y(_0344_),
    .A(_0245_),
    .B(_0343_));
 sg13g2_xor2_1 _2118_ (.B(_0329_),
    .A(_0328_),
    .X(_0345_));
 sg13g2_nand2b_1 _2119_ (.Y(_0346_),
    .B(_0345_),
    .A_N(_0344_));
 sg13g2_xnor2_1 _2120_ (.Y(_0347_),
    .A(_0224_),
    .B(_0332_));
 sg13g2_nor2b_1 _2121_ (.A(_0346_),
    .B_N(_0347_),
    .Y(_0348_));
 sg13g2_xor2_1 _2122_ (.B(_0334_),
    .A(_0323_),
    .X(_0349_));
 sg13g2_nand2_1 _2123_ (.Y(_0350_),
    .A(net333),
    .B(net294));
 sg13g2_xnor2_1 _2124_ (.Y(_0351_),
    .A(_0348_),
    .B(_0349_));
 sg13g2_nor2_1 _2125_ (.A(_0350_),
    .B(_0351_),
    .Y(_0352_));
 sg13g2_a21oi_1 _2126_ (.A1(_0348_),
    .A2(_0349_),
    .Y(_0353_),
    .B1(_0352_));
 sg13g2_xor2_1 _2127_ (.B(_0338_),
    .A(_0337_),
    .X(_0354_));
 sg13g2_nor2b_1 _2128_ (.A(_0353_),
    .B_N(_0354_),
    .Y(_0355_));
 sg13g2_nand2_1 _2129_ (.Y(_0356_),
    .A(net333),
    .B(net293));
 sg13g2_xnor2_1 _2130_ (.Y(_0357_),
    .A(_0346_),
    .B(_0347_));
 sg13g2_nor2b_1 _2131_ (.A(_0356_),
    .B_N(_0357_),
    .Y(_0358_));
 sg13g2_and2_1 _2132_ (.A(net333),
    .B(net292),
    .X(_0359_));
 sg13g2_xnor2_1 _2133_ (.Y(_0360_),
    .A(_0344_),
    .B(_0345_));
 sg13g2_nand2_1 _2134_ (.Y(_0361_),
    .A(net331),
    .B(net290));
 sg13g2_nand2_2 _2135_ (.Y(_0362_),
    .A(net328),
    .B(net289));
 sg13g2_a22oi_1 _2136_ (.Y(_0363_),
    .B1(_0362_),
    .B2(_0325_),
    .A2(_0343_),
    .A1(_0245_));
 sg13g2_nor2b_1 _2137_ (.A(_0361_),
    .B_N(_0363_),
    .Y(_0364_));
 sg13g2_nand2_2 _2138_ (.Y(_0365_),
    .A(net331),
    .B(net287));
 sg13g2_nor2_1 _2139_ (.A(_0362_),
    .B(_0365_),
    .Y(_0366_));
 sg13g2_xnor2_1 _2140_ (.Y(_0367_),
    .A(_0361_),
    .B(_0363_));
 sg13g2_a21oi_1 _2141_ (.A1(_0366_),
    .A2(_0367_),
    .Y(_0368_),
    .B1(_0364_));
 sg13g2_xor2_1 _2142_ (.B(_0360_),
    .A(_0359_),
    .X(_0369_));
 sg13g2_nor2b_1 _2143_ (.A(_0368_),
    .B_N(_0369_),
    .Y(_0370_));
 sg13g2_a21oi_1 _2144_ (.A1(_0359_),
    .A2(_0360_),
    .Y(_0371_),
    .B1(_0370_));
 sg13g2_xnor2_1 _2145_ (.Y(_0372_),
    .A(_0356_),
    .B(_0357_));
 sg13g2_nor2b_1 _2146_ (.A(_0371_),
    .B_N(_0372_),
    .Y(_0373_));
 sg13g2_nor2_1 _2147_ (.A(_0358_),
    .B(_0373_),
    .Y(_0374_));
 sg13g2_xor2_1 _2148_ (.B(_0351_),
    .A(_0350_),
    .X(_0375_));
 sg13g2_nor2b_1 _2149_ (.A(_0374_),
    .B_N(_0375_),
    .Y(_0376_));
 sg13g2_xnor2_1 _2150_ (.Y(_0377_),
    .A(_0353_),
    .B(_0354_));
 sg13g2_a21o_1 _2151_ (.A2(_0377_),
    .A1(_0376_),
    .B1(_0355_),
    .X(_0378_));
 sg13g2_xnor2_1 _2152_ (.Y(_0379_),
    .A(_0340_),
    .B(_0341_));
 sg13g2_a21oi_2 _2153_ (.B1(_0342_),
    .Y(_0380_),
    .A2(_0379_),
    .A1(_0378_));
 sg13g2_xnor2_1 _2154_ (.Y(_0381_),
    .A(_0284_),
    .B(_0320_));
 sg13g2_nand2b_1 _2155_ (.Y(_0382_),
    .B(_0381_),
    .A_N(_0380_));
 sg13g2_o21ai_1 _2156_ (.B1(_0382_),
    .Y(_0383_),
    .A1(_0284_),
    .A2(_0321_));
 sg13g2_o21ai_1 _2157_ (.B1(_0319_),
    .Y(_0384_),
    .A1(_0286_),
    .A2(_0317_));
 sg13g2_a21oi_1 _2158_ (.A1(_0287_),
    .A2(_0316_),
    .Y(_0385_),
    .B1(_0315_));
 sg13g2_a21oi_1 _2159_ (.A1(_0302_),
    .A2(_0313_),
    .Y(_0386_),
    .B1(_0301_));
 sg13g2_a21oi_1 _2160_ (.A1(_0303_),
    .A2(_0312_),
    .Y(_0387_),
    .B1(_0311_));
 sg13g2_xnor2_1 _2161_ (.Y(_0388_),
    .A(_0386_),
    .B(_0387_));
 sg13g2_o21ai_1 _2162_ (.B1(_0309_),
    .Y(_0389_),
    .A1(_0260_),
    .A2(_0307_));
 sg13g2_nand2_1 _2163_ (.Y(_0390_),
    .A(net320),
    .B(net294));
 sg13g2_nand2_1 _2164_ (.Y(_0391_),
    .A(net317),
    .B(net293));
 sg13g2_xnor2_1 _2165_ (.Y(_0392_),
    .A(_0295_),
    .B(_0391_));
 sg13g2_xnor2_1 _2166_ (.Y(_0393_),
    .A(_0390_),
    .B(_0392_));
 sg13g2_xnor2_1 _2167_ (.Y(_0394_),
    .A(_0389_),
    .B(_0393_));
 sg13g2_nor3_1 _2168_ (.A(_0568_),
    .B(_0582_),
    .C(_0289_),
    .Y(_0395_));
 sg13g2_a21oi_1 _2169_ (.A1(_0582_),
    .A2(_0289_),
    .Y(_0396_),
    .B1(_0395_));
 sg13g2_nand2_1 _2170_ (.Y(_0397_),
    .A(\inst_calculator.reg_arg[9] ),
    .B(net286));
 sg13g2_xor2_1 _2171_ (.B(_0397_),
    .A(_0288_),
    .X(_0398_));
 sg13g2_xnor2_1 _2172_ (.Y(_0399_),
    .A(_0396_),
    .B(_0398_));
 sg13g2_xnor2_1 _2173_ (.Y(_0400_),
    .A(_0296_),
    .B(_0299_));
 sg13g2_o21ai_1 _2174_ (.B1(_0400_),
    .Y(_0401_),
    .A1(_0292_),
    .A2(_0297_));
 sg13g2_nand2_1 _2175_ (.Y(_0402_),
    .A(net326),
    .B(net296));
 sg13g2_xor2_1 _2176_ (.B(_0402_),
    .A(_0306_),
    .X(_0403_));
 sg13g2_nand2_1 _2177_ (.Y(_0404_),
    .A(net331),
    .B(\inst_calculator.reg_result[9] ));
 sg13g2_nand2_1 _2178_ (.Y(_0405_),
    .A(net330),
    .B(\inst_calculator.reg_result[8] ));
 sg13g2_xnor2_1 _2179_ (.Y(_0406_),
    .A(_0404_),
    .B(_0405_));
 sg13g2_xnor2_1 _2180_ (.Y(_0407_),
    .A(_0403_),
    .B(_0406_));
 sg13g2_xnor2_1 _2181_ (.Y(_0408_),
    .A(_0399_),
    .B(_0407_));
 sg13g2_xnor2_1 _2182_ (.Y(_0409_),
    .A(_0394_),
    .B(_0408_));
 sg13g2_xnor2_1 _2183_ (.Y(_0410_),
    .A(_0401_),
    .B(_0409_));
 sg13g2_xnor2_1 _2184_ (.Y(_0411_),
    .A(_0388_),
    .B(_0410_));
 sg13g2_xor2_1 _2185_ (.B(_0411_),
    .A(_0385_),
    .X(_0412_));
 sg13g2_xnor2_1 _2186_ (.Y(_0413_),
    .A(_0384_),
    .B(_0412_));
 sg13g2_o21ai_1 _2187_ (.B1(net304),
    .Y(_0414_),
    .A1(_0383_),
    .A2(_0413_));
 sg13g2_a21oi_1 _2188_ (.A1(_0383_),
    .A2(_0413_),
    .Y(_0415_),
    .B1(_0414_));
 sg13g2_xnor2_1 _2189_ (.Y(_0416_),
    .A(\inst_calculator.reg_arg[9] ),
    .B(\inst_calculator.reg_result[9] ));
 sg13g2_nand2b_1 _2190_ (.Y(_0417_),
    .B(\inst_calculator.reg_result[8] ),
    .A_N(\inst_calculator.reg_arg[8] ));
 sg13g2_xor2_1 _2191_ (.B(\inst_calculator.reg_result[8] ),
    .A(\inst_calculator.reg_arg[8] ),
    .X(_0418_));
 sg13g2_xnor2_1 _2192_ (.Y(_0419_),
    .A(\inst_calculator.reg_arg[7] ),
    .B(net296));
 sg13g2_xor2_1 _2193_ (.B(\inst_calculator.reg_result[7] ),
    .A(net314),
    .X(_0420_));
 sg13g2_xor2_1 _2194_ (.B(\inst_calculator.reg_result[6] ),
    .A(net316),
    .X(_0421_));
 sg13g2_inv_1 _2195_ (.Y(_0422_),
    .A(_0421_));
 sg13g2_nand2_1 _2196_ (.Y(_0423_),
    .A(net319),
    .B(net294));
 sg13g2_xor2_1 _2197_ (.B(\inst_calculator.reg_result[5] ),
    .A(net319),
    .X(_0424_));
 sg13g2_xor2_1 _2198_ (.B(net293),
    .A(net320),
    .X(_0425_));
 sg13g2_inv_1 _2199_ (.Y(_0426_),
    .A(_0425_));
 sg13g2_xor2_1 _2200_ (.B(\inst_calculator.reg_result[3] ),
    .A(net322),
    .X(_0427_));
 sg13g2_nor2_1 _2201_ (.A(net327),
    .B(_0582_),
    .Y(_0428_));
 sg13g2_xor2_1 _2202_ (.B(net291),
    .A(net327),
    .X(_0429_));
 sg13g2_inv_1 _2203_ (.Y(_0430_),
    .A(_0429_));
 sg13g2_xor2_1 _2204_ (.B(net289),
    .A(net329),
    .X(_0431_));
 sg13g2_nor2b_1 _2205_ (.A(net287),
    .B_N(net331),
    .Y(_0432_));
 sg13g2_nand2b_1 _2206_ (.Y(_0433_),
    .B(net289),
    .A_N(net329));
 sg13g2_o21ai_1 _2207_ (.B1(_0433_),
    .Y(_0434_),
    .A1(_0431_),
    .A2(_0432_));
 sg13g2_a21oi_1 _2208_ (.A1(_0430_),
    .A2(_0434_),
    .Y(_0435_),
    .B1(_0428_));
 sg13g2_nor2_1 _2209_ (.A(_0427_),
    .B(_0435_),
    .Y(_0436_));
 sg13g2_a21oi_1 _2210_ (.A1(_0572_),
    .A2(\inst_calculator.reg_result[3] ),
    .Y(_0437_),
    .B1(_0436_));
 sg13g2_nor2_1 _2211_ (.A(_0425_),
    .B(_0437_),
    .Y(_0438_));
 sg13g2_a21oi_1 _2212_ (.A1(_0571_),
    .A2(\inst_calculator.reg_result[4] ),
    .Y(_0439_),
    .B1(_0438_));
 sg13g2_nor2_1 _2213_ (.A(_0424_),
    .B(_0439_),
    .Y(_0440_));
 sg13g2_a21oi_1 _2214_ (.A1(_0570_),
    .A2(net294),
    .Y(_0441_),
    .B1(_0440_));
 sg13g2_nor2_1 _2215_ (.A(_0421_),
    .B(_0441_),
    .Y(_0442_));
 sg13g2_a21oi_1 _2216_ (.A1(_0569_),
    .A2(net295),
    .Y(_0443_),
    .B1(_0442_));
 sg13g2_nor2_1 _2217_ (.A(_0420_),
    .B(_0443_),
    .Y(_0444_));
 sg13g2_a21oi_1 _2218_ (.A1(_0568_),
    .A2(net296),
    .Y(_0445_),
    .B1(_0444_));
 sg13g2_o21ai_1 _2219_ (.B1(_0417_),
    .Y(_0446_),
    .A1(_0418_),
    .A2(_0445_));
 sg13g2_xnor2_1 _2220_ (.Y(_0447_),
    .A(_0416_),
    .B(_0446_));
 sg13g2_nand2b_1 _2221_ (.Y(_0448_),
    .B(_0431_),
    .A_N(_0365_));
 sg13g2_a21oi_1 _2222_ (.A1(_0362_),
    .A2(_0448_),
    .Y(_0449_),
    .B1(_0430_));
 sg13g2_o21ai_1 _2223_ (.B1(_0427_),
    .Y(_0450_),
    .A1(_0217_),
    .A2(_0449_));
 sg13g2_a21oi_1 _2224_ (.A1(_0215_),
    .A2(_0450_),
    .Y(_0451_),
    .B1(_0426_));
 sg13g2_o21ai_1 _2225_ (.B1(_0424_),
    .Y(_0452_),
    .A1(_0293_),
    .A2(_0451_));
 sg13g2_a21oi_1 _2226_ (.A1(_0423_),
    .A2(_0452_),
    .Y(_0453_),
    .B1(_0422_));
 sg13g2_a21oi_1 _2227_ (.A1(net316),
    .A2(\inst_calculator.reg_result[6] ),
    .Y(_0454_),
    .B1(_0453_));
 sg13g2_nor2_1 _2228_ (.A(_0419_),
    .B(_0454_),
    .Y(_0455_));
 sg13g2_a21oi_1 _2229_ (.A1(\inst_calculator.reg_arg[7] ),
    .A2(\inst_calculator.reg_result[7] ),
    .Y(_0456_),
    .B1(_0455_));
 sg13g2_nor2b_1 _2230_ (.A(_0456_),
    .B_N(_0418_),
    .Y(_0457_));
 sg13g2_a21oi_1 _2231_ (.A1(net313),
    .A2(\inst_calculator.reg_result[8] ),
    .Y(_0458_),
    .B1(_0457_));
 sg13g2_nor2_1 _2232_ (.A(\inst_calculator.reg_operator[1] ),
    .B(\inst_calculator.reg_operator[0] ),
    .Y(_0459_));
 sg13g2_xnor2_1 _2233_ (.Y(_0460_),
    .A(_0416_),
    .B(_0458_));
 sg13g2_a221oi_1 _2234_ (.B2(_0460_),
    .C1(_0415_),
    .B1(net278),
    .A1(net279),
    .Y(_0461_),
    .A2(_0447_));
 sg13g2_a22oi_1 _2235_ (.Y(_0462_),
    .B1(_0461_),
    .B2(net297),
    .A2(net148),
    .A1(net302));
 sg13g2_nand3b_1 _2236_ (.B(\inst_calculator.reg_operator[0] ),
    .C(net305),
    .Y(_0463_),
    .A_N(_0046_));
 sg13g2_nor2_1 _2237_ (.A(net303),
    .B(\inst_calculator.state[0] ),
    .Y(_0464_));
 sg13g2_nand2_1 _2238_ (.Y(_0465_),
    .A(_0046_),
    .B(_0464_));
 sg13g2_nand4_1 _2239_ (.B(_0631_),
    .C(_0463_),
    .A(net343),
    .Y(_0466_),
    .D(_0465_));
 sg13g2_nand2b_2 _2240_ (.Y(_0467_),
    .B(_0203_),
    .A_N(net274));
 sg13g2_nand2_1 _2241_ (.Y(_0468_),
    .A(net404),
    .B(net274));
 sg13g2_o21ai_1 _2242_ (.B1(_0468_),
    .Y(_0163_),
    .A1(_0462_),
    .A2(_0467_));
 sg13g2_nand2_1 _2243_ (.Y(_0469_),
    .A(\inst_calculator.reg_result[8] ),
    .B(net273));
 sg13g2_xor2_1 _2244_ (.B(_0381_),
    .A(_0380_),
    .X(_0470_));
 sg13g2_xor2_1 _2245_ (.B(_0456_),
    .A(_0418_),
    .X(_0471_));
 sg13g2_and2_1 _2246_ (.A(net278),
    .B(_0471_),
    .X(_0472_));
 sg13g2_xnor2_1 _2247_ (.Y(_0473_),
    .A(_0418_),
    .B(_0445_));
 sg13g2_a221oi_1 _2248_ (.B2(_0201_),
    .C1(_0472_),
    .B1(_0473_),
    .A1(net304),
    .Y(_0474_),
    .A2(_0470_));
 sg13g2_a22oi_1 _2249_ (.Y(_0475_),
    .B1(_0474_),
    .B2(net299),
    .A2(net383),
    .A1(net303));
 sg13g2_o21ai_1 _2250_ (.B1(_0469_),
    .Y(_0164_),
    .A1(_0467_),
    .A2(net384));
 sg13g2_nand2_1 _2251_ (.Y(_0476_),
    .A(net296),
    .B(net274));
 sg13g2_xnor2_1 _2252_ (.Y(_0477_),
    .A(_0378_),
    .B(_0379_));
 sg13g2_xnor2_1 _2253_ (.Y(_0478_),
    .A(_0420_),
    .B(_0443_));
 sg13g2_and2_1 _2254_ (.A(net279),
    .B(_0478_),
    .X(_0479_));
 sg13g2_xnor2_1 _2255_ (.Y(_0480_),
    .A(_0419_),
    .B(_0454_));
 sg13g2_a221oi_1 _2256_ (.B2(_0459_),
    .C1(_0479_),
    .B1(_0480_),
    .A1(net305),
    .Y(_0481_),
    .A2(_0477_));
 sg13g2_a22oi_1 _2257_ (.Y(_0482_),
    .B1(_0481_),
    .B2(net297),
    .A2(net234),
    .A1(net303));
 sg13g2_o21ai_1 _2258_ (.B1(_0476_),
    .Y(_0165_),
    .A1(_0467_),
    .A2(_0482_));
 sg13g2_nand2_1 _2259_ (.Y(_0483_),
    .A(net295),
    .B(net274));
 sg13g2_xnor2_1 _2260_ (.Y(_0484_),
    .A(_0376_),
    .B(_0377_));
 sg13g2_nand3_1 _2261_ (.B(_0423_),
    .C(_0452_),
    .A(_0422_),
    .Y(_0485_));
 sg13g2_nor2b_1 _2262_ (.A(_0453_),
    .B_N(_0485_),
    .Y(_0486_));
 sg13g2_nor2b_1 _2263_ (.A(_0486_),
    .B_N(net278),
    .Y(_0487_));
 sg13g2_xnor2_1 _2264_ (.Y(_0488_),
    .A(_0421_),
    .B(_0441_));
 sg13g2_a221oi_1 _2265_ (.B2(_0201_),
    .C1(_0487_),
    .B1(_0488_),
    .A1(net304),
    .Y(_0489_),
    .A2(_0484_));
 sg13g2_a22oi_1 _2266_ (.Y(_0490_),
    .B1(_0489_),
    .B2(net297),
    .A2(net153),
    .A1(net302));
 sg13g2_o21ai_1 _2267_ (.B1(_0483_),
    .Y(_0166_),
    .A1(_0467_),
    .A2(_0490_));
 sg13g2_nor2b_1 _2268_ (.A(_0375_),
    .B_N(_0374_),
    .Y(_0491_));
 sg13g2_o21ai_1 _2269_ (.B1(net304),
    .Y(_0492_),
    .A1(_0376_),
    .A2(_0491_));
 sg13g2_xnor2_1 _2270_ (.Y(_0493_),
    .A(_0424_),
    .B(_0439_));
 sg13g2_or3_1 _2271_ (.A(_0293_),
    .B(_0424_),
    .C(_0451_),
    .X(_0494_));
 sg13g2_nand2_1 _2272_ (.Y(_0495_),
    .A(_0452_),
    .B(_0494_));
 sg13g2_a22oi_1 _2273_ (.Y(_0496_),
    .B1(_0495_),
    .B2(net278),
    .A2(_0493_),
    .A1(net279));
 sg13g2_nand3_1 _2274_ (.B(_0492_),
    .C(_0496_),
    .A(net297),
    .Y(_0497_));
 sg13g2_a21oi_1 _2275_ (.A1(net302),
    .A2(net182),
    .Y(_0498_),
    .B1(net272));
 sg13g2_a22oi_1 _2276_ (.Y(_0167_),
    .B1(_0497_),
    .B2(_0498_),
    .A2(net272),
    .A1(_0579_));
 sg13g2_nor2b_1 _2277_ (.A(_0372_),
    .B_N(_0371_),
    .Y(_0499_));
 sg13g2_o21ai_1 _2278_ (.B1(net304),
    .Y(_0500_),
    .A1(_0373_),
    .A2(_0499_));
 sg13g2_xnor2_1 _2279_ (.Y(_0501_),
    .A(_0425_),
    .B(_0437_));
 sg13g2_nand3_1 _2280_ (.B(_0426_),
    .C(_0450_),
    .A(_0215_),
    .Y(_0502_));
 sg13g2_nand2b_1 _2281_ (.Y(_0503_),
    .B(_0502_),
    .A_N(_0451_));
 sg13g2_a22oi_1 _2282_ (.Y(_0504_),
    .B1(_0503_),
    .B2(net278),
    .A2(_0501_),
    .A1(net279));
 sg13g2_nand3_1 _2283_ (.B(_0500_),
    .C(_0504_),
    .A(net297),
    .Y(_0505_));
 sg13g2_a21oi_1 _2284_ (.A1(net302),
    .A2(net158),
    .Y(_0506_),
    .B1(net272));
 sg13g2_a22oi_1 _2285_ (.Y(_0168_),
    .B1(_0505_),
    .B2(_0506_),
    .A2(net272),
    .A1(_0580_));
 sg13g2_nor2b_1 _2286_ (.A(_0369_),
    .B_N(_0368_),
    .Y(_0507_));
 sg13g2_o21ai_1 _2287_ (.B1(net304),
    .Y(_0508_),
    .A1(_0370_),
    .A2(_0507_));
 sg13g2_or3_1 _2288_ (.A(_0217_),
    .B(_0427_),
    .C(_0449_),
    .X(_0509_));
 sg13g2_nand2_1 _2289_ (.Y(_0510_),
    .A(_0450_),
    .B(_0509_));
 sg13g2_xnor2_1 _2290_ (.Y(_0511_),
    .A(_0427_),
    .B(_0435_));
 sg13g2_a22oi_1 _2291_ (.Y(_0512_),
    .B1(_0511_),
    .B2(net279),
    .A2(_0510_),
    .A1(net278));
 sg13g2_nand3_1 _2292_ (.B(_0508_),
    .C(_0512_),
    .A(net297),
    .Y(_0513_));
 sg13g2_a21oi_1 _2293_ (.A1(net302),
    .A2(net184),
    .Y(_0514_),
    .B1(net272));
 sg13g2_a22oi_1 _2294_ (.Y(_0169_),
    .B1(_0513_),
    .B2(_0514_),
    .A2(net273),
    .A1(_0581_));
 sg13g2_xnor2_1 _2295_ (.Y(_0515_),
    .A(_0366_),
    .B(_0367_));
 sg13g2_nand2_1 _2296_ (.Y(_0516_),
    .A(net304),
    .B(_0515_));
 sg13g2_xnor2_1 _2297_ (.Y(_0517_),
    .A(_0430_),
    .B(_0434_));
 sg13g2_nand3_1 _2298_ (.B(_0430_),
    .C(_0448_),
    .A(_0362_),
    .Y(_0518_));
 sg13g2_nand2b_1 _2299_ (.Y(_0519_),
    .B(_0518_),
    .A_N(_0449_));
 sg13g2_a22oi_1 _2300_ (.Y(_0520_),
    .B1(_0519_),
    .B2(net278),
    .A2(_0517_),
    .A1(net279));
 sg13g2_nand3_1 _2301_ (.B(_0516_),
    .C(_0520_),
    .A(net297),
    .Y(_0521_));
 sg13g2_a21oi_1 _2302_ (.A1(net302),
    .A2(net209),
    .Y(_0522_),
    .B1(net272));
 sg13g2_a22oi_1 _2303_ (.Y(_0170_),
    .B1(_0521_),
    .B2(_0522_),
    .A2(net274),
    .A1(_0582_));
 sg13g2_xor2_1 _2304_ (.B(_0431_),
    .A(_0365_),
    .X(_0523_));
 sg13g2_a21oi_1 _2305_ (.A1(net333),
    .A2(net288),
    .Y(_0524_),
    .B1(_0343_));
 sg13g2_o21ai_1 _2306_ (.B1(net304),
    .Y(_0525_),
    .A1(_0366_),
    .A2(_0524_));
 sg13g2_xnor2_1 _2307_ (.Y(_0526_),
    .A(_0431_),
    .B(_0432_));
 sg13g2_a22oi_1 _2308_ (.Y(_0527_),
    .B1(_0526_),
    .B2(net279),
    .A2(_0523_),
    .A1(net278));
 sg13g2_nand3_1 _2309_ (.B(_0525_),
    .C(_0527_),
    .A(net297),
    .Y(_0528_));
 sg13g2_a21oi_1 _2310_ (.A1(net302),
    .A2(net430),
    .Y(_0529_),
    .B1(net272));
 sg13g2_a22oi_1 _2311_ (.Y(_0171_),
    .B1(_0528_),
    .B2(_0529_),
    .A2(net272),
    .A1(_0583_));
 sg13g2_nor2b_1 _2312_ (.A(_0610_),
    .B_N(_0365_),
    .Y(_0530_));
 sg13g2_o21ai_1 _2313_ (.B1(_0530_),
    .Y(_0531_),
    .A1(net331),
    .A2(net287));
 sg13g2_o21ai_1 _2314_ (.B1(_0531_),
    .Y(_0532_),
    .A1(_0632_),
    .A2(_0365_));
 sg13g2_a21oi_1 _2315_ (.A1(net302),
    .A2(net436),
    .Y(_0533_),
    .B1(_0532_));
 sg13g2_nand2_1 _2316_ (.Y(_0534_),
    .A(net287),
    .B(net273));
 sg13g2_o21ai_1 _2317_ (.B1(_0534_),
    .Y(_0172_),
    .A1(net273),
    .A2(_0533_));
 sg13g2_nor2b_1 _2318_ (.A(_0613_),
    .B_N(net339),
    .Y(_0535_));
 sg13g2_a22oi_1 _2319_ (.Y(_0536_),
    .B1(\inst_calculator.reg_result[9] ),
    .B2(\inst_calculator.state[4] ),
    .A2(\inst_calculator.reg_arg[9] ),
    .A1(\inst_calculator.state[7] ));
 sg13g2_nor2_1 _2320_ (.A(net251),
    .B(net275),
    .Y(_0537_));
 sg13g2_a21oi_1 _2321_ (.A1(net275),
    .A2(_0536_),
    .Y(_0173_),
    .B1(_0537_));
 sg13g2_a22oi_1 _2322_ (.Y(_0538_),
    .B1(\inst_calculator.reg_result[8] ),
    .B2(\inst_calculator.state[4] ),
    .A2(net313),
    .A1(\inst_calculator.state[7] ));
 sg13g2_nor2_1 _2323_ (.A(net428),
    .B(net275),
    .Y(_0539_));
 sg13g2_a21oi_1 _2324_ (.A1(net275),
    .A2(_0538_),
    .Y(_0174_),
    .B1(_0539_));
 sg13g2_a22oi_1 _2325_ (.Y(_0540_),
    .B1(net296),
    .B2(net301),
    .A2(net314),
    .A1(net300));
 sg13g2_nor2_1 _2326_ (.A(net434),
    .B(net275),
    .Y(_0541_));
 sg13g2_a21oi_1 _2327_ (.A1(net275),
    .A2(_0540_),
    .Y(_0175_),
    .B1(_0541_));
 sg13g2_a22oi_1 _2328_ (.Y(_0542_),
    .B1(net295),
    .B2(net301),
    .A2(net316),
    .A1(net300));
 sg13g2_nor2_1 _2329_ (.A(net230),
    .B(net275),
    .Y(_0543_));
 sg13g2_a21oi_1 _2330_ (.A1(net275),
    .A2(_0542_),
    .Y(_0176_),
    .B1(_0543_));
 sg13g2_a22oi_1 _2331_ (.Y(_0544_),
    .B1(net294),
    .B2(net301),
    .A2(net317),
    .A1(net300));
 sg13g2_nor2_1 _2332_ (.A(net375),
    .B(net277),
    .Y(_0545_));
 sg13g2_a21oi_1 _2333_ (.A1(net277),
    .A2(_0544_),
    .Y(_0177_),
    .B1(_0545_));
 sg13g2_a22oi_1 _2334_ (.Y(_0546_),
    .B1(net293),
    .B2(net301),
    .A2(net321),
    .A1(net300));
 sg13g2_nor2_1 _2335_ (.A(net193),
    .B(net277),
    .Y(_0547_));
 sg13g2_a21oi_1 _2336_ (.A1(net276),
    .A2(_0546_),
    .Y(_0178_),
    .B1(_0547_));
 sg13g2_a22oi_1 _2337_ (.Y(_0548_),
    .B1(net292),
    .B2(net301),
    .A2(net323),
    .A1(net300));
 sg13g2_nor2_1 _2338_ (.A(net192),
    .B(net276),
    .Y(_0549_));
 sg13g2_a21oi_1 _2339_ (.A1(net276),
    .A2(_0548_),
    .Y(_0179_),
    .B1(_0549_));
 sg13g2_a22oi_1 _2340_ (.Y(_0550_),
    .B1(net290),
    .B2(net301),
    .A2(net326),
    .A1(net300));
 sg13g2_nor2_1 _2341_ (.A(net181),
    .B(net277),
    .Y(_0551_));
 sg13g2_a21oi_1 _2342_ (.A1(net276),
    .A2(_0550_),
    .Y(_0180_),
    .B1(_0551_));
 sg13g2_a22oi_1 _2343_ (.Y(_0552_),
    .B1(net288),
    .B2(net301),
    .A2(net329),
    .A1(net300));
 sg13g2_nor2_1 _2344_ (.A(net205),
    .B(net276),
    .Y(_0553_));
 sg13g2_a21oi_1 _2345_ (.A1(net276),
    .A2(_0552_),
    .Y(_0181_),
    .B1(_0553_));
 sg13g2_a22oi_1 _2346_ (.Y(_0554_),
    .B1(net286),
    .B2(net301),
    .A2(net331),
    .A1(net300));
 sg13g2_nor2_1 _2347_ (.A(net177),
    .B(net276),
    .Y(_0555_));
 sg13g2_a21oi_1 _2348_ (.A1(net276),
    .A2(_0554_),
    .Y(_0182_),
    .B1(_0555_));
 sg13g2_o21ai_1 _2349_ (.B1(net348),
    .Y(_0556_),
    .A1(\inst_calculator.state[5] ),
    .A2(net174));
 sg13g2_and2_1 _2350_ (.A(net347),
    .B(_0016_),
    .X(_0557_));
 sg13g2_o21ai_1 _2351_ (.B1(net175),
    .Y(_0183_),
    .A1(_0559_),
    .A2(_0557_));
 sg13g2_o21ai_1 _2352_ (.B1(net347),
    .Y(_0558_),
    .A1(net187),
    .A2(\inst_calculator.state[5] ));
 sg13g2_o21ai_1 _2353_ (.B1(net188),
    .Y(_0184_),
    .A1(_0560_),
    .A2(_0557_));
 sg13g2_dfrbp_1 _2354_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net27),
    .D(_0069_),
    .Q_N(_1187_),
    .Q(\inst_calculator.reg_arg[0] ));
 sg13g2_dfrbp_1 _2355_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net60),
    .D(_0070_),
    .Q_N(_1186_),
    .Q(\inst_calculator.reg_arg[1] ));
 sg13g2_dfrbp_1 _2356_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net58),
    .D(_0071_),
    .Q_N(_1185_),
    .Q(\inst_calculator.reg_arg[2] ));
 sg13g2_dfrbp_1 _2357_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net56),
    .D(_0072_),
    .Q_N(_1184_),
    .Q(\inst_calculator.reg_arg[3] ));
 sg13g2_dfrbp_1 _2358_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net54),
    .D(_0073_),
    .Q_N(_1183_),
    .Q(\inst_calculator.reg_arg[4] ));
 sg13g2_dfrbp_1 _2359_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net52),
    .D(_0074_),
    .Q_N(_1182_),
    .Q(\inst_calculator.reg_arg[5] ));
 sg13g2_dfrbp_1 _2360_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net50),
    .D(_0075_),
    .Q_N(_1181_),
    .Q(\inst_calculator.reg_arg[6] ));
 sg13g2_dfrbp_1 _2361_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net48),
    .D(_0076_),
    .Q_N(_1180_),
    .Q(\inst_calculator.reg_arg[7] ));
 sg13g2_dfrbp_1 _2362_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net46),
    .D(_0077_),
    .Q_N(_1179_),
    .Q(\inst_calculator.reg_arg[8] ));
 sg13g2_dfrbp_1 _2363_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net44),
    .D(_0078_),
    .Q_N(_1178_),
    .Q(\inst_calculator.reg_arg[9] ));
 sg13g2_dfrbp_1 _2364_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net42),
    .D(_0079_),
    .Q_N(_0055_),
    .Q(\inst_calculator.inst_keypad_poller.clk_counter[0] ));
 sg13g2_dfrbp_1 _2365_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net40),
    .D(net201),
    .Q_N(_1177_),
    .Q(\inst_calculator.inst_keypad_poller.clk_counter[1] ));
 sg13g2_dfrbp_1 _2366_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net38),
    .D(_0081_),
    .Q_N(_1176_),
    .Q(\inst_calculator.inst_keypad_poller.clk_counter[2] ));
 sg13g2_dfrbp_1 _2367_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net36),
    .D(_0082_),
    .Q_N(_1175_),
    .Q(\inst_calculator.inst_keypad_poller.clk_counter[3] ));
 sg13g2_dfrbp_1 _2368_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net35),
    .D(net241),
    .Q_N(_1174_),
    .Q(\inst_calculator.inst_keypad_poller.clk_counter[4] ));
 sg13g2_dfrbp_1 _2369_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net33),
    .D(_0084_),
    .Q_N(_1173_),
    .Q(\inst_calculator.inst_keypad_poller.clk_counter[5] ));
 sg13g2_dfrbp_1 _2370_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net31),
    .D(net213),
    .Q_N(_1172_),
    .Q(\inst_calculator.inst_keypad_poller.clk_counter[6] ));
 sg13g2_dfrbp_1 _2371_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net29),
    .D(_0086_),
    .Q_N(_1171_),
    .Q(\inst_calculator.inst_keypad_poller.clk_counter[7] ));
 sg13g2_dfrbp_1 _2372_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net26),
    .D(_0087_),
    .Q_N(_1170_),
    .Q(\inst_calculator.inst_keypad_poller.clk_counter[8] ));
 sg13g2_dfrbp_1 _2373_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net24),
    .D(_0088_),
    .Q_N(_1169_),
    .Q(\inst_calculator.inst_keypad_poller.clk_counter[9] ));
 sg13g2_dfrbp_1 _2374_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net22),
    .D(net371),
    .Q_N(_1168_),
    .Q(\inst_calculator.inst_keypad_poller.clk_counter[10] ));
 sg13g2_dfrbp_1 _2375_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net20),
    .D(_0090_),
    .Q_N(_1167_),
    .Q(\inst_calculator.inst_keypad_poller.clk_counter[11] ));
 sg13g2_dfrbp_1 _2376_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net18),
    .D(_0091_),
    .Q_N(_1166_),
    .Q(\inst_calculator.inst_keypad_poller.clk_counter[12] ));
 sg13g2_dfrbp_1 _2377_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net16),
    .D(net394),
    .Q_N(_1165_),
    .Q(\inst_calculator.inst_keypad_poller.clk_counter[13] ));
 sg13g2_dfrbp_1 _2378_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net14),
    .D(_0093_),
    .Q_N(_1164_),
    .Q(\inst_calculator.inst_keypad_poller.clk_counter[14] ));
 sg13g2_dfrbp_1 _2379_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net12),
    .D(_0094_),
    .Q_N(_1163_),
    .Q(\inst_calculator.inst_keypad_poller.clk_counter[15] ));
 sg13g2_dfrbp_1 _2380_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net10),
    .D(_0095_),
    .Q_N(_1162_),
    .Q(\inst_calculator.inst_keypad_poller.clk_counter[16] ));
 sg13g2_dfrbp_1 _2381_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net349),
    .D(_0063_),
    .Q_N(\inst_calculator.inst_keypad_poller.state[0] ),
    .Q(_0056_));
 sg13g2_dfrbp_1 _2382_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net353),
    .D(net180),
    .Q_N(_1188_),
    .Q(\inst_calculator.inst_keypad_poller.state[1] ));
 sg13g2_dfrbp_1 _2383_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net353),
    .D(net264),
    .Q_N(_1189_),
    .Q(\inst_calculator.inst_keypad_poller.state[2] ));
 sg13g2_dfrbp_1 _2384_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net350),
    .D(net103),
    .Q_N(_1190_),
    .Q(\inst_calculator.inst_keypad_poller.state[3] ));
 sg13g2_dfrbp_1 _2385_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net353),
    .D(net157),
    .Q_N(_0047_),
    .Q(\inst_calculator.inst_keypad_poller.state[4] ));
 sg13g2_dfrbp_1 _2386_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net352),
    .D(net161),
    .Q_N(_0048_),
    .Q(\inst_calculator.inst_keypad_poller.state[5] ));
 sg13g2_dfrbp_1 _2387_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net340),
    .D(_0052_),
    .Q_N(_1161_),
    .Q(\inst_calculator.inst_drive.flag ));
 sg13g2_dfrbp_1 _2388_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net340),
    .D(_0064_),
    .Q_N(uio_out[1]),
    .Q(_0057_));
 sg13g2_dfrbp_1 _2389_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net337),
    .D(_0065_),
    .Q_N(uio_out[2]),
    .Q(_0058_));
 sg13g2_dfrbp_1 _2390_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net340),
    .D(_0066_),
    .Q_N(uio_out[3]),
    .Q(_0059_));
 sg13g2_dfrbp_1 _2391_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net337),
    .D(_0185_),
    .Q_N(_1191_),
    .Q(\inst_calculator.inst_drive.num_disp[0] ));
 sg13g2_dfrbp_1 _2392_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net337),
    .D(net167),
    .Q_N(_0050_),
    .Q(\inst_calculator.inst_drive.num_disp[1] ));
 sg13g2_dfrbp_1 _2393_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net337),
    .D(_0187_),
    .Q_N(_0049_),
    .Q(\inst_calculator.inst_drive.num_disp[2] ));
 sg13g2_dfrbp_1 _2394_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net340),
    .D(_0188_),
    .Q_N(_1192_),
    .Q(\inst_calculator.inst_drive.num_disp[3] ));
 sg13g2_dfrbp_1 _2395_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net336),
    .D(_0022_),
    .Q_N(_1193_),
    .Q(\inst_calculator.inst_drive.cnt0[0] ));
 sg13g2_dfrbp_1 _2396_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net336),
    .D(_0027_),
    .Q_N(_1194_),
    .Q(\inst_calculator.inst_drive.cnt0[1] ));
 sg13g2_dfrbp_1 _2397_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net336),
    .D(net131),
    .Q_N(_1195_),
    .Q(\inst_calculator.inst_drive.cnt0[2] ));
 sg13g2_dfrbp_1 _2398_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net334),
    .D(_0029_),
    .Q_N(_1196_),
    .Q(\inst_calculator.inst_drive.cnt0[3] ));
 sg13g2_dfrbp_1 _2399_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net334),
    .D(_0030_),
    .Q_N(_1197_),
    .Q(\inst_calculator.inst_drive.cnt0[4] ));
 sg13g2_dfrbp_1 _2400_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net335),
    .D(_0031_),
    .Q_N(_1198_),
    .Q(\inst_calculator.inst_drive.cnt0[5] ));
 sg13g2_dfrbp_1 _2401_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net335),
    .D(net170),
    .Q_N(_1199_),
    .Q(\inst_calculator.inst_drive.cnt0[6] ));
 sg13g2_dfrbp_1 _2402_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net334),
    .D(_0033_),
    .Q_N(_1200_),
    .Q(\inst_calculator.inst_drive.cnt0[7] ));
 sg13g2_dfrbp_1 _2403_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net334),
    .D(net222),
    .Q_N(_1201_),
    .Q(\inst_calculator.inst_drive.cnt0[8] ));
 sg13g2_dfrbp_1 _2404_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net334),
    .D(_0035_),
    .Q_N(_1202_),
    .Q(\inst_calculator.inst_drive.cnt0[9] ));
 sg13g2_dfrbp_1 _2405_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net334),
    .D(_0023_),
    .Q_N(_1203_),
    .Q(\inst_calculator.inst_drive.cnt0[10] ));
 sg13g2_dfrbp_1 _2406_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net334),
    .D(_0024_),
    .Q_N(_0051_),
    .Q(\inst_calculator.inst_drive.cnt0[11] ));
 sg13g2_dfrbp_1 _2407_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net334),
    .D(net199),
    .Q_N(_1204_),
    .Q(\inst_calculator.inst_drive.cnt0[12] ));
 sg13g2_dfrbp_1 _2408_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net335),
    .D(net387),
    .Q_N(_1160_),
    .Q(\inst_calculator.inst_drive.cnt0[13] ));
 sg13g2_dfrbp_1 _2409_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net342),
    .D(net101),
    .Q_N(_0054_),
    .Q(\inst_calculator.inst_divider.q[0] ));
 sg13g2_dfrbp_1 _2410_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net342),
    .D(_0097_),
    .Q_N(_1159_),
    .Q(\inst_calculator.inst_divider.q[1] ));
 sg13g2_dfrbp_1 _2411_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net342),
    .D(net210),
    .Q_N(_1158_),
    .Q(\inst_calculator.inst_divider.q[2] ));
 sg13g2_dfrbp_1 _2412_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net341),
    .D(net185),
    .Q_N(_1157_),
    .Q(\inst_calculator.inst_divider.q[3] ));
 sg13g2_dfrbp_1 _2413_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net341),
    .D(net159),
    .Q_N(_1156_),
    .Q(\inst_calculator.inst_divider.q[4] ));
 sg13g2_dfrbp_1 _2414_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net342),
    .D(_0101_),
    .Q_N(_1155_),
    .Q(\inst_calculator.inst_divider.q[5] ));
 sg13g2_dfrbp_1 _2415_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net342),
    .D(net155),
    .Q_N(_1154_),
    .Q(\inst_calculator.inst_divider.q[6] ));
 sg13g2_dfrbp_1 _2416_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net342),
    .D(_0103_),
    .Q_N(_1153_),
    .Q(\inst_calculator.inst_divider.q[7] ));
 sg13g2_dfrbp_1 _2417_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net342),
    .D(_0104_),
    .Q_N(_1152_),
    .Q(\inst_calculator.inst_divider.q[8] ));
 sg13g2_dfrbp_1 _2418_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net342),
    .D(net149),
    .Q_N(_1205_),
    .Q(\inst_calculator.inst_divider.q[9] ));
 sg13g2_dfrbp_1 _2419_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net349),
    .D(net443),
    .Q_N(_1206_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _2420_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net349),
    .D(net427),
    .Q_N(_1207_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _2421_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net349),
    .D(net109),
    .Q_N(_1208_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _2422_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net338),
    .D(_0003_),
    .Q_N(_1209_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _2423_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net338),
    .D(net106),
    .Q_N(_1210_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _2424_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net338),
    .D(net419),
    .Q_N(_1151_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _2425_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net338),
    .D(net91),
    .Q_N(uo_out[6]),
    .Q(_0060_));
 sg13g2_dfrbp_1 _2426_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net78),
    .D(_0106_),
    .Q_N(_1150_),
    .Q(\inst_calculator.inst_divider.busy ));
 sg13g2_dfrbp_1 _2427_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net76),
    .D(_0107_),
    .Q_N(_1149_),
    .Q(\inst_calculator.denominator[0] ));
 sg13g2_dfrbp_1 _2428_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net75),
    .D(_0108_),
    .Q_N(_1148_),
    .Q(\inst_calculator.denominator[1] ));
 sg13g2_dfrbp_1 _2429_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net74),
    .D(_0109_),
    .Q_N(_1147_),
    .Q(\inst_calculator.denominator[2] ));
 sg13g2_dfrbp_1 _2430_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net73),
    .D(net125),
    .Q_N(_1146_),
    .Q(\inst_calculator.denominator[3] ));
 sg13g2_dfrbp_1 _2431_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net72),
    .D(_0111_),
    .Q_N(_1145_),
    .Q(\inst_calculator.denominator[4] ));
 sg13g2_dfrbp_1 _2432_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net71),
    .D(net113),
    .Q_N(_1144_),
    .Q(\inst_calculator.denominator[5] ));
 sg13g2_dfrbp_1 _2433_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net70),
    .D(net116),
    .Q_N(_1143_),
    .Q(\inst_calculator.denominator[6] ));
 sg13g2_dfrbp_1 _2434_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net69),
    .D(net141),
    .Q_N(_1142_),
    .Q(\inst_calculator.denominator[7] ));
 sg13g2_dfrbp_1 _2435_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net68),
    .D(_0115_),
    .Q_N(_1141_),
    .Q(\inst_calculator.denominator[8] ));
 sg13g2_dfrbp_1 _2436_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net67),
    .D(net260),
    .Q_N(_1140_),
    .Q(\inst_calculator.denominator[9] ));
 sg13g2_dfrbp_1 _2437_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net352),
    .D(net97),
    .Q_N(_1139_),
    .Q(\inst_calculator.divider_done ));
 sg13g2_dfrbp_1 _2438_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net344),
    .D(net246),
    .Q_N(_1138_),
    .Q(\inst_calculator.inst_divider.d[0] ));
 sg13g2_dfrbp_1 _2439_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net344),
    .D(net229),
    .Q_N(_1137_),
    .Q(\inst_calculator.inst_divider.d[1] ));
 sg13g2_dfrbp_1 _2440_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net345),
    .D(net238),
    .Q_N(_1136_),
    .Q(\inst_calculator.inst_divider.d[2] ));
 sg13g2_dfrbp_1 _2441_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net344),
    .D(_0121_),
    .Q_N(_1135_),
    .Q(\inst_calculator.inst_divider.d[3] ));
 sg13g2_dfrbp_1 _2442_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net344),
    .D(_0122_),
    .Q_N(_1134_),
    .Q(\inst_calculator.inst_divider.d[4] ));
 sg13g2_dfrbp_1 _2443_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net346),
    .D(_0123_),
    .Q_N(_1133_),
    .Q(\inst_calculator.inst_divider.d[5] ));
 sg13g2_dfrbp_1 _2444_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net345),
    .D(_0124_),
    .Q_N(_1132_),
    .Q(\inst_calculator.inst_divider.d[6] ));
 sg13g2_dfrbp_1 _2445_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net345),
    .D(_0125_),
    .Q_N(_1131_),
    .Q(\inst_calculator.inst_divider.d[7] ));
 sg13g2_dfrbp_1 _2446_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net352),
    .D(net236),
    .Q_N(_1130_),
    .Q(\inst_calculator.inst_divider.d[8] ));
 sg13g2_dfrbp_1 _2447_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net352),
    .D(net219),
    .Q_N(_1129_),
    .Q(\inst_calculator.inst_divider.d[9] ));
 sg13g2_dfrbp_1 _2448_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net344),
    .D(net144),
    .Q_N(_1128_),
    .Q(\inst_calculator.inst_divider.n[0] ));
 sg13g2_dfrbp_1 _2449_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net344),
    .D(net215),
    .Q_N(_1127_),
    .Q(\inst_calculator.inst_divider.n[1] ));
 sg13g2_dfrbp_1 _2450_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net344),
    .D(net378),
    .Q_N(_1126_),
    .Q(\inst_calculator.inst_divider.n[2] ));
 sg13g2_dfrbp_1 _2451_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net344),
    .D(net258),
    .Q_N(_1125_),
    .Q(\inst_calculator.inst_divider.n[3] ));
 sg13g2_dfrbp_1 _2452_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net345),
    .D(net250),
    .Q_N(_1124_),
    .Q(\inst_calculator.inst_divider.n[4] ));
 sg13g2_dfrbp_1 _2453_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net345),
    .D(_0133_),
    .Q_N(_1123_),
    .Q(\inst_calculator.inst_divider.n[5] ));
 sg13g2_dfrbp_1 _2454_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net345),
    .D(net262),
    .Q_N(_1122_),
    .Q(\inst_calculator.inst_divider.n[6] ));
 sg13g2_dfrbp_1 _2455_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net345),
    .D(net374),
    .Q_N(_1121_),
    .Q(\inst_calculator.inst_divider.n[7] ));
 sg13g2_dfrbp_1 _2456_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net352),
    .D(net400),
    .Q_N(_1120_),
    .Q(\inst_calculator.inst_divider.n[8] ));
 sg13g2_dfrbp_1 _2457_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net352),
    .D(net227),
    .Q_N(_1211_),
    .Q(\inst_calculator.inst_divider.n[9] ));
 sg13g2_dfrbp_1 _2458_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net349),
    .D(_0189_),
    .Q_N(_1212_),
    .Q(\inst_calculator.inst_keypad_encoder.key[0] ));
 sg13g2_dfrbp_1 _2459_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net349),
    .D(_0190_),
    .Q_N(_1213_),
    .Q(\inst_calculator.inst_keypad_encoder.key[1] ));
 sg13g2_dfrbp_1 _2460_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net349),
    .D(_0191_),
    .Q_N(_1214_),
    .Q(\inst_calculator.inst_keypad_encoder.key[2] ));
 sg13g2_dfrbp_1 _2461_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net337),
    .D(_0192_),
    .Q_N(_0045_),
    .Q(\inst_calculator.inst_keypad_encoder.key[3] ));
 sg13g2_dfrbp_1 _2462_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net353),
    .D(_0138_),
    .Q_N(_1119_),
    .Q(\inst_calculator.inst_keypad_encoder.rows[0] ));
 sg13g2_dfrbp_1 _2463_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net350),
    .D(_0139_),
    .Q_N(_1118_),
    .Q(\inst_calculator.inst_keypad_encoder.rows[1] ));
 sg13g2_dfrbp_1 _2464_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net353),
    .D(_0140_),
    .Q_N(_1117_),
    .Q(\inst_calculator.inst_keypad_encoder.rows[2] ));
 sg13g2_dfrbp_1 _2465_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net350),
    .D(_0141_),
    .Q_N(_1116_),
    .Q(\inst_calculator.inst_keypad_encoder.rows[3] ));
 sg13g2_dfrbp_1 _2466_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net340),
    .D(_0142_),
    .Q_N(_1115_),
    .Q(\inst_calculator.inst_drive.cnt_sel[0] ));
 sg13g2_dfrbp_1 _2467_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net340),
    .D(net118),
    .Q_N(_1114_),
    .Q(\inst_calculator.inst_drive.cnt_sel[1] ));
 sg13g2_dfrbp_1 _2468_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net338),
    .D(net99),
    .Q_N(uio_out[4]),
    .Q(_0061_));
 sg13g2_dfrbp_1 _2469_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net337),
    .D(_0145_),
    .Q_N(_1113_),
    .Q(uio_out[5]));
 sg13g2_dfrbp_1 _2470_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net337),
    .D(_0146_),
    .Q_N(_1112_),
    .Q(uio_out[6]));
 sg13g2_dfrbp_1 _2471_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net338),
    .D(net422),
    .Q_N(_0053_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _2472_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net350),
    .D(_0148_),
    .Q_N(_1111_),
    .Q(\inst_calculator.inst_keypad_poller.key_pressed ));
 sg13g2_dfrbp_1 _2473_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net64),
    .D(net121),
    .Q_N(_1110_),
    .Q(\inst_calculator.key_pressed_prev ));
 sg13g2_dfrbp_1 _2474_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net63),
    .D(net93),
    .Q_N(_0020_),
    .Q(\inst_calculator.divider_start ));
 sg13g2_dfrbp_1 _2475_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net62),
    .D(_0151_),
    .Q_N(_1109_),
    .Q(\inst_calculator.reg_operator[0] ));
 sg13g2_dfrbp_1 _2476_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net59),
    .D(_0152_),
    .Q_N(_1108_),
    .Q(\inst_calculator.reg_operator[1] ));
 sg13g2_dfrbp_1 _2477_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net55),
    .D(net137),
    .Q_N(_1107_),
    .Q(\inst_calculator.inst_divider.numerator[0] ));
 sg13g2_dfrbp_1 _2478_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net53),
    .D(net139),
    .Q_N(_1106_),
    .Q(\inst_calculator.inst_divider.numerator[1] ));
 sg13g2_dfrbp_1 _2479_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net51),
    .D(net123),
    .Q_N(_1105_),
    .Q(\inst_calculator.inst_divider.numerator[2] ));
 sg13g2_dfrbp_1 _2480_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net49),
    .D(net133),
    .Q_N(_1104_),
    .Q(\inst_calculator.inst_divider.numerator[3] ));
 sg13g2_dfrbp_1 _2481_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net47),
    .D(net147),
    .Q_N(_1103_),
    .Q(\inst_calculator.inst_divider.numerator[4] ));
 sg13g2_dfrbp_1 _2482_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net45),
    .D(net127),
    .Q_N(_1102_),
    .Q(\inst_calculator.inst_divider.numerator[5] ));
 sg13g2_dfrbp_1 _2483_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net43),
    .D(net217),
    .Q_N(_1101_),
    .Q(\inst_calculator.inst_divider.numerator[6] ));
 sg13g2_dfrbp_1 _2484_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net41),
    .D(net224),
    .Q_N(_1100_),
    .Q(\inst_calculator.inst_divider.numerator[7] ));
 sg13g2_dfrbp_1 _2485_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net39),
    .D(net361),
    .Q_N(_1099_),
    .Q(\inst_calculator.inst_divider.numerator[8] ));
 sg13g2_dfrbp_1 _2486_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net37),
    .D(net256),
    .Q_N(_1098_),
    .Q(\inst_calculator.inst_divider.numerator[9] ));
 sg13g2_dfrbp_1 _2487_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net347),
    .D(_0068_),
    .Q_N(\inst_calculator.state[0] ),
    .Q(_0062_));
 sg13g2_dfrbp_1 _2488_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net343),
    .D(net411),
    .Q_N(_0021_),
    .Q(\inst_calculator.state[1] ));
 sg13g2_dfrbp_1 _2489_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net347),
    .D(_0008_),
    .Q_N(_1215_),
    .Q(\inst_calculator.state[2] ));
 sg13g2_dfrbp_1 _2490_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net339),
    .D(_0009_),
    .Q_N(_1216_),
    .Q(\inst_calculator.state[3] ));
 sg13g2_dfrbp_1 _2491_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net343),
    .D(net415),
    .Q_N(_1217_),
    .Q(\inst_calculator.state[4] ));
 sg13g2_dfrbp_1 _2492_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net347),
    .D(_0010_),
    .Q_N(_1218_),
    .Q(\inst_calculator.state[5] ));
 sg13g2_dfrbp_1 _2493_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net337),
    .D(net173),
    .Q_N(_1219_),
    .Q(\inst_calculator.state[6] ));
 sg13g2_dfrbp_1 _2494_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net339),
    .D(net89),
    .Q_N(_1220_),
    .Q(\inst_calculator.state[7] ));
 sg13g2_dfrbp_1 _2495_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net347),
    .D(net191),
    .Q_N(_1221_),
    .Q(\inst_calculator.state[8] ));
 sg13g2_dfrbp_1 _2496_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net347),
    .D(net111),
    .Q_N(_1222_),
    .Q(\inst_calculator.state[9] ));
 sg13g2_dfrbp_1 _2497_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net348),
    .D(net391),
    .Q_N(_0046_),
    .Q(\inst_calculator.state[10] ));
 sg13g2_dfrbp_1 _2498_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net32),
    .D(_0163_),
    .Q_N(_1097_),
    .Q(\inst_calculator.reg_result[9] ));
 sg13g2_dfrbp_1 _2499_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net28),
    .D(net385),
    .Q_N(_1096_),
    .Q(\inst_calculator.reg_result[8] ));
 sg13g2_dfrbp_1 _2500_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net23),
    .D(_0165_),
    .Q_N(_1095_),
    .Q(\inst_calculator.reg_result[7] ));
 sg13g2_dfrbp_1 _2501_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net19),
    .D(_0166_),
    .Q_N(_1094_),
    .Q(\inst_calculator.reg_result[6] ));
 sg13g2_dfrbp_1 _2502_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net15),
    .D(_0167_),
    .Q_N(_1093_),
    .Q(\inst_calculator.reg_result[5] ));
 sg13g2_dfrbp_1 _2503_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net11),
    .D(_0168_),
    .Q_N(_1092_),
    .Q(\inst_calculator.reg_result[4] ));
 sg13g2_dfrbp_1 _2504_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net8),
    .D(_0169_),
    .Q_N(_1091_),
    .Q(\inst_calculator.reg_result[3] ));
 sg13g2_dfrbp_1 _2505_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net7),
    .D(net440),
    .Q_N(_1090_),
    .Q(\inst_calculator.reg_result[2] ));
 sg13g2_dfrbp_1 _2506_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net79),
    .D(net431),
    .Q_N(_1089_),
    .Q(\inst_calculator.reg_result[1] ));
 sg13g2_dfrbp_1 _2507_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net66),
    .D(net437),
    .Q_N(_1088_),
    .Q(\inst_calculator.reg_result[0] ));
 sg13g2_dfrbp_1 _2508_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net61),
    .D(net252),
    .Q_N(_0037_),
    .Q(\inst_calculator.inst_bin2bcd.bin_in[9] ));
 sg13g2_dfrbp_1 _2509_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net34),
    .D(net429),
    .Q_N(_0038_),
    .Q(\inst_calculator.inst_bin2bcd.bin_in[8] ));
 sg13g2_dfrbp_1 _2510_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net25),
    .D(net435),
    .Q_N(_0036_),
    .Q(\inst_calculator.inst_bin2bcd.bin_in[7] ));
 sg13g2_dfrbp_1 _2511_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net17),
    .D(net231),
    .Q_N(_0039_),
    .Q(\inst_calculator.inst_bin2bcd.bin_in[6] ));
 sg13g2_dfrbp_1 _2512_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net9),
    .D(net376),
    .Q_N(_0040_),
    .Q(\inst_calculator.inst_bin2bcd.bin_in[5] ));
 sg13g2_dfrbp_1 _2513_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net6),
    .D(net194),
    .Q_N(_0041_),
    .Q(\inst_calculator.inst_bin2bcd.bin_in[4] ));
 sg13g2_dfrbp_1 _2514_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net65),
    .D(_0179_),
    .Q_N(_0042_),
    .Q(\inst_calculator.inst_bin2bcd.bin_in[3] ));
 sg13g2_dfrbp_1 _2515_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net30),
    .D(_0180_),
    .Q_N(_0043_),
    .Q(\inst_calculator.inst_bin2bcd.bin_in[2] ));
 sg13g2_dfrbp_1 _2516_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net13),
    .D(_0181_),
    .Q_N(_0044_),
    .Q(\inst_calculator.inst_bin2bcd.bin_in[1] ));
 sg13g2_dfrbp_1 _2517_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net77),
    .D(_0182_),
    .Q_N(_1087_),
    .Q(\inst_calculator.bcd[0] ));
 sg13g2_dfrbp_1 _2518_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net21),
    .D(net176),
    .Q_N(_1086_),
    .Q(\inst_calculator.reg_operator_next[1] ));
 sg13g2_dfrbp_1 _2519_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net57),
    .D(net189),
    .Q_N(_1085_),
    .Q(\inst_calculator.reg_operator_next[0] ));
 sg13g2_tiehi _2505__7 (.L_HI(net7));
 sg13g2_tiehi _2504__8 (.L_HI(net8));
 sg13g2_tiehi _2512__9 (.L_HI(net9));
 sg13g2_tiehi _2380__10 (.L_HI(net10));
 sg13g2_tiehi _2503__11 (.L_HI(net11));
 sg13g2_tiehi _2379__12 (.L_HI(net12));
 sg13g2_tiehi _2516__13 (.L_HI(net13));
 sg13g2_tiehi _2378__14 (.L_HI(net14));
 sg13g2_tiehi _2502__15 (.L_HI(net15));
 sg13g2_tiehi _2377__16 (.L_HI(net16));
 sg13g2_tiehi _2511__17 (.L_HI(net17));
 sg13g2_tiehi _2376__18 (.L_HI(net18));
 sg13g2_tiehi _2501__19 (.L_HI(net19));
 sg13g2_tiehi _2375__20 (.L_HI(net20));
 sg13g2_tiehi _2518__21 (.L_HI(net21));
 sg13g2_tiehi _2374__22 (.L_HI(net22));
 sg13g2_tiehi _2500__23 (.L_HI(net23));
 sg13g2_tiehi _2373__24 (.L_HI(net24));
 sg13g2_tiehi _2510__25 (.L_HI(net25));
 sg13g2_tiehi _2372__26 (.L_HI(net26));
 sg13g2_tiehi _2354__27 (.L_HI(net27));
 sg13g2_tiehi _2499__28 (.L_HI(net28));
 sg13g2_tiehi _2371__29 (.L_HI(net29));
 sg13g2_tiehi _2515__30 (.L_HI(net30));
 sg13g2_tiehi _2370__31 (.L_HI(net31));
 sg13g2_tiehi _2498__32 (.L_HI(net32));
 sg13g2_tiehi _2369__33 (.L_HI(net33));
 sg13g2_tiehi _2509__34 (.L_HI(net34));
 sg13g2_tiehi _2368__35 (.L_HI(net35));
 sg13g2_tiehi _2367__36 (.L_HI(net36));
 sg13g2_tiehi _2486__37 (.L_HI(net37));
 sg13g2_tiehi _2366__38 (.L_HI(net38));
 sg13g2_tiehi _2485__39 (.L_HI(net39));
 sg13g2_tiehi _2365__40 (.L_HI(net40));
 sg13g2_tiehi _2484__41 (.L_HI(net41));
 sg13g2_tiehi _2364__42 (.L_HI(net42));
 sg13g2_tiehi _2483__43 (.L_HI(net43));
 sg13g2_tiehi _2363__44 (.L_HI(net44));
 sg13g2_tiehi _2482__45 (.L_HI(net45));
 sg13g2_tiehi _2362__46 (.L_HI(net46));
 sg13g2_tiehi _2481__47 (.L_HI(net47));
 sg13g2_tiehi _2361__48 (.L_HI(net48));
 sg13g2_tiehi _2480__49 (.L_HI(net49));
 sg13g2_tiehi _2360__50 (.L_HI(net50));
 sg13g2_tiehi _2479__51 (.L_HI(net51));
 sg13g2_tiehi _2359__52 (.L_HI(net52));
 sg13g2_tiehi _2478__53 (.L_HI(net53));
 sg13g2_tiehi _2358__54 (.L_HI(net54));
 sg13g2_tiehi _2477__55 (.L_HI(net55));
 sg13g2_tiehi _2357__56 (.L_HI(net56));
 sg13g2_tiehi _2519__57 (.L_HI(net57));
 sg13g2_tiehi _2356__58 (.L_HI(net58));
 sg13g2_tiehi _2476__59 (.L_HI(net59));
 sg13g2_tiehi _2355__60 (.L_HI(net60));
 sg13g2_tiehi _2508__61 (.L_HI(net61));
 sg13g2_tiehi _2475__62 (.L_HI(net62));
 sg13g2_tiehi _2474__63 (.L_HI(net63));
 sg13g2_tiehi _2473__64 (.L_HI(net64));
 sg13g2_tiehi _2514__65 (.L_HI(net65));
 sg13g2_tiehi _2507__66 (.L_HI(net66));
 sg13g2_tiehi _2436__67 (.L_HI(net67));
 sg13g2_tiehi _2435__68 (.L_HI(net68));
 sg13g2_tiehi _2434__69 (.L_HI(net69));
 sg13g2_tiehi _2433__70 (.L_HI(net70));
 sg13g2_tiehi _2432__71 (.L_HI(net71));
 sg13g2_tiehi _2431__72 (.L_HI(net72));
 sg13g2_tiehi _2430__73 (.L_HI(net73));
 sg13g2_tiehi _2429__74 (.L_HI(net74));
 sg13g2_tiehi _2428__75 (.L_HI(net75));
 sg13g2_tiehi _2427__76 (.L_HI(net76));
 sg13g2_tiehi _2517__77 (.L_HI(net77));
 sg13g2_tiehi _2426__78 (.L_HI(net78));
 sg13g2_tiehi _2506__79 (.L_HI(net79));
 sg13g2_tiehi tt_um_shuangyu_top_80 (.L_HI(net80));
 sg13g2_tiehi tt_um_shuangyu_top_81 (.L_HI(net81));
 sg13g2_tiehi tt_um_shuangyu_top_82 (.L_HI(net82));
 sg13g2_tiehi tt_um_shuangyu_top_83 (.L_HI(net83));
 sg13g2_tiehi tt_um_shuangyu_top_84 (.L_HI(net84));
 sg13g2_tiehi tt_um_shuangyu_top_85 (.L_HI(net85));
 sg13g2_tiehi tt_um_shuangyu_top_86 (.L_HI(net86));
 sg13g2_tiehi tt_um_shuangyu_top_87 (.L_HI(net87));
 sg13g2_tiehi tt_um_shuangyu_top_88 (.L_HI(net88));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _2513__6 (.L_HI(net6));
 sg13g2_buf_4 fanout265 (.X(net265),
    .A(_1051_));
 sg13g2_buf_2 fanout266 (.A(net267),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_0052_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_0900_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(net270),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_0980_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_0899_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(net273),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(net274),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_0466_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(net277),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(net277),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_0535_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_0459_),
    .X(net278));
 sg13g2_buf_4 fanout279 (.X(net279),
    .A(_0201_));
 sg13g2_buf_2 fanout280 (.A(net281),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(net285),
    .X(net281));
 sg13g2_buf_1 fanout282 (.A(net285),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(net285),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(net285),
    .X(net284));
 sg13g2_buf_1 fanout285 (.A(_1053_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(net287),
    .X(net286));
 sg13g2_buf_4 fanout287 (.X(net287),
    .A(\inst_calculator.reg_result[0] ));
 sg13g2_buf_2 fanout288 (.A(net289),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(\inst_calculator.reg_result[1] ),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(net291),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(net439),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(\inst_calculator.reg_result[3] ),
    .X(net292));
 sg13g2_buf_4 fanout293 (.X(net293),
    .A(\inst_calculator.reg_result[4] ));
 sg13g2_buf_4 fanout294 (.X(net294),
    .A(\inst_calculator.reg_result[5] ));
 sg13g2_buf_4 fanout295 (.X(net295),
    .A(net417));
 sg13g2_buf_4 fanout296 (.X(net296),
    .A(net432));
 sg13g2_buf_2 fanout297 (.A(net299),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(net299),
    .X(net298));
 sg13g2_buf_1 fanout299 (.A(\inst_calculator.state[10] ),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(\inst_calculator.state[7] ),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(\inst_calculator.state[4] ),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(net303),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(net414),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(net305),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(\inst_calculator.reg_operator[1] ),
    .X(net305));
 sg13g2_buf_4 fanout306 (.X(net306),
    .A(net307));
 sg13g2_buf_2 fanout307 (.A(\inst_calculator.divider_start ),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(net310),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(net310),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(\inst_calculator.divider_start ),
    .X(net310));
 sg13g2_buf_4 fanout311 (.X(net311),
    .A(net166));
 sg13g2_buf_2 fanout312 (.A(net110),
    .X(net312));
 sg13g2_buf_4 fanout313 (.X(net313),
    .A(net366));
 sg13g2_buf_4 fanout314 (.X(net314),
    .A(net449));
 sg13g2_buf_4 fanout315 (.X(net315),
    .A(net316));
 sg13g2_buf_2 fanout316 (.A(\inst_calculator.reg_arg[6] ),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(net318),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(net319),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(\inst_calculator.reg_arg[5] ),
    .X(net319));
 sg13g2_buf_4 fanout320 (.X(net320),
    .A(\inst_calculator.reg_arg[4] ));
 sg13g2_buf_2 fanout321 (.A(net448),
    .X(net321));
 sg13g2_buf_4 fanout322 (.X(net322),
    .A(net324));
 sg13g2_buf_2 fanout323 (.A(net324),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(\inst_calculator.reg_arg[3] ),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(net326),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(net327),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(net242),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(net330),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(net330),
    .X(net329));
 sg13g2_buf_4 fanout330 (.X(net330),
    .A(net253));
 sg13g2_buf_4 fanout331 (.X(net331),
    .A(\inst_calculator.reg_arg[0] ));
 sg13g2_buf_1 fanout332 (.A(\inst_calculator.reg_arg[0] ),
    .X(net332));
 sg13g2_buf_4 fanout333 (.X(net333),
    .A(net254));
 sg13g2_buf_4 fanout334 (.X(net334),
    .A(net335));
 sg13g2_buf_2 fanout335 (.A(net336),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(net341),
    .X(net336));
 sg13g2_buf_4 fanout337 (.X(net337),
    .A(net339));
 sg13g2_buf_4 fanout338 (.X(net338),
    .A(net339));
 sg13g2_buf_2 fanout339 (.A(net340),
    .X(net339));
 sg13g2_buf_4 fanout340 (.X(net340),
    .A(net341));
 sg13g2_buf_4 fanout341 (.X(net341),
    .A(rst_n));
 sg13g2_buf_4 fanout342 (.X(net342),
    .A(net346));
 sg13g2_buf_2 fanout343 (.A(net346),
    .X(net343));
 sg13g2_buf_4 fanout344 (.X(net344),
    .A(net345));
 sg13g2_buf_4 fanout345 (.X(net345),
    .A(net346));
 sg13g2_buf_2 fanout346 (.A(net354),
    .X(net346));
 sg13g2_buf_4 fanout347 (.X(net347),
    .A(net351));
 sg13g2_buf_1 fanout348 (.A(net351),
    .X(net348));
 sg13g2_buf_4 fanout349 (.X(net349),
    .A(net351));
 sg13g2_buf_2 fanout350 (.A(net351),
    .X(net350));
 sg13g2_buf_1 fanout351 (.A(net354),
    .X(net351));
 sg13g2_buf_4 fanout352 (.X(net352),
    .A(net354));
 sg13g2_buf_4 fanout353 (.X(net353),
    .A(net354));
 sg13g2_buf_2 fanout354 (.A(rst_n),
    .X(net354));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_tielo tt_um_shuangyu_top_5 (.L_LO(net5));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_25__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\inst_calculator.state[3] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0050_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0067_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0021_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0150_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0055_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0976_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0020_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0117_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0053_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0144_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0054_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0096_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold14 (.A(\inst_calculator.inst_keypad_poller.state[0] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0015_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0049_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0633_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0004_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold19 (.A(\inst_calculator.inst_keypad_poller.state[4] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold20 (.A(\inst_calculator.inst_drive.num_disp[1] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0002_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold22 (.A(\inst_calculator.inst_keypad_encoder.key[1] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0012_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold24 (.A(\inst_calculator.denominator[5] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0112_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold26 (.A(\inst_calculator.inst_drive.cnt0[0] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold27 (.A(\inst_calculator.denominator[6] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0113_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold29 (.A(\inst_calculator.inst_drive.flag ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0143_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold31 (.A(\inst_calculator.key_pressed_prev ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0200_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0149_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold34 (.A(\inst_calculator.inst_divider.numerator[2] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0155_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold36 (.A(\inst_calculator.denominator[3] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0110_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold38 (.A(\inst_calculator.inst_divider.numerator[5] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0158_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold40 (.A(\inst_calculator.denominator[4] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold41 (.A(\inst_calculator.inst_drive.cnt0[2] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0651_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0028_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold44 (.A(\inst_calculator.inst_divider.numerator[3] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0156_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold46 (.A(\inst_calculator.reg_operator_next[1] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0208_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold48 (.A(\inst_calculator.inst_divider.numerator[0] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0153_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold50 (.A(\inst_calculator.inst_divider.numerator[1] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0154_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold52 (.A(\inst_calculator.denominator[7] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0114_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold54 (.A(\inst_calculator.inst_divider.n[0] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold55 (.A(_1063_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0128_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold57 (.A(\inst_calculator.inst_keypad_poller.key_pressed ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold58 (.A(\inst_calculator.inst_divider.numerator[4] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0157_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold60 (.A(\inst_calculator.inst_divider.q[9] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0105_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold62 (.A(\inst_calculator.inst_divider.d[4] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold63 (.A(\inst_calculator.reg_operator_next[0] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0207_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold65 (.A(\inst_calculator.inst_divider.q[6] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold66 (.A(_1048_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0102_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold68 (.A(\inst_calculator.inst_keypad_poller.state[1] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0006_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold70 (.A(\inst_calculator.inst_divider.q[4] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0100_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold72 (.A(\inst_calculator.inst_keypad_poller.state[2] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0007_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold74 (.A(\inst_calculator.inst_divider.d[6] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold75 (.A(\inst_calculator.inst_keypad_poller.clk_counter[2] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0979_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold77 (.A(\inst_calculator.inst_divider.d[7] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold78 (.A(\inst_calculator.inst_drive.cnt_sel[0] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0186_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold80 (.A(\inst_calculator.inst_drive.cnt0[6] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0655_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0032_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold83 (.A(\inst_calculator.state[6] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0615_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0019_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold86 (.A(\inst_calculator.state[8] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0556_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0183_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold89 (.A(\inst_calculator.bcd[0] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0047_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0630_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0013_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold93 (.A(\inst_calculator.inst_bin2bcd.bin_in[2] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold94 (.A(\inst_calculator.inst_divider.q[5] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold95 (.A(\inst_calculator.inst_drive.cnt0[1] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold96 (.A(\inst_calculator.inst_divider.q[3] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0099_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold98 (.A(\inst_calculator.inst_drive.cnt0[3] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold99 (.A(\inst_calculator.state[2] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0558_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0184_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold102 (.A(\inst_calculator.inst_keypad_encoder.key[0] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0011_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold104 (.A(\inst_calculator.inst_bin2bcd.bin_in[3] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold105 (.A(\inst_calculator.inst_bin2bcd.bin_in[4] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0178_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold107 (.A(\inst_calculator.inst_keypad_encoder.rows[0] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold108 (.A(_1084_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold109 (.A(\inst_calculator.inst_drive.cnt0[12] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0667_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0025_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold112 (.A(\inst_calculator.inst_keypad_poller.clk_counter[1] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0080_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold114 (.A(\inst_calculator.inst_keypad_encoder.rows[3] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0195_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold116 (.A(\inst_calculator.inst_divider.d[3] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold117 (.A(\inst_calculator.inst_bin2bcd.bin_in[1] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold118 (.A(\inst_calculator.state[0] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0901_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold120 (.A(\inst_calculator.inst_divider.d[5] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold121 (.A(\inst_calculator.inst_divider.q[2] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0098_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold123 (.A(\inst_calculator.inst_keypad_poller.clk_counter[6] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0989_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0085_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold126 (.A(\inst_calculator.inst_divider.n[1] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0129_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold128 (.A(\inst_calculator.inst_divider.numerator[6] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0159_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold130 (.A(\inst_calculator.inst_divider.d[9] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0127_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold132 (.A(\inst_calculator.inst_drive.cnt0[8] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0660_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0034_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold135 (.A(\inst_calculator.inst_divider.numerator[7] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0160_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold137 (.A(\inst_calculator.inst_divider.n[9] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold138 (.A(_1082_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0137_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold140 (.A(\inst_calculator.denominator[1] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0119_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold142 (.A(\inst_calculator.inst_bin2bcd.bin_in[6] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0176_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold144 (.A(\inst_calculator.inst_keypad_poller.clk_counter[8] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0993_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold146 (.A(\inst_calculator.inst_divider.q[7] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold147 (.A(\inst_calculator.denominator[8] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0126_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold149 (.A(\inst_calculator.denominator[2] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0120_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold151 (.A(\inst_calculator.inst_keypad_poller.clk_counter[4] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0985_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0083_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold154 (.A(\inst_calculator.reg_arg[2] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold155 (.A(\inst_calculator.inst_keypad_poller.clk_counter[5] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold156 (.A(\inst_calculator.inst_divider.n[5] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold157 (.A(\inst_calculator.denominator[0] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0118_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold159 (.A(\inst_calculator.inst_keypad_poller.clk_counter[3] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0983_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold161 (.A(\inst_calculator.inst_divider.n[4] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0132_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold163 (.A(\inst_calculator.inst_bin2bcd.bin_in[9] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0173_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold165 (.A(\inst_calculator.reg_arg[1] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold166 (.A(\inst_calculator.reg_arg[0] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold167 (.A(\inst_calculator.inst_divider.numerator[9] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0162_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold169 (.A(\inst_calculator.inst_divider.n[3] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0131_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold171 (.A(\inst_calculator.denominator[9] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0116_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold173 (.A(\inst_calculator.inst_divider.n[6] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0134_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold175 (.A(\inst_calculator.inst_keypad_poller.state[3] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0014_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0051_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0665_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0045_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0597_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold181 (.A(\inst_calculator.inst_divider.busy ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold182 (.A(\inst_calculator.inst_divider.numerator[8] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0161_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold184 (.A(\inst_calculator.inst_drive.cnt0[7] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0657_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold186 (.A(\inst_calculator.inst_keypad_encoder.key[3] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0602_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold188 (.A(\inst_calculator.reg_arg[8] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold189 (.A(\inst_calculator.inst_drive.cnt0[10] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0663_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold191 (.A(\inst_calculator.inst_keypad_poller.clk_counter[10] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0997_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0089_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold194 (.A(\inst_calculator.inst_drive.cnt0[9] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold195 (.A(\inst_calculator.inst_divider.n[7] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0135_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold197 (.A(\inst_calculator.inst_bin2bcd.bin_in[5] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0177_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold199 (.A(\inst_calculator.inst_divider.n[2] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0130_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold201 (.A(\inst_calculator.inst_keypad_encoder.rows[1] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0193_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold203 (.A(\inst_calculator.inst_keypad_encoder.key[2] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold204 (.A(\inst_calculator.inst_keypad_poller.clk_counter[9] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold205 (.A(\inst_calculator.inst_divider.q[8] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0475_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0164_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold208 (.A(\inst_calculator.inst_drive.cnt0[13] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0026_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold210 (.A(\inst_calculator.inst_keypad_poller.clk_counter[14] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold211 (.A(_1005_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold212 (.A(\inst_calculator.state[9] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0016_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold214 (.A(\inst_calculator.inst_keypad_poller.clk_counter[13] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold215 (.A(_1003_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0092_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold217 (.A(\inst_calculator.inst_keypad_poller.clk_counter[12] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold218 (.A(_1001_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold219 (.A(\inst_calculator.inst_keypad_poller.clk_counter[15] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold220 (.A(\inst_calculator.inst_keypad_poller.clk_counter[11] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold221 (.A(\inst_calculator.inst_divider.n[8] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0136_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold223 (.A(\inst_calculator.inst_drive.cnt0[9] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold224 (.A(\inst_calculator.inst_keypad_encoder.rows[2] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0194_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold226 (.A(\inst_calculator.reg_result[9] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold227 (.A(\inst_calculator.inst_drive.cnt_sel[1] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold228 (.A(\inst_calculator.inst_drive.cnt0[4] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold229 (.A(\inst_calculator.inst_keypad_poller.clk_counter[7] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold230 (.A(\inst_calculator.inst_keypad_encoder.key[2] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold231 (.A(\inst_calculator.divider_done ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0631_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0017_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold234 (.A(\inst_calculator.inst_keypad_poller.clk_counter[16] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold235 (.A(\inst_calculator.inst_drive.cnt0[5] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold236 (.A(\inst_calculator.state[1] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0018_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold238 (.A(\inst_calculator.reg_result[4] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold239 (.A(\inst_calculator.reg_result[6] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold240 (.A(\inst_calculator.inst_drive.num_disp[3] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0005_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0044_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold243 (.A(uio_out[6]),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0147_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold245 (.A(\inst_calculator.reg_arg[9] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold246 (.A(uio_out[5]),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold247 (.A(\inst_calculator.reg_result[5] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold248 (.A(\inst_calculator.inst_drive.num_disp[2] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0001_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold250 (.A(\inst_calculator.inst_bin2bcd.bin_in[8] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0174_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold252 (.A(\inst_calculator.inst_divider.q[1] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0171_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold254 (.A(\inst_calculator.reg_result[7] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold255 (.A(uio_out[4]),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold256 (.A(\inst_calculator.inst_bin2bcd.bin_in[7] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0175_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold258 (.A(\inst_calculator.inst_divider.q[0] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold259 (.A(_0172_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold260 (.A(\inst_calculator.reg_result[3] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold261 (.A(\inst_calculator.reg_result[2] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0170_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold263 (.A(\inst_calculator.inst_drive.num_disp[0] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0635_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold265 (.A(_0000_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold266 (.A(uio_out[7]),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0878_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0880_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0881_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold270 (.A(\inst_calculator.reg_arg[4] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold271 (.A(\inst_calculator.reg_arg[7] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold272 (.A(\inst_calculator.inst_divider.n[4] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold273 (.A(uio_out[4]),
    .X(net451));
 sg13g2_fill_2 FILLER_0_0 ();
 sg13g2_fill_1 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_72 ();
 sg13g2_decap_8 FILLER_0_79 ();
 sg13g2_decap_8 FILLER_0_86 ();
 sg13g2_decap_8 FILLER_0_93 ();
 sg13g2_decap_8 FILLER_0_100 ();
 sg13g2_decap_8 FILLER_0_107 ();
 sg13g2_decap_8 FILLER_0_114 ();
 sg13g2_decap_8 FILLER_0_121 ();
 sg13g2_decap_8 FILLER_0_128 ();
 sg13g2_decap_8 FILLER_0_135 ();
 sg13g2_decap_8 FILLER_0_142 ();
 sg13g2_decap_8 FILLER_0_149 ();
 sg13g2_decap_8 FILLER_0_156 ();
 sg13g2_decap_8 FILLER_0_163 ();
 sg13g2_decap_8 FILLER_0_170 ();
 sg13g2_decap_8 FILLER_0_177 ();
 sg13g2_decap_8 FILLER_0_184 ();
 sg13g2_decap_8 FILLER_0_191 ();
 sg13g2_decap_8 FILLER_0_198 ();
 sg13g2_decap_8 FILLER_0_205 ();
 sg13g2_decap_8 FILLER_0_212 ();
 sg13g2_decap_8 FILLER_0_219 ();
 sg13g2_decap_8 FILLER_0_226 ();
 sg13g2_decap_8 FILLER_0_233 ();
 sg13g2_decap_8 FILLER_0_279 ();
 sg13g2_decap_8 FILLER_0_286 ();
 sg13g2_decap_8 FILLER_0_293 ();
 sg13g2_decap_8 FILLER_0_300 ();
 sg13g2_decap_8 FILLER_0_307 ();
 sg13g2_fill_1 FILLER_0_314 ();
 sg13g2_fill_2 FILLER_0_327 ();
 sg13g2_fill_1 FILLER_0_329 ();
 sg13g2_fill_2 FILLER_0_338 ();
 sg13g2_fill_1 FILLER_0_349 ();
 sg13g2_decap_8 FILLER_0_355 ();
 sg13g2_decap_8 FILLER_0_362 ();
 sg13g2_decap_8 FILLER_0_369 ();
 sg13g2_decap_8 FILLER_0_376 ();
 sg13g2_decap_8 FILLER_0_383 ();
 sg13g2_decap_8 FILLER_0_390 ();
 sg13g2_decap_8 FILLER_0_397 ();
 sg13g2_decap_4 FILLER_0_404 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_fill_1 FILLER_1_0 ();
 sg13g2_fill_1 FILLER_1_39 ();
 sg13g2_fill_2 FILLER_1_49 ();
 sg13g2_fill_1 FILLER_1_51 ();
 sg13g2_decap_8 FILLER_1_82 ();
 sg13g2_decap_8 FILLER_1_89 ();
 sg13g2_decap_8 FILLER_1_96 ();
 sg13g2_decap_8 FILLER_1_103 ();
 sg13g2_decap_8 FILLER_1_110 ();
 sg13g2_decap_8 FILLER_1_117 ();
 sg13g2_decap_8 FILLER_1_124 ();
 sg13g2_decap_8 FILLER_1_131 ();
 sg13g2_decap_8 FILLER_1_138 ();
 sg13g2_decap_8 FILLER_1_145 ();
 sg13g2_decap_8 FILLER_1_152 ();
 sg13g2_decap_8 FILLER_1_159 ();
 sg13g2_decap_8 FILLER_1_166 ();
 sg13g2_decap_8 FILLER_1_173 ();
 sg13g2_decap_8 FILLER_1_180 ();
 sg13g2_decap_8 FILLER_1_187 ();
 sg13g2_decap_8 FILLER_1_194 ();
 sg13g2_decap_8 FILLER_1_201 ();
 sg13g2_decap_8 FILLER_1_208 ();
 sg13g2_decap_8 FILLER_1_215 ();
 sg13g2_decap_8 FILLER_1_222 ();
 sg13g2_fill_2 FILLER_1_229 ();
 sg13g2_fill_1 FILLER_1_231 ();
 sg13g2_fill_1 FILLER_1_259 ();
 sg13g2_fill_2 FILLER_1_319 ();
 sg13g2_fill_2 FILLER_1_325 ();
 sg13g2_fill_1 FILLER_1_327 ();
 sg13g2_fill_1 FILLER_1_341 ();
 sg13g2_fill_2 FILLER_1_365 ();
 sg13g2_fill_1 FILLER_1_367 ();
 sg13g2_decap_4 FILLER_1_373 ();
 sg13g2_fill_1 FILLER_1_387 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_fill_1 FILLER_2_61 ();
 sg13g2_decap_8 FILLER_2_88 ();
 sg13g2_decap_8 FILLER_2_95 ();
 sg13g2_decap_8 FILLER_2_102 ();
 sg13g2_decap_8 FILLER_2_109 ();
 sg13g2_decap_8 FILLER_2_116 ();
 sg13g2_decap_4 FILLER_2_123 ();
 sg13g2_fill_2 FILLER_2_127 ();
 sg13g2_decap_8 FILLER_2_141 ();
 sg13g2_decap_8 FILLER_2_156 ();
 sg13g2_decap_8 FILLER_2_163 ();
 sg13g2_decap_4 FILLER_2_170 ();
 sg13g2_fill_2 FILLER_2_179 ();
 sg13g2_decap_8 FILLER_2_188 ();
 sg13g2_decap_8 FILLER_2_195 ();
 sg13g2_decap_8 FILLER_2_202 ();
 sg13g2_fill_1 FILLER_2_209 ();
 sg13g2_decap_8 FILLER_2_214 ();
 sg13g2_fill_2 FILLER_2_272 ();
 sg13g2_fill_1 FILLER_2_274 ();
 sg13g2_fill_2 FILLER_2_290 ();
 sg13g2_decap_4 FILLER_2_403 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_fill_1 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_3_27 ();
 sg13g2_fill_2 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_97 ();
 sg13g2_decap_8 FILLER_3_104 ();
 sg13g2_decap_8 FILLER_3_111 ();
 sg13g2_fill_2 FILLER_3_118 ();
 sg13g2_decap_4 FILLER_3_164 ();
 sg13g2_fill_1 FILLER_3_168 ();
 sg13g2_fill_1 FILLER_3_190 ();
 sg13g2_fill_1 FILLER_3_230 ();
 sg13g2_fill_2 FILLER_3_260 ();
 sg13g2_fill_1 FILLER_3_262 ();
 sg13g2_fill_2 FILLER_3_350 ();
 sg13g2_fill_1 FILLER_3_352 ();
 sg13g2_fill_2 FILLER_3_385 ();
 sg13g2_fill_1 FILLER_3_387 ();
 sg13g2_fill_2 FILLER_3_393 ();
 sg13g2_fill_1 FILLER_3_395 ();
 sg13g2_fill_1 FILLER_4_35 ();
 sg13g2_fill_2 FILLER_4_46 ();
 sg13g2_fill_1 FILLER_4_48 ();
 sg13g2_fill_1 FILLER_4_96 ();
 sg13g2_fill_1 FILLER_4_102 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_fill_1 FILLER_4_126 ();
 sg13g2_fill_2 FILLER_4_131 ();
 sg13g2_decap_8 FILLER_4_142 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_fill_2 FILLER_4_161 ();
 sg13g2_fill_1 FILLER_4_163 ();
 sg13g2_fill_1 FILLER_4_169 ();
 sg13g2_decap_8 FILLER_4_186 ();
 sg13g2_decap_4 FILLER_4_193 ();
 sg13g2_fill_1 FILLER_4_197 ();
 sg13g2_fill_2 FILLER_4_208 ();
 sg13g2_fill_2 FILLER_4_254 ();
 sg13g2_fill_1 FILLER_4_256 ();
 sg13g2_fill_1 FILLER_4_288 ();
 sg13g2_fill_1 FILLER_5_23 ();
 sg13g2_fill_1 FILLER_5_32 ();
 sg13g2_fill_2 FILLER_5_40 ();
 sg13g2_fill_1 FILLER_5_42 ();
 sg13g2_fill_2 FILLER_5_61 ();
 sg13g2_fill_1 FILLER_5_63 ();
 sg13g2_fill_2 FILLER_5_99 ();
 sg13g2_fill_1 FILLER_5_101 ();
 sg13g2_decap_4 FILLER_5_121 ();
 sg13g2_fill_2 FILLER_5_125 ();
 sg13g2_decap_8 FILLER_5_148 ();
 sg13g2_decap_8 FILLER_5_155 ();
 sg13g2_fill_1 FILLER_5_162 ();
 sg13g2_decap_4 FILLER_5_171 ();
 sg13g2_decap_8 FILLER_5_180 ();
 sg13g2_fill_2 FILLER_5_214 ();
 sg13g2_fill_1 FILLER_5_233 ();
 sg13g2_fill_2 FILLER_5_252 ();
 sg13g2_fill_1 FILLER_5_254 ();
 sg13g2_fill_1 FILLER_5_302 ();
 sg13g2_fill_1 FILLER_5_317 ();
 sg13g2_fill_2 FILLER_5_375 ();
 sg13g2_fill_1 FILLER_5_377 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_fill_2 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_33 ();
 sg13g2_fill_2 FILLER_6_60 ();
 sg13g2_fill_1 FILLER_6_62 ();
 sg13g2_decap_4 FILLER_6_81 ();
 sg13g2_decap_4 FILLER_6_109 ();
 sg13g2_fill_1 FILLER_6_113 ();
 sg13g2_decap_4 FILLER_6_133 ();
 sg13g2_fill_2 FILLER_6_137 ();
 sg13g2_fill_2 FILLER_6_165 ();
 sg13g2_decap_8 FILLER_6_185 ();
 sg13g2_fill_2 FILLER_6_192 ();
 sg13g2_fill_1 FILLER_6_194 ();
 sg13g2_fill_1 FILLER_6_209 ();
 sg13g2_fill_2 FILLER_6_255 ();
 sg13g2_fill_1 FILLER_6_306 ();
 sg13g2_fill_2 FILLER_6_364 ();
 sg13g2_fill_1 FILLER_6_366 ();
 sg13g2_fill_2 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_28 ();
 sg13g2_fill_2 FILLER_7_56 ();
 sg13g2_fill_1 FILLER_7_67 ();
 sg13g2_fill_2 FILLER_7_90 ();
 sg13g2_fill_1 FILLER_7_92 ();
 sg13g2_fill_2 FILLER_7_105 ();
 sg13g2_fill_2 FILLER_7_118 ();
 sg13g2_fill_1 FILLER_7_138 ();
 sg13g2_decap_4 FILLER_7_164 ();
 sg13g2_fill_2 FILLER_7_168 ();
 sg13g2_decap_4 FILLER_7_189 ();
 sg13g2_fill_2 FILLER_7_234 ();
 sg13g2_fill_1 FILLER_7_236 ();
 sg13g2_fill_2 FILLER_7_269 ();
 sg13g2_fill_1 FILLER_7_276 ();
 sg13g2_fill_1 FILLER_7_316 ();
 sg13g2_fill_2 FILLER_7_382 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_fill_1 FILLER_8_86 ();
 sg13g2_decap_4 FILLER_8_111 ();
 sg13g2_fill_1 FILLER_8_115 ();
 sg13g2_fill_1 FILLER_8_125 ();
 sg13g2_fill_2 FILLER_8_168 ();
 sg13g2_fill_2 FILLER_8_180 ();
 sg13g2_fill_1 FILLER_8_190 ();
 sg13g2_fill_2 FILLER_8_218 ();
 sg13g2_fill_1 FILLER_8_234 ();
 sg13g2_fill_2 FILLER_8_245 ();
 sg13g2_fill_1 FILLER_8_247 ();
 sg13g2_fill_2 FILLER_8_253 ();
 sg13g2_fill_1 FILLER_8_318 ();
 sg13g2_fill_1 FILLER_8_363 ();
 sg13g2_fill_1 FILLER_9_26 ();
 sg13g2_fill_2 FILLER_9_50 ();
 sg13g2_fill_1 FILLER_9_74 ();
 sg13g2_decap_4 FILLER_9_90 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_114 ();
 sg13g2_fill_1 FILLER_9_136 ();
 sg13g2_decap_8 FILLER_9_141 ();
 sg13g2_fill_2 FILLER_9_148 ();
 sg13g2_fill_2 FILLER_9_164 ();
 sg13g2_fill_1 FILLER_9_166 ();
 sg13g2_decap_8 FILLER_9_193 ();
 sg13g2_decap_4 FILLER_9_200 ();
 sg13g2_fill_2 FILLER_9_213 ();
 sg13g2_fill_1 FILLER_9_215 ();
 sg13g2_fill_1 FILLER_9_225 ();
 sg13g2_fill_1 FILLER_9_284 ();
 sg13g2_fill_1 FILLER_9_294 ();
 sg13g2_fill_2 FILLER_9_325 ();
 sg13g2_fill_2 FILLER_9_336 ();
 sg13g2_fill_1 FILLER_9_338 ();
 sg13g2_fill_2 FILLER_9_349 ();
 sg13g2_fill_1 FILLER_9_351 ();
 sg13g2_fill_2 FILLER_9_372 ();
 sg13g2_fill_1 FILLER_9_374 ();
 sg13g2_fill_2 FILLER_9_397 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_4 ();
 sg13g2_fill_2 FILLER_10_86 ();
 sg13g2_fill_1 FILLER_10_88 ();
 sg13g2_fill_2 FILLER_10_113 ();
 sg13g2_fill_2 FILLER_10_133 ();
 sg13g2_decap_4 FILLER_10_151 ();
 sg13g2_decap_8 FILLER_10_159 ();
 sg13g2_decap_4 FILLER_10_166 ();
 sg13g2_fill_2 FILLER_10_170 ();
 sg13g2_fill_2 FILLER_10_180 ();
 sg13g2_fill_1 FILLER_10_201 ();
 sg13g2_decap_8 FILLER_10_211 ();
 sg13g2_decap_8 FILLER_10_218 ();
 sg13g2_decap_4 FILLER_10_225 ();
 sg13g2_fill_2 FILLER_10_247 ();
 sg13g2_fill_2 FILLER_10_310 ();
 sg13g2_fill_2 FILLER_10_381 ();
 sg13g2_fill_1 FILLER_10_383 ();
 sg13g2_fill_2 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_7 ();
 sg13g2_fill_2 FILLER_11_24 ();
 sg13g2_fill_2 FILLER_11_31 ();
 sg13g2_fill_2 FILLER_11_55 ();
 sg13g2_fill_1 FILLER_11_72 ();
 sg13g2_decap_8 FILLER_11_82 ();
 sg13g2_fill_1 FILLER_11_89 ();
 sg13g2_fill_1 FILLER_11_100 ();
 sg13g2_decap_8 FILLER_11_110 ();
 sg13g2_fill_1 FILLER_11_122 ();
 sg13g2_decap_8 FILLER_11_135 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_fill_1 FILLER_11_154 ();
 sg13g2_fill_2 FILLER_11_160 ();
 sg13g2_fill_1 FILLER_11_162 ();
 sg13g2_fill_2 FILLER_11_168 ();
 sg13g2_fill_2 FILLER_11_174 ();
 sg13g2_fill_1 FILLER_11_176 ();
 sg13g2_fill_2 FILLER_11_187 ();
 sg13g2_fill_1 FILLER_11_189 ();
 sg13g2_decap_4 FILLER_11_216 ();
 sg13g2_fill_1 FILLER_11_238 ();
 sg13g2_fill_2 FILLER_11_251 ();
 sg13g2_fill_2 FILLER_11_258 ();
 sg13g2_fill_2 FILLER_11_294 ();
 sg13g2_fill_1 FILLER_11_296 ();
 sg13g2_fill_1 FILLER_11_307 ();
 sg13g2_fill_1 FILLER_11_340 ();
 sg13g2_fill_2 FILLER_12_72 ();
 sg13g2_fill_2 FILLER_12_87 ();
 sg13g2_fill_2 FILLER_12_113 ();
 sg13g2_fill_1 FILLER_12_115 ();
 sg13g2_fill_2 FILLER_12_124 ();
 sg13g2_fill_1 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_132 ();
 sg13g2_fill_1 FILLER_12_139 ();
 sg13g2_decap_4 FILLER_12_145 ();
 sg13g2_fill_1 FILLER_12_149 ();
 sg13g2_fill_2 FILLER_12_155 ();
 sg13g2_decap_8 FILLER_12_179 ();
 sg13g2_fill_2 FILLER_12_196 ();
 sg13g2_fill_1 FILLER_12_198 ();
 sg13g2_decap_4 FILLER_12_209 ();
 sg13g2_fill_1 FILLER_12_213 ();
 sg13g2_fill_1 FILLER_12_238 ();
 sg13g2_fill_2 FILLER_12_274 ();
 sg13g2_fill_1 FILLER_12_276 ();
 sg13g2_fill_2 FILLER_12_291 ();
 sg13g2_fill_1 FILLER_12_293 ();
 sg13g2_fill_1 FILLER_12_382 ();
 sg13g2_decap_4 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_4 ();
 sg13g2_decap_4 FILLER_13_63 ();
 sg13g2_decap_4 FILLER_13_87 ();
 sg13g2_decap_4 FILLER_13_111 ();
 sg13g2_decap_8 FILLER_13_123 ();
 sg13g2_fill_1 FILLER_13_130 ();
 sg13g2_fill_2 FILLER_13_139 ();
 sg13g2_fill_1 FILLER_13_141 ();
 sg13g2_fill_1 FILLER_13_161 ();
 sg13g2_decap_4 FILLER_13_166 ();
 sg13g2_fill_1 FILLER_13_170 ();
 sg13g2_decap_8 FILLER_13_181 ();
 sg13g2_decap_4 FILLER_13_209 ();
 sg13g2_fill_2 FILLER_13_213 ();
 sg13g2_fill_2 FILLER_13_222 ();
 sg13g2_decap_8 FILLER_13_234 ();
 sg13g2_decap_4 FILLER_13_241 ();
 sg13g2_fill_1 FILLER_13_245 ();
 sg13g2_fill_2 FILLER_13_260 ();
 sg13g2_fill_2 FILLER_13_309 ();
 sg13g2_fill_1 FILLER_13_311 ();
 sg13g2_fill_1 FILLER_13_329 ();
 sg13g2_fill_1 FILLER_13_390 ();
 sg13g2_fill_2 FILLER_14_26 ();
 sg13g2_decap_4 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_fill_1 FILLER_14_112 ();
 sg13g2_fill_2 FILLER_14_136 ();
 sg13g2_fill_1 FILLER_14_138 ();
 sg13g2_decap_4 FILLER_14_143 ();
 sg13g2_fill_2 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_fill_2 FILLER_14_170 ();
 sg13g2_fill_1 FILLER_14_172 ();
 sg13g2_fill_2 FILLER_14_181 ();
 sg13g2_fill_1 FILLER_14_183 ();
 sg13g2_decap_8 FILLER_14_197 ();
 sg13g2_decap_8 FILLER_14_204 ();
 sg13g2_fill_2 FILLER_14_226 ();
 sg13g2_fill_2 FILLER_14_244 ();
 sg13g2_fill_1 FILLER_14_256 ();
 sg13g2_fill_1 FILLER_14_301 ();
 sg13g2_decap_4 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_44 ();
 sg13g2_fill_1 FILLER_15_66 ();
 sg13g2_fill_1 FILLER_15_136 ();
 sg13g2_fill_1 FILLER_15_158 ();
 sg13g2_decap_4 FILLER_15_177 ();
 sg13g2_decap_8 FILLER_15_185 ();
 sg13g2_decap_8 FILLER_15_192 ();
 sg13g2_decap_4 FILLER_15_207 ();
 sg13g2_fill_1 FILLER_15_211 ();
 sg13g2_fill_2 FILLER_15_225 ();
 sg13g2_fill_1 FILLER_15_227 ();
 sg13g2_decap_8 FILLER_15_235 ();
 sg13g2_fill_2 FILLER_15_264 ();
 sg13g2_fill_1 FILLER_15_277 ();
 sg13g2_fill_1 FILLER_15_291 ();
 sg13g2_fill_1 FILLER_15_301 ();
 sg13g2_fill_2 FILLER_15_311 ();
 sg13g2_fill_2 FILLER_15_343 ();
 sg13g2_fill_1 FILLER_15_345 ();
 sg13g2_fill_2 FILLER_15_355 ();
 sg13g2_fill_1 FILLER_15_357 ();
 sg13g2_fill_2 FILLER_15_366 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_11 ();
 sg13g2_fill_1 FILLER_16_40 ();
 sg13g2_fill_2 FILLER_16_46 ();
 sg13g2_decap_4 FILLER_16_72 ();
 sg13g2_decap_8 FILLER_16_103 ();
 sg13g2_decap_8 FILLER_16_110 ();
 sg13g2_fill_2 FILLER_16_117 ();
 sg13g2_decap_8 FILLER_16_129 ();
 sg13g2_fill_2 FILLER_16_150 ();
 sg13g2_fill_1 FILLER_16_156 ();
 sg13g2_fill_1 FILLER_16_173 ();
 sg13g2_decap_8 FILLER_16_209 ();
 sg13g2_decap_8 FILLER_16_216 ();
 sg13g2_fill_2 FILLER_16_249 ();
 sg13g2_fill_1 FILLER_16_266 ();
 sg13g2_fill_2 FILLER_16_316 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_28 ();
 sg13g2_fill_2 FILLER_17_37 ();
 sg13g2_fill_2 FILLER_17_43 ();
 sg13g2_decap_4 FILLER_17_72 ();
 sg13g2_fill_2 FILLER_17_76 ();
 sg13g2_decap_4 FILLER_17_102 ();
 sg13g2_fill_2 FILLER_17_106 ();
 sg13g2_fill_1 FILLER_17_117 ();
 sg13g2_decap_4 FILLER_17_124 ();
 sg13g2_fill_1 FILLER_17_128 ();
 sg13g2_fill_2 FILLER_17_141 ();
 sg13g2_fill_1 FILLER_17_143 ();
 sg13g2_fill_2 FILLER_17_155 ();
 sg13g2_fill_2 FILLER_17_183 ();
 sg13g2_fill_2 FILLER_17_197 ();
 sg13g2_fill_2 FILLER_17_203 ();
 sg13g2_fill_1 FILLER_17_205 ();
 sg13g2_fill_1 FILLER_17_226 ();
 sg13g2_fill_2 FILLER_17_259 ();
 sg13g2_fill_2 FILLER_17_270 ();
 sg13g2_fill_1 FILLER_17_272 ();
 sg13g2_fill_1 FILLER_17_317 ();
 sg13g2_fill_2 FILLER_17_332 ();
 sg13g2_fill_1 FILLER_17_353 ();
 sg13g2_fill_1 FILLER_17_363 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_7 ();
 sg13g2_fill_2 FILLER_18_30 ();
 sg13g2_fill_1 FILLER_18_32 ();
 sg13g2_fill_2 FILLER_18_68 ();
 sg13g2_decap_8 FILLER_18_79 ();
 sg13g2_fill_1 FILLER_18_86 ();
 sg13g2_decap_4 FILLER_18_93 ();
 sg13g2_fill_2 FILLER_18_102 ();
 sg13g2_decap_4 FILLER_18_121 ();
 sg13g2_fill_1 FILLER_18_125 ();
 sg13g2_fill_1 FILLER_18_131 ();
 sg13g2_fill_2 FILLER_18_152 ();
 sg13g2_fill_1 FILLER_18_154 ();
 sg13g2_fill_1 FILLER_18_165 ();
 sg13g2_fill_2 FILLER_18_181 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_fill_2 FILLER_18_203 ();
 sg13g2_fill_1 FILLER_18_213 ();
 sg13g2_decap_4 FILLER_18_219 ();
 sg13g2_fill_2 FILLER_18_239 ();
 sg13g2_fill_1 FILLER_18_249 ();
 sg13g2_fill_1 FILLER_18_275 ();
 sg13g2_fill_1 FILLER_18_342 ();
 sg13g2_fill_1 FILLER_18_370 ();
 sg13g2_fill_1 FILLER_18_382 ();
 sg13g2_decap_4 FILLER_19_26 ();
 sg13g2_fill_1 FILLER_19_37 ();
 sg13g2_fill_1 FILLER_19_47 ();
 sg13g2_decap_4 FILLER_19_104 ();
 sg13g2_fill_2 FILLER_19_124 ();
 sg13g2_fill_1 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_149 ();
 sg13g2_decap_4 FILLER_19_156 ();
 sg13g2_fill_1 FILLER_19_166 ();
 sg13g2_fill_2 FILLER_19_172 ();
 sg13g2_decap_8 FILLER_19_179 ();
 sg13g2_decap_8 FILLER_19_186 ();
 sg13g2_fill_2 FILLER_19_255 ();
 sg13g2_fill_1 FILLER_19_257 ();
 sg13g2_fill_2 FILLER_19_272 ();
 sg13g2_fill_1 FILLER_19_332 ();
 sg13g2_fill_1 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_4 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_15 ();
 sg13g2_decap_8 FILLER_20_22 ();
 sg13g2_fill_2 FILLER_20_29 ();
 sg13g2_fill_1 FILLER_20_31 ();
 sg13g2_fill_1 FILLER_20_50 ();
 sg13g2_fill_2 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_73 ();
 sg13g2_fill_2 FILLER_20_80 ();
 sg13g2_fill_2 FILLER_20_87 ();
 sg13g2_decap_8 FILLER_20_93 ();
 sg13g2_decap_4 FILLER_20_100 ();
 sg13g2_fill_1 FILLER_20_104 ();
 sg13g2_fill_2 FILLER_20_110 ();
 sg13g2_fill_1 FILLER_20_112 ();
 sg13g2_decap_4 FILLER_20_148 ();
 sg13g2_fill_2 FILLER_20_152 ();
 sg13g2_fill_2 FILLER_20_176 ();
 sg13g2_fill_1 FILLER_20_178 ();
 sg13g2_fill_1 FILLER_20_188 ();
 sg13g2_fill_2 FILLER_20_263 ();
 sg13g2_fill_2 FILLER_20_276 ();
 sg13g2_fill_1 FILLER_20_278 ();
 sg13g2_fill_2 FILLER_20_305 ();
 sg13g2_fill_1 FILLER_20_307 ();
 sg13g2_fill_2 FILLER_20_353 ();
 sg13g2_fill_1 FILLER_20_355 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_4 FILLER_21_75 ();
 sg13g2_decap_8 FILLER_21_83 ();
 sg13g2_decap_4 FILLER_21_90 ();
 sg13g2_fill_1 FILLER_21_98 ();
 sg13g2_fill_1 FILLER_21_123 ();
 sg13g2_fill_2 FILLER_21_132 ();
 sg13g2_fill_1 FILLER_21_138 ();
 sg13g2_decap_8 FILLER_21_143 ();
 sg13g2_decap_4 FILLER_21_150 ();
 sg13g2_fill_1 FILLER_21_162 ();
 sg13g2_fill_1 FILLER_21_168 ();
 sg13g2_fill_2 FILLER_21_177 ();
 sg13g2_fill_1 FILLER_21_205 ();
 sg13g2_fill_2 FILLER_21_240 ();
 sg13g2_fill_1 FILLER_21_242 ();
 sg13g2_fill_1 FILLER_21_271 ();
 sg13g2_fill_2 FILLER_21_318 ();
 sg13g2_fill_1 FILLER_21_320 ();
 sg13g2_fill_1 FILLER_21_382 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_4 ();
 sg13g2_fill_1 FILLER_22_42 ();
 sg13g2_fill_2 FILLER_22_80 ();
 sg13g2_fill_1 FILLER_22_82 ();
 sg13g2_fill_1 FILLER_22_109 ();
 sg13g2_fill_1 FILLER_22_117 ();
 sg13g2_fill_1 FILLER_22_185 ();
 sg13g2_fill_1 FILLER_22_207 ();
 sg13g2_fill_2 FILLER_22_221 ();
 sg13g2_fill_1 FILLER_22_223 ();
 sg13g2_fill_2 FILLER_22_263 ();
 sg13g2_fill_2 FILLER_22_340 ();
 sg13g2_fill_1 FILLER_22_342 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_7 ();
 sg13g2_decap_4 FILLER_23_18 ();
 sg13g2_fill_2 FILLER_23_22 ();
 sg13g2_fill_2 FILLER_23_29 ();
 sg13g2_fill_2 FILLER_23_45 ();
 sg13g2_fill_1 FILLER_23_47 ();
 sg13g2_decap_4 FILLER_23_64 ();
 sg13g2_fill_1 FILLER_23_68 ();
 sg13g2_decap_8 FILLER_23_86 ();
 sg13g2_decap_8 FILLER_23_93 ();
 sg13g2_fill_1 FILLER_23_100 ();
 sg13g2_fill_2 FILLER_23_110 ();
 sg13g2_fill_1 FILLER_23_133 ();
 sg13g2_decap_4 FILLER_23_138 ();
 sg13g2_fill_2 FILLER_23_142 ();
 sg13g2_decap_8 FILLER_23_149 ();
 sg13g2_decap_4 FILLER_23_160 ();
 sg13g2_fill_2 FILLER_23_164 ();
 sg13g2_fill_2 FILLER_23_313 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_2 ();
 sg13g2_decap_8 FILLER_24_20 ();
 sg13g2_fill_2 FILLER_24_44 ();
 sg13g2_fill_1 FILLER_24_46 ();
 sg13g2_fill_1 FILLER_24_54 ();
 sg13g2_fill_1 FILLER_24_62 ();
 sg13g2_fill_2 FILLER_24_116 ();
 sg13g2_fill_1 FILLER_24_118 ();
 sg13g2_fill_2 FILLER_24_145 ();
 sg13g2_decap_4 FILLER_24_151 ();
 sg13g2_fill_1 FILLER_24_155 ();
 sg13g2_fill_1 FILLER_24_178 ();
 sg13g2_fill_2 FILLER_24_205 ();
 sg13g2_fill_1 FILLER_24_237 ();
 sg13g2_fill_1 FILLER_24_255 ();
 sg13g2_fill_1 FILLER_24_261 ();
 sg13g2_fill_2 FILLER_24_279 ();
 sg13g2_fill_2 FILLER_24_331 ();
 sg13g2_fill_1 FILLER_24_333 ();
 sg13g2_fill_2 FILLER_24_358 ();
 sg13g2_fill_1 FILLER_24_360 ();
 sg13g2_fill_2 FILLER_24_371 ();
 sg13g2_fill_1 FILLER_24_382 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_27 ();
 sg13g2_fill_2 FILLER_25_34 ();
 sg13g2_fill_1 FILLER_25_36 ();
 sg13g2_fill_2 FILLER_25_44 ();
 sg13g2_fill_2 FILLER_25_56 ();
 sg13g2_fill_1 FILLER_25_58 ();
 sg13g2_decap_8 FILLER_25_78 ();
 sg13g2_fill_1 FILLER_25_85 ();
 sg13g2_fill_1 FILLER_25_98 ();
 sg13g2_fill_1 FILLER_25_108 ();
 sg13g2_fill_2 FILLER_25_114 ();
 sg13g2_decap_4 FILLER_25_124 ();
 sg13g2_fill_2 FILLER_25_128 ();
 sg13g2_fill_2 FILLER_25_134 ();
 sg13g2_fill_2 FILLER_25_162 ();
 sg13g2_fill_1 FILLER_25_294 ();
 sg13g2_fill_2 FILLER_25_305 ();
 sg13g2_fill_2 FILLER_25_337 ();
 sg13g2_fill_2 FILLER_25_365 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_2 ();
 sg13g2_decap_8 FILLER_26_24 ();
 sg13g2_decap_8 FILLER_26_31 ();
 sg13g2_decap_4 FILLER_26_38 ();
 sg13g2_fill_1 FILLER_26_42 ();
 sg13g2_decap_4 FILLER_26_48 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_fill_1 FILLER_26_63 ();
 sg13g2_fill_2 FILLER_26_76 ();
 sg13g2_fill_1 FILLER_26_78 ();
 sg13g2_decap_4 FILLER_26_96 ();
 sg13g2_fill_1 FILLER_26_100 ();
 sg13g2_decap_4 FILLER_26_131 ();
 sg13g2_fill_2 FILLER_26_151 ();
 sg13g2_fill_2 FILLER_26_178 ();
 sg13g2_fill_1 FILLER_26_185 ();
 sg13g2_fill_1 FILLER_26_191 ();
 sg13g2_fill_1 FILLER_26_200 ();
 sg13g2_fill_2 FILLER_26_271 ();
 sg13g2_fill_2 FILLER_26_303 ();
 sg13g2_fill_2 FILLER_26_391 ();
 sg13g2_fill_1 FILLER_26_393 ();
 sg13g2_fill_2 FILLER_26_398 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_7 ();
 sg13g2_fill_1 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_54 ();
 sg13g2_fill_1 FILLER_27_124 ();
 sg13g2_fill_2 FILLER_27_139 ();
 sg13g2_fill_1 FILLER_27_141 ();
 sg13g2_fill_2 FILLER_27_177 ();
 sg13g2_fill_1 FILLER_27_200 ();
 sg13g2_fill_1 FILLER_27_269 ();
 sg13g2_fill_1 FILLER_27_302 ();
 sg13g2_fill_2 FILLER_27_352 ();
 sg13g2_fill_2 FILLER_27_368 ();
 sg13g2_fill_1 FILLER_27_370 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_2 ();
 sg13g2_fill_2 FILLER_28_31 ();
 sg13g2_fill_1 FILLER_28_33 ();
 sg13g2_fill_1 FILLER_28_41 ();
 sg13g2_decap_8 FILLER_28_52 ();
 sg13g2_decap_4 FILLER_28_59 ();
 sg13g2_fill_1 FILLER_28_63 ();
 sg13g2_decap_4 FILLER_28_74 ();
 sg13g2_fill_1 FILLER_28_100 ();
 sg13g2_fill_1 FILLER_28_106 ();
 sg13g2_fill_2 FILLER_28_147 ();
 sg13g2_fill_1 FILLER_28_149 ();
 sg13g2_fill_2 FILLER_28_185 ();
 sg13g2_fill_1 FILLER_28_214 ();
 sg13g2_fill_2 FILLER_28_241 ();
 sg13g2_fill_2 FILLER_28_262 ();
 sg13g2_fill_1 FILLER_28_273 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_20 ();
 sg13g2_fill_1 FILLER_29_22 ();
 sg13g2_fill_2 FILLER_29_28 ();
 sg13g2_fill_1 FILLER_29_30 ();
 sg13g2_fill_1 FILLER_29_42 ();
 sg13g2_fill_2 FILLER_29_77 ();
 sg13g2_fill_2 FILLER_29_84 ();
 sg13g2_fill_1 FILLER_29_98 ();
 sg13g2_fill_2 FILLER_29_112 ();
 sg13g2_fill_2 FILLER_29_175 ();
 sg13g2_fill_2 FILLER_29_212 ();
 sg13g2_fill_1 FILLER_29_263 ();
 sg13g2_fill_1 FILLER_29_347 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_7 ();
 sg13g2_decap_4 FILLER_30_49 ();
 sg13g2_fill_1 FILLER_30_53 ();
 sg13g2_fill_1 FILLER_30_73 ();
 sg13g2_fill_2 FILLER_30_86 ();
 sg13g2_fill_1 FILLER_30_162 ();
 sg13g2_fill_1 FILLER_30_193 ();
 sg13g2_fill_2 FILLER_30_221 ();
 sg13g2_fill_2 FILLER_30_298 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_23 ();
 sg13g2_fill_2 FILLER_31_32 ();
 sg13g2_fill_1 FILLER_31_34 ();
 sg13g2_fill_1 FILLER_31_41 ();
 sg13g2_decap_4 FILLER_31_47 ();
 sg13g2_fill_1 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_71 ();
 sg13g2_fill_1 FILLER_31_81 ();
 sg13g2_fill_2 FILLER_31_113 ();
 sg13g2_fill_2 FILLER_31_144 ();
 sg13g2_fill_2 FILLER_31_154 ();
 sg13g2_fill_1 FILLER_31_165 ();
 sg13g2_fill_2 FILLER_31_184 ();
 sg13g2_fill_1 FILLER_31_213 ();
 sg13g2_fill_1 FILLER_31_220 ();
 sg13g2_fill_1 FILLER_31_256 ();
 sg13g2_fill_1 FILLER_31_262 ();
 sg13g2_fill_2 FILLER_31_322 ();
 sg13g2_fill_1 FILLER_31_329 ();
 sg13g2_fill_1 FILLER_31_382 ();
 sg13g2_fill_1 FILLER_32_139 ();
 sg13g2_fill_1 FILLER_32_170 ();
 sg13g2_fill_1 FILLER_32_176 ();
 sg13g2_fill_2 FILLER_32_287 ();
 sg13g2_fill_2 FILLER_32_298 ();
 sg13g2_fill_1 FILLER_32_338 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_38 ();
 sg13g2_fill_1 FILLER_33_93 ();
 sg13g2_fill_2 FILLER_33_151 ();
 sg13g2_fill_1 FILLER_33_283 ();
 sg13g2_fill_1 FILLER_33_328 ();
 sg13g2_fill_1 FILLER_33_355 ();
 sg13g2_fill_2 FILLER_34_26 ();
 sg13g2_fill_1 FILLER_34_54 ();
 sg13g2_fill_2 FILLER_34_108 ();
 sg13g2_fill_1 FILLER_34_125 ();
 sg13g2_fill_1 FILLER_34_131 ();
 sg13g2_fill_1 FILLER_34_171 ();
 sg13g2_fill_2 FILLER_34_179 ();
 sg13g2_fill_1 FILLER_34_190 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_4 ();
 sg13g2_fill_1 FILLER_35_62 ();
 sg13g2_fill_1 FILLER_35_102 ();
 sg13g2_fill_1 FILLER_35_176 ();
 sg13g2_fill_1 FILLER_35_226 ();
 sg13g2_fill_2 FILLER_35_256 ();
 sg13g2_fill_1 FILLER_35_331 ();
 sg13g2_fill_2 FILLER_35_358 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_fill_1 FILLER_36_26 ();
 sg13g2_fill_1 FILLER_36_71 ();
 sg13g2_fill_1 FILLER_36_95 ();
 sg13g2_fill_2 FILLER_36_149 ();
 sg13g2_fill_1 FILLER_36_160 ();
 sg13g2_fill_2 FILLER_36_170 ();
 sg13g2_fill_2 FILLER_36_209 ();
 sg13g2_fill_2 FILLER_36_222 ();
 sg13g2_fill_1 FILLER_36_337 ();
 sg13g2_fill_1 FILLER_36_343 ();
 sg13g2_fill_1 FILLER_36_366 ();
 sg13g2_fill_1 FILLER_36_382 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_35 ();
 sg13g2_fill_1 FILLER_37_92 ();
 sg13g2_fill_1 FILLER_37_132 ();
 sg13g2_fill_1 FILLER_37_175 ();
 sg13g2_fill_1 FILLER_37_186 ();
 sg13g2_fill_1 FILLER_37_213 ();
 sg13g2_fill_2 FILLER_37_228 ();
 sg13g2_fill_1 FILLER_37_264 ();
 sg13g2_fill_2 FILLER_37_291 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_125 ();
 sg13g2_fill_1 FILLER_38_157 ();
 sg13g2_fill_1 FILLER_38_165 ();
 sg13g2_fill_2 FILLER_38_171 ();
 sg13g2_fill_1 FILLER_38_183 ();
 sg13g2_fill_1 FILLER_38_189 ();
 sg13g2_fill_1 FILLER_38_205 ();
 sg13g2_fill_2 FILLER_38_226 ();
 sg13g2_fill_2 FILLER_38_303 ();
 sg13g2_fill_1 FILLER_38_314 ();
 sg13g2_fill_1 FILLER_38_351 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net80;
 assign uio_oe[1] = net81;
 assign uio_oe[2] = net82;
 assign uio_oe[3] = net83;
 assign uio_oe[4] = net84;
 assign uio_oe[5] = net85;
 assign uio_oe[6] = net86;
 assign uio_oe[7] = net87;
 assign uio_out[0] = net5;
 assign uo_out[7] = net88;
endmodule

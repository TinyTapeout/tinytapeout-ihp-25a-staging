module tt_um_frequency_counter (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire clk_regs;
 wire \counter.cnt_ref_enable ;
 wire \counter.cnt_x_digits[0] ;
 wire \counter.cnt_x_digits[10] ;
 wire \counter.cnt_x_digits[11] ;
 wire \counter.cnt_x_digits[12] ;
 wire \counter.cnt_x_digits[13] ;
 wire \counter.cnt_x_digits[14] ;
 wire \counter.cnt_x_digits[15] ;
 wire \counter.cnt_x_digits[16] ;
 wire \counter.cnt_x_digits[17] ;
 wire \counter.cnt_x_digits[18] ;
 wire \counter.cnt_x_digits[19] ;
 wire \counter.cnt_x_digits[1] ;
 wire \counter.cnt_x_digits[20] ;
 wire \counter.cnt_x_digits[21] ;
 wire \counter.cnt_x_digits[22] ;
 wire \counter.cnt_x_digits[23] ;
 wire \counter.cnt_x_digits[2] ;
 wire \counter.cnt_x_digits[3] ;
 wire \counter.cnt_x_digits[4] ;
 wire \counter.cnt_x_digits[5] ;
 wire \counter.cnt_x_digits[6] ;
 wire \counter.cnt_x_digits[7] ;
 wire \counter.cnt_x_digits[8] ;
 wire \counter.cnt_x_digits[9] ;
 wire \counter.counter_ref.digit_0.digit_out[0] ;
 wire \counter.counter_ref.digit_0.digit_out[1] ;
 wire \counter.counter_ref.digit_0.digit_out[2] ;
 wire \counter.counter_ref.digit_0.digit_out[3] ;
 wire \counter.counter_ref.digits_out[10] ;
 wire \counter.counter_ref.digits_out[11] ;
 wire \counter.counter_ref.digits_out[12] ;
 wire \counter.counter_ref.digits_out[13] ;
 wire \counter.counter_ref.digits_out[14] ;
 wire \counter.counter_ref.digits_out[15] ;
 wire \counter.counter_ref.digits_out[16] ;
 wire \counter.counter_ref.digits_out[17] ;
 wire \counter.counter_ref.digits_out[18] ;
 wire \counter.counter_ref.digits_out[19] ;
 wire \counter.counter_ref.digits_out[20] ;
 wire \counter.counter_ref.digits_out[21] ;
 wire \counter.counter_ref.digits_out[22] ;
 wire \counter.counter_ref.digits_out[23] ;
 wire \counter.counter_ref.digits_out[4] ;
 wire \counter.counter_ref.digits_out[5] ;
 wire \counter.counter_ref.digits_out[6] ;
 wire \counter.counter_ref.digits_out[7] ;
 wire \counter.counter_ref.digits_out[8] ;
 wire \counter.counter_ref.digits_out[9] ;
 wire \counter.oled_clk_out ;
 wire \counter.oled_csn_out ;
 wire \counter.oled_dc_out ;
 wire \counter.oled_driver.mc_exec.delay_cnt[0] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[10] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[11] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[12] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[13] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[14] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[15] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[16] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[1] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[2] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[3] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[4] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[5] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[6] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[7] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[8] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[9] ;
 wire \counter.oled_driver.mc_exec.microcode_rom.address[0] ;
 wire \counter.oled_driver.mc_exec.microcode_rom.address[1] ;
 wire \counter.oled_driver.mc_exec.microcode_rom.address[2] ;
 wire \counter.oled_driver.mc_exec.microcode_rom.address[3] ;
 wire \counter.oled_driver.mc_exec.microcode_rom.address[4] ;
 wire \counter.oled_driver.mc_exec.microcode_rom.address[5] ;
 wire \counter.oled_driver.mc_exec.oled_dc_out ;
 wire \counter.oled_driver.mc_exec.oled_rstn_out ;
 wire \counter.oled_driver.mc_exec.oled_vbatn_out ;
 wire \counter.oled_driver.mc_exec.oled_vcdn_out ;
 wire \counter.oled_driver.mc_exec.procedure_done_out ;
 wire \counter.oled_driver.mc_exec.procedure_offset_in[0] ;
 wire \counter.oled_driver.mc_exec.procedure_start_in ;
 wire \counter.oled_driver.mc_exec.reset_in ;
 wire \counter.oled_driver.mc_exec.spi_tx_trigger_out ;
 wire \counter.oled_driver.mc_exec.state_r[0] ;
 wire \counter.oled_driver.mc_exec.state_r[2] ;
 wire \counter.oled_driver.mc_exec.state_r[3] ;
 wire \counter.oled_driver.mc_exec.state_r[5] ;
 wire \counter.oled_driver.mc_exec.state_r[6] ;
 wire \counter.oled_driver.oled_mosi_out ;
 wire \counter.oled_driver.ready_out ;
 wire \counter.oled_driver.spi_data[0] ;
 wire \counter.oled_driver.spi_data[1] ;
 wire \counter.oled_driver.spi_data[2] ;
 wire \counter.oled_driver.spi_data[3] ;
 wire \counter.oled_driver.spi_data[4] ;
 wire \counter.oled_driver.spi_data[5] ;
 wire \counter.oled_driver.spi_data[6] ;
 wire \counter.oled_driver.spi_data[7] ;
 wire \counter.oled_driver.spi_deactivate_cs ;
 wire \counter.oled_driver.spi_driver.deactivate_cs_r ;
 wire \counter.oled_driver.spi_driver.shift_reg.bit_counter_r[0] ;
 wire \counter.oled_driver.spi_driver.shift_reg.bit_counter_r[1] ;
 wire \counter.oled_driver.spi_driver.shift_reg.bit_counter_r[2] ;
 wire \counter.oled_driver.spi_driver.shift_reg.bit_counter_r[3] ;
 wire \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[0] ;
 wire \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[1] ;
 wire \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[2] ;
 wire \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[3] ;
 wire \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[4] ;
 wire \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[5] ;
 wire \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[6] ;
 wire \counter.oled_driver.spi_driver.shift_reg.start_in ;
 wire \counter.oled_driver.spi_driver.state_r[0] ;
 wire \counter.oled_driver.spi_driver.state_r[1] ;
 wire \counter.oled_driver.state_r[0] ;
 wire \counter.oled_driver.state_r[2] ;
 wire \counter.oled_driver.state_r[4] ;
 wire \counter.oled_driver.sync_stb_in ;
 wire \counter.oled_driver.write_stb_in ;
 wire \counter.refresh_display ;
 wire \counter.state[0] ;
 wire \counter.state[1] ;
 wire \counter.streamer.digit_cnt_r[0] ;
 wire \counter.streamer.digit_cnt_r[1] ;
 wire \counter.streamer.digit_cnt_r[2] ;
 wire \counter.streamer.digits_r[0] ;
 wire \counter.streamer.digits_r[10] ;
 wire \counter.streamer.digits_r[11] ;
 wire \counter.streamer.digits_r[12] ;
 wire \counter.streamer.digits_r[13] ;
 wire \counter.streamer.digits_r[14] ;
 wire \counter.streamer.digits_r[15] ;
 wire \counter.streamer.digits_r[16] ;
 wire \counter.streamer.digits_r[17] ;
 wire \counter.streamer.digits_r[18] ;
 wire \counter.streamer.digits_r[19] ;
 wire \counter.streamer.digits_r[1] ;
 wire \counter.streamer.digits_r[20] ;
 wire \counter.streamer.digits_r[21] ;
 wire \counter.streamer.digits_r[22] ;
 wire \counter.streamer.digits_r[23] ;
 wire \counter.streamer.digits_r[2] ;
 wire \counter.streamer.digits_r[3] ;
 wire \counter.streamer.digits_r[4] ;
 wire \counter.streamer.digits_r[5] ;
 wire \counter.streamer.digits_r[6] ;
 wire \counter.streamer.digits_r[7] ;
 wire \counter.streamer.digits_r[8] ;
 wire \counter.streamer.digits_r[9] ;
 wire \counter.streamer.graphical_decoder.index_x_in[0] ;
 wire \counter.streamer.graphical_decoder.index_x_in[1] ;
 wire \counter.streamer.graphical_decoder.index_x_in[2] ;
 wire \counter.streamer.graphical_decoder.index_x_in[3] ;
 wire \counter.streamer.graphical_decoder.index_x_in[4] ;
 wire \counter.streamer.graphical_decoder.index_y_in[0] ;
 wire \counter.streamer.graphical_decoder.index_y_in[1] ;
 wire \counter.streamer.graphical_decoder.pattern_adg[1] ;
 wire \counter.streamer.graphical_decoder.pattern_adg[2] ;
 wire \counter.streamer.graphical_decoder.pattern_adg[3] ;
 wire \counter.streamer.graphical_decoder.pattern_adg[4] ;
 wire \counter.streamer.ready_out ;
 wire \counter.streamer.state_r[4] ;
 wire \counter.streamer.state_r[5] ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net1;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire clknet_5_0__leaf_clk_regs;
 wire clknet_5_1__leaf_clk_regs;
 wire clknet_5_2__leaf_clk_regs;
 wire clknet_5_3__leaf_clk_regs;
 wire clknet_5_4__leaf_clk_regs;
 wire clknet_5_5__leaf_clk_regs;
 wire clknet_5_6__leaf_clk_regs;
 wire clknet_5_7__leaf_clk_regs;
 wire clknet_5_8__leaf_clk_regs;
 wire clknet_5_9__leaf_clk_regs;
 wire clknet_5_10__leaf_clk_regs;
 wire clknet_5_11__leaf_clk_regs;
 wire clknet_5_12__leaf_clk_regs;
 wire clknet_5_13__leaf_clk_regs;
 wire clknet_5_14__leaf_clk_regs;
 wire clknet_5_15__leaf_clk_regs;
 wire clknet_5_16__leaf_clk_regs;
 wire clknet_5_17__leaf_clk_regs;
 wire clknet_5_18__leaf_clk_regs;
 wire clknet_5_19__leaf_clk_regs;
 wire clknet_5_20__leaf_clk_regs;
 wire clknet_5_21__leaf_clk_regs;
 wire clknet_5_22__leaf_clk_regs;
 wire clknet_5_23__leaf_clk_regs;
 wire clknet_5_24__leaf_clk_regs;
 wire clknet_5_25__leaf_clk_regs;
 wire clknet_5_26__leaf_clk_regs;
 wire clknet_5_27__leaf_clk_regs;
 wire clknet_5_28__leaf_clk_regs;
 wire clknet_5_29__leaf_clk_regs;
 wire clknet_5_30__leaf_clk_regs;
 wire clknet_5_31__leaf_clk_regs;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;

 sg13g2_inv_1 _1296_ (.Y(_0529_),
    .A(net314));
 sg13g2_inv_1 _1297_ (.Y(_0530_),
    .A(net448));
 sg13g2_inv_1 _1298_ (.Y(_0531_),
    .A(\counter.counter_ref.digits_out[12] ));
 sg13g2_inv_1 _1299_ (.Y(_0532_),
    .A(net168));
 sg13g2_inv_1 _1300_ (.Y(_0533_),
    .A(\counter.cnt_x_digits[19] ));
 sg13g2_inv_1 _1301_ (.Y(_0534_),
    .A(\counter.cnt_x_digits[18] ));
 sg13g2_inv_1 _1302_ (.Y(_0535_),
    .A(\counter.cnt_x_digits[17] ));
 sg13g2_inv_1 _1303_ (.Y(_0536_),
    .A(\counter.cnt_x_digits[16] ));
 sg13g2_inv_1 _1304_ (.Y(_0537_),
    .A(\counter.cnt_x_digits[15] ));
 sg13g2_inv_1 _1305_ (.Y(_0538_),
    .A(\counter.cnt_x_digits[14] ));
 sg13g2_inv_1 _1306_ (.Y(_0539_),
    .A(\counter.cnt_x_digits[13] ));
 sg13g2_inv_1 _1307_ (.Y(_0540_),
    .A(\counter.cnt_x_digits[12] ));
 sg13g2_inv_1 _1308_ (.Y(_0541_),
    .A(\counter.cnt_x_digits[11] ));
 sg13g2_inv_1 _1309_ (.Y(_0542_),
    .A(\counter.cnt_x_digits[10] ));
 sg13g2_inv_1 _1310_ (.Y(_0543_),
    .A(\counter.cnt_x_digits[9] ));
 sg13g2_inv_1 _1311_ (.Y(_0544_),
    .A(\counter.cnt_x_digits[8] ));
 sg13g2_inv_1 _1312_ (.Y(_0545_),
    .A(\counter.cnt_x_digits[7] ));
 sg13g2_inv_1 _1313_ (.Y(_0546_),
    .A(\counter.cnt_x_digits[6] ));
 sg13g2_inv_1 _1314_ (.Y(_0547_),
    .A(\counter.cnt_x_digits[5] ));
 sg13g2_inv_1 _1315_ (.Y(_0548_),
    .A(\counter.cnt_x_digits[4] ));
 sg13g2_inv_2 _1316_ (.Y(_0549_),
    .A(\counter.cnt_x_digits[3] ));
 sg13g2_inv_1 _1317_ (.Y(_0550_),
    .A(\counter.cnt_x_digits[2] ));
 sg13g2_inv_1 _1318_ (.Y(_0551_),
    .A(\counter.cnt_x_digits[1] ));
 sg13g2_inv_1 _1319_ (.Y(_0552_),
    .A(\counter.cnt_x_digits[0] ));
 sg13g2_inv_1 _1320_ (.Y(_0553_),
    .A(net164));
 sg13g2_inv_1 _1321_ (.Y(_0554_),
    .A(net286));
 sg13g2_inv_1 _1322_ (.Y(_0555_),
    .A(\counter.cnt_x_digits[23] ));
 sg13g2_inv_1 _1323_ (.Y(_0556_),
    .A(\counter.cnt_x_digits[22] ));
 sg13g2_inv_1 _1324_ (.Y(_0557_),
    .A(\counter.cnt_x_digits[21] ));
 sg13g2_inv_1 _1325_ (.Y(_0558_),
    .A(\counter.cnt_x_digits[20] ));
 sg13g2_inv_2 _1326_ (.Y(_0559_),
    .A(net246));
 sg13g2_inv_1 _1327_ (.Y(_0560_),
    .A(\counter.streamer.graphical_decoder.index_y_in[0] ));
 sg13g2_inv_1 _1328_ (.Y(_0561_),
    .A(net431));
 sg13g2_inv_1 _1329_ (.Y(_0562_),
    .A(\counter.streamer.digit_cnt_r[2] ));
 sg13g2_inv_2 _1330_ (.Y(_0563_),
    .A(\counter.oled_driver.ready_out ));
 sg13g2_inv_1 _1331_ (.Y(_0564_),
    .A(_0033_));
 sg13g2_inv_1 _1332_ (.Y(\counter.oled_driver.mc_exec.reset_in ),
    .A(net276));
 sg13g2_inv_1 _1333_ (.Y(_0565_),
    .A(net401));
 sg13g2_inv_1 _1334_ (.Y(_0566_),
    .A(net357));
 sg13g2_inv_1 _1335_ (.Y(_0567_),
    .A(_0034_));
 sg13g2_inv_2 _1336_ (.Y(_0568_),
    .A(_0035_));
 sg13g2_inv_2 _1337_ (.Y(_0569_),
    .A(_0036_));
 sg13g2_inv_1 _1338_ (.Y(_0570_),
    .A(_0037_));
 sg13g2_inv_2 _1339_ (.Y(_0571_),
    .A(net258));
 sg13g2_inv_1 _1340_ (.Y(_0572_),
    .A(\counter.oled_driver.mc_exec.state_r[3] ));
 sg13g2_inv_1 _1341_ (.Y(_0573_),
    .A(net296));
 sg13g2_inv_1 _1342_ (.Y(_0574_),
    .A(net360));
 sg13g2_inv_1 _1343_ (.Y(_0575_),
    .A(net354));
 sg13g2_inv_1 _1344_ (.Y(_0576_),
    .A(\counter.oled_driver.state_r[0] ));
 sg13g2_inv_1 _1345_ (.Y(_0577_),
    .A(net186));
 sg13g2_inv_1 _1346_ (.Y(_0578_),
    .A(\counter.oled_driver.spi_deactivate_cs ));
 sg13g2_inv_1 _1347_ (.Y(_0579_),
    .A(net184));
 sg13g2_inv_2 _1348_ (.Y(_0580_),
    .A(_0066_));
 sg13g2_inv_1 _1349_ (.Y(_0581_),
    .A(_0077_));
 sg13g2_inv_1 _1350_ (.Y(_0582_),
    .A(_0043_));
 sg13g2_inv_1 _1351_ (.Y(_0583_),
    .A(_0044_));
 sg13g2_inv_1 _1352_ (.Y(_0584_),
    .A(_0045_));
 sg13g2_inv_1 _1353_ (.Y(_0585_),
    .A(_0052_));
 sg13g2_nand2_1 _1354_ (.Y(_0586_),
    .A(net260),
    .B(\counter.cnt_x_digits[0] ));
 sg13g2_nor4_2 _1355_ (.A(_0549_),
    .B(\counter.cnt_x_digits[2] ),
    .C(\counter.cnt_x_digits[1] ),
    .Y(_0587_),
    .D(_0586_));
 sg13g2_and2_1 _1356_ (.A(\counter.cnt_x_digits[4] ),
    .B(_0587_),
    .X(_0588_));
 sg13g2_nand2_1 _1357_ (.Y(_0589_),
    .A(\counter.cnt_x_digits[7] ),
    .B(_0546_));
 sg13g2_and4_2 _1358_ (.A(\counter.cnt_x_digits[7] ),
    .B(_0546_),
    .C(_0547_),
    .D(_0588_),
    .X(_0590_));
 sg13g2_and2_1 _1359_ (.A(\counter.cnt_x_digits[8] ),
    .B(_0590_),
    .X(_0591_));
 sg13g2_nand2_2 _1360_ (.Y(_0592_),
    .A(\counter.cnt_x_digits[8] ),
    .B(_0590_));
 sg13g2_nand2_2 _1361_ (.Y(_0593_),
    .A(\counter.cnt_x_digits[11] ),
    .B(_0542_));
 sg13g2_nor4_2 _1362_ (.A(_0540_),
    .B(\counter.cnt_x_digits[9] ),
    .C(_0592_),
    .Y(_0594_),
    .D(_0593_));
 sg13g2_inv_1 _1363_ (.Y(_0595_),
    .A(_0594_));
 sg13g2_nand2_2 _1364_ (.Y(_0596_),
    .A(\counter.cnt_x_digits[15] ),
    .B(_0538_));
 sg13g2_nor3_2 _1365_ (.A(\counter.cnt_x_digits[13] ),
    .B(_0595_),
    .C(_0596_),
    .Y(_0597_));
 sg13g2_and2_1 _1366_ (.A(\counter.cnt_x_digits[16] ),
    .B(_0597_),
    .X(_0598_));
 sg13g2_nor3_2 _1367_ (.A(\counter.cnt_x_digits[9] ),
    .B(_0592_),
    .C(_0593_),
    .Y(_0599_));
 sg13g2_nand2_1 _1368_ (.Y(_0600_),
    .A(\counter.cnt_x_digits[12] ),
    .B(_0599_));
 sg13g2_nor3_2 _1369_ (.A(\counter.cnt_x_digits[13] ),
    .B(_0596_),
    .C(_0600_),
    .Y(_0601_));
 sg13g2_nand2_1 _1370_ (.Y(_0602_),
    .A(\counter.cnt_x_digits[16] ),
    .B(_0601_));
 sg13g2_nand4_1 _1371_ (.B(\counter.cnt_x_digits[17] ),
    .C(\counter.cnt_x_digits[16] ),
    .A(\counter.cnt_x_digits[18] ),
    .Y(_0603_),
    .D(_0601_));
 sg13g2_nand2_1 _1372_ (.Y(_0604_),
    .A(\counter.cnt_x_digits[19] ),
    .B(_0534_));
 sg13g2_nor3_2 _1373_ (.A(\counter.cnt_x_digits[17] ),
    .B(_0602_),
    .C(_0604_),
    .Y(_0605_));
 sg13g2_xnor2_1 _1374_ (.Y(_0606_),
    .A(_0533_),
    .B(_0603_));
 sg13g2_nor2_1 _1375_ (.A(_0605_),
    .B(_0606_),
    .Y(_0212_));
 sg13g2_o21ai_1 _1376_ (.B1(_0534_),
    .Y(_0607_),
    .A1(_0535_),
    .A2(_0602_));
 sg13g2_and2_1 _1377_ (.A(_0603_),
    .B(_0607_),
    .X(_0211_));
 sg13g2_a21oi_1 _1378_ (.A1(_0598_),
    .A2(_0604_),
    .Y(_0608_),
    .B1(\counter.cnt_x_digits[17] ));
 sg13g2_a21oi_1 _1379_ (.A1(\counter.cnt_x_digits[17] ),
    .A2(_0598_),
    .Y(_0210_),
    .B1(_0608_));
 sg13g2_xnor2_1 _1380_ (.Y(_0209_),
    .A(_0536_),
    .B(_0597_));
 sg13g2_nand4_1 _1381_ (.B(\counter.cnt_x_digits[13] ),
    .C(\counter.cnt_x_digits[12] ),
    .A(\counter.cnt_x_digits[14] ),
    .Y(_0609_),
    .D(_0599_));
 sg13g2_xnor2_1 _1382_ (.Y(_0610_),
    .A(_0537_),
    .B(_0609_));
 sg13g2_nor2_1 _1383_ (.A(_0601_),
    .B(_0610_),
    .Y(_0208_));
 sg13g2_o21ai_1 _1384_ (.B1(_0538_),
    .Y(_0611_),
    .A1(_0539_),
    .A2(_0595_));
 sg13g2_and2_1 _1385_ (.A(_0609_),
    .B(_0611_),
    .X(_0207_));
 sg13g2_a21oi_1 _1386_ (.A1(_0594_),
    .A2(_0596_),
    .Y(_0612_),
    .B1(\counter.cnt_x_digits[13] ));
 sg13g2_a21oi_1 _1387_ (.A1(\counter.cnt_x_digits[13] ),
    .A2(_0594_),
    .Y(_0206_),
    .B1(_0612_));
 sg13g2_xnor2_1 _1388_ (.Y(_0205_),
    .A(_0540_),
    .B(_0599_));
 sg13g2_nor2_1 _1389_ (.A(_0543_),
    .B(_0592_),
    .Y(_0613_));
 sg13g2_nand2_1 _1390_ (.Y(_0614_),
    .A(\counter.cnt_x_digits[10] ),
    .B(_0613_));
 sg13g2_xnor2_1 _1391_ (.Y(_0615_),
    .A(_0541_),
    .B(_0614_));
 sg13g2_nor2_1 _1392_ (.A(_0599_),
    .B(_0615_),
    .Y(_0204_));
 sg13g2_xnor2_1 _1393_ (.Y(_0203_),
    .A(_0542_),
    .B(_0613_));
 sg13g2_a21oi_1 _1394_ (.A1(_0591_),
    .A2(_0593_),
    .Y(_0616_),
    .B1(\counter.cnt_x_digits[9] ));
 sg13g2_nor2_1 _1395_ (.A(_0613_),
    .B(_0616_),
    .Y(_0202_));
 sg13g2_xnor2_1 _1396_ (.Y(_0201_),
    .A(_0544_),
    .B(_0590_));
 sg13g2_nand3_1 _1397_ (.B(\counter.cnt_x_digits[5] ),
    .C(_0588_),
    .A(\counter.cnt_x_digits[6] ),
    .Y(_0617_));
 sg13g2_xnor2_1 _1398_ (.Y(_0618_),
    .A(_0545_),
    .B(_0617_));
 sg13g2_nor2_1 _1399_ (.A(_0590_),
    .B(_0618_),
    .Y(_0200_));
 sg13g2_a21o_1 _1400_ (.A2(_0588_),
    .A1(\counter.cnt_x_digits[5] ),
    .B1(\counter.cnt_x_digits[6] ),
    .X(_0619_));
 sg13g2_and2_1 _1401_ (.A(_0617_),
    .B(_0619_),
    .X(_0199_));
 sg13g2_a21oi_1 _1402_ (.A1(_0588_),
    .A2(_0589_),
    .Y(_0620_),
    .B1(\counter.cnt_x_digits[5] ));
 sg13g2_a21oi_1 _1403_ (.A1(\counter.cnt_x_digits[5] ),
    .A2(_0588_),
    .Y(_0198_),
    .B1(_0620_));
 sg13g2_xnor2_1 _1404_ (.Y(_0197_),
    .A(_0548_),
    .B(_0587_));
 sg13g2_nor2_1 _1405_ (.A(_0551_),
    .B(_0586_),
    .Y(_0621_));
 sg13g2_nand2_1 _1406_ (.Y(_0622_),
    .A(\counter.cnt_x_digits[2] ),
    .B(_0621_));
 sg13g2_xnor2_1 _1407_ (.Y(_0623_),
    .A(_0549_),
    .B(_0622_));
 sg13g2_nor2_1 _1408_ (.A(_0587_),
    .B(_0623_),
    .Y(_0196_));
 sg13g2_xnor2_1 _1409_ (.Y(_0195_),
    .A(_0550_),
    .B(_0621_));
 sg13g2_a21oi_1 _1410_ (.A1(net260),
    .A2(\counter.cnt_x_digits[0] ),
    .Y(_0624_),
    .B1(\counter.cnt_x_digits[1] ));
 sg13g2_nor3_1 _1411_ (.A(_0587_),
    .B(_0621_),
    .C(_0624_),
    .Y(_0194_));
 sg13g2_xor2_1 _1412_ (.B(\counter.cnt_x_digits[0] ),
    .A(net260),
    .X(_0193_));
 sg13g2_xor2_1 _1413_ (.B(\counter.cnt_x_digits[21] ),
    .A(\counter.cnt_x_digits[22] ),
    .X(_0625_));
 sg13g2_nand2_2 _1414_ (.Y(_0626_),
    .A(\counter.cnt_x_digits[20] ),
    .B(_0605_));
 sg13g2_nor2_1 _1415_ (.A(_0625_),
    .B(_0626_),
    .Y(_0627_));
 sg13g2_o21ai_1 _1416_ (.B1(\counter.cnt_x_digits[23] ),
    .Y(_0628_),
    .A1(_0625_),
    .A2(_0626_));
 sg13g2_nand4_1 _1417_ (.B(\counter.cnt_x_digits[21] ),
    .C(\counter.cnt_x_digits[20] ),
    .A(\counter.cnt_x_digits[22] ),
    .Y(_0629_),
    .D(_0605_));
 sg13g2_o21ai_1 _1418_ (.B1(_0628_),
    .Y(_0106_),
    .A1(\counter.cnt_x_digits[23] ),
    .A2(_0629_));
 sg13g2_a21oi_1 _1419_ (.A1(_0556_),
    .A2(_0626_),
    .Y(_0105_),
    .B1(_0627_));
 sg13g2_a21oi_1 _1420_ (.A1(\counter.cnt_x_digits[23] ),
    .A2(_0556_),
    .Y(_0630_),
    .B1(\counter.cnt_x_digits[21] ));
 sg13g2_mux2_1 _1421_ (.A0(_0630_),
    .A1(\counter.cnt_x_digits[21] ),
    .S(_0626_),
    .X(_0104_));
 sg13g2_xnor2_1 _1422_ (.Y(_0103_),
    .A(_0558_),
    .B(_0605_));
 sg13g2_nand2_1 _1423_ (.Y(_0631_),
    .A(net278),
    .B(\counter.oled_driver.mc_exec.state_r[2] ));
 sg13g2_a21o_2 _1424_ (.A2(\counter.oled_driver.mc_exec.microcode_rom.address[2] ),
    .A1(\counter.oled_driver.mc_exec.microcode_rom.address[3] ),
    .B1(\counter.oled_driver.mc_exec.microcode_rom.address[4] ),
    .X(_0632_));
 sg13g2_nand2_1 _1425_ (.Y(_0633_),
    .A(\counter.oled_driver.mc_exec.microcode_rom.address[5] ),
    .B(_0632_));
 sg13g2_and2_2 _1426_ (.A(_0042_),
    .B(net229),
    .X(_0634_));
 sg13g2_nand2_2 _1427_ (.Y(_0635_),
    .A(_0042_),
    .B(net229));
 sg13g2_nand2b_1 _1428_ (.Y(_0636_),
    .B(_0634_),
    .A_N(_0631_));
 sg13g2_nor2_1 _1429_ (.A(_0040_),
    .B(_0636_),
    .Y(_0637_));
 sg13g2_nand2_2 _1430_ (.Y(_0638_),
    .A(_0033_),
    .B(net230));
 sg13g2_and2_2 _1431_ (.A(_0038_),
    .B(_0633_),
    .X(_0639_));
 sg13g2_nand2_1 _1432_ (.Y(_0640_),
    .A(_0038_),
    .B(net229));
 sg13g2_a21oi_2 _1433_ (.B1(_0570_),
    .Y(_0641_),
    .A2(_0632_),
    .A1(net245));
 sg13g2_nor4_1 _1434_ (.A(_0034_),
    .B(_0037_),
    .C(_0638_),
    .D(_0639_),
    .Y(_0642_));
 sg13g2_a21oi_2 _1435_ (.B1(_0569_),
    .Y(_0643_),
    .A2(_0632_),
    .A1(\counter.oled_driver.mc_exec.microcode_rom.address[5] ));
 sg13g2_a21oi_2 _1436_ (.B1(_0568_),
    .Y(_0644_),
    .A2(_0632_),
    .A1(net245));
 sg13g2_a21o_1 _1437_ (.A2(_0632_),
    .A1(\counter.oled_driver.mc_exec.microcode_rom.address[5] ),
    .B1(_0568_),
    .X(_0645_));
 sg13g2_nor2_1 _1438_ (.A(_0643_),
    .B(_0644_),
    .Y(_0646_));
 sg13g2_a22oi_1 _1439_ (.Y(_0647_),
    .B1(_0632_),
    .B2(net245),
    .A2(_0569_),
    .A1(_0568_));
 sg13g2_nand2_2 _1440_ (.Y(_0648_),
    .A(_0039_),
    .B(net230));
 sg13g2_nand2_1 _1441_ (.Y(_0649_),
    .A(_0040_),
    .B(net230));
 sg13g2_o21ai_1 _1442_ (.B1(net229),
    .Y(_0650_),
    .A1(_0040_),
    .A2(_0039_));
 sg13g2_nand3_1 _1443_ (.B(_0646_),
    .C(_0650_),
    .A(_0642_),
    .Y(_0651_));
 sg13g2_or3_1 _1444_ (.A(_0040_),
    .B(_0636_),
    .C(_0651_),
    .X(_0652_));
 sg13g2_nand4_1 _1445_ (.B(net278),
    .C(net441),
    .A(net245),
    .Y(_0653_),
    .D(_0632_));
 sg13g2_nand2_1 _1446_ (.Y(_0654_),
    .A(net271),
    .B(net257));
 sg13g2_a21oi_1 _1447_ (.A1(\counter.oled_driver.spi_driver.state_r[0] ),
    .A2(net357),
    .Y(_0655_),
    .B1(_0654_));
 sg13g2_a21oi_1 _1448_ (.A1(net271),
    .A2(net320),
    .Y(_0656_),
    .B1(_0655_));
 sg13g2_nand3_1 _1449_ (.B(net442),
    .C(_0656_),
    .A(_0652_),
    .Y(_0019_));
 sg13g2_and2_1 _1450_ (.A(net270),
    .B(\counter.oled_driver.spi_driver.state_r[0] ),
    .X(_0657_));
 sg13g2_nand2_1 _1451_ (.Y(_0658_),
    .A(net270),
    .B(\counter.oled_driver.spi_driver.state_r[0] ));
 sg13g2_nand2_1 _1452_ (.Y(_0659_),
    .A(net296),
    .B(_0657_));
 sg13g2_nor2_2 _1453_ (.A(_0563_),
    .B(net265),
    .Y(_0660_));
 sg13g2_nand3_1 _1454_ (.B(_0575_),
    .C(_0660_),
    .A(_0574_),
    .Y(_0661_));
 sg13g2_nand3_1 _1455_ (.B(net257),
    .C(net397),
    .A(net270),
    .Y(_0662_));
 sg13g2_nand3_1 _1456_ (.B(_0661_),
    .C(_0662_),
    .A(_0659_),
    .Y(_0026_));
 sg13g2_nor2_1 _1457_ (.A(net379),
    .B(_0658_),
    .Y(_0663_));
 sg13g2_nand2_1 _1458_ (.Y(_0664_),
    .A(net354),
    .B(_0660_));
 sg13g2_a22oi_1 _1459_ (.Y(_0665_),
    .B1(_0663_),
    .B2(\counter.oled_driver.state_r[0] ),
    .A2(_0660_),
    .A1(net354));
 sg13g2_o21ai_1 _1460_ (.B1(_0665_),
    .Y(_0025_),
    .A1(_0566_),
    .A2(_0654_));
 sg13g2_and3_1 _1461_ (.X(_0666_),
    .A(_0570_),
    .B(_0639_),
    .C(_0650_));
 sg13g2_a22oi_1 _1462_ (.Y(_0667_),
    .B1(_0632_),
    .B2(net245),
    .A2(_0567_),
    .A1(_0564_));
 sg13g2_or2_1 _1463_ (.X(_0668_),
    .B(_0667_),
    .A(_0647_));
 sg13g2_nor3_1 _1464_ (.A(_0641_),
    .B(_0647_),
    .C(_0667_),
    .Y(_0669_));
 sg13g2_and2_1 _1465_ (.A(_0640_),
    .B(_0669_),
    .X(_0670_));
 sg13g2_a21oi_1 _1466_ (.A1(_0650_),
    .A2(_0670_),
    .Y(_0671_),
    .B1(_0666_));
 sg13g2_a21oi_1 _1467_ (.A1(_0649_),
    .A2(_0671_),
    .Y(_0672_),
    .B1(_0636_));
 sg13g2_nor2_1 _1468_ (.A(net369),
    .B(\counter.oled_driver.mc_exec.delay_cnt[0] ),
    .Y(_0673_));
 sg13g2_nor4_2 _1469_ (.A(net343),
    .B(net284),
    .C(net369),
    .Y(_0674_),
    .D(\counter.oled_driver.mc_exec.delay_cnt[0] ));
 sg13g2_inv_1 _1470_ (.Y(_0675_),
    .A(_0674_));
 sg13g2_nor3_2 _1471_ (.A(\counter.oled_driver.mc_exec.delay_cnt[5] ),
    .B(net189),
    .C(_0675_),
    .Y(_0676_));
 sg13g2_nor2_1 _1472_ (.A(\counter.oled_driver.mc_exec.delay_cnt[7] ),
    .B(\counter.oled_driver.mc_exec.delay_cnt[6] ),
    .Y(_0677_));
 sg13g2_nand2_1 _1473_ (.Y(_0678_),
    .A(_0676_),
    .B(_0677_));
 sg13g2_or3_1 _1474_ (.A(\counter.oled_driver.mc_exec.delay_cnt[9] ),
    .B(\counter.oled_driver.mc_exec.delay_cnt[8] ),
    .C(_0678_),
    .X(_0679_));
 sg13g2_nor3_1 _1475_ (.A(\counter.oled_driver.mc_exec.delay_cnt[11] ),
    .B(net174),
    .C(_0679_),
    .Y(_0680_));
 sg13g2_nor2b_1 _1476_ (.A(\counter.oled_driver.mc_exec.delay_cnt[12] ),
    .B_N(_0680_),
    .Y(_0681_));
 sg13g2_nor2b_2 _1477_ (.A(net204),
    .B_N(_0681_),
    .Y(_0682_));
 sg13g2_nor2_1 _1478_ (.A(\counter.oled_driver.mc_exec.delay_cnt[15] ),
    .B(\counter.oled_driver.mc_exec.delay_cnt[14] ),
    .Y(_0683_));
 sg13g2_nand3_1 _1479_ (.B(_0682_),
    .C(_0683_),
    .A(net306),
    .Y(_0684_));
 sg13g2_nand2_1 _1480_ (.Y(_0685_),
    .A(net271),
    .B(net372));
 sg13g2_a21oi_1 _1481_ (.A1(net198),
    .A2(_0657_),
    .Y(_0686_),
    .B1(_0672_));
 sg13g2_o21ai_1 _1482_ (.B1(_0686_),
    .Y(_0018_),
    .A1(net307),
    .A2(_0685_));
 sg13g2_nand2_1 _1483_ (.Y(_0687_),
    .A(net206),
    .B(_0657_));
 sg13g2_o21ai_1 _1484_ (.B1(net207),
    .Y(_0016_),
    .A1(_0631_),
    .A2(_0634_));
 sg13g2_nand4_1 _1485_ (.B(_0648_),
    .C(_0651_),
    .A(_0637_),
    .Y(_0688_),
    .D(_0671_));
 sg13g2_nand3_1 _1486_ (.B(net441),
    .C(net230),
    .A(net271),
    .Y(_0689_));
 sg13g2_nand4_1 _1487_ (.B(net449),
    .C(net357),
    .A(net270),
    .Y(_0690_),
    .D(net257));
 sg13g2_nand3_1 _1488_ (.B(_0689_),
    .C(_0690_),
    .A(_0688_),
    .Y(_0017_));
 sg13g2_nand2_1 _1489_ (.Y(_0691_),
    .A(net360),
    .B(_0660_));
 sg13g2_o21ai_1 _1490_ (.B1(_0691_),
    .Y(_0024_),
    .A1(_0578_),
    .A2(_0658_));
 sg13g2_nand2b_1 _1491_ (.Y(_0692_),
    .B(\counter.streamer.ready_out ),
    .A_N(\counter.refresh_display ));
 sg13g2_nand3_1 _1492_ (.B(net186),
    .C(_0692_),
    .A(net273),
    .Y(_0693_));
 sg13g2_nor2b_1 _1493_ (.A(net359),
    .B_N(net353),
    .Y(_0694_));
 sg13g2_nor2b_1 _1494_ (.A(net201),
    .B_N(\counter.counter_ref.digits_out[11] ),
    .Y(_0695_));
 sg13g2_and2_1 _1495_ (.A(_0694_),
    .B(_0695_),
    .X(_0696_));
 sg13g2_nand2b_1 _1496_ (.Y(_0697_),
    .B(net191),
    .A_N(\counter.counter_ref.digits_out[6] ));
 sg13g2_nor3_2 _1497_ (.A(\counter.counter_ref.digits_out[5] ),
    .B(_0532_),
    .C(_0697_),
    .Y(_0698_));
 sg13g2_nand2b_1 _1498_ (.Y(_0699_),
    .B(net273),
    .A_N(net179));
 sg13g2_inv_2 _1499_ (.Y(_0079_),
    .A(net243));
 sg13g2_nand2_1 _1500_ (.Y(_0700_),
    .A(\counter.counter_ref.digit_0.digit_out[3] ),
    .B(\counter.counter_ref.digit_0.digit_out[0] ));
 sg13g2_nor3_2 _1501_ (.A(\counter.counter_ref.digit_0.digit_out[2] ),
    .B(net464),
    .C(_0700_),
    .Y(_0701_));
 sg13g2_nand2_1 _1502_ (.Y(_0702_),
    .A(net259),
    .B(net465));
 sg13g2_nor2_1 _1503_ (.A(net239),
    .B(_0702_),
    .Y(_0703_));
 sg13g2_and4_1 _1504_ (.A(net259),
    .B(_0698_),
    .C(net228),
    .D(_0701_),
    .X(_0704_));
 sg13g2_and2_1 _1505_ (.A(_0696_),
    .B(_0704_),
    .X(_0705_));
 sg13g2_nand2b_1 _1506_ (.Y(_0706_),
    .B(\counter.counter_ref.digits_out[16] ),
    .A_N(\counter.counter_ref.digits_out[17] ));
 sg13g2_nor3_1 _1507_ (.A(\counter.counter_ref.digits_out[13] ),
    .B(_0531_),
    .C(_0706_),
    .Y(_0707_));
 sg13g2_nand2b_1 _1508_ (.Y(_0708_),
    .B(\counter.counter_ref.digits_out[23] ),
    .A_N(net323));
 sg13g2_nand2b_2 _1509_ (.Y(_0709_),
    .B(net288),
    .A_N(net439));
 sg13g2_nor2_1 _1510_ (.A(_0708_),
    .B(_0709_),
    .Y(_0710_));
 sg13g2_nand2b_2 _1511_ (.Y(_0711_),
    .B(\counter.counter_ref.digits_out[19] ),
    .A_N(\counter.counter_ref.digits_out[18] ));
 sg13g2_nor3_1 _1512_ (.A(\counter.counter_ref.digits_out[21] ),
    .B(_0529_),
    .C(_0711_),
    .Y(_0712_));
 sg13g2_and4_1 _1513_ (.A(_0705_),
    .B(_0707_),
    .C(_0710_),
    .D(_0712_),
    .X(_0713_));
 sg13g2_and3_1 _1514_ (.X(_0714_),
    .A(_0694_),
    .B(_0695_),
    .C(net228));
 sg13g2_and4_1 _1515_ (.A(net259),
    .B(_0698_),
    .C(_0701_),
    .D(_0714_),
    .X(_0715_));
 sg13g2_nor4_1 _1516_ (.A(\counter.counter_ref.digits_out[21] ),
    .B(_0529_),
    .C(\counter.counter_ref.digits_out[13] ),
    .D(_0531_),
    .Y(_0716_));
 sg13g2_nand2_1 _1517_ (.Y(_0717_),
    .A(_0710_),
    .B(_0716_));
 sg13g2_nor3_2 _1518_ (.A(_0706_),
    .B(_0711_),
    .C(_0717_),
    .Y(_0718_));
 sg13g2_nand2_1 _1519_ (.Y(_0719_),
    .A(_0715_),
    .B(_0718_));
 sg13g2_and4_1 _1520_ (.A(_0696_),
    .B(_0698_),
    .C(net227),
    .D(_0701_),
    .X(_0720_));
 sg13g2_nand2_1 _1521_ (.Y(_0028_),
    .A(net187),
    .B(_0719_));
 sg13g2_or2_1 _1522_ (.X(_0721_),
    .B(_0692_),
    .A(net261));
 sg13g2_a21o_1 _1523_ (.A2(\counter.streamer.ready_out ),
    .A1(net273),
    .B1(_0079_),
    .X(_0722_));
 sg13g2_o21ai_1 _1524_ (.B1(_0722_),
    .Y(_0027_),
    .A1(net166),
    .A2(_0721_));
 sg13g2_a21oi_1 _1525_ (.A1(net270),
    .A2(_0576_),
    .Y(_0023_),
    .B1(net380));
 sg13g2_nor3_1 _1526_ (.A(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[2] ),
    .B(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[1] ),
    .C(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[0] ),
    .Y(_0723_));
 sg13g2_nor2b_2 _1527_ (.A(net388),
    .B_N(_0723_),
    .Y(_0724_));
 sg13g2_nand2_1 _1528_ (.Y(_0725_),
    .A(net280),
    .B(_0724_));
 sg13g2_nor2b_1 _1529_ (.A(net253),
    .B_N(\counter.oled_driver.mc_exec.spi_tx_trigger_out ),
    .Y(_0726_));
 sg13g2_a21oi_1 _1530_ (.A1(net254),
    .A2(\counter.oled_driver.spi_deactivate_cs ),
    .Y(_0727_),
    .B1(_0726_));
 sg13g2_nor2_1 _1531_ (.A(net226),
    .B(_0727_),
    .Y(_0728_));
 sg13g2_nand2_1 _1532_ (.Y(_0729_),
    .A(net449),
    .B(_0728_));
 sg13g2_nand3_1 _1533_ (.B(net364),
    .C(_0724_),
    .A(net280),
    .Y(_0730_));
 sg13g2_nand2_1 _1534_ (.Y(_0022_),
    .A(_0729_),
    .B(net225));
 sg13g2_nand2_1 _1535_ (.Y(_0731_),
    .A(net401),
    .B(_0660_));
 sg13g2_nor3_1 _1536_ (.A(\counter.streamer.graphical_decoder.index_x_in[3] ),
    .B(net248),
    .C(\counter.streamer.graphical_decoder.index_x_in[0] ),
    .Y(_0732_));
 sg13g2_nand3_1 _1537_ (.B(\counter.streamer.graphical_decoder.index_x_in[2] ),
    .C(_0732_),
    .A(\counter.streamer.graphical_decoder.index_x_in[4] ),
    .Y(_0733_));
 sg13g2_nand2_2 _1538_ (.Y(_0734_),
    .A(net247),
    .B(\counter.streamer.graphical_decoder.index_y_in[0] ));
 sg13g2_nor2_1 _1539_ (.A(net249),
    .B(net251),
    .Y(_0735_));
 sg13g2_nor3_1 _1540_ (.A(\counter.streamer.digit_cnt_r[2] ),
    .B(net249),
    .C(net251),
    .Y(_0736_));
 sg13g2_nor2b_1 _1541_ (.A(_0733_),
    .B_N(_0736_),
    .Y(_0737_));
 sg13g2_nand2b_1 _1542_ (.Y(_0738_),
    .B(_0737_),
    .A_N(_0734_));
 sg13g2_o21ai_1 _1543_ (.B1(_0664_),
    .Y(_0030_),
    .A1(_0731_),
    .A2(_0738_));
 sg13g2_nand2_1 _1544_ (.Y(_0739_),
    .A(net347),
    .B(net389));
 sg13g2_nand2b_2 _1545_ (.Y(_0740_),
    .B(net280),
    .A_N(\counter.oled_driver.spi_driver.state_r[0] ));
 sg13g2_inv_1 _1546_ (.Y(_0741_),
    .A(_0740_));
 sg13g2_o21ai_1 _1547_ (.B1(_0739_),
    .Y(_0021_),
    .A1(_0728_),
    .A2(_0741_));
 sg13g2_nand3_1 _1548_ (.B(\counter.streamer.ready_out ),
    .C(net179),
    .A(net273),
    .Y(_0742_));
 sg13g2_nand2_1 _1549_ (.Y(_0743_),
    .A(net260),
    .B(net273));
 sg13g2_and4_1 _1550_ (.A(_0698_),
    .B(_0701_),
    .C(_0714_),
    .D(_0718_),
    .X(_0744_));
 sg13g2_o21ai_1 _1551_ (.B1(net180),
    .Y(_0029_),
    .A1(_0743_),
    .A2(_0744_));
 sg13g2_nand2b_1 _1552_ (.Y(_0745_),
    .B(_0738_),
    .A_N(_0731_));
 sg13g2_and2_1 _1553_ (.A(\counter.refresh_display ),
    .B(\counter.streamer.ready_out ),
    .X(_0746_));
 sg13g2_nand2_1 _1554_ (.Y(_0747_),
    .A(net273),
    .B(net235));
 sg13g2_nand3_1 _1555_ (.B(_0745_),
    .C(_0747_),
    .A(_0691_),
    .Y(_0031_));
 sg13g2_nor4_2 _1556_ (.A(_0040_),
    .B(_0571_),
    .C(_0635_),
    .Y(_0748_),
    .D(_0648_));
 sg13g2_a21oi_1 _1557_ (.A1(net372),
    .A2(_0684_),
    .Y(_0749_),
    .B1(_0748_));
 sg13g2_nor2_1 _1558_ (.A(net261),
    .B(net373),
    .Y(_0020_));
 sg13g2_a22oi_1 _1559_ (.Y(_0750_),
    .B1(net184),
    .B2(_0660_),
    .A2(net320),
    .A1(net276));
 sg13g2_nand2_1 _1560_ (.Y(_0032_),
    .A(_0721_),
    .B(_0750_));
 sg13g2_nand3b_1 _1561_ (.B(_0634_),
    .C(_0040_),
    .Y(_0751_),
    .A_N(_0056_));
 sg13g2_o21ai_1 _1562_ (.B1(_0643_),
    .Y(_0752_),
    .A1(_0644_),
    .A2(_0667_));
 sg13g2_xnor2_1 _1563_ (.Y(_0753_),
    .A(_0645_),
    .B(_0667_));
 sg13g2_a21oi_1 _1564_ (.A1(_0668_),
    .A2(_0752_),
    .Y(_0754_),
    .B1(_0753_));
 sg13g2_xnor2_1 _1565_ (.Y(_0755_),
    .A(_0641_),
    .B(_0668_));
 sg13g2_xnor2_1 _1566_ (.Y(_0756_),
    .A(_0640_),
    .B(_0669_));
 sg13g2_o21ai_1 _1567_ (.B1(_0756_),
    .Y(_0757_),
    .A1(_0754_),
    .A2(_0755_));
 sg13g2_xor2_1 _1568_ (.B(_0670_),
    .A(_0648_),
    .X(_0758_));
 sg13g2_a21oi_1 _1569_ (.A1(_0757_),
    .A2(_0758_),
    .Y(_0759_),
    .B1(_0751_));
 sg13g2_a21o_1 _1570_ (.A2(_0758_),
    .A1(_0757_),
    .B1(_0751_),
    .X(_0760_));
 sg13g2_nor3_1 _1571_ (.A(_0040_),
    .B(_0056_),
    .C(_0635_),
    .Y(_0761_));
 sg13g2_nor2_2 _1572_ (.A(\counter.oled_driver.mc_exec.state_r[0] ),
    .B(net258),
    .Y(_0762_));
 sg13g2_nor3_1 _1573_ (.A(\counter.oled_driver.mc_exec.state_r[0] ),
    .B(net258),
    .C(\counter.oled_driver.mc_exec.state_r[3] ),
    .Y(_0763_));
 sg13g2_o21ai_1 _1574_ (.B1(_0690_),
    .Y(_0764_),
    .A1(net257),
    .A2(_0763_));
 sg13g2_o21ai_1 _1575_ (.B1(_0764_),
    .Y(_0765_),
    .A1(_0057_),
    .A2(net230));
 sg13g2_a21oi_1 _1576_ (.A1(\counter.oled_driver.mc_exec.state_r[2] ),
    .A2(_0635_),
    .Y(_0766_),
    .B1(_0765_));
 sg13g2_nor2b_2 _1577_ (.A(_0761_),
    .B_N(_0766_),
    .Y(_0767_));
 sg13g2_inv_1 _1578_ (.Y(_0768_),
    .A(_0767_));
 sg13g2_nor2_2 _1579_ (.A(net221),
    .B(_0768_),
    .Y(_0769_));
 sg13g2_and3_2 _1580_ (.X(_0770_),
    .A(_0571_),
    .B(_0572_),
    .C(_0054_));
 sg13g2_nand3_1 _1581_ (.B(_0572_),
    .C(net379),
    .A(_0571_),
    .Y(_0771_));
 sg13g2_nand2_1 _1582_ (.Y(_0772_),
    .A(\counter.oled_driver.mc_exec.microcode_rom.address[1] ),
    .B(\counter.oled_driver.mc_exec.microcode_rom.address[0] ));
 sg13g2_and4_1 _1583_ (.A(\counter.oled_driver.mc_exec.microcode_rom.address[3] ),
    .B(\counter.oled_driver.mc_exec.microcode_rom.address[2] ),
    .C(\counter.oled_driver.mc_exec.microcode_rom.address[1] ),
    .D(\counter.oled_driver.mc_exec.microcode_rom.address[0] ),
    .X(_0773_));
 sg13g2_a21oi_1 _1584_ (.A1(\counter.oled_driver.mc_exec.microcode_rom.address[4] ),
    .A2(_0773_),
    .Y(_0774_),
    .B1(net245));
 sg13g2_nand3_1 _1585_ (.B(\counter.oled_driver.mc_exec.microcode_rom.address[4] ),
    .C(_0773_),
    .A(net245),
    .Y(_0775_));
 sg13g2_nor2_1 _1586_ (.A(_0572_),
    .B(_0774_),
    .Y(_0776_));
 sg13g2_a22oi_1 _1587_ (.Y(_0777_),
    .B1(_0775_),
    .B2(_0776_),
    .A2(net257),
    .A1(\counter.oled_driver.mc_exec.procedure_offset_in[0] ));
 sg13g2_nor2_1 _1588_ (.A(_0770_),
    .B(_0777_),
    .Y(_0778_));
 sg13g2_a21oi_1 _1589_ (.A1(\counter.oled_driver.mc_exec.state_r[2] ),
    .A2(_0756_),
    .Y(_0779_),
    .B1(_0778_));
 sg13g2_o21ai_1 _1590_ (.B1(net278),
    .Y(_0780_),
    .A1(net245),
    .A2(_0769_));
 sg13g2_a21oi_2 _1591_ (.B1(_0780_),
    .Y(_0168_),
    .A2(_0779_),
    .A1(_0769_));
 sg13g2_inv_2 _1592_ (.Y(_0781_),
    .A(_0168_));
 sg13g2_nor2_1 _1593_ (.A(_0056_),
    .B(_0770_),
    .Y(_0782_));
 sg13g2_a21oi_1 _1594_ (.A1(_0668_),
    .A2(_0752_),
    .Y(_0783_),
    .B1(_0056_));
 sg13g2_nor2_2 _1595_ (.A(_0057_),
    .B(_0770_),
    .Y(_0784_));
 sg13g2_o21ai_1 _1596_ (.B1(_0061_),
    .Y(_0785_),
    .A1(_0060_),
    .A2(_0772_));
 sg13g2_nor3_1 _1597_ (.A(_0060_),
    .B(_0061_),
    .C(_0772_),
    .Y(_0786_));
 sg13g2_nor2_1 _1598_ (.A(_0057_),
    .B(_0786_),
    .Y(_0787_));
 sg13g2_a21oi_1 _1599_ (.A1(_0785_),
    .A2(_0787_),
    .Y(_0788_),
    .B1(_0783_));
 sg13g2_or4_1 _1600_ (.A(net221),
    .B(net220),
    .C(_0770_),
    .D(_0788_),
    .X(_0789_));
 sg13g2_o21ai_1 _1601_ (.B1(_0789_),
    .Y(_0790_),
    .A1(_0061_),
    .A2(_0769_));
 sg13g2_and2_1 _1602_ (.A(net277),
    .B(net219),
    .X(_0791_));
 sg13g2_nand2_2 _1603_ (.Y(_0792_),
    .A(net277),
    .B(net219));
 sg13g2_a22oi_1 _1604_ (.Y(_0793_),
    .B1(net258),
    .B2(_0638_),
    .A2(net257),
    .A1(\counter.oled_driver.mc_exec.procedure_offset_in[0] ));
 sg13g2_o21ai_1 _1605_ (.B1(_0793_),
    .Y(_0794_),
    .A1(\counter.oled_driver.mc_exec.microcode_rom.address[0] ),
    .A2(_0572_));
 sg13g2_nand2_1 _1606_ (.Y(_0795_),
    .A(_0771_),
    .B(_0794_));
 sg13g2_nor3_1 _1607_ (.A(_0759_),
    .B(net220),
    .C(_0795_),
    .Y(_0796_));
 sg13g2_nand3b_1 _1608_ (.B(_0760_),
    .C(_0767_),
    .Y(_0797_),
    .A_N(_0795_));
 sg13g2_a21oi_1 _1609_ (.A1(_0760_),
    .A2(_0767_),
    .Y(_0798_),
    .B1(_0064_));
 sg13g2_or2_2 _1610_ (.X(_0799_),
    .B(_0798_),
    .A(_0796_));
 sg13g2_o21ai_1 _1611_ (.B1(_0667_),
    .Y(_0800_),
    .A1(_0564_),
    .A2(_0567_));
 sg13g2_xor2_1 _1612_ (.B(\counter.oled_driver.mc_exec.microcode_rom.address[0] ),
    .A(\counter.oled_driver.mc_exec.microcode_rom.address[1] ),
    .X(_0801_));
 sg13g2_a22oi_1 _1613_ (.Y(_0802_),
    .B1(_0801_),
    .B2(_0784_),
    .A2(_0800_),
    .A1(net258));
 sg13g2_nor3_2 _1614_ (.A(net221),
    .B(net220),
    .C(_0802_),
    .Y(_0803_));
 sg13g2_nand2b_1 _1615_ (.Y(_0804_),
    .B(_0769_),
    .A_N(_0802_));
 sg13g2_a21oi_2 _1616_ (.B1(_0063_),
    .Y(_0805_),
    .A2(_0767_),
    .A1(_0760_));
 sg13g2_nor2_2 _1617_ (.A(_0803_),
    .B(_0805_),
    .Y(_0806_));
 sg13g2_or2_2 _1618_ (.X(_0807_),
    .B(_0805_),
    .A(_0803_));
 sg13g2_nor2_1 _1619_ (.A(net264),
    .B(_0806_),
    .Y(_0808_));
 sg13g2_o21ai_1 _1620_ (.B1(net278),
    .Y(_0809_),
    .A1(_0803_),
    .A2(_0805_));
 sg13g2_or2_1 _1621_ (.X(_0810_),
    .B(_0809_),
    .A(net218));
 sg13g2_nor2_1 _1622_ (.A(_0571_),
    .B(_0753_),
    .Y(_0811_));
 sg13g2_xor2_1 _1623_ (.B(_0772_),
    .A(_0060_),
    .X(_0812_));
 sg13g2_a21oi_1 _1624_ (.A1(_0784_),
    .A2(_0812_),
    .Y(_0813_),
    .B1(_0811_));
 sg13g2_or3_2 _1625_ (.A(net221),
    .B(net220),
    .C(_0813_),
    .X(_0814_));
 sg13g2_a21o_1 _1626_ (.A2(_0767_),
    .A1(_0760_),
    .B1(_0060_),
    .X(_0815_));
 sg13g2_nand2_2 _1627_ (.Y(_0816_),
    .A(_0814_),
    .B(_0815_));
 sg13g2_nor3_2 _1628_ (.A(net218),
    .B(_0809_),
    .C(_0816_),
    .Y(_0817_));
 sg13g2_o21ai_1 _1629_ (.B1(net278),
    .Y(_0818_),
    .A1(_0796_),
    .A2(_0798_));
 sg13g2_or2_1 _1630_ (.X(_0819_),
    .B(_0818_),
    .A(_0807_));
 sg13g2_or2_1 _1631_ (.X(_0820_),
    .B(_0818_),
    .A(_0816_));
 sg13g2_nor3_2 _1632_ (.A(_0807_),
    .B(_0816_),
    .C(_0818_),
    .Y(_0821_));
 sg13g2_nor2_1 _1633_ (.A(_0817_),
    .B(_0821_),
    .Y(_0822_));
 sg13g2_o21ai_1 _1634_ (.B1(net215),
    .Y(_0823_),
    .A1(_0817_),
    .A2(_0821_));
 sg13g2_a21oi_2 _1635_ (.B1(net264),
    .Y(_0824_),
    .A2(_0815_),
    .A1(_0814_));
 sg13g2_nand2_1 _1636_ (.Y(_0825_),
    .A(net277),
    .B(_0816_));
 sg13g2_nand2_2 _1637_ (.Y(_0826_),
    .A(net218),
    .B(_0824_));
 sg13g2_nand3_1 _1638_ (.B(net218),
    .C(_0824_),
    .A(net219),
    .Y(_0827_));
 sg13g2_nand2_1 _1639_ (.Y(_0828_),
    .A(_0823_),
    .B(_0827_));
 sg13g2_or2_1 _1640_ (.X(_0829_),
    .B(_0769_),
    .A(\counter.oled_driver.mc_exec.microcode_rom.address[4] ));
 sg13g2_xnor2_1 _1641_ (.Y(_0830_),
    .A(_0062_),
    .B(_0773_));
 sg13g2_a22oi_1 _1642_ (.Y(_0831_),
    .B1(_0784_),
    .B2(_0830_),
    .A2(_0782_),
    .A1(_0755_));
 sg13g2_nand2_1 _1643_ (.Y(_0832_),
    .A(_0769_),
    .B(_0831_));
 sg13g2_nand3_1 _1644_ (.B(_0829_),
    .C(_0832_),
    .A(net278),
    .Y(_0833_));
 sg13g2_inv_2 _1645_ (.Y(_0167_),
    .A(net213));
 sg13g2_nand2_2 _1646_ (.Y(_0834_),
    .A(_0792_),
    .B(_0826_));
 sg13g2_nor2_1 _1647_ (.A(_0808_),
    .B(_0824_),
    .Y(_0835_));
 sg13g2_o21ai_1 _1648_ (.B1(net213),
    .Y(_0836_),
    .A1(_0834_),
    .A2(_0835_));
 sg13g2_nor2b_2 _1649_ (.A(net218),
    .B_N(_0824_),
    .Y(_0837_));
 sg13g2_nand2b_1 _1650_ (.Y(_0838_),
    .B(_0824_),
    .A_N(net218));
 sg13g2_nand2b_2 _1651_ (.Y(_0839_),
    .B(_0816_),
    .A_N(_0809_));
 sg13g2_nand3_1 _1652_ (.B(_0819_),
    .C(_0824_),
    .A(_0810_),
    .Y(_0840_));
 sg13g2_nand2b_1 _1653_ (.Y(_0841_),
    .B(_0799_),
    .A_N(_0809_));
 sg13g2_a21o_1 _1654_ (.A2(_0841_),
    .A1(_0825_),
    .B1(net215),
    .X(_0842_));
 sg13g2_nand3_1 _1655_ (.B(_0840_),
    .C(_0842_),
    .A(_0167_),
    .Y(_0843_));
 sg13g2_o21ai_1 _1656_ (.B1(_0843_),
    .Y(_0844_),
    .A1(_0828_),
    .A2(_0836_));
 sg13g2_a21oi_2 _1657_ (.B1(_0824_),
    .Y(_0845_),
    .A2(net218),
    .A1(net277));
 sg13g2_nor2_1 _1658_ (.A(_0781_),
    .B(_0790_),
    .Y(_0846_));
 sg13g2_nor3_1 _1659_ (.A(_0781_),
    .B(_0790_),
    .C(_0845_),
    .Y(_0847_));
 sg13g2_a22oi_1 _1660_ (.Y(_0000_),
    .B1(_0847_),
    .B2(_0840_),
    .A2(_0844_),
    .A1(_0781_));
 sg13g2_nand2_1 _1661_ (.Y(_0848_),
    .A(net219),
    .B(_0807_));
 sg13g2_or2_1 _1662_ (.X(_0849_),
    .B(_0848_),
    .A(_0826_));
 sg13g2_nand2_1 _1663_ (.Y(_0850_),
    .A(_0167_),
    .B(_0849_));
 sg13g2_nor2_1 _1664_ (.A(net214),
    .B(_0817_),
    .Y(_0851_));
 sg13g2_a21oi_1 _1665_ (.A1(_0822_),
    .A2(_0840_),
    .Y(_0852_),
    .B1(_0851_));
 sg13g2_nand4_1 _1666_ (.B(net218),
    .C(_0806_),
    .A(net214),
    .Y(_0853_),
    .D(_0824_));
 sg13g2_nand3_1 _1667_ (.B(_0833_),
    .C(_0853_),
    .A(_0823_),
    .Y(_0854_));
 sg13g2_o21ai_1 _1668_ (.B1(_0854_),
    .Y(_0855_),
    .A1(_0850_),
    .A2(_0852_));
 sg13g2_nand3_1 _1669_ (.B(_0820_),
    .C(_0846_),
    .A(_0810_),
    .Y(_0856_));
 sg13g2_o21ai_1 _1670_ (.B1(_0856_),
    .Y(_0001_),
    .A1(net216),
    .A2(_0855_));
 sg13g2_nor2_1 _1671_ (.A(_0792_),
    .B(_0799_),
    .Y(_0857_));
 sg13g2_nor2_1 _1672_ (.A(_0808_),
    .B(_0834_),
    .Y(_0858_));
 sg13g2_o21ai_1 _1673_ (.B1(_0168_),
    .Y(_0859_),
    .A1(_0857_),
    .A2(_0858_));
 sg13g2_nand3_1 _1674_ (.B(_0806_),
    .C(_0837_),
    .A(net214),
    .Y(_0860_));
 sg13g2_nand4_1 _1675_ (.B(_0827_),
    .C(_0167_),
    .A(_0823_),
    .Y(_0861_),
    .D(_0860_));
 sg13g2_nand2_2 _1676_ (.Y(_0862_),
    .A(_0807_),
    .B(_0837_));
 sg13g2_nand3_1 _1677_ (.B(_0833_),
    .C(_0862_),
    .A(_0819_),
    .Y(_0863_));
 sg13g2_nand3_1 _1678_ (.B(_0861_),
    .C(_0863_),
    .A(_0781_),
    .Y(_0864_));
 sg13g2_nand2_1 _1679_ (.Y(_0002_),
    .A(_0859_),
    .B(_0864_));
 sg13g2_or2_1 _1680_ (.X(_0865_),
    .B(_0819_),
    .A(net219));
 sg13g2_nand3_1 _1681_ (.B(_0806_),
    .C(_0838_),
    .A(net215),
    .Y(_0866_));
 sg13g2_nand3_1 _1682_ (.B(_0865_),
    .C(_0866_),
    .A(net213),
    .Y(_0867_));
 sg13g2_a21oi_1 _1683_ (.A1(_0808_),
    .A2(_0826_),
    .Y(_0868_),
    .B1(_0791_));
 sg13g2_o21ai_1 _1684_ (.B1(_0867_),
    .Y(_0869_),
    .A1(_0850_),
    .A2(_0868_));
 sg13g2_o21ai_1 _1685_ (.B1(_0859_),
    .Y(_0003_),
    .A1(net216),
    .A2(_0869_));
 sg13g2_or2_1 _1686_ (.X(_0870_),
    .B(_0860_),
    .A(_0781_));
 sg13g2_nand3_1 _1687_ (.B(net213),
    .C(_0862_),
    .A(_0823_),
    .Y(_0871_));
 sg13g2_nand3_1 _1688_ (.B(_0839_),
    .C(_0865_),
    .A(_0167_),
    .Y(_0872_));
 sg13g2_nand2_1 _1689_ (.Y(_0873_),
    .A(_0871_),
    .B(_0872_));
 sg13g2_o21ai_1 _1690_ (.B1(_0870_),
    .Y(_0004_),
    .A1(net216),
    .A2(_0873_));
 sg13g2_and2_1 _1691_ (.A(net214),
    .B(_0839_),
    .X(_0874_));
 sg13g2_o21ai_1 _1692_ (.B1(_0841_),
    .Y(_0875_),
    .A1(_0857_),
    .A2(_0874_));
 sg13g2_nand2_1 _1693_ (.Y(_0876_),
    .A(_0809_),
    .B(_0845_));
 sg13g2_nand2_1 _1694_ (.Y(_0877_),
    .A(_0840_),
    .B(_0876_));
 sg13g2_a21o_1 _1695_ (.A2(_0876_),
    .A1(_0840_),
    .B1(net214),
    .X(_0878_));
 sg13g2_a21oi_1 _1696_ (.A1(_0792_),
    .A2(_0862_),
    .Y(_0879_),
    .B1(net213));
 sg13g2_nor2_1 _1697_ (.A(net216),
    .B(net213),
    .Y(_0880_));
 sg13g2_nand3_1 _1698_ (.B(_0809_),
    .C(_0845_),
    .A(net215),
    .Y(_0881_));
 sg13g2_nand4_1 _1699_ (.B(_0810_),
    .C(_0838_),
    .A(net214),
    .Y(_0882_),
    .D(_0839_));
 sg13g2_nand3_1 _1700_ (.B(_0881_),
    .C(_0882_),
    .A(_0849_),
    .Y(_0883_));
 sg13g2_a221oi_1 _1701_ (.B2(net213),
    .C1(_0168_),
    .B1(_0883_),
    .A1(_0878_),
    .Y(_0884_),
    .A2(_0879_));
 sg13g2_a21oi_1 _1702_ (.A1(net216),
    .A2(_0875_),
    .Y(_0005_),
    .B1(_0884_));
 sg13g2_nand3_1 _1703_ (.B(_0826_),
    .C(_0839_),
    .A(net214),
    .Y(_0885_));
 sg13g2_nand3_1 _1704_ (.B(_0862_),
    .C(_0876_),
    .A(net215),
    .Y(_0886_));
 sg13g2_o21ai_1 _1705_ (.B1(_0880_),
    .Y(_0887_),
    .A1(_0835_),
    .A2(_0885_));
 sg13g2_nand2b_1 _1706_ (.Y(_0888_),
    .B(_0886_),
    .A_N(_0887_));
 sg13g2_nor2_2 _1707_ (.A(net216),
    .B(_0167_),
    .Y(_0889_));
 sg13g2_a21oi_1 _1708_ (.A1(_0837_),
    .A2(_0848_),
    .Y(_0890_),
    .B1(_0817_));
 sg13g2_nand2b_1 _1709_ (.Y(_0891_),
    .B(_0889_),
    .A_N(_0890_));
 sg13g2_nand3_1 _1710_ (.B(_0888_),
    .C(_0891_),
    .A(_0870_),
    .Y(_0006_));
 sg13g2_o21ai_1 _1711_ (.B1(_0823_),
    .Y(_0892_),
    .A1(net215),
    .A2(_0817_));
 sg13g2_nand2_1 _1712_ (.Y(_0893_),
    .A(_0880_),
    .B(_0892_));
 sg13g2_nand3b_1 _1713_ (.B(net215),
    .C(_0826_),
    .Y(_0894_),
    .A_N(_0845_));
 sg13g2_nand3_1 _1714_ (.B(_0889_),
    .C(_0894_),
    .A(_0885_),
    .Y(_0895_));
 sg13g2_nand3_1 _1715_ (.B(_0845_),
    .C(_0846_),
    .A(_0809_),
    .Y(_0896_));
 sg13g2_nand3_1 _1716_ (.B(_0895_),
    .C(_0896_),
    .A(_0893_),
    .Y(_0007_));
 sg13g2_a221oi_1 _1717_ (.B2(_0825_),
    .C1(net214),
    .B1(_0841_),
    .A1(_0806_),
    .Y(_0897_),
    .A2(_0837_));
 sg13g2_o21ai_1 _1718_ (.B1(_0880_),
    .Y(_0898_),
    .A1(net219),
    .A2(_0818_));
 sg13g2_nand4_1 _1719_ (.B(_0820_),
    .C(_0838_),
    .A(net215),
    .Y(_0899_),
    .D(_0839_));
 sg13g2_and2_1 _1720_ (.A(_0889_),
    .B(_0899_),
    .X(_0900_));
 sg13g2_a22oi_1 _1721_ (.Y(_0901_),
    .B1(_0900_),
    .B2(_0834_),
    .A2(_0877_),
    .A1(_0846_));
 sg13g2_o21ai_1 _1722_ (.B1(_0901_),
    .Y(_0008_),
    .A1(_0897_),
    .A2(_0898_));
 sg13g2_and2_1 _1723_ (.A(net213),
    .B(_0885_),
    .X(_0902_));
 sg13g2_o21ai_1 _1724_ (.B1(_0862_),
    .Y(_0903_),
    .A1(_0807_),
    .A2(_0826_));
 sg13g2_a21oi_1 _1725_ (.A1(net219),
    .A2(_0903_),
    .Y(_0904_),
    .B1(_0889_));
 sg13g2_o21ai_1 _1726_ (.B1(net216),
    .Y(_0905_),
    .A1(net219),
    .A2(_0821_));
 sg13g2_o21ai_1 _1727_ (.B1(_0905_),
    .Y(_0009_),
    .A1(_0902_),
    .A2(_0904_));
 sg13g2_nor2_1 _1728_ (.A(net198),
    .B(\counter.oled_driver.mc_exec.spi_tx_trigger_out ),
    .Y(_0906_));
 sg13g2_nor2_1 _1729_ (.A(_0740_),
    .B(net199),
    .Y(_0010_));
 sg13g2_a21oi_1 _1730_ (.A1(_0573_),
    .A2(_0578_),
    .Y(_0013_),
    .B1(_0740_));
 sg13g2_nand2_1 _1731_ (.Y(_0907_),
    .A(_0563_),
    .B(net270));
 sg13g2_a21oi_1 _1732_ (.A1(_0565_),
    .A2(_0574_),
    .Y(_0015_),
    .B1(_0907_));
 sg13g2_a21oi_1 _1733_ (.A1(_0575_),
    .A2(_0579_),
    .Y(_0014_),
    .B1(_0907_));
 sg13g2_o21ai_1 _1734_ (.B1(net270),
    .Y(_0908_),
    .A1(net357),
    .A2(net397));
 sg13g2_nor2_1 _1735_ (.A(net257),
    .B(_0908_),
    .Y(_0012_));
 sg13g2_or2_1 _1736_ (.X(\counter.oled_dc_out ),
    .B(net256),
    .A(\counter.oled_driver.mc_exec.oled_dc_out ));
 sg13g2_nor2_1 _1737_ (.A(net347),
    .B(net364),
    .Y(_0909_));
 sg13g2_nand2b_1 _1738_ (.Y(_0910_),
    .B(net277),
    .A_N(_0724_));
 sg13g2_nor2_1 _1739_ (.A(_0909_),
    .B(_0910_),
    .Y(_0011_));
 sg13g2_nor2_1 _1740_ (.A(clknet_1_0__leaf_clk),
    .B(_0910_),
    .Y(\counter.oled_clk_out ));
 sg13g2_and2_1 _1741_ (.A(_0565_),
    .B(net235),
    .X(_0911_));
 sg13g2_and3_1 _1742_ (.X(_0912_),
    .A(\counter.oled_driver.ready_out ),
    .B(\counter.streamer.state_r[5] ),
    .C(_0692_));
 sg13g2_nor2_1 _1743_ (.A(_0911_),
    .B(_0912_),
    .Y(_0913_));
 sg13g2_a21o_1 _1744_ (.A2(_0734_),
    .A1(\counter.streamer.state_r[5] ),
    .B1(_0913_),
    .X(_0914_));
 sg13g2_and2_1 _1745_ (.A(net274),
    .B(net224),
    .X(_0915_));
 sg13g2_nand2_1 _1746_ (.Y(_0916_),
    .A(net274),
    .B(net224));
 sg13g2_nor2_1 _1747_ (.A(_0561_),
    .B(_0916_),
    .Y(_0917_));
 sg13g2_nand2_1 _1748_ (.Y(_0918_),
    .A(\counter.streamer.state_r[5] ),
    .B(_0733_));
 sg13g2_nor3_1 _1749_ (.A(net261),
    .B(net224),
    .C(_0918_),
    .Y(_0919_));
 sg13g2_nand2_1 _1750_ (.Y(_0920_),
    .A(net248),
    .B(\counter.streamer.graphical_decoder.index_x_in[0] ));
 sg13g2_nand3_1 _1751_ (.B(net248),
    .C(\counter.streamer.graphical_decoder.index_x_in[0] ),
    .A(\counter.streamer.graphical_decoder.index_x_in[2] ),
    .Y(_0921_));
 sg13g2_nand4_1 _1752_ (.B(\counter.streamer.graphical_decoder.index_x_in[2] ),
    .C(net248),
    .A(\counter.streamer.graphical_decoder.index_x_in[3] ),
    .Y(_0922_),
    .D(\counter.streamer.graphical_decoder.index_x_in[0] ));
 sg13g2_xor2_1 _1753_ (.B(_0922_),
    .A(net461),
    .X(_0923_));
 sg13g2_a21o_1 _1754_ (.A2(_0923_),
    .A1(_0919_),
    .B1(_0917_),
    .X(_0124_));
 sg13g2_nor2_1 _1755_ (.A(net224),
    .B(_0921_),
    .Y(_0924_));
 sg13g2_nor2_1 _1756_ (.A(net455),
    .B(_0924_),
    .Y(_0925_));
 sg13g2_a21oi_1 _1757_ (.A1(net401),
    .A2(_0922_),
    .Y(_0926_),
    .B1(net224));
 sg13g2_nor3_2 _1758_ (.A(net261),
    .B(net456),
    .C(_0926_),
    .Y(_0123_));
 sg13g2_inv_1 _1759_ (.Y(_0927_),
    .A(_0123_));
 sg13g2_xnor2_1 _1760_ (.Y(_0928_),
    .A(_0580_),
    .B(_0920_));
 sg13g2_a22oi_1 _1761_ (.Y(_0929_),
    .B1(_0919_),
    .B2(_0928_),
    .A2(_0915_),
    .A1(net458));
 sg13g2_inv_1 _1762_ (.Y(_0122_),
    .A(_0929_));
 sg13g2_a21oi_1 _1763_ (.A1(_0927_),
    .A2(_0929_),
    .Y(_0107_),
    .B1(_0124_));
 sg13g2_o21ai_1 _1764_ (.B1(\counter.streamer.state_r[5] ),
    .Y(_0930_),
    .A1(net248),
    .A2(\counter.streamer.graphical_decoder.index_x_in[0] ));
 sg13g2_nand2b_1 _1765_ (.Y(_0931_),
    .B(_0920_),
    .A_N(_0930_));
 sg13g2_nand2_1 _1766_ (.Y(_0932_),
    .A(net248),
    .B(net224));
 sg13g2_o21ai_1 _1767_ (.B1(_0932_),
    .Y(_0933_),
    .A1(net224),
    .A2(_0931_));
 sg13g2_nand2_1 _1768_ (.Y(_0934_),
    .A(_0122_),
    .B(_0933_));
 sg13g2_xnor2_1 _1769_ (.Y(_0935_),
    .A(_0927_),
    .B(_0934_));
 sg13g2_nor2_1 _1770_ (.A(_0124_),
    .B(_0935_),
    .Y(_0239_));
 sg13g2_nor2_1 _1771_ (.A(_0734_),
    .B(_0918_),
    .Y(_0936_));
 sg13g2_nor2_1 _1772_ (.A(\counter.streamer.graphical_decoder.index_x_in[0] ),
    .B(_0913_),
    .Y(_0937_));
 sg13g2_a22oi_1 _1773_ (.Y(_0938_),
    .B1(_0936_),
    .B2(_0937_),
    .A2(net224),
    .A1(net463));
 sg13g2_nor2_1 _1774_ (.A(_0934_),
    .B(_0938_),
    .Y(_0939_));
 sg13g2_nor2_1 _1775_ (.A(net261),
    .B(_0938_),
    .Y(_0120_));
 sg13g2_nor2_1 _1776_ (.A(_0933_),
    .B(_0120_),
    .Y(_0940_));
 sg13g2_nor2_1 _1777_ (.A(_0929_),
    .B(_0940_),
    .Y(_0941_));
 sg13g2_inv_1 _1778_ (.Y(_0942_),
    .A(_0941_));
 sg13g2_nor2_1 _1779_ (.A(_0939_),
    .B(_0942_),
    .Y(_0943_));
 sg13g2_nor2b_1 _1780_ (.A(_0943_),
    .B_N(_0239_),
    .Y(_0108_));
 sg13g2_a21oi_1 _1781_ (.A1(_0034_),
    .A2(net229),
    .Y(_0944_),
    .B1(net255));
 sg13g2_nor2b_1 _1782_ (.A(net196),
    .B_N(net253),
    .Y(_0945_));
 sg13g2_nor3_1 _1783_ (.A(net225),
    .B(_0944_),
    .C(_0945_),
    .Y(_0946_));
 sg13g2_nor2_1 _1784_ (.A(\counter.oled_driver.spi_driver.shift_reg.start_in ),
    .B(net226),
    .Y(_0947_));
 sg13g2_a221oi_1 _1785_ (.B2(net440),
    .C1(_0946_),
    .B1(net223),
    .A1(net291),
    .Y(_0948_),
    .A2(net226));
 sg13g2_nor2_1 _1786_ (.A(net263),
    .B(_0948_),
    .Y(_0109_));
 sg13g2_a22oi_1 _1787_ (.Y(_0949_),
    .B1(net223),
    .B2(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[2] ),
    .A2(net226),
    .A1(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[1] ));
 sg13g2_a21oi_1 _1788_ (.A1(net253),
    .A2(net300),
    .Y(_0950_),
    .B1(net225));
 sg13g2_o21ai_1 _1789_ (.B1(_0950_),
    .Y(_0951_),
    .A1(net253),
    .A2(_0644_));
 sg13g2_a21oi_1 _1790_ (.A1(_0949_),
    .A2(net301),
    .Y(_0110_),
    .B1(net262));
 sg13g2_nor2_1 _1791_ (.A(net255),
    .B(_0643_),
    .Y(_0952_));
 sg13g2_nor2b_1 _1792_ (.A(net178),
    .B_N(net254),
    .Y(_0953_));
 sg13g2_nor3_1 _1793_ (.A(net225),
    .B(_0952_),
    .C(_0953_),
    .Y(_0954_));
 sg13g2_a221oi_1 _1794_ (.B2(net435),
    .C1(_0954_),
    .B1(net223),
    .A1(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[2] ),
    .Y(_0955_),
    .A2(net226));
 sg13g2_nor2_1 _1795_ (.A(net263),
    .B(net436),
    .Y(_0111_));
 sg13g2_a21oi_1 _1796_ (.A1(net253),
    .A2(net333),
    .Y(_0956_),
    .B1(net225));
 sg13g2_o21ai_1 _1797_ (.B1(_0956_),
    .Y(_0957_),
    .A1(net255),
    .A2(_0641_));
 sg13g2_a22oi_1 _1798_ (.Y(_0958_),
    .B1(net223),
    .B2(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[4] ),
    .A2(net226),
    .A1(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[3] ));
 sg13g2_a21oi_1 _1799_ (.A1(net334),
    .A2(_0958_),
    .Y(_0112_),
    .B1(net262));
 sg13g2_a22oi_1 _1800_ (.Y(_0959_),
    .B1(net223),
    .B2(net317),
    .A2(net226),
    .A1(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[4] ));
 sg13g2_a21oi_1 _1801_ (.A1(_0554_),
    .A2(net254),
    .Y(_0960_),
    .B1(net225));
 sg13g2_o21ai_1 _1802_ (.B1(_0960_),
    .Y(_0961_),
    .A1(net253),
    .A2(_0639_));
 sg13g2_a21oi_1 _1803_ (.A1(net318),
    .A2(_0961_),
    .Y(_0113_),
    .B1(net263));
 sg13g2_a21oi_1 _1804_ (.A1(_0039_),
    .A2(net229),
    .Y(_0962_),
    .B1(net255));
 sg13g2_nor2b_1 _1805_ (.A(net212),
    .B_N(net254),
    .Y(_0963_));
 sg13g2_nor3_1 _1806_ (.A(_0730_),
    .B(_0962_),
    .C(_0963_),
    .Y(_0964_));
 sg13g2_a221oi_1 _1807_ (.B2(net430),
    .C1(_0964_),
    .B1(net223),
    .A1(net317),
    .Y(_0965_),
    .A2(_0725_));
 sg13g2_nor2_1 _1808_ (.A(net265),
    .B(_0965_),
    .Y(_0114_));
 sg13g2_a22oi_1 _1809_ (.Y(_0966_),
    .B1(_0947_),
    .B2(net309),
    .A2(net226),
    .A1(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[6] ));
 sg13g2_nand2b_1 _1810_ (.Y(_0967_),
    .B(_0649_),
    .A_N(net255));
 sg13g2_a21oi_1 _1811_ (.A1(net253),
    .A2(_0048_),
    .Y(_0968_),
    .B1(net225));
 sg13g2_nand2_1 _1812_ (.Y(_0969_),
    .A(_0967_),
    .B(_0968_));
 sg13g2_a21oi_1 _1813_ (.A1(net310),
    .A2(_0969_),
    .Y(_0115_),
    .B1(net265));
 sg13g2_a21oi_1 _1814_ (.A1(\counter.oled_driver.ready_out ),
    .A2(\counter.oled_driver.sync_stb_in ),
    .Y(_0970_),
    .B1(net293));
 sg13g2_o21ai_1 _1815_ (.B1(net270),
    .Y(_0971_),
    .A1(\counter.oled_driver.ready_out ),
    .A2(_0576_));
 sg13g2_nor2_1 _1816_ (.A(net294),
    .B(_0971_),
    .Y(_0116_));
 sg13g2_nor2_2 _1817_ (.A(_0914_),
    .B(_0936_),
    .Y(_0972_));
 sg13g2_o21ai_1 _1818_ (.B1(_0972_),
    .Y(_0973_),
    .A1(net453),
    .A2(_0736_));
 sg13g2_nand2_1 _1819_ (.Y(_0974_),
    .A(net274),
    .B(_0973_));
 sg13g2_nor2b_1 _1820_ (.A(_0972_),
    .B_N(net251),
    .Y(_0975_));
 sg13g2_a21oi_1 _1821_ (.A1(net182),
    .A2(_0972_),
    .Y(_0976_),
    .B1(_0975_));
 sg13g2_nand2b_1 _1822_ (.Y(_0117_),
    .B(_0976_),
    .A_N(_0974_));
 sg13g2_and2_1 _1823_ (.A(net249),
    .B(net251),
    .X(_0977_));
 sg13g2_nor3_1 _1824_ (.A(net249),
    .B(net251),
    .C(net438),
    .Y(_0978_));
 sg13g2_o21ai_1 _1825_ (.B1(net401),
    .Y(_0979_),
    .A1(_0977_),
    .A2(_0978_));
 sg13g2_o21ai_1 _1826_ (.B1(net275),
    .Y(_0980_),
    .A1(net249),
    .A2(_0972_));
 sg13g2_a21oi_1 _1827_ (.A1(_0972_),
    .A2(_0979_),
    .Y(_0118_),
    .B1(_0980_));
 sg13g2_a21oi_1 _1828_ (.A1(_0735_),
    .A2(_0972_),
    .Y(_0981_),
    .B1(_0562_));
 sg13g2_or2_1 _1829_ (.X(_0119_),
    .B(_0981_),
    .A(_0974_));
 sg13g2_and2_1 _1830_ (.A(net274),
    .B(_0933_),
    .X(_0121_));
 sg13g2_o21ai_1 _1831_ (.B1(net459),
    .Y(_0982_),
    .A1(_0911_),
    .A2(_0912_));
 sg13g2_o21ai_1 _1832_ (.B1(_0982_),
    .Y(_0983_),
    .A1(net459),
    .A2(_0912_));
 sg13g2_nor2_1 _1833_ (.A(net261),
    .B(net460),
    .Y(_0125_));
 sg13g2_a21oi_1 _1834_ (.A1(_0559_),
    .A2(_0982_),
    .Y(_0126_),
    .B1(_0916_));
 sg13g2_o21ai_1 _1835_ (.B1(net275),
    .Y(_0984_),
    .A1(net366),
    .A2(net232));
 sg13g2_a21oi_1 _1836_ (.A1(_0552_),
    .A2(net232),
    .Y(_0127_),
    .B1(_0984_));
 sg13g2_o21ai_1 _1837_ (.B1(net272),
    .Y(_0985_),
    .A1(net415),
    .A2(net232));
 sg13g2_a21oi_1 _1838_ (.A1(_0551_),
    .A2(net232),
    .Y(_0128_),
    .B1(_0985_));
 sg13g2_o21ai_1 _1839_ (.B1(net272),
    .Y(_0986_),
    .A1(net421),
    .A2(net232));
 sg13g2_a21oi_1 _1840_ (.A1(_0550_),
    .A2(net232),
    .Y(_0129_),
    .B1(_0986_));
 sg13g2_o21ai_1 _1841_ (.B1(net272),
    .Y(_0987_),
    .A1(net327),
    .A2(net232));
 sg13g2_a21oi_1 _1842_ (.A1(_0549_),
    .A2(net232),
    .Y(_0130_),
    .B1(_0987_));
 sg13g2_o21ai_1 _1843_ (.B1(net272),
    .Y(_0988_),
    .A1(net418),
    .A2(net231));
 sg13g2_a21oi_1 _1844_ (.A1(_0548_),
    .A2(net231),
    .Y(_0131_),
    .B1(_0988_));
 sg13g2_o21ai_1 _1845_ (.B1(net272),
    .Y(_0989_),
    .A1(net407),
    .A2(net231));
 sg13g2_a21oi_1 _1846_ (.A1(_0547_),
    .A2(net231),
    .Y(_0132_),
    .B1(_0989_));
 sg13g2_o21ai_1 _1847_ (.B1(net272),
    .Y(_0990_),
    .A1(net447),
    .A2(net231));
 sg13g2_a21oi_1 _1848_ (.A1(_0546_),
    .A2(net231),
    .Y(_0133_),
    .B1(_0990_));
 sg13g2_o21ai_1 _1849_ (.B1(net272),
    .Y(_0991_),
    .A1(net342),
    .A2(net231));
 sg13g2_a21oi_1 _1850_ (.A1(_0545_),
    .A2(net231),
    .Y(_0134_),
    .B1(_0991_));
 sg13g2_o21ai_1 _1851_ (.B1(net272),
    .Y(_0992_),
    .A1(net419),
    .A2(net233));
 sg13g2_a21oi_1 _1852_ (.A1(_0544_),
    .A2(net233),
    .Y(_0135_),
    .B1(_0992_));
 sg13g2_o21ai_1 _1853_ (.B1(net275),
    .Y(_0993_),
    .A1(net349),
    .A2(net233));
 sg13g2_a21oi_1 _1854_ (.A1(_0543_),
    .A2(net234),
    .Y(_0136_),
    .B1(_0993_));
 sg13g2_o21ai_1 _1855_ (.B1(net274),
    .Y(_0994_),
    .A1(net426),
    .A2(net233));
 sg13g2_a21oi_1 _1856_ (.A1(_0542_),
    .A2(net234),
    .Y(_0137_),
    .B1(_0994_));
 sg13g2_o21ai_1 _1857_ (.B1(net274),
    .Y(_0995_),
    .A1(net363),
    .A2(net234));
 sg13g2_a21oi_1 _1858_ (.A1(_0541_),
    .A2(net233),
    .Y(_0138_),
    .B1(_0995_));
 sg13g2_o21ai_1 _1859_ (.B1(net275),
    .Y(_0996_),
    .A1(net362),
    .A2(net234));
 sg13g2_a21oi_1 _1860_ (.A1(_0540_),
    .A2(net233),
    .Y(_0139_),
    .B1(_0996_));
 sg13g2_o21ai_1 _1861_ (.B1(net274),
    .Y(_0997_),
    .A1(net410),
    .A2(net238));
 sg13g2_a21oi_1 _1862_ (.A1(_0539_),
    .A2(net238),
    .Y(_0140_),
    .B1(_0997_));
 sg13g2_o21ai_1 _1863_ (.B1(net274),
    .Y(_0998_),
    .A1(net405),
    .A2(net238));
 sg13g2_a21oi_1 _1864_ (.A1(_0538_),
    .A2(net238),
    .Y(_0141_),
    .B1(_0998_));
 sg13g2_o21ai_1 _1865_ (.B1(net279),
    .Y(_0999_),
    .A1(net322),
    .A2(net238));
 sg13g2_a21oi_1 _1866_ (.A1(_0537_),
    .A2(net238),
    .Y(_0142_),
    .B1(_0999_));
 sg13g2_o21ai_1 _1867_ (.B1(net279),
    .Y(_1000_),
    .A1(net352),
    .A2(net237));
 sg13g2_a21oi_1 _1868_ (.A1(_0536_),
    .A2(net237),
    .Y(_0143_),
    .B1(_1000_));
 sg13g2_o21ai_1 _1869_ (.B1(net279),
    .Y(_1001_),
    .A1(net374),
    .A2(net237));
 sg13g2_a21oi_1 _1870_ (.A1(_0535_),
    .A2(net237),
    .Y(_0144_),
    .B1(_1001_));
 sg13g2_o21ai_1 _1871_ (.B1(net279),
    .Y(_1002_),
    .A1(net356),
    .A2(net237));
 sg13g2_a21oi_1 _1872_ (.A1(_0534_),
    .A2(net237),
    .Y(_0145_),
    .B1(_1002_));
 sg13g2_o21ai_1 _1873_ (.B1(net280),
    .Y(_1003_),
    .A1(net305),
    .A2(net237));
 sg13g2_a21oi_1 _1874_ (.A1(_0533_),
    .A2(net237),
    .Y(_0146_),
    .B1(_1003_));
 sg13g2_o21ai_1 _1875_ (.B1(net279),
    .Y(_1004_),
    .A1(net387),
    .A2(net236));
 sg13g2_a21oi_1 _1876_ (.A1(_0558_),
    .A2(net236),
    .Y(_0147_),
    .B1(_1004_));
 sg13g2_o21ai_1 _1877_ (.B1(net279),
    .Y(_1005_),
    .A1(net420),
    .A2(net236));
 sg13g2_a21oi_1 _1878_ (.A1(_0557_),
    .A2(net236),
    .Y(_0148_),
    .B1(_1005_));
 sg13g2_o21ai_1 _1879_ (.B1(net279),
    .Y(_1006_),
    .A1(net412),
    .A2(net236));
 sg13g2_a21oi_1 _1880_ (.A1(_0556_),
    .A2(net236),
    .Y(_0149_),
    .B1(_1006_));
 sg13g2_o21ai_1 _1881_ (.B1(net279),
    .Y(_1007_),
    .A1(net406),
    .A2(net236));
 sg13g2_a21oi_1 _1882_ (.A1(_0555_),
    .A2(net236),
    .Y(_0150_),
    .B1(_1007_));
 sg13g2_nor2_1 _1883_ (.A(\counter.oled_driver.ready_out ),
    .B(\counter.oled_driver.state_r[0] ),
    .Y(_1008_));
 sg13g2_o21ai_1 _1884_ (.B1(_0659_),
    .Y(_1009_),
    .A1(\counter.oled_driver.state_r[4] ),
    .A2(_1008_));
 sg13g2_o21ai_1 _1885_ (.B1(\counter.oled_driver.ready_out ),
    .Y(_1010_),
    .A1(_0574_),
    .A2(\counter.oled_driver.sync_stb_in ));
 sg13g2_nand2_2 _1886_ (.Y(_1011_),
    .A(_1009_),
    .B(_1010_));
 sg13g2_nor2_2 _1887_ (.A(_0563_),
    .B(net222),
    .Y(_1012_));
 sg13g2_nor2_1 _1888_ (.A(\counter.streamer.digits_r[17] ),
    .B(\counter.streamer.digit_cnt_r[0] ),
    .Y(_1013_));
 sg13g2_nand2b_2 _1889_ (.Y(_0240_),
    .B(\counter.streamer.digit_cnt_r[2] ),
    .A_N(net250));
 sg13g2_nor2b_1 _1890_ (.A(\counter.streamer.digits_r[21] ),
    .B_N(\counter.streamer.digit_cnt_r[0] ),
    .Y(_0241_));
 sg13g2_nor3_2 _1891_ (.A(_1013_),
    .B(_0240_),
    .C(_0241_),
    .Y(_0242_));
 sg13g2_mux4_1 _1892_ (.S0(net251),
    .A0(\counter.streamer.digits_r[1] ),
    .A1(\counter.streamer.digits_r[5] ),
    .A2(\counter.streamer.digits_r[9] ),
    .A3(\counter.streamer.digits_r[13] ),
    .S1(net250),
    .X(_0243_));
 sg13g2_and2_2 _1893_ (.A(_0562_),
    .B(_0243_),
    .X(_0244_));
 sg13g2_nor2_1 _1894_ (.A(_0242_),
    .B(_0244_),
    .Y(_0245_));
 sg13g2_or2_1 _1895_ (.X(_0246_),
    .B(_0244_),
    .A(_0242_));
 sg13g2_mux4_1 _1896_ (.S0(net251),
    .A0(\counter.streamer.digits_r[0] ),
    .A1(\counter.streamer.digits_r[4] ),
    .A2(\counter.streamer.digits_r[8] ),
    .A3(\counter.streamer.digits_r[12] ),
    .S1(net250),
    .X(_0247_));
 sg13g2_and2_1 _1897_ (.A(_0562_),
    .B(_0247_),
    .X(_0248_));
 sg13g2_nor2_1 _1898_ (.A(\counter.streamer.digits_r[16] ),
    .B(net252),
    .Y(_0249_));
 sg13g2_nor2b_1 _1899_ (.A(\counter.streamer.digits_r[20] ),
    .B_N(net252),
    .Y(_0250_));
 sg13g2_nor3_2 _1900_ (.A(_0240_),
    .B(_0249_),
    .C(_0250_),
    .Y(_0251_));
 sg13g2_nor2_1 _1901_ (.A(_0248_),
    .B(_0251_),
    .Y(_0252_));
 sg13g2_or2_2 _1902_ (.X(_0253_),
    .B(_0251_),
    .A(_0248_));
 sg13g2_nor4_2 _1903_ (.A(_0242_),
    .B(_0244_),
    .C(_0248_),
    .Y(_0254_),
    .D(_0251_));
 sg13g2_mux4_1 _1904_ (.S0(net252),
    .A0(\counter.streamer.digits_r[2] ),
    .A1(\counter.streamer.digits_r[6] ),
    .A2(\counter.streamer.digits_r[10] ),
    .A3(\counter.streamer.digits_r[14] ),
    .S1(net249),
    .X(_0255_));
 sg13g2_and2_1 _1905_ (.A(_0562_),
    .B(_0255_),
    .X(_0256_));
 sg13g2_nor2_1 _1906_ (.A(\counter.streamer.digits_r[18] ),
    .B(net252),
    .Y(_0257_));
 sg13g2_nor2b_1 _1907_ (.A(\counter.streamer.digits_r[22] ),
    .B_N(net252),
    .Y(_0258_));
 sg13g2_nor3_2 _1908_ (.A(_0240_),
    .B(_0257_),
    .C(_0258_),
    .Y(_0259_));
 sg13g2_nor2_2 _1909_ (.A(_0256_),
    .B(_0259_),
    .Y(_0260_));
 sg13g2_or2_1 _1910_ (.X(_0261_),
    .B(_0259_),
    .A(_0256_));
 sg13g2_nand2_1 _1911_ (.Y(_0262_),
    .A(_0246_),
    .B(_0253_));
 sg13g2_o21ai_1 _1912_ (.B1(_0261_),
    .Y(_0263_),
    .A1(_0245_),
    .A2(_0252_));
 sg13g2_nor2b_1 _1913_ (.A(_0074_),
    .B_N(net250),
    .Y(_0264_));
 sg13g2_nor2_1 _1914_ (.A(net249),
    .B(_0072_),
    .Y(_0265_));
 sg13g2_nor3_1 _1915_ (.A(net251),
    .B(_0264_),
    .C(_0265_),
    .Y(_0266_));
 sg13g2_nor2b_1 _1916_ (.A(_0075_),
    .B_N(net250),
    .Y(_0267_));
 sg13g2_o21ai_1 _1917_ (.B1(net252),
    .Y(_0268_),
    .A1(net249),
    .A2(_0073_));
 sg13g2_o21ai_1 _1918_ (.B1(_0562_),
    .Y(_0269_),
    .A1(_0267_),
    .A2(_0268_));
 sg13g2_mux2_1 _1919_ (.A0(\counter.streamer.digits_r[19] ),
    .A1(\counter.streamer.digits_r[23] ),
    .S(net252),
    .X(_0270_));
 sg13g2_nand3_1 _1920_ (.B(_0071_),
    .C(_0270_),
    .A(\counter.streamer.digit_cnt_r[2] ),
    .Y(_0271_));
 sg13g2_o21ai_1 _1921_ (.B1(_0271_),
    .Y(_0272_),
    .A1(_0266_),
    .A2(_0269_));
 sg13g2_inv_1 _1922_ (.Y(_0273_),
    .A(_0272_));
 sg13g2_nor2_1 _1923_ (.A(_0254_),
    .B(_0272_),
    .Y(_0274_));
 sg13g2_nor2_1 _1924_ (.A(_0246_),
    .B(_0260_),
    .Y(_0275_));
 sg13g2_and2_1 _1925_ (.A(_0253_),
    .B(_0272_),
    .X(_0276_));
 sg13g2_o21ai_1 _1926_ (.B1(\counter.streamer.graphical_decoder.index_x_in[3] ),
    .Y(_0277_),
    .A1(\counter.streamer.graphical_decoder.index_x_in[2] ),
    .A2(net248));
 sg13g2_nand2_1 _1927_ (.Y(_0278_),
    .A(_0065_),
    .B(_0277_));
 sg13g2_nand3_1 _1928_ (.B(_0065_),
    .C(_0277_),
    .A(_0559_),
    .Y(_0279_));
 sg13g2_a221oi_1 _1929_ (.B2(_0276_),
    .C1(_0279_),
    .B1(_0275_),
    .A1(_0263_),
    .Y(_0280_),
    .A2(_0274_));
 sg13g2_a21oi_1 _1930_ (.A1(_0245_),
    .A2(_0261_),
    .Y(_0281_),
    .B1(_0253_));
 sg13g2_or2_1 _1931_ (.X(_0282_),
    .B(_0278_),
    .A(_0076_));
 sg13g2_nor4_1 _1932_ (.A(_0242_),
    .B(_0244_),
    .C(_0256_),
    .D(_0259_),
    .Y(_0283_));
 sg13g2_a21oi_1 _1933_ (.A1(_0253_),
    .A2(_0283_),
    .Y(_0284_),
    .B1(_0282_));
 sg13g2_o21ai_1 _1934_ (.B1(_0284_),
    .Y(_0285_),
    .A1(_0272_),
    .A2(_0281_));
 sg13g2_nand2b_2 _1935_ (.Y(_0286_),
    .B(_0285_),
    .A_N(_0280_));
 sg13g2_inv_1 _1936_ (.Y(_0287_),
    .A(_0286_));
 sg13g2_and3_1 _1937_ (.X(_0288_),
    .A(_0245_),
    .B(_0253_),
    .C(_0272_));
 sg13g2_a21oi_1 _1938_ (.A1(_0260_),
    .A2(_0262_),
    .Y(_0289_),
    .B1(_0288_));
 sg13g2_o21ai_1 _1939_ (.B1(_0273_),
    .Y(_0290_),
    .A1(_0254_),
    .A2(_0263_));
 sg13g2_nand2_1 _1940_ (.Y(_0291_),
    .A(_0076_),
    .B(_0278_));
 sg13g2_a21o_1 _1941_ (.A2(_0290_),
    .A1(_0289_),
    .B1(_0291_),
    .X(_0292_));
 sg13g2_a21oi_1 _1942_ (.A1(_0260_),
    .A2(_0272_),
    .Y(_0293_),
    .B1(_0288_));
 sg13g2_nand3_1 _1943_ (.B(_0252_),
    .C(_0260_),
    .A(_0246_),
    .Y(_0294_));
 sg13g2_nand2_1 _1944_ (.Y(_0295_),
    .A(_0273_),
    .B(_0294_));
 sg13g2_nand2b_1 _1945_ (.Y(_0296_),
    .B(_0278_),
    .A_N(_0076_));
 sg13g2_a21o_1 _1946_ (.A2(_0295_),
    .A1(_0293_),
    .B1(_0296_),
    .X(_0297_));
 sg13g2_and2_1 _1947_ (.A(_0292_),
    .B(_0297_),
    .X(_0298_));
 sg13g2_nor2b_1 _1948_ (.A(_0280_),
    .B_N(_0292_),
    .Y(_0299_));
 sg13g2_nand3b_1 _1949_ (.B(_0292_),
    .C(_0297_),
    .Y(_0300_),
    .A_N(_0286_));
 sg13g2_a21oi_1 _1950_ (.A1(_0285_),
    .A2(_0297_),
    .Y(_0301_),
    .B1(_0581_));
 sg13g2_mux2_1 _1951_ (.A0(\counter.streamer.graphical_decoder.index_y_in[0] ),
    .A1(_0301_),
    .S(_0299_),
    .X(_0302_));
 sg13g2_nand2_1 _1952_ (.Y(_0303_),
    .A(\counter.streamer.graphical_decoder.index_x_in[1] ),
    .B(_0286_));
 sg13g2_a21oi_1 _1953_ (.A1(_0292_),
    .A2(_0297_),
    .Y(_0304_),
    .B1(_0582_));
 sg13g2_a21o_1 _1954_ (.A2(_0297_),
    .A1(_0292_),
    .B1(_0582_),
    .X(_0305_));
 sg13g2_a22oi_1 _1955_ (.Y(_0306_),
    .B1(_0303_),
    .B2(_0305_),
    .A2(_0300_),
    .A1(_0580_));
 sg13g2_and4_1 _1956_ (.A(_0580_),
    .B(_0300_),
    .C(_0303_),
    .D(_0305_),
    .X(_0307_));
 sg13g2_a221oi_1 _1957_ (.B2(_0305_),
    .C1(_0066_),
    .B1(_0303_),
    .A1(_0287_),
    .Y(_0308_),
    .A2(_0298_));
 sg13g2_a221oi_1 _1958_ (.B2(_0580_),
    .C1(_0304_),
    .B1(_0300_),
    .A1(net248),
    .Y(_0309_),
    .A2(_0286_));
 sg13g2_nor2_1 _1959_ (.A(_0308_),
    .B(_0309_),
    .Y(_0310_));
 sg13g2_o21ai_1 _1960_ (.B1(_0302_),
    .Y(_0311_),
    .A1(_0306_),
    .A2(_0307_));
 sg13g2_nand2b_1 _1961_ (.Y(_0312_),
    .B(_0559_),
    .A_N(_0311_));
 sg13g2_nor3_2 _1962_ (.A(_0302_),
    .B(_0308_),
    .C(_0309_),
    .Y(_0313_));
 sg13g2_nand2_1 _1963_ (.Y(_0314_),
    .A(_0246_),
    .B(_0260_));
 sg13g2_nand3_1 _1964_ (.B(_0273_),
    .C(_0314_),
    .A(_0263_),
    .Y(_0315_));
 sg13g2_nor2_1 _1965_ (.A(\counter.streamer.graphical_decoder.index_x_in[3] ),
    .B(\counter.streamer.graphical_decoder.index_x_in[2] ),
    .Y(_0316_));
 sg13g2_nor3_2 _1966_ (.A(_0561_),
    .B(_0732_),
    .C(_0316_),
    .Y(_0317_));
 sg13g2_nor2_1 _1967_ (.A(_0253_),
    .B(_0273_),
    .Y(_0318_));
 sg13g2_a21oi_1 _1968_ (.A1(_0275_),
    .A2(_0318_),
    .Y(_0319_),
    .B1(_0317_));
 sg13g2_nand4_1 _1969_ (.B(_0560_),
    .C(_0315_),
    .A(net247),
    .Y(_0320_),
    .D(_0319_));
 sg13g2_nor2_1 _1970_ (.A(_0070_),
    .B(_0320_),
    .Y(_0321_));
 sg13g2_a21oi_1 _1971_ (.A1(net246),
    .A2(_0313_),
    .Y(_0322_),
    .B1(_0321_));
 sg13g2_nand2_1 _1972_ (.Y(_0323_),
    .A(_0312_),
    .B(_0322_));
 sg13g2_a22oi_1 _1973_ (.Y(_0324_),
    .B1(_1012_),
    .B2(_0323_),
    .A2(_1011_),
    .A1(net298));
 sg13g2_nor2_1 _1974_ (.A(net263),
    .B(net299),
    .Y(_0151_));
 sg13g2_nand2_1 _1975_ (.Y(_0325_),
    .A(\counter.streamer.graphical_decoder.index_x_in[0] ),
    .B(_0286_));
 sg13g2_o21ai_1 _1976_ (.B1(_0325_),
    .Y(_0326_),
    .A1(_0584_),
    .A2(_0298_));
 sg13g2_and2_1 _1977_ (.A(_0306_),
    .B(_0326_),
    .X(_0327_));
 sg13g2_nand2_1 _1978_ (.Y(_0328_),
    .A(_0306_),
    .B(_0326_));
 sg13g2_o21ai_1 _1979_ (.B1(net246),
    .Y(_0329_),
    .A1(_0313_),
    .A2(_0327_));
 sg13g2_nor2_1 _1980_ (.A(_0044_),
    .B(_0320_),
    .Y(_0330_));
 sg13g2_nor2_1 _1981_ (.A(_0252_),
    .B(_0283_),
    .Y(_0331_));
 sg13g2_nor3_2 _1982_ (.A(_0272_),
    .B(_0281_),
    .C(_0331_),
    .Y(_0332_));
 sg13g2_or2_1 _1983_ (.X(_0333_),
    .B(_0317_),
    .A(\counter.streamer.graphical_decoder.index_y_in[0] ));
 sg13g2_a21oi_1 _1984_ (.A1(_0260_),
    .A2(_0262_),
    .Y(_0334_),
    .B1(_0293_));
 sg13g2_nor4_2 _1985_ (.A(net247),
    .B(_0332_),
    .C(_0333_),
    .Y(_0335_),
    .D(_0334_));
 sg13g2_inv_1 _1986_ (.Y(_0336_),
    .A(_0335_));
 sg13g2_a21oi_1 _1987_ (.A1(\counter.streamer.graphical_decoder.pattern_adg[1] ),
    .A2(_0335_),
    .Y(_0337_),
    .B1(_0330_));
 sg13g2_nand3_1 _1988_ (.B(_0329_),
    .C(_0337_),
    .A(_0312_),
    .Y(_0338_));
 sg13g2_a22oi_1 _1989_ (.Y(_0339_),
    .B1(_1012_),
    .B2(_0338_),
    .A2(net222),
    .A1(net196));
 sg13g2_nor2_1 _1990_ (.A(net263),
    .B(net197),
    .Y(_0152_));
 sg13g2_nand2_1 _1991_ (.Y(_0340_),
    .A(net172),
    .B(net222));
 sg13g2_nand3_1 _1992_ (.B(_0300_),
    .C(_0326_),
    .A(_0580_),
    .Y(_0341_));
 sg13g2_nand2_1 _1993_ (.Y(_0342_),
    .A(_0310_),
    .B(_0341_));
 sg13g2_a21oi_1 _1994_ (.A1(_0310_),
    .A2(_0341_),
    .Y(_0343_),
    .B1(_0313_));
 sg13g2_nor2_1 _1995_ (.A(_0559_),
    .B(_0343_),
    .Y(_0344_));
 sg13g2_o21ai_1 _1996_ (.B1(_0312_),
    .Y(_0345_),
    .A1(_0070_),
    .A2(_0336_));
 sg13g2_o21ai_1 _1997_ (.B1(_1012_),
    .Y(_0346_),
    .A1(_0344_),
    .A2(_0345_));
 sg13g2_a21oi_1 _1998_ (.A1(_0340_),
    .A2(_0346_),
    .Y(_0153_),
    .B1(net262));
 sg13g2_nand2_1 _1999_ (.Y(_0347_),
    .A(net178),
    .B(net222));
 sg13g2_a21oi_1 _2000_ (.A1(_0311_),
    .A2(_0342_),
    .Y(_0348_),
    .B1(_0559_));
 sg13g2_a21oi_1 _2001_ (.A1(_0311_),
    .A2(_0328_),
    .Y(_0349_),
    .B1(net246));
 sg13g2_nor2_1 _2002_ (.A(_0734_),
    .B(_0317_),
    .Y(_0350_));
 sg13g2_o21ai_1 _2003_ (.B1(_0350_),
    .Y(_0351_),
    .A1(_0260_),
    .A2(_0262_));
 sg13g2_nor2_1 _2004_ (.A(_0273_),
    .B(_0294_),
    .Y(_0352_));
 sg13g2_nor3_2 _2005_ (.A(_0332_),
    .B(_0351_),
    .C(_0352_),
    .Y(_0353_));
 sg13g2_a22oi_1 _2006_ (.Y(_0354_),
    .B1(_0353_),
    .B2(\counter.streamer.graphical_decoder.pattern_adg[4] ),
    .A2(_0335_),
    .A1(_0583_));
 sg13g2_nand2b_1 _2007_ (.Y(_0355_),
    .B(_0354_),
    .A_N(_0349_));
 sg13g2_o21ai_1 _2008_ (.B1(_1012_),
    .Y(_0356_),
    .A1(_0348_),
    .A2(_0355_));
 sg13g2_a21oi_1 _2009_ (.A1(_0347_),
    .A2(_0356_),
    .Y(_0154_),
    .B1(net262));
 sg13g2_nand2_1 _2010_ (.Y(_0357_),
    .A(net169),
    .B(net222));
 sg13g2_a21oi_1 _2011_ (.A1(_0311_),
    .A2(_0342_),
    .Y(_0358_),
    .B1(net246));
 sg13g2_a21oi_1 _2012_ (.A1(_0311_),
    .A2(_0328_),
    .Y(_0359_),
    .B1(_0559_));
 sg13g2_a22oi_1 _2013_ (.Y(_0360_),
    .B1(_0353_),
    .B2(\counter.streamer.graphical_decoder.pattern_adg[3] ),
    .A2(_0335_),
    .A1(\counter.streamer.graphical_decoder.pattern_adg[4] ));
 sg13g2_nand2b_1 _2014_ (.Y(_0361_),
    .B(_0360_),
    .A_N(_0359_));
 sg13g2_o21ai_1 _2015_ (.B1(_1012_),
    .Y(_0362_),
    .A1(_0358_),
    .A2(_0361_));
 sg13g2_a21oi_1 _2016_ (.A1(_0357_),
    .A2(_0362_),
    .Y(_0155_),
    .B1(net262));
 sg13g2_nand2_1 _2017_ (.Y(_0363_),
    .A(net286),
    .B(net222));
 sg13g2_and2_1 _2018_ (.A(_0920_),
    .B(_0316_),
    .X(_0364_));
 sg13g2_nor3_1 _2019_ (.A(\counter.streamer.digit_cnt_r[2] ),
    .B(_0065_),
    .C(_0734_),
    .Y(_0365_));
 sg13g2_nand2_1 _2020_ (.Y(_0366_),
    .A(_0977_),
    .B(_0365_));
 sg13g2_nor3_1 _2021_ (.A(_0317_),
    .B(_0364_),
    .C(_0366_),
    .Y(_0367_));
 sg13g2_inv_1 _2022_ (.Y(_0368_),
    .A(_0367_));
 sg13g2_o21ai_1 _2023_ (.B1(_0368_),
    .Y(_0369_),
    .A1(_0559_),
    .A2(_0311_));
 sg13g2_nand2b_1 _2024_ (.Y(_0370_),
    .B(_0353_),
    .A_N(_0070_));
 sg13g2_o21ai_1 _2025_ (.B1(_0370_),
    .Y(_0371_),
    .A1(net246),
    .A2(_0343_));
 sg13g2_o21ai_1 _2026_ (.B1(_1012_),
    .Y(_0372_),
    .A1(_0369_),
    .A2(_0371_));
 sg13g2_a21oi_1 _2027_ (.A1(_0363_),
    .A2(_0372_),
    .Y(_0156_),
    .B1(net262));
 sg13g2_o21ai_1 _2028_ (.B1(_0559_),
    .Y(_0373_),
    .A1(_0313_),
    .A2(_0327_));
 sg13g2_and3_1 _2029_ (.X(_0374_),
    .A(\counter.streamer.graphical_decoder.index_y_in[0] ),
    .B(_0315_),
    .C(_0319_));
 sg13g2_nor2b_1 _2030_ (.A(net246),
    .B_N(\counter.streamer.graphical_decoder.pattern_adg[3] ),
    .Y(_0375_));
 sg13g2_a22oi_1 _2031_ (.Y(_0376_),
    .B1(_0374_),
    .B2(_0375_),
    .A2(_0353_),
    .A1(\counter.streamer.graphical_decoder.pattern_adg[1] ));
 sg13g2_nand3b_1 _2032_ (.B(_0373_),
    .C(_0376_),
    .Y(_0377_),
    .A_N(_0369_));
 sg13g2_a22oi_1 _2033_ (.Y(_0378_),
    .B1(_1012_),
    .B2(_0377_),
    .A2(net222),
    .A1(net212));
 sg13g2_nor2_1 _2034_ (.A(net262),
    .B(net281),
    .Y(_0157_));
 sg13g2_nand2_1 _2035_ (.Y(_0379_),
    .A(net170),
    .B(net222));
 sg13g2_a21oi_1 _2036_ (.A1(\counter.streamer.graphical_decoder.pattern_adg[2] ),
    .A2(_0374_),
    .Y(_0380_),
    .B1(_0313_));
 sg13g2_nor2_1 _2037_ (.A(net246),
    .B(_0380_),
    .Y(_0381_));
 sg13g2_o21ai_1 _2038_ (.B1(_1012_),
    .Y(_0382_),
    .A1(_0369_),
    .A2(_0381_));
 sg13g2_a21oi_1 _2039_ (.A1(_0379_),
    .A2(_0382_),
    .Y(_0158_),
    .B1(net262));
 sg13g2_nand2_2 _2040_ (.Y(_0383_),
    .A(net258),
    .B(_0666_));
 sg13g2_nor4_2 _2041_ (.A(_0035_),
    .B(_0569_),
    .C(_0635_),
    .Y(_0384_),
    .D(_0383_));
 sg13g2_nand2b_1 _2042_ (.Y(_0385_),
    .B(net336),
    .A_N(_0384_));
 sg13g2_nand2b_1 _2043_ (.Y(_0386_),
    .B(_0384_),
    .A_N(_0638_));
 sg13g2_nand3_1 _2044_ (.B(net337),
    .C(_0386_),
    .A(net277),
    .Y(_0159_));
 sg13g2_nor3_1 _2045_ (.A(_0568_),
    .B(_0635_),
    .C(_0383_),
    .Y(_0387_));
 sg13g2_inv_1 _2046_ (.Y(_0388_),
    .A(_0387_));
 sg13g2_nand4_1 _2047_ (.B(_0569_),
    .C(net230),
    .A(_0033_),
    .Y(_0389_),
    .D(_0387_));
 sg13g2_o21ai_1 _2048_ (.B1(net394),
    .Y(_0390_),
    .A1(_0036_),
    .A2(_0388_));
 sg13g2_nand3_1 _2049_ (.B(_0389_),
    .C(net395),
    .A(net277),
    .Y(_0160_));
 sg13g2_nor2b_1 _2050_ (.A(_0039_),
    .B_N(_0761_),
    .Y(_0391_));
 sg13g2_inv_1 _2051_ (.Y(_0392_),
    .A(_0391_));
 sg13g2_o21ai_1 _2052_ (.B1(_0751_),
    .Y(_0393_),
    .A1(_0571_),
    .A2(_0634_));
 sg13g2_a21oi_1 _2053_ (.A1(_0646_),
    .A2(_0666_),
    .Y(_0394_),
    .B1(_0392_));
 sg13g2_nor4_1 _2054_ (.A(_0748_),
    .B(_0762_),
    .C(_0393_),
    .D(_0394_),
    .Y(_0395_));
 sg13g2_or2_1 _2055_ (.X(_0396_),
    .B(_0638_),
    .A(_0056_));
 sg13g2_o21ai_1 _2056_ (.B1(net278),
    .Y(_0397_),
    .A1(net403),
    .A2(_0395_));
 sg13g2_a21oi_1 _2057_ (.A1(_0395_),
    .A2(_0396_),
    .Y(_0161_),
    .B1(_0397_));
 sg13g2_nor2_1 _2058_ (.A(_0569_),
    .B(_0388_),
    .Y(_0398_));
 sg13g2_o21ai_1 _2059_ (.B1(net277),
    .Y(_0399_),
    .A1(net384),
    .A2(_0398_));
 sg13g2_a21oi_1 _2060_ (.A1(_0638_),
    .A2(_0398_),
    .Y(_0162_),
    .B1(net385));
 sg13g2_o21ai_1 _2061_ (.B1(net434),
    .Y(_0400_),
    .A1(net221),
    .A2(net220));
 sg13g2_a21oi_1 _2062_ (.A1(_0797_),
    .A2(_0400_),
    .Y(_0163_),
    .B1(net264));
 sg13g2_o21ai_1 _2063_ (.B1(net413),
    .Y(_0401_),
    .A1(net221),
    .A2(net220));
 sg13g2_a21oi_1 _2064_ (.A1(_0804_),
    .A2(_0401_),
    .Y(_0164_),
    .B1(net264));
 sg13g2_o21ai_1 _2065_ (.B1(net346),
    .Y(_0402_),
    .A1(net221),
    .A2(net220));
 sg13g2_a21oi_1 _2066_ (.A1(_0814_),
    .A2(_0402_),
    .Y(_0165_),
    .B1(net264));
 sg13g2_o21ai_1 _2067_ (.B1(net399),
    .Y(_0403_),
    .A1(net221),
    .A2(net220));
 sg13g2_a21oi_1 _2068_ (.A1(_0789_),
    .A2(_0403_),
    .Y(_0166_),
    .B1(net264));
 sg13g2_or2_2 _2069_ (.X(_0404_),
    .B(_0393_),
    .A(_0391_));
 sg13g2_a21oi_2 _2070_ (.B1(_0404_),
    .Y(_0405_),
    .A2(_0762_),
    .A1(_0058_));
 sg13g2_a21o_2 _2071_ (.A2(_0762_),
    .A1(_0058_),
    .B1(_0404_),
    .X(_0406_));
 sg13g2_nor3_1 _2072_ (.A(net437),
    .B(_0685_),
    .C(_0406_),
    .Y(_0407_));
 sg13g2_nor2_2 _2073_ (.A(net261),
    .B(_0405_),
    .Y(_0408_));
 sg13g2_a21o_1 _2074_ (.A2(net217),
    .A1(net437),
    .B1(_0407_),
    .X(_0169_));
 sg13g2_o21ai_1 _2075_ (.B1(net271),
    .Y(_0409_),
    .A1(net258),
    .A2(\counter.oled_driver.mc_exec.state_r[6] ));
 sg13g2_nor2_2 _2076_ (.A(_0058_),
    .B(_0409_),
    .Y(_0410_));
 sg13g2_nor2b_2 _2077_ (.A(_0404_),
    .B_N(_0410_),
    .Y(_0411_));
 sg13g2_nand2b_2 _2078_ (.Y(_0412_),
    .B(_0410_),
    .A_N(_0404_));
 sg13g2_nand2_1 _2079_ (.Y(_0413_),
    .A(_0673_),
    .B(_0411_));
 sg13g2_nor2_2 _2080_ (.A(_0408_),
    .B(_0410_),
    .Y(_0414_));
 sg13g2_o21ai_1 _2081_ (.B1(net369),
    .Y(_0415_),
    .A1(\counter.oled_driver.mc_exec.delay_cnt[0] ),
    .A2(_0406_));
 sg13g2_o21ai_1 _2082_ (.B1(_0413_),
    .Y(_0170_),
    .A1(_0414_),
    .A2(net370));
 sg13g2_and2_1 _2083_ (.A(_0049_),
    .B(_0673_),
    .X(_0416_));
 sg13g2_xor2_1 _2084_ (.B(_0673_),
    .A(_0049_),
    .X(_0417_));
 sg13g2_nand2_1 _2085_ (.Y(_0418_),
    .A(net284),
    .B(net217));
 sg13g2_o21ai_1 _2086_ (.B1(_0418_),
    .Y(_0171_),
    .A1(_0412_),
    .A2(_0417_));
 sg13g2_and3_1 _2087_ (.X(_0419_),
    .A(net343),
    .B(_0405_),
    .C(_0416_));
 sg13g2_a21oi_1 _2088_ (.A1(_0405_),
    .A2(_0416_),
    .Y(_0420_),
    .B1(net343));
 sg13g2_nor3_1 _2089_ (.A(_0414_),
    .B(_0419_),
    .C(net344),
    .Y(_0172_));
 sg13g2_xor2_1 _2090_ (.B(_0674_),
    .A(_0050_),
    .X(_0421_));
 sg13g2_nand2_1 _2091_ (.Y(_0422_),
    .A(net189),
    .B(net217));
 sg13g2_o21ai_1 _2092_ (.B1(_0422_),
    .Y(_0173_),
    .A1(_0412_),
    .A2(_0421_));
 sg13g2_nand3_1 _2093_ (.B(_0674_),
    .C(_0405_),
    .A(_0050_),
    .Y(_0423_));
 sg13g2_xor2_1 _2094_ (.B(_0423_),
    .A(net416),
    .X(_0424_));
 sg13g2_nor2_1 _2095_ (.A(_0414_),
    .B(net417),
    .Y(_0174_));
 sg13g2_xor2_1 _2096_ (.B(_0676_),
    .A(_0051_),
    .X(_0425_));
 sg13g2_nand2_1 _2097_ (.Y(_0426_),
    .A(net176),
    .B(net217));
 sg13g2_o21ai_1 _2098_ (.B1(_0426_),
    .Y(_0175_),
    .A1(_0412_),
    .A2(_0425_));
 sg13g2_nand3_1 _2099_ (.B(_0676_),
    .C(_0405_),
    .A(_0051_),
    .Y(_0427_));
 sg13g2_xor2_1 _2100_ (.B(_0427_),
    .A(net423),
    .X(_0428_));
 sg13g2_nor2_1 _2101_ (.A(_0414_),
    .B(net424),
    .Y(_0176_));
 sg13g2_nor3_1 _2102_ (.A(net452),
    .B(_0678_),
    .C(_0406_),
    .Y(_0429_));
 sg13g2_o21ai_1 _2103_ (.B1(net452),
    .Y(_0430_),
    .A1(_0678_),
    .A2(_0406_));
 sg13g2_nor2b_1 _2104_ (.A(_0429_),
    .B_N(_0430_),
    .Y(_0431_));
 sg13g2_nor2_1 _2105_ (.A(_0414_),
    .B(_0431_),
    .Y(_0177_));
 sg13g2_xnor2_1 _2106_ (.Y(_0432_),
    .A(net367),
    .B(_0429_));
 sg13g2_nor2_1 _2107_ (.A(_0414_),
    .B(net368),
    .Y(_0178_));
 sg13g2_nor2_1 _2108_ (.A(_0585_),
    .B(_0679_),
    .Y(_0433_));
 sg13g2_xnor2_1 _2109_ (.Y(_0434_),
    .A(_0052_),
    .B(_0679_));
 sg13g2_nand2_1 _2110_ (.Y(_0435_),
    .A(net174),
    .B(_0408_));
 sg13g2_o21ai_1 _2111_ (.B1(_0435_),
    .Y(_0179_),
    .A1(_0412_),
    .A2(_0434_));
 sg13g2_xnor2_1 _2112_ (.Y(_0436_),
    .A(net350),
    .B(_0433_));
 sg13g2_o21ai_1 _2113_ (.B1(_0396_),
    .Y(_0437_),
    .A1(_0058_),
    .A2(_0436_));
 sg13g2_nor2_1 _2114_ (.A(_0406_),
    .B(_0409_),
    .Y(_0438_));
 sg13g2_a22oi_1 _2115_ (.Y(_0439_),
    .B1(_0437_),
    .B2(_0438_),
    .A2(net217),
    .A1(net350));
 sg13g2_inv_1 _2116_ (.Y(_0180_),
    .A(net351));
 sg13g2_nor3_2 _2117_ (.A(_0056_),
    .B(_0406_),
    .C(_0409_),
    .Y(_0440_));
 sg13g2_nand3_1 _2118_ (.B(net230),
    .C(_0440_),
    .A(_0034_),
    .Y(_0441_));
 sg13g2_xor2_1 _2119_ (.B(_0680_),
    .A(net427),
    .X(_0442_));
 sg13g2_a22oi_1 _2120_ (.Y(_0443_),
    .B1(_0411_),
    .B2(_0442_),
    .A2(net217),
    .A1(net427));
 sg13g2_nand2_1 _2121_ (.Y(_0181_),
    .A(_0441_),
    .B(net428));
 sg13g2_nor2_1 _2122_ (.A(_0681_),
    .B(_0412_),
    .Y(_0444_));
 sg13g2_o21ai_1 _2123_ (.B1(net204),
    .Y(_0445_),
    .A1(net217),
    .A2(_0444_));
 sg13g2_nor3_2 _2124_ (.A(_0631_),
    .B(_0645_),
    .C(_0404_),
    .Y(_0446_));
 sg13g2_a21oi_1 _2125_ (.A1(_0682_),
    .A2(_0411_),
    .Y(_0447_),
    .B1(_0446_));
 sg13g2_nand2_1 _2126_ (.Y(_0182_),
    .A(_0445_),
    .B(_0447_));
 sg13g2_xor2_1 _2127_ (.B(_0682_),
    .A(_0053_),
    .X(_0448_));
 sg13g2_a22oi_1 _2128_ (.Y(_0449_),
    .B1(_0440_),
    .B2(_0643_),
    .A2(_0408_),
    .A1(net391));
 sg13g2_o21ai_1 _2129_ (.B1(net392),
    .Y(_0183_),
    .A1(_0412_),
    .A2(_0448_));
 sg13g2_nand3_1 _2130_ (.B(_0682_),
    .C(_0405_),
    .A(_0053_),
    .Y(_0450_));
 sg13g2_xor2_1 _2131_ (.B(_0450_),
    .A(net444),
    .X(_0451_));
 sg13g2_nand4_1 _2132_ (.B(net258),
    .C(_0641_),
    .A(net271),
    .Y(_0452_),
    .D(_0405_));
 sg13g2_o21ai_1 _2133_ (.B1(_0452_),
    .Y(_0184_),
    .A1(_0414_),
    .A2(net445));
 sg13g2_a21o_1 _2134_ (.A2(_0683_),
    .A1(_0682_),
    .B1(net306),
    .X(_0453_));
 sg13g2_a21oi_1 _2135_ (.A1(_0684_),
    .A2(_0453_),
    .Y(_0454_),
    .B1(_0412_));
 sg13g2_a22oi_1 _2136_ (.Y(_0455_),
    .B1(_0440_),
    .B2(_0639_),
    .A2(net217),
    .A1(net339));
 sg13g2_nand2b_1 _2137_ (.Y(_0185_),
    .B(net340),
    .A_N(_0454_));
 sg13g2_a21oi_1 _2138_ (.A1(_0033_),
    .A2(net229),
    .Y(_0456_),
    .B1(net256));
 sg13g2_nor2b_1 _2139_ (.A(\counter.oled_driver.spi_data[0] ),
    .B_N(net253),
    .Y(_0457_));
 sg13g2_nor3_1 _2140_ (.A(net225),
    .B(_0456_),
    .C(_0457_),
    .Y(_0458_));
 sg13g2_a21o_1 _2141_ (.A2(net223),
    .A1(net291),
    .B1(_0458_),
    .X(_0186_));
 sg13g2_a21o_1 _2142_ (.A2(_0723_),
    .A1(net388),
    .B1(net263),
    .X(_0459_));
 sg13g2_nor3_1 _2143_ (.A(_0553_),
    .B(net223),
    .C(_0459_),
    .Y(_0187_));
 sg13g2_o21ai_1 _2144_ (.B1(net280),
    .Y(_0460_),
    .A1(net312),
    .A2(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[0] ));
 sg13g2_a21oi_1 _2145_ (.A1(net312),
    .A2(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[0] ),
    .Y(_0188_),
    .B1(_0460_));
 sg13g2_nand3_1 _2146_ (.B(net312),
    .C(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[0] ),
    .A(net432),
    .Y(_0461_));
 sg13g2_a21oi_1 _2147_ (.A1(net312),
    .A2(net451),
    .Y(_0462_),
    .B1(net432));
 sg13g2_nor2_1 _2148_ (.A(_0459_),
    .B(_0462_),
    .Y(_0463_));
 sg13g2_and2_1 _2149_ (.A(net433),
    .B(_0463_),
    .X(_0189_));
 sg13g2_xor2_1 _2150_ (.B(net433),
    .A(net388),
    .X(_0464_));
 sg13g2_nor2_1 _2151_ (.A(_0459_),
    .B(_0464_),
    .Y(_0190_));
 sg13g2_o21ai_1 _2152_ (.B1(_0729_),
    .Y(_0465_),
    .A1(_0739_),
    .A2(_0740_));
 sg13g2_nor3_1 _2153_ (.A(\counter.oled_csn_out ),
    .B(net263),
    .C(_0465_),
    .Y(_0466_));
 sg13g2_nand2_1 _2154_ (.Y(_0467_),
    .A(net193),
    .B(net347));
 sg13g2_a21oi_1 _2155_ (.A1(_0465_),
    .A2(_0467_),
    .Y(_0191_),
    .B1(_0466_));
 sg13g2_a21oi_1 _2156_ (.A1(\counter.oled_driver.spi_driver.state_r[0] ),
    .A2(_0728_),
    .Y(_0468_),
    .B1(net193));
 sg13g2_a221oi_1 _2157_ (.B2(net229),
    .C1(_0729_),
    .B1(_0041_),
    .A1(net256),
    .Y(_0469_),
    .A2(\counter.oled_driver.spi_deactivate_cs ));
 sg13g2_nor3_1 _2158_ (.A(net264),
    .B(net194),
    .C(_0469_),
    .Y(_0192_));
 sg13g2_xnor2_1 _2159_ (.Y(_0470_),
    .A(net259),
    .B(net408));
 sg13g2_nor2_1 _2160_ (.A(net239),
    .B(net409),
    .Y(_0213_));
 sg13g2_nand2_1 _2161_ (.Y(_0471_),
    .A(net227),
    .B(_0702_));
 sg13g2_and3_1 _2162_ (.X(_0472_),
    .A(net259),
    .B(net209),
    .C(\counter.counter_ref.digit_0.digit_out[0] ));
 sg13g2_a21oi_1 _2163_ (.A1(net259),
    .A2(\counter.counter_ref.digit_0.digit_out[0] ),
    .Y(_0473_),
    .B1(net209));
 sg13g2_nor3_1 _2164_ (.A(_0471_),
    .B(_0472_),
    .C(net210),
    .Y(_0214_));
 sg13g2_nor2_1 _2165_ (.A(net377),
    .B(_0472_),
    .Y(_0474_));
 sg13g2_and2_1 _2166_ (.A(net377),
    .B(_0472_),
    .X(_0475_));
 sg13g2_nor3_1 _2167_ (.A(net239),
    .B(net378),
    .C(_0475_),
    .Y(_0215_));
 sg13g2_xnor2_1 _2168_ (.Y(_0476_),
    .A(net331),
    .B(_0475_));
 sg13g2_nor2_1 _2169_ (.A(_0471_),
    .B(net332),
    .Y(_0216_));
 sg13g2_nor2_1 _2170_ (.A(net168),
    .B(_0703_),
    .Y(_0477_));
 sg13g2_a21oi_1 _2171_ (.A1(net168),
    .A2(_0471_),
    .Y(_0217_),
    .B1(_0477_));
 sg13g2_nor3_1 _2172_ (.A(_0532_),
    .B(net239),
    .C(_0702_),
    .Y(_0478_));
 sg13g2_a21oi_1 _2173_ (.A1(_0697_),
    .A2(_0478_),
    .Y(_0479_),
    .B1(net303));
 sg13g2_and2_1 _2174_ (.A(net303),
    .B(_0478_),
    .X(_0480_));
 sg13g2_nor3_1 _2175_ (.A(net239),
    .B(net304),
    .C(_0480_),
    .Y(_0218_));
 sg13g2_and2_1 _2176_ (.A(net422),
    .B(_0480_),
    .X(_0481_));
 sg13g2_o21ai_1 _2177_ (.B1(net227),
    .Y(_0482_),
    .A1(net422),
    .A2(_0480_));
 sg13g2_nor2_1 _2178_ (.A(_0481_),
    .B(_0482_),
    .Y(_0219_));
 sg13g2_o21ai_1 _2179_ (.B1(net227),
    .Y(_0483_),
    .A1(net191),
    .A2(_0481_));
 sg13g2_a221oi_1 _2180_ (.B2(net191),
    .C1(_0483_),
    .B1(_0481_),
    .A1(_0698_),
    .Y(_0220_),
    .A2(_0703_));
 sg13g2_nor2_1 _2181_ (.A(net353),
    .B(_0704_),
    .Y(_0484_));
 sg13g2_and2_1 _2182_ (.A(net353),
    .B(_0704_),
    .X(_0485_));
 sg13g2_nor2_1 _2183_ (.A(net240),
    .B(_0485_),
    .Y(_0486_));
 sg13g2_nor3_1 _2184_ (.A(net239),
    .B(_0484_),
    .C(_0485_),
    .Y(_0221_));
 sg13g2_nor2b_1 _2185_ (.A(_0695_),
    .B_N(_0694_),
    .Y(_0487_));
 sg13g2_a22oi_1 _2186_ (.Y(_0488_),
    .B1(_0487_),
    .B2(_0704_),
    .A2(_0486_),
    .A1(net359));
 sg13g2_inv_1 _2187_ (.Y(_0222_),
    .A(_0488_));
 sg13g2_a21oi_1 _2188_ (.A1(\counter.counter_ref.digits_out[9] ),
    .A2(_0485_),
    .Y(_0489_),
    .B1(net201));
 sg13g2_and3_1 _2189_ (.X(_0490_),
    .A(net201),
    .B(net359),
    .C(_0485_));
 sg13g2_nor3_1 _2190_ (.A(net239),
    .B(net202),
    .C(_0490_),
    .Y(_0223_));
 sg13g2_o21ai_1 _2191_ (.B1(net228),
    .Y(_0491_),
    .A1(net425),
    .A2(_0490_));
 sg13g2_a21oi_1 _2192_ (.A1(net425),
    .A2(_0490_),
    .Y(_0492_),
    .B1(_0715_));
 sg13g2_nor2b_1 _2193_ (.A(_0491_),
    .B_N(_0492_),
    .Y(_0224_));
 sg13g2_nand2_1 _2194_ (.Y(_0493_),
    .A(net390),
    .B(_0705_));
 sg13g2_nand3_1 _2195_ (.B(net259),
    .C(_0720_),
    .A(net390),
    .Y(_0494_));
 sg13g2_nand2_1 _2196_ (.Y(_0495_),
    .A(net227),
    .B(_0494_));
 sg13g2_nor2_1 _2197_ (.A(net390),
    .B(_0705_),
    .Y(_0496_));
 sg13g2_nor2_1 _2198_ (.A(_0495_),
    .B(_0496_),
    .Y(_0225_));
 sg13g2_nor2_1 _2199_ (.A(net448),
    .B(_0494_),
    .Y(_0497_));
 sg13g2_nand3_1 _2200_ (.B(_0709_),
    .C(_0497_),
    .A(net227),
    .Y(_0498_));
 sg13g2_o21ai_1 _2201_ (.B1(_0498_),
    .Y(_0226_),
    .A1(_0530_),
    .A2(_0495_));
 sg13g2_nor2_1 _2202_ (.A(_0530_),
    .B(_0493_),
    .Y(_0499_));
 sg13g2_a21oi_1 _2203_ (.A1(net439),
    .A2(_0499_),
    .Y(_0500_),
    .B1(net239));
 sg13g2_o21ai_1 _2204_ (.B1(_0500_),
    .Y(_0501_),
    .A1(net439),
    .A2(_0499_));
 sg13g2_inv_1 _2205_ (.Y(_0227_),
    .A(_0501_));
 sg13g2_a21oi_1 _2206_ (.A1(\counter.counter_ref.digits_out[14] ),
    .A2(_0499_),
    .Y(_0502_),
    .B1(net288));
 sg13g2_nor3_1 _2207_ (.A(\counter.counter_ref.digits_out[13] ),
    .B(_0709_),
    .C(_0493_),
    .Y(_0503_));
 sg13g2_nor3_2 _2208_ (.A(\counter.counter_ref.digits_out[13] ),
    .B(_0709_),
    .C(_0494_),
    .Y(_0504_));
 sg13g2_and3_1 _2209_ (.X(_0505_),
    .A(net288),
    .B(\counter.counter_ref.digits_out[14] ),
    .C(_0499_));
 sg13g2_nor4_1 _2210_ (.A(net242),
    .B(net289),
    .C(_0504_),
    .D(_0505_),
    .Y(_0228_));
 sg13g2_or2_1 _2211_ (.X(_0506_),
    .B(_0504_),
    .A(net457));
 sg13g2_nand2_1 _2212_ (.Y(_0507_),
    .A(net457),
    .B(_0503_));
 sg13g2_and3_1 _2213_ (.X(_0229_),
    .A(net227),
    .B(_0506_),
    .C(_0507_));
 sg13g2_nand3_1 _2214_ (.B(net228),
    .C(_0507_),
    .A(net328),
    .Y(_0508_));
 sg13g2_nand2_1 _2215_ (.Y(_0509_),
    .A(net227),
    .B(_0711_));
 sg13g2_or2_1 _2216_ (.X(_0510_),
    .B(_0507_),
    .A(net328));
 sg13g2_o21ai_1 _2217_ (.B1(net329),
    .Y(_0230_),
    .A1(_0509_),
    .A2(_0510_));
 sg13g2_and2_1 _2218_ (.A(\counter.counter_ref.digits_out[17] ),
    .B(\counter.counter_ref.digits_out[16] ),
    .X(_0511_));
 sg13g2_a21oi_1 _2219_ (.A1(_0504_),
    .A2(_0511_),
    .Y(_0512_),
    .B1(net282));
 sg13g2_and3_1 _2220_ (.X(_0513_),
    .A(net282),
    .B(_0504_),
    .C(_0511_));
 sg13g2_nor3_1 _2221_ (.A(net240),
    .B(net283),
    .C(_0513_),
    .Y(_0231_));
 sg13g2_nor2_1 _2222_ (.A(net382),
    .B(_0513_),
    .Y(_0514_));
 sg13g2_nor2_1 _2223_ (.A(_0711_),
    .B(_0510_),
    .Y(_0515_));
 sg13g2_and2_1 _2224_ (.A(net382),
    .B(_0513_),
    .X(_0516_));
 sg13g2_nor4_1 _2225_ (.A(net240),
    .B(_0514_),
    .C(_0515_),
    .D(_0516_),
    .Y(_0232_));
 sg13g2_nor2_1 _2226_ (.A(net314),
    .B(_0515_),
    .Y(_0517_));
 sg13g2_nor3_1 _2227_ (.A(_0529_),
    .B(_0711_),
    .C(_0510_),
    .Y(_0518_));
 sg13g2_nor3_1 _2228_ (.A(net240),
    .B(net315),
    .C(_0518_),
    .Y(_0233_));
 sg13g2_a21oi_1 _2229_ (.A1(_0708_),
    .A2(_0518_),
    .Y(_0519_),
    .B1(net325));
 sg13g2_and2_1 _2230_ (.A(net325),
    .B(_0518_),
    .X(_0520_));
 sg13g2_nor3_1 _2231_ (.A(net240),
    .B(net326),
    .C(_0520_),
    .Y(_0234_));
 sg13g2_nor2_1 _2232_ (.A(net323),
    .B(_0520_),
    .Y(_0521_));
 sg13g2_and2_1 _2233_ (.A(net323),
    .B(_0520_),
    .X(_0522_));
 sg13g2_nor3_1 _2234_ (.A(net240),
    .B(net324),
    .C(_0522_),
    .Y(_0235_));
 sg13g2_nor2_1 _2235_ (.A(net375),
    .B(_0522_),
    .Y(_0523_));
 sg13g2_and2_1 _2236_ (.A(net375),
    .B(_0522_),
    .X(_0524_));
 sg13g2_nor4_1 _2237_ (.A(net240),
    .B(_0713_),
    .C(_0523_),
    .D(_0524_),
    .Y(_0236_));
 sg13g2_o21ai_1 _2238_ (.B1(_0719_),
    .Y(_0525_),
    .A1(net259),
    .A2(_0577_));
 sg13g2_nor2_1 _2239_ (.A(net166),
    .B(net235),
    .Y(_0526_));
 sg13g2_o21ai_1 _2240_ (.B1(net273),
    .Y(_0527_),
    .A1(net376),
    .A2(_0525_));
 sg13g2_a21oi_1 _2241_ (.A1(_0525_),
    .A2(_0526_),
    .Y(_0237_),
    .B1(_0527_));
 sg13g2_a21o_1 _2242_ (.A2(_0939_),
    .A1(_0123_),
    .B1(_0124_),
    .X(_0528_));
 sg13g2_a21oi_1 _2243_ (.A1(_0927_),
    .A2(_0942_),
    .Y(_0238_),
    .B1(_0528_));
 sg13g2_inv_1 _2244_ (.Y(_0080_),
    .A(net243));
 sg13g2_inv_1 _2245_ (.Y(_0081_),
    .A(net243));
 sg13g2_inv_1 _2246_ (.Y(_0082_),
    .A(net243));
 sg13g2_inv_1 _2247_ (.Y(_0083_),
    .A(net241));
 sg13g2_inv_1 _2248_ (.Y(_0084_),
    .A(net241));
 sg13g2_inv_1 _2249_ (.Y(_0085_),
    .A(net241));
 sg13g2_inv_1 _2250_ (.Y(_0086_),
    .A(net241));
 sg13g2_inv_1 _2251_ (.Y(_0087_),
    .A(net242));
 sg13g2_inv_1 _2252_ (.Y(_0088_),
    .A(net241));
 sg13g2_inv_1 _2253_ (.Y(_0089_),
    .A(net241));
 sg13g2_inv_1 _2254_ (.Y(_0090_),
    .A(net241));
 sg13g2_inv_1 _2255_ (.Y(_0091_),
    .A(net241));
 sg13g2_inv_1 _2256_ (.Y(_0092_),
    .A(net244));
 sg13g2_inv_1 _2257_ (.Y(_0093_),
    .A(net244));
 sg13g2_inv_1 _2258_ (.Y(_0094_),
    .A(net244));
 sg13g2_inv_1 _2259_ (.Y(_0095_),
    .A(net244));
 sg13g2_inv_1 _2260_ (.Y(_0096_),
    .A(net244));
 sg13g2_inv_1 _2261_ (.Y(_0097_),
    .A(net244));
 sg13g2_inv_1 _2262_ (.Y(_0098_),
    .A(net243));
 sg13g2_inv_1 _2263_ (.Y(_0099_),
    .A(net243));
 sg13g2_inv_1 _2264_ (.Y(_0100_),
    .A(net243));
 sg13g2_inv_1 _2265_ (.Y(_0101_),
    .A(net243));
 sg13g2_inv_1 _2266_ (.Y(_0102_),
    .A(net244));
 sg13g2_dfrbp_1 _2267_ (.CLK(net269),
    .RESET_B(_0079_),
    .D(_0103_),
    .Q_N(_1119_),
    .Q(\counter.cnt_x_digits[20] ));
 sg13g2_dfrbp_1 _2268_ (.CLK(net269),
    .RESET_B(_0080_),
    .D(_0104_),
    .Q_N(_1118_),
    .Q(\counter.cnt_x_digits[21] ));
 sg13g2_dfrbp_1 _2269_ (.CLK(net268),
    .RESET_B(_0081_),
    .D(_0105_),
    .Q_N(_1117_),
    .Q(\counter.cnt_x_digits[22] ));
 sg13g2_dfrbp_1 _2270_ (.CLK(net268),
    .RESET_B(_0082_),
    .D(_0106_),
    .Q_N(_1116_),
    .Q(\counter.cnt_x_digits[23] ));
 sg13g2_dfrbp_1 _2271_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net79),
    .D(_0107_),
    .Q_N(_1115_),
    .Q(\counter.streamer.graphical_decoder.pattern_adg[1] ));
 sg13g2_dfrbp_1 _2272_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net23),
    .D(_0108_),
    .Q_N(_1120_),
    .Q(\counter.streamer.graphical_decoder.pattern_adg[4] ));
 sg13g2_dfrbp_1 _2273_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net24),
    .D(net167),
    .Q_N(_1121_),
    .Q(\counter.state[0] ));
 sg13g2_dfrbp_1 _2274_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net25),
    .D(net188),
    .Q_N(_0059_),
    .Q(\counter.state[1] ));
 sg13g2_dfrbp_1 _2275_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net26),
    .D(net181),
    .Q_N(_1122_),
    .Q(\counter.cnt_ref_enable ));
 sg13g2_dfrbp_1 _2276_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net27),
    .D(net208),
    .Q_N(_1123_),
    .Q(\counter.oled_driver.mc_exec.spi_tx_trigger_out ));
 sg13g2_dfrbp_1 _2277_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net28),
    .D(net450),
    .Q_N(_0056_),
    .Q(\counter.oled_driver.mc_exec.state_r[2] ));
 sg13g2_dfrbp_1 _2278_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net29),
    .D(net308),
    .Q_N(_0057_),
    .Q(\counter.oled_driver.mc_exec.state_r[3] ));
 sg13g2_dfrbp_1 _2279_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net30),
    .D(net443),
    .Q_N(_0054_),
    .Q(\counter.oled_driver.mc_exec.procedure_done_out ));
 sg13g2_dfrbp_1 _2280_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net31),
    .D(net200),
    .Q_N(_1124_),
    .Q(\counter.oled_driver.mc_exec.state_r[5] ));
 sg13g2_dfrbp_1 _2281_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net32),
    .D(_0020_),
    .Q_N(_0058_),
    .Q(\counter.oled_driver.mc_exec.state_r[6] ));
 sg13g2_dfrbp_1 _2282_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net33),
    .D(_0000_),
    .Q_N(_1125_),
    .Q(_0033_));
 sg13g2_dfrbp_1 _2283_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net34),
    .D(_0001_),
    .Q_N(_1126_),
    .Q(_0034_));
 sg13g2_dfrbp_1 _2284_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net35),
    .D(_0002_),
    .Q_N(_1127_),
    .Q(_0035_));
 sg13g2_dfrbp_1 _2285_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net36),
    .D(_0003_),
    .Q_N(_1128_),
    .Q(_0036_));
 sg13g2_dfrbp_1 _2286_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net37),
    .D(_0004_),
    .Q_N(_1129_),
    .Q(_0037_));
 sg13g2_dfrbp_1 _2287_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net38),
    .D(_0005_),
    .Q_N(_1130_),
    .Q(_0038_));
 sg13g2_dfrbp_1 _2288_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net39),
    .D(_0006_),
    .Q_N(_1131_),
    .Q(_0039_));
 sg13g2_dfrbp_1 _2289_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net40),
    .D(_0007_),
    .Q_N(_1132_),
    .Q(_0040_));
 sg13g2_dfrbp_1 _2290_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net85),
    .D(_0008_),
    .Q_N(_1133_),
    .Q(_0041_));
 sg13g2_dfrbp_1 _2291_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net78),
    .D(_0009_),
    .Q_N(_1114_),
    .Q(_0042_));
 sg13g2_dfrbp_1 _2292_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net77),
    .D(_0109_),
    .Q_N(_1113_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[1] ));
 sg13g2_dfrbp_1 _2293_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net75),
    .D(net302),
    .Q_N(_1112_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[2] ));
 sg13g2_dfrbp_1 _2294_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net74),
    .D(_0111_),
    .Q_N(_1111_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[3] ));
 sg13g2_dfrbp_1 _2295_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net72),
    .D(net335),
    .Q_N(_1110_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[4] ));
 sg13g2_dfrbp_1 _2296_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net70),
    .D(net319),
    .Q_N(_1109_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[5] ));
 sg13g2_dfrbp_1 _2297_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net68),
    .D(_0114_),
    .Q_N(_1108_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[6] ));
 sg13g2_dfrbp_1 _2298_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net67),
    .D(net311),
    .Q_N(_1107_),
    .Q(\counter.oled_driver.oled_mosi_out ));
 sg13g2_dfrbp_1 _2299_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net65),
    .D(net295),
    .Q_N(_1106_),
    .Q(\counter.oled_driver.mc_exec.procedure_offset_in[0] ));
 sg13g2_dfrbp_1 _2300_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net63),
    .D(net183),
    .Q_N(_0068_),
    .Q(\counter.streamer.digit_cnt_r[0] ));
 sg13g2_dfrbp_1 _2301_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net61),
    .D(_0118_),
    .Q_N(_0071_),
    .Q(\counter.streamer.digit_cnt_r[1] ));
 sg13g2_dfrbp_1 _2302_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net60),
    .D(net454),
    .Q_N(_0069_),
    .Q(\counter.streamer.digit_cnt_r[2] ));
 sg13g2_dfrbp_1 _2303_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net58),
    .D(_0120_),
    .Q_N(_0045_),
    .Q(\counter.streamer.graphical_decoder.index_x_in[0] ));
 sg13g2_dfrbp_1 _2304_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net56),
    .D(_0121_),
    .Q_N(_0043_),
    .Q(\counter.streamer.graphical_decoder.index_x_in[1] ));
 sg13g2_dfrbp_1 _2305_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net54),
    .D(_0122_),
    .Q_N(_0066_),
    .Q(\counter.streamer.graphical_decoder.index_x_in[2] ));
 sg13g2_dfrbp_1 _2306_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net53),
    .D(_0123_),
    .Q_N(_1105_),
    .Q(\counter.streamer.graphical_decoder.index_x_in[3] ));
 sg13g2_dfrbp_1 _2307_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net51),
    .D(net462),
    .Q_N(_0065_),
    .Q(\counter.streamer.graphical_decoder.index_x_in[4] ));
 sg13g2_dfrbp_1 _2308_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net49),
    .D(_0125_),
    .Q_N(_0077_),
    .Q(\counter.streamer.graphical_decoder.index_y_in[0] ));
 sg13g2_dfrbp_1 _2309_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net47),
    .D(_0126_),
    .Q_N(_0076_),
    .Q(\counter.streamer.graphical_decoder.index_y_in[1] ));
 sg13g2_dfrbp_1 _2310_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net46),
    .D(_0127_),
    .Q_N(_1104_),
    .Q(\counter.streamer.digits_r[0] ));
 sg13g2_dfrbp_1 _2311_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net44),
    .D(_0128_),
    .Q_N(_1103_),
    .Q(\counter.streamer.digits_r[1] ));
 sg13g2_dfrbp_1 _2312_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net42),
    .D(_0129_),
    .Q_N(_1102_),
    .Q(\counter.streamer.digits_r[2] ));
 sg13g2_dfrbp_1 _2313_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net22),
    .D(_0130_),
    .Q_N(_0072_),
    .Q(\counter.streamer.digits_r[3] ));
 sg13g2_dfrbp_1 _2314_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net20),
    .D(_0131_),
    .Q_N(_1101_),
    .Q(\counter.streamer.digits_r[4] ));
 sg13g2_dfrbp_1 _2315_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net18),
    .D(_0132_),
    .Q_N(_1100_),
    .Q(\counter.streamer.digits_r[5] ));
 sg13g2_dfrbp_1 _2316_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net163),
    .D(_0133_),
    .Q_N(_1099_),
    .Q(\counter.streamer.digits_r[6] ));
 sg13g2_dfrbp_1 _2317_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net161),
    .D(_0134_),
    .Q_N(_0073_),
    .Q(\counter.streamer.digits_r[7] ));
 sg13g2_dfrbp_1 _2318_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net156),
    .D(_0135_),
    .Q_N(_1098_),
    .Q(\counter.streamer.digits_r[8] ));
 sg13g2_dfrbp_1 _2319_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net154),
    .D(_0136_),
    .Q_N(_1097_),
    .Q(\counter.streamer.digits_r[9] ));
 sg13g2_dfrbp_1 _2320_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net152),
    .D(_0137_),
    .Q_N(_1096_),
    .Q(\counter.streamer.digits_r[10] ));
 sg13g2_dfrbp_1 _2321_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net150),
    .D(_0138_),
    .Q_N(_0074_),
    .Q(\counter.streamer.digits_r[11] ));
 sg13g2_dfrbp_1 _2322_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net148),
    .D(_0139_),
    .Q_N(_1095_),
    .Q(\counter.streamer.digits_r[12] ));
 sg13g2_dfrbp_1 _2323_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net146),
    .D(_0140_),
    .Q_N(_1094_),
    .Q(\counter.streamer.digits_r[13] ));
 sg13g2_dfrbp_1 _2324_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net144),
    .D(_0141_),
    .Q_N(_1093_),
    .Q(\counter.streamer.digits_r[14] ));
 sg13g2_dfrbp_1 _2325_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net142),
    .D(_0142_),
    .Q_N(_0075_),
    .Q(\counter.streamer.digits_r[15] ));
 sg13g2_dfrbp_1 _2326_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net140),
    .D(_0143_),
    .Q_N(_1092_),
    .Q(\counter.streamer.digits_r[16] ));
 sg13g2_dfrbp_1 _2327_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net138),
    .D(_0144_),
    .Q_N(_1091_),
    .Q(\counter.streamer.digits_r[17] ));
 sg13g2_dfrbp_1 _2328_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net136),
    .D(_0145_),
    .Q_N(_1090_),
    .Q(\counter.streamer.digits_r[18] ));
 sg13g2_dfrbp_1 _2329_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net135),
    .D(_0146_),
    .Q_N(_1089_),
    .Q(\counter.streamer.digits_r[19] ));
 sg13g2_dfrbp_1 _2330_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net133),
    .D(_0147_),
    .Q_N(_1088_),
    .Q(\counter.streamer.digits_r[20] ));
 sg13g2_dfrbp_1 _2331_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net132),
    .D(_0148_),
    .Q_N(_1087_),
    .Q(\counter.streamer.digits_r[21] ));
 sg13g2_dfrbp_1 _2332_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net130),
    .D(_0149_),
    .Q_N(_1086_),
    .Q(\counter.streamer.digits_r[22] ));
 sg13g2_dfrbp_1 _2333_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net129),
    .D(_0150_),
    .Q_N(_1085_),
    .Q(\counter.streamer.digits_r[23] ));
 sg13g2_dfrbp_1 _2334_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net127),
    .D(_0151_),
    .Q_N(_1084_),
    .Q(\counter.oled_driver.spi_data[0] ));
 sg13g2_dfrbp_1 _2335_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net126),
    .D(_0152_),
    .Q_N(_1083_),
    .Q(\counter.oled_driver.spi_data[1] ));
 sg13g2_dfrbp_1 _2336_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net124),
    .D(net173),
    .Q_N(_0046_),
    .Q(\counter.oled_driver.spi_data[2] ));
 sg13g2_dfrbp_1 _2337_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net123),
    .D(_0154_),
    .Q_N(_1082_),
    .Q(\counter.oled_driver.spi_data[3] ));
 sg13g2_dfrbp_1 _2338_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net121),
    .D(_0155_),
    .Q_N(_0047_),
    .Q(\counter.oled_driver.spi_data[4] ));
 sg13g2_dfrbp_1 _2339_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net120),
    .D(net287),
    .Q_N(_1081_),
    .Q(\counter.oled_driver.spi_data[5] ));
 sg13g2_dfrbp_1 _2340_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net112),
    .D(_0157_),
    .Q_N(_1080_),
    .Q(\counter.oled_driver.spi_data[6] ));
 sg13g2_dfrbp_1 _2341_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net111),
    .D(net171),
    .Q_N(_0048_),
    .Q(\counter.oled_driver.spi_data[7] ));
 sg13g2_dfrbp_1 _2342_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net109),
    .D(net338),
    .Q_N(_1079_),
    .Q(\counter.oled_driver.mc_exec.oled_vcdn_out ));
 sg13g2_dfrbp_1 _2343_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net108),
    .D(net396),
    .Q_N(_1078_),
    .Q(\counter.oled_driver.mc_exec.oled_vbatn_out ));
 sg13g2_dfrbp_1 _2344_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net86),
    .D(net404),
    .Q_N(_1134_),
    .Q(\counter.oled_driver.mc_exec.oled_rstn_out ));
 sg13g2_dfrbp_1 _2345_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net87),
    .D(net381),
    .Q_N(_1135_),
    .Q(\counter.oled_driver.state_r[0] ));
 sg13g2_dfrbp_1 _2346_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net88),
    .D(net361),
    .Q_N(_1136_),
    .Q(\counter.oled_driver.spi_deactivate_cs ));
 sg13g2_dfrbp_1 _2347_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net89),
    .D(net398),
    .Q_N(_1137_),
    .Q(\counter.oled_driver.state_r[2] ));
 sg13g2_dfrbp_1 _2348_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net90),
    .D(net358),
    .Q_N(_1138_),
    .Q(\counter.oled_driver.mc_exec.procedure_start_in ));
 sg13g2_dfrbp_1 _2349_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net114),
    .D(net297),
    .Q_N(_1139_),
    .Q(\counter.oled_driver.state_r[4] ));
 sg13g2_dfrbp_1 _2350_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net106),
    .D(_0026_),
    .Q_N(_1077_),
    .Q(\counter.oled_driver.ready_out ));
 sg13g2_dfrbp_1 _2351_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net105),
    .D(net386),
    .Q_N(_1076_),
    .Q(\counter.oled_driver.mc_exec.oled_dc_out ));
 sg13g2_dfrbp_1 _2352_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net103),
    .D(_0163_),
    .Q_N(_0064_),
    .Q(\counter.oled_driver.mc_exec.microcode_rom.address[0] ));
 sg13g2_dfrbp_1 _2353_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net102),
    .D(net414),
    .Q_N(_0063_),
    .Q(\counter.oled_driver.mc_exec.microcode_rom.address[1] ));
 sg13g2_dfrbp_1 _2354_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net100),
    .D(_0165_),
    .Q_N(_0060_),
    .Q(\counter.oled_driver.mc_exec.microcode_rom.address[2] ));
 sg13g2_dfrbp_1 _2355_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net99),
    .D(net400),
    .Q_N(_0061_),
    .Q(\counter.oled_driver.mc_exec.microcode_rom.address[3] ));
 sg13g2_dfrbp_1 _2356_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net97),
    .D(_0167_),
    .Q_N(_0062_),
    .Q(\counter.oled_driver.mc_exec.microcode_rom.address[4] ));
 sg13g2_dfrbp_1 _2357_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net96),
    .D(net216),
    .Q_N(_1075_),
    .Q(\counter.oled_driver.mc_exec.microcode_rom.address[5] ));
 sg13g2_dfrbp_1 _2358_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net94),
    .D(_0169_),
    .Q_N(_1074_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[0] ));
 sg13g2_dfrbp_1 _2359_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net93),
    .D(net371),
    .Q_N(_1073_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[1] ));
 sg13g2_dfrbp_1 _2360_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net91),
    .D(net285),
    .Q_N(_0049_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[2] ));
 sg13g2_dfrbp_1 _2361_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net84),
    .D(net345),
    .Q_N(_1072_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[3] ));
 sg13g2_dfrbp_1 _2362_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net82),
    .D(net190),
    .Q_N(_0050_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[4] ));
 sg13g2_dfrbp_1 _2363_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net81),
    .D(_0174_),
    .Q_N(_1071_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[5] ));
 sg13g2_dfrbp_1 _2364_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net76),
    .D(net177),
    .Q_N(_0051_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[6] ));
 sg13g2_dfrbp_1 _2365_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net73),
    .D(_0176_),
    .Q_N(_1070_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[7] ));
 sg13g2_dfrbp_1 _2366_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net69),
    .D(_0177_),
    .Q_N(_1069_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[8] ));
 sg13g2_dfrbp_1 _2367_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net66),
    .D(_0178_),
    .Q_N(_1068_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[9] ));
 sg13g2_dfrbp_1 _2368_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net62),
    .D(net175),
    .Q_N(_0052_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[10] ));
 sg13g2_dfrbp_1 _2369_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net59),
    .D(_0180_),
    .Q_N(_1067_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[11] ));
 sg13g2_dfrbp_1 _2370_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net55),
    .D(net429),
    .Q_N(_1066_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[12] ));
 sg13g2_dfrbp_1 _2371_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net52),
    .D(net205),
    .Q_N(_1065_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[13] ));
 sg13g2_dfrbp_1 _2372_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net48),
    .D(net393),
    .Q_N(_0053_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[14] ));
 sg13g2_dfrbp_1 _2373_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net45),
    .D(net446),
    .Q_N(_1064_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[15] ));
 sg13g2_dfrbp_1 _2374_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net41),
    .D(net341),
    .Q_N(_0055_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[16] ));
 sg13g2_dfrbp_1 _2375_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net19),
    .D(net292),
    .Q_N(_1063_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[0] ));
 sg13g2_dfrbp_1 _2376_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net162),
    .D(net165),
    .Q_N(_0078_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[0] ));
 sg13g2_dfrbp_1 _2377_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net155),
    .D(net313),
    .Q_N(_1062_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[1] ));
 sg13g2_dfrbp_1 _2378_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net151),
    .D(_0189_),
    .Q_N(_1061_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[2] ));
 sg13g2_dfrbp_1 _2379_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net147),
    .D(_0190_),
    .Q_N(_1060_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[3] ));
 sg13g2_dfrbp_1 _2380_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net143),
    .D(net348),
    .Q_N(_1059_),
    .Q(\counter.oled_csn_out ));
 sg13g2_dfrbp_1 _2381_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net115),
    .D(net195),
    .Q_N(_1140_),
    .Q(\counter.oled_driver.spi_driver.deactivate_cs_r ));
 sg13g2_dfrbp_1 _2382_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net116),
    .D(net261),
    .Q_N(_1141_),
    .Q(\counter.oled_driver.mc_exec.state_r[0] ));
 sg13g2_dfrbp_1 _2383_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net117),
    .D(net355),
    .Q_N(_1142_),
    .Q(\counter.oled_driver.sync_stb_in ));
 sg13g2_dfrbp_1 _2384_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net118),
    .D(_0031_),
    .Q_N(_1143_),
    .Q(\counter.oled_driver.write_stb_in ));
 sg13g2_dfrbp_1 _2385_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net119),
    .D(net321),
    .Q_N(_1144_),
    .Q(\counter.streamer.ready_out ));
 sg13g2_dfrbp_1 _2386_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net158),
    .D(net185),
    .Q_N(_1145_),
    .Q(\counter.streamer.state_r[4] ));
 sg13g2_dfrbp_1 _2387_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net139),
    .D(net402),
    .Q_N(_0067_),
    .Q(\counter.streamer.state_r[5] ));
 sg13g2_dfrbp_1 _2388_ (.CLK(net266),
    .RESET_B(_0083_),
    .D(_0193_),
    .Q_N(_1058_),
    .Q(\counter.cnt_x_digits[0] ));
 sg13g2_dfrbp_1 _2389_ (.CLK(net266),
    .RESET_B(_0084_),
    .D(_0194_),
    .Q_N(_1057_),
    .Q(\counter.cnt_x_digits[1] ));
 sg13g2_dfrbp_1 _2390_ (.CLK(net266),
    .RESET_B(_0085_),
    .D(_0195_),
    .Q_N(_1056_),
    .Q(\counter.cnt_x_digits[2] ));
 sg13g2_dfrbp_1 _2391_ (.CLK(net266),
    .RESET_B(_0086_),
    .D(_0196_),
    .Q_N(_1055_),
    .Q(\counter.cnt_x_digits[3] ));
 sg13g2_dfrbp_1 _2392_ (.CLK(net266),
    .RESET_B(_0087_),
    .D(_0197_),
    .Q_N(_1054_),
    .Q(\counter.cnt_x_digits[4] ));
 sg13g2_dfrbp_1 _2393_ (.CLK(net267),
    .RESET_B(_0088_),
    .D(_0198_),
    .Q_N(_1053_),
    .Q(\counter.cnt_x_digits[5] ));
 sg13g2_dfrbp_1 _2394_ (.CLK(net266),
    .RESET_B(_0089_),
    .D(_0199_),
    .Q_N(_1052_),
    .Q(\counter.cnt_x_digits[6] ));
 sg13g2_dfrbp_1 _2395_ (.CLK(net266),
    .RESET_B(_0090_),
    .D(_0200_),
    .Q_N(_1051_),
    .Q(\counter.cnt_x_digits[7] ));
 sg13g2_dfrbp_1 _2396_ (.CLK(net266),
    .RESET_B(_0091_),
    .D(_0201_),
    .Q_N(_1050_),
    .Q(\counter.cnt_x_digits[8] ));
 sg13g2_dfrbp_1 _2397_ (.CLK(net267),
    .RESET_B(_0092_),
    .D(_0202_),
    .Q_N(_1049_),
    .Q(\counter.cnt_x_digits[9] ));
 sg13g2_dfrbp_1 _2398_ (.CLK(net267),
    .RESET_B(_0093_),
    .D(_0203_),
    .Q_N(_1048_),
    .Q(\counter.cnt_x_digits[10] ));
 sg13g2_dfrbp_1 _2399_ (.CLK(net267),
    .RESET_B(_0094_),
    .D(_0204_),
    .Q_N(_1047_),
    .Q(\counter.cnt_x_digits[11] ));
 sg13g2_dfrbp_1 _2400_ (.CLK(net268),
    .RESET_B(_0095_),
    .D(_0205_),
    .Q_N(_1046_),
    .Q(\counter.cnt_x_digits[12] ));
 sg13g2_dfrbp_1 _2401_ (.CLK(net268),
    .RESET_B(_0096_),
    .D(_0206_),
    .Q_N(_1045_),
    .Q(\counter.cnt_x_digits[13] ));
 sg13g2_dfrbp_1 _2402_ (.CLK(net268),
    .RESET_B(_0097_),
    .D(_0207_),
    .Q_N(_1044_),
    .Q(\counter.cnt_x_digits[14] ));
 sg13g2_dfrbp_1 _2403_ (.CLK(net268),
    .RESET_B(_0098_),
    .D(_0208_),
    .Q_N(_1043_),
    .Q(\counter.cnt_x_digits[15] ));
 sg13g2_dfrbp_1 _2404_ (.CLK(net269),
    .RESET_B(_0099_),
    .D(_0209_),
    .Q_N(_1042_),
    .Q(\counter.cnt_x_digits[16] ));
 sg13g2_dfrbp_1 _2405_ (.CLK(net268),
    .RESET_B(_0100_),
    .D(_0210_),
    .Q_N(_1041_),
    .Q(\counter.cnt_x_digits[17] ));
 sg13g2_dfrbp_1 _2406_ (.CLK(net268),
    .RESET_B(_0101_),
    .D(_0211_),
    .Q_N(_1040_),
    .Q(\counter.cnt_x_digits[18] ));
 sg13g2_dfrbp_1 _2407_ (.CLK(net269),
    .RESET_B(_0102_),
    .D(_0212_),
    .Q_N(_1039_),
    .Q(\counter.cnt_x_digits[19] ));
 sg13g2_dfrbp_1 _2408_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net21),
    .D(_0213_),
    .Q_N(_1038_),
    .Q(\counter.counter_ref.digit_0.digit_out[0] ));
 sg13g2_dfrbp_1 _2409_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net157),
    .D(net211),
    .Q_N(_1037_),
    .Q(\counter.counter_ref.digit_0.digit_out[1] ));
 sg13g2_dfrbp_1 _2410_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net149),
    .D(_0215_),
    .Q_N(_1036_),
    .Q(\counter.counter_ref.digit_0.digit_out[2] ));
 sg13g2_dfrbp_1 _2411_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net141),
    .D(_0216_),
    .Q_N(_1035_),
    .Q(\counter.counter_ref.digit_0.digit_out[3] ));
 sg13g2_dfrbp_1 _2412_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net134),
    .D(_0217_),
    .Q_N(_1034_),
    .Q(\counter.counter_ref.digits_out[4] ));
 sg13g2_dfrbp_1 _2413_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net128),
    .D(_0218_),
    .Q_N(_1033_),
    .Q(\counter.counter_ref.digits_out[5] ));
 sg13g2_dfrbp_1 _2414_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net122),
    .D(_0219_),
    .Q_N(_1032_),
    .Q(\counter.counter_ref.digits_out[6] ));
 sg13g2_dfrbp_1 _2415_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net110),
    .D(net192),
    .Q_N(_1031_),
    .Q(\counter.counter_ref.digits_out[7] ));
 sg13g2_dfrbp_1 _2416_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net104),
    .D(_0221_),
    .Q_N(_1030_),
    .Q(\counter.counter_ref.digits_out[8] ));
 sg13g2_dfrbp_1 _2417_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net98),
    .D(_0222_),
    .Q_N(_1029_),
    .Q(\counter.counter_ref.digits_out[9] ));
 sg13g2_dfrbp_1 _2418_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net92),
    .D(net203),
    .Q_N(_1028_),
    .Q(\counter.counter_ref.digits_out[10] ));
 sg13g2_dfrbp_1 _2419_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net80),
    .D(_0224_),
    .Q_N(_1027_),
    .Q(\counter.counter_ref.digits_out[11] ));
 sg13g2_dfrbp_1 _2420_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net64),
    .D(_0225_),
    .Q_N(_1026_),
    .Q(\counter.counter_ref.digits_out[12] ));
 sg13g2_dfrbp_1 _2421_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net50),
    .D(_0226_),
    .Q_N(_1025_),
    .Q(\counter.counter_ref.digits_out[13] ));
 sg13g2_dfrbp_1 _2422_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net17),
    .D(_0227_),
    .Q_N(_1024_),
    .Q(\counter.counter_ref.digits_out[14] ));
 sg13g2_dfrbp_1 _2423_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net145),
    .D(net290),
    .Q_N(_1023_),
    .Q(\counter.counter_ref.digits_out[15] ));
 sg13g2_dfrbp_1 _2424_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net131),
    .D(_0229_),
    .Q_N(_1022_),
    .Q(\counter.counter_ref.digits_out[16] ));
 sg13g2_dfrbp_1 _2425_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net113),
    .D(net330),
    .Q_N(_1021_),
    .Q(\counter.counter_ref.digits_out[17] ));
 sg13g2_dfrbp_1 _2426_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net101),
    .D(_0231_),
    .Q_N(_1020_),
    .Q(\counter.counter_ref.digits_out[18] ));
 sg13g2_dfrbp_1 _2427_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net83),
    .D(net383),
    .Q_N(_1019_),
    .Q(\counter.counter_ref.digits_out[19] ));
 sg13g2_dfrbp_1 _2428_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net57),
    .D(net316),
    .Q_N(_1018_),
    .Q(\counter.counter_ref.digits_out[20] ));
 sg13g2_dfrbp_1 _2429_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net153),
    .D(_0234_),
    .Q_N(_1017_),
    .Q(\counter.counter_ref.digits_out[21] ));
 sg13g2_dfrbp_1 _2430_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net125),
    .D(_0235_),
    .Q_N(_1016_),
    .Q(\counter.counter_ref.digits_out[22] ));
 sg13g2_dfrbp_1 _2431_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net159),
    .D(_0236_),
    .Q_N(_1146_),
    .Q(\counter.counter_ref.digits_out[23] ));
 sg13g2_dfrbp_1 _2432_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net160),
    .D(_0021_),
    .Q_N(_1147_),
    .Q(\counter.oled_driver.spi_driver.state_r[0] ));
 sg13g2_dfrbp_1 _2433_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net137),
    .D(net365),
    .Q_N(_1148_),
    .Q(\counter.oled_driver.spi_driver.state_r[1] ));
 sg13g2_dfrbp_1 _2434_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net95),
    .D(_0022_),
    .Q_N(_1015_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.start_in ));
 sg13g2_dfrbp_1 _2435_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net43),
    .D(_0237_),
    .Q_N(_1014_),
    .Q(\counter.refresh_display ));
 sg13g2_dfrbp_1 _2436_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net107),
    .D(_0238_),
    .Q_N(_0070_),
    .Q(\counter.streamer.graphical_decoder.pattern_adg[2] ));
 sg13g2_dfrbp_1 _2437_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net71),
    .D(_0239_),
    .Q_N(_0044_),
    .Q(\counter.streamer.graphical_decoder.pattern_adg[3] ));
 sg13g2_tiehi _2315__18 (.L_HI(net18));
 sg13g2_tiehi _2375__19 (.L_HI(net19));
 sg13g2_tiehi _2314__20 (.L_HI(net20));
 sg13g2_tiehi _2408__21 (.L_HI(net21));
 sg13g2_tiehi _2313__22 (.L_HI(net22));
 sg13g2_tiehi _2272__23 (.L_HI(net23));
 sg13g2_tiehi _2273__24 (.L_HI(net24));
 sg13g2_tiehi _2274__25 (.L_HI(net25));
 sg13g2_tiehi _2275__26 (.L_HI(net26));
 sg13g2_tiehi _2276__27 (.L_HI(net27));
 sg13g2_tiehi _2277__28 (.L_HI(net28));
 sg13g2_tiehi _2278__29 (.L_HI(net29));
 sg13g2_tiehi _2279__30 (.L_HI(net30));
 sg13g2_tiehi _2280__31 (.L_HI(net31));
 sg13g2_tiehi _2281__32 (.L_HI(net32));
 sg13g2_tiehi _2282__33 (.L_HI(net33));
 sg13g2_tiehi _2283__34 (.L_HI(net34));
 sg13g2_tiehi _2284__35 (.L_HI(net35));
 sg13g2_tiehi _2285__36 (.L_HI(net36));
 sg13g2_tiehi _2286__37 (.L_HI(net37));
 sg13g2_tiehi _2287__38 (.L_HI(net38));
 sg13g2_tiehi _2288__39 (.L_HI(net39));
 sg13g2_tiehi _2289__40 (.L_HI(net40));
 sg13g2_tiehi _2374__41 (.L_HI(net41));
 sg13g2_tiehi _2312__42 (.L_HI(net42));
 sg13g2_tiehi _2435__43 (.L_HI(net43));
 sg13g2_tiehi _2311__44 (.L_HI(net44));
 sg13g2_tiehi _2373__45 (.L_HI(net45));
 sg13g2_tiehi _2310__46 (.L_HI(net46));
 sg13g2_tiehi _2309__47 (.L_HI(net47));
 sg13g2_tiehi _2372__48 (.L_HI(net48));
 sg13g2_tiehi _2308__49 (.L_HI(net49));
 sg13g2_tiehi _2421__50 (.L_HI(net50));
 sg13g2_tiehi _2307__51 (.L_HI(net51));
 sg13g2_tiehi _2371__52 (.L_HI(net52));
 sg13g2_tiehi _2306__53 (.L_HI(net53));
 sg13g2_tiehi _2305__54 (.L_HI(net54));
 sg13g2_tiehi _2370__55 (.L_HI(net55));
 sg13g2_tiehi _2304__56 (.L_HI(net56));
 sg13g2_tiehi _2428__57 (.L_HI(net57));
 sg13g2_tiehi _2303__58 (.L_HI(net58));
 sg13g2_tiehi _2369__59 (.L_HI(net59));
 sg13g2_tiehi _2302__60 (.L_HI(net60));
 sg13g2_tiehi _2301__61 (.L_HI(net61));
 sg13g2_tiehi _2368__62 (.L_HI(net62));
 sg13g2_tiehi _2300__63 (.L_HI(net63));
 sg13g2_tiehi _2420__64 (.L_HI(net64));
 sg13g2_tiehi _2299__65 (.L_HI(net65));
 sg13g2_tiehi _2367__66 (.L_HI(net66));
 sg13g2_tiehi _2298__67 (.L_HI(net67));
 sg13g2_tiehi _2297__68 (.L_HI(net68));
 sg13g2_tiehi _2366__69 (.L_HI(net69));
 sg13g2_tiehi _2296__70 (.L_HI(net70));
 sg13g2_tiehi _2437__71 (.L_HI(net71));
 sg13g2_tiehi _2295__72 (.L_HI(net72));
 sg13g2_tiehi _2365__73 (.L_HI(net73));
 sg13g2_tiehi _2294__74 (.L_HI(net74));
 sg13g2_tiehi _2293__75 (.L_HI(net75));
 sg13g2_tiehi _2364__76 (.L_HI(net76));
 sg13g2_tiehi _2292__77 (.L_HI(net77));
 sg13g2_tiehi _2291__78 (.L_HI(net78));
 sg13g2_tiehi _2271__79 (.L_HI(net79));
 sg13g2_tiehi _2419__80 (.L_HI(net80));
 sg13g2_tiehi _2363__81 (.L_HI(net81));
 sg13g2_tiehi _2362__82 (.L_HI(net82));
 sg13g2_tiehi _2427__83 (.L_HI(net83));
 sg13g2_tiehi _2361__84 (.L_HI(net84));
 sg13g2_tiehi _2290__85 (.L_HI(net85));
 sg13g2_tiehi _2344__86 (.L_HI(net86));
 sg13g2_tiehi _2345__87 (.L_HI(net87));
 sg13g2_tiehi _2346__88 (.L_HI(net88));
 sg13g2_tiehi _2347__89 (.L_HI(net89));
 sg13g2_tiehi _2348__90 (.L_HI(net90));
 sg13g2_tiehi _2360__91 (.L_HI(net91));
 sg13g2_tiehi _2418__92 (.L_HI(net92));
 sg13g2_tiehi _2359__93 (.L_HI(net93));
 sg13g2_tiehi _2358__94 (.L_HI(net94));
 sg13g2_tiehi _2434__95 (.L_HI(net95));
 sg13g2_tiehi _2357__96 (.L_HI(net96));
 sg13g2_tiehi _2356__97 (.L_HI(net97));
 sg13g2_tiehi _2417__98 (.L_HI(net98));
 sg13g2_tiehi _2355__99 (.L_HI(net99));
 sg13g2_tiehi _2354__100 (.L_HI(net100));
 sg13g2_tiehi _2426__101 (.L_HI(net101));
 sg13g2_tiehi _2353__102 (.L_HI(net102));
 sg13g2_tiehi _2352__103 (.L_HI(net103));
 sg13g2_tiehi _2416__104 (.L_HI(net104));
 sg13g2_tiehi _2351__105 (.L_HI(net105));
 sg13g2_tiehi _2350__106 (.L_HI(net106));
 sg13g2_tiehi _2436__107 (.L_HI(net107));
 sg13g2_tiehi _2343__108 (.L_HI(net108));
 sg13g2_tiehi _2342__109 (.L_HI(net109));
 sg13g2_tiehi _2415__110 (.L_HI(net110));
 sg13g2_tiehi _2341__111 (.L_HI(net111));
 sg13g2_tiehi _2340__112 (.L_HI(net112));
 sg13g2_tiehi _2425__113 (.L_HI(net113));
 sg13g2_tiehi _2349__114 (.L_HI(net114));
 sg13g2_tiehi _2381__115 (.L_HI(net115));
 sg13g2_tiehi _2382__116 (.L_HI(net116));
 sg13g2_tiehi _2383__117 (.L_HI(net117));
 sg13g2_tiehi _2384__118 (.L_HI(net118));
 sg13g2_tiehi _2385__119 (.L_HI(net119));
 sg13g2_tiehi _2339__120 (.L_HI(net120));
 sg13g2_tiehi _2338__121 (.L_HI(net121));
 sg13g2_tiehi _2414__122 (.L_HI(net122));
 sg13g2_tiehi _2337__123 (.L_HI(net123));
 sg13g2_tiehi _2336__124 (.L_HI(net124));
 sg13g2_tiehi _2430__125 (.L_HI(net125));
 sg13g2_tiehi _2335__126 (.L_HI(net126));
 sg13g2_tiehi _2334__127 (.L_HI(net127));
 sg13g2_tiehi _2413__128 (.L_HI(net128));
 sg13g2_tiehi _2333__129 (.L_HI(net129));
 sg13g2_tiehi _2332__130 (.L_HI(net130));
 sg13g2_tiehi _2424__131 (.L_HI(net131));
 sg13g2_tiehi _2331__132 (.L_HI(net132));
 sg13g2_tiehi _2330__133 (.L_HI(net133));
 sg13g2_tiehi _2412__134 (.L_HI(net134));
 sg13g2_tiehi _2329__135 (.L_HI(net135));
 sg13g2_tiehi _2328__136 (.L_HI(net136));
 sg13g2_tiehi _2433__137 (.L_HI(net137));
 sg13g2_tiehi _2327__138 (.L_HI(net138));
 sg13g2_tiehi _2387__139 (.L_HI(net139));
 sg13g2_tiehi _2326__140 (.L_HI(net140));
 sg13g2_tiehi _2411__141 (.L_HI(net141));
 sg13g2_tiehi _2325__142 (.L_HI(net142));
 sg13g2_tiehi _2380__143 (.L_HI(net143));
 sg13g2_tiehi _2324__144 (.L_HI(net144));
 sg13g2_tiehi _2423__145 (.L_HI(net145));
 sg13g2_tiehi _2323__146 (.L_HI(net146));
 sg13g2_tiehi _2379__147 (.L_HI(net147));
 sg13g2_tiehi _2322__148 (.L_HI(net148));
 sg13g2_tiehi _2410__149 (.L_HI(net149));
 sg13g2_tiehi _2321__150 (.L_HI(net150));
 sg13g2_tiehi _2378__151 (.L_HI(net151));
 sg13g2_tiehi _2320__152 (.L_HI(net152));
 sg13g2_tiehi _2429__153 (.L_HI(net153));
 sg13g2_tiehi _2319__154 (.L_HI(net154));
 sg13g2_tiehi _2377__155 (.L_HI(net155));
 sg13g2_tiehi _2318__156 (.L_HI(net156));
 sg13g2_tiehi _2409__157 (.L_HI(net157));
 sg13g2_tiehi _2386__158 (.L_HI(net158));
 sg13g2_tiehi _2431__159 (.L_HI(net159));
 sg13g2_tiehi _2432__160 (.L_HI(net160));
 sg13g2_tiehi _2317__161 (.L_HI(net161));
 sg13g2_tiehi _2376__162 (.L_HI(net162));
 sg13g2_tiehi _2316__163 (.L_HI(net163));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_tielo tt_um_frequency_counter_2 (.L_LO(net2));
 sg13g2_tielo tt_um_frequency_counter_3 (.L_LO(net3));
 sg13g2_tielo tt_um_frequency_counter_4 (.L_LO(net4));
 sg13g2_tielo tt_um_frequency_counter_5 (.L_LO(net5));
 sg13g2_tielo tt_um_frequency_counter_6 (.L_LO(net6));
 sg13g2_tielo tt_um_frequency_counter_7 (.L_LO(net7));
 sg13g2_tielo tt_um_frequency_counter_8 (.L_LO(net8));
 sg13g2_tielo tt_um_frequency_counter_9 (.L_LO(net9));
 sg13g2_tielo tt_um_frequency_counter_10 (.L_LO(net10));
 sg13g2_tielo tt_um_frequency_counter_11 (.L_LO(net11));
 sg13g2_tielo tt_um_frequency_counter_12 (.L_LO(net12));
 sg13g2_tielo tt_um_frequency_counter_13 (.L_LO(net13));
 sg13g2_tielo tt_um_frequency_counter_14 (.L_LO(net14));
 sg13g2_tielo tt_um_frequency_counter_15 (.L_LO(net15));
 sg13g2_tielo tt_um_frequency_counter_16 (.L_LO(net16));
 sg13g2_tiehi _2422__17 (.L_HI(net17));
 sg13g2_buf_2 _2601_ (.A(\counter.oled_driver.mc_exec.oled_rstn_out ),
    .X(uo_out[0]));
 sg13g2_buf_1 _2602_ (.A(\counter.oled_driver.mc_exec.oled_vbatn_out ),
    .X(uo_out[1]));
 sg13g2_buf_1 _2603_ (.A(\counter.oled_driver.mc_exec.oled_vcdn_out ),
    .X(uo_out[2]));
 sg13g2_buf_1 _2604_ (.A(\counter.oled_csn_out ),
    .X(uo_out[3]));
 sg13g2_buf_1 _2605_ (.A(\counter.oled_dc_out ),
    .X(uo_out[4]));
 sg13g2_buf_1 _2606_ (.A(\counter.oled_clk_out ),
    .X(uo_out[5]));
 sg13g2_buf_1 _2607_ (.A(\counter.oled_driver.oled_mosi_out ),
    .X(uo_out[6]));
 sg13g2_buf_1 _2608_ (.A(ui_in[7]),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout213 (.A(_0833_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_0792_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_0791_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_0168_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_0408_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_0799_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_0790_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_0768_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_0759_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_1011_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_0947_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_0914_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_0730_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_0725_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(net228),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_0079_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(net230),
    .X(net229));
 sg13g2_buf_4 fanout230 (.X(net230),
    .A(_0633_));
 sg13g2_buf_2 fanout231 (.A(net233),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(net233),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(net235),
    .X(net233));
 sg13g2_buf_1 fanout234 (.A(net235),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_0746_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(net238),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(net238),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_0746_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(net240),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(net242),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(net242),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_0699_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(net244),
    .X(net243));
 sg13g2_buf_4 fanout244 (.X(net244),
    .A(_0699_));
 sg13g2_buf_4 fanout245 (.X(net245),
    .A(\counter.oled_driver.mc_exec.microcode_rom.address[5] ));
 sg13g2_buf_2 fanout246 (.A(net247),
    .X(net246));
 sg13g2_buf_1 fanout247 (.A(\counter.streamer.graphical_decoder.index_y_in[1] ),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(\counter.streamer.graphical_decoder.index_x_in[1] ),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(net250),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(\counter.streamer.digit_cnt_r[1] ),
    .X(net250));
 sg13g2_buf_4 fanout251 (.X(net251),
    .A(net252));
 sg13g2_buf_4 fanout252 (.X(net252),
    .A(\counter.streamer.digit_cnt_r[0] ));
 sg13g2_buf_2 fanout253 (.A(net255),
    .X(net253));
 sg13g2_buf_1 fanout254 (.A(net255),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(net256),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(net257),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(net411),
    .X(net257));
 sg13g2_buf_4 fanout258 (.X(net258),
    .A(\counter.oled_driver.mc_exec.state_r[2] ));
 sg13g2_buf_2 fanout259 (.A(\counter.cnt_ref_enable ),
    .X(net259));
 sg13g2_buf_1 fanout260 (.A(\counter.cnt_ref_enable ),
    .X(net260));
 sg13g2_buf_4 fanout261 (.X(net261),
    .A(net265));
 sg13g2_buf_2 fanout262 (.A(net263),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(net264),
    .X(net263));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(net265));
 sg13g2_buf_2 fanout265 (.A(\counter.oled_driver.mc_exec.reset_in ),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(net267),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(ui_in[0]),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(ui_in[0]),
    .X(net268));
 sg13g2_buf_1 fanout269 (.A(ui_in[0]),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(net271),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(net276),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(net273),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(net275),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(net275),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(net276),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(rst_n),
    .X(net276));
 sg13g2_buf_4 fanout277 (.X(net277),
    .A(net278));
 sg13g2_buf_2 fanout278 (.A(net280),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(net280),
    .X(net279));
 sg13g2_buf_4 fanout280 (.X(net280),
    .A(rst_n));
 sg13g2_tielo tt_um_frequency_counter_1 (.L_LO(net1));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_buf_2 clkbuf_5_0__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_1__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_2__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_2__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_3__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_4__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_4__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_5__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_6__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_6__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_7__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_8__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_8__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_9__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_10__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_10__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_11__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_12__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_12__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_13__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_14__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_14__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_15__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_15__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_16__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_16__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_17__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_18__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_18__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_19__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_20__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_20__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_21__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_22__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_22__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_23__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_23__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_24__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_24__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_25__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_26__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_26__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_27__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_28__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_28__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_29__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_29__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_30__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_30__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_31__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_31__leaf_clk_regs));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk_regs));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk_regs));
 sg13g2_inv_1 clkload3 (.A(clknet_5_11__leaf_clk_regs));
 sg13g2_inv_1 clkload4 (.A(clknet_5_13__leaf_clk_regs));
 sg13g2_inv_1 clkload5 (.A(clknet_5_15__leaf_clk_regs));
 sg13g2_inv_1 clkload6 (.A(clknet_5_19__leaf_clk_regs));
 sg13g2_inv_1 clkload7 (.A(clknet_5_21__leaf_clk_regs));
 sg13g2_inv_1 clkload8 (.A(clknet_5_23__leaf_clk_regs));
 sg13g2_inv_1 clkload9 (.A(clknet_5_25__leaf_clk_regs));
 sg13g2_inv_1 clkload10 (.A(clknet_5_27__leaf_clk_regs));
 sg13g2_inv_1 clkload11 (.A(clknet_5_29__leaf_clk_regs));
 sg13g2_inv_1 clkload12 (.A(clknet_5_31__leaf_clk_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0078_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0187_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0059_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0027_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold5 (.A(\counter.counter_ref.digits_out[4] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold6 (.A(\counter.oled_driver.spi_data[4] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold7 (.A(\counter.oled_driver.spi_data[7] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0158_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold9 (.A(\counter.oled_driver.spi_data[2] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0153_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold11 (.A(\counter.oled_driver.mc_exec.delay_cnt[10] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0179_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold13 (.A(\counter.oled_driver.mc_exec.delay_cnt[6] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0175_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold15 (.A(\counter.oled_driver.spi_data[3] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold16 (.A(\counter.state[0] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0742_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0029_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0068_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0117_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold21 (.A(\counter.streamer.state_r[4] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0014_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold23 (.A(\counter.state[1] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0693_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0028_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold26 (.A(\counter.oled_driver.mc_exec.delay_cnt[4] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0173_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold28 (.A(\counter.counter_ref.digits_out[7] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0220_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold30 (.A(\counter.oled_driver.spi_driver.deactivate_cs_r ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0468_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0192_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold33 (.A(\counter.oled_driver.spi_data[1] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0339_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold35 (.A(\counter.oled_driver.mc_exec.state_r[5] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0906_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0010_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold38 (.A(\counter.counter_ref.digits_out[10] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0489_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0223_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold41 (.A(\counter.oled_driver.mc_exec.delay_cnt[13] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0182_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold43 (.A(\counter.oled_driver.mc_exec.spi_tx_trigger_out ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0687_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0016_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold46 (.A(\counter.counter_ref.digit_0.digit_out[1] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0473_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0214_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold49 (.A(\counter.oled_driver.spi_data[6] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0378_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold51 (.A(\counter.counter_ref.digits_out[18] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0512_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold53 (.A(\counter.oled_driver.mc_exec.delay_cnt[2] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0171_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold55 (.A(\counter.oled_driver.spi_data[5] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0156_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold57 (.A(\counter.counter_ref.digits_out[15] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0502_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0228_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold60 (.A(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[0] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0186_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold62 (.A(\counter.oled_driver.mc_exec.procedure_offset_in[0] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0970_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0116_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold65 (.A(\counter.oled_driver.state_r[4] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0013_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold67 (.A(\counter.oled_driver.spi_data[0] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0324_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0046_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0951_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0110_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold72 (.A(\counter.counter_ref.digits_out[5] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0479_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold74 (.A(\counter.streamer.digits_r[19] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0055_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0684_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0018_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold78 (.A(\counter.oled_driver.oled_mosi_out ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0966_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0115_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold81 (.A(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[1] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0188_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold83 (.A(\counter.counter_ref.digits_out[20] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0517_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0233_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold86 (.A(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[5] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0959_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0113_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold89 (.A(\counter.oled_driver.mc_exec.state_r[0] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0032_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold91 (.A(\counter.streamer.digits_r[15] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold92 (.A(\counter.counter_ref.digits_out[22] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0521_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold94 (.A(\counter.counter_ref.digits_out[21] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0519_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold96 (.A(\counter.streamer.digits_r[3] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold97 (.A(\counter.counter_ref.digits_out[17] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0508_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0230_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold100 (.A(\counter.counter_ref.digit_0.digit_out[3] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0476_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0047_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0957_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0112_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold105 (.A(\counter.oled_driver.mc_exec.oled_vcdn_out ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0385_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0159_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold108 (.A(\counter.oled_driver.mc_exec.delay_cnt[16] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0455_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0185_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold111 (.A(\counter.streamer.digits_r[7] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold112 (.A(\counter.oled_driver.mc_exec.delay_cnt[3] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0420_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0172_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold115 (.A(\counter.oled_driver.mc_exec.microcode_rom.address[2] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold116 (.A(\counter.oled_driver.spi_driver.state_r[1] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0191_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold118 (.A(\counter.streamer.digits_r[9] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold119 (.A(\counter.oled_driver.mc_exec.delay_cnt[11] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0439_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold121 (.A(\counter.streamer.digits_r[16] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold122 (.A(\counter.counter_ref.digits_out[8] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold123 (.A(\counter.oled_driver.sync_stb_in ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0030_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold125 (.A(\counter.streamer.digits_r[18] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold126 (.A(\counter.oled_driver.mc_exec.procedure_start_in ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0025_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold128 (.A(\counter.counter_ref.digits_out[9] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold129 (.A(\counter.oled_driver.write_stb_in ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0024_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold131 (.A(\counter.streamer.digits_r[12] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold132 (.A(\counter.streamer.digits_r[11] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold133 (.A(\counter.oled_driver.spi_driver.shift_reg.start_in ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0011_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold135 (.A(\counter.streamer.digits_r[0] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold136 (.A(\counter.oled_driver.mc_exec.delay_cnt[9] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0432_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold138 (.A(\counter.oled_driver.mc_exec.delay_cnt[1] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0415_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0170_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold141 (.A(\counter.oled_driver.mc_exec.state_r[6] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0749_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold143 (.A(\counter.streamer.digits_r[17] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold144 (.A(\counter.counter_ref.digits_out[23] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold145 (.A(\counter.refresh_display ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold146 (.A(\counter.counter_ref.digit_0.digit_out[2] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0474_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0054_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0663_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0023_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold151 (.A(\counter.counter_ref.digits_out[19] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0232_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold153 (.A(\counter.oled_driver.mc_exec.oled_dc_out ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0399_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0162_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold156 (.A(\counter.streamer.digits_r[20] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold157 (.A(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[3] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0724_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold159 (.A(\counter.counter_ref.digits_out[12] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold160 (.A(\counter.oled_driver.mc_exec.delay_cnt[14] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0449_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0183_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold163 (.A(\counter.oled_driver.mc_exec.oled_vbatn_out ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0390_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0160_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold166 (.A(\counter.oled_driver.state_r[2] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0012_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold168 (.A(\counter.oled_driver.mc_exec.microcode_rom.address[3] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0166_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold170 (.A(\counter.streamer.state_r[5] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0015_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold172 (.A(\counter.oled_driver.mc_exec.oled_rstn_out ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0161_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold174 (.A(\counter.streamer.digits_r[14] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold175 (.A(\counter.streamer.digits_r[23] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold176 (.A(\counter.streamer.digits_r[5] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold177 (.A(\counter.counter_ref.digit_0.digit_out[0] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0470_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold179 (.A(\counter.streamer.digits_r[13] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold180 (.A(\counter.oled_driver.mc_exec.procedure_done_out ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold181 (.A(\counter.streamer.digits_r[22] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold182 (.A(\counter.oled_driver.mc_exec.microcode_rom.address[1] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0164_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold184 (.A(\counter.streamer.digits_r[1] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold185 (.A(\counter.oled_driver.mc_exec.delay_cnt[5] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0424_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold187 (.A(\counter.streamer.digits_r[4] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold188 (.A(\counter.streamer.digits_r[8] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold189 (.A(\counter.streamer.digits_r[21] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold190 (.A(\counter.streamer.digits_r[2] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold191 (.A(\counter.counter_ref.digits_out[6] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold192 (.A(\counter.oled_driver.mc_exec.delay_cnt[7] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0428_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold194 (.A(\counter.counter_ref.digits_out[11] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold195 (.A(\counter.streamer.digits_r[10] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold196 (.A(\counter.oled_driver.mc_exec.delay_cnt[12] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0443_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0181_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold199 (.A(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[6] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold200 (.A(\counter.streamer.graphical_decoder.index_x_in[4] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold201 (.A(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[2] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0461_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold203 (.A(\counter.oled_driver.mc_exec.microcode_rom.address[0] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold204 (.A(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[3] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0955_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold206 (.A(\counter.oled_driver.mc_exec.delay_cnt[0] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0069_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold208 (.A(\counter.counter_ref.digits_out[14] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold209 (.A(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[1] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold210 (.A(\counter.oled_driver.mc_exec.state_r[3] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0653_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0019_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold213 (.A(\counter.oled_driver.mc_exec.delay_cnt[15] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0451_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0184_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold216 (.A(\counter.streamer.digits_r[6] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold217 (.A(\counter.counter_ref.digits_out[13] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold218 (.A(\counter.oled_driver.spi_driver.state_r[0] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0017_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold220 (.A(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[0] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold221 (.A(\counter.oled_driver.mc_exec.delay_cnt[8] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0067_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0119_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold224 (.A(\counter.streamer.graphical_decoder.index_x_in[3] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0925_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold226 (.A(\counter.counter_ref.digits_out[16] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold227 (.A(\counter.streamer.graphical_decoder.index_x_in[2] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold228 (.A(\counter.streamer.graphical_decoder.index_y_in[0] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0983_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0065_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0124_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold232 (.A(\counter.streamer.graphical_decoder.index_x_in[0] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold233 (.A(\counter.counter_ref.digit_0.digit_out[1] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0701_),
    .X(net465));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_4 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_295 ();
 sg13g2_decap_8 FILLER_14_302 ();
 sg13g2_decap_8 FILLER_14_309 ();
 sg13g2_decap_8 FILLER_14_316 ();
 sg13g2_decap_8 FILLER_14_323 ();
 sg13g2_decap_8 FILLER_14_330 ();
 sg13g2_decap_8 FILLER_14_337 ();
 sg13g2_decap_8 FILLER_14_344 ();
 sg13g2_decap_8 FILLER_14_351 ();
 sg13g2_decap_8 FILLER_14_358 ();
 sg13g2_decap_8 FILLER_14_365 ();
 sg13g2_decap_8 FILLER_14_372 ();
 sg13g2_decap_8 FILLER_14_379 ();
 sg13g2_decap_8 FILLER_14_386 ();
 sg13g2_decap_8 FILLER_14_393 ();
 sg13g2_decap_8 FILLER_14_400 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_fill_2 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_311 ();
 sg13g2_decap_8 FILLER_15_318 ();
 sg13g2_decap_8 FILLER_15_325 ();
 sg13g2_decap_8 FILLER_15_332 ();
 sg13g2_decap_8 FILLER_15_339 ();
 sg13g2_decap_8 FILLER_15_346 ();
 sg13g2_decap_8 FILLER_15_353 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_decap_8 FILLER_15_367 ();
 sg13g2_decap_8 FILLER_15_374 ();
 sg13g2_decap_8 FILLER_15_381 ();
 sg13g2_decap_8 FILLER_15_388 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_4 FILLER_16_266 ();
 sg13g2_fill_2 FILLER_16_270 ();
 sg13g2_fill_1 FILLER_16_307 ();
 sg13g2_decap_8 FILLER_16_334 ();
 sg13g2_decap_8 FILLER_16_341 ();
 sg13g2_decap_8 FILLER_16_348 ();
 sg13g2_decap_8 FILLER_16_355 ();
 sg13g2_decap_8 FILLER_16_362 ();
 sg13g2_decap_8 FILLER_16_369 ();
 sg13g2_decap_8 FILLER_16_376 ();
 sg13g2_decap_8 FILLER_16_383 ();
 sg13g2_decap_8 FILLER_16_390 ();
 sg13g2_decap_8 FILLER_16_397 ();
 sg13g2_decap_4 FILLER_16_404 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_fill_1 FILLER_17_266 ();
 sg13g2_fill_1 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_341 ();
 sg13g2_decap_8 FILLER_17_348 ();
 sg13g2_decap_8 FILLER_17_355 ();
 sg13g2_decap_8 FILLER_17_362 ();
 sg13g2_decap_8 FILLER_17_369 ();
 sg13g2_decap_8 FILLER_17_376 ();
 sg13g2_decap_8 FILLER_17_383 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_4 FILLER_18_245 ();
 sg13g2_fill_1 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_334 ();
 sg13g2_decap_8 FILLER_18_341 ();
 sg13g2_decap_8 FILLER_18_348 ();
 sg13g2_decap_8 FILLER_18_355 ();
 sg13g2_decap_8 FILLER_18_362 ();
 sg13g2_decap_8 FILLER_18_369 ();
 sg13g2_decap_8 FILLER_18_376 ();
 sg13g2_decap_8 FILLER_18_383 ();
 sg13g2_decap_8 FILLER_18_390 ();
 sg13g2_decap_8 FILLER_18_397 ();
 sg13g2_decap_4 FILLER_18_404 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_fill_2 FILLER_19_285 ();
 sg13g2_fill_1 FILLER_19_287 ();
 sg13g2_fill_1 FILLER_19_307 ();
 sg13g2_decap_8 FILLER_19_339 ();
 sg13g2_decap_8 FILLER_19_346 ();
 sg13g2_decap_8 FILLER_19_353 ();
 sg13g2_decap_8 FILLER_19_360 ();
 sg13g2_decap_8 FILLER_19_367 ();
 sg13g2_decap_8 FILLER_19_374 ();
 sg13g2_decap_8 FILLER_19_381 ();
 sg13g2_decap_8 FILLER_19_388 ();
 sg13g2_decap_8 FILLER_19_395 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_fill_1 FILLER_20_238 ();
 sg13g2_fill_1 FILLER_20_243 ();
 sg13g2_fill_2 FILLER_20_300 ();
 sg13g2_fill_1 FILLER_20_302 ();
 sg13g2_fill_2 FILLER_20_308 ();
 sg13g2_fill_1 FILLER_20_310 ();
 sg13g2_decap_8 FILLER_20_334 ();
 sg13g2_decap_8 FILLER_20_341 ();
 sg13g2_decap_8 FILLER_20_348 ();
 sg13g2_decap_8 FILLER_20_355 ();
 sg13g2_decap_8 FILLER_20_362 ();
 sg13g2_decap_8 FILLER_20_369 ();
 sg13g2_decap_8 FILLER_20_376 ();
 sg13g2_decap_8 FILLER_20_383 ();
 sg13g2_decap_8 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_397 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_4 FILLER_21_224 ();
 sg13g2_fill_1 FILLER_21_262 ();
 sg13g2_fill_2 FILLER_21_277 ();
 sg13g2_decap_8 FILLER_21_339 ();
 sg13g2_decap_8 FILLER_21_346 ();
 sg13g2_decap_8 FILLER_21_353 ();
 sg13g2_decap_8 FILLER_21_360 ();
 sg13g2_decap_8 FILLER_21_367 ();
 sg13g2_decap_8 FILLER_21_374 ();
 sg13g2_decap_8 FILLER_21_381 ();
 sg13g2_decap_8 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_fill_2 FILLER_22_224 ();
 sg13g2_fill_1 FILLER_22_296 ();
 sg13g2_fill_1 FILLER_22_312 ();
 sg13g2_decap_8 FILLER_22_348 ();
 sg13g2_decap_8 FILLER_22_355 ();
 sg13g2_decap_8 FILLER_22_362 ();
 sg13g2_decap_8 FILLER_22_369 ();
 sg13g2_decap_8 FILLER_22_376 ();
 sg13g2_decap_8 FILLER_22_383 ();
 sg13g2_decap_8 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_4 FILLER_23_168 ();
 sg13g2_fill_1 FILLER_23_176 ();
 sg13g2_decap_8 FILLER_23_185 ();
 sg13g2_decap_8 FILLER_23_192 ();
 sg13g2_decap_8 FILLER_23_199 ();
 sg13g2_decap_8 FILLER_23_206 ();
 sg13g2_decap_8 FILLER_23_213 ();
 sg13g2_fill_2 FILLER_23_220 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_4 FILLER_24_154 ();
 sg13g2_fill_2 FILLER_24_158 ();
 sg13g2_decap_4 FILLER_24_164 ();
 sg13g2_decap_8 FILLER_24_194 ();
 sg13g2_decap_8 FILLER_24_201 ();
 sg13g2_decap_8 FILLER_24_208 ();
 sg13g2_decap_4 FILLER_24_215 ();
 sg13g2_fill_2 FILLER_24_219 ();
 sg13g2_fill_1 FILLER_24_247 ();
 sg13g2_fill_1 FILLER_24_284 ();
 sg13g2_fill_2 FILLER_24_297 ();
 sg13g2_decap_8 FILLER_24_334 ();
 sg13g2_decap_8 FILLER_24_341 ();
 sg13g2_decap_8 FILLER_24_348 ();
 sg13g2_decap_8 FILLER_24_355 ();
 sg13g2_decap_8 FILLER_24_362 ();
 sg13g2_decap_8 FILLER_24_369 ();
 sg13g2_decap_8 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_24_383 ();
 sg13g2_decap_8 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_4 FILLER_25_147 ();
 sg13g2_fill_2 FILLER_25_164 ();
 sg13g2_fill_2 FILLER_25_176 ();
 sg13g2_fill_1 FILLER_25_187 ();
 sg13g2_decap_8 FILLER_25_205 ();
 sg13g2_decap_8 FILLER_25_212 ();
 sg13g2_decap_8 FILLER_25_219 ();
 sg13g2_decap_8 FILLER_25_226 ();
 sg13g2_fill_1 FILLER_25_240 ();
 sg13g2_fill_2 FILLER_25_263 ();
 sg13g2_fill_2 FILLER_25_304 ();
 sg13g2_decap_8 FILLER_25_320 ();
 sg13g2_decap_8 FILLER_25_327 ();
 sg13g2_decap_8 FILLER_25_334 ();
 sg13g2_decap_8 FILLER_25_341 ();
 sg13g2_decap_8 FILLER_25_348 ();
 sg13g2_decap_8 FILLER_25_355 ();
 sg13g2_decap_8 FILLER_25_362 ();
 sg13g2_decap_8 FILLER_25_369 ();
 sg13g2_decap_8 FILLER_25_376 ();
 sg13g2_decap_8 FILLER_25_383 ();
 sg13g2_decap_8 FILLER_25_390 ();
 sg13g2_decap_8 FILLER_25_397 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_4 FILLER_26_140 ();
 sg13g2_fill_2 FILLER_26_144 ();
 sg13g2_fill_2 FILLER_26_172 ();
 sg13g2_fill_1 FILLER_26_183 ();
 sg13g2_decap_8 FILLER_26_206 ();
 sg13g2_decap_8 FILLER_26_213 ();
 sg13g2_decap_4 FILLER_26_220 ();
 sg13g2_fill_2 FILLER_26_224 ();
 sg13g2_decap_4 FILLER_26_265 ();
 sg13g2_fill_2 FILLER_26_269 ();
 sg13g2_fill_2 FILLER_26_279 ();
 sg13g2_fill_1 FILLER_26_281 ();
 sg13g2_fill_2 FILLER_26_300 ();
 sg13g2_decap_8 FILLER_26_334 ();
 sg13g2_decap_8 FILLER_26_341 ();
 sg13g2_decap_8 FILLER_26_348 ();
 sg13g2_decap_8 FILLER_26_355 ();
 sg13g2_decap_8 FILLER_26_362 ();
 sg13g2_decap_8 FILLER_26_369 ();
 sg13g2_decap_8 FILLER_26_376 ();
 sg13g2_decap_8 FILLER_26_383 ();
 sg13g2_decap_8 FILLER_26_390 ();
 sg13g2_decap_8 FILLER_26_397 ();
 sg13g2_decap_4 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_fill_2 FILLER_27_166 ();
 sg13g2_fill_1 FILLER_27_199 ();
 sg13g2_decap_8 FILLER_27_212 ();
 sg13g2_decap_8 FILLER_27_219 ();
 sg13g2_decap_8 FILLER_27_226 ();
 sg13g2_fill_2 FILLER_27_233 ();
 sg13g2_fill_1 FILLER_27_235 ();
 sg13g2_decap_8 FILLER_27_240 ();
 sg13g2_decap_4 FILLER_27_247 ();
 sg13g2_fill_2 FILLER_27_251 ();
 sg13g2_decap_8 FILLER_27_257 ();
 sg13g2_decap_8 FILLER_27_264 ();
 sg13g2_fill_2 FILLER_27_298 ();
 sg13g2_decap_8 FILLER_27_344 ();
 sg13g2_decap_8 FILLER_27_351 ();
 sg13g2_decap_8 FILLER_27_358 ();
 sg13g2_decap_8 FILLER_27_365 ();
 sg13g2_decap_8 FILLER_27_372 ();
 sg13g2_decap_8 FILLER_27_379 ();
 sg13g2_decap_8 FILLER_27_386 ();
 sg13g2_decap_8 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_4 FILLER_28_140 ();
 sg13g2_fill_2 FILLER_28_144 ();
 sg13g2_fill_1 FILLER_28_180 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_4 FILLER_28_231 ();
 sg13g2_fill_1 FILLER_28_235 ();
 sg13g2_fill_2 FILLER_28_240 ();
 sg13g2_fill_1 FILLER_28_242 ();
 sg13g2_fill_2 FILLER_28_247 ();
 sg13g2_fill_2 FILLER_28_258 ();
 sg13g2_fill_1 FILLER_28_260 ();
 sg13g2_fill_2 FILLER_28_303 ();
 sg13g2_decap_8 FILLER_28_335 ();
 sg13g2_decap_8 FILLER_28_342 ();
 sg13g2_decap_8 FILLER_28_349 ();
 sg13g2_decap_8 FILLER_28_356 ();
 sg13g2_decap_8 FILLER_28_363 ();
 sg13g2_decap_8 FILLER_28_370 ();
 sg13g2_decap_8 FILLER_28_377 ();
 sg13g2_decap_8 FILLER_28_384 ();
 sg13g2_decap_8 FILLER_28_391 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_fill_1 FILLER_29_154 ();
 sg13g2_fill_2 FILLER_29_167 ();
 sg13g2_fill_1 FILLER_29_169 ();
 sg13g2_decap_8 FILLER_29_194 ();
 sg13g2_decap_8 FILLER_29_201 ();
 sg13g2_decap_8 FILLER_29_208 ();
 sg13g2_decap_8 FILLER_29_215 ();
 sg13g2_fill_2 FILLER_29_222 ();
 sg13g2_fill_1 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_324 ();
 sg13g2_decap_8 FILLER_29_331 ();
 sg13g2_decap_8 FILLER_29_342 ();
 sg13g2_decap_8 FILLER_29_349 ();
 sg13g2_decap_8 FILLER_29_356 ();
 sg13g2_decap_8 FILLER_29_363 ();
 sg13g2_decap_8 FILLER_29_370 ();
 sg13g2_decap_8 FILLER_29_377 ();
 sg13g2_decap_8 FILLER_29_384 ();
 sg13g2_decap_8 FILLER_29_391 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_fill_2 FILLER_30_154 ();
 sg13g2_fill_1 FILLER_30_170 ();
 sg13g2_fill_2 FILLER_30_179 ();
 sg13g2_fill_1 FILLER_30_181 ();
 sg13g2_fill_1 FILLER_30_194 ();
 sg13g2_decap_8 FILLER_30_213 ();
 sg13g2_fill_1 FILLER_30_220 ();
 sg13g2_decap_4 FILLER_30_314 ();
 sg13g2_fill_1 FILLER_30_326 ();
 sg13g2_decap_4 FILLER_30_353 ();
 sg13g2_fill_2 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_362 ();
 sg13g2_decap_8 FILLER_30_369 ();
 sg13g2_decap_8 FILLER_30_376 ();
 sg13g2_decap_8 FILLER_30_383 ();
 sg13g2_decap_8 FILLER_30_390 ();
 sg13g2_decap_8 FILLER_30_397 ();
 sg13g2_decap_4 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_fill_1 FILLER_31_140 ();
 sg13g2_fill_1 FILLER_31_185 ();
 sg13g2_decap_8 FILLER_31_212 ();
 sg13g2_decap_4 FILLER_31_219 ();
 sg13g2_fill_1 FILLER_31_223 ();
 sg13g2_fill_2 FILLER_31_250 ();
 sg13g2_fill_2 FILLER_31_279 ();
 sg13g2_fill_1 FILLER_31_281 ();
 sg13g2_fill_2 FILLER_31_336 ();
 sg13g2_fill_1 FILLER_31_338 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_4 FILLER_32_133 ();
 sg13g2_fill_1 FILLER_32_163 ();
 sg13g2_decap_8 FILLER_32_208 ();
 sg13g2_decap_8 FILLER_32_215 ();
 sg13g2_decap_8 FILLER_32_222 ();
 sg13g2_fill_2 FILLER_32_229 ();
 sg13g2_fill_2 FILLER_32_276 ();
 sg13g2_fill_1 FILLER_32_278 ();
 sg13g2_fill_1 FILLER_32_328 ();
 sg13g2_fill_1 FILLER_32_337 ();
 sg13g2_decap_8 FILLER_32_381 ();
 sg13g2_decap_8 FILLER_32_388 ();
 sg13g2_decap_8 FILLER_32_395 ();
 sg13g2_decap_8 FILLER_32_402 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_fill_2 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_212 ();
 sg13g2_decap_8 FILLER_33_219 ();
 sg13g2_decap_8 FILLER_33_226 ();
 sg13g2_fill_1 FILLER_33_233 ();
 sg13g2_fill_2 FILLER_33_267 ();
 sg13g2_fill_1 FILLER_33_269 ();
 sg13g2_fill_2 FILLER_33_302 ();
 sg13g2_fill_1 FILLER_33_304 ();
 sg13g2_fill_1 FILLER_33_321 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_4 FILLER_34_133 ();
 sg13g2_fill_2 FILLER_34_137 ();
 sg13g2_fill_1 FILLER_34_192 ();
 sg13g2_decap_8 FILLER_34_201 ();
 sg13g2_decap_8 FILLER_34_208 ();
 sg13g2_decap_8 FILLER_34_215 ();
 sg13g2_decap_8 FILLER_34_222 ();
 sg13g2_decap_8 FILLER_34_229 ();
 sg13g2_fill_2 FILLER_34_236 ();
 sg13g2_fill_1 FILLER_34_324 ();
 sg13g2_fill_1 FILLER_34_335 ();
 sg13g2_decap_8 FILLER_34_377 ();
 sg13g2_decap_8 FILLER_34_384 ();
 sg13g2_decap_8 FILLER_34_391 ();
 sg13g2_decap_8 FILLER_34_398 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_fill_2 FILLER_35_159 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_decap_4 FILLER_35_245 ();
 sg13g2_decap_4 FILLER_35_253 ();
 sg13g2_fill_1 FILLER_35_257 ();
 sg13g2_fill_1 FILLER_35_349 ();
 sg13g2_decap_8 FILLER_35_383 ();
 sg13g2_decap_8 FILLER_35_390 ();
 sg13g2_decap_8 FILLER_35_397 ();
 sg13g2_decap_4 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_fill_1 FILLER_36_147 ();
 sg13g2_fill_2 FILLER_36_174 ();
 sg13g2_fill_1 FILLER_36_197 ();
 sg13g2_fill_1 FILLER_36_207 ();
 sg13g2_decap_8 FILLER_36_213 ();
 sg13g2_decap_8 FILLER_36_220 ();
 sg13g2_decap_8 FILLER_36_227 ();
 sg13g2_decap_8 FILLER_36_234 ();
 sg13g2_decap_8 FILLER_36_241 ();
 sg13g2_decap_8 FILLER_36_248 ();
 sg13g2_decap_8 FILLER_36_255 ();
 sg13g2_decap_8 FILLER_36_262 ();
 sg13g2_fill_2 FILLER_36_269 ();
 sg13g2_fill_1 FILLER_36_271 ();
 sg13g2_decap_4 FILLER_36_294 ();
 sg13g2_fill_1 FILLER_36_298 ();
 sg13g2_fill_2 FILLER_36_302 ();
 sg13g2_decap_4 FILLER_36_307 ();
 sg13g2_decap_8 FILLER_36_319 ();
 sg13g2_fill_1 FILLER_36_326 ();
 sg13g2_decap_4 FILLER_36_331 ();
 sg13g2_fill_1 FILLER_36_335 ();
 sg13g2_decap_8 FILLER_36_355 ();
 sg13g2_fill_1 FILLER_36_362 ();
 sg13g2_decap_8 FILLER_36_366 ();
 sg13g2_decap_8 FILLER_36_373 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_fill_2 FILLER_37_147 ();
 sg13g2_fill_1 FILLER_37_149 ();
 sg13g2_decap_8 FILLER_37_211 ();
 sg13g2_decap_8 FILLER_37_218 ();
 sg13g2_decap_8 FILLER_37_225 ();
 sg13g2_decap_8 FILLER_37_232 ();
 sg13g2_decap_8 FILLER_37_239 ();
 sg13g2_decap_8 FILLER_37_246 ();
 sg13g2_decap_8 FILLER_37_253 ();
 sg13g2_decap_8 FILLER_37_260 ();
 sg13g2_decap_8 FILLER_37_267 ();
 sg13g2_decap_8 FILLER_37_274 ();
 sg13g2_decap_4 FILLER_37_281 ();
 sg13g2_fill_1 FILLER_37_285 ();
 sg13g2_fill_2 FILLER_37_300 ();
 sg13g2_fill_1 FILLER_37_312 ();
 sg13g2_decap_8 FILLER_37_325 ();
 sg13g2_fill_1 FILLER_37_358 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_4 FILLER_38_133 ();
 sg13g2_fill_2 FILLER_38_137 ();
 sg13g2_decap_8 FILLER_38_206 ();
 sg13g2_decap_8 FILLER_38_213 ();
 sg13g2_decap_8 FILLER_38_220 ();
 sg13g2_decap_4 FILLER_38_227 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_250 ();
 sg13g2_decap_8 FILLER_38_257 ();
 sg13g2_decap_8 FILLER_38_264 ();
 sg13g2_fill_2 FILLER_38_330 ();
 sg13g2_fill_1 FILLER_38_351 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_4 FILLER_39_133 ();
 sg13g2_fill_2 FILLER_39_137 ();
 sg13g2_fill_2 FILLER_39_184 ();
 sg13g2_fill_1 FILLER_39_186 ();
 sg13g2_decap_8 FILLER_39_206 ();
 sg13g2_decap_8 FILLER_39_213 ();
 sg13g2_decap_8 FILLER_39_220 ();
 sg13g2_decap_8 FILLER_39_227 ();
 sg13g2_decap_8 FILLER_39_234 ();
 sg13g2_decap_8 FILLER_39_241 ();
 sg13g2_decap_8 FILLER_39_248 ();
 sg13g2_decap_4 FILLER_39_321 ();
 sg13g2_fill_1 FILLER_39_325 ();
 sg13g2_decap_8 FILLER_39_377 ();
 sg13g2_decap_8 FILLER_39_384 ();
 sg13g2_decap_8 FILLER_39_391 ();
 sg13g2_decap_8 FILLER_39_398 ();
 sg13g2_decap_4 FILLER_39_405 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_fill_1 FILLER_40_165 ();
 sg13g2_decap_8 FILLER_40_205 ();
 sg13g2_decap_8 FILLER_40_212 ();
 sg13g2_decap_8 FILLER_40_219 ();
 sg13g2_decap_8 FILLER_40_226 ();
 sg13g2_decap_8 FILLER_40_233 ();
 sg13g2_decap_8 FILLER_40_240 ();
 sg13g2_decap_8 FILLER_40_247 ();
 sg13g2_fill_2 FILLER_40_254 ();
 sg13g2_decap_8 FILLER_40_312 ();
 sg13g2_fill_1 FILLER_40_319 ();
 sg13g2_decap_8 FILLER_40_324 ();
 sg13g2_decap_8 FILLER_40_331 ();
 sg13g2_fill_1 FILLER_40_338 ();
 sg13g2_decap_8 FILLER_40_352 ();
 sg13g2_decap_8 FILLER_40_359 ();
 sg13g2_decap_8 FILLER_40_392 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_fill_2 FILLER_40_406 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_4 FILLER_41_147 ();
 sg13g2_fill_2 FILLER_41_151 ();
 sg13g2_decap_4 FILLER_41_166 ();
 sg13g2_fill_2 FILLER_41_178 ();
 sg13g2_decap_8 FILLER_41_222 ();
 sg13g2_decap_8 FILLER_41_229 ();
 sg13g2_decap_8 FILLER_41_236 ();
 sg13g2_decap_8 FILLER_41_243 ();
 sg13g2_decap_8 FILLER_41_250 ();
 sg13g2_decap_8 FILLER_41_257 ();
 sg13g2_fill_2 FILLER_41_264 ();
 sg13g2_fill_2 FILLER_41_306 ();
 sg13g2_fill_1 FILLER_41_308 ();
 sg13g2_fill_1 FILLER_41_345 ();
 sg13g2_decap_4 FILLER_41_350 ();
 sg13g2_fill_1 FILLER_41_354 ();
 sg13g2_fill_1 FILLER_41_363 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_fill_2 FILLER_41_406 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_4 FILLER_42_133 ();
 sg13g2_fill_1 FILLER_42_137 ();
 sg13g2_fill_2 FILLER_42_175 ();
 sg13g2_fill_1 FILLER_42_177 ();
 sg13g2_fill_1 FILLER_42_210 ();
 sg13g2_decap_8 FILLER_42_224 ();
 sg13g2_decap_8 FILLER_42_231 ();
 sg13g2_decap_8 FILLER_42_238 ();
 sg13g2_decap_8 FILLER_42_245 ();
 sg13g2_decap_8 FILLER_42_252 ();
 sg13g2_decap_8 FILLER_42_259 ();
 sg13g2_fill_2 FILLER_42_266 ();
 sg13g2_fill_1 FILLER_42_268 ();
 sg13g2_fill_1 FILLER_42_273 ();
 sg13g2_fill_2 FILLER_42_308 ();
 sg13g2_decap_8 FILLER_42_389 ();
 sg13g2_decap_8 FILLER_42_396 ();
 sg13g2_decap_4 FILLER_42_403 ();
 sg13g2_fill_2 FILLER_42_407 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_4 FILLER_43_140 ();
 sg13g2_fill_1 FILLER_43_144 ();
 sg13g2_fill_1 FILLER_43_152 ();
 sg13g2_decap_8 FILLER_43_217 ();
 sg13g2_decap_8 FILLER_43_224 ();
 sg13g2_decap_8 FILLER_43_231 ();
 sg13g2_decap_8 FILLER_43_238 ();
 sg13g2_decap_8 FILLER_43_245 ();
 sg13g2_decap_8 FILLER_43_252 ();
 sg13g2_fill_1 FILLER_43_322 ();
 sg13g2_fill_2 FILLER_43_362 ();
 sg13g2_fill_1 FILLER_43_364 ();
 sg13g2_decap_8 FILLER_43_388 ();
 sg13g2_decap_8 FILLER_43_395 ();
 sg13g2_decap_8 FILLER_43_402 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_decap_4 FILLER_44_140 ();
 sg13g2_fill_2 FILLER_44_144 ();
 sg13g2_fill_1 FILLER_44_168 ();
 sg13g2_fill_1 FILLER_44_184 ();
 sg13g2_fill_1 FILLER_44_194 ();
 sg13g2_decap_8 FILLER_44_216 ();
 sg13g2_fill_2 FILLER_44_223 ();
 sg13g2_fill_2 FILLER_44_234 ();
 sg13g2_decap_4 FILLER_44_241 ();
 sg13g2_fill_1 FILLER_44_245 ();
 sg13g2_decap_4 FILLER_44_249 ();
 sg13g2_fill_1 FILLER_44_253 ();
 sg13g2_fill_2 FILLER_44_322 ();
 sg13g2_fill_1 FILLER_44_371 ();
 sg13g2_decap_4 FILLER_44_404 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_fill_2 FILLER_45_147 ();
 sg13g2_fill_2 FILLER_45_210 ();
 sg13g2_decap_4 FILLER_45_215 ();
 sg13g2_fill_1 FILLER_45_219 ();
 sg13g2_fill_1 FILLER_45_250 ();
 sg13g2_fill_1 FILLER_45_255 ();
 sg13g2_fill_1 FILLER_45_273 ();
 sg13g2_fill_2 FILLER_45_279 ();
 sg13g2_fill_1 FILLER_45_298 ();
 sg13g2_fill_2 FILLER_45_330 ();
 sg13g2_fill_1 FILLER_45_332 ();
 sg13g2_fill_2 FILLER_45_342 ();
 sg13g2_fill_1 FILLER_45_344 ();
 sg13g2_decap_8 FILLER_45_363 ();
 sg13g2_fill_1 FILLER_45_386 ();
 sg13g2_decap_8 FILLER_45_390 ();
 sg13g2_decap_8 FILLER_45_397 ();
 sg13g2_decap_4 FILLER_45_404 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_fill_2 FILLER_46_119 ();
 sg13g2_fill_1 FILLER_46_121 ();
 sg13g2_fill_2 FILLER_46_131 ();
 sg13g2_fill_1 FILLER_46_163 ();
 sg13g2_fill_1 FILLER_46_262 ();
 sg13g2_fill_2 FILLER_46_268 ();
 sg13g2_decap_4 FILLER_46_281 ();
 sg13g2_fill_2 FILLER_46_320 ();
 sg13g2_decap_4 FILLER_46_370 ();
 sg13g2_fill_2 FILLER_46_374 ();
 sg13g2_decap_8 FILLER_46_384 ();
 sg13g2_fill_1 FILLER_46_391 ();
 sg13g2_decap_8 FILLER_46_395 ();
 sg13g2_decap_8 FILLER_46_402 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_fill_2 FILLER_47_168 ();
 sg13g2_fill_2 FILLER_47_190 ();
 sg13g2_fill_1 FILLER_47_288 ();
 sg13g2_decap_4 FILLER_47_298 ();
 sg13g2_fill_2 FILLER_47_302 ();
 sg13g2_decap_4 FILLER_47_348 ();
 sg13g2_fill_1 FILLER_47_378 ();
 sg13g2_fill_1 FILLER_47_382 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_fill_2 FILLER_48_98 ();
 sg13g2_fill_2 FILLER_48_126 ();
 sg13g2_fill_2 FILLER_48_152 ();
 sg13g2_fill_1 FILLER_48_154 ();
 sg13g2_fill_2 FILLER_48_195 ();
 sg13g2_fill_2 FILLER_48_220 ();
 sg13g2_fill_2 FILLER_48_236 ();
 sg13g2_fill_1 FILLER_48_263 ();
 sg13g2_fill_1 FILLER_48_341 ();
 sg13g2_decap_8 FILLER_48_377 ();
 sg13g2_decap_8 FILLER_48_384 ();
 sg13g2_fill_1 FILLER_48_391 ();
 sg13g2_decap_8 FILLER_48_395 ();
 sg13g2_decap_8 FILLER_48_402 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_4 FILLER_49_98 ();
 sg13g2_fill_1 FILLER_49_155 ();
 sg13g2_fill_1 FILLER_49_182 ();
 sg13g2_fill_1 FILLER_49_193 ();
 sg13g2_fill_2 FILLER_49_253 ();
 sg13g2_decap_8 FILLER_49_317 ();
 sg13g2_decap_8 FILLER_49_324 ();
 sg13g2_fill_1 FILLER_49_331 ();
 sg13g2_fill_2 FILLER_49_336 ();
 sg13g2_decap_4 FILLER_49_343 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_fill_2 FILLER_50_112 ();
 sg13g2_fill_2 FILLER_50_137 ();
 sg13g2_fill_2 FILLER_50_144 ();
 sg13g2_fill_1 FILLER_50_146 ();
 sg13g2_fill_2 FILLER_50_169 ();
 sg13g2_fill_1 FILLER_50_171 ();
 sg13g2_fill_1 FILLER_50_230 ();
 sg13g2_fill_2 FILLER_50_245 ();
 sg13g2_fill_2 FILLER_50_265 ();
 sg13g2_fill_2 FILLER_50_281 ();
 sg13g2_fill_1 FILLER_50_297 ();
 sg13g2_fill_2 FILLER_50_311 ();
 sg13g2_fill_1 FILLER_50_313 ();
 sg13g2_decap_8 FILLER_50_317 ();
 sg13g2_decap_4 FILLER_50_324 ();
 sg13g2_fill_2 FILLER_50_328 ();
 sg13g2_decap_8 FILLER_50_339 ();
 sg13g2_fill_1 FILLER_50_346 ();
 sg13g2_fill_2 FILLER_50_352 ();
 sg13g2_fill_2 FILLER_50_363 ();
 sg13g2_fill_2 FILLER_50_369 ();
 sg13g2_decap_8 FILLER_50_400 ();
 sg13g2_fill_2 FILLER_50_407 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_4 FILLER_51_91 ();
 sg13g2_fill_1 FILLER_51_126 ();
 sg13g2_fill_2 FILLER_51_143 ();
 sg13g2_fill_2 FILLER_51_150 ();
 sg13g2_fill_1 FILLER_51_152 ();
 sg13g2_fill_2 FILLER_51_244 ();
 sg13g2_fill_1 FILLER_51_287 ();
 sg13g2_fill_1 FILLER_51_305 ();
 sg13g2_decap_4 FILLER_51_328 ();
 sg13g2_fill_2 FILLER_51_332 ();
 sg13g2_decap_4 FILLER_51_360 ();
 sg13g2_fill_2 FILLER_51_364 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_fill_1 FILLER_52_91 ();
 sg13g2_fill_2 FILLER_52_114 ();
 sg13g2_fill_1 FILLER_52_116 ();
 sg13g2_fill_1 FILLER_52_143 ();
 sg13g2_fill_1 FILLER_52_154 ();
 sg13g2_fill_2 FILLER_52_166 ();
 sg13g2_fill_1 FILLER_52_168 ();
 sg13g2_fill_1 FILLER_52_204 ();
 sg13g2_fill_1 FILLER_52_227 ();
 sg13g2_fill_1 FILLER_52_287 ();
 sg13g2_fill_2 FILLER_52_331 ();
 sg13g2_fill_2 FILLER_52_377 ();
 sg13g2_fill_1 FILLER_52_379 ();
 sg13g2_fill_2 FILLER_52_389 ();
 sg13g2_fill_1 FILLER_52_391 ();
 sg13g2_decap_8 FILLER_52_395 ();
 sg13g2_decap_8 FILLER_52_402 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_4 FILLER_53_91 ();
 sg13g2_fill_2 FILLER_53_149 ();
 sg13g2_fill_2 FILLER_53_159 ();
 sg13g2_fill_1 FILLER_53_161 ();
 sg13g2_fill_1 FILLER_53_192 ();
 sg13g2_fill_2 FILLER_53_208 ();
 sg13g2_fill_2 FILLER_53_227 ();
 sg13g2_fill_1 FILLER_53_242 ();
 sg13g2_fill_2 FILLER_53_257 ();
 sg13g2_fill_1 FILLER_53_259 ();
 sg13g2_fill_2 FILLER_53_351 ();
 sg13g2_fill_1 FILLER_53_353 ();
 sg13g2_fill_2 FILLER_53_373 ();
 sg13g2_fill_1 FILLER_53_375 ();
 sg13g2_decap_8 FILLER_53_391 ();
 sg13g2_decap_8 FILLER_53_398 ();
 sg13g2_decap_4 FILLER_53_405 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_fill_1 FILLER_54_105 ();
 sg13g2_decap_4 FILLER_54_110 ();
 sg13g2_fill_1 FILLER_54_155 ();
 sg13g2_fill_1 FILLER_54_168 ();
 sg13g2_fill_2 FILLER_54_187 ();
 sg13g2_fill_1 FILLER_54_189 ();
 sg13g2_fill_1 FILLER_54_281 ();
 sg13g2_fill_1 FILLER_54_312 ();
 sg13g2_fill_2 FILLER_54_381 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_4 FILLER_55_105 ();
 sg13g2_fill_1 FILLER_55_109 ();
 sg13g2_fill_2 FILLER_55_135 ();
 sg13g2_fill_1 FILLER_55_159 ();
 sg13g2_fill_2 FILLER_55_252 ();
 sg13g2_fill_1 FILLER_55_254 ();
 sg13g2_fill_2 FILLER_55_262 ();
 sg13g2_fill_2 FILLER_55_271 ();
 sg13g2_fill_1 FILLER_55_273 ();
 sg13g2_fill_2 FILLER_55_290 ();
 sg13g2_fill_2 FILLER_55_332 ();
 sg13g2_decap_4 FILLER_55_371 ();
 sg13g2_fill_2 FILLER_55_375 ();
 sg13g2_fill_1 FILLER_55_391 ();
 sg13g2_decap_8 FILLER_55_395 ();
 sg13g2_decap_8 FILLER_55_402 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_fill_2 FILLER_56_123 ();
 sg13g2_fill_1 FILLER_56_164 ();
 sg13g2_decap_4 FILLER_56_241 ();
 sg13g2_decap_8 FILLER_56_360 ();
 sg13g2_decap_8 FILLER_56_367 ();
 sg13g2_fill_2 FILLER_56_374 ();
 sg13g2_fill_1 FILLER_56_376 ();
 sg13g2_fill_2 FILLER_56_389 ();
 sg13g2_decap_8 FILLER_56_399 ();
 sg13g2_fill_2 FILLER_56_406 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_4 FILLER_57_98 ();
 sg13g2_fill_2 FILLER_57_153 ();
 sg13g2_fill_1 FILLER_57_155 ();
 sg13g2_fill_2 FILLER_57_161 ();
 sg13g2_fill_1 FILLER_57_199 ();
 sg13g2_fill_2 FILLER_57_231 ();
 sg13g2_fill_1 FILLER_57_233 ();
 sg13g2_decap_4 FILLER_57_242 ();
 sg13g2_fill_1 FILLER_57_276 ();
 sg13g2_fill_2 FILLER_57_312 ();
 sg13g2_fill_1 FILLER_57_314 ();
 sg13g2_fill_1 FILLER_57_341 ();
 sg13g2_fill_2 FILLER_57_350 ();
 sg13g2_fill_1 FILLER_57_352 ();
 sg13g2_fill_1 FILLER_57_382 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_4 FILLER_58_98 ();
 sg13g2_fill_2 FILLER_58_102 ();
 sg13g2_decap_8 FILLER_58_113 ();
 sg13g2_decap_4 FILLER_58_120 ();
 sg13g2_fill_2 FILLER_58_124 ();
 sg13g2_decap_4 FILLER_58_145 ();
 sg13g2_fill_2 FILLER_58_170 ();
 sg13g2_fill_1 FILLER_58_172 ();
 sg13g2_fill_2 FILLER_58_178 ();
 sg13g2_fill_1 FILLER_58_180 ();
 sg13g2_fill_2 FILLER_58_191 ();
 sg13g2_fill_1 FILLER_58_193 ();
 sg13g2_fill_1 FILLER_58_207 ();
 sg13g2_decap_8 FILLER_58_220 ();
 sg13g2_fill_1 FILLER_58_227 ();
 sg13g2_decap_4 FILLER_58_245 ();
 sg13g2_fill_1 FILLER_58_249 ();
 sg13g2_fill_1 FILLER_58_268 ();
 sg13g2_fill_2 FILLER_58_304 ();
 sg13g2_fill_1 FILLER_58_306 ();
 sg13g2_fill_2 FILLER_58_340 ();
 sg13g2_fill_1 FILLER_58_382 ();
 sg13g2_decap_8 FILLER_58_401 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_4 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_113 ();
 sg13g2_decap_8 FILLER_59_120 ();
 sg13g2_decap_8 FILLER_59_127 ();
 sg13g2_decap_8 FILLER_59_134 ();
 sg13g2_decap_4 FILLER_59_141 ();
 sg13g2_fill_2 FILLER_59_145 ();
 sg13g2_fill_1 FILLER_59_158 ();
 sg13g2_fill_1 FILLER_59_164 ();
 sg13g2_decap_4 FILLER_59_170 ();
 sg13g2_fill_1 FILLER_59_174 ();
 sg13g2_fill_1 FILLER_59_181 ();
 sg13g2_fill_2 FILLER_59_187 ();
 sg13g2_decap_8 FILLER_59_209 ();
 sg13g2_decap_4 FILLER_59_216 ();
 sg13g2_fill_1 FILLER_59_220 ();
 sg13g2_decap_8 FILLER_59_229 ();
 sg13g2_decap_8 FILLER_59_236 ();
 sg13g2_decap_8 FILLER_59_243 ();
 sg13g2_decap_8 FILLER_59_250 ();
 sg13g2_decap_8 FILLER_59_261 ();
 sg13g2_decap_8 FILLER_59_268 ();
 sg13g2_fill_1 FILLER_59_275 ();
 sg13g2_fill_2 FILLER_59_279 ();
 sg13g2_fill_1 FILLER_59_281 ();
 sg13g2_fill_2 FILLER_59_286 ();
 sg13g2_decap_4 FILLER_59_338 ();
 sg13g2_fill_2 FILLER_59_342 ();
 sg13g2_fill_1 FILLER_59_382 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_fill_2 FILLER_60_91 ();
 sg13g2_fill_1 FILLER_60_93 ();
 sg13g2_decap_8 FILLER_60_120 ();
 sg13g2_decap_8 FILLER_60_127 ();
 sg13g2_decap_4 FILLER_60_134 ();
 sg13g2_decap_8 FILLER_60_142 ();
 sg13g2_decap_4 FILLER_60_149 ();
 sg13g2_fill_1 FILLER_60_153 ();
 sg13g2_decap_8 FILLER_60_157 ();
 sg13g2_fill_2 FILLER_60_164 ();
 sg13g2_fill_1 FILLER_60_166 ();
 sg13g2_decap_8 FILLER_60_201 ();
 sg13g2_fill_1 FILLER_60_208 ();
 sg13g2_fill_1 FILLER_60_239 ();
 sg13g2_fill_2 FILLER_60_244 ();
 sg13g2_decap_8 FILLER_60_329 ();
 sg13g2_decap_8 FILLER_60_336 ();
 sg13g2_fill_2 FILLER_60_343 ();
 sg13g2_fill_2 FILLER_60_354 ();
 sg13g2_fill_1 FILLER_60_378 ();
 sg13g2_decap_8 FILLER_60_401 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_4 FILLER_61_84 ();
 sg13g2_fill_2 FILLER_61_125 ();
 sg13g2_decap_8 FILLER_61_153 ();
 sg13g2_fill_2 FILLER_61_160 ();
 sg13g2_fill_2 FILLER_61_194 ();
 sg13g2_fill_1 FILLER_61_196 ();
 sg13g2_fill_1 FILLER_61_280 ();
 sg13g2_decap_8 FILLER_61_285 ();
 sg13g2_decap_8 FILLER_61_292 ();
 sg13g2_decap_8 FILLER_61_299 ();
 sg13g2_fill_2 FILLER_61_306 ();
 sg13g2_fill_1 FILLER_61_331 ();
 sg13g2_fill_2 FILLER_61_367 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_fill_2 FILLER_62_91 ();
 sg13g2_fill_1 FILLER_62_134 ();
 sg13g2_fill_1 FILLER_62_181 ();
 sg13g2_fill_1 FILLER_62_225 ();
 sg13g2_fill_2 FILLER_62_249 ();
 sg13g2_decap_4 FILLER_62_277 ();
 sg13g2_fill_1 FILLER_62_281 ();
 sg13g2_decap_8 FILLER_62_290 ();
 sg13g2_fill_1 FILLER_62_297 ();
 sg13g2_decap_4 FILLER_62_307 ();
 sg13g2_fill_1 FILLER_62_311 ();
 sg13g2_fill_1 FILLER_62_321 ();
 sg13g2_fill_2 FILLER_62_359 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_4 FILLER_63_84 ();
 sg13g2_fill_1 FILLER_63_115 ();
 sg13g2_fill_1 FILLER_63_122 ();
 sg13g2_fill_1 FILLER_63_133 ();
 sg13g2_fill_2 FILLER_63_178 ();
 sg13g2_fill_1 FILLER_63_180 ();
 sg13g2_decap_4 FILLER_63_191 ();
 sg13g2_fill_1 FILLER_63_195 ();
 sg13g2_fill_2 FILLER_63_255 ();
 sg13g2_fill_2 FILLER_63_261 ();
 sg13g2_fill_2 FILLER_63_283 ();
 sg13g2_fill_1 FILLER_63_285 ();
 sg13g2_fill_1 FILLER_63_290 ();
 sg13g2_fill_2 FILLER_63_314 ();
 sg13g2_fill_2 FILLER_63_345 ();
 sg13g2_decap_8 FILLER_63_400 ();
 sg13g2_fill_2 FILLER_63_407 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_fill_1 FILLER_64_98 ();
 sg13g2_fill_2 FILLER_64_104 ();
 sg13g2_fill_1 FILLER_64_106 ();
 sg13g2_fill_2 FILLER_64_119 ();
 sg13g2_fill_1 FILLER_64_121 ();
 sg13g2_decap_4 FILLER_64_137 ();
 sg13g2_fill_2 FILLER_64_141 ();
 sg13g2_fill_2 FILLER_64_148 ();
 sg13g2_decap_8 FILLER_64_158 ();
 sg13g2_decap_4 FILLER_64_165 ();
 sg13g2_decap_4 FILLER_64_183 ();
 sg13g2_fill_1 FILLER_64_274 ();
 sg13g2_fill_2 FILLER_64_313 ();
 sg13g2_fill_1 FILLER_64_327 ();
 sg13g2_fill_1 FILLER_64_363 ();
 sg13g2_decap_8 FILLER_64_388 ();
 sg13g2_decap_8 FILLER_64_395 ();
 sg13g2_decap_8 FILLER_64_402 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_4 FILLER_65_84 ();
 sg13g2_fill_1 FILLER_65_110 ();
 sg13g2_fill_2 FILLER_65_115 ();
 sg13g2_fill_1 FILLER_65_117 ();
 sg13g2_decap_4 FILLER_65_127 ();
 sg13g2_fill_2 FILLER_65_131 ();
 sg13g2_fill_2 FILLER_65_224 ();
 sg13g2_fill_1 FILLER_65_226 ();
 sg13g2_fill_1 FILLER_65_301 ();
 sg13g2_decap_8 FILLER_65_347 ();
 sg13g2_decap_8 FILLER_65_389 ();
 sg13g2_decap_8 FILLER_65_396 ();
 sg13g2_decap_4 FILLER_65_403 ();
 sg13g2_fill_2 FILLER_65_407 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_4 FILLER_66_84 ();
 sg13g2_fill_2 FILLER_66_113 ();
 sg13g2_fill_1 FILLER_66_115 ();
 sg13g2_decap_8 FILLER_66_136 ();
 sg13g2_decap_4 FILLER_66_143 ();
 sg13g2_decap_8 FILLER_66_151 ();
 sg13g2_fill_2 FILLER_66_158 ();
 sg13g2_fill_1 FILLER_66_193 ();
 sg13g2_fill_2 FILLER_66_208 ();
 sg13g2_fill_1 FILLER_66_210 ();
 sg13g2_fill_2 FILLER_66_242 ();
 sg13g2_decap_8 FILLER_66_297 ();
 sg13g2_decap_8 FILLER_66_304 ();
 sg13g2_fill_2 FILLER_66_311 ();
 sg13g2_fill_1 FILLER_66_313 ();
 sg13g2_fill_1 FILLER_66_325 ();
 sg13g2_decap_8 FILLER_66_340 ();
 sg13g2_decap_8 FILLER_66_347 ();
 sg13g2_decap_8 FILLER_66_354 ();
 sg13g2_decap_4 FILLER_66_361 ();
 sg13g2_decap_8 FILLER_66_369 ();
 sg13g2_decap_8 FILLER_66_402 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_fill_1 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_130 ();
 sg13g2_decap_8 FILLER_67_163 ();
 sg13g2_fill_1 FILLER_67_170 ();
 sg13g2_fill_2 FILLER_67_197 ();
 sg13g2_fill_2 FILLER_67_208 ();
 sg13g2_fill_1 FILLER_67_266 ();
 sg13g2_decap_4 FILLER_67_281 ();
 sg13g2_fill_2 FILLER_67_285 ();
 sg13g2_fill_2 FILLER_67_296 ();
 sg13g2_decap_4 FILLER_67_307 ();
 sg13g2_decap_8 FILLER_67_316 ();
 sg13g2_decap_8 FILLER_67_331 ();
 sg13g2_decap_8 FILLER_67_338 ();
 sg13g2_fill_2 FILLER_67_345 ();
 sg13g2_fill_1 FILLER_67_347 ();
 sg13g2_decap_8 FILLER_67_352 ();
 sg13g2_fill_1 FILLER_67_359 ();
 sg13g2_decap_8 FILLER_67_387 ();
 sg13g2_decap_8 FILLER_67_394 ();
 sg13g2_decap_8 FILLER_67_401 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_4 FILLER_68_98 ();
 sg13g2_fill_1 FILLER_68_102 ();
 sg13g2_fill_1 FILLER_68_114 ();
 sg13g2_fill_2 FILLER_68_136 ();
 sg13g2_decap_8 FILLER_68_169 ();
 sg13g2_fill_2 FILLER_68_176 ();
 sg13g2_fill_2 FILLER_68_218 ();
 sg13g2_fill_1 FILLER_68_230 ();
 sg13g2_decap_4 FILLER_68_251 ();
 sg13g2_fill_1 FILLER_68_255 ();
 sg13g2_fill_1 FILLER_68_307 ();
 sg13g2_decap_8 FILLER_68_326 ();
 sg13g2_fill_2 FILLER_68_378 ();
 sg13g2_decap_8 FILLER_68_398 ();
 sg13g2_decap_4 FILLER_68_405 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_4 FILLER_69_91 ();
 sg13g2_fill_1 FILLER_69_117 ();
 sg13g2_decap_8 FILLER_69_123 ();
 sg13g2_decap_8 FILLER_69_130 ();
 sg13g2_fill_2 FILLER_69_137 ();
 sg13g2_decap_4 FILLER_69_143 ();
 sg13g2_fill_2 FILLER_69_151 ();
 sg13g2_decap_4 FILLER_69_160 ();
 sg13g2_fill_1 FILLER_69_164 ();
 sg13g2_fill_2 FILLER_69_181 ();
 sg13g2_fill_1 FILLER_69_183 ();
 sg13g2_fill_2 FILLER_69_198 ();
 sg13g2_fill_1 FILLER_69_200 ();
 sg13g2_fill_2 FILLER_69_242 ();
 sg13g2_fill_1 FILLER_69_244 ();
 sg13g2_fill_1 FILLER_69_265 ();
 sg13g2_fill_2 FILLER_69_291 ();
 sg13g2_fill_1 FILLER_69_293 ();
 sg13g2_decap_8 FILLER_69_324 ();
 sg13g2_fill_2 FILLER_69_331 ();
 sg13g2_fill_2 FILLER_69_373 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_4 FILLER_70_84 ();
 sg13g2_fill_1 FILLER_70_128 ();
 sg13g2_fill_2 FILLER_70_155 ();
 sg13g2_fill_1 FILLER_70_157 ();
 sg13g2_decap_4 FILLER_70_176 ();
 sg13g2_fill_1 FILLER_70_270 ();
 sg13g2_fill_2 FILLER_70_283 ();
 sg13g2_decap_8 FILLER_70_328 ();
 sg13g2_fill_2 FILLER_70_370 ();
 sg13g2_fill_1 FILLER_70_372 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_4 FILLER_71_84 ();
 sg13g2_fill_1 FILLER_71_88 ();
 sg13g2_fill_2 FILLER_71_120 ();
 sg13g2_fill_1 FILLER_71_122 ();
 sg13g2_fill_2 FILLER_71_137 ();
 sg13g2_fill_1 FILLER_71_139 ();
 sg13g2_fill_2 FILLER_71_200 ();
 sg13g2_fill_1 FILLER_71_202 ();
 sg13g2_fill_1 FILLER_71_260 ();
 sg13g2_fill_2 FILLER_71_281 ();
 sg13g2_fill_2 FILLER_71_304 ();
 sg13g2_decap_8 FILLER_71_318 ();
 sg13g2_decap_8 FILLER_71_325 ();
 sg13g2_fill_2 FILLER_71_332 ();
 sg13g2_decap_8 FILLER_71_339 ();
 sg13g2_fill_1 FILLER_71_350 ();
 sg13g2_fill_1 FILLER_71_360 ();
 sg13g2_fill_2 FILLER_71_381 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_fill_2 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_132 ();
 sg13g2_decap_8 FILLER_72_139 ();
 sg13g2_decap_4 FILLER_72_146 ();
 sg13g2_fill_1 FILLER_72_150 ();
 sg13g2_fill_1 FILLER_72_155 ();
 sg13g2_fill_1 FILLER_72_160 ();
 sg13g2_fill_2 FILLER_72_208 ();
 sg13g2_fill_1 FILLER_72_219 ();
 sg13g2_fill_2 FILLER_72_232 ();
 sg13g2_fill_2 FILLER_72_238 ();
 sg13g2_fill_1 FILLER_72_275 ();
 sg13g2_decap_8 FILLER_72_297 ();
 sg13g2_decap_8 FILLER_72_304 ();
 sg13g2_decap_8 FILLER_72_311 ();
 sg13g2_decap_8 FILLER_72_318 ();
 sg13g2_decap_8 FILLER_72_325 ();
 sg13g2_decap_8 FILLER_72_332 ();
 sg13g2_decap_8 FILLER_72_339 ();
 sg13g2_fill_2 FILLER_72_346 ();
 sg13g2_decap_8 FILLER_72_400 ();
 sg13g2_fill_2 FILLER_72_407 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_4 FILLER_73_103 ();
 sg13g2_fill_1 FILLER_73_107 ();
 sg13g2_fill_2 FILLER_73_113 ();
 sg13g2_fill_1 FILLER_73_115 ();
 sg13g2_fill_2 FILLER_73_121 ();
 sg13g2_fill_1 FILLER_73_123 ();
 sg13g2_fill_1 FILLER_73_154 ();
 sg13g2_fill_2 FILLER_73_169 ();
 sg13g2_fill_2 FILLER_73_176 ();
 sg13g2_fill_1 FILLER_73_178 ();
 sg13g2_fill_1 FILLER_73_221 ();
 sg13g2_decap_8 FILLER_73_292 ();
 sg13g2_decap_8 FILLER_73_299 ();
 sg13g2_decap_8 FILLER_73_306 ();
 sg13g2_decap_8 FILLER_73_313 ();
 sg13g2_decap_8 FILLER_73_320 ();
 sg13g2_decap_8 FILLER_73_327 ();
 sg13g2_decap_8 FILLER_73_334 ();
 sg13g2_decap_8 FILLER_73_341 ();
 sg13g2_decap_8 FILLER_73_348 ();
 sg13g2_decap_4 FILLER_73_355 ();
 sg13g2_decap_4 FILLER_73_363 ();
 sg13g2_fill_1 FILLER_73_367 ();
 sg13g2_decap_8 FILLER_73_381 ();
 sg13g2_decap_8 FILLER_73_388 ();
 sg13g2_decap_8 FILLER_73_395 ();
 sg13g2_decap_8 FILLER_73_402 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_4 FILLER_74_119 ();
 sg13g2_fill_2 FILLER_74_123 ();
 sg13g2_fill_1 FILLER_74_151 ();
 sg13g2_fill_2 FILLER_74_209 ();
 sg13g2_fill_1 FILLER_74_211 ();
 sg13g2_fill_2 FILLER_74_285 ();
 sg13g2_fill_1 FILLER_74_287 ();
 sg13g2_decap_8 FILLER_74_317 ();
 sg13g2_decap_8 FILLER_74_324 ();
 sg13g2_decap_8 FILLER_74_331 ();
 sg13g2_decap_8 FILLER_74_338 ();
 sg13g2_decap_8 FILLER_74_345 ();
 sg13g2_decap_8 FILLER_74_352 ();
 sg13g2_decap_8 FILLER_74_359 ();
 sg13g2_decap_8 FILLER_74_366 ();
 sg13g2_decap_8 FILLER_74_373 ();
 sg13g2_decap_8 FILLER_74_380 ();
 sg13g2_decap_8 FILLER_74_387 ();
 sg13g2_decap_8 FILLER_74_394 ();
 sg13g2_decap_8 FILLER_74_401 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_fill_1 FILLER_75_133 ();
 sg13g2_fill_2 FILLER_75_187 ();
 sg13g2_fill_1 FILLER_75_189 ();
 sg13g2_fill_1 FILLER_75_199 ();
 sg13g2_decap_8 FILLER_75_281 ();
 sg13g2_decap_8 FILLER_75_288 ();
 sg13g2_decap_4 FILLER_75_295 ();
 sg13g2_decap_8 FILLER_75_303 ();
 sg13g2_decap_8 FILLER_75_310 ();
 sg13g2_decap_8 FILLER_75_317 ();
 sg13g2_decap_8 FILLER_75_324 ();
 sg13g2_decap_8 FILLER_75_331 ();
 sg13g2_decap_8 FILLER_75_338 ();
 sg13g2_decap_8 FILLER_75_345 ();
 sg13g2_decap_8 FILLER_75_352 ();
 sg13g2_decap_8 FILLER_75_359 ();
 sg13g2_decap_8 FILLER_75_366 ();
 sg13g2_decap_8 FILLER_75_373 ();
 sg13g2_decap_8 FILLER_75_380 ();
 sg13g2_decap_8 FILLER_75_387 ();
 sg13g2_decap_8 FILLER_75_394 ();
 sg13g2_decap_8 FILLER_75_401 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_4 FILLER_76_133 ();
 sg13g2_fill_1 FILLER_76_137 ();
 sg13g2_fill_2 FILLER_76_160 ();
 sg13g2_fill_2 FILLER_76_176 ();
 sg13g2_fill_1 FILLER_76_178 ();
 sg13g2_fill_1 FILLER_76_188 ();
 sg13g2_fill_2 FILLER_76_203 ();
 sg13g2_fill_1 FILLER_76_205 ();
 sg13g2_fill_2 FILLER_76_220 ();
 sg13g2_fill_1 FILLER_76_240 ();
 sg13g2_decap_8 FILLER_76_273 ();
 sg13g2_decap_8 FILLER_76_280 ();
 sg13g2_decap_8 FILLER_76_287 ();
 sg13g2_decap_8 FILLER_76_294 ();
 sg13g2_decap_8 FILLER_76_301 ();
 sg13g2_decap_8 FILLER_76_308 ();
 sg13g2_decap_8 FILLER_76_315 ();
 sg13g2_decap_8 FILLER_76_322 ();
 sg13g2_decap_8 FILLER_76_329 ();
 sg13g2_decap_8 FILLER_76_336 ();
 sg13g2_decap_8 FILLER_76_343 ();
 sg13g2_decap_8 FILLER_76_350 ();
 sg13g2_decap_8 FILLER_76_357 ();
 sg13g2_decap_8 FILLER_76_364 ();
 sg13g2_decap_8 FILLER_76_371 ();
 sg13g2_decap_8 FILLER_76_378 ();
 sg13g2_decap_8 FILLER_76_385 ();
 sg13g2_decap_8 FILLER_76_392 ();
 sg13g2_decap_8 FILLER_76_399 ();
 sg13g2_fill_2 FILLER_76_406 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_fill_2 FILLER_77_140 ();
 sg13g2_fill_1 FILLER_77_142 ();
 sg13g2_fill_2 FILLER_77_146 ();
 sg13g2_fill_1 FILLER_77_175 ();
 sg13g2_fill_2 FILLER_77_190 ();
 sg13g2_fill_1 FILLER_77_192 ();
 sg13g2_fill_2 FILLER_77_219 ();
 sg13g2_fill_2 FILLER_77_247 ();
 sg13g2_decap_8 FILLER_77_284 ();
 sg13g2_decap_8 FILLER_77_291 ();
 sg13g2_decap_8 FILLER_77_298 ();
 sg13g2_decap_8 FILLER_77_305 ();
 sg13g2_decap_8 FILLER_77_312 ();
 sg13g2_decap_8 FILLER_77_319 ();
 sg13g2_decap_8 FILLER_77_326 ();
 sg13g2_decap_8 FILLER_77_333 ();
 sg13g2_decap_8 FILLER_77_340 ();
 sg13g2_decap_8 FILLER_77_347 ();
 sg13g2_decap_8 FILLER_77_354 ();
 sg13g2_decap_8 FILLER_77_361 ();
 sg13g2_decap_8 FILLER_77_368 ();
 sg13g2_decap_8 FILLER_77_375 ();
 sg13g2_decap_8 FILLER_77_382 ();
 sg13g2_decap_8 FILLER_77_389 ();
 sg13g2_decap_8 FILLER_77_396 ();
 sg13g2_decap_4 FILLER_77_403 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_4 FILLER_78_154 ();
 sg13g2_fill_1 FILLER_78_158 ();
 sg13g2_fill_1 FILLER_78_185 ();
 sg13g2_decap_8 FILLER_78_273 ();
 sg13g2_decap_8 FILLER_78_280 ();
 sg13g2_decap_8 FILLER_78_287 ();
 sg13g2_decap_8 FILLER_78_294 ();
 sg13g2_decap_8 FILLER_78_301 ();
 sg13g2_decap_8 FILLER_78_308 ();
 sg13g2_decap_8 FILLER_78_315 ();
 sg13g2_decap_8 FILLER_78_322 ();
 sg13g2_decap_8 FILLER_78_329 ();
 sg13g2_decap_8 FILLER_78_336 ();
 sg13g2_decap_8 FILLER_78_343 ();
 sg13g2_decap_8 FILLER_78_350 ();
 sg13g2_decap_8 FILLER_78_357 ();
 sg13g2_decap_8 FILLER_78_364 ();
 sg13g2_decap_8 FILLER_78_371 ();
 sg13g2_decap_8 FILLER_78_378 ();
 sg13g2_decap_8 FILLER_78_385 ();
 sg13g2_decap_8 FILLER_78_392 ();
 sg13g2_decap_8 FILLER_78_399 ();
 sg13g2_fill_2 FILLER_78_406 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_fill_1 FILLER_79_231 ();
 sg13g2_fill_2 FILLER_79_259 ();
 sg13g2_fill_1 FILLER_79_261 ();
 sg13g2_decap_8 FILLER_79_275 ();
 sg13g2_decap_8 FILLER_79_282 ();
 sg13g2_decap_8 FILLER_79_289 ();
 sg13g2_decap_4 FILLER_79_296 ();
 sg13g2_decap_8 FILLER_79_304 ();
 sg13g2_decap_8 FILLER_79_311 ();
 sg13g2_decap_8 FILLER_79_318 ();
 sg13g2_decap_8 FILLER_79_325 ();
 sg13g2_decap_8 FILLER_79_332 ();
 sg13g2_decap_8 FILLER_79_339 ();
 sg13g2_decap_8 FILLER_79_346 ();
 sg13g2_decap_8 FILLER_79_353 ();
 sg13g2_decap_8 FILLER_79_360 ();
 sg13g2_decap_8 FILLER_79_367 ();
 sg13g2_decap_8 FILLER_79_374 ();
 sg13g2_decap_8 FILLER_79_381 ();
 sg13g2_decap_8 FILLER_79_388 ();
 sg13g2_decap_8 FILLER_79_395 ();
 sg13g2_decap_8 FILLER_79_402 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_fill_2 FILLER_80_156 ();
 sg13g2_fill_1 FILLER_80_198 ();
 sg13g2_fill_2 FILLER_80_218 ();
 sg13g2_decap_8 FILLER_80_239 ();
 sg13g2_decap_4 FILLER_80_255 ();
 sg13g2_fill_1 FILLER_80_259 ();
 sg13g2_decap_8 FILLER_80_264 ();
 sg13g2_decap_8 FILLER_80_271 ();
 sg13g2_decap_8 FILLER_80_278 ();
 sg13g2_decap_8 FILLER_80_285 ();
 sg13g2_decap_8 FILLER_80_292 ();
 sg13g2_decap_8 FILLER_80_299 ();
 sg13g2_decap_8 FILLER_80_306 ();
 sg13g2_decap_8 FILLER_80_313 ();
 sg13g2_decap_8 FILLER_80_320 ();
 sg13g2_decap_8 FILLER_80_327 ();
 sg13g2_decap_8 FILLER_80_334 ();
 sg13g2_decap_8 FILLER_80_341 ();
 sg13g2_decap_8 FILLER_80_348 ();
 sg13g2_decap_8 FILLER_80_355 ();
 sg13g2_decap_8 FILLER_80_362 ();
 sg13g2_decap_8 FILLER_80_369 ();
 sg13g2_decap_8 FILLER_80_376 ();
 sg13g2_decap_8 FILLER_80_383 ();
 sg13g2_decap_8 FILLER_80_390 ();
 sg13g2_decap_8 FILLER_80_397 ();
 sg13g2_decap_4 FILLER_80_404 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net1;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net3;
 assign uio_oe[3] = net4;
 assign uio_oe[4] = net5;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net8;
 assign uio_out[0] = net9;
 assign uio_out[1] = net10;
 assign uio_out[2] = net11;
 assign uio_out[3] = net12;
 assign uio_out[4] = net13;
 assign uio_out[5] = net14;
 assign uio_out[6] = net15;
 assign uio_out[7] = net16;
endmodule

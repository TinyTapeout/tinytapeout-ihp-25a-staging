module tt_um_kailinsley (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire clknet_0_clk;
 wire \hidden_lif_0.spike_n ;
 wire \hidden_lif_0.state_r[0] ;
 wire \hidden_lif_0.state_r[1] ;
 wire \hidden_lif_0.state_r[2] ;
 wire \hidden_lif_0.state_r[3] ;
 wire \hidden_lif_0.state_r[4] ;
 wire \hidden_lif_0.state_r[5] ;
 wire \hidden_lif_0.state_r[6] ;
 wire \hidden_lif_0.state_r[7] ;
 wire \hidden_lif_0.variant_threshold[0] ;
 wire \hidden_lif_0.variant_threshold[1] ;
 wire \hidden_lif_0.variant_threshold[2] ;
 wire \hidden_lif_0.variant_threshold[3] ;
 wire \hidden_lif_0.variant_threshold[4] ;
 wire \hidden_lif_0.variant_threshold[5] ;
 wire \hidden_lif_0.variant_threshold[6] ;
 wire \hidden_lif_0.variant_threshold[7] ;
 wire \hidden_lif_1.spike_n ;
 wire \hidden_lif_1.state_r[0] ;
 wire \hidden_lif_1.state_r[1] ;
 wire \hidden_lif_1.state_r[2] ;
 wire \hidden_lif_1.state_r[3] ;
 wire \hidden_lif_1.state_r[4] ;
 wire \hidden_lif_1.state_r[5] ;
 wire \hidden_lif_1.state_r[6] ;
 wire \hidden_lif_1.state_r[7] ;
 wire \hidden_lif_1.variant_threshold[0] ;
 wire \hidden_lif_1.variant_threshold[1] ;
 wire \hidden_lif_1.variant_threshold[2] ;
 wire \hidden_lif_1.variant_threshold[3] ;
 wire \hidden_lif_1.variant_threshold[4] ;
 wire \hidden_lif_1.variant_threshold[5] ;
 wire \hidden_lif_1.variant_threshold[6] ;
 wire \hidden_lif_1.variant_threshold[7] ;
 wire \hidden_lif_2.spike_n ;
 wire \hidden_lif_2.state_r[0] ;
 wire \hidden_lif_2.state_r[1] ;
 wire \hidden_lif_2.state_r[2] ;
 wire \hidden_lif_2.state_r[3] ;
 wire \hidden_lif_2.state_r[4] ;
 wire \hidden_lif_2.state_r[5] ;
 wire \hidden_lif_2.state_r[6] ;
 wire \hidden_lif_2.state_r[7] ;
 wire \hidden_lif_2.variant_threshold[0] ;
 wire \hidden_lif_2.variant_threshold[1] ;
 wire \hidden_lif_2.variant_threshold[2] ;
 wire \hidden_lif_2.variant_threshold[3] ;
 wire \hidden_lif_2.variant_threshold[4] ;
 wire \hidden_lif_2.variant_threshold[5] ;
 wire \hidden_lif_2.variant_threshold[6] ;
 wire \hidden_lif_2.variant_threshold[7] ;
 wire \hidden_weight_0[0] ;
 wire \hidden_weight_0[1] ;
 wire \hidden_weight_0[2] ;
 wire \hidden_weight_1[0] ;
 wire \output_lif_0.spike_n ;
 wire \output_lif_0.state_r[0] ;
 wire \output_lif_0.state_r[1] ;
 wire \output_lif_0.state_r[2] ;
 wire \output_lif_0.state_r[3] ;
 wire \output_lif_0.state_r[4] ;
 wire \output_lif_0.state_r[5] ;
 wire \output_lif_0.state_r[6] ;
 wire \output_lif_0.state_r[7] ;
 wire \output_lif_0.variant_threshold[0] ;
 wire \output_lif_0.variant_threshold[1] ;
 wire \output_lif_0.variant_threshold[2] ;
 wire \output_lif_0.variant_threshold[3] ;
 wire \output_lif_0.variant_threshold[4] ;
 wire \output_lif_0.variant_threshold[5] ;
 wire \output_lif_0.variant_threshold[6] ;
 wire \output_lif_0.variant_threshold[7] ;
 wire \output_weight_0[0] ;
 wire \output_weight_0[1] ;
 wire \output_weight_0[2] ;
 wire \output_weight_1[0] ;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;

 sg13g2_inv_1 _0871_ (.Y(_0104_),
    .A(net166));
 sg13g2_inv_1 _0872_ (.Y(_0105_),
    .A(net101));
 sg13g2_inv_1 _0873_ (.Y(_0106_),
    .A(net220));
 sg13g2_inv_1 _0874_ (.Y(_0107_),
    .A(net136));
 sg13g2_inv_1 _0875_ (.Y(_0108_),
    .A(\hidden_lif_0.variant_threshold[0] ));
 sg13g2_inv_1 _0876_ (.Y(_0109_),
    .A(net143));
 sg13g2_inv_1 _0877_ (.Y(_0110_),
    .A(net210));
 sg13g2_inv_1 _0878_ (.Y(_0111_),
    .A(net227));
 sg13g2_inv_1 _0879_ (.Y(_0112_),
    .A(net230));
 sg13g2_inv_1 _0880_ (.Y(_0113_),
    .A(\hidden_lif_0.variant_threshold[4] ));
 sg13g2_inv_1 _0881_ (.Y(_0114_),
    .A(\hidden_lif_0.variant_threshold[3] ));
 sg13g2_inv_1 _0882_ (.Y(_0115_),
    .A(\hidden_lif_0.variant_threshold[2] ));
 sg13g2_inv_1 _0883_ (.Y(_0116_),
    .A(\hidden_lif_0.variant_threshold[1] ));
 sg13g2_inv_1 _0884_ (.Y(_0117_),
    .A(\hidden_lif_1.variant_threshold[0] ));
 sg13g2_inv_1 _0885_ (.Y(_0118_),
    .A(\output_lif_0.variant_threshold[7] ));
 sg13g2_inv_1 _0886_ (.Y(_0119_),
    .A(net236));
 sg13g2_inv_1 _0887_ (.Y(_0120_),
    .A(net237));
 sg13g2_inv_1 _0888_ (.Y(_0121_),
    .A(\output_lif_0.variant_threshold[4] ));
 sg13g2_inv_1 _0889_ (.Y(_0122_),
    .A(\output_lif_0.variant_threshold[3] ));
 sg13g2_inv_1 _0890_ (.Y(_0123_),
    .A(\output_lif_0.variant_threshold[2] ));
 sg13g2_inv_1 _0891_ (.Y(_0124_),
    .A(net173));
 sg13g2_inv_1 _0892_ (.Y(_0125_),
    .A(\hidden_lif_2.variant_threshold[6] ));
 sg13g2_inv_1 _0893_ (.Y(_0126_),
    .A(net234));
 sg13g2_inv_1 _0894_ (.Y(_0127_),
    .A(\hidden_lif_2.variant_threshold[4] ));
 sg13g2_inv_1 _0895_ (.Y(_0128_),
    .A(\hidden_lif_2.variant_threshold[3] ));
 sg13g2_inv_1 _0896_ (.Y(_0129_),
    .A(\hidden_lif_2.variant_threshold[2] ));
 sg13g2_inv_1 _0897_ (.Y(_0130_),
    .A(net213));
 sg13g2_inv_1 _0898_ (.Y(_0131_),
    .A(net191));
 sg13g2_inv_1 _0899_ (.Y(_0132_),
    .A(net97));
 sg13g2_inv_1 _0900_ (.Y(_0133_),
    .A(net103));
 sg13g2_inv_1 _0901_ (.Y(_0134_),
    .A(net197));
 sg13g2_inv_1 _0902_ (.Y(_0135_),
    .A(\hidden_lif_0.state_r[6] ));
 sg13g2_inv_1 _0903_ (.Y(_0136_),
    .A(\hidden_lif_0.state_r[5] ));
 sg13g2_inv_1 _0904_ (.Y(_0137_),
    .A(\hidden_lif_0.state_r[4] ));
 sg13g2_inv_1 _0905_ (.Y(_0138_),
    .A(\hidden_lif_0.state_r[3] ));
 sg13g2_inv_2 _0906_ (.Y(_0139_),
    .A(net106));
 sg13g2_inv_1 _0907_ (.Y(_0140_),
    .A(net190));
 sg13g2_inv_1 _0908_ (.Y(_0141_),
    .A(\hidden_lif_1.state_r[6] ));
 sg13g2_inv_1 _0909_ (.Y(_0142_),
    .A(\hidden_lif_1.state_r[5] ));
 sg13g2_inv_1 _0910_ (.Y(_0143_),
    .A(\hidden_lif_1.state_r[4] ));
 sg13g2_inv_2 _0911_ (.Y(_0144_),
    .A(\hidden_lif_1.state_r[3] ));
 sg13g2_inv_1 _0912_ (.Y(_0145_),
    .A(\hidden_lif_1.state_r[1] ));
 sg13g2_inv_1 _0913_ (.Y(_0146_),
    .A(net254));
 sg13g2_inv_1 _0914_ (.Y(_0147_),
    .A(net100));
 sg13g2_inv_1 _0915_ (.Y(_0148_),
    .A(net231));
 sg13g2_inv_1 _0916_ (.Y(_0149_),
    .A(\hidden_lif_2.state_r[6] ));
 sg13g2_inv_1 _0917_ (.Y(_0150_),
    .A(\hidden_lif_2.state_r[5] ));
 sg13g2_inv_1 _0918_ (.Y(_0151_),
    .A(\hidden_lif_2.state_r[4] ));
 sg13g2_inv_1 _0919_ (.Y(_0152_),
    .A(\hidden_lif_2.state_r[3] ));
 sg13g2_inv_1 _0920_ (.Y(_0153_),
    .A(\hidden_lif_2.state_r[2] ));
 sg13g2_inv_1 _0921_ (.Y(_0154_),
    .A(\output_lif_0.state_r[3] ));
 sg13g2_inv_1 _0922_ (.Y(_0155_),
    .A(\output_lif_0.state_r[2] ));
 sg13g2_inv_1 _0923_ (.Y(_0156_),
    .A(\output_lif_0.state_r[5] ));
 sg13g2_inv_1 _0924_ (.Y(_0157_),
    .A(\output_lif_0.state_r[4] ));
 sg13g2_inv_1 _0925_ (.Y(_0158_),
    .A(net239));
 sg13g2_inv_1 _0926_ (.Y(_0159_),
    .A(net92));
 sg13g2_inv_1 _0927_ (.Y(_0160_),
    .A(net158));
 sg13g2_inv_1 _0928_ (.Y(_0161_),
    .A(_0005_));
 sg13g2_inv_1 _0929_ (.Y(_0162_),
    .A(_0008_));
 sg13g2_inv_1 _0930_ (.Y(_0163_),
    .A(_0009_));
 sg13g2_inv_1 _0931_ (.Y(_0164_),
    .A(_0012_));
 sg13g2_inv_1 _0932_ (.Y(_0165_),
    .A(_0013_));
 sg13g2_inv_1 _0933_ (.Y(_0166_),
    .A(_0016_));
 sg13g2_or2_1 _0934_ (.X(_0167_),
    .B(\hidden_lif_1.variant_threshold[1] ),
    .A(\hidden_lif_1.variant_threshold[0] ));
 sg13g2_o21ai_1 _0935_ (.B1(\hidden_lif_1.variant_threshold[3] ),
    .Y(_0168_),
    .A1(\hidden_lif_1.variant_threshold[2] ),
    .A2(_0167_));
 sg13g2_nor4_1 _0936_ (.A(\hidden_lif_1.variant_threshold[7] ),
    .B(\hidden_lif_1.variant_threshold[6] ),
    .C(\hidden_lif_1.variant_threshold[5] ),
    .D(\hidden_lif_1.variant_threshold[4] ),
    .Y(_0169_));
 sg13g2_and2_1 _0937_ (.A(_0168_),
    .B(_0169_),
    .X(_0170_));
 sg13g2_and2_1 _0938_ (.A(net140),
    .B(_0170_),
    .X(_0171_));
 sg13g2_nand2_1 _0939_ (.Y(_0172_),
    .A(net140),
    .B(_0170_));
 sg13g2_a21oi_1 _0940_ (.A1(_0132_),
    .A2(_0167_),
    .Y(_0173_),
    .B1(_0171_));
 sg13g2_nor2_1 _0941_ (.A(net218),
    .B(_0173_),
    .Y(_0174_));
 sg13g2_nor2_1 _0942_ (.A(\hidden_lif_1.variant_threshold[0] ),
    .B(net97),
    .Y(_0175_));
 sg13g2_a22oi_1 _0943_ (.Y(_0176_),
    .B1(_0175_),
    .B2(net218),
    .A2(_0162_),
    .A1(net97));
 sg13g2_o21ai_1 _0944_ (.B1(net107),
    .Y(_0177_),
    .A1(_0171_),
    .A2(_0176_));
 sg13g2_nor2_1 _0945_ (.A(_0174_),
    .B(_0177_),
    .Y(_0020_));
 sg13g2_nand2b_1 _0946_ (.Y(_0178_),
    .B(net97),
    .A_N(net253));
 sg13g2_and3_1 _0947_ (.X(_0179_),
    .A(net212),
    .B(_0173_),
    .C(_0178_));
 sg13g2_a21oi_1 _0948_ (.A1(_0173_),
    .A2(_0178_),
    .Y(_0180_),
    .B1(net212));
 sg13g2_nor3_1 _0949_ (.A(net105),
    .B(_0179_),
    .C(_0180_),
    .Y(_0021_));
 sg13g2_nor3_2 _0950_ (.A(\hidden_lif_1.variant_threshold[3] ),
    .B(\hidden_lif_1.variant_threshold[2] ),
    .C(_0167_),
    .Y(_0181_));
 sg13g2_inv_1 _0951_ (.Y(_0182_),
    .A(_0181_));
 sg13g2_a21oi_1 _0952_ (.A1(_0168_),
    .A2(_0182_),
    .Y(_0183_),
    .B1(net98));
 sg13g2_nand3_1 _0953_ (.B(\hidden_lif_1.variant_threshold[2] ),
    .C(\hidden_lif_1.variant_threshold[1] ),
    .A(\hidden_lif_1.variant_threshold[3] ),
    .Y(_0184_));
 sg13g2_nand2_1 _0954_ (.Y(_0185_),
    .A(net97),
    .B(_0184_));
 sg13g2_nand4_1 _0955_ (.B(\hidden_lif_1.variant_threshold[1] ),
    .C(net98),
    .A(\hidden_lif_1.variant_threshold[2] ),
    .Y(_0186_),
    .D(_0184_));
 sg13g2_nor2b_1 _0956_ (.A(_0183_),
    .B_N(_0186_),
    .Y(_0187_));
 sg13g2_nand2_2 _0957_ (.Y(_0188_),
    .A(net107),
    .B(_0172_));
 sg13g2_nand2_1 _0958_ (.Y(_0189_),
    .A(_0172_),
    .B(_0185_));
 sg13g2_nand3_1 _0959_ (.B(net107),
    .C(_0189_),
    .A(net193),
    .Y(_0190_));
 sg13g2_o21ai_1 _0960_ (.B1(_0190_),
    .Y(_0022_),
    .A1(_0187_),
    .A2(_0188_));
 sg13g2_o21ai_1 _0961_ (.B1(_0185_),
    .Y(_0191_),
    .A1(net97),
    .A2(_0181_));
 sg13g2_xnor2_1 _0962_ (.Y(_0192_),
    .A(_0131_),
    .B(_0191_));
 sg13g2_o21ai_1 _0963_ (.B1(net107),
    .Y(_0023_),
    .A1(_0171_),
    .A2(_0192_));
 sg13g2_nor2_1 _0964_ (.A(_0131_),
    .B(_0184_),
    .Y(_0193_));
 sg13g2_nor2_1 _0965_ (.A(\hidden_lif_1.variant_threshold[4] ),
    .B(net97),
    .Y(_0194_));
 sg13g2_nand2_1 _0966_ (.Y(_0195_),
    .A(_0181_),
    .B(_0194_));
 sg13g2_a22oi_1 _0967_ (.Y(_0196_),
    .B1(_0194_),
    .B2(_0181_),
    .A2(_0193_),
    .A1(net97));
 sg13g2_xor2_1 _0968_ (.B(_0196_),
    .A(net214),
    .X(_0197_));
 sg13g2_nor2_1 _0969_ (.A(_0188_),
    .B(_0197_),
    .Y(_0024_));
 sg13g2_nand3_1 _0970_ (.B(net98),
    .C(_0193_),
    .A(\hidden_lif_1.variant_threshold[5] ),
    .Y(_0198_));
 sg13g2_nor2_1 _0971_ (.A(\hidden_lif_1.variant_threshold[5] ),
    .B(_0195_),
    .Y(_0199_));
 sg13g2_o21ai_1 _0972_ (.B1(_0198_),
    .Y(_0200_),
    .A1(\hidden_lif_1.variant_threshold[5] ),
    .A2(_0195_));
 sg13g2_xnor2_1 _0973_ (.Y(_0201_),
    .A(net195),
    .B(_0200_));
 sg13g2_nor2_1 _0974_ (.A(_0188_),
    .B(net196),
    .Y(_0025_));
 sg13g2_nand2_1 _0975_ (.Y(_0202_),
    .A(net195),
    .B(_0198_));
 sg13g2_o21ai_1 _0976_ (.B1(_0202_),
    .Y(_0203_),
    .A1(net195),
    .A2(_0199_));
 sg13g2_xnor2_1 _0977_ (.Y(_0204_),
    .A(_0130_),
    .B(_0203_));
 sg13g2_nor2_1 _0978_ (.A(_0188_),
    .B(_0204_),
    .Y(_0026_));
 sg13g2_or2_1 _0979_ (.X(_0205_),
    .B(\hidden_lif_2.variant_threshold[1] ),
    .A(\hidden_lif_2.variant_threshold[0] ));
 sg13g2_o21ai_1 _0980_ (.B1(\hidden_lif_2.variant_threshold[3] ),
    .Y(_0206_),
    .A1(\hidden_lif_2.variant_threshold[2] ),
    .A2(_0205_));
 sg13g2_nor4_1 _0981_ (.A(\hidden_lif_2.variant_threshold[7] ),
    .B(\hidden_lif_2.variant_threshold[6] ),
    .C(\hidden_lif_2.variant_threshold[5] ),
    .D(\hidden_lif_2.variant_threshold[4] ),
    .Y(_0207_));
 sg13g2_and2_1 _0982_ (.A(_0206_),
    .B(_0207_),
    .X(_0208_));
 sg13g2_nand2_2 _0983_ (.Y(_0209_),
    .A(net148),
    .B(_0208_));
 sg13g2_a22oi_1 _0984_ (.Y(_0210_),
    .B1(_0208_),
    .B2(net148),
    .A2(_0205_),
    .A1(_0133_));
 sg13g2_nor2_1 _0985_ (.A(net143),
    .B(net103),
    .Y(_0211_));
 sg13g2_a22oi_1 _0986_ (.Y(_0212_),
    .B1(_0211_),
    .B2(\hidden_lif_2.variant_threshold[1] ),
    .A2(_0164_),
    .A1(net103));
 sg13g2_inv_1 _0987_ (.Y(_0213_),
    .A(_0212_));
 sg13g2_o21ai_1 _0988_ (.B1(net106),
    .Y(_0214_),
    .A1(\hidden_lif_2.variant_threshold[1] ),
    .A2(_0210_));
 sg13g2_a21oi_1 _0989_ (.A1(_0209_),
    .A2(_0213_),
    .Y(_0027_),
    .B1(_0214_));
 sg13g2_nand2b_1 _0990_ (.Y(_0215_),
    .B(net103),
    .A_N(\hidden_lif_2.variant_threshold[1] ));
 sg13g2_and3_1 _0991_ (.X(_0216_),
    .A(net189),
    .B(_0210_),
    .C(_0215_));
 sg13g2_a21oi_1 _0992_ (.A1(_0210_),
    .A2(_0215_),
    .Y(_0217_),
    .B1(net189));
 sg13g2_nor3_1 _0993_ (.A(net105),
    .B(_0216_),
    .C(_0217_),
    .Y(_0028_));
 sg13g2_nor3_1 _0994_ (.A(\hidden_lif_2.variant_threshold[3] ),
    .B(\hidden_lif_2.variant_threshold[2] ),
    .C(_0205_),
    .Y(_0218_));
 sg13g2_inv_1 _0995_ (.Y(_0219_),
    .A(_0218_));
 sg13g2_a21oi_1 _0996_ (.A1(_0206_),
    .A2(_0219_),
    .Y(_0220_),
    .B1(net104));
 sg13g2_nand3_1 _0997_ (.B(\hidden_lif_2.variant_threshold[2] ),
    .C(\hidden_lif_2.variant_threshold[1] ),
    .A(\hidden_lif_2.variant_threshold[3] ),
    .Y(_0221_));
 sg13g2_nand2_1 _0998_ (.Y(_0222_),
    .A(net104),
    .B(_0221_));
 sg13g2_nand4_1 _0999_ (.B(\hidden_lif_2.variant_threshold[2] ),
    .C(\hidden_lif_2.variant_threshold[1] ),
    .A(_0128_),
    .Y(_0223_),
    .D(net104));
 sg13g2_nor2b_1 _1000_ (.A(_0220_),
    .B_N(_0223_),
    .Y(_0224_));
 sg13g2_nand2_2 _1001_ (.Y(_0225_),
    .A(net109),
    .B(_0209_));
 sg13g2_nand2_1 _1002_ (.Y(_0226_),
    .A(_0209_),
    .B(_0222_));
 sg13g2_nand3_1 _1003_ (.B(net106),
    .C(_0226_),
    .A(net185),
    .Y(_0227_));
 sg13g2_o21ai_1 _1004_ (.B1(_0227_),
    .Y(_0029_),
    .A1(_0224_),
    .A2(_0225_));
 sg13g2_nor2_1 _1005_ (.A(net104),
    .B(_0218_),
    .Y(_0228_));
 sg13g2_a21oi_1 _1006_ (.A1(net104),
    .A2(_0221_),
    .Y(_0229_),
    .B1(_0228_));
 sg13g2_and2_1 _1007_ (.A(net233),
    .B(_0229_),
    .X(_0230_));
 sg13g2_o21ai_1 _1008_ (.B1(_0209_),
    .Y(_0231_),
    .A1(net233),
    .A2(_0229_));
 sg13g2_o21ai_1 _1009_ (.B1(net109),
    .Y(_0030_),
    .A1(_0230_),
    .A2(_0231_));
 sg13g2_nor2_1 _1010_ (.A(_0127_),
    .B(_0221_),
    .Y(_0232_));
 sg13g2_nand2_1 _1011_ (.Y(_0233_),
    .A(_0127_),
    .B(_0218_));
 sg13g2_nor2_1 _1012_ (.A(net103),
    .B(_0233_),
    .Y(_0234_));
 sg13g2_a21oi_1 _1013_ (.A1(net103),
    .A2(_0232_),
    .Y(_0235_),
    .B1(_0234_));
 sg13g2_xnor2_1 _1014_ (.Y(_0236_),
    .A(_0126_),
    .B(_0235_));
 sg13g2_nor2_1 _1015_ (.A(_0225_),
    .B(_0236_),
    .Y(_0031_));
 sg13g2_nand3_1 _1016_ (.B(net103),
    .C(_0232_),
    .A(\hidden_lif_2.variant_threshold[5] ),
    .Y(_0237_));
 sg13g2_nand2_1 _1017_ (.Y(_0238_),
    .A(_0126_),
    .B(_0133_));
 sg13g2_a21oi_1 _1018_ (.A1(_0126_),
    .A2(_0234_),
    .Y(_0239_),
    .B1(\hidden_lif_2.variant_threshold[6] ));
 sg13g2_o21ai_1 _1019_ (.B1(_0237_),
    .Y(_0240_),
    .A1(_0233_),
    .A2(_0238_));
 sg13g2_xnor2_1 _1020_ (.Y(_0241_),
    .A(net200),
    .B(_0240_));
 sg13g2_nor2_1 _1021_ (.A(_0225_),
    .B(net201),
    .Y(_0032_));
 sg13g2_a21oi_1 _1022_ (.A1(\hidden_lif_2.variant_threshold[6] ),
    .A2(_0237_),
    .Y(_0242_),
    .B1(_0239_));
 sg13g2_xnor2_1 _1023_ (.Y(_0243_),
    .A(net173),
    .B(_0242_));
 sg13g2_nor2_1 _1024_ (.A(_0225_),
    .B(net174),
    .Y(_0033_));
 sg13g2_nor2_1 _1025_ (.A(\output_lif_0.variant_threshold[0] ),
    .B(\output_lif_0.variant_threshold[1] ),
    .Y(_0244_));
 sg13g2_nand2_1 _1026_ (.Y(_0245_),
    .A(_0123_),
    .B(_0244_));
 sg13g2_nand2_1 _1027_ (.Y(_0246_),
    .A(\output_lif_0.variant_threshold[3] ),
    .B(_0245_));
 sg13g2_nor4_1 _1028_ (.A(\output_lif_0.variant_threshold[7] ),
    .B(\output_lif_0.variant_threshold[6] ),
    .C(\output_lif_0.variant_threshold[5] ),
    .D(\output_lif_0.variant_threshold[4] ),
    .Y(_0247_));
 sg13g2_and2_1 _1029_ (.A(_0246_),
    .B(_0247_),
    .X(_0248_));
 sg13g2_and2_1 _1030_ (.A(net175),
    .B(_0248_),
    .X(_0249_));
 sg13g2_nand2_1 _1031_ (.Y(_0250_),
    .A(net175),
    .B(_0248_));
 sg13g2_nor2_1 _1032_ (.A(net101),
    .B(_0244_),
    .Y(_0251_));
 sg13g2_nor2_1 _1033_ (.A(_0249_),
    .B(_0251_),
    .Y(_0252_));
 sg13g2_nor2_1 _1034_ (.A(net101),
    .B(net188),
    .Y(_0253_));
 sg13g2_a22oi_1 _1035_ (.Y(_0254_),
    .B1(_0253_),
    .B2(\output_lif_0.variant_threshold[1] ),
    .A2(_0166_),
    .A1(net101));
 sg13g2_inv_1 _1036_ (.Y(_0255_),
    .A(_0254_));
 sg13g2_o21ai_1 _1037_ (.B1(net108),
    .Y(_0256_),
    .A1(\output_lif_0.variant_threshold[1] ),
    .A2(_0252_));
 sg13g2_a21oi_1 _1038_ (.A1(_0250_),
    .A2(_0255_),
    .Y(_0034_),
    .B1(_0256_));
 sg13g2_nand2b_1 _1039_ (.Y(_0257_),
    .B(net102),
    .A_N(\output_lif_0.variant_threshold[1] ));
 sg13g2_and3_1 _1040_ (.X(_0258_),
    .A(net171),
    .B(_0252_),
    .C(_0257_));
 sg13g2_a21oi_1 _1041_ (.A1(_0252_),
    .A2(_0257_),
    .Y(_0259_),
    .B1(net171));
 sg13g2_nor3_1 _1042_ (.A(net105),
    .B(_0258_),
    .C(net172),
    .Y(_0035_));
 sg13g2_nand2_2 _1043_ (.Y(_0260_),
    .A(net108),
    .B(_0250_));
 sg13g2_nor2_1 _1044_ (.A(net101),
    .B(_0246_),
    .Y(_0261_));
 sg13g2_nand3_1 _1045_ (.B(\output_lif_0.variant_threshold[2] ),
    .C(\output_lif_0.variant_threshold[1] ),
    .A(\output_lif_0.variant_threshold[3] ),
    .Y(_0262_));
 sg13g2_and4_1 _1046_ (.A(net101),
    .B(_0122_),
    .C(\output_lif_0.variant_threshold[2] ),
    .D(\output_lif_0.variant_threshold[1] ),
    .X(_0263_));
 sg13g2_nor3_2 _1047_ (.A(net101),
    .B(\output_lif_0.variant_threshold[3] ),
    .C(_0245_),
    .Y(_0264_));
 sg13g2_nor3_1 _1048_ (.A(_0261_),
    .B(_0263_),
    .C(_0264_),
    .Y(_0265_));
 sg13g2_a21o_1 _1049_ (.A2(_0262_),
    .A1(net101),
    .B1(_0249_),
    .X(_0266_));
 sg13g2_nand3_1 _1050_ (.B(net108),
    .C(_0266_),
    .A(net186),
    .Y(_0267_));
 sg13g2_o21ai_1 _1051_ (.B1(_0267_),
    .Y(_0036_),
    .A1(_0260_),
    .A2(_0265_));
 sg13g2_nor2_1 _1052_ (.A(_0105_),
    .B(_0262_),
    .Y(_0268_));
 sg13g2_nor3_1 _1053_ (.A(net243),
    .B(_0264_),
    .C(_0268_),
    .Y(_0269_));
 sg13g2_o21ai_1 _1054_ (.B1(net243),
    .Y(_0270_),
    .A1(_0264_),
    .A2(_0268_));
 sg13g2_nand2_1 _1055_ (.Y(_0271_),
    .A(_0250_),
    .B(_0270_));
 sg13g2_o21ai_1 _1056_ (.B1(net108),
    .Y(_0037_),
    .A1(_0269_),
    .A2(_0271_));
 sg13g2_and2_1 _1057_ (.A(_0121_),
    .B(_0264_),
    .X(_0272_));
 sg13g2_a21oi_1 _1058_ (.A1(\output_lif_0.variant_threshold[4] ),
    .A2(_0268_),
    .Y(_0273_),
    .B1(_0272_));
 sg13g2_xnor2_1 _1059_ (.Y(_0274_),
    .A(_0120_),
    .B(_0273_));
 sg13g2_nor2_1 _1060_ (.A(_0260_),
    .B(net238),
    .Y(_0038_));
 sg13g2_nor4_1 _1061_ (.A(_0105_),
    .B(_0120_),
    .C(_0121_),
    .D(_0262_),
    .Y(_0275_));
 sg13g2_and2_1 _1062_ (.A(_0120_),
    .B(_0272_),
    .X(_0276_));
 sg13g2_nor2_1 _1063_ (.A(_0275_),
    .B(_0276_),
    .Y(_0277_));
 sg13g2_xnor2_1 _1064_ (.Y(_0278_),
    .A(_0119_),
    .B(_0277_));
 sg13g2_nor2_1 _1065_ (.A(_0260_),
    .B(_0278_),
    .Y(_0039_));
 sg13g2_mux2_1 _1066_ (.A0(_0275_),
    .A1(_0276_),
    .S(_0119_),
    .X(_0279_));
 sg13g2_xnor2_1 _1067_ (.Y(_0280_),
    .A(net179),
    .B(_0279_));
 sg13g2_nor2_1 _1068_ (.A(_0260_),
    .B(_0280_),
    .Y(_0040_));
 sg13g2_nand2b_1 _1069_ (.Y(_0281_),
    .B(\hidden_lif_2.state_r[1] ),
    .A_N(\hidden_lif_2.variant_threshold[1] ));
 sg13g2_nand3b_1 _1070_ (.B(_0281_),
    .C(\hidden_lif_2.variant_threshold[0] ),
    .Y(_0282_),
    .A_N(\hidden_lif_2.state_r[0] ));
 sg13g2_nand2b_1 _1071_ (.Y(_0283_),
    .B(\hidden_lif_2.variant_threshold[1] ),
    .A_N(\hidden_lif_2.state_r[1] ));
 sg13g2_a22oi_1 _1072_ (.Y(_0284_),
    .B1(_0282_),
    .B2(_0283_),
    .A2(\hidden_lif_2.state_r[2] ),
    .A1(_0129_));
 sg13g2_a221oi_1 _1073_ (.B2(\hidden_lif_2.variant_threshold[2] ),
    .C1(_0284_),
    .B1(_0153_),
    .A1(\hidden_lif_2.variant_threshold[3] ),
    .Y(_0285_),
    .A2(_0152_));
 sg13g2_a221oi_1 _1074_ (.B2(_0128_),
    .C1(_0285_),
    .B1(\hidden_lif_2.state_r[3] ),
    .A1(_0127_),
    .Y(_0286_),
    .A2(\hidden_lif_2.state_r[4] ));
 sg13g2_a221oi_1 _1075_ (.B2(\hidden_lif_2.variant_threshold[4] ),
    .C1(_0286_),
    .B1(_0151_),
    .A1(\hidden_lif_2.variant_threshold[5] ),
    .Y(_0287_),
    .A2(_0150_));
 sg13g2_a221oi_1 _1076_ (.B2(_0126_),
    .C1(_0287_),
    .B1(\hidden_lif_2.state_r[5] ),
    .A1(_0125_),
    .Y(_0288_),
    .A2(\hidden_lif_2.state_r[6] ));
 sg13g2_a221oi_1 _1077_ (.B2(\hidden_lif_2.variant_threshold[6] ),
    .C1(_0288_),
    .B1(_0149_),
    .A1(net173),
    .Y(_0289_),
    .A2(_0148_));
 sg13g2_a21oi_2 _1078_ (.B1(_0289_),
    .Y(_0290_),
    .A2(net231),
    .A1(_0124_));
 sg13g2_nor2_1 _1079_ (.A(net105),
    .B(_0290_),
    .Y(_0041_));
 sg13g2_nand2b_1 _1080_ (.Y(_0291_),
    .B(\output_lif_0.state_r[1] ),
    .A_N(\output_lif_0.variant_threshold[1] ));
 sg13g2_nor2b_1 _1081_ (.A(\output_lif_0.state_r[0] ),
    .B_N(\output_lif_0.variant_threshold[0] ),
    .Y(_0292_));
 sg13g2_nor2b_1 _1082_ (.A(\output_lif_0.state_r[1] ),
    .B_N(\output_lif_0.variant_threshold[1] ),
    .Y(_0293_));
 sg13g2_a221oi_1 _1083_ (.B2(_0292_),
    .C1(_0293_),
    .B1(_0291_),
    .A1(\output_lif_0.variant_threshold[2] ),
    .Y(_0294_),
    .A2(_0155_));
 sg13g2_a221oi_1 _1084_ (.B2(_0123_),
    .C1(_0294_),
    .B1(\output_lif_0.state_r[2] ),
    .A1(_0122_),
    .Y(_0295_),
    .A2(\output_lif_0.state_r[3] ));
 sg13g2_a221oi_1 _1085_ (.B2(\output_lif_0.variant_threshold[4] ),
    .C1(_0295_),
    .B1(_0157_),
    .A1(\output_lif_0.variant_threshold[3] ),
    .Y(_0296_),
    .A2(_0154_));
 sg13g2_a221oi_1 _1086_ (.B2(_0121_),
    .C1(_0296_),
    .B1(\output_lif_0.state_r[4] ),
    .A1(_0120_),
    .Y(_0297_),
    .A2(\output_lif_0.state_r[5] ));
 sg13g2_a221oi_1 _1087_ (.B2(\output_lif_0.variant_threshold[6] ),
    .C1(_0297_),
    .B1(_0159_),
    .A1(\output_lif_0.variant_threshold[5] ),
    .Y(_0298_),
    .A2(_0156_));
 sg13g2_a221oi_1 _1088_ (.B2(_0119_),
    .C1(_0298_),
    .B1(net92),
    .A1(_0118_),
    .Y(_0299_),
    .A2(net239));
 sg13g2_a21oi_1 _1089_ (.A1(net179),
    .A2(_0158_),
    .Y(_0300_),
    .B1(net240));
 sg13g2_and2_1 _1090_ (.A(net108),
    .B(_0300_),
    .X(_0042_));
 sg13g2_nand2b_1 _1091_ (.Y(_0301_),
    .B(net140),
    .A_N(_0170_));
 sg13g2_o21ai_1 _1092_ (.B1(net107),
    .Y(_0302_),
    .A1(_0175_),
    .A2(_0301_));
 sg13g2_a21oi_1 _1093_ (.A1(_0117_),
    .A2(_0301_),
    .Y(_0043_),
    .B1(_0302_));
 sg13g2_xnor2_1 _1094_ (.Y(_0303_),
    .A(net7),
    .B(net8));
 sg13g2_and2_1 _1095_ (.A(net1),
    .B(net2),
    .X(_0304_));
 sg13g2_or2_1 _1096_ (.X(_0305_),
    .B(net2),
    .A(net1));
 sg13g2_xnor2_1 _1097_ (.Y(_0306_),
    .A(net1),
    .B(net2));
 sg13g2_xnor2_1 _1098_ (.Y(_0307_),
    .A(net3),
    .B(_0306_));
 sg13g2_or2_1 _1099_ (.X(_0308_),
    .B(net5),
    .A(net4));
 sg13g2_a21o_1 _1100_ (.A2(net5),
    .A1(net4),
    .B1(net6),
    .X(_0309_));
 sg13g2_and2_1 _1101_ (.A(_0308_),
    .B(_0309_),
    .X(_0310_));
 sg13g2_xnor2_1 _1102_ (.Y(_0311_),
    .A(net4),
    .B(net5));
 sg13g2_xnor2_1 _1103_ (.Y(_0312_),
    .A(net6),
    .B(_0311_));
 sg13g2_xnor2_1 _1104_ (.Y(_0313_),
    .A(_0307_),
    .B(_0312_));
 sg13g2_nor2_1 _1105_ (.A(_0303_),
    .B(_0313_),
    .Y(_0314_));
 sg13g2_xor2_1 _1106_ (.B(_0313_),
    .A(_0303_),
    .X(_0315_));
 sg13g2_and2_2 _1107_ (.A(net96),
    .B(_0315_),
    .X(_0316_));
 sg13g2_and2_1 _1108_ (.A(net96),
    .B(_0314_),
    .X(_0317_));
 sg13g2_and2_1 _1109_ (.A(net8),
    .B(\hidden_weight_0[1] ),
    .X(_0318_));
 sg13g2_nand2_1 _1110_ (.Y(_0319_),
    .A(net7),
    .B(\hidden_weight_0[1] ));
 sg13g2_nand3_1 _1111_ (.B(_0308_),
    .C(_0309_),
    .A(net95),
    .Y(_0320_));
 sg13g2_nand2_1 _1112_ (.Y(_0321_),
    .A(net95),
    .B(net7));
 sg13g2_xor2_1 _1113_ (.B(_0320_),
    .A(_0319_),
    .X(_0322_));
 sg13g2_nand2_1 _1114_ (.Y(_0323_),
    .A(_0318_),
    .B(_0322_));
 sg13g2_xor2_1 _1115_ (.B(_0322_),
    .A(_0318_),
    .X(_0324_));
 sg13g2_inv_1 _1116_ (.Y(_0325_),
    .A(_0324_));
 sg13g2_nand2_1 _1117_ (.Y(_0326_),
    .A(net94),
    .B(_0312_));
 sg13g2_and2_1 _1118_ (.A(net94),
    .B(_0307_),
    .X(_0327_));
 sg13g2_nand2_1 _1119_ (.Y(_0328_),
    .A(\hidden_weight_0[1] ),
    .B(_0312_));
 sg13g2_a21o_2 _1120_ (.A2(_0305_),
    .A1(net3),
    .B1(_0304_),
    .X(_0329_));
 sg13g2_and4_1 _1121_ (.A(net95),
    .B(net3),
    .C(\hidden_weight_0[1] ),
    .D(_0304_),
    .X(_0330_));
 sg13g2_a22oi_1 _1122_ (.Y(_0331_),
    .B1(_0329_),
    .B2(net94),
    .A2(_0307_),
    .A1(\hidden_weight_0[1] ));
 sg13g2_or3_1 _1123_ (.A(_0328_),
    .B(_0330_),
    .C(_0331_),
    .X(_0332_));
 sg13g2_o21ai_1 _1124_ (.B1(_0328_),
    .Y(_0333_),
    .A1(_0330_),
    .A2(_0331_));
 sg13g2_nand2_1 _1125_ (.Y(_0334_),
    .A(_0332_),
    .B(_0333_));
 sg13g2_and4_1 _1126_ (.A(net94),
    .B(_0307_),
    .C(_0312_),
    .D(_0329_),
    .X(_0335_));
 sg13g2_nand4_1 _1127_ (.B(_0307_),
    .C(_0312_),
    .A(net94),
    .Y(_0336_),
    .D(_0329_));
 sg13g2_a22oi_1 _1128_ (.Y(_0337_),
    .B1(_0332_),
    .B2(_0333_),
    .A2(_0327_),
    .A1(_0312_));
 sg13g2_nand3b_1 _1129_ (.B(_0324_),
    .C(_0336_),
    .Y(_0338_),
    .A_N(_0337_));
 sg13g2_o21ai_1 _1130_ (.B1(_0325_),
    .Y(_0339_),
    .A1(_0335_),
    .A2(_0337_));
 sg13g2_and3_1 _1131_ (.X(_0340_),
    .A(_0317_),
    .B(_0338_),
    .C(_0339_));
 sg13g2_nand3_1 _1132_ (.B(_0338_),
    .C(_0339_),
    .A(_0317_),
    .Y(_0341_));
 sg13g2_nand2_1 _1133_ (.Y(_0342_),
    .A(net95),
    .B(net8));
 sg13g2_and3_2 _1134_ (.X(_0343_),
    .A(net96),
    .B(net7),
    .C(net8));
 sg13g2_a21o_2 _1135_ (.A2(_0339_),
    .A1(_0338_),
    .B1(_0317_),
    .X(_0344_));
 sg13g2_and3_1 _1136_ (.X(_0345_),
    .A(_0341_),
    .B(_0343_),
    .C(_0344_));
 sg13g2_nand3_1 _1137_ (.B(_0343_),
    .C(_0344_),
    .A(_0341_),
    .Y(_0346_));
 sg13g2_a21oi_1 _1138_ (.A1(_0343_),
    .A2(_0344_),
    .Y(_0347_),
    .B1(_0340_));
 sg13g2_nand2_1 _1139_ (.Y(_0348_),
    .A(_0336_),
    .B(_0338_));
 sg13g2_nand2_1 _1140_ (.Y(_0349_),
    .A(\hidden_weight_0[2] ),
    .B(_0315_));
 sg13g2_o21ai_1 _1141_ (.B1(\hidden_weight_0[1] ),
    .Y(_0350_),
    .A1(_0310_),
    .A2(_0329_));
 sg13g2_a21oi_1 _1142_ (.A1(_0310_),
    .A2(_0329_),
    .Y(_0351_),
    .B1(_0350_));
 sg13g2_xnor2_1 _1143_ (.Y(_0352_),
    .A(_0349_),
    .B(_0351_));
 sg13g2_o21ai_1 _1144_ (.B1(_0323_),
    .Y(_0353_),
    .A1(_0319_),
    .A2(_0320_));
 sg13g2_nor2b_1 _1145_ (.A(_0330_),
    .B_N(_0332_),
    .Y(_0354_));
 sg13g2_xor2_1 _1146_ (.B(_0354_),
    .A(_0353_),
    .X(_0355_));
 sg13g2_xnor2_1 _1147_ (.Y(_0356_),
    .A(_0352_),
    .B(_0355_));
 sg13g2_xnor2_1 _1148_ (.Y(_0357_),
    .A(_0348_),
    .B(_0356_));
 sg13g2_xnor2_1 _1149_ (.Y(_0358_),
    .A(_0347_),
    .B(_0357_));
 sg13g2_a21oi_2 _1150_ (.B1(_0343_),
    .Y(_0359_),
    .A2(_0344_),
    .A1(_0341_));
 sg13g2_a21o_1 _1151_ (.A2(_0344_),
    .A1(_0341_),
    .B1(_0343_),
    .X(_0360_));
 sg13g2_o21ai_1 _1152_ (.B1(_0358_),
    .Y(_0361_),
    .A1(_0345_),
    .A2(_0359_));
 sg13g2_nor2_1 _1153_ (.A(_0316_),
    .B(_0361_),
    .Y(_0362_));
 sg13g2_or2_2 _1154_ (.X(_0363_),
    .B(_0361_),
    .A(_0316_));
 sg13g2_nor2_1 _1155_ (.A(_0138_),
    .B(\hidden_lif_0.state_r[0] ),
    .Y(_0364_));
 sg13g2_xnor2_1 _1156_ (.Y(_0365_),
    .A(\hidden_lif_0.state_r[3] ),
    .B(net207));
 sg13g2_nor2_1 _1157_ (.A(\hidden_lif_0.state_r[1] ),
    .B(_0316_),
    .Y(_0366_));
 sg13g2_nand2b_1 _1158_ (.Y(_0367_),
    .B(\hidden_lif_0.variant_threshold[1] ),
    .A_N(\hidden_lif_0.state_r[1] ));
 sg13g2_o21ai_1 _1159_ (.B1(_0367_),
    .Y(_0368_),
    .A1(_0108_),
    .A2(\hidden_lif_0.state_r[0] ));
 sg13g2_a22oi_1 _1160_ (.Y(_0369_),
    .B1(\hidden_lif_0.state_r[1] ),
    .B2(_0116_),
    .A2(\hidden_lif_0.state_r[2] ),
    .A1(_0115_));
 sg13g2_nor2_1 _1161_ (.A(_0115_),
    .B(\hidden_lif_0.state_r[2] ),
    .Y(_0370_));
 sg13g2_a221oi_1 _1162_ (.B2(_0369_),
    .C1(_0370_),
    .B1(_0368_),
    .A1(\hidden_lif_0.variant_threshold[3] ),
    .Y(_0371_),
    .A2(_0138_));
 sg13g2_a221oi_1 _1163_ (.B2(_0114_),
    .C1(_0371_),
    .B1(\hidden_lif_0.state_r[3] ),
    .A1(_0113_),
    .Y(_0372_),
    .A2(\hidden_lif_0.state_r[4] ));
 sg13g2_a221oi_1 _1164_ (.B2(\hidden_lif_0.variant_threshold[4] ),
    .C1(_0372_),
    .B1(_0137_),
    .A1(\hidden_lif_0.variant_threshold[5] ),
    .Y(_0373_),
    .A2(_0136_));
 sg13g2_a221oi_1 _1165_ (.B2(_0112_),
    .C1(_0373_),
    .B1(\hidden_lif_0.state_r[5] ),
    .A1(_0111_),
    .Y(_0374_),
    .A2(\hidden_lif_0.state_r[6] ));
 sg13g2_a221oi_1 _1166_ (.B2(\hidden_lif_0.variant_threshold[6] ),
    .C1(_0374_),
    .B1(_0135_),
    .A1(net210),
    .Y(_0375_),
    .A2(_0134_));
 sg13g2_a21oi_2 _1167_ (.B1(_0375_),
    .Y(_0376_),
    .A2(net197),
    .A1(_0110_));
 sg13g2_nand2_2 _1168_ (.Y(_0377_),
    .A(net110),
    .B(_0376_));
 sg13g2_nand2_1 _1169_ (.Y(_0378_),
    .A(net252),
    .B(_0316_));
 sg13g2_nand3_1 _1170_ (.B(_0376_),
    .C(_0378_),
    .A(net110),
    .Y(_0379_));
 sg13g2_a221oi_1 _1171_ (.B2(_0361_),
    .C1(_0379_),
    .B1(_0366_),
    .A1(net87),
    .Y(_0044_),
    .A2(net208));
 sg13g2_nor3_2 _1172_ (.A(_0005_),
    .B(_0345_),
    .C(_0359_),
    .Y(_0380_));
 sg13g2_a21oi_1 _1173_ (.A1(_0346_),
    .A2(_0360_),
    .Y(_0381_),
    .B1(_0161_));
 sg13g2_nor3_1 _1174_ (.A(_0378_),
    .B(_0380_),
    .C(_0381_),
    .Y(_0382_));
 sg13g2_or3_1 _1175_ (.A(net87),
    .B(_0380_),
    .C(_0381_),
    .X(_0383_));
 sg13g2_a21oi_1 _1176_ (.A1(_0378_),
    .A2(_0383_),
    .Y(_0384_),
    .B1(_0382_));
 sg13g2_nor2b_1 _1177_ (.A(\hidden_lif_0.state_r[4] ),
    .B_N(\hidden_lif_0.state_r[1] ),
    .Y(_0385_));
 sg13g2_xor2_1 _1178_ (.B(\hidden_lif_0.state_r[1] ),
    .A(\hidden_lif_0.state_r[4] ),
    .X(_0386_));
 sg13g2_nor2_1 _1179_ (.A(_0364_),
    .B(_0386_),
    .Y(_0387_));
 sg13g2_xor2_1 _1180_ (.B(_0386_),
    .A(_0364_),
    .X(_0388_));
 sg13g2_a21oi_1 _1181_ (.A1(net86),
    .A2(_0388_),
    .Y(_0389_),
    .B1(_0384_));
 sg13g2_nor2_1 _1182_ (.A(_0377_),
    .B(_0389_),
    .Y(_0045_));
 sg13g2_nand2b_1 _1183_ (.Y(_0390_),
    .B(\hidden_lif_0.state_r[3] ),
    .A_N(_0358_));
 sg13g2_xnor2_1 _1184_ (.Y(_0391_),
    .A(\hidden_lif_0.state_r[3] ),
    .B(_0358_));
 sg13g2_o21ai_1 _1185_ (.B1(_0391_),
    .Y(_0392_),
    .A1(_0380_),
    .A2(_0382_));
 sg13g2_or3_1 _1186_ (.A(_0380_),
    .B(_0382_),
    .C(_0391_),
    .X(_0393_));
 sg13g2_nand2_1 _1187_ (.Y(_0394_),
    .A(_0136_),
    .B(\hidden_lif_0.state_r[2] ));
 sg13g2_xnor2_1 _1188_ (.Y(_0395_),
    .A(\hidden_lif_0.state_r[5] ),
    .B(\hidden_lif_0.state_r[2] ));
 sg13g2_o21ai_1 _1189_ (.B1(_0395_),
    .Y(_0396_),
    .A1(_0385_),
    .A2(_0387_));
 sg13g2_or3_1 _1190_ (.A(_0385_),
    .B(_0387_),
    .C(_0395_),
    .X(_0397_));
 sg13g2_a21oi_1 _1191_ (.A1(_0396_),
    .A2(_0397_),
    .Y(_0398_),
    .B1(_0363_));
 sg13g2_a21oi_1 _1192_ (.A1(_0392_),
    .A2(_0393_),
    .Y(_0399_),
    .B1(net87));
 sg13g2_nor3_1 _1193_ (.A(_0377_),
    .B(_0398_),
    .C(_0399_),
    .Y(_0046_));
 sg13g2_nor2_1 _1194_ (.A(\hidden_lif_0.state_r[6] ),
    .B(_0138_),
    .Y(_0400_));
 sg13g2_xor2_1 _1195_ (.B(\hidden_lif_0.state_r[3] ),
    .A(\hidden_lif_0.state_r[6] ),
    .X(_0401_));
 sg13g2_and3_1 _1196_ (.X(_0402_),
    .A(_0394_),
    .B(_0396_),
    .C(_0401_));
 sg13g2_a21oi_2 _1197_ (.B1(_0401_),
    .Y(_0403_),
    .A2(_0396_),
    .A1(_0394_));
 sg13g2_nor2_1 _1198_ (.A(_0402_),
    .B(_0403_),
    .Y(_0404_));
 sg13g2_nand3_1 _1199_ (.B(_0390_),
    .C(_0392_),
    .A(net192),
    .Y(_0405_));
 sg13g2_a21oi_2 _1200_ (.B1(net192),
    .Y(_0406_),
    .A2(_0392_),
    .A1(_0390_));
 sg13g2_nor2_1 _1201_ (.A(net86),
    .B(_0406_),
    .Y(_0407_));
 sg13g2_a22oi_1 _1202_ (.Y(_0408_),
    .B1(_0405_),
    .B2(_0407_),
    .A2(_0404_),
    .A1(net86));
 sg13g2_nor2_1 _1203_ (.A(_0377_),
    .B(_0408_),
    .Y(_0047_));
 sg13g2_nand2_1 _1204_ (.Y(_0409_),
    .A(_0134_),
    .B(\hidden_lif_0.state_r[4] ));
 sg13g2_xnor2_1 _1205_ (.Y(_0410_),
    .A(\hidden_lif_0.state_r[7] ),
    .B(\hidden_lif_0.state_r[4] ));
 sg13g2_nor3_1 _1206_ (.A(_0400_),
    .B(_0403_),
    .C(_0410_),
    .Y(_0411_));
 sg13g2_o21ai_1 _1207_ (.B1(_0410_),
    .Y(_0412_),
    .A1(_0400_),
    .A2(_0403_));
 sg13g2_nand2b_1 _1208_ (.Y(_0413_),
    .B(_0412_),
    .A_N(_0411_));
 sg13g2_xor2_1 _1209_ (.B(_0406_),
    .A(net161),
    .X(_0414_));
 sg13g2_a21o_1 _1210_ (.A2(_0413_),
    .A1(net86),
    .B1(_0377_),
    .X(_0415_));
 sg13g2_a21oi_1 _1211_ (.A1(_0363_),
    .A2(net162),
    .Y(_0048_),
    .B1(_0415_));
 sg13g2_a21o_1 _1212_ (.A2(_0406_),
    .A1(net250),
    .B1(\hidden_lif_0.state_r[6] ),
    .X(_0416_));
 sg13g2_nor2_1 _1213_ (.A(_0135_),
    .B(_0136_),
    .Y(_0417_));
 sg13g2_a21oi_1 _1214_ (.A1(_0406_),
    .A2(_0417_),
    .Y(_0418_),
    .B1(net86));
 sg13g2_nand2_1 _1215_ (.Y(_0419_),
    .A(_0409_),
    .B(_0412_));
 sg13g2_xnor2_1 _1216_ (.Y(_0420_),
    .A(net250),
    .B(_0419_));
 sg13g2_a22oi_1 _1217_ (.Y(_0421_),
    .B1(_0420_),
    .B2(net86),
    .A2(_0418_),
    .A1(_0416_));
 sg13g2_nor2_1 _1218_ (.A(_0377_),
    .B(net251),
    .Y(_0049_));
 sg13g2_nand3_1 _1219_ (.B(_0406_),
    .C(_0417_),
    .A(_0134_),
    .Y(_0422_));
 sg13g2_a21oi_1 _1220_ (.A1(_0406_),
    .A2(_0417_),
    .Y(_0423_),
    .B1(_0134_));
 sg13g2_nor2_1 _1221_ (.A(net86),
    .B(_0423_),
    .Y(_0424_));
 sg13g2_and2_1 _1222_ (.A(net161),
    .B(_0409_),
    .X(_0425_));
 sg13g2_o21ai_1 _1223_ (.B1(_0425_),
    .Y(_0426_),
    .A1(\hidden_lif_0.state_r[5] ),
    .A2(_0412_));
 sg13g2_nor2_1 _1224_ (.A(\hidden_lif_0.state_r[6] ),
    .B(_0426_),
    .Y(_0427_));
 sg13g2_xnor2_1 _1225_ (.Y(_0428_),
    .A(_0135_),
    .B(_0426_));
 sg13g2_a221oi_1 _1226_ (.B2(net86),
    .C1(_0377_),
    .B1(_0428_),
    .A1(_0422_),
    .Y(_0050_),
    .A2(_0424_));
 sg13g2_xnor2_1 _1227_ (.Y(_0429_),
    .A(net197),
    .B(_0427_));
 sg13g2_nor3_1 _1228_ (.A(_0377_),
    .B(_0418_),
    .C(net198),
    .Y(_0051_));
 sg13g2_nor2_1 _1229_ (.A(_0139_),
    .B(net211),
    .Y(_0052_));
 sg13g2_or2_1 _1230_ (.X(_0430_),
    .B(\hidden_lif_0.variant_threshold[1] ),
    .A(\hidden_lif_0.variant_threshold[0] ));
 sg13g2_o21ai_1 _1231_ (.B1(\hidden_lif_0.variant_threshold[3] ),
    .Y(_0431_),
    .A1(\hidden_lif_0.variant_threshold[2] ),
    .A2(_0430_));
 sg13g2_nor2_1 _1232_ (.A(net228),
    .B(\hidden_lif_0.variant_threshold[5] ),
    .Y(_0432_));
 sg13g2_and4_1 _1233_ (.A(_0110_),
    .B(_0113_),
    .C(_0431_),
    .D(_0432_),
    .X(_0433_));
 sg13g2_nand2_2 _1234_ (.Y(_0434_),
    .A(net156),
    .B(_0433_));
 sg13g2_a22oi_1 _1235_ (.Y(_0435_),
    .B1(_0433_),
    .B2(net156),
    .A2(_0430_),
    .A1(_0147_));
 sg13g2_nor2_1 _1236_ (.A(\hidden_lif_0.variant_threshold[0] ),
    .B(net99),
    .Y(_0436_));
 sg13g2_a22oi_1 _1237_ (.Y(_0437_),
    .B1(_0436_),
    .B2(\hidden_lif_0.variant_threshold[1] ),
    .A2(_0160_),
    .A1(net99));
 sg13g2_inv_1 _1238_ (.Y(_0438_),
    .A(net159));
 sg13g2_o21ai_1 _1239_ (.B1(net111),
    .Y(_0439_),
    .A1(\hidden_lif_0.variant_threshold[1] ),
    .A2(_0435_));
 sg13g2_a21oi_1 _1240_ (.A1(_0434_),
    .A2(_0438_),
    .Y(_0053_),
    .B1(_0439_));
 sg13g2_nand2b_1 _1241_ (.Y(_0440_),
    .B(net99),
    .A_N(\hidden_lif_0.variant_threshold[1] ));
 sg13g2_and3_1 _1242_ (.X(_0441_),
    .A(net165),
    .B(_0435_),
    .C(_0440_));
 sg13g2_a21oi_1 _1243_ (.A1(_0435_),
    .A2(_0440_),
    .Y(_0442_),
    .B1(net165));
 sg13g2_nor3_1 _1244_ (.A(_0139_),
    .B(_0441_),
    .C(_0442_),
    .Y(_0054_));
 sg13g2_nand3b_1 _1245_ (.B(_0115_),
    .C(_0114_),
    .Y(_0443_),
    .A_N(_0430_));
 sg13g2_a21oi_1 _1246_ (.A1(_0431_),
    .A2(_0443_),
    .Y(_0444_),
    .B1(net99));
 sg13g2_nand3_1 _1247_ (.B(\hidden_lif_0.variant_threshold[2] ),
    .C(\hidden_lif_0.variant_threshold[1] ),
    .A(\hidden_lif_0.variant_threshold[3] ),
    .Y(_0445_));
 sg13g2_nand2_1 _1248_ (.Y(_0446_),
    .A(net99),
    .B(_0445_));
 sg13g2_nand4_1 _1249_ (.B(net165),
    .C(\hidden_lif_0.variant_threshold[1] ),
    .A(_0114_),
    .Y(_0447_),
    .D(net99));
 sg13g2_nor2b_1 _1250_ (.A(_0444_),
    .B_N(_0447_),
    .Y(_0448_));
 sg13g2_nand2_2 _1251_ (.Y(_0449_),
    .A(net110),
    .B(_0434_));
 sg13g2_nand2_1 _1252_ (.Y(_0450_),
    .A(_0434_),
    .B(_0446_));
 sg13g2_nand3_1 _1253_ (.B(net110),
    .C(_0450_),
    .A(net168),
    .Y(_0451_));
 sg13g2_o21ai_1 _1254_ (.B1(_0451_),
    .Y(_0055_),
    .A1(_0448_),
    .A2(_0449_));
 sg13g2_nand2_1 _1255_ (.Y(_0452_),
    .A(_0147_),
    .B(_0443_));
 sg13g2_nand3_1 _1256_ (.B(_0446_),
    .C(_0452_),
    .A(net187),
    .Y(_0453_));
 sg13g2_a21oi_1 _1257_ (.A1(_0446_),
    .A2(_0452_),
    .Y(_0454_),
    .B1(net187));
 sg13g2_nand2_1 _1258_ (.Y(_0455_),
    .A(_0434_),
    .B(_0453_));
 sg13g2_o21ai_1 _1259_ (.B1(net110),
    .Y(_0056_),
    .A1(_0454_),
    .A2(_0455_));
 sg13g2_nor2_1 _1260_ (.A(_0113_),
    .B(_0445_),
    .Y(_0456_));
 sg13g2_nor3_1 _1261_ (.A(\hidden_lif_0.variant_threshold[4] ),
    .B(net99),
    .C(_0443_),
    .Y(_0457_));
 sg13g2_a21oi_1 _1262_ (.A1(net99),
    .A2(_0456_),
    .Y(_0458_),
    .B1(_0457_));
 sg13g2_xnor2_1 _1263_ (.Y(_0459_),
    .A(_0112_),
    .B(_0458_));
 sg13g2_nor2_1 _1264_ (.A(_0449_),
    .B(_0459_),
    .Y(_0057_));
 sg13g2_nor4_1 _1265_ (.A(_0112_),
    .B(_0113_),
    .C(_0147_),
    .D(_0445_),
    .Y(_0460_));
 sg13g2_a21oi_1 _1266_ (.A1(_0112_),
    .A2(_0457_),
    .Y(_0461_),
    .B1(_0460_));
 sg13g2_xnor2_1 _1267_ (.Y(_0462_),
    .A(_0111_),
    .B(_0461_));
 sg13g2_nor2_1 _1268_ (.A(_0449_),
    .B(_0462_),
    .Y(_0058_));
 sg13g2_a22oi_1 _1269_ (.Y(_0463_),
    .B1(_0460_),
    .B2(net227),
    .A2(_0457_),
    .A1(net229));
 sg13g2_xnor2_1 _1270_ (.Y(_0464_),
    .A(_0110_),
    .B(_0463_));
 sg13g2_nor2_1 _1271_ (.A(_0449_),
    .B(_0464_),
    .Y(_0059_));
 sg13g2_nand2b_1 _1272_ (.Y(_0465_),
    .B(_0001_),
    .A_N(_0208_));
 sg13g2_o21ai_1 _1273_ (.B1(net106),
    .Y(_0466_),
    .A1(_0211_),
    .A2(_0465_));
 sg13g2_a21oi_1 _1274_ (.A1(_0109_),
    .A2(_0465_),
    .Y(_0060_),
    .B1(_0466_));
 sg13g2_and2_1 _1275_ (.A(net93),
    .B(_0314_),
    .X(_0467_));
 sg13g2_nand2_1 _1276_ (.Y(_0468_),
    .A(\hidden_weight_1[0] ),
    .B(_0310_));
 sg13g2_or2_1 _1277_ (.X(_0469_),
    .B(_0468_),
    .A(_0321_));
 sg13g2_and2_1 _1278_ (.A(_0321_),
    .B(_0468_),
    .X(_0470_));
 sg13g2_xor2_1 _1279_ (.B(_0468_),
    .A(_0321_),
    .X(_0471_));
 sg13g2_xnor2_1 _1280_ (.Y(_0472_),
    .A(_0342_),
    .B(_0471_));
 sg13g2_and3_1 _1281_ (.X(_0473_),
    .A(\hidden_weight_1[0] ),
    .B(_0307_),
    .C(_0312_));
 sg13g2_and4_1 _1282_ (.A(net94),
    .B(net3),
    .C(net93),
    .D(_0304_),
    .X(_0474_));
 sg13g2_a22oi_1 _1283_ (.Y(_0475_),
    .B1(_0329_),
    .B2(net93),
    .A2(_0307_),
    .A1(net94));
 sg13g2_or3_1 _1284_ (.A(_0326_),
    .B(_0474_),
    .C(_0475_),
    .X(_0476_));
 sg13g2_o21ai_1 _1285_ (.B1(_0326_),
    .Y(_0477_),
    .A1(_0474_),
    .A2(_0475_));
 sg13g2_nand3_1 _1286_ (.B(_0476_),
    .C(_0477_),
    .A(_0473_),
    .Y(_0478_));
 sg13g2_a21o_1 _1287_ (.A2(_0477_),
    .A1(_0476_),
    .B1(_0473_),
    .X(_0479_));
 sg13g2_nand3_1 _1288_ (.B(_0478_),
    .C(_0479_),
    .A(_0472_),
    .Y(_0480_));
 sg13g2_a21o_1 _1289_ (.A2(_0479_),
    .A1(_0478_),
    .B1(_0472_),
    .X(_0481_));
 sg13g2_and3_1 _1290_ (.X(_0482_),
    .A(_0467_),
    .B(_0480_),
    .C(_0481_));
 sg13g2_nand3_1 _1291_ (.B(_0480_),
    .C(_0481_),
    .A(_0467_),
    .Y(_0483_));
 sg13g2_and3_1 _1292_ (.X(_0484_),
    .A(net7),
    .B(net8),
    .C(net93));
 sg13g2_a21o_1 _1293_ (.A2(_0481_),
    .A1(_0480_),
    .B1(_0467_),
    .X(_0485_));
 sg13g2_nand3_1 _1294_ (.B(_0484_),
    .C(_0485_),
    .A(_0483_),
    .Y(_0486_));
 sg13g2_a21oi_1 _1295_ (.A1(_0484_),
    .A2(_0485_),
    .Y(_0487_),
    .B1(_0482_));
 sg13g2_nand2_1 _1296_ (.Y(_0488_),
    .A(_0478_),
    .B(_0480_));
 sg13g2_o21ai_1 _1297_ (.B1(_0469_),
    .Y(_0489_),
    .A1(_0342_),
    .A2(_0470_));
 sg13g2_nor2b_1 _1298_ (.A(_0474_),
    .B_N(_0476_),
    .Y(_0490_));
 sg13g2_xor2_1 _1299_ (.B(_0490_),
    .A(_0489_),
    .X(_0491_));
 sg13g2_xnor2_1 _1300_ (.Y(_0492_),
    .A(_0324_),
    .B(_0334_));
 sg13g2_xnor2_1 _1301_ (.Y(_0493_),
    .A(_0491_),
    .B(_0492_));
 sg13g2_xnor2_1 _1302_ (.Y(_0494_),
    .A(_0488_),
    .B(_0493_));
 sg13g2_xor2_1 _1303_ (.B(_0494_),
    .A(_0487_),
    .X(_0495_));
 sg13g2_a21o_1 _1304_ (.A2(_0485_),
    .A1(_0483_),
    .B1(_0484_),
    .X(_0496_));
 sg13g2_a221oi_1 _1305_ (.B2(_0496_),
    .C1(_0495_),
    .B1(_0486_),
    .A1(net93),
    .Y(_0497_),
    .A2(_0315_));
 sg13g2_inv_1 _1306_ (.Y(_0498_),
    .A(net88));
 sg13g2_nand2_1 _1307_ (.Y(_0499_),
    .A(\hidden_lif_1.state_r[3] ),
    .B(_0146_));
 sg13g2_nand2_1 _1308_ (.Y(_0500_),
    .A(_0144_),
    .B(net241));
 sg13g2_nand3_1 _1309_ (.B(_0499_),
    .C(_0500_),
    .A(net89),
    .Y(_0501_));
 sg13g2_a21oi_1 _1310_ (.A1(net93),
    .A2(_0315_),
    .Y(_0502_),
    .B1(\hidden_lif_1.state_r[1] ));
 sg13g2_nand2b_1 _1311_ (.Y(_0503_),
    .B(\hidden_lif_1.state_r[6] ),
    .A_N(\hidden_lif_1.variant_threshold[6] ));
 sg13g2_nor2b_1 _1312_ (.A(\hidden_lif_1.state_r[5] ),
    .B_N(\hidden_lif_1.variant_threshold[5] ),
    .Y(_0504_));
 sg13g2_nand2b_1 _1313_ (.Y(_0505_),
    .B(\hidden_lif_1.state_r[2] ),
    .A_N(\hidden_lif_1.variant_threshold[2] ));
 sg13g2_a22oi_1 _1314_ (.Y(_0506_),
    .B1(_0146_),
    .B2(\hidden_lif_1.variant_threshold[0] ),
    .A2(_0145_),
    .A1(\hidden_lif_1.variant_threshold[1] ));
 sg13g2_o21ai_1 _1315_ (.B1(_0505_),
    .Y(_0507_),
    .A1(\hidden_lif_1.variant_threshold[1] ),
    .A2(_0145_));
 sg13g2_nand2b_1 _1316_ (.Y(_0508_),
    .B(\hidden_lif_1.variant_threshold[2] ),
    .A_N(\hidden_lif_1.state_r[2] ));
 sg13g2_o21ai_1 _1317_ (.B1(_0508_),
    .Y(_0509_),
    .A1(_0506_),
    .A2(_0507_));
 sg13g2_o21ai_1 _1318_ (.B1(_0509_),
    .Y(_0510_),
    .A1(\hidden_lif_1.variant_threshold[3] ),
    .A2(_0144_));
 sg13g2_a22oi_1 _1319_ (.Y(_0511_),
    .B1(_0144_),
    .B2(\hidden_lif_1.variant_threshold[3] ),
    .A2(_0143_),
    .A1(\hidden_lif_1.variant_threshold[4] ));
 sg13g2_nor2_1 _1320_ (.A(\hidden_lif_1.variant_threshold[5] ),
    .B(_0142_),
    .Y(_0512_));
 sg13g2_a221oi_1 _1321_ (.B2(_0511_),
    .C1(_0512_),
    .B1(_0510_),
    .A1(_0131_),
    .Y(_0513_),
    .A2(\hidden_lif_1.state_r[4] ));
 sg13g2_o21ai_1 _1322_ (.B1(_0503_),
    .Y(_0514_),
    .A1(_0504_),
    .A2(_0513_));
 sg13g2_a22oi_1 _1323_ (.Y(_0515_),
    .B1(_0141_),
    .B2(net244),
    .A2(_0140_),
    .A1(net213));
 sg13g2_a22oi_1 _1324_ (.Y(_0516_),
    .B1(_0514_),
    .B2(_0515_),
    .A2(net190),
    .A1(_0130_));
 sg13g2_nand2_2 _1325_ (.Y(_0517_),
    .A(net107),
    .B(_0516_));
 sg13g2_nand3_1 _1326_ (.B(net93),
    .C(_0315_),
    .A(\hidden_lif_1.state_r[1] ),
    .Y(_0518_));
 sg13g2_nor2b_1 _1327_ (.A(_0502_),
    .B_N(_0518_),
    .Y(_0519_));
 sg13g2_o21ai_1 _1328_ (.B1(_0501_),
    .Y(_0520_),
    .A1(net89),
    .A2(_0519_));
 sg13g2_nor2_1 _1329_ (.A(_0517_),
    .B(net242),
    .Y(_0061_));
 sg13g2_and3_1 _1330_ (.X(_0521_),
    .A(_0163_),
    .B(_0486_),
    .C(_0496_));
 sg13g2_a21oi_1 _1331_ (.A1(_0486_),
    .A2(_0496_),
    .Y(_0522_),
    .B1(_0163_));
 sg13g2_or2_1 _1332_ (.X(_0523_),
    .B(_0522_),
    .A(_0521_));
 sg13g2_nor3_2 _1333_ (.A(_0518_),
    .B(_0521_),
    .C(_0522_),
    .Y(_0524_));
 sg13g2_inv_1 _1334_ (.Y(_0525_),
    .A(_0524_));
 sg13g2_o21ai_1 _1335_ (.B1(_0518_),
    .Y(_0526_),
    .A1(net89),
    .A2(_0523_));
 sg13g2_nor2b_1 _1336_ (.A(\hidden_lif_1.state_r[4] ),
    .B_N(\hidden_lif_1.state_r[1] ),
    .Y(_0527_));
 sg13g2_xnor2_1 _1337_ (.Y(_0528_),
    .A(\hidden_lif_1.state_r[4] ),
    .B(\hidden_lif_1.state_r[1] ));
 sg13g2_xor2_1 _1338_ (.B(_0528_),
    .A(_0499_),
    .X(_0529_));
 sg13g2_a22oi_1 _1339_ (.Y(_0530_),
    .B1(_0529_),
    .B2(net88),
    .A2(_0526_),
    .A1(_0525_));
 sg13g2_nor2_1 _1340_ (.A(_0517_),
    .B(_0530_),
    .Y(_0062_));
 sg13g2_nand2_1 _1341_ (.Y(_0531_),
    .A(\hidden_lif_1.state_r[3] ),
    .B(_0495_));
 sg13g2_xnor2_1 _1342_ (.Y(_0532_),
    .A(_0144_),
    .B(_0495_));
 sg13g2_o21ai_1 _1343_ (.B1(_0532_),
    .Y(_0533_),
    .A1(_0521_),
    .A2(_0524_));
 sg13g2_or3_1 _1344_ (.A(_0521_),
    .B(_0524_),
    .C(_0532_),
    .X(_0534_));
 sg13g2_nand3_1 _1345_ (.B(_0533_),
    .C(_0534_),
    .A(_0498_),
    .Y(_0535_));
 sg13g2_xnor2_1 _1346_ (.Y(_0536_),
    .A(\hidden_lif_1.state_r[5] ),
    .B(\hidden_lif_1.state_r[2] ));
 sg13g2_a21oi_1 _1347_ (.A1(_0499_),
    .A2(_0528_),
    .Y(_0537_),
    .B1(_0527_));
 sg13g2_nor2b_1 _1348_ (.A(_0537_),
    .B_N(_0536_),
    .Y(_0538_));
 sg13g2_nand2b_1 _1349_ (.Y(_0539_),
    .B(_0537_),
    .A_N(_0536_));
 sg13g2_nand3b_1 _1350_ (.B(_0539_),
    .C(net88),
    .Y(_0540_),
    .A_N(_0538_));
 sg13g2_a21oi_1 _1351_ (.A1(_0535_),
    .A2(_0540_),
    .Y(_0063_),
    .B1(_0517_));
 sg13g2_nand2_1 _1352_ (.Y(_0541_),
    .A(_0141_),
    .B(\hidden_lif_1.state_r[3] ));
 sg13g2_xor2_1 _1353_ (.B(\hidden_lif_1.state_r[3] ),
    .A(\hidden_lif_1.state_r[6] ),
    .X(_0542_));
 sg13g2_a21oi_1 _1354_ (.A1(_0142_),
    .A2(\hidden_lif_1.state_r[2] ),
    .Y(_0543_),
    .B1(_0538_));
 sg13g2_xor2_1 _1355_ (.B(_0543_),
    .A(_0542_),
    .X(_0544_));
 sg13g2_nand3_1 _1356_ (.B(_0531_),
    .C(_0533_),
    .A(net184),
    .Y(_0545_));
 sg13g2_a21oi_2 _1357_ (.B1(net184),
    .Y(_0546_),
    .A2(_0533_),
    .A1(_0531_));
 sg13g2_nor2_1 _1358_ (.A(net89),
    .B(_0546_),
    .Y(_0547_));
 sg13g2_a22oi_1 _1359_ (.Y(_0548_),
    .B1(_0545_),
    .B2(_0547_),
    .A2(_0544_),
    .A1(net88));
 sg13g2_nor2_1 _1360_ (.A(_0517_),
    .B(_0548_),
    .Y(_0064_));
 sg13g2_nand2_1 _1361_ (.Y(_0549_),
    .A(\hidden_lif_1.state_r[7] ),
    .B(_0143_));
 sg13g2_nor2_1 _1362_ (.A(\hidden_lif_1.state_r[7] ),
    .B(_0143_),
    .Y(_0550_));
 sg13g2_nand2_1 _1363_ (.Y(_0551_),
    .A(_0140_),
    .B(\hidden_lif_1.state_r[4] ));
 sg13g2_and2_1 _1364_ (.A(_0549_),
    .B(_0551_),
    .X(_0552_));
 sg13g2_o21ai_1 _1365_ (.B1(_0541_),
    .Y(_0553_),
    .A1(_0542_),
    .A2(_0543_));
 sg13g2_xnor2_1 _1366_ (.Y(_0554_),
    .A(_0552_),
    .B(_0553_));
 sg13g2_xor2_1 _1367_ (.B(_0546_),
    .A(net169),
    .X(_0555_));
 sg13g2_a21o_1 _1368_ (.A2(_0554_),
    .A1(net88),
    .B1(_0517_),
    .X(_0556_));
 sg13g2_a21oi_1 _1369_ (.A1(_0498_),
    .A2(net170),
    .Y(_0065_),
    .B1(_0556_));
 sg13g2_a21o_1 _1370_ (.A2(_0546_),
    .A1(net246),
    .B1(net245),
    .X(_0557_));
 sg13g2_nor2_1 _1371_ (.A(_0141_),
    .B(_0142_),
    .Y(_0558_));
 sg13g2_nand2_1 _1372_ (.Y(_0559_),
    .A(_0546_),
    .B(_0558_));
 sg13g2_a21oi_1 _1373_ (.A1(_0546_),
    .A2(_0558_),
    .Y(_0560_),
    .B1(net88));
 sg13g2_a21oi_1 _1374_ (.A1(_0549_),
    .A2(_0553_),
    .Y(_0561_),
    .B1(_0550_));
 sg13g2_xnor2_1 _1375_ (.Y(_0562_),
    .A(_0142_),
    .B(_0561_));
 sg13g2_a22oi_1 _1376_ (.Y(_0563_),
    .B1(_0562_),
    .B2(net88),
    .A2(_0560_),
    .A1(_0557_));
 sg13g2_nor2_1 _1377_ (.A(_0517_),
    .B(net247),
    .Y(_0066_));
 sg13g2_xnor2_1 _1378_ (.Y(_0564_),
    .A(_0140_),
    .B(_0559_));
 sg13g2_a21oi_1 _1379_ (.A1(\hidden_lif_1.state_r[5] ),
    .A2(_0551_),
    .Y(_0565_),
    .B1(_0561_));
 sg13g2_nor2b_1 _1380_ (.A(_0565_),
    .B_N(net169),
    .Y(_0566_));
 sg13g2_and2_1 _1381_ (.A(_0141_),
    .B(_0566_),
    .X(_0567_));
 sg13g2_xnor2_1 _1382_ (.Y(_0568_),
    .A(net245),
    .B(_0566_));
 sg13g2_a21o_1 _1383_ (.A2(_0568_),
    .A1(net88),
    .B1(_0517_),
    .X(_0569_));
 sg13g2_a21oi_1 _1384_ (.A1(_0498_),
    .A2(_0564_),
    .Y(_0067_),
    .B1(_0569_));
 sg13g2_xnor2_1 _1385_ (.Y(_0570_),
    .A(net190),
    .B(_0567_));
 sg13g2_nor3_1 _1386_ (.A(_0517_),
    .B(_0560_),
    .C(_0570_),
    .Y(_0068_));
 sg13g2_nor2_1 _1387_ (.A(net105),
    .B(_0516_),
    .Y(_0069_));
 sg13g2_nor2b_1 _1388_ (.A(_0248_),
    .B_N(net175),
    .Y(_0571_));
 sg13g2_nand2b_1 _1389_ (.Y(_0572_),
    .B(_0571_),
    .A_N(_0253_));
 sg13g2_o21ai_1 _1390_ (.B1(net108),
    .Y(_0573_),
    .A1(net188),
    .A2(_0571_));
 sg13g2_nor2b_1 _1391_ (.A(_0573_),
    .B_N(_0572_),
    .Y(_0070_));
 sg13g2_nor2_1 _1392_ (.A(_0152_),
    .B(\hidden_lif_2.state_r[0] ),
    .Y(_0574_));
 sg13g2_xnor2_1 _1393_ (.Y(_0575_),
    .A(\hidden_lif_2.state_r[3] ),
    .B(net215));
 sg13g2_nor2_1 _1394_ (.A(\hidden_lif_2.state_r[1] ),
    .B(_0316_),
    .Y(_0576_));
 sg13g2_nand2_2 _1395_ (.Y(_0577_),
    .A(net110),
    .B(_0290_));
 sg13g2_nand2_1 _1396_ (.Y(_0578_),
    .A(\hidden_lif_2.state_r[1] ),
    .B(_0316_));
 sg13g2_nand3_1 _1397_ (.B(_0290_),
    .C(_0578_),
    .A(net110),
    .Y(_0579_));
 sg13g2_a221oi_1 _1398_ (.B2(_0361_),
    .C1(_0579_),
    .B1(_0576_),
    .A1(net85),
    .Y(_0071_),
    .A2(net216));
 sg13g2_nor3_2 _1399_ (.A(_0013_),
    .B(_0345_),
    .C(_0359_),
    .Y(_0580_));
 sg13g2_a21oi_1 _1400_ (.A1(_0346_),
    .A2(_0360_),
    .Y(_0581_),
    .B1(_0165_));
 sg13g2_nor2_1 _1401_ (.A(_0580_),
    .B(_0581_),
    .Y(_0582_));
 sg13g2_nor3_2 _1402_ (.A(_0578_),
    .B(_0580_),
    .C(_0581_),
    .Y(_0583_));
 sg13g2_a22oi_1 _1403_ (.Y(_0584_),
    .B1(_0363_),
    .B2(_0582_),
    .A2(_0316_),
    .A1(net249));
 sg13g2_nor2b_1 _1404_ (.A(\hidden_lif_2.state_r[4] ),
    .B_N(\hidden_lif_2.state_r[1] ),
    .Y(_0585_));
 sg13g2_xor2_1 _1405_ (.B(\hidden_lif_2.state_r[1] ),
    .A(\hidden_lif_2.state_r[4] ),
    .X(_0586_));
 sg13g2_nand2_1 _1406_ (.Y(_0587_),
    .A(_0574_),
    .B(_0586_));
 sg13g2_nor2_1 _1407_ (.A(_0574_),
    .B(_0586_),
    .Y(_0588_));
 sg13g2_nand3b_1 _1408_ (.B(net87),
    .C(_0587_),
    .Y(_0589_),
    .A_N(_0588_));
 sg13g2_o21ai_1 _1409_ (.B1(_0589_),
    .Y(_0590_),
    .A1(_0583_),
    .A2(_0584_));
 sg13g2_nor2b_1 _1410_ (.A(_0577_),
    .B_N(_0590_),
    .Y(_0072_));
 sg13g2_nand2b_1 _1411_ (.Y(_0591_),
    .B(\hidden_lif_2.state_r[3] ),
    .A_N(_0358_));
 sg13g2_xnor2_1 _1412_ (.Y(_0592_),
    .A(\hidden_lif_2.state_r[3] ),
    .B(_0358_));
 sg13g2_nor2_1 _1413_ (.A(_0580_),
    .B(_0583_),
    .Y(_0593_));
 sg13g2_o21ai_1 _1414_ (.B1(_0592_),
    .Y(_0594_),
    .A1(_0580_),
    .A2(_0583_));
 sg13g2_nand2_1 _1415_ (.Y(_0595_),
    .A(_0150_),
    .B(\hidden_lif_2.state_r[2] ));
 sg13g2_xnor2_1 _1416_ (.Y(_0596_),
    .A(\hidden_lif_2.state_r[5] ),
    .B(\hidden_lif_2.state_r[2] ));
 sg13g2_o21ai_1 _1417_ (.B1(_0596_),
    .Y(_0597_),
    .A1(_0585_),
    .A2(_0588_));
 sg13g2_or3_1 _1418_ (.A(_0585_),
    .B(_0588_),
    .C(_0596_),
    .X(_0598_));
 sg13g2_a21o_1 _1419_ (.A2(_0598_),
    .A1(_0597_),
    .B1(_0363_),
    .X(_0599_));
 sg13g2_xnor2_1 _1420_ (.Y(_0600_),
    .A(_0592_),
    .B(_0593_));
 sg13g2_o21ai_1 _1421_ (.B1(_0599_),
    .Y(_0601_),
    .A1(net85),
    .A2(_0600_));
 sg13g2_nor2_1 _1422_ (.A(_0577_),
    .B(_0601_),
    .Y(_0073_));
 sg13g2_nor2_1 _1423_ (.A(\hidden_lif_2.state_r[6] ),
    .B(_0152_),
    .Y(_0602_));
 sg13g2_xor2_1 _1424_ (.B(\hidden_lif_2.state_r[3] ),
    .A(\hidden_lif_2.state_r[6] ),
    .X(_0603_));
 sg13g2_nand3_1 _1425_ (.B(_0597_),
    .C(_0603_),
    .A(_0595_),
    .Y(_0604_));
 sg13g2_a21oi_1 _1426_ (.A1(_0595_),
    .A2(_0597_),
    .Y(_0605_),
    .B1(_0603_));
 sg13g2_nand3b_1 _1427_ (.B(net85),
    .C(_0604_),
    .Y(_0606_),
    .A_N(_0605_));
 sg13g2_nand3_1 _1428_ (.B(_0591_),
    .C(_0594_),
    .A(net203),
    .Y(_0607_));
 sg13g2_a21oi_2 _1429_ (.B1(net203),
    .Y(_0608_),
    .A2(_0594_),
    .A1(_0591_));
 sg13g2_nor2_1 _1430_ (.A(net85),
    .B(_0608_),
    .Y(_0609_));
 sg13g2_nand2_1 _1431_ (.Y(_0610_),
    .A(_0607_),
    .B(_0609_));
 sg13g2_a21oi_1 _1432_ (.A1(_0606_),
    .A2(_0610_),
    .Y(_0074_),
    .B1(_0577_));
 sg13g2_nand2_1 _1433_ (.Y(_0611_),
    .A(_0148_),
    .B(\hidden_lif_2.state_r[4] ));
 sg13g2_xnor2_1 _1434_ (.Y(_0612_),
    .A(\hidden_lif_2.state_r[7] ),
    .B(\hidden_lif_2.state_r[4] ));
 sg13g2_nor3_1 _1435_ (.A(_0602_),
    .B(_0605_),
    .C(_0612_),
    .Y(_0613_));
 sg13g2_o21ai_1 _1436_ (.B1(_0612_),
    .Y(_0614_),
    .A1(_0602_),
    .A2(_0605_));
 sg13g2_nand2b_1 _1437_ (.Y(_0615_),
    .B(_0614_),
    .A_N(_0613_));
 sg13g2_xor2_1 _1438_ (.B(_0608_),
    .A(net177),
    .X(_0616_));
 sg13g2_a21o_1 _1439_ (.A2(_0615_),
    .A1(net85),
    .B1(_0577_),
    .X(_0617_));
 sg13g2_a21oi_1 _1440_ (.A1(_0363_),
    .A2(net178),
    .Y(_0075_),
    .B1(_0617_));
 sg13g2_a21o_1 _1441_ (.A2(_0608_),
    .A1(\hidden_lif_2.state_r[5] ),
    .B1(net222),
    .X(_0618_));
 sg13g2_nand3_1 _1442_ (.B(\hidden_lif_2.state_r[5] ),
    .C(_0608_),
    .A(net222),
    .Y(_0619_));
 sg13g2_nand3_1 _1443_ (.B(_0618_),
    .C(_0619_),
    .A(_0363_),
    .Y(_0620_));
 sg13g2_nand2_1 _1444_ (.Y(_0621_),
    .A(_0611_),
    .B(_0614_));
 sg13g2_xnor2_1 _1445_ (.Y(_0622_),
    .A(\hidden_lif_2.state_r[5] ),
    .B(_0621_));
 sg13g2_nand2_1 _1446_ (.Y(_0623_),
    .A(net85),
    .B(_0622_));
 sg13g2_a21oi_1 _1447_ (.A1(_0620_),
    .A2(_0623_),
    .Y(_0076_),
    .B1(_0577_));
 sg13g2_nand2b_1 _1448_ (.Y(_0624_),
    .B(_0148_),
    .A_N(_0619_));
 sg13g2_a21oi_1 _1449_ (.A1(net231),
    .A2(_0619_),
    .Y(_0625_),
    .B1(net85));
 sg13g2_and2_1 _1450_ (.A(_0015_),
    .B(_0611_),
    .X(_0626_));
 sg13g2_o21ai_1 _1451_ (.B1(_0626_),
    .Y(_0627_),
    .A1(\hidden_lif_2.state_r[5] ),
    .A2(_0614_));
 sg13g2_nor2_1 _1452_ (.A(\hidden_lif_2.state_r[6] ),
    .B(_0627_),
    .Y(_0628_));
 sg13g2_xnor2_1 _1453_ (.Y(_0629_),
    .A(_0149_),
    .B(_0627_));
 sg13g2_a221oi_1 _1454_ (.B2(net85),
    .C1(_0577_),
    .B1(_0629_),
    .A1(_0624_),
    .Y(_0077_),
    .A2(_0625_));
 sg13g2_xnor2_1 _1455_ (.Y(_0630_),
    .A(_0148_),
    .B(_0628_));
 sg13g2_nand2b_1 _1456_ (.Y(_0631_),
    .B(_0630_),
    .A_N(_0577_));
 sg13g2_a21oi_1 _1457_ (.A1(_0363_),
    .A2(net223),
    .Y(_0078_),
    .B1(_0631_));
 sg13g2_xnor2_1 _1458_ (.Y(_0632_),
    .A(net150),
    .B(net93));
 sg13g2_nor2_1 _1459_ (.A(_0139_),
    .B(_0632_),
    .Y(_0079_));
 sg13g2_and2_1 _1460_ (.A(net111),
    .B(net94),
    .X(_0080_));
 sg13g2_nand2b_1 _1461_ (.Y(_0081_),
    .B(net111),
    .A_N(net183));
 sg13g2_nand2b_1 _1462_ (.Y(_0082_),
    .B(net111),
    .A_N(net150));
 sg13g2_nand2b_1 _1463_ (.Y(_0633_),
    .B(net156),
    .A_N(_0433_));
 sg13g2_o21ai_1 _1464_ (.B1(net110),
    .Y(_0634_),
    .A1(_0436_),
    .A2(_0633_));
 sg13g2_a21oi_1 _1465_ (.A1(_0108_),
    .A2(_0633_),
    .Y(_0083_),
    .B1(_0634_));
 sg13g2_nand2_1 _1466_ (.Y(_0635_),
    .A(net98),
    .B(net100));
 sg13g2_xnor2_1 _1467_ (.Y(_0636_),
    .A(net98),
    .B(net100));
 sg13g2_xnor2_1 _1468_ (.Y(_0637_),
    .A(net103),
    .B(_0636_));
 sg13g2_nand2_1 _1469_ (.Y(_0638_),
    .A(net139),
    .B(_0637_));
 sg13g2_inv_1 _1470_ (.Y(_0639_),
    .A(_0638_));
 sg13g2_nand2_1 _1471_ (.Y(_0640_),
    .A(\output_weight_0[2] ),
    .B(_0637_));
 sg13g2_o21ai_1 _1472_ (.B1(_0635_),
    .Y(_0641_),
    .A1(_0133_),
    .A2(_0636_));
 sg13g2_nand3_1 _1473_ (.B(_0638_),
    .C(_0641_),
    .A(\output_weight_0[1] ),
    .Y(_0642_));
 sg13g2_xor2_1 _1474_ (.B(_0642_),
    .A(_0640_),
    .X(_0643_));
 sg13g2_nand2_1 _1475_ (.Y(_0644_),
    .A(\output_weight_0[1] ),
    .B(_0637_));
 sg13g2_nand2_1 _1476_ (.Y(_0645_),
    .A(\output_weight_0[0] ),
    .B(_0641_));
 sg13g2_xor2_1 _1477_ (.B(_0645_),
    .A(_0644_),
    .X(_0646_));
 sg13g2_nor3_1 _1478_ (.A(_0639_),
    .B(_0643_),
    .C(_0646_),
    .Y(_0647_));
 sg13g2_nor2_1 _1479_ (.A(net235),
    .B(_0154_),
    .Y(_0648_));
 sg13g2_nand2_1 _1480_ (.Y(_0649_),
    .A(net235),
    .B(_0154_));
 sg13g2_nand3b_1 _1481_ (.B(_0649_),
    .C(net91),
    .Y(_0650_),
    .A_N(_0648_));
 sg13g2_nand2b_2 _1482_ (.Y(_0651_),
    .B(net108),
    .A_N(_0300_));
 sg13g2_nand2_1 _1483_ (.Y(_0652_),
    .A(\output_lif_0.state_r[1] ),
    .B(_0639_));
 sg13g2_xnor2_1 _1484_ (.Y(_0653_),
    .A(\output_lif_0.state_r[1] ),
    .B(_0638_));
 sg13g2_o21ai_1 _1485_ (.B1(_0650_),
    .Y(_0654_),
    .A1(net91),
    .A2(_0653_));
 sg13g2_nor2_1 _1486_ (.A(_0651_),
    .B(_0654_),
    .Y(_0084_));
 sg13g2_nand2_1 _1487_ (.Y(_0655_),
    .A(\output_lif_0.state_r[2] ),
    .B(_0646_));
 sg13g2_xnor2_1 _1488_ (.Y(_0656_),
    .A(\output_lif_0.state_r[2] ),
    .B(_0646_));
 sg13g2_or2_1 _1489_ (.X(_0657_),
    .B(_0656_),
    .A(_0652_));
 sg13g2_a21oi_1 _1490_ (.A1(_0652_),
    .A2(_0656_),
    .Y(_0658_),
    .B1(net91));
 sg13g2_xnor2_1 _1491_ (.Y(_0659_),
    .A(\output_lif_0.state_r[1] ),
    .B(\output_lif_0.state_r[4] ));
 sg13g2_nor2b_1 _1492_ (.A(_0648_),
    .B_N(_0659_),
    .Y(_0660_));
 sg13g2_xnor2_1 _1493_ (.Y(_0661_),
    .A(_0648_),
    .B(_0659_));
 sg13g2_a22oi_1 _1494_ (.Y(_0662_),
    .B1(_0661_),
    .B2(net91),
    .A2(_0658_),
    .A1(_0657_));
 sg13g2_nor2_1 _1495_ (.A(_0651_),
    .B(_0662_),
    .Y(_0085_));
 sg13g2_and2_1 _1496_ (.A(\output_lif_0.state_r[3] ),
    .B(_0643_),
    .X(_0663_));
 sg13g2_nand2_1 _1497_ (.Y(_0664_),
    .A(\output_lif_0.state_r[3] ),
    .B(_0643_));
 sg13g2_xnor2_1 _1498_ (.Y(_0665_),
    .A(\output_lif_0.state_r[3] ),
    .B(_0643_));
 sg13g2_a21oi_2 _1499_ (.B1(_0665_),
    .Y(_0666_),
    .A2(_0657_),
    .A1(_0655_));
 sg13g2_and3_1 _1500_ (.X(_0667_),
    .A(_0655_),
    .B(_0657_),
    .C(_0665_));
 sg13g2_nor3_1 _1501_ (.A(net91),
    .B(_0666_),
    .C(_0667_),
    .Y(_0668_));
 sg13g2_xnor2_1 _1502_ (.Y(_0669_),
    .A(\output_lif_0.state_r[2] ),
    .B(\output_lif_0.state_r[5] ));
 sg13g2_a21oi_1 _1503_ (.A1(\output_lif_0.state_r[1] ),
    .A2(_0157_),
    .Y(_0670_),
    .B1(_0660_));
 sg13g2_nor2b_1 _1504_ (.A(_0670_),
    .B_N(_0669_),
    .Y(_0671_));
 sg13g2_xnor2_1 _1505_ (.Y(_0672_),
    .A(_0669_),
    .B(_0670_));
 sg13g2_a21oi_1 _1506_ (.A1(net90),
    .A2(_0672_),
    .Y(_0673_),
    .B1(_0668_));
 sg13g2_nor2_1 _1507_ (.A(_0651_),
    .B(_0673_),
    .Y(_0086_));
 sg13g2_o21ai_1 _1508_ (.B1(net154),
    .Y(_0674_),
    .A1(_0663_),
    .A2(_0666_));
 sg13g2_nor3_1 _1509_ (.A(net154),
    .B(_0663_),
    .C(_0666_),
    .Y(_0675_));
 sg13g2_nor2_1 _1510_ (.A(net91),
    .B(_0675_),
    .Y(_0676_));
 sg13g2_nor2_1 _1511_ (.A(_0154_),
    .B(\output_lif_0.state_r[6] ),
    .Y(_0677_));
 sg13g2_xnor2_1 _1512_ (.Y(_0678_),
    .A(\output_lif_0.state_r[3] ),
    .B(net92));
 sg13g2_a21oi_1 _1513_ (.A1(\output_lif_0.state_r[2] ),
    .A2(_0156_),
    .Y(_0679_),
    .B1(_0671_));
 sg13g2_nor2b_1 _1514_ (.A(_0679_),
    .B_N(_0678_),
    .Y(_0680_));
 sg13g2_xor2_1 _1515_ (.B(_0679_),
    .A(_0678_),
    .X(_0681_));
 sg13g2_a221oi_1 _1516_ (.B2(net90),
    .C1(_0651_),
    .B1(_0681_),
    .A1(_0674_),
    .Y(_0087_),
    .A2(_0676_));
 sg13g2_nand2_1 _1517_ (.Y(_0682_),
    .A(\output_lif_0.state_r[4] ),
    .B(_0666_));
 sg13g2_o21ai_1 _1518_ (.B1(_0682_),
    .Y(_0683_),
    .A1(_0017_),
    .A2(_0664_));
 sg13g2_nand2_1 _1519_ (.Y(_0684_),
    .A(\output_lif_0.state_r[4] ),
    .B(_0158_));
 sg13g2_xnor2_1 _1520_ (.Y(_0685_),
    .A(\output_lif_0.state_r[4] ),
    .B(\output_lif_0.state_r[7] ));
 sg13g2_o21ai_1 _1521_ (.B1(_0685_),
    .Y(_0686_),
    .A1(_0677_),
    .A2(_0680_));
 sg13g2_or3_1 _1522_ (.A(_0677_),
    .B(_0680_),
    .C(_0685_),
    .X(_0687_));
 sg13g2_nand2_1 _1523_ (.Y(_0688_),
    .A(_0686_),
    .B(_0687_));
 sg13g2_xnor2_1 _1524_ (.Y(_0689_),
    .A(net205),
    .B(_0683_));
 sg13g2_a21oi_1 _1525_ (.A1(net90),
    .A2(_0688_),
    .Y(_0690_),
    .B1(_0651_));
 sg13g2_o21ai_1 _1526_ (.B1(_0690_),
    .Y(_0691_),
    .A1(net90),
    .A2(net206));
 sg13g2_inv_1 _1527_ (.Y(_0088_),
    .A(_0691_));
 sg13g2_and2_1 _1528_ (.A(\output_lif_0.state_r[5] ),
    .B(_0683_),
    .X(_0692_));
 sg13g2_nand2_1 _1529_ (.Y(_0693_),
    .A(net92),
    .B(_0692_));
 sg13g2_a21oi_1 _1530_ (.A1(net92),
    .A2(_0692_),
    .Y(_0694_),
    .B1(net90));
 sg13g2_o21ai_1 _1531_ (.B1(_0694_),
    .Y(_0695_),
    .A1(net92),
    .A2(_0692_));
 sg13g2_nand2_1 _1532_ (.Y(_0696_),
    .A(_0684_),
    .B(_0686_));
 sg13g2_xnor2_1 _1533_ (.Y(_0697_),
    .A(net248),
    .B(_0696_));
 sg13g2_nand2_1 _1534_ (.Y(_0698_),
    .A(net90),
    .B(_0697_));
 sg13g2_a21oi_1 _1535_ (.A1(_0695_),
    .A2(_0698_),
    .Y(_0089_),
    .B1(_0651_));
 sg13g2_nand2_1 _1536_ (.Y(_0699_),
    .A(net205),
    .B(_0684_));
 sg13g2_a21o_1 _1537_ (.A2(_0696_),
    .A1(_0156_),
    .B1(_0699_),
    .X(_0700_));
 sg13g2_nor2_1 _1538_ (.A(net92),
    .B(_0700_),
    .Y(_0701_));
 sg13g2_xnor2_1 _1539_ (.Y(_0702_),
    .A(net92),
    .B(_0700_));
 sg13g2_xnor2_1 _1540_ (.Y(_0703_),
    .A(_0158_),
    .B(_0693_));
 sg13g2_nor2_1 _1541_ (.A(net90),
    .B(_0703_),
    .Y(_0704_));
 sg13g2_a21oi_1 _1542_ (.A1(net90),
    .A2(_0702_),
    .Y(_0705_),
    .B1(_0704_));
 sg13g2_nor2_1 _1543_ (.A(_0651_),
    .B(_0705_),
    .Y(_0090_));
 sg13g2_xnor2_1 _1544_ (.Y(_0706_),
    .A(net180),
    .B(_0701_));
 sg13g2_nor3_1 _1545_ (.A(_0651_),
    .B(_0694_),
    .C(net181),
    .Y(_0091_));
 sg13g2_xnor2_1 _1546_ (.Y(_0707_),
    .A(net142),
    .B(net155));
 sg13g2_nand2_1 _1547_ (.Y(_0092_),
    .A(net106),
    .B(_0707_));
 sg13g2_nand2b_1 _1548_ (.Y(_0093_),
    .B(net106),
    .A_N(net139));
 sg13g2_and2_1 _1549_ (.A(net106),
    .B(net138),
    .X(_0094_));
 sg13g2_and2_1 _1550_ (.A(net106),
    .B(net142),
    .X(_0095_));
 sg13g2_o21ai_1 _1551_ (.B1(net111),
    .Y(_0708_),
    .A1(net102),
    .A2(uo_out[0]));
 sg13g2_a21oi_1 _1552_ (.A1(net102),
    .A2(_0107_),
    .Y(_0096_),
    .B1(_0708_));
 sg13g2_a21oi_1 _1553_ (.A1(net102),
    .A2(uo_out[0]),
    .Y(_0709_),
    .B1(net145));
 sg13g2_nand3_1 _1554_ (.B(net145),
    .C(uo_out[0]),
    .A(net102),
    .Y(_0710_));
 sg13g2_nand2_1 _1555_ (.Y(_0711_),
    .A(net111),
    .B(_0710_));
 sg13g2_nor2_1 _1556_ (.A(net146),
    .B(_0711_),
    .Y(_0097_));
 sg13g2_and2_1 _1557_ (.A(_0106_),
    .B(_0710_),
    .X(_0712_));
 sg13g2_nor2_1 _1558_ (.A(_0106_),
    .B(_0710_),
    .Y(_0713_));
 sg13g2_nor3_1 _1559_ (.A(net105),
    .B(net221),
    .C(_0713_),
    .Y(_0098_));
 sg13g2_nor2_1 _1560_ (.A(net163),
    .B(_0713_),
    .Y(_0714_));
 sg13g2_and2_2 _1561_ (.A(net163),
    .B(_0713_),
    .X(_0715_));
 sg13g2_nor3_1 _1562_ (.A(net105),
    .B(net164),
    .C(_0715_),
    .Y(_0099_));
 sg13g2_xnor2_1 _1563_ (.Y(_0716_),
    .A(net202),
    .B(_0715_));
 sg13g2_nor2_1 _1564_ (.A(net105),
    .B(_0716_),
    .Y(_0100_));
 sg13g2_a21oi_1 _1565_ (.A1(uo_out[4]),
    .A2(_0715_),
    .Y(_0717_),
    .B1(net151));
 sg13g2_nand3_1 _1566_ (.B(net202),
    .C(_0715_),
    .A(net151),
    .Y(_0718_));
 sg13g2_nand2_1 _1567_ (.Y(_0719_),
    .A(net109),
    .B(_0718_));
 sg13g2_nor2_1 _1568_ (.A(net152),
    .B(_0719_),
    .Y(_0101_));
 sg13g2_nand2b_1 _1569_ (.Y(_0720_),
    .B(_0718_),
    .A_N(net225));
 sg13g2_nand4_1 _1570_ (.B(net151),
    .C(uo_out[4]),
    .A(net225),
    .Y(_0721_),
    .D(_0715_));
 sg13g2_and3_1 _1571_ (.X(_0102_),
    .A(net107),
    .B(_0720_),
    .C(_0721_));
 sg13g2_o21ai_1 _1572_ (.B1(net107),
    .Y(_0722_),
    .A1(_0104_),
    .A2(_0721_));
 sg13g2_a21oi_1 _1573_ (.A1(_0104_),
    .A2(_0721_),
    .Y(_0103_),
    .B1(_0722_));
 sg13g2_dfrbp_1 _1574_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net77),
    .D(net219),
    .Q_N(_0008_),
    .Q(\hidden_lif_1.variant_threshold[1] ));
 sg13g2_dfrbp_1 _1575_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net51),
    .D(_0021_),
    .Q_N(_0786_),
    .Q(\hidden_lif_1.variant_threshold[2] ));
 sg13g2_dfrbp_1 _1576_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net49),
    .D(net194),
    .Q_N(_0785_),
    .Q(\hidden_lif_1.variant_threshold[3] ));
 sg13g2_dfrbp_1 _1577_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net47),
    .D(_0023_),
    .Q_N(_0784_),
    .Q(\hidden_lif_1.variant_threshold[4] ));
 sg13g2_dfrbp_1 _1578_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net45),
    .D(_0024_),
    .Q_N(_0783_),
    .Q(\hidden_lif_1.variant_threshold[5] ));
 sg13g2_dfrbp_1 _1579_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net43),
    .D(_0025_),
    .Q_N(_0782_),
    .Q(\hidden_lif_1.variant_threshold[6] ));
 sg13g2_dfrbp_1 _1580_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net41),
    .D(_0026_),
    .Q_N(_0781_),
    .Q(\hidden_lif_1.variant_threshold[7] ));
 sg13g2_dfrbp_1 _1581_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net39),
    .D(net149),
    .Q_N(_0012_),
    .Q(\hidden_lif_2.variant_threshold[1] ));
 sg13g2_dfrbp_1 _1582_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net37),
    .D(_0028_),
    .Q_N(_0780_),
    .Q(\hidden_lif_2.variant_threshold[2] ));
 sg13g2_dfrbp_1 _1583_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net35),
    .D(_0029_),
    .Q_N(_0779_),
    .Q(\hidden_lif_2.variant_threshold[3] ));
 sg13g2_dfrbp_1 _1584_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net33),
    .D(_0030_),
    .Q_N(_0778_),
    .Q(\hidden_lif_2.variant_threshold[4] ));
 sg13g2_dfrbp_1 _1585_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net31),
    .D(_0031_),
    .Q_N(_0777_),
    .Q(\hidden_lif_2.variant_threshold[5] ));
 sg13g2_dfrbp_1 _1586_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net29),
    .D(_0032_),
    .Q_N(_0776_),
    .Q(\hidden_lif_2.variant_threshold[6] ));
 sg13g2_dfrbp_1 _1587_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net27),
    .D(_0033_),
    .Q_N(_0775_),
    .Q(\hidden_lif_2.variant_threshold[7] ));
 sg13g2_dfrbp_1 _1588_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net25),
    .D(net176),
    .Q_N(_0016_),
    .Q(\output_lif_0.variant_threshold[1] ));
 sg13g2_dfrbp_1 _1589_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net134),
    .D(_0035_),
    .Q_N(_0774_),
    .Q(\output_lif_0.variant_threshold[2] ));
 sg13g2_dfrbp_1 _1590_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net132),
    .D(_0036_),
    .Q_N(_0773_),
    .Q(\output_lif_0.variant_threshold[3] ));
 sg13g2_dfrbp_1 _1591_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net130),
    .D(_0037_),
    .Q_N(_0772_),
    .Q(\output_lif_0.variant_threshold[4] ));
 sg13g2_dfrbp_1 _1592_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net128),
    .D(_0038_),
    .Q_N(_0771_),
    .Q(\output_lif_0.variant_threshold[5] ));
 sg13g2_dfrbp_1 _1593_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net126),
    .D(_0039_),
    .Q_N(_0770_),
    .Q(\output_lif_0.variant_threshold[6] ));
 sg13g2_dfrbp_1 _1594_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net124),
    .D(_0040_),
    .Q_N(_0769_),
    .Q(\output_lif_0.variant_threshold[7] ));
 sg13g2_dfrbp_1 _1595_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net122),
    .D(_0041_),
    .Q_N(_0001_),
    .Q(\hidden_lif_2.spike_n ));
 sg13g2_dfrbp_1 _1596_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net121),
    .D(_0042_),
    .Q_N(_0002_),
    .Q(\output_lif_0.spike_n ));
 sg13g2_dfrbp_1 _1597_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net120),
    .D(net141),
    .Q_N(_0768_),
    .Q(\hidden_lif_1.variant_threshold[0] ));
 sg13g2_dfrbp_1 _1598_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net118),
    .D(net209),
    .Q_N(_0767_),
    .Q(\hidden_lif_0.state_r[0] ));
 sg13g2_dfrbp_1 _1599_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net117),
    .D(_0045_),
    .Q_N(_0766_),
    .Q(\hidden_lif_0.state_r[1] ));
 sg13g2_dfrbp_1 _1600_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net116),
    .D(_0046_),
    .Q_N(_0005_),
    .Q(\hidden_lif_0.state_r[2] ));
 sg13g2_dfrbp_1 _1601_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net115),
    .D(_0047_),
    .Q_N(_0765_),
    .Q(\hidden_lif_0.state_r[3] ));
 sg13g2_dfrbp_1 _1602_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net114),
    .D(_0048_),
    .Q_N(_0006_),
    .Q(\hidden_lif_0.state_r[4] ));
 sg13g2_dfrbp_1 _1603_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net113),
    .D(_0049_),
    .Q_N(_0007_),
    .Q(\hidden_lif_0.state_r[5] ));
 sg13g2_dfrbp_1 _1604_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net112),
    .D(_0050_),
    .Q_N(_0764_),
    .Q(\hidden_lif_0.state_r[6] ));
 sg13g2_dfrbp_1 _1605_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net84),
    .D(_0051_),
    .Q_N(_0763_),
    .Q(\hidden_lif_0.state_r[7] ));
 sg13g2_dfrbp_1 _1606_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net83),
    .D(_0052_),
    .Q_N(_0003_),
    .Q(\hidden_lif_0.spike_n ));
 sg13g2_dfrbp_1 _1607_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net82),
    .D(net160),
    .Q_N(_0004_),
    .Q(\hidden_lif_0.variant_threshold[1] ));
 sg13g2_dfrbp_1 _1608_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net80),
    .D(_0054_),
    .Q_N(_0762_),
    .Q(\hidden_lif_0.variant_threshold[2] ));
 sg13g2_dfrbp_1 _1609_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net78),
    .D(_0055_),
    .Q_N(_0761_),
    .Q(\hidden_lif_0.variant_threshold[3] ));
 sg13g2_dfrbp_1 _1610_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net76),
    .D(_0056_),
    .Q_N(_0760_),
    .Q(\hidden_lif_0.variant_threshold[4] ));
 sg13g2_dfrbp_1 _1611_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net74),
    .D(_0057_),
    .Q_N(_0759_),
    .Q(\hidden_lif_0.variant_threshold[5] ));
 sg13g2_dfrbp_1 _1612_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net72),
    .D(_0058_),
    .Q_N(_0758_),
    .Q(\hidden_lif_0.variant_threshold[6] ));
 sg13g2_dfrbp_1 _1613_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net70),
    .D(_0059_),
    .Q_N(_0757_),
    .Q(\hidden_lif_0.variant_threshold[7] ));
 sg13g2_dfrbp_1 _1614_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net68),
    .D(net144),
    .Q_N(_0756_),
    .Q(\hidden_lif_2.variant_threshold[0] ));
 sg13g2_dfrbp_1 _1615_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net66),
    .D(_0061_),
    .Q_N(_0755_),
    .Q(\hidden_lif_1.state_r[0] ));
 sg13g2_dfrbp_1 _1616_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net65),
    .D(_0062_),
    .Q_N(_0754_),
    .Q(\hidden_lif_1.state_r[1] ));
 sg13g2_dfrbp_1 _1617_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net64),
    .D(_0063_),
    .Q_N(_0009_),
    .Q(\hidden_lif_1.state_r[2] ));
 sg13g2_dfrbp_1 _1618_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net63),
    .D(_0064_),
    .Q_N(_0753_),
    .Q(\hidden_lif_1.state_r[3] ));
 sg13g2_dfrbp_1 _1619_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net62),
    .D(_0065_),
    .Q_N(_0010_),
    .Q(\hidden_lif_1.state_r[4] ));
 sg13g2_dfrbp_1 _1620_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net61),
    .D(_0066_),
    .Q_N(_0011_),
    .Q(\hidden_lif_1.state_r[5] ));
 sg13g2_dfrbp_1 _1621_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net60),
    .D(_0067_),
    .Q_N(_0752_),
    .Q(\hidden_lif_1.state_r[6] ));
 sg13g2_dfrbp_1 _1622_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net59),
    .D(_0068_),
    .Q_N(_0751_),
    .Q(\hidden_lif_1.state_r[7] ));
 sg13g2_dfrbp_1 _1623_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net58),
    .D(_0069_),
    .Q_N(_0000_),
    .Q(\hidden_lif_1.spike_n ));
 sg13g2_dfrbp_1 _1624_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net57),
    .D(_0070_),
    .Q_N(_0750_),
    .Q(\output_lif_0.variant_threshold[0] ));
 sg13g2_dfrbp_1 _1625_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net55),
    .D(net217),
    .Q_N(_0749_),
    .Q(\hidden_lif_2.state_r[0] ));
 sg13g2_dfrbp_1 _1626_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net54),
    .D(_0072_),
    .Q_N(_0748_),
    .Q(\hidden_lif_2.state_r[1] ));
 sg13g2_dfrbp_1 _1627_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net53),
    .D(_0073_),
    .Q_N(_0013_),
    .Q(\hidden_lif_2.state_r[2] ));
 sg13g2_dfrbp_1 _1628_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net52),
    .D(net204),
    .Q_N(_0747_),
    .Q(\hidden_lif_2.state_r[3] ));
 sg13g2_dfrbp_1 _1629_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net50),
    .D(_0075_),
    .Q_N(_0014_),
    .Q(\hidden_lif_2.state_r[4] ));
 sg13g2_dfrbp_1 _1630_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net48),
    .D(_0076_),
    .Q_N(_0015_),
    .Q(\hidden_lif_2.state_r[5] ));
 sg13g2_dfrbp_1 _1631_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net46),
    .D(net232),
    .Q_N(_0746_),
    .Q(\hidden_lif_2.state_r[6] ));
 sg13g2_dfrbp_1 _1632_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net44),
    .D(net224),
    .Q_N(_0745_),
    .Q(\hidden_lif_2.state_r[7] ));
 sg13g2_dfrbp_1 _1633_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net42),
    .D(_0079_),
    .Q_N(_0744_),
    .Q(\hidden_weight_0[0] ));
 sg13g2_dfrbp_1 _1634_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net40),
    .D(_0080_),
    .Q_N(_0743_),
    .Q(\hidden_weight_0[1] ));
 sg13g2_dfrbp_1 _1635_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net38),
    .D(_0081_),
    .Q_N(_0742_),
    .Q(\hidden_weight_0[2] ));
 sg13g2_dfrbp_1 _1636_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net36),
    .D(_0082_),
    .Q_N(_0741_),
    .Q(\hidden_weight_1[0] ));
 sg13g2_dfrbp_1 _1637_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net34),
    .D(net157),
    .Q_N(_0740_),
    .Q(\hidden_lif_0.variant_threshold[0] ));
 sg13g2_dfrbp_1 _1638_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net30),
    .D(_0084_),
    .Q_N(_0739_),
    .Q(\output_lif_0.state_r[0] ));
 sg13g2_dfrbp_1 _1639_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net28),
    .D(_0085_),
    .Q_N(_0738_),
    .Q(\output_lif_0.state_r[1] ));
 sg13g2_dfrbp_1 _1640_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net26),
    .D(_0086_),
    .Q_N(_0737_),
    .Q(\output_lif_0.state_r[2] ));
 sg13g2_dfrbp_1 _1641_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net135),
    .D(_0087_),
    .Q_N(_0736_),
    .Q(\output_lif_0.state_r[3] ));
 sg13g2_dfrbp_1 _1642_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net133),
    .D(_0088_),
    .Q_N(_0017_),
    .Q(\output_lif_0.state_r[4] ));
 sg13g2_dfrbp_1 _1643_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net131),
    .D(_0089_),
    .Q_N(_0018_),
    .Q(\output_lif_0.state_r[5] ));
 sg13g2_dfrbp_1 _1644_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net129),
    .D(_0090_),
    .Q_N(_0735_),
    .Q(\output_lif_0.state_r[6] ));
 sg13g2_dfrbp_1 _1645_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net127),
    .D(net182),
    .Q_N(_0734_),
    .Q(\output_lif_0.state_r[7] ));
 sg13g2_dfrbp_1 _1646_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net125),
    .D(_0092_),
    .Q_N(_0733_),
    .Q(\output_weight_0[0] ));
 sg13g2_dfrbp_1 _1647_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net123),
    .D(_0093_),
    .Q_N(_0732_),
    .Q(\output_weight_0[1] ));
 sg13g2_dfrbp_1 _1648_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net119),
    .D(_0094_),
    .Q_N(_0731_),
    .Q(\output_weight_0[2] ));
 sg13g2_dfrbp_1 _1649_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net81),
    .D(_0095_),
    .Q_N(_0730_),
    .Q(\output_weight_1[0] ));
 sg13g2_dfrbp_1 _1650_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net79),
    .D(net137),
    .Q_N(_0019_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _1651_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net75),
    .D(net147),
    .Q_N(_0729_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _1652_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net71),
    .D(_0098_),
    .Q_N(_0728_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _1653_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net67),
    .D(_0099_),
    .Q_N(_0727_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _1654_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net32),
    .D(_0100_),
    .Q_N(_0726_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _1655_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net73),
    .D(net153),
    .Q_N(_0725_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _1656_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net56),
    .D(net226),
    .Q_N(_0724_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _1657_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net69),
    .D(net167),
    .Q_N(_0723_),
    .Q(uo_out[7]));
 sg13g2_tiehi _1640__26 (.L_HI(net26));
 sg13g2_tiehi _1587__27 (.L_HI(net27));
 sg13g2_tiehi _1639__28 (.L_HI(net28));
 sg13g2_tiehi _1586__29 (.L_HI(net29));
 sg13g2_tiehi _1638__30 (.L_HI(net30));
 sg13g2_tiehi _1585__31 (.L_HI(net31));
 sg13g2_tiehi _1654__32 (.L_HI(net32));
 sg13g2_tiehi _1584__33 (.L_HI(net33));
 sg13g2_tiehi _1637__34 (.L_HI(net34));
 sg13g2_tiehi _1583__35 (.L_HI(net35));
 sg13g2_tiehi _1636__36 (.L_HI(net36));
 sg13g2_tiehi _1582__37 (.L_HI(net37));
 sg13g2_tiehi _1635__38 (.L_HI(net38));
 sg13g2_tiehi _1581__39 (.L_HI(net39));
 sg13g2_tiehi _1634__40 (.L_HI(net40));
 sg13g2_tiehi _1580__41 (.L_HI(net41));
 sg13g2_tiehi _1633__42 (.L_HI(net42));
 sg13g2_tiehi _1579__43 (.L_HI(net43));
 sg13g2_tiehi _1632__44 (.L_HI(net44));
 sg13g2_tiehi _1578__45 (.L_HI(net45));
 sg13g2_tiehi _1631__46 (.L_HI(net46));
 sg13g2_tiehi _1577__47 (.L_HI(net47));
 sg13g2_tiehi _1630__48 (.L_HI(net48));
 sg13g2_tiehi _1576__49 (.L_HI(net49));
 sg13g2_tiehi _1629__50 (.L_HI(net50));
 sg13g2_tiehi _1575__51 (.L_HI(net51));
 sg13g2_tiehi _1628__52 (.L_HI(net52));
 sg13g2_tiehi _1627__53 (.L_HI(net53));
 sg13g2_tiehi _1626__54 (.L_HI(net54));
 sg13g2_tiehi _1625__55 (.L_HI(net55));
 sg13g2_tiehi _1656__56 (.L_HI(net56));
 sg13g2_tiehi _1624__57 (.L_HI(net57));
 sg13g2_tiehi _1623__58 (.L_HI(net58));
 sg13g2_tiehi _1622__59 (.L_HI(net59));
 sg13g2_tiehi _1621__60 (.L_HI(net60));
 sg13g2_tiehi _1620__61 (.L_HI(net61));
 sg13g2_tiehi _1619__62 (.L_HI(net62));
 sg13g2_tiehi _1618__63 (.L_HI(net63));
 sg13g2_tiehi _1617__64 (.L_HI(net64));
 sg13g2_tiehi _1616__65 (.L_HI(net65));
 sg13g2_tiehi _1615__66 (.L_HI(net66));
 sg13g2_tiehi _1653__67 (.L_HI(net67));
 sg13g2_tiehi _1614__68 (.L_HI(net68));
 sg13g2_tiehi _1657__69 (.L_HI(net69));
 sg13g2_tiehi _1613__70 (.L_HI(net70));
 sg13g2_tiehi _1652__71 (.L_HI(net71));
 sg13g2_tiehi _1612__72 (.L_HI(net72));
 sg13g2_tiehi _1655__73 (.L_HI(net73));
 sg13g2_tiehi _1611__74 (.L_HI(net74));
 sg13g2_tiehi _1651__75 (.L_HI(net75));
 sg13g2_tiehi _1610__76 (.L_HI(net76));
 sg13g2_tiehi _1574__77 (.L_HI(net77));
 sg13g2_tiehi _1609__78 (.L_HI(net78));
 sg13g2_tiehi _1650__79 (.L_HI(net79));
 sg13g2_tiehi _1608__80 (.L_HI(net80));
 sg13g2_tiehi _1649__81 (.L_HI(net81));
 sg13g2_tiehi _1607__82 (.L_HI(net82));
 sg13g2_tiehi _1606__83 (.L_HI(net83));
 sg13g2_tiehi _1605__84 (.L_HI(net84));
 sg13g2_tiehi _1604__85 (.L_HI(net112));
 sg13g2_tiehi _1603__86 (.L_HI(net113));
 sg13g2_tiehi _1602__87 (.L_HI(net114));
 sg13g2_tiehi _1601__88 (.L_HI(net115));
 sg13g2_tiehi _1600__89 (.L_HI(net116));
 sg13g2_tiehi _1599__90 (.L_HI(net117));
 sg13g2_tiehi _1598__91 (.L_HI(net118));
 sg13g2_tiehi _1648__92 (.L_HI(net119));
 sg13g2_tiehi _1597__93 (.L_HI(net120));
 sg13g2_tiehi _1596__94 (.L_HI(net121));
 sg13g2_tiehi _1595__95 (.L_HI(net122));
 sg13g2_tiehi _1647__96 (.L_HI(net123));
 sg13g2_tiehi _1594__97 (.L_HI(net124));
 sg13g2_tiehi _1646__98 (.L_HI(net125));
 sg13g2_tiehi _1593__99 (.L_HI(net126));
 sg13g2_tiehi _1645__100 (.L_HI(net127));
 sg13g2_tiehi _1592__101 (.L_HI(net128));
 sg13g2_tiehi _1644__102 (.L_HI(net129));
 sg13g2_tiehi _1591__103 (.L_HI(net130));
 sg13g2_tiehi _1643__104 (.L_HI(net131));
 sg13g2_tiehi _1590__105 (.L_HI(net132));
 sg13g2_tiehi _1642__106 (.L_HI(net133));
 sg13g2_tiehi _1589__107 (.L_HI(net134));
 sg13g2_tiehi _1641__108 (.L_HI(net135));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_kailinsley_10 (.L_LO(net10));
 sg13g2_tielo tt_um_kailinsley_11 (.L_LO(net11));
 sg13g2_tielo tt_um_kailinsley_12 (.L_LO(net12));
 sg13g2_tielo tt_um_kailinsley_13 (.L_LO(net13));
 sg13g2_tielo tt_um_kailinsley_14 (.L_LO(net14));
 sg13g2_tielo tt_um_kailinsley_15 (.L_LO(net15));
 sg13g2_tielo tt_um_kailinsley_16 (.L_LO(net16));
 sg13g2_tielo tt_um_kailinsley_17 (.L_LO(net17));
 sg13g2_tielo tt_um_kailinsley_18 (.L_LO(net18));
 sg13g2_tielo tt_um_kailinsley_19 (.L_LO(net19));
 sg13g2_tielo tt_um_kailinsley_20 (.L_LO(net20));
 sg13g2_tielo tt_um_kailinsley_21 (.L_LO(net21));
 sg13g2_tielo tt_um_kailinsley_22 (.L_LO(net22));
 sg13g2_tielo tt_um_kailinsley_23 (.L_LO(net23));
 sg13g2_tielo tt_um_kailinsley_24 (.L_LO(net24));
 sg13g2_tiehi _1588__25 (.L_HI(net25));
 sg13g2_buf_2 fanout85 (.A(net87),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(net87),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_0362_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_0497_),
    .X(net88));
 sg13g2_buf_1 fanout89 (.A(_0497_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_0647_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_0647_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(\output_lif_0.state_r[6] ),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(net199),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(net95),
    .X(net94));
 sg13g2_buf_1 fanout95 (.A(net96),
    .X(net95));
 sg13g2_buf_1 fanout96 (.A(\hidden_weight_0[0] ),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(net98),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(\hidden_lif_1.spike_n ),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(net100),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(\hidden_lif_0.spike_n ),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(net102),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(\output_lif_0.spike_n ),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(\hidden_lif_2.spike_n ),
    .X(net103));
 sg13g2_buf_1 fanout104 (.A(\hidden_lif_2.spike_n ),
    .X(net104));
 sg13g2_buf_4 fanout105 (.X(net105),
    .A(_0139_));
 sg13g2_buf_2 fanout106 (.A(net109),
    .X(net106));
 sg13g2_buf_4 fanout107 (.X(net107),
    .A(net108));
 sg13g2_buf_4 fanout108 (.X(net108),
    .A(net109));
 sg13g2_buf_2 fanout109 (.A(rst_n),
    .X(net109));
 sg13g2_buf_4 fanout110 (.X(net110),
    .A(net111));
 sg13g2_buf_4 fanout111 (.X(net111),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_kailinsley_9 (.L_LO(net9));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0019_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0096_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold3 (.A(\output_weight_0[1] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold4 (.A(\output_weight_0[0] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0000_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0043_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold7 (.A(\output_weight_0[2] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold8 (.A(\hidden_lif_2.variant_threshold[0] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0060_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold10 (.A(uo_out[1]),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0709_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0097_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0001_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0027_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold15 (.A(\hidden_weight_0[2] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold16 (.A(uo_out[5]),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0717_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0101_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0017_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold20 (.A(\output_weight_1[0] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0003_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0083_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0004_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0437_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0053_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0007_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0414_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold28 (.A(uo_out[3]),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0714_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold30 (.A(\hidden_lif_0.variant_threshold[2] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold31 (.A(uo_out[7]),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0103_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold33 (.A(\hidden_lif_0.variant_threshold[3] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0011_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0555_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold36 (.A(\output_lif_0.variant_threshold[2] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0259_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold38 (.A(\hidden_lif_2.variant_threshold[7] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0243_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0002_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0034_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0015_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0616_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold44 (.A(\output_lif_0.variant_threshold[7] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold45 (.A(\output_lif_0.state_r[7] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0706_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0091_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold48 (.A(\hidden_weight_0[1] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0010_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold50 (.A(\hidden_lif_2.variant_threshold[3] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold51 (.A(\output_lif_0.variant_threshold[3] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold52 (.A(\hidden_lif_0.variant_threshold[4] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold53 (.A(\output_lif_0.variant_threshold[0] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold54 (.A(\hidden_lif_2.variant_threshold[2] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold55 (.A(\hidden_lif_1.state_r[7] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold56 (.A(\hidden_lif_1.variant_threshold[4] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0006_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold58 (.A(\hidden_lif_1.variant_threshold[3] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0022_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold60 (.A(\hidden_lif_1.variant_threshold[6] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0201_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold62 (.A(\hidden_lif_0.state_r[7] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0429_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold64 (.A(\hidden_weight_1[0] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold65 (.A(\hidden_lif_2.variant_threshold[6] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0241_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold67 (.A(uo_out[4]),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0014_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0074_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0018_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0689_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold72 (.A(\hidden_lif_0.state_r[0] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0365_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0044_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold75 (.A(\hidden_lif_0.variant_threshold[7] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0376_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold77 (.A(\hidden_lif_1.variant_threshold[2] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold78 (.A(\hidden_lif_1.variant_threshold[7] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold79 (.A(\hidden_lif_1.variant_threshold[5] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold80 (.A(\hidden_lif_2.state_r[0] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0575_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0071_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold83 (.A(\hidden_lif_1.variant_threshold[1] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0020_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold85 (.A(uo_out[2]),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0712_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold87 (.A(\hidden_lif_2.state_r[6] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0619_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0078_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold90 (.A(uo_out[6]),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0102_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold92 (.A(\hidden_lif_0.variant_threshold[6] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold93 (.A(\hidden_lif_0.variant_threshold[6] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0432_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold95 (.A(\hidden_lif_0.variant_threshold[5] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold96 (.A(\hidden_lif_2.state_r[7] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0077_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold98 (.A(\hidden_lif_2.variant_threshold[4] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold99 (.A(\hidden_lif_2.variant_threshold[5] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold100 (.A(\output_lif_0.state_r[0] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold101 (.A(\output_lif_0.variant_threshold[6] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold102 (.A(\output_lif_0.variant_threshold[5] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0274_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold104 (.A(\output_lif_0.state_r[7] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0299_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold106 (.A(\hidden_lif_1.state_r[0] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0520_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold108 (.A(\output_lif_0.variant_threshold[4] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold109 (.A(\hidden_lif_1.variant_threshold[6] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold110 (.A(\hidden_lif_1.state_r[6] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold111 (.A(\hidden_lif_1.state_r[5] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0563_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold113 (.A(\output_lif_0.state_r[5] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold114 (.A(\hidden_lif_2.state_r[1] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold115 (.A(\hidden_lif_0.state_r[5] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0421_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold117 (.A(\hidden_lif_0.state_r[1] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold118 (.A(\hidden_lif_1.variant_threshold[1] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold119 (.A(\hidden_lif_1.state_r[0] ),
    .X(net254));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_4 FILLER_12_322 ();
 sg13g2_fill_1 FILLER_12_326 ();
 sg13g2_decap_8 FILLER_12_331 ();
 sg13g2_decap_8 FILLER_12_338 ();
 sg13g2_decap_8 FILLER_12_345 ();
 sg13g2_fill_1 FILLER_12_352 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_fill_2 FILLER_13_140 ();
 sg13g2_fill_1 FILLER_13_142 ();
 sg13g2_fill_2 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_153 ();
 sg13g2_decap_8 FILLER_13_160 ();
 sg13g2_decap_4 FILLER_13_167 ();
 sg13g2_fill_1 FILLER_13_171 ();
 sg13g2_decap_8 FILLER_13_176 ();
 sg13g2_decap_8 FILLER_13_183 ();
 sg13g2_decap_4 FILLER_13_190 ();
 sg13g2_decap_8 FILLER_13_197 ();
 sg13g2_fill_2 FILLER_13_204 ();
 sg13g2_decap_4 FILLER_13_237 ();
 sg13g2_fill_1 FILLER_13_241 ();
 sg13g2_decap_8 FILLER_13_251 ();
 sg13g2_decap_8 FILLER_13_258 ();
 sg13g2_decap_8 FILLER_13_265 ();
 sg13g2_decap_8 FILLER_13_272 ();
 sg13g2_decap_8 FILLER_13_279 ();
 sg13g2_fill_2 FILLER_13_286 ();
 sg13g2_fill_1 FILLER_13_288 ();
 sg13g2_fill_1 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_368 ();
 sg13g2_decap_8 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_4 FILLER_13_403 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_4 FILLER_14_133 ();
 sg13g2_fill_1 FILLER_14_137 ();
 sg13g2_decap_4 FILLER_14_164 ();
 sg13g2_decap_4 FILLER_14_205 ();
 sg13g2_decap_8 FILLER_14_257 ();
 sg13g2_decap_8 FILLER_14_264 ();
 sg13g2_decap_8 FILLER_14_271 ();
 sg13g2_fill_2 FILLER_14_278 ();
 sg13g2_fill_1 FILLER_14_280 ();
 sg13g2_fill_2 FILLER_14_285 ();
 sg13g2_fill_1 FILLER_14_287 ();
 sg13g2_fill_2 FILLER_14_323 ();
 sg13g2_fill_1 FILLER_14_325 ();
 sg13g2_fill_1 FILLER_14_354 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_4 FILLER_15_77 ();
 sg13g2_fill_2 FILLER_15_81 ();
 sg13g2_decap_8 FILLER_15_87 ();
 sg13g2_decap_8 FILLER_15_94 ();
 sg13g2_decap_8 FILLER_15_101 ();
 sg13g2_decap_8 FILLER_15_108 ();
 sg13g2_fill_2 FILLER_15_115 ();
 sg13g2_fill_2 FILLER_15_147 ();
 sg13g2_fill_2 FILLER_15_178 ();
 sg13g2_fill_2 FILLER_15_193 ();
 sg13g2_fill_1 FILLER_15_195 ();
 sg13g2_fill_2 FILLER_15_207 ();
 sg13g2_fill_2 FILLER_15_217 ();
 sg13g2_decap_4 FILLER_15_228 ();
 sg13g2_fill_1 FILLER_15_269 ();
 sg13g2_fill_1 FILLER_15_331 ();
 sg13g2_fill_2 FILLER_15_348 ();
 sg13g2_fill_1 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_368 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_fill_2 FILLER_15_386 ();
 sg13g2_fill_1 FILLER_15_388 ();
 sg13g2_fill_2 FILLER_15_392 ();
 sg13g2_fill_2 FILLER_15_398 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_4 FILLER_16_49 ();
 sg13g2_fill_2 FILLER_16_53 ();
 sg13g2_decap_8 FILLER_16_59 ();
 sg13g2_decap_8 FILLER_16_66 ();
 sg13g2_decap_8 FILLER_16_108 ();
 sg13g2_fill_2 FILLER_16_115 ();
 sg13g2_decap_4 FILLER_16_121 ();
 sg13g2_fill_1 FILLER_16_125 ();
 sg13g2_fill_2 FILLER_16_140 ();
 sg13g2_fill_1 FILLER_16_142 ();
 sg13g2_fill_2 FILLER_16_169 ();
 sg13g2_fill_1 FILLER_16_171 ();
 sg13g2_fill_1 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_201 ();
 sg13g2_decap_4 FILLER_16_208 ();
 sg13g2_fill_2 FILLER_16_225 ();
 sg13g2_fill_1 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_276 ();
 sg13g2_decap_4 FILLER_16_283 ();
 sg13g2_fill_1 FILLER_16_287 ();
 sg13g2_fill_2 FILLER_16_307 ();
 sg13g2_fill_1 FILLER_16_309 ();
 sg13g2_fill_2 FILLER_16_326 ();
 sg13g2_fill_2 FILLER_16_342 ();
 sg13g2_fill_1 FILLER_16_349 ();
 sg13g2_fill_1 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_fill_2 FILLER_17_42 ();
 sg13g2_fill_1 FILLER_17_105 ();
 sg13g2_fill_2 FILLER_17_132 ();
 sg13g2_fill_1 FILLER_17_134 ();
 sg13g2_fill_1 FILLER_17_185 ();
 sg13g2_decap_8 FILLER_17_197 ();
 sg13g2_fill_2 FILLER_17_212 ();
 sg13g2_fill_2 FILLER_17_241 ();
 sg13g2_fill_1 FILLER_17_259 ();
 sg13g2_decap_4 FILLER_17_357 ();
 sg13g2_fill_2 FILLER_17_361 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_4 FILLER_18_42 ();
 sg13g2_fill_2 FILLER_18_46 ();
 sg13g2_decap_8 FILLER_18_109 ();
 sg13g2_fill_1 FILLER_18_116 ();
 sg13g2_decap_4 FILLER_18_130 ();
 sg13g2_fill_1 FILLER_18_134 ();
 sg13g2_fill_1 FILLER_18_159 ();
 sg13g2_decap_8 FILLER_18_173 ();
 sg13g2_decap_8 FILLER_18_187 ();
 sg13g2_fill_2 FILLER_18_194 ();
 sg13g2_decap_4 FILLER_18_199 ();
 sg13g2_fill_2 FILLER_18_207 ();
 sg13g2_fill_2 FILLER_18_231 ();
 sg13g2_fill_1 FILLER_18_233 ();
 sg13g2_fill_1 FILLER_18_247 ();
 sg13g2_fill_2 FILLER_18_262 ();
 sg13g2_fill_1 FILLER_18_281 ();
 sg13g2_decap_8 FILLER_18_290 ();
 sg13g2_fill_2 FILLER_18_297 ();
 sg13g2_decap_4 FILLER_18_309 ();
 sg13g2_decap_4 FILLER_18_350 ();
 sg13g2_fill_2 FILLER_18_365 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_4 FILLER_19_69 ();
 sg13g2_fill_1 FILLER_19_73 ();
 sg13g2_fill_2 FILLER_19_79 ();
 sg13g2_fill_1 FILLER_19_81 ();
 sg13g2_fill_2 FILLER_19_86 ();
 sg13g2_fill_1 FILLER_19_88 ();
 sg13g2_decap_4 FILLER_19_101 ();
 sg13g2_fill_2 FILLER_19_105 ();
 sg13g2_fill_1 FILLER_19_155 ();
 sg13g2_fill_2 FILLER_19_177 ();
 sg13g2_fill_1 FILLER_19_199 ();
 sg13g2_fill_1 FILLER_19_212 ();
 sg13g2_fill_1 FILLER_19_218 ();
 sg13g2_fill_2 FILLER_19_226 ();
 sg13g2_fill_1 FILLER_19_228 ();
 sg13g2_fill_2 FILLER_19_234 ();
 sg13g2_fill_1 FILLER_19_236 ();
 sg13g2_fill_1 FILLER_19_251 ();
 sg13g2_fill_1 FILLER_19_322 ();
 sg13g2_fill_2 FILLER_19_337 ();
 sg13g2_fill_1 FILLER_19_354 ();
 sg13g2_fill_2 FILLER_19_362 ();
 sg13g2_fill_2 FILLER_19_372 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_33 ();
 sg13g2_decap_4 FILLER_20_49 ();
 sg13g2_fill_2 FILLER_20_53 ();
 sg13g2_fill_2 FILLER_20_81 ();
 sg13g2_decap_8 FILLER_20_107 ();
 sg13g2_decap_8 FILLER_20_118 ();
 sg13g2_fill_1 FILLER_20_125 ();
 sg13g2_fill_2 FILLER_20_150 ();
 sg13g2_fill_1 FILLER_20_157 ();
 sg13g2_fill_2 FILLER_20_180 ();
 sg13g2_fill_1 FILLER_20_185 ();
 sg13g2_fill_2 FILLER_20_194 ();
 sg13g2_decap_8 FILLER_20_202 ();
 sg13g2_fill_1 FILLER_20_209 ();
 sg13g2_decap_8 FILLER_20_218 ();
 sg13g2_fill_1 FILLER_20_225 ();
 sg13g2_fill_2 FILLER_20_278 ();
 sg13g2_fill_1 FILLER_20_280 ();
 sg13g2_fill_1 FILLER_20_290 ();
 sg13g2_fill_2 FILLER_20_308 ();
 sg13g2_fill_1 FILLER_20_328 ();
 sg13g2_fill_1 FILLER_20_339 ();
 sg13g2_fill_1 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_4 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_22 ();
 sg13g2_fill_2 FILLER_21_29 ();
 sg13g2_fill_2 FILLER_21_60 ();
 sg13g2_fill_1 FILLER_21_62 ();
 sg13g2_decap_8 FILLER_21_76 ();
 sg13g2_fill_1 FILLER_21_83 ();
 sg13g2_fill_2 FILLER_21_96 ();
 sg13g2_decap_4 FILLER_21_129 ();
 sg13g2_fill_1 FILLER_21_133 ();
 sg13g2_fill_2 FILLER_21_150 ();
 sg13g2_fill_2 FILLER_21_199 ();
 sg13g2_fill_1 FILLER_21_201 ();
 sg13g2_decap_4 FILLER_21_231 ();
 sg13g2_fill_2 FILLER_21_239 ();
 sg13g2_fill_2 FILLER_21_262 ();
 sg13g2_fill_1 FILLER_21_320 ();
 sg13g2_fill_2 FILLER_21_347 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_4 ();
 sg13g2_decap_4 FILLER_22_78 ();
 sg13g2_decap_8 FILLER_22_108 ();
 sg13g2_fill_2 FILLER_22_115 ();
 sg13g2_fill_1 FILLER_22_161 ();
 sg13g2_fill_1 FILLER_22_171 ();
 sg13g2_decap_4 FILLER_22_203 ();
 sg13g2_fill_2 FILLER_22_215 ();
 sg13g2_decap_4 FILLER_22_241 ();
 sg13g2_fill_2 FILLER_22_245 ();
 sg13g2_fill_2 FILLER_22_289 ();
 sg13g2_fill_1 FILLER_22_291 ();
 sg13g2_fill_2 FILLER_22_314 ();
 sg13g2_fill_1 FILLER_22_316 ();
 sg13g2_fill_2 FILLER_22_321 ();
 sg13g2_fill_1 FILLER_22_330 ();
 sg13g2_decap_8 FILLER_22_386 ();
 sg13g2_decap_8 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_14 ();
 sg13g2_fill_2 FILLER_23_54 ();
 sg13g2_fill_1 FILLER_23_56 ();
 sg13g2_decap_4 FILLER_23_69 ();
 sg13g2_fill_1 FILLER_23_73 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_fill_1 FILLER_23_126 ();
 sg13g2_decap_4 FILLER_23_131 ();
 sg13g2_fill_2 FILLER_23_190 ();
 sg13g2_fill_2 FILLER_23_218 ();
 sg13g2_fill_1 FILLER_23_220 ();
 sg13g2_decap_4 FILLER_23_225 ();
 sg13g2_fill_2 FILLER_23_234 ();
 sg13g2_fill_1 FILLER_23_236 ();
 sg13g2_decap_4 FILLER_23_241 ();
 sg13g2_fill_1 FILLER_23_245 ();
 sg13g2_fill_1 FILLER_23_255 ();
 sg13g2_fill_2 FILLER_23_271 ();
 sg13g2_fill_1 FILLER_23_273 ();
 sg13g2_fill_1 FILLER_23_306 ();
 sg13g2_fill_2 FILLER_23_327 ();
 sg13g2_fill_1 FILLER_23_329 ();
 sg13g2_fill_1 FILLER_23_338 ();
 sg13g2_fill_1 FILLER_23_369 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_fill_1 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_fill_1 FILLER_24_91 ();
 sg13g2_fill_2 FILLER_24_106 ();
 sg13g2_fill_1 FILLER_24_108 ();
 sg13g2_decap_8 FILLER_24_135 ();
 sg13g2_fill_2 FILLER_24_142 ();
 sg13g2_fill_1 FILLER_24_144 ();
 sg13g2_fill_2 FILLER_24_154 ();
 sg13g2_fill_1 FILLER_24_156 ();
 sg13g2_fill_1 FILLER_24_162 ();
 sg13g2_fill_2 FILLER_24_172 ();
 sg13g2_fill_1 FILLER_24_174 ();
 sg13g2_decap_8 FILLER_24_179 ();
 sg13g2_fill_2 FILLER_24_186 ();
 sg13g2_fill_1 FILLER_24_188 ();
 sg13g2_decap_8 FILLER_24_193 ();
 sg13g2_fill_2 FILLER_24_200 ();
 sg13g2_fill_1 FILLER_24_202 ();
 sg13g2_decap_4 FILLER_24_207 ();
 sg13g2_fill_1 FILLER_24_211 ();
 sg13g2_decap_8 FILLER_24_216 ();
 sg13g2_fill_2 FILLER_24_223 ();
 sg13g2_fill_1 FILLER_24_225 ();
 sg13g2_fill_2 FILLER_24_252 ();
 sg13g2_fill_1 FILLER_24_254 ();
 sg13g2_fill_1 FILLER_24_276 ();
 sg13g2_decap_8 FILLER_24_282 ();
 sg13g2_fill_1 FILLER_24_289 ();
 sg13g2_decap_4 FILLER_24_302 ();
 sg13g2_fill_1 FILLER_24_306 ();
 sg13g2_fill_2 FILLER_24_312 ();
 sg13g2_fill_1 FILLER_24_314 ();
 sg13g2_fill_2 FILLER_24_320 ();
 sg13g2_decap_4 FILLER_24_337 ();
 sg13g2_fill_2 FILLER_24_346 ();
 sg13g2_fill_1 FILLER_24_359 ();
 sg13g2_fill_2 FILLER_24_374 ();
 sg13g2_fill_1 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_24_386 ();
 sg13g2_fill_1 FILLER_24_393 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_9 ();
 sg13g2_fill_2 FILLER_25_22 ();
 sg13g2_fill_1 FILLER_25_75 ();
 sg13g2_decap_4 FILLER_25_79 ();
 sg13g2_fill_2 FILLER_25_83 ();
 sg13g2_decap_4 FILLER_25_109 ();
 sg13g2_fill_1 FILLER_25_113 ();
 sg13g2_fill_1 FILLER_25_123 ();
 sg13g2_decap_8 FILLER_25_158 ();
 sg13g2_decap_4 FILLER_25_165 ();
 sg13g2_fill_2 FILLER_25_169 ();
 sg13g2_fill_2 FILLER_25_175 ();
 sg13g2_fill_2 FILLER_25_194 ();
 sg13g2_fill_1 FILLER_25_240 ();
 sg13g2_fill_1 FILLER_25_262 ();
 sg13g2_fill_2 FILLER_25_280 ();
 sg13g2_fill_1 FILLER_25_282 ();
 sg13g2_fill_1 FILLER_25_297 ();
 sg13g2_fill_2 FILLER_25_313 ();
 sg13g2_fill_1 FILLER_25_315 ();
 sg13g2_fill_1 FILLER_25_342 ();
 sg13g2_decap_8 FILLER_25_348 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_fill_2 FILLER_26_26 ();
 sg13g2_decap_4 FILLER_26_54 ();
 sg13g2_fill_2 FILLER_26_58 ();
 sg13g2_decap_4 FILLER_26_66 ();
 sg13g2_fill_2 FILLER_26_88 ();
 sg13g2_fill_2 FILLER_26_98 ();
 sg13g2_fill_1 FILLER_26_100 ();
 sg13g2_fill_2 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_fill_1 FILLER_26_140 ();
 sg13g2_decap_4 FILLER_26_153 ();
 sg13g2_fill_2 FILLER_26_187 ();
 sg13g2_fill_1 FILLER_26_189 ();
 sg13g2_fill_2 FILLER_26_233 ();
 sg13g2_decap_8 FILLER_26_261 ();
 sg13g2_decap_8 FILLER_26_268 ();
 sg13g2_fill_1 FILLER_26_280 ();
 sg13g2_fill_2 FILLER_26_296 ();
 sg13g2_fill_1 FILLER_26_298 ();
 sg13g2_fill_2 FILLER_26_309 ();
 sg13g2_fill_1 FILLER_26_311 ();
 sg13g2_decap_8 FILLER_26_333 ();
 sg13g2_fill_1 FILLER_26_340 ();
 sg13g2_decap_8 FILLER_26_376 ();
 sg13g2_decap_8 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_42 ();
 sg13g2_decap_4 FILLER_27_62 ();
 sg13g2_fill_2 FILLER_27_74 ();
 sg13g2_decap_4 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_102 ();
 sg13g2_decap_4 FILLER_27_109 ();
 sg13g2_fill_2 FILLER_27_139 ();
 sg13g2_fill_1 FILLER_27_141 ();
 sg13g2_fill_2 FILLER_27_176 ();
 sg13g2_fill_1 FILLER_27_178 ();
 sg13g2_fill_2 FILLER_27_188 ();
 sg13g2_fill_1 FILLER_27_214 ();
 sg13g2_fill_2 FILLER_27_225 ();
 sg13g2_fill_1 FILLER_27_227 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_fill_1 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_272 ();
 sg13g2_decap_4 FILLER_27_299 ();
 sg13g2_fill_2 FILLER_27_303 ();
 sg13g2_decap_4 FILLER_27_331 ();
 sg13g2_fill_1 FILLER_27_335 ();
 sg13g2_decap_8 FILLER_27_344 ();
 sg13g2_fill_1 FILLER_27_351 ();
 sg13g2_fill_2 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_370 ();
 sg13g2_decap_8 FILLER_27_377 ();
 sg13g2_decap_8 FILLER_27_384 ();
 sg13g2_decap_8 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_fill_2 FILLER_28_16 ();
 sg13g2_fill_1 FILLER_28_27 ();
 sg13g2_fill_1 FILLER_28_63 ();
 sg13g2_decap_4 FILLER_28_75 ();
 sg13g2_fill_1 FILLER_28_79 ();
 sg13g2_fill_2 FILLER_28_84 ();
 sg13g2_fill_1 FILLER_28_98 ();
 sg13g2_fill_2 FILLER_28_108 ();
 sg13g2_decap_8 FILLER_28_136 ();
 sg13g2_decap_8 FILLER_28_143 ();
 sg13g2_decap_4 FILLER_28_150 ();
 sg13g2_fill_2 FILLER_28_190 ();
 sg13g2_fill_1 FILLER_28_192 ();
 sg13g2_decap_4 FILLER_28_216 ();
 sg13g2_fill_1 FILLER_28_220 ();
 sg13g2_fill_1 FILLER_28_230 ();
 sg13g2_decap_4 FILLER_28_253 ();
 sg13g2_fill_2 FILLER_28_261 ();
 sg13g2_fill_1 FILLER_28_263 ();
 sg13g2_decap_8 FILLER_28_269 ();
 sg13g2_decap_8 FILLER_28_276 ();
 sg13g2_fill_1 FILLER_28_290 ();
 sg13g2_decap_8 FILLER_28_317 ();
 sg13g2_fill_2 FILLER_28_324 ();
 sg13g2_fill_1 FILLER_28_326 ();
 sg13g2_decap_8 FILLER_28_385 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_fill_2 FILLER_29_64 ();
 sg13g2_fill_1 FILLER_29_91 ();
 sg13g2_decap_4 FILLER_29_97 ();
 sg13g2_fill_2 FILLER_29_109 ();
 sg13g2_fill_1 FILLER_29_111 ();
 sg13g2_fill_2 FILLER_29_121 ();
 sg13g2_fill_1 FILLER_29_123 ();
 sg13g2_fill_2 FILLER_29_160 ();
 sg13g2_fill_2 FILLER_29_185 ();
 sg13g2_fill_2 FILLER_29_198 ();
 sg13g2_fill_1 FILLER_29_200 ();
 sg13g2_fill_1 FILLER_29_206 ();
 sg13g2_fill_2 FILLER_29_211 ();
 sg13g2_fill_1 FILLER_29_213 ();
 sg13g2_fill_1 FILLER_29_222 ();
 sg13g2_fill_1 FILLER_29_228 ();
 sg13g2_fill_1 FILLER_29_258 ();
 sg13g2_fill_1 FILLER_29_283 ();
 sg13g2_decap_8 FILLER_29_319 ();
 sg13g2_fill_2 FILLER_29_326 ();
 sg13g2_fill_1 FILLER_29_328 ();
 sg13g2_fill_2 FILLER_29_352 ();
 sg13g2_decap_8 FILLER_29_369 ();
 sg13g2_decap_4 FILLER_29_376 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_9 ();
 sg13g2_fill_2 FILLER_30_51 ();
 sg13g2_fill_1 FILLER_30_103 ();
 sg13g2_fill_2 FILLER_30_149 ();
 sg13g2_fill_1 FILLER_30_151 ();
 sg13g2_fill_1 FILLER_30_186 ();
 sg13g2_fill_2 FILLER_30_218 ();
 sg13g2_decap_8 FILLER_30_223 ();
 sg13g2_fill_2 FILLER_30_258 ();
 sg13g2_fill_2 FILLER_30_269 ();
 sg13g2_fill_1 FILLER_30_284 ();
 sg13g2_fill_2 FILLER_30_328 ();
 sg13g2_decap_4 FILLER_30_370 ();
 sg13g2_fill_2 FILLER_30_374 ();
 sg13g2_fill_2 FILLER_30_381 ();
 sg13g2_fill_1 FILLER_30_383 ();
 sg13g2_fill_1 FILLER_30_388 ();
 sg13g2_decap_8 FILLER_30_398 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_7 ();
 sg13g2_decap_4 FILLER_31_82 ();
 sg13g2_fill_1 FILLER_31_86 ();
 sg13g2_fill_2 FILLER_31_125 ();
 sg13g2_fill_1 FILLER_31_127 ();
 sg13g2_decap_4 FILLER_31_141 ();
 sg13g2_decap_8 FILLER_31_149 ();
 sg13g2_decap_8 FILLER_31_156 ();
 sg13g2_fill_2 FILLER_31_163 ();
 sg13g2_fill_2 FILLER_31_190 ();
 sg13g2_fill_1 FILLER_31_192 ();
 sg13g2_fill_1 FILLER_31_236 ();
 sg13g2_fill_2 FILLER_31_247 ();
 sg13g2_fill_1 FILLER_31_266 ();
 sg13g2_fill_2 FILLER_31_277 ();
 sg13g2_fill_1 FILLER_31_279 ();
 sg13g2_decap_8 FILLER_31_284 ();
 sg13g2_fill_2 FILLER_31_291 ();
 sg13g2_fill_1 FILLER_31_293 ();
 sg13g2_decap_8 FILLER_31_309 ();
 sg13g2_fill_1 FILLER_31_321 ();
 sg13g2_fill_1 FILLER_31_332 ();
 sg13g2_fill_2 FILLER_31_337 ();
 sg13g2_fill_1 FILLER_31_339 ();
 sg13g2_fill_2 FILLER_31_344 ();
 sg13g2_fill_1 FILLER_31_346 ();
 sg13g2_fill_2 FILLER_31_355 ();
 sg13g2_fill_1 FILLER_31_362 ();
 sg13g2_fill_2 FILLER_31_380 ();
 sg13g2_fill_1 FILLER_31_382 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_fill_2 FILLER_32_28 ();
 sg13g2_fill_1 FILLER_32_30 ();
 sg13g2_fill_2 FILLER_32_57 ();
 sg13g2_fill_1 FILLER_32_59 ();
 sg13g2_fill_2 FILLER_32_70 ();
 sg13g2_fill_1 FILLER_32_72 ();
 sg13g2_fill_1 FILLER_32_99 ();
 sg13g2_fill_1 FILLER_32_150 ();
 sg13g2_fill_2 FILLER_32_177 ();
 sg13g2_fill_1 FILLER_32_205 ();
 sg13g2_decap_4 FILLER_32_226 ();
 sg13g2_fill_1 FILLER_32_230 ();
 sg13g2_fill_2 FILLER_32_253 ();
 sg13g2_fill_2 FILLER_32_268 ();
 sg13g2_fill_2 FILLER_32_277 ();
 sg13g2_decap_8 FILLER_32_318 ();
 sg13g2_decap_4 FILLER_32_325 ();
 sg13g2_decap_4 FILLER_32_379 ();
 sg13g2_fill_1 FILLER_32_383 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_46 ();
 sg13g2_decap_8 FILLER_33_53 ();
 sg13g2_decap_4 FILLER_33_60 ();
 sg13g2_fill_2 FILLER_33_64 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_88 ();
 sg13g2_decap_8 FILLER_33_124 ();
 sg13g2_fill_1 FILLER_33_131 ();
 sg13g2_decap_8 FILLER_33_141 ();
 sg13g2_fill_2 FILLER_33_148 ();
 sg13g2_fill_1 FILLER_33_162 ();
 sg13g2_decap_8 FILLER_33_201 ();
 sg13g2_fill_1 FILLER_33_208 ();
 sg13g2_fill_1 FILLER_33_214 ();
 sg13g2_fill_2 FILLER_33_223 ();
 sg13g2_fill_1 FILLER_33_225 ();
 sg13g2_fill_1 FILLER_33_248 ();
 sg13g2_decap_8 FILLER_33_273 ();
 sg13g2_decap_4 FILLER_33_280 ();
 sg13g2_fill_2 FILLER_33_284 ();
 sg13g2_fill_2 FILLER_33_306 ();
 sg13g2_fill_1 FILLER_33_308 ();
 sg13g2_decap_8 FILLER_33_326 ();
 sg13g2_decap_8 FILLER_33_333 ();
 sg13g2_decap_8 FILLER_33_340 ();
 sg13g2_fill_2 FILLER_33_347 ();
 sg13g2_fill_2 FILLER_33_374 ();
 sg13g2_fill_1 FILLER_33_376 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_fill_2 FILLER_34_126 ();
 sg13g2_fill_1 FILLER_34_128 ();
 sg13g2_fill_2 FILLER_34_204 ();
 sg13g2_fill_1 FILLER_34_206 ();
 sg13g2_decap_4 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_327 ();
 sg13g2_decap_4 FILLER_34_334 ();
 sg13g2_fill_1 FILLER_34_343 ();
 sg13g2_fill_2 FILLER_34_351 ();
 sg13g2_fill_1 FILLER_34_361 ();
 sg13g2_fill_2 FILLER_34_371 ();
 sg13g2_fill_1 FILLER_34_373 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_4 FILLER_35_112 ();
 sg13g2_fill_2 FILLER_35_116 ();
 sg13g2_fill_2 FILLER_35_149 ();
 sg13g2_fill_1 FILLER_35_151 ();
 sg13g2_fill_1 FILLER_35_184 ();
 sg13g2_decap_4 FILLER_35_202 ();
 sg13g2_fill_2 FILLER_35_206 ();
 sg13g2_fill_2 FILLER_35_283 ();
 sg13g2_fill_1 FILLER_35_285 ();
 sg13g2_decap_4 FILLER_35_321 ();
 sg13g2_fill_2 FILLER_35_325 ();
 sg13g2_decap_4 FILLER_35_339 ();
 sg13g2_decap_4 FILLER_35_372 ();
 sg13g2_fill_2 FILLER_35_376 ();
 sg13g2_fill_2 FILLER_35_392 ();
 sg13g2_fill_1 FILLER_35_394 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_fill_2 FILLER_36_126 ();
 sg13g2_fill_2 FILLER_36_132 ();
 sg13g2_fill_1 FILLER_36_150 ();
 sg13g2_fill_1 FILLER_36_196 ();
 sg13g2_fill_2 FILLER_36_254 ();
 sg13g2_fill_1 FILLER_36_279 ();
 sg13g2_fill_2 FILLER_36_289 ();
 sg13g2_fill_2 FILLER_36_337 ();
 sg13g2_fill_2 FILLER_36_348 ();
 sg13g2_decap_4 FILLER_36_356 ();
 sg13g2_fill_2 FILLER_36_373 ();
 sg13g2_fill_1 FILLER_36_375 ();
 sg13g2_fill_2 FILLER_36_381 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_4 FILLER_37_126 ();
 sg13g2_fill_2 FILLER_37_130 ();
 sg13g2_fill_2 FILLER_37_186 ();
 sg13g2_fill_1 FILLER_37_213 ();
 sg13g2_fill_2 FILLER_37_267 ();
 sg13g2_fill_2 FILLER_37_283 ();
 sg13g2_fill_1 FILLER_37_307 ();
 sg13g2_fill_2 FILLER_37_333 ();
 sg13g2_fill_1 FILLER_37_335 ();
 sg13g2_fill_2 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_fill_1 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_fill_1 FILLER_38_124 ();
 sg13g2_fill_1 FILLER_38_232 ();
 sg13g2_fill_2 FILLER_38_246 ();
 sg13g2_fill_1 FILLER_38_330 ();
 sg13g2_decap_8 FILLER_38_398 ();
 sg13g2_decap_4 FILLER_38_405 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule

module tt_um_synth_simple_mm (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire pwm_out_i;
 wire pwm_out_right;
 wire \sm_i.adsr_i.dout[0] ;
 wire \sm_i.adsr_i.dout[1] ;
 wire \sm_i.adsr_i.dout[2] ;
 wire \sm_i.adsr_i.dout[3] ;
 wire \sm_i.adsr_i.dout[4] ;
 wire \sm_i.adsr_i.dout[5] ;
 wire \sm_i.adsr_i.scnt_pwl[0] ;
 wire \sm_i.adsr_i.scnt_pwl[1] ;
 wire \sm_i.adsr_i.scnt_pwl[2] ;
 wire \sm_i.adsr_i.scnt_step[0] ;
 wire \sm_i.adsr_i.scnt_step[10] ;
 wire \sm_i.adsr_i.scnt_step[11] ;
 wire \sm_i.adsr_i.scnt_step[12] ;
 wire \sm_i.adsr_i.scnt_step[13] ;
 wire \sm_i.adsr_i.scnt_step[14] ;
 wire \sm_i.adsr_i.scnt_step[15] ;
 wire \sm_i.adsr_i.scnt_step[16] ;
 wire \sm_i.adsr_i.scnt_step[17] ;
 wire \sm_i.adsr_i.scnt_step[18] ;
 wire \sm_i.adsr_i.scnt_step[19] ;
 wire \sm_i.adsr_i.scnt_step[1] ;
 wire \sm_i.adsr_i.scnt_step[20] ;
 wire \sm_i.adsr_i.scnt_step[21] ;
 wire \sm_i.adsr_i.scnt_step[22] ;
 wire \sm_i.adsr_i.scnt_step[23] ;
 wire \sm_i.adsr_i.scnt_step[24] ;
 wire \sm_i.adsr_i.scnt_step[25] ;
 wire \sm_i.adsr_i.scnt_step[26] ;
 wire \sm_i.adsr_i.scnt_step[27] ;
 wire \sm_i.adsr_i.scnt_step[2] ;
 wire \sm_i.adsr_i.scnt_step[3] ;
 wire \sm_i.adsr_i.scnt_step[4] ;
 wire \sm_i.adsr_i.scnt_step[5] ;
 wire \sm_i.adsr_i.scnt_step[6] ;
 wire \sm_i.adsr_i.scnt_step[7] ;
 wire \sm_i.adsr_i.scnt_step[8] ;
 wire \sm_i.adsr_i.scnt_step[9] ;
 wire \sm_i.adsr_i.sstate[0] ;
 wire \sm_i.adsr_i.sstate[1] ;
 wire \sm_i.adsr_i.sstate[2] ;
 wire \sm_i.adsr_i.vout ;
 wire \sm_i.sadsr_sel[0] ;
 wire \sm_i.sadsr_sel[1] ;
 wire \sm_i.scnt_pwm[0] ;
 wire \sm_i.scnt_pwm[1] ;
 wire \sm_i.scnt_pwm[2] ;
 wire \sm_i.scnt_pwm[3] ;
 wire \sm_i.scnt_pwm[4] ;
 wire \sm_i.scnt_pwm[5] ;
 wire \sm_i.scnt_pwm[6] ;
 wire \sm_i.scnt_pwm[7] ;
 wire \sm_i.scnt_pwm_on[0] ;
 wire \sm_i.scnt_pwm_on[1] ;
 wire \sm_i.scnt_pwm_on[2] ;
 wire \sm_i.scnt_pwm_on[3] ;
 wire \sm_i.scnt_pwm_on[4] ;
 wire \sm_i.scnt_pwm_on[5] ;
 wire \sm_i.scnt_pwm_on[6] ;
 wire \sm_i.scnt_pwm_on[7] ;
 wire \sm_i.scnt_pwm_on_en ;
 wire \sm_i.snote_synch[0][0] ;
 wire \sm_i.snote_synch[0][1] ;
 wire \sm_i.snote_synch[0][2] ;
 wire \sm_i.snote_synch[0][3] ;
 wire \sm_i.snote_synch[0][4] ;
 wire \sm_i.snote_synch[1][0] ;
 wire \sm_i.snote_synch[1][1] ;
 wire \sm_i.snote_synch[1][2] ;
 wire \sm_i.snote_synch[1][3] ;
 wire \sm_i.snote_synch[1][4] ;
 wire \sm_i.snote_synch[2][0] ;
 wire \sm_i.snote_synch[2][1] ;
 wire \sm_i.snote_synch[2][2] ;
 wire \sm_i.snote_synch[2][3] ;
 wire \sm_i.snote_synch[2][4] ;
 wire \sm_i.snotes_sel[0] ;
 wire \sm_i.snotes_sel[1] ;
 wire \sm_i.snotes_sel[2] ;
 wire \sm_i.snotes_sel[3] ;
 wire \sm_i.ssw_reg[0][0] ;
 wire \sm_i.ssw_reg[0][1] ;
 wire \sm_i.ssw_reg[0][2] ;
 wire \sm_i.ssw_reg[0][3] ;
 wire \sm_i.ssw_reg[0][4] ;
 wire \sm_i.ssw_reg[0][5] ;
 wire \sm_i.ssw_reg[0][6] ;
 wire \sm_i.ssw_reg[0][7] ;
 wire \sm_i.ssw_reg[1][0] ;
 wire \sm_i.ssw_reg[1][1] ;
 wire \sm_i.ssw_reg[1][2] ;
 wire \sm_i.ssw_reg[1][3] ;
 wire \sm_i.ssw_reg[1][4] ;
 wire \sm_i.ssw_reg[1][5] ;
 wire \sm_i.ssw_reg[1][6] ;
 wire \sm_i.ssw_reg[1][7] ;
 wire \sm_i.ssw_reg[2][0] ;
 wire \sm_i.ssw_reg[2][1] ;
 wire \sm_i.wav_gen_1.rom_ampl_sin_i.addr[0] ;
 wire \sm_i.wav_gen_1.rom_ampl_sin_i.data_out[0] ;
 wire \sm_i.wav_gen_1.rom_ampl_sin_i.data_out[1] ;
 wire \sm_i.wav_gen_1.rom_ampl_sin_i.data_out[2] ;
 wire \sm_i.wav_gen_1.rom_ampl_sin_i.data_out[3] ;
 wire \sm_i.wav_gen_1.rom_ampl_sin_i.data_out[4] ;
 wire \sm_i.wav_gen_1.rom_ampl_sin_i.en ;
 wire \sm_i.wav_gen_1.rom_freq_saw_i.data_out[0] ;
 wire \sm_i.wav_gen_1.rom_freq_saw_i.data_out[10] ;
 wire \sm_i.wav_gen_1.rom_freq_saw_i.data_out[11] ;
 wire \sm_i.wav_gen_1.rom_freq_saw_i.data_out[12] ;
 wire \sm_i.wav_gen_1.rom_freq_saw_i.data_out[1] ;
 wire \sm_i.wav_gen_1.rom_freq_saw_i.data_out[2] ;
 wire \sm_i.wav_gen_1.rom_freq_saw_i.data_out[3] ;
 wire \sm_i.wav_gen_1.rom_freq_saw_i.data_out[4] ;
 wire \sm_i.wav_gen_1.rom_freq_saw_i.data_out[5] ;
 wire \sm_i.wav_gen_1.rom_freq_saw_i.data_out[6] ;
 wire \sm_i.wav_gen_1.rom_freq_saw_i.data_out[7] ;
 wire \sm_i.wav_gen_1.rom_freq_saw_i.data_out[8] ;
 wire \sm_i.wav_gen_1.rom_freq_saw_i.data_out[9] ;
 wire \sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[0] ;
 wire \sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[10] ;
 wire \sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[1] ;
 wire \sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[2] ;
 wire \sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[3] ;
 wire \sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[4] ;
 wire \sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[5] ;
 wire \sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[6] ;
 wire \sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[7] ;
 wire \sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[8] ;
 wire \sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[9] ;
 wire \sm_i.wav_gen_1.smem_rom_ampl_sin_val_is_neg ;
 wire \sm_i.wav_gen_1.snote_enable ;
 wire \sm_i.wav_gen_1.sstep_cnt[0] ;
 wire \sm_i.wav_gen_1.sstep_cnt[10] ;
 wire \sm_i.wav_gen_1.sstep_cnt[11] ;
 wire \sm_i.wav_gen_1.sstep_cnt[12] ;
 wire \sm_i.wav_gen_1.sstep_cnt[13] ;
 wire \sm_i.wav_gen_1.sstep_cnt[14] ;
 wire \sm_i.wav_gen_1.sstep_cnt[15] ;
 wire \sm_i.wav_gen_1.sstep_cnt[1] ;
 wire \sm_i.wav_gen_1.sstep_cnt[2] ;
 wire \sm_i.wav_gen_1.sstep_cnt[3] ;
 wire \sm_i.wav_gen_1.sstep_cnt[4] ;
 wire \sm_i.wav_gen_1.sstep_cnt[5] ;
 wire \sm_i.wav_gen_1.sstep_cnt[6] ;
 wire \sm_i.wav_gen_1.sstep_cnt[7] ;
 wire \sm_i.wav_gen_1.sstep_cnt[8] ;
 wire \sm_i.wav_gen_1.sstep_cnt[9] ;
 wire \sm_i.wav_gen_1.swave_cnt_tri[1] ;
 wire \sm_i.wav_gen_1.swave_cnt_tri[2] ;
 wire \sm_i.wav_gen_1.swave_cnt_tri[3] ;
 wire \sm_i.wav_gen_1.swave_cnt_tri[4] ;
 wire \sm_i.wav_gen_1.swave_cnt_tri[5] ;
 wire \sm_i.wav_gen_1.swave_cnt_tri_down_up_n ;
 wire \sm_i.wav_gen_1.swave_saw[0] ;
 wire \sm_i.wav_gen_1.swave_saw[1] ;
 wire \sm_i.wav_gen_1.swave_saw[2] ;
 wire \sm_i.wav_gen_1.swave_saw[3] ;
 wire \sm_i.wav_gen_1.swave_saw[4] ;
 wire \sm_i.wav_gen_1.swave_saw[5] ;
 wire \sm_i.wav_gen_1.swave_squ[0] ;
 wire \sm_i.wav_gen_1.swave_squ[1] ;
 wire \sm_i.wav_gen_1.swave_squ[5] ;
 wire \sm_i.wav_gen_1.swave_squ_sel ;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire clknet_0_clk;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;

 sg13g2_inv_1 _1258_ (.Y(_0103_),
    .A(net58));
 sg13g2_inv_1 _1259_ (.Y(_0102_),
    .A(net46));
 sg13g2_inv_1 _1260_ (.Y(_0101_),
    .A(net1));
 sg13g2_inv_1 _1261_ (.Y(_0557_),
    .A(net84));
 sg13g2_inv_1 _1262_ (.Y(_0558_),
    .A(net83));
 sg13g2_inv_1 _1263_ (.Y(_0559_),
    .A(net165));
 sg13g2_inv_1 _1264_ (.Y(_0560_),
    .A(net193));
 sg13g2_inv_1 _1265_ (.Y(_0561_),
    .A(\sm_i.adsr_i.scnt_step[20] ));
 sg13g2_inv_1 _1266_ (.Y(_0562_),
    .A(net140));
 sg13g2_inv_1 _1267_ (.Y(_0563_),
    .A(\sm_i.adsr_i.dout[1] ));
 sg13g2_inv_1 _1268_ (.Y(_0564_),
    .A(net304));
 sg13g2_inv_1 _1269_ (.Y(_0565_),
    .A(net205));
 sg13g2_inv_1 _1270_ (.Y(_0566_),
    .A(net284));
 sg13g2_inv_1 _1271_ (.Y(_0567_),
    .A(net301));
 sg13g2_inv_1 _1272_ (.Y(_0568_),
    .A(net209));
 sg13g2_inv_2 _1273_ (.Y(_0569_),
    .A(net305));
 sg13g2_inv_1 _1274_ (.Y(_0570_),
    .A(net282));
 sg13g2_inv_1 _1275_ (.Y(_0571_),
    .A(net202));
 sg13g2_inv_1 _1276_ (.Y(_0572_),
    .A(net66));
 sg13g2_inv_1 _1277_ (.Y(_0573_),
    .A(_0065_));
 sg13g2_inv_1 _1278_ (.Y(_0574_),
    .A(\sm_i.wav_gen_1.sstep_cnt[1] ));
 sg13g2_inv_1 _1279_ (.Y(_0575_),
    .A(\sm_i.wav_gen_1.sstep_cnt[2] ));
 sg13g2_inv_1 _1280_ (.Y(_0576_),
    .A(net191));
 sg13g2_inv_1 _1281_ (.Y(_0577_),
    .A(\sm_i.wav_gen_1.sstep_cnt[5] ));
 sg13g2_inv_1 _1282_ (.Y(_0578_),
    .A(net210));
 sg13g2_inv_1 _1283_ (.Y(_0579_),
    .A(\sm_i.wav_gen_1.sstep_cnt[9] ));
 sg13g2_inv_1 _1284_ (.Y(_0580_),
    .A(\sm_i.wav_gen_1.sstep_cnt[11] ));
 sg13g2_inv_1 _1285_ (.Y(_0581_),
    .A(\sm_i.wav_gen_1.sstep_cnt[14] ));
 sg13g2_inv_2 _1286_ (.Y(_0582_),
    .A(net299));
 sg13g2_inv_2 _1287_ (.Y(_0583_),
    .A(_0053_));
 sg13g2_inv_1 _1288_ (.Y(_0584_),
    .A(net97));
 sg13g2_inv_1 _1289_ (.Y(_0585_),
    .A(net90));
 sg13g2_inv_1 _1290_ (.Y(_0586_),
    .A(net127));
 sg13g2_inv_1 _1291_ (.Y(_0000_),
    .A(net68));
 sg13g2_inv_1 _1292_ (.Y(_0587_),
    .A(\sm_i.scnt_pwm[3] ));
 sg13g2_inv_1 _1293_ (.Y(_0588_),
    .A(_0069_));
 sg13g2_inv_1 _1294_ (.Y(_0589_),
    .A(_0066_));
 sg13g2_inv_1 _1295_ (.Y(_0590_),
    .A(\sm_i.snote_synch[2][4] ));
 sg13g2_inv_2 _1296_ (.Y(_0591_),
    .A(\sm_i.snotes_sel[1] ));
 sg13g2_inv_2 _1297_ (.Y(_0592_),
    .A(\sm_i.snotes_sel[0] ));
 sg13g2_inv_1 _1298_ (.Y(_0593_),
    .A(net114));
 sg13g2_inv_1 _1299_ (.Y(_0594_),
    .A(net143));
 sg13g2_inv_1 _1300_ (.Y(_0595_),
    .A(net175));
 sg13g2_inv_1 _1301_ (.Y(_0596_),
    .A(net158));
 sg13g2_inv_1 _1302_ (.Y(_0597_),
    .A(net120));
 sg13g2_inv_1 _1303_ (.Y(_0598_),
    .A(net162));
 sg13g2_inv_1 _1304_ (.Y(_0599_),
    .A(net125));
 sg13g2_inv_1 _1305_ (.Y(_0600_),
    .A(net117));
 sg13g2_inv_1 _1306_ (.Y(_0601_),
    .A(_0084_));
 sg13g2_inv_1 _1307_ (.Y(_0602_),
    .A(\sm_i.sadsr_sel[0] ));
 sg13g2_and2_1 _1308_ (.A(net66),
    .B(net67),
    .X(_0030_));
 sg13g2_nor2_1 _1309_ (.A(_0572_),
    .B(net67),
    .Y(_0031_));
 sg13g2_nor2_1 _1310_ (.A(_0569_),
    .B(net239),
    .Y(_0024_));
 sg13g2_nor2_1 _1311_ (.A(_0570_),
    .B(net239),
    .Y(_0025_));
 sg13g2_nor2_1 _1312_ (.A(_0571_),
    .B(net239),
    .Y(_0026_));
 sg13g2_and2_1 _1313_ (.A(net123),
    .B(net66),
    .X(_0027_));
 sg13g2_and2_1 _1314_ (.A(net169),
    .B(net66),
    .X(_0028_));
 sg13g2_and2_1 _1315_ (.A(net245),
    .B(net66),
    .X(_0029_));
 sg13g2_nor2b_2 _1316_ (.A(net240),
    .B_N(\sm_i.ssw_reg[2][1] ),
    .Y(_0603_));
 sg13g2_nand2b_1 _1317_ (.Y(_0604_),
    .B(\sm_i.ssw_reg[2][1] ),
    .A_N(\sm_i.ssw_reg[2][0] ));
 sg13g2_mux2_2 _1318_ (.A0(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[0] ),
    .A1(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[0] ),
    .S(net237),
    .X(_0605_));
 sg13g2_mux2_2 _1319_ (.A0(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[1] ),
    .A1(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[1] ),
    .S(net237),
    .X(_0606_));
 sg13g2_mux2_1 _1320_ (.A0(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[2] ),
    .A1(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[2] ),
    .S(net237),
    .X(_0607_));
 sg13g2_nor3_1 _1321_ (.A(_0605_),
    .B(_0606_),
    .C(_0607_),
    .Y(_0608_));
 sg13g2_mux2_1 _1322_ (.A0(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[3] ),
    .A1(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[3] ),
    .S(net237),
    .X(_0609_));
 sg13g2_nor4_2 _1323_ (.A(_0605_),
    .B(_0606_),
    .C(_0607_),
    .Y(_0610_),
    .D(_0609_));
 sg13g2_nor2_1 _1324_ (.A(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[4] ),
    .B(_0603_),
    .Y(_0611_));
 sg13g2_a21oi_2 _1325_ (.B1(_0611_),
    .Y(_0612_),
    .A2(net238),
    .A1(_0598_));
 sg13g2_nand2b_2 _1326_ (.Y(_0613_),
    .B(_0610_),
    .A_N(_0612_));
 sg13g2_nor2_1 _1327_ (.A(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[5] ),
    .B(net238),
    .Y(_0614_));
 sg13g2_a21oi_2 _1328_ (.B1(_0614_),
    .Y(_0615_),
    .A2(net238),
    .A1(_0596_));
 sg13g2_mux2_1 _1329_ (.A0(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[6] ),
    .A1(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[6] ),
    .S(net236),
    .X(_0616_));
 sg13g2_nor3_2 _1330_ (.A(_0613_),
    .B(_0615_),
    .C(_0616_),
    .Y(_0617_));
 sg13g2_nor2_1 _1331_ (.A(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[7] ),
    .B(net238),
    .Y(_0618_));
 sg13g2_a21oi_1 _1332_ (.A1(_0595_),
    .A2(net238),
    .Y(_0619_),
    .B1(_0618_));
 sg13g2_nor2b_1 _1333_ (.A(_0619_),
    .B_N(_0617_),
    .Y(_0620_));
 sg13g2_mux2_1 _1334_ (.A0(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[8] ),
    .A1(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[8] ),
    .S(net236),
    .X(_0621_));
 sg13g2_inv_1 _1335_ (.Y(_0622_),
    .A(_0621_));
 sg13g2_nand2_1 _1336_ (.Y(_0623_),
    .A(_0620_),
    .B(_0622_));
 sg13g2_mux2_1 _1337_ (.A0(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[9] ),
    .A1(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[9] ),
    .S(net236),
    .X(_0624_));
 sg13g2_nor2_1 _1338_ (.A(_0623_),
    .B(_0624_),
    .Y(_0625_));
 sg13g2_nor2_1 _1339_ (.A(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[10] ),
    .B(net236),
    .Y(_0626_));
 sg13g2_a21oi_2 _1340_ (.B1(_0626_),
    .Y(_0627_),
    .A2(net236),
    .A1(_0600_));
 sg13g2_nand2b_1 _1341_ (.Y(_0628_),
    .B(_0625_),
    .A_N(_0627_));
 sg13g2_nand2_1 _1342_ (.Y(_0629_),
    .A(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[11] ),
    .B(net238));
 sg13g2_nor2b_2 _1343_ (.A(_0628_),
    .B_N(_0629_),
    .Y(_0630_));
 sg13g2_and2_1 _1344_ (.A(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[12] ),
    .B(net236),
    .X(_0631_));
 sg13g2_nor2_1 _1345_ (.A(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[12] ),
    .B(_0630_),
    .Y(_0632_));
 sg13g2_or3_1 _1346_ (.A(\sm_i.wav_gen_1.sstep_cnt[15] ),
    .B(_0631_),
    .C(_0632_),
    .X(_0633_));
 sg13g2_nor2_1 _1347_ (.A(_0059_),
    .B(net236),
    .Y(_0634_));
 sg13g2_xor2_1 _1348_ (.B(_0634_),
    .A(_0630_),
    .X(_0635_));
 sg13g2_a21oi_1 _1349_ (.A1(net236),
    .A2(_0630_),
    .Y(_0636_),
    .B1(_0059_));
 sg13g2_a21o_1 _1350_ (.A2(_0630_),
    .A1(_0059_),
    .B1(_0636_),
    .X(_0637_));
 sg13g2_xor2_1 _1351_ (.B(_0637_),
    .A(_0081_),
    .X(_0638_));
 sg13g2_o21ai_1 _1352_ (.B1(_0638_),
    .Y(_0639_),
    .A1(_0080_),
    .A2(_0635_));
 sg13g2_and2_1 _1353_ (.A(_0080_),
    .B(_0635_),
    .X(_0640_));
 sg13g2_xnor2_1 _1354_ (.Y(_0641_),
    .A(_0628_),
    .B(_0629_));
 sg13g2_nand2_1 _1355_ (.Y(_0642_),
    .A(\sm_i.wav_gen_1.sstep_cnt[11] ),
    .B(_0641_));
 sg13g2_xnor2_1 _1356_ (.Y(_0643_),
    .A(_0623_),
    .B(_0624_));
 sg13g2_xnor2_1 _1357_ (.Y(_0644_),
    .A(_0617_),
    .B(_0619_));
 sg13g2_nand2_1 _1358_ (.Y(_0645_),
    .A(\sm_i.wav_gen_1.sstep_cnt[7] ),
    .B(_0644_));
 sg13g2_xnor2_1 _1359_ (.Y(_0646_),
    .A(_0613_),
    .B(_0615_));
 sg13g2_xnor2_1 _1360_ (.Y(_0647_),
    .A(_0610_),
    .B(_0612_));
 sg13g2_nand2b_1 _1361_ (.Y(_0648_),
    .B(_0074_),
    .A_N(_0647_));
 sg13g2_xnor2_1 _1362_ (.Y(_0649_),
    .A(_0608_),
    .B(_0609_));
 sg13g2_a22oi_1 _1363_ (.Y(_0650_),
    .B1(_0649_),
    .B2(\sm_i.wav_gen_1.sstep_cnt[3] ),
    .A2(_0647_),
    .A1(_0576_));
 sg13g2_inv_1 _1364_ (.Y(_0651_),
    .A(_0650_));
 sg13g2_nor2_1 _1365_ (.A(\sm_i.wav_gen_1.sstep_cnt[3] ),
    .B(_0649_),
    .Y(_0652_));
 sg13g2_o21ai_1 _1366_ (.B1(_0607_),
    .Y(_0653_),
    .A1(_0605_),
    .A2(_0606_));
 sg13g2_nand2b_1 _1367_ (.Y(_0654_),
    .B(_0653_),
    .A_N(_0608_));
 sg13g2_nand2_1 _1368_ (.Y(_0655_),
    .A(\sm_i.wav_gen_1.sstep_cnt[0] ),
    .B(_0605_));
 sg13g2_xnor2_1 _1369_ (.Y(_0656_),
    .A(_0605_),
    .B(_0606_));
 sg13g2_o21ai_1 _1370_ (.B1(_0655_),
    .Y(_0657_),
    .A1(_0574_),
    .A2(_0656_));
 sg13g2_nand2_1 _1371_ (.Y(_0658_),
    .A(_0574_),
    .B(_0656_));
 sg13g2_nand2_1 _1372_ (.Y(_0659_),
    .A(_0657_),
    .B(_0658_));
 sg13g2_xor2_1 _1373_ (.B(_0654_),
    .A(_0073_),
    .X(_0660_));
 sg13g2_a221oi_1 _1374_ (.B2(_0660_),
    .C1(_0652_),
    .B1(_0659_),
    .A1(_0575_),
    .Y(_0661_),
    .A2(_0654_));
 sg13g2_nand3_1 _1375_ (.B(_0650_),
    .C(_0660_),
    .A(_0648_),
    .Y(_0662_));
 sg13g2_o21ai_1 _1376_ (.B1(_0648_),
    .Y(_0663_),
    .A1(_0651_),
    .A2(_0661_));
 sg13g2_xor2_1 _1377_ (.B(_0646_),
    .A(_0075_),
    .X(_0664_));
 sg13g2_a22oi_1 _1378_ (.Y(_0665_),
    .B1(_0663_),
    .B2(_0664_),
    .A2(_0646_),
    .A1(_0577_));
 sg13g2_o21ai_1 _1379_ (.B1(_0616_),
    .Y(_0666_),
    .A1(_0613_),
    .A2(_0615_));
 sg13g2_nor2b_1 _1380_ (.A(_0617_),
    .B_N(_0666_),
    .Y(_0667_));
 sg13g2_xor2_1 _1381_ (.B(_0667_),
    .A(_0076_),
    .X(_0668_));
 sg13g2_or2_1 _1382_ (.X(_0669_),
    .B(_0667_),
    .A(\sm_i.wav_gen_1.sstep_cnt[6] ));
 sg13g2_o21ai_1 _1383_ (.B1(_0669_),
    .Y(_0670_),
    .A1(_0665_),
    .A2(_0668_));
 sg13g2_xnor2_1 _1384_ (.Y(_0671_),
    .A(_0620_),
    .B(_0622_));
 sg13g2_nor2_1 _1385_ (.A(\sm_i.wav_gen_1.sstep_cnt[7] ),
    .B(_0644_),
    .Y(_0672_));
 sg13g2_a21o_1 _1386_ (.A2(_0671_),
    .A1(_0077_),
    .B1(_0672_),
    .X(_0673_));
 sg13g2_a21o_1 _1387_ (.A2(_0670_),
    .A1(_0645_),
    .B1(_0673_),
    .X(_0674_));
 sg13g2_nor2_1 _1388_ (.A(_0077_),
    .B(_0671_),
    .Y(_0675_));
 sg13g2_xnor2_1 _1389_ (.Y(_0676_),
    .A(_0078_),
    .B(_0643_));
 sg13g2_nor2_1 _1390_ (.A(_0675_),
    .B(_0676_),
    .Y(_0677_));
 sg13g2_a22oi_1 _1391_ (.Y(_0678_),
    .B1(_0674_),
    .B2(_0677_),
    .A2(_0643_),
    .A1(_0579_));
 sg13g2_xnor2_1 _1392_ (.Y(_0679_),
    .A(_0625_),
    .B(_0627_));
 sg13g2_xor2_1 _1393_ (.B(_0679_),
    .A(_0079_),
    .X(_0680_));
 sg13g2_nor2_1 _1394_ (.A(_0678_),
    .B(_0680_),
    .Y(_0681_));
 sg13g2_or2_1 _1395_ (.X(_0682_),
    .B(_0641_),
    .A(\sm_i.wav_gen_1.sstep_cnt[11] ));
 sg13g2_o21ai_1 _1396_ (.B1(_0682_),
    .Y(_0683_),
    .A1(\sm_i.wav_gen_1.sstep_cnt[10] ),
    .A2(_0679_));
 sg13g2_o21ai_1 _1397_ (.B1(_0642_),
    .Y(_0684_),
    .A1(_0681_),
    .A2(_0683_));
 sg13g2_nor2b_1 _1398_ (.A(_0640_),
    .B_N(_0684_),
    .Y(_0685_));
 sg13g2_nand2b_1 _1399_ (.Y(_0686_),
    .B(_0637_),
    .A_N(\sm_i.wav_gen_1.sstep_cnt[13] ));
 sg13g2_o21ai_1 _1400_ (.B1(_0686_),
    .Y(_0687_),
    .A1(_0639_),
    .A2(_0685_));
 sg13g2_a21oi_1 _1401_ (.A1(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[12] ),
    .A2(net238),
    .Y(_0688_),
    .B1(_0632_));
 sg13g2_xor2_1 _1402_ (.B(_0688_),
    .A(_0082_),
    .X(_0689_));
 sg13g2_a22oi_1 _1403_ (.Y(_0690_),
    .B1(_0689_),
    .B2(_0687_),
    .A2(_0688_),
    .A1(_0581_));
 sg13g2_o21ai_1 _1404_ (.B1(\sm_i.wav_gen_1.sstep_cnt[15] ),
    .Y(_0691_),
    .A1(_0631_),
    .A2(_0632_));
 sg13g2_a21oi_1 _1405_ (.A1(\sm_i.wav_gen_1.sstep_cnt[11] ),
    .A2(_0641_),
    .Y(_0692_),
    .B1(_0680_));
 sg13g2_or2_1 _1406_ (.X(_0693_),
    .B(_0605_),
    .A(\sm_i.wav_gen_1.sstep_cnt[0] ));
 sg13g2_nor2b_1 _1407_ (.A(_0657_),
    .B_N(_0658_),
    .Y(_0694_));
 sg13g2_nor4_1 _1408_ (.A(_0652_),
    .B(_0662_),
    .C(_0668_),
    .D(_0672_),
    .Y(_0695_));
 sg13g2_and4_1 _1409_ (.A(_0645_),
    .B(_0664_),
    .C(_0693_),
    .D(_0694_),
    .X(_0696_));
 sg13g2_xnor2_1 _1410_ (.Y(_0697_),
    .A(_0578_),
    .B(_0671_));
 sg13g2_nand3_1 _1411_ (.B(_0696_),
    .C(_0697_),
    .A(_0695_),
    .Y(_0698_));
 sg13g2_nor3_1 _1412_ (.A(_0640_),
    .B(_0676_),
    .C(_0698_),
    .Y(_0699_));
 sg13g2_nand4_1 _1413_ (.B(_0689_),
    .C(_0692_),
    .A(_0682_),
    .Y(_0700_),
    .D(_0699_));
 sg13g2_o21ai_1 _1414_ (.B1(_0691_),
    .Y(_0701_),
    .A1(_0639_),
    .A2(_0700_));
 sg13g2_o21ai_1 _1415_ (.B1(_0633_),
    .Y(_0702_),
    .A1(_0690_),
    .A2(_0701_));
 sg13g2_nand2_2 _1416_ (.Y(_0703_),
    .A(net65),
    .B(_0702_));
 sg13g2_nor2_1 _1417_ (.A(net113),
    .B(net211),
    .Y(_0008_));
 sg13g2_nor2_1 _1418_ (.A(net113),
    .B(net148),
    .Y(_0704_));
 sg13g2_and2_1 _1419_ (.A(net113),
    .B(net148),
    .X(_0705_));
 sg13g2_nor3_1 _1420_ (.A(net212),
    .B(_0704_),
    .C(_0705_),
    .Y(_0015_));
 sg13g2_xor2_1 _1421_ (.B(_0705_),
    .A(net178),
    .X(_0706_));
 sg13g2_nor2_1 _1422_ (.A(net211),
    .B(_0706_),
    .Y(_0016_));
 sg13g2_a21oi_1 _1423_ (.A1(\sm_i.wav_gen_1.sstep_cnt[2] ),
    .A2(_0705_),
    .Y(_0707_),
    .B1(net137));
 sg13g2_and3_1 _1424_ (.X(_0708_),
    .A(\sm_i.wav_gen_1.sstep_cnt[2] ),
    .B(net137),
    .C(_0705_));
 sg13g2_nor3_1 _1425_ (.A(net211),
    .B(net138),
    .C(_0708_),
    .Y(_0017_));
 sg13g2_nand2_1 _1426_ (.Y(_0709_),
    .A(_0576_),
    .B(_0708_));
 sg13g2_xnor2_1 _1427_ (.Y(_0710_),
    .A(_0576_),
    .B(_0708_));
 sg13g2_nor2_1 _1428_ (.A(net211),
    .B(net192),
    .Y(_0018_));
 sg13g2_xnor2_1 _1429_ (.Y(_0711_),
    .A(net135),
    .B(_0709_));
 sg13g2_nor2_1 _1430_ (.A(net211),
    .B(net136),
    .Y(_0019_));
 sg13g2_and3_1 _1431_ (.X(_0712_),
    .A(\sm_i.wav_gen_1.sstep_cnt[4] ),
    .B(\sm_i.wav_gen_1.sstep_cnt[5] ),
    .C(_0708_));
 sg13g2_xor2_1 _1432_ (.B(_0712_),
    .A(net170),
    .X(_0713_));
 sg13g2_nor2_1 _1433_ (.A(net211),
    .B(net171),
    .Y(_0020_));
 sg13g2_a21oi_1 _1434_ (.A1(\sm_i.wav_gen_1.sstep_cnt[6] ),
    .A2(_0712_),
    .Y(_0714_),
    .B1(net159));
 sg13g2_and3_2 _1435_ (.X(_0715_),
    .A(\sm_i.wav_gen_1.sstep_cnt[6] ),
    .B(net159),
    .C(_0712_));
 sg13g2_nor3_1 _1436_ (.A(net211),
    .B(net160),
    .C(_0715_),
    .Y(_0021_));
 sg13g2_nor2_1 _1437_ (.A(_0578_),
    .B(_0715_),
    .Y(_0716_));
 sg13g2_and2_1 _1438_ (.A(_0578_),
    .B(_0715_),
    .X(_0717_));
 sg13g2_nor3_1 _1439_ (.A(net211),
    .B(net278),
    .C(_0717_),
    .Y(_0022_));
 sg13g2_xor2_1 _1440_ (.B(_0717_),
    .A(net179),
    .X(_0718_));
 sg13g2_nor2_1 _1441_ (.A(net212),
    .B(net180),
    .Y(_0023_));
 sg13g2_nand3_1 _1442_ (.B(\sm_i.wav_gen_1.sstep_cnt[9] ),
    .C(_0715_),
    .A(\sm_i.wav_gen_1.sstep_cnt[8] ),
    .Y(_0719_));
 sg13g2_xnor2_1 _1443_ (.Y(_0720_),
    .A(net149),
    .B(_0719_));
 sg13g2_nor2_1 _1444_ (.A(net212),
    .B(net150),
    .Y(_0009_));
 sg13g2_nand4_1 _1445_ (.B(\sm_i.wav_gen_1.sstep_cnt[9] ),
    .C(\sm_i.wav_gen_1.sstep_cnt[10] ),
    .A(\sm_i.wav_gen_1.sstep_cnt[8] ),
    .Y(_0721_),
    .D(_0715_));
 sg13g2_nand4_1 _1446_ (.B(\sm_i.wav_gen_1.sstep_cnt[9] ),
    .C(\sm_i.wav_gen_1.sstep_cnt[10] ),
    .A(net294),
    .Y(_0722_),
    .D(_0715_));
 sg13g2_and2_1 _1447_ (.A(_0580_),
    .B(net295),
    .X(_0723_));
 sg13g2_nor2_1 _1448_ (.A(_0580_),
    .B(net295),
    .Y(_0724_));
 sg13g2_nor3_1 _1449_ (.A(net212),
    .B(net296),
    .C(_0724_),
    .Y(_0010_));
 sg13g2_nor2b_1 _1450_ (.A(_0724_),
    .B_N(net206),
    .Y(_0725_));
 sg13g2_nor3_1 _1451_ (.A(_0580_),
    .B(net206),
    .C(_0721_),
    .Y(_0726_));
 sg13g2_nor3_1 _1452_ (.A(net212),
    .B(net207),
    .C(_0726_),
    .Y(_0011_));
 sg13g2_xor2_1 _1453_ (.B(_0726_),
    .A(net146),
    .X(_0727_));
 sg13g2_nor2_1 _1454_ (.A(net212),
    .B(net147),
    .Y(_0012_));
 sg13g2_nand3_1 _1455_ (.B(\sm_i.wav_gen_1.sstep_cnt[12] ),
    .C(_0724_),
    .A(\sm_i.wav_gen_1.sstep_cnt[13] ),
    .Y(_0728_));
 sg13g2_xnor2_1 _1456_ (.Y(_0729_),
    .A(net128),
    .B(_0728_));
 sg13g2_nor2_1 _1457_ (.A(net212),
    .B(net129),
    .Y(_0013_));
 sg13g2_or2_1 _1458_ (.X(_0730_),
    .B(_0728_),
    .A(_0581_));
 sg13g2_xor2_1 _1459_ (.B(_0730_),
    .A(net181),
    .X(_0731_));
 sg13g2_nor2_1 _1460_ (.A(net212),
    .B(net182),
    .Y(_0014_));
 sg13g2_nor2_1 _1461_ (.A(net244),
    .B(_0061_),
    .Y(_0732_));
 sg13g2_nor2_2 _1462_ (.A(\sm_i.wav_gen_1.rom_ampl_sin_i.addr[0] ),
    .B(\sm_i.wav_gen_1.swave_cnt_tri[1] ),
    .Y(_0733_));
 sg13g2_nor2_1 _1463_ (.A(\sm_i.wav_gen_1.swave_cnt_tri[2] ),
    .B(\sm_i.wav_gen_1.swave_cnt_tri[3] ),
    .Y(_0734_));
 sg13g2_nor3_1 _1464_ (.A(\sm_i.wav_gen_1.rom_ampl_sin_i.addr[0] ),
    .B(\sm_i.wav_gen_1.swave_cnt_tri[1] ),
    .C(\sm_i.wav_gen_1.swave_cnt_tri[2] ),
    .Y(_0735_));
 sg13g2_nand2_1 _1465_ (.Y(_0736_),
    .A(_0571_),
    .B(_0733_));
 sg13g2_nand2_2 _1466_ (.Y(_0737_),
    .A(_0733_),
    .B(_0734_));
 sg13g2_nor2_1 _1467_ (.A(\sm_i.wav_gen_1.swave_cnt_tri[4] ),
    .B(_0737_),
    .Y(_0738_));
 sg13g2_xor2_1 _1468_ (.B(_0737_),
    .A(\sm_i.wav_gen_1.swave_cnt_tri[4] ),
    .X(_0739_));
 sg13g2_a21oi_1 _1469_ (.A1(net245),
    .A2(_0739_),
    .Y(_0740_),
    .B1(_0732_));
 sg13g2_a21o_1 _1470_ (.A2(_0739_),
    .A1(net245),
    .B1(_0732_),
    .X(_0741_));
 sg13g2_o21ai_1 _1471_ (.B1(\sm_i.wav_gen_1.swave_cnt_tri[2] ),
    .Y(_0742_),
    .A1(\sm_i.wav_gen_1.rom_ampl_sin_i.addr[0] ),
    .A2(\sm_i.wav_gen_1.swave_cnt_tri[1] ));
 sg13g2_nand3_1 _1472_ (.B(_0736_),
    .C(_0742_),
    .A(net244),
    .Y(_0743_));
 sg13g2_o21ai_1 _1473_ (.B1(_0743_),
    .Y(_0744_),
    .A1(net245),
    .A2(_0063_));
 sg13g2_nand2_1 _1474_ (.Y(_0745_),
    .A(\sm_i.wav_gen_1.swave_cnt_tri[3] ),
    .B(_0736_));
 sg13g2_nand3_1 _1475_ (.B(_0737_),
    .C(_0745_),
    .A(net244),
    .Y(_0746_));
 sg13g2_o21ai_1 _1476_ (.B1(_0746_),
    .Y(_0747_),
    .A1(net244),
    .A2(_0062_));
 sg13g2_and2_2 _1477_ (.A(_0744_),
    .B(_0747_),
    .X(_0748_));
 sg13g2_nand2_1 _1478_ (.Y(_0749_),
    .A(_0744_),
    .B(_0747_));
 sg13g2_nor2_1 _1479_ (.A(net245),
    .B(_0064_),
    .Y(_0750_));
 sg13g2_nor2_1 _1480_ (.A(_0569_),
    .B(_0570_),
    .Y(_0751_));
 sg13g2_nor2_1 _1481_ (.A(_0733_),
    .B(_0751_),
    .Y(_0752_));
 sg13g2_a21oi_2 _1482_ (.B1(_0750_),
    .Y(_0753_),
    .A2(_0752_),
    .A1(net244));
 sg13g2_nand2b_1 _1483_ (.Y(_0754_),
    .B(\sm_i.wav_gen_1.rom_ampl_sin_i.addr[0] ),
    .A_N(_0753_));
 sg13g2_nand2_1 _1484_ (.Y(_0755_),
    .A(_0748_),
    .B(_0754_));
 sg13g2_o21ai_1 _1485_ (.B1(_0748_),
    .Y(_0756_),
    .A1(_0573_),
    .A2(_0754_));
 sg13g2_nor2b_1 _1486_ (.A(_0744_),
    .B_N(_0747_),
    .Y(_0757_));
 sg13g2_and2_1 _1487_ (.A(_0569_),
    .B(_0753_),
    .X(_0758_));
 sg13g2_nand2_1 _1488_ (.Y(_0759_),
    .A(_0569_),
    .B(_0753_));
 sg13g2_and2_1 _1489_ (.A(_0757_),
    .B(_0758_),
    .X(_0760_));
 sg13g2_nand2b_1 _1490_ (.Y(_0761_),
    .B(_0744_),
    .A_N(_0747_));
 sg13g2_inv_1 _1491_ (.Y(_0762_),
    .A(_0761_));
 sg13g2_and2_1 _1492_ (.A(_0753_),
    .B(_0762_),
    .X(_0763_));
 sg13g2_a21oi_1 _1493_ (.A1(\sm_i.wav_gen_1.rom_ampl_sin_i.addr[0] ),
    .A2(_0763_),
    .Y(_0764_),
    .B1(_0760_));
 sg13g2_a21o_1 _1494_ (.A2(_0764_),
    .A1(_0756_),
    .B1(net232),
    .X(_0765_));
 sg13g2_nand3_1 _1495_ (.B(_0748_),
    .C(_0753_),
    .A(\sm_i.wav_gen_1.rom_ampl_sin_i.addr[0] ),
    .Y(_0766_));
 sg13g2_nor2_2 _1496_ (.A(_0065_),
    .B(_0753_),
    .Y(_0767_));
 sg13g2_nand2_1 _1497_ (.Y(_0768_),
    .A(_0762_),
    .B(_0767_));
 sg13g2_nand2_1 _1498_ (.Y(_0769_),
    .A(_0766_),
    .B(_0768_));
 sg13g2_nand3_1 _1499_ (.B(_0748_),
    .C(_0767_),
    .A(net232),
    .Y(_0770_));
 sg13g2_nor2_2 _1500_ (.A(_0744_),
    .B(_0747_),
    .Y(_0771_));
 sg13g2_nand2_1 _1501_ (.Y(_0772_),
    .A(_0767_),
    .B(_0771_));
 sg13g2_nor2_1 _1502_ (.A(\sm_i.wav_gen_1.rom_ampl_sin_i.addr[0] ),
    .B(_0753_),
    .Y(_0773_));
 sg13g2_and2_1 _1503_ (.A(_0749_),
    .B(_0773_),
    .X(_0774_));
 sg13g2_o21ai_1 _1504_ (.B1(_0774_),
    .Y(_0775_),
    .A1(net232),
    .A2(_0771_));
 sg13g2_nand3_1 _1505_ (.B(_0772_),
    .C(_0775_),
    .A(_0770_),
    .Y(_0776_));
 sg13g2_a21oi_1 _1506_ (.A1(_0740_),
    .A2(_0769_),
    .Y(_0777_),
    .B1(_0776_));
 sg13g2_a21oi_1 _1507_ (.A1(_0765_),
    .A2(_0777_),
    .Y(_0032_),
    .B1(net239));
 sg13g2_nand2_1 _1508_ (.Y(_0778_),
    .A(_0757_),
    .B(_0767_));
 sg13g2_nand3_1 _1509_ (.B(_0757_),
    .C(_0759_),
    .A(_0754_),
    .Y(_0779_));
 sg13g2_nand3_1 _1510_ (.B(_0778_),
    .C(_0779_),
    .A(_0756_),
    .Y(_0780_));
 sg13g2_o21ai_1 _1511_ (.B1(_0741_),
    .Y(_0781_),
    .A1(_0763_),
    .A2(_0780_));
 sg13g2_nand3_1 _1512_ (.B(_0748_),
    .C(_0758_),
    .A(net232),
    .Y(_0782_));
 sg13g2_nand3_1 _1513_ (.B(_0758_),
    .C(_0771_),
    .A(_0741_),
    .Y(_0783_));
 sg13g2_nand3_1 _1514_ (.B(_0759_),
    .C(_0771_),
    .A(_0754_),
    .Y(_0784_));
 sg13g2_or2_1 _1515_ (.X(_0785_),
    .B(_0784_),
    .A(_0741_));
 sg13g2_o21ai_1 _1516_ (.B1(_0779_),
    .Y(_0786_),
    .A1(_0759_),
    .A2(_0761_));
 sg13g2_nand2_1 _1517_ (.Y(_0787_),
    .A(net232),
    .B(_0786_));
 sg13g2_o21ai_1 _1518_ (.B1(_0740_),
    .Y(_0788_),
    .A1(_0769_),
    .A2(_0786_));
 sg13g2_and4_1 _1519_ (.A(_0782_),
    .B(_0783_),
    .C(_0785_),
    .D(_0788_),
    .X(_0789_));
 sg13g2_a21oi_1 _1520_ (.A1(_0781_),
    .A2(_0789_),
    .Y(_0033_),
    .B1(net239));
 sg13g2_o21ai_1 _1521_ (.B1(_0762_),
    .Y(_0790_),
    .A1(_0767_),
    .A2(_0773_));
 sg13g2_nand2b_1 _1522_ (.Y(_0791_),
    .B(_0790_),
    .A_N(_0760_));
 sg13g2_nor2_1 _1523_ (.A(_0780_),
    .B(_0791_),
    .Y(_0792_));
 sg13g2_nor2_1 _1524_ (.A(net232),
    .B(_0792_),
    .Y(_0793_));
 sg13g2_a21oi_1 _1525_ (.A1(_0748_),
    .A2(_0773_),
    .Y(_0794_),
    .B1(_0760_));
 sg13g2_a21oi_1 _1526_ (.A1(_0772_),
    .A2(_0794_),
    .Y(_0795_),
    .B1(_0741_));
 sg13g2_nand2_1 _1527_ (.Y(_0796_),
    .A(_0770_),
    .B(_0783_));
 sg13g2_nor3_1 _1528_ (.A(_0793_),
    .B(_0795_),
    .C(_0796_),
    .Y(_0797_));
 sg13g2_a21oi_1 _1529_ (.A1(_0787_),
    .A2(_0797_),
    .Y(_0034_),
    .B1(net239));
 sg13g2_nand3_1 _1530_ (.B(_0779_),
    .C(_0790_),
    .A(_0764_),
    .Y(_0798_));
 sg13g2_nand2_1 _1531_ (.Y(_0799_),
    .A(net232),
    .B(_0798_));
 sg13g2_nand3b_1 _1532_ (.B(_0772_),
    .C(_0784_),
    .Y(_0800_),
    .A_N(_0763_));
 sg13g2_a21oi_1 _1533_ (.A1(_0741_),
    .A2(_0800_),
    .Y(_0801_),
    .B1(_0793_));
 sg13g2_a21oi_1 _1534_ (.A1(_0799_),
    .A2(_0801_),
    .Y(_0035_),
    .B1(net239));
 sg13g2_nand2_1 _1535_ (.Y(_0802_),
    .A(_0755_),
    .B(_0778_));
 sg13g2_a21oi_1 _1536_ (.A1(net232),
    .A2(_0802_),
    .Y(_0803_),
    .B1(_0796_));
 sg13g2_a21oi_1 _1537_ (.A1(_0801_),
    .A2(_0803_),
    .Y(_0036_),
    .B1(net239));
 sg13g2_xor2_1 _1538_ (.B(net99),
    .A(net68),
    .X(_0001_));
 sg13g2_nand3_1 _1539_ (.B(net99),
    .C(net281),
    .A(net68),
    .Y(_0804_));
 sg13g2_a21o_1 _1540_ (.A2(net99),
    .A1(net68),
    .B1(net281),
    .X(_0805_));
 sg13g2_and2_1 _1541_ (.A(_0804_),
    .B(_0805_),
    .X(_0002_));
 sg13g2_nor2_1 _1542_ (.A(_0587_),
    .B(_0804_),
    .Y(_0806_));
 sg13g2_xnor2_1 _1543_ (.Y(_0003_),
    .A(net88),
    .B(_0804_));
 sg13g2_and2_1 _1544_ (.A(net81),
    .B(_0806_),
    .X(_0807_));
 sg13g2_xor2_1 _1545_ (.B(_0806_),
    .A(net81),
    .X(_0004_));
 sg13g2_xor2_1 _1546_ (.B(_0807_),
    .A(net112),
    .X(_0005_));
 sg13g2_and3_2 _1547_ (.X(_0808_),
    .A(net112),
    .B(net72),
    .C(_0807_));
 sg13g2_a21oi_1 _1548_ (.A1(\sm_i.scnt_pwm[5] ),
    .A2(_0807_),
    .Y(_0809_),
    .B1(net72));
 sg13g2_nor2_1 _1549_ (.A(_0808_),
    .B(net73),
    .Y(_0006_));
 sg13g2_and2_2 _1550_ (.A(net124),
    .B(_0808_),
    .X(_0810_));
 sg13g2_nand2_2 _1551_ (.Y(_0811_),
    .A(net124),
    .B(_0808_));
 sg13g2_xor2_1 _1552_ (.B(_0808_),
    .A(net124),
    .X(_0007_));
 sg13g2_nor2_2 _1553_ (.A(\sm_i.adsr_i.sstate[0] ),
    .B(\sm_i.adsr_i.sstate[1] ),
    .Y(_0812_));
 sg13g2_and2_1 _1554_ (.A(\sm_i.adsr_i.sstate[2] ),
    .B(_0812_),
    .X(_0813_));
 sg13g2_nand2_2 _1555_ (.Y(_0814_),
    .A(\sm_i.adsr_i.sstate[2] ),
    .B(_0812_));
 sg13g2_nand2_1 _1556_ (.Y(_0815_),
    .A(\sm_i.adsr_i.sstate[0] ),
    .B(_0084_));
 sg13g2_nand2b_1 _1557_ (.Y(_0816_),
    .B(\sm_i.adsr_i.sstate[1] ),
    .A_N(\sm_i.adsr_i.sstate[0] ));
 sg13g2_or2_2 _1558_ (.X(_0817_),
    .B(_0816_),
    .A(_0601_));
 sg13g2_and2_1 _1559_ (.A(_0814_),
    .B(_0817_),
    .X(_0818_));
 sg13g2_nand2_2 _1560_ (.Y(_0819_),
    .A(_0814_),
    .B(_0817_));
 sg13g2_and2_1 _1561_ (.A(_0815_),
    .B(_0818_),
    .X(_0820_));
 sg13g2_inv_1 _1562_ (.Y(\sm_i.adsr_i.vout ),
    .A(net229));
 sg13g2_or2_2 _1563_ (.X(_0821_),
    .B(\sm_i.scnt_pwm_on[1] ),
    .A(net185));
 sg13g2_nor3_2 _1564_ (.A(net298),
    .B(net155),
    .C(_0821_),
    .Y(_0822_));
 sg13g2_nand2b_2 _1565_ (.Y(_0823_),
    .B(_0822_),
    .A_N(net153));
 sg13g2_nor2_1 _1566_ (.A(net174),
    .B(_0823_),
    .Y(_0824_));
 sg13g2_nor3_2 _1567_ (.A(net174),
    .B(net204),
    .C(_0823_),
    .Y(_0825_));
 sg13g2_nand2b_2 _1568_ (.Y(\sm_i.scnt_pwm_on_en ),
    .B(_0825_),
    .A_N(net85));
 sg13g2_nand3b_1 _1569_ (.B(_0569_),
    .C(\sm_i.wav_gen_1.swave_cnt_tri[1] ),
    .Y(_0826_),
    .A_N(net214));
 sg13g2_nand3b_1 _1570_ (.B(_0734_),
    .C(net244),
    .Y(_0827_),
    .A_N(\sm_i.wav_gen_1.swave_cnt_tri[4] ));
 sg13g2_or2_1 _1571_ (.X(_0828_),
    .B(_0827_),
    .A(net130));
 sg13g2_o21ai_1 _1572_ (.B1(net67),
    .Y(_0829_),
    .A1(_0826_),
    .A2(_0828_));
 sg13g2_nand2_1 _1573_ (.Y(_0830_),
    .A(net123),
    .B(net169));
 sg13g2_nor3_2 _1574_ (.A(_0571_),
    .B(net244),
    .C(_0830_),
    .Y(_0831_));
 sg13g2_nand2b_1 _1575_ (.Y(_0832_),
    .B(_0831_),
    .A_N(_0826_));
 sg13g2_o21ai_1 _1576_ (.B1(net131),
    .Y(_0104_),
    .A1(net247),
    .A2(_0832_));
 sg13g2_a21oi_1 _1577_ (.A1(_0751_),
    .A2(_0831_),
    .Y(_0833_),
    .B1(net247));
 sg13g2_and3_2 _1578_ (.X(_0834_),
    .A(net238),
    .B(_0751_),
    .C(_0831_));
 sg13g2_nor3_1 _1579_ (.A(_0569_),
    .B(net282),
    .C(_0827_),
    .Y(_0835_));
 sg13g2_nor3_1 _1580_ (.A(_0833_),
    .B(_0834_),
    .C(_0835_),
    .Y(_0105_));
 sg13g2_nor4_1 _1581_ (.A(\sm_i.adsr_i.dout[3] ),
    .B(\sm_i.adsr_i.dout[2] ),
    .C(\sm_i.adsr_i.dout[5] ),
    .D(\sm_i.adsr_i.dout[4] ),
    .Y(_0836_));
 sg13g2_nand3_1 _1582_ (.B(_0564_),
    .C(_0836_),
    .A(_0563_),
    .Y(_0837_));
 sg13g2_nand3b_1 _1583_ (.B(\sm_i.snote_synch[2][1] ),
    .C(\sm_i.snote_synch[2][0] ),
    .Y(_0838_),
    .A_N(_0086_));
 sg13g2_nor3_2 _1584_ (.A(_0087_),
    .B(_0590_),
    .C(_0838_),
    .Y(_0839_));
 sg13g2_nor2_1 _1585_ (.A(\sm_i.adsr_i.sstate[1] ),
    .B(_0601_),
    .Y(_0840_));
 sg13g2_nand2_1 _1586_ (.Y(_0841_),
    .A(_0084_),
    .B(_0812_));
 sg13g2_a22oi_1 _1587_ (.Y(_0842_),
    .B1(_0813_),
    .B2(_0837_),
    .A2(_0812_),
    .A1(_0084_));
 sg13g2_nand3_1 _1588_ (.B(\sm_i.adsr_i.sstate[1] ),
    .C(_0084_),
    .A(\sm_i.adsr_i.sstate[0] ),
    .Y(_0843_));
 sg13g2_nor2b_1 _1589_ (.A(_0839_),
    .B_N(_0843_),
    .Y(_0844_));
 sg13g2_nand4_1 _1590_ (.B(\sm_i.adsr_i.dout[2] ),
    .C(\sm_i.adsr_i.dout[5] ),
    .A(\sm_i.adsr_i.dout[3] ),
    .Y(_0845_),
    .D(\sm_i.adsr_i.dout[4] ));
 sg13g2_nor3_1 _1591_ (.A(_0563_),
    .B(_0564_),
    .C(_0845_),
    .Y(_0846_));
 sg13g2_nor3_1 _1592_ (.A(\sm_i.sadsr_sel[0] ),
    .B(_0817_),
    .C(_0846_),
    .Y(_0847_));
 sg13g2_nor2_1 _1593_ (.A(_0602_),
    .B(_0817_),
    .Y(_0848_));
 sg13g2_a21oi_1 _1594_ (.A1(_0837_),
    .A2(_0848_),
    .Y(_0849_),
    .B1(_0847_));
 sg13g2_a22oi_1 _1595_ (.Y(_0850_),
    .B1(_0844_),
    .B2(_0849_),
    .A2(_0842_),
    .A1(_0839_));
 sg13g2_nor2_1 _1596_ (.A(\sm_i.adsr_i.sstate[1] ),
    .B(_0815_),
    .Y(_0851_));
 sg13g2_nand2_1 _1597_ (.Y(_0852_),
    .A(\sm_i.adsr_i.sstate[0] ),
    .B(_0840_));
 sg13g2_nor2_1 _1598_ (.A(_0839_),
    .B(_0852_),
    .Y(_0853_));
 sg13g2_nor2b_2 _1599_ (.A(net242),
    .B_N(\sm_i.adsr_i.scnt_pwl[1] ),
    .Y(_0854_));
 sg13g2_nand2_1 _1600_ (.Y(_0855_),
    .A(\sm_i.adsr_i.scnt_pwl[1] ),
    .B(\sm_i.adsr_i.scnt_pwl[2] ));
 sg13g2_nor2_1 _1601_ (.A(net242),
    .B(_0855_),
    .Y(_0856_));
 sg13g2_nand2_2 _1602_ (.Y(_0857_),
    .A(\sm_i.adsr_i.scnt_pwl[2] ),
    .B(_0854_));
 sg13g2_nor2_1 _1603_ (.A(_0582_),
    .B(net242),
    .Y(_0858_));
 sg13g2_a21oi_1 _1604_ (.A1(\sm_i.adsr_i.scnt_pwl[0] ),
    .A2(_0037_),
    .Y(_0859_),
    .B1(_0858_));
 sg13g2_nand2_2 _1605_ (.Y(_0860_),
    .A(_0582_),
    .B(_0854_));
 sg13g2_nor2b_2 _1606_ (.A(\sm_i.adsr_i.scnt_pwl[1] ),
    .B_N(net242),
    .Y(_0861_));
 sg13g2_nand2_2 _1607_ (.Y(_0862_),
    .A(\sm_i.adsr_i.scnt_pwl[2] ),
    .B(_0861_));
 sg13g2_o21ai_1 _1608_ (.B1(\sm_i.adsr_i.scnt_pwl[2] ),
    .Y(_0863_),
    .A1(_0854_),
    .A2(_0861_));
 sg13g2_nor3_2 _1609_ (.A(\sm_i.adsr_i.scnt_pwl[1] ),
    .B(_0582_),
    .C(net242),
    .Y(_0864_));
 sg13g2_inv_1 _1610_ (.Y(_0865_),
    .A(_0864_));
 sg13g2_nand3_1 _1611_ (.B(net242),
    .C(_0085_),
    .A(\sm_i.adsr_i.scnt_pwl[1] ),
    .Y(_0866_));
 sg13g2_nand2_1 _1612_ (.Y(_0867_),
    .A(_0863_),
    .B(_0866_));
 sg13g2_nor2_2 _1613_ (.A(_0864_),
    .B(_0867_),
    .Y(_0868_));
 sg13g2_nand2_1 _1614_ (.Y(_0869_),
    .A(_0085_),
    .B(_0861_));
 sg13g2_inv_1 _1615_ (.Y(_0870_),
    .A(_0869_));
 sg13g2_nand2_2 _1616_ (.Y(_0871_),
    .A(_0860_),
    .B(_0868_));
 sg13g2_nand2_1 _1617_ (.Y(_0872_),
    .A(_0860_),
    .B(_0869_));
 sg13g2_nor2_2 _1618_ (.A(_0870_),
    .B(_0871_),
    .Y(_0873_));
 sg13g2_xnor2_1 _1619_ (.Y(_0874_),
    .A(_0818_),
    .B(_0873_));
 sg13g2_nand2_1 _1620_ (.Y(_0875_),
    .A(_0859_),
    .B(_0874_));
 sg13g2_o21ai_1 _1621_ (.B1(_0875_),
    .Y(_0876_),
    .A1(_0819_),
    .A2(_0859_));
 sg13g2_xor2_1 _1622_ (.B(_0874_),
    .A(_0038_),
    .X(_0877_));
 sg13g2_nor2_2 _1623_ (.A(_0085_),
    .B(_0862_),
    .Y(_0878_));
 sg13g2_a21oi_1 _1624_ (.A1(\sm_i.sadsr_sel[0] ),
    .A2(_0878_),
    .Y(_0879_),
    .B1(_0864_));
 sg13g2_nor3_1 _1625_ (.A(net242),
    .B(_0813_),
    .C(_0879_),
    .Y(_0880_));
 sg13g2_a21oi_1 _1626_ (.A1(_0813_),
    .A2(_0879_),
    .Y(_0881_),
    .B1(_0880_));
 sg13g2_xor2_1 _1627_ (.B(_0817_),
    .A(_0042_),
    .X(_0882_));
 sg13g2_xnor2_1 _1628_ (.Y(_0883_),
    .A(_0881_),
    .B(_0882_));
 sg13g2_xor2_1 _1629_ (.B(_0878_),
    .A(_0817_),
    .X(_0884_));
 sg13g2_nor2_1 _1630_ (.A(\sm_i.sadsr_sel[0] ),
    .B(_0814_),
    .Y(_0885_));
 sg13g2_xnor2_1 _1631_ (.Y(_0886_),
    .A(_0043_),
    .B(_0885_));
 sg13g2_xnor2_1 _1632_ (.Y(_0887_),
    .A(_0884_),
    .B(_0886_));
 sg13g2_xnor2_1 _1633_ (.Y(_0888_),
    .A(_0039_),
    .B(_0819_));
 sg13g2_xnor2_1 _1634_ (.Y(_0889_),
    .A(_0871_),
    .B(_0888_));
 sg13g2_nand2_1 _1635_ (.Y(_0890_),
    .A(_0868_),
    .B(_0872_));
 sg13g2_xnor2_1 _1636_ (.Y(_0891_),
    .A(_0040_),
    .B(_0819_));
 sg13g2_xnor2_1 _1637_ (.Y(_0892_),
    .A(_0890_),
    .B(_0891_));
 sg13g2_nand4_1 _1638_ (.B(_0887_),
    .C(_0889_),
    .A(_0883_),
    .Y(_0893_),
    .D(_0892_));
 sg13g2_xnor2_1 _1639_ (.Y(_0894_),
    .A(net243),
    .B(_0876_));
 sg13g2_a21oi_2 _1640_ (.B1(_0848_),
    .Y(_0895_),
    .A2(net234),
    .A1(\sm_i.sadsr_sel[1] ));
 sg13g2_a21o_2 _1641_ (.A2(net234),
    .A1(\sm_i.sadsr_sel[1] ),
    .B1(_0848_),
    .X(_0896_));
 sg13g2_nand3_1 _1642_ (.B(_0869_),
    .C(net228),
    .A(_0868_),
    .Y(_0897_));
 sg13g2_nor2b_2 _1643_ (.A(_0897_),
    .B_N(_0860_),
    .Y(_0898_));
 sg13g2_a21oi_2 _1644_ (.B1(_0873_),
    .Y(_0899_),
    .A2(net227),
    .A1(_0870_));
 sg13g2_nand2_1 _1645_ (.Y(_0900_),
    .A(_0858_),
    .B(net227));
 sg13g2_nor2_1 _1646_ (.A(_0865_),
    .B(net228),
    .Y(_0901_));
 sg13g2_nand2b_1 _1647_ (.Y(_0902_),
    .B(net227),
    .A_N(_0862_));
 sg13g2_a21o_1 _1648_ (.A2(_0862_),
    .A1(_0860_),
    .B1(_0895_),
    .X(_0903_));
 sg13g2_nand2_1 _1649_ (.Y(_0904_),
    .A(_0857_),
    .B(_0903_));
 sg13g2_nor2_1 _1650_ (.A(_0901_),
    .B(_0904_),
    .Y(_0905_));
 sg13g2_a21oi_1 _1651_ (.A1(_0899_),
    .A2(_0905_),
    .Y(_0906_),
    .B1(_0898_));
 sg13g2_xnor2_1 _1652_ (.Y(_0907_),
    .A(_0048_),
    .B(_0906_));
 sg13g2_and2_1 _1653_ (.A(_0900_),
    .B(_0903_),
    .X(_0908_));
 sg13g2_nor2_2 _1654_ (.A(_0868_),
    .B(_0872_),
    .Y(_0909_));
 sg13g2_a21oi_1 _1655_ (.A1(_0865_),
    .A2(_0866_),
    .Y(_0910_),
    .B1(net228));
 sg13g2_a21o_1 _1656_ (.A2(_0866_),
    .A1(_0865_),
    .B1(net228),
    .X(_0911_));
 sg13g2_nor2_1 _1657_ (.A(_0864_),
    .B(_0910_),
    .Y(_0912_));
 sg13g2_nand3_1 _1658_ (.B(_0909_),
    .C(_0912_),
    .A(_0863_),
    .Y(_0913_));
 sg13g2_nand2_1 _1659_ (.Y(_0914_),
    .A(_0856_),
    .B(net227));
 sg13g2_o21ai_1 _1660_ (.B1(net228),
    .Y(_0915_),
    .A1(_0856_),
    .A2(_0873_));
 sg13g2_nand2_1 _1661_ (.Y(_0916_),
    .A(_0867_),
    .B(net227));
 sg13g2_xnor2_1 _1662_ (.Y(_0917_),
    .A(_0561_),
    .B(_0916_));
 sg13g2_a21o_1 _1663_ (.A2(_0869_),
    .A1(_0868_),
    .B1(net228),
    .X(_0918_));
 sg13g2_nor2_1 _1664_ (.A(\sm_i.adsr_i.scnt_step[18] ),
    .B(_0918_),
    .Y(_0919_));
 sg13g2_o21ai_1 _1665_ (.B1(_0058_),
    .Y(_0920_),
    .A1(_0860_),
    .A2(net227));
 sg13g2_nor3_1 _1666_ (.A(_0058_),
    .B(_0860_),
    .C(net227),
    .Y(_0921_));
 sg13g2_xor2_1 _1667_ (.B(_0898_),
    .A(\sm_i.adsr_i.scnt_step[0] ),
    .X(_0922_));
 sg13g2_nand4_1 _1668_ (.B(_0863_),
    .C(_0899_),
    .A(_0860_),
    .Y(_0923_),
    .D(_0912_));
 sg13g2_nor2b_1 _1669_ (.A(_0898_),
    .B_N(_0923_),
    .Y(_0924_));
 sg13g2_nand4_1 _1670_ (.B(_0899_),
    .C(_0911_),
    .A(_0862_),
    .Y(_0925_),
    .D(_0914_));
 sg13g2_nor2b_1 _1671_ (.A(_0898_),
    .B_N(_0925_),
    .Y(_0926_));
 sg13g2_xnor2_1 _1672_ (.Y(_0927_),
    .A(_0049_),
    .B(_0926_));
 sg13g2_nor2_1 _1673_ (.A(_0873_),
    .B(_0904_),
    .Y(_0928_));
 sg13g2_a21oi_1 _1674_ (.A1(_0912_),
    .A2(_0928_),
    .Y(_0929_),
    .B1(_0898_));
 sg13g2_xor2_1 _1675_ (.B(_0929_),
    .A(_0050_),
    .X(_0930_));
 sg13g2_o21ai_1 _1676_ (.B1(_0916_),
    .Y(_0931_),
    .A1(_0895_),
    .A2(_0909_));
 sg13g2_nand2_1 _1677_ (.Y(_0932_),
    .A(_0582_),
    .B(_0870_));
 sg13g2_a21oi_1 _1678_ (.A1(_0896_),
    .A2(_0932_),
    .Y(_0933_),
    .B1(_0045_));
 sg13g2_nor2_1 _1679_ (.A(_0867_),
    .B(_0901_),
    .Y(_0934_));
 sg13g2_and2_1 _1680_ (.A(_0909_),
    .B(_0934_),
    .X(_0935_));
 sg13g2_nand2b_1 _1681_ (.Y(_0936_),
    .B(_0935_),
    .A_N(_0056_));
 sg13g2_nand2b_1 _1682_ (.Y(_0937_),
    .B(_0056_),
    .A_N(_0935_));
 sg13g2_nand2_1 _1683_ (.Y(_0938_),
    .A(\sm_i.adsr_i.scnt_step[18] ),
    .B(_0918_));
 sg13g2_xor2_1 _1684_ (.B(_0902_),
    .A(\sm_i.adsr_i.scnt_step[22] ),
    .X(_0939_));
 sg13g2_nand2_1 _1685_ (.Y(_0940_),
    .A(_0878_),
    .B(net228));
 sg13g2_or2_1 _1686_ (.X(_0941_),
    .B(_0940_),
    .A(_0055_));
 sg13g2_nor2_1 _1687_ (.A(_0896_),
    .B(_0932_),
    .Y(_0942_));
 sg13g2_o21ai_1 _1688_ (.B1(_0942_),
    .Y(_0943_),
    .A1(\sm_i.adsr_i.scnt_step[1] ),
    .A2(_0583_));
 sg13g2_nand3_1 _1689_ (.B(_0896_),
    .C(_0932_),
    .A(_0045_),
    .Y(_0944_));
 sg13g2_a21oi_1 _1690_ (.A1(\sm_i.adsr_i.scnt_step[1] ),
    .A2(_0583_),
    .Y(_0945_),
    .B1(_0942_));
 sg13g2_or4_1 _1691_ (.A(\sm_i.adsr_i.scnt_step[25] ),
    .B(\sm_i.adsr_i.scnt_step[24] ),
    .C(\sm_i.adsr_i.scnt_step[27] ),
    .D(\sm_i.adsr_i.scnt_step[26] ),
    .X(_0946_));
 sg13g2_a21oi_1 _1692_ (.A1(_0857_),
    .A2(_0909_),
    .Y(_0947_),
    .B1(net228));
 sg13g2_nor2_1 _1693_ (.A(_0910_),
    .B(_0947_),
    .Y(_0948_));
 sg13g2_nand2_1 _1694_ (.Y(_0949_),
    .A(_0872_),
    .B(net227));
 sg13g2_and2_1 _1695_ (.A(_0911_),
    .B(_0949_),
    .X(_0950_));
 sg13g2_a21oi_1 _1696_ (.A1(_0902_),
    .A2(_0950_),
    .Y(_0951_),
    .B1(\sm_i.adsr_i.scnt_step[16] ));
 sg13g2_nand3_1 _1697_ (.B(_0902_),
    .C(_0950_),
    .A(\sm_i.adsr_i.scnt_step[16] ),
    .Y(_0952_));
 sg13g2_and2_1 _1698_ (.A(_0934_),
    .B(_0949_),
    .X(_0953_));
 sg13g2_xnor2_1 _1699_ (.Y(_0954_),
    .A(_0046_),
    .B(_0948_));
 sg13g2_xor2_1 _1700_ (.B(_0913_),
    .A(_0057_),
    .X(_0955_));
 sg13g2_o21ai_1 _1701_ (.B1(_0943_),
    .Y(_0956_),
    .A1(\sm_i.adsr_i.scnt_step[21] ),
    .A2(_0900_));
 sg13g2_xnor2_1 _1702_ (.Y(_0957_),
    .A(\sm_i.adsr_i.scnt_step[23] ),
    .B(_0914_));
 sg13g2_nor4_1 _1703_ (.A(_0945_),
    .B(_0946_),
    .C(_0956_),
    .D(_0957_),
    .Y(_0958_));
 sg13g2_or2_1 _1704_ (.X(_0959_),
    .B(_0908_),
    .A(\sm_i.adsr_i.scnt_step[19] ));
 sg13g2_nand2_1 _1705_ (.Y(_0960_),
    .A(\sm_i.adsr_i.scnt_step[19] ),
    .B(_0908_));
 sg13g2_nand2_1 _1706_ (.Y(_0961_),
    .A(_0051_),
    .B(_0924_));
 sg13g2_o21ai_1 _1707_ (.B1(_0937_),
    .Y(_0962_),
    .A1(\sm_i.adsr_i.scnt_step[10] ),
    .A2(_0953_));
 sg13g2_a221oi_1 _1708_ (.B2(_0055_),
    .C1(_0962_),
    .B1(_0940_),
    .A1(_0047_),
    .Y(_0963_),
    .A2(_0931_));
 sg13g2_nand4_1 _1709_ (.B(_0958_),
    .C(_0959_),
    .A(_0936_),
    .Y(_0964_),
    .D(_0960_));
 sg13g2_o21ai_1 _1710_ (.B1(_0938_),
    .Y(_0965_),
    .A1(_0052_),
    .A2(_0897_));
 sg13g2_nor3_1 _1711_ (.A(_0919_),
    .B(_0951_),
    .C(_0965_),
    .Y(_0966_));
 sg13g2_a21oi_1 _1712_ (.A1(\sm_i.adsr_i.scnt_step[21] ),
    .A2(_0900_),
    .Y(_0967_),
    .B1(_0933_));
 sg13g2_and4_1 _1713_ (.A(_0917_),
    .B(_0939_),
    .C(_0944_),
    .D(_0967_),
    .X(_0968_));
 sg13g2_nand4_1 _1714_ (.B(_0952_),
    .C(_0966_),
    .A(_0920_),
    .Y(_0969_),
    .D(_0968_));
 sg13g2_a21oi_1 _1715_ (.A1(_0052_),
    .A2(_0897_),
    .Y(_0970_),
    .B1(_0921_));
 sg13g2_nand4_1 _1716_ (.B(_0954_),
    .C(_0955_),
    .A(_0922_),
    .Y(_0971_),
    .D(_0970_));
 sg13g2_nor4_1 _1717_ (.A(_0907_),
    .B(_0964_),
    .C(_0969_),
    .D(_0971_),
    .Y(_0972_));
 sg13g2_o21ai_1 _1718_ (.B1(_0961_),
    .Y(_0973_),
    .A1(_0054_),
    .A2(_0915_));
 sg13g2_a21oi_1 _1719_ (.A1(_0054_),
    .A2(_0915_),
    .Y(_0974_),
    .B1(_0973_));
 sg13g2_o21ai_1 _1720_ (.B1(_0941_),
    .Y(_0975_),
    .A1(_0047_),
    .A2(_0931_));
 sg13g2_a21oi_1 _1721_ (.A1(\sm_i.adsr_i.scnt_step[10] ),
    .A2(_0953_),
    .Y(_0976_),
    .B1(_0975_));
 sg13g2_and2_1 _1722_ (.A(_0963_),
    .B(_0976_),
    .X(_0977_));
 sg13g2_o21ai_1 _1723_ (.B1(_0930_),
    .Y(_0978_),
    .A1(_0051_),
    .A2(_0924_));
 sg13g2_nor2_1 _1724_ (.A(_0927_),
    .B(_0978_),
    .Y(_0979_));
 sg13g2_nand4_1 _1725_ (.B(_0974_),
    .C(_0977_),
    .A(_0972_),
    .Y(_0980_),
    .D(_0979_));
 sg13g2_or4_1 _1726_ (.A(_0877_),
    .B(_0893_),
    .C(_0894_),
    .D(_0980_),
    .X(_0981_));
 sg13g2_o21ai_1 _1727_ (.B1(_0853_),
    .Y(_0982_),
    .A1(_0857_),
    .A2(_0981_));
 sg13g2_nand2b_2 _1728_ (.Y(_0983_),
    .B(_0982_),
    .A_N(_0850_));
 sg13g2_o21ai_1 _1729_ (.B1(_0841_),
    .Y(_0984_),
    .A1(_0818_),
    .A2(_0839_));
 sg13g2_mux2_1 _1730_ (.A0(_0984_),
    .A1(net285),
    .S(_0983_),
    .X(_0106_));
 sg13g2_a21oi_1 _1731_ (.A1(_0817_),
    .A2(_0852_),
    .Y(_0985_),
    .B1(_0839_));
 sg13g2_mux2_1 _1732_ (.A0(_0985_),
    .A1(net289),
    .S(_0983_),
    .X(_0107_));
 sg13g2_nor3_1 _1733_ (.A(_0601_),
    .B(_0812_),
    .C(_0844_),
    .Y(_0986_));
 sg13g2_mux2_1 _1734_ (.A0(_0986_),
    .A1(net197),
    .S(_0983_),
    .X(_0108_));
 sg13g2_nor3_2 _1735_ (.A(_0087_),
    .B(\sm_i.snote_synch[2][4] ),
    .C(_0838_),
    .Y(_0987_));
 sg13g2_nand2_2 _1736_ (.Y(_0988_),
    .A(\sm_i.snotes_sel[3] ),
    .B(\sm_i.snotes_sel[2] ));
 sg13g2_nor2_2 _1737_ (.A(\sm_i.snotes_sel[1] ),
    .B(\sm_i.snotes_sel[0] ),
    .Y(_0989_));
 sg13g2_nor2b_1 _1738_ (.A(_0988_),
    .B_N(_0989_),
    .Y(_0990_));
 sg13g2_nor2_2 _1739_ (.A(\sm_i.snotes_sel[3] ),
    .B(\sm_i.snotes_sel[2] ),
    .Y(_0991_));
 sg13g2_nor2_2 _1740_ (.A(_0591_),
    .B(_0592_),
    .Y(_0992_));
 sg13g2_a21oi_2 _1741_ (.B1(_0990_),
    .Y(_0993_),
    .A2(_0992_),
    .A1(_0991_));
 sg13g2_nor2_2 _1742_ (.A(\sm_i.snotes_sel[1] ),
    .B(_0592_),
    .Y(_0994_));
 sg13g2_nor2b_2 _1743_ (.A(\sm_i.snotes_sel[2] ),
    .B_N(\sm_i.snotes_sel[3] ),
    .Y(_0995_));
 sg13g2_nand2_1 _1744_ (.Y(_0996_),
    .A(_0994_),
    .B(_0995_));
 sg13g2_nand2_1 _1745_ (.Y(_0997_),
    .A(_0993_),
    .B(_0996_));
 sg13g2_nor2_1 _1746_ (.A(_0591_),
    .B(\sm_i.snotes_sel[0] ),
    .Y(_0998_));
 sg13g2_nand2_1 _1747_ (.Y(_0999_),
    .A(\sm_i.snotes_sel[3] ),
    .B(_0998_));
 sg13g2_nor2_1 _1748_ (.A(\sm_i.snotes_sel[2] ),
    .B(_0999_),
    .Y(_1000_));
 sg13g2_a21oi_1 _1749_ (.A1(_0991_),
    .A2(_0994_),
    .Y(_1001_),
    .B1(_1000_));
 sg13g2_nor3_2 _1750_ (.A(_0591_),
    .B(\sm_i.snotes_sel[0] ),
    .C(_0988_),
    .Y(_1002_));
 sg13g2_a21oi_1 _1751_ (.A1(_0992_),
    .A2(_0995_),
    .Y(_1003_),
    .B1(_1002_));
 sg13g2_and2_1 _1752_ (.A(_1001_),
    .B(_1003_),
    .X(_1004_));
 sg13g2_nor2b_1 _1753_ (.A(_0998_),
    .B_N(_0991_),
    .Y(_1005_));
 sg13g2_o21ai_1 _1754_ (.B1(_0988_),
    .Y(_1006_),
    .A1(_0989_),
    .A2(_0991_));
 sg13g2_o21ai_1 _1755_ (.B1(_1004_),
    .Y(_1007_),
    .A1(_1005_),
    .A2(_1006_));
 sg13g2_nor2_1 _1756_ (.A(\sm_i.snotes_sel[1] ),
    .B(_1007_),
    .Y(_1008_));
 sg13g2_o21ai_1 _1757_ (.B1(_0987_),
    .Y(_1009_),
    .A1(_0997_),
    .A2(_1008_));
 sg13g2_nand2b_1 _1758_ (.Y(_1010_),
    .B(\sm_i.snote_synch[2][0] ),
    .A_N(\sm_i.snote_synch[2][1] ));
 sg13g2_nand2_1 _1759_ (.Y(_1011_),
    .A(_0086_),
    .B(_1010_));
 sg13g2_a21oi_1 _1760_ (.A1(_0087_),
    .A2(_1011_),
    .Y(_1012_),
    .B1(\sm_i.snote_synch[2][4] ));
 sg13g2_nor3_2 _1761_ (.A(\sm_i.snote_synch[2][3] ),
    .B(_0838_),
    .C(_1012_),
    .Y(_1013_));
 sg13g2_nand4_1 _1762_ (.B(\sm_i.snote_synch[2][1] ),
    .C(_0086_),
    .A(\sm_i.snote_synch[2][0] ),
    .Y(_1014_),
    .D(\sm_i.snote_synch[2][4] ));
 sg13g2_or3_2 _1763_ (.A(_0087_),
    .B(_0590_),
    .C(_1010_),
    .X(_1015_));
 sg13g2_nor2_1 _1764_ (.A(_0987_),
    .B(_1013_),
    .Y(_1016_));
 sg13g2_nand3_1 _1765_ (.B(_1015_),
    .C(_1016_),
    .A(_1014_),
    .Y(_1017_));
 sg13g2_inv_1 _1766_ (.Y(_1018_),
    .A(_1017_));
 sg13g2_nand2_1 _1767_ (.Y(_1019_),
    .A(\sm_i.snotes_sel[2] ),
    .B(_0992_));
 sg13g2_nand2b_1 _1768_ (.Y(_1020_),
    .B(\sm_i.snotes_sel[2] ),
    .A_N(\sm_i.snotes_sel[3] ));
 sg13g2_nand2_1 _1769_ (.Y(_1021_),
    .A(_1019_),
    .B(_1020_));
 sg13g2_o21ai_1 _1770_ (.B1(_1019_),
    .Y(_1022_),
    .A1(\sm_i.snotes_sel[0] ),
    .A2(_1020_));
 sg13g2_nand2_1 _1771_ (.Y(_1023_),
    .A(_1013_),
    .B(_1022_));
 sg13g2_and2_1 _1772_ (.A(_1017_),
    .B(_1023_),
    .X(_1024_));
 sg13g2_nand3b_1 _1773_ (.B(_0994_),
    .C(_1013_),
    .Y(_1025_),
    .A_N(\sm_i.snotes_sel[3] ));
 sg13g2_nor3_1 _1774_ (.A(_0990_),
    .B(_1000_),
    .C(_1021_),
    .Y(_1026_));
 sg13g2_nor2_1 _1775_ (.A(_1015_),
    .B(_1026_),
    .Y(_1027_));
 sg13g2_a22oi_1 _1776_ (.Y(_1028_),
    .B1(_0995_),
    .B2(_0591_),
    .A2(_0991_),
    .A1(_0592_));
 sg13g2_a21oi_1 _1777_ (.A1(_0991_),
    .A2(_0992_),
    .Y(_1029_),
    .B1(_1002_));
 sg13g2_a21oi_1 _1778_ (.A1(_1028_),
    .A2(_1029_),
    .Y(_1030_),
    .B1(_1014_));
 sg13g2_nor2_1 _1779_ (.A(_1027_),
    .B(_1030_),
    .Y(_1031_));
 sg13g2_nand4_1 _1780_ (.B(_1024_),
    .C(_1025_),
    .A(_1009_),
    .Y(_1032_),
    .D(_1031_));
 sg13g2_nand2b_1 _1781_ (.Y(_1033_),
    .B(_0994_),
    .A_N(_0988_));
 sg13g2_nand2_1 _1782_ (.Y(_1034_),
    .A(_0989_),
    .B(_0995_));
 sg13g2_nand4_1 _1783_ (.B(_1029_),
    .C(_1033_),
    .A(_1018_),
    .Y(_1035_),
    .D(_1034_));
 sg13g2_and2_2 _1784_ (.A(_1032_),
    .B(_1035_),
    .X(_1036_));
 sg13g2_nor2b_1 _1785_ (.A(_1022_),
    .B_N(_1028_),
    .Y(_1037_));
 sg13g2_a21oi_2 _1786_ (.B1(_1014_),
    .Y(_1038_),
    .A2(_1037_),
    .A1(_0993_));
 sg13g2_o21ai_1 _1787_ (.B1(_1023_),
    .Y(_1039_),
    .A1(_1002_),
    .A2(_1015_));
 sg13g2_nor3_2 _1788_ (.A(_1018_),
    .B(_1038_),
    .C(_1039_),
    .Y(_1040_));
 sg13g2_nor2_1 _1789_ (.A(\sm_i.snotes_sel[1] ),
    .B(_0997_),
    .Y(_1041_));
 sg13g2_o21ai_1 _1790_ (.B1(_0987_),
    .Y(_1042_),
    .A1(_1007_),
    .A2(_1041_));
 sg13g2_or3_1 _1791_ (.A(_0591_),
    .B(_0592_),
    .C(_1020_),
    .X(_1043_));
 sg13g2_nand3_1 _1792_ (.B(_1033_),
    .C(_1043_),
    .A(_1001_),
    .Y(_1044_));
 sg13g2_a21o_1 _1793_ (.A2(_1019_),
    .A1(_0993_),
    .B1(_1014_),
    .X(_1045_));
 sg13g2_a21oi_1 _1794_ (.A1(\sm_i.snotes_sel[3] ),
    .A2(_0989_),
    .Y(_1046_),
    .B1(_0992_));
 sg13g2_a21oi_1 _1795_ (.A1(_1020_),
    .A2(_1046_),
    .Y(_1047_),
    .B1(_1015_));
 sg13g2_a21oi_1 _1796_ (.A1(_1013_),
    .A2(_1044_),
    .Y(_1048_),
    .B1(_1047_));
 sg13g2_nand4_1 _1797_ (.B(_1042_),
    .C(_1045_),
    .A(_1017_),
    .Y(_1049_),
    .D(_1048_));
 sg13g2_or2_1 _1798_ (.X(_1050_),
    .B(_1017_),
    .A(_0999_));
 sg13g2_and2_2 _1799_ (.A(_1049_),
    .B(_1050_),
    .X(_1051_));
 sg13g2_nor2_1 _1800_ (.A(_1040_),
    .B(_1051_),
    .Y(_1052_));
 sg13g2_inv_1 _1801_ (.Y(_1053_),
    .A(_1052_));
 sg13g2_and2_1 _1802_ (.A(_1036_),
    .B(_1052_),
    .X(_1054_));
 sg13g2_nor2b_2 _1803_ (.A(_1036_),
    .B_N(_1051_),
    .Y(_1055_));
 sg13g2_nor2b_2 _1804_ (.A(_1004_),
    .B_N(_0987_),
    .Y(_1056_));
 sg13g2_a21oi_1 _1805_ (.A1(\sm_i.snotes_sel[2] ),
    .A2(_1033_),
    .Y(_1057_),
    .B1(_1015_));
 sg13g2_nand2b_1 _1806_ (.Y(_1058_),
    .B(_1013_),
    .A_N(_1003_));
 sg13g2_and2_1 _1807_ (.A(_1023_),
    .B(net224),
    .X(_1059_));
 sg13g2_nand2_1 _1808_ (.Y(_1060_),
    .A(_1050_),
    .B(_1059_));
 sg13g2_nor4_2 _1809_ (.A(_1038_),
    .B(_1056_),
    .C(_1057_),
    .Y(_1061_),
    .D(_1060_));
 sg13g2_nor2b_2 _1810_ (.A(_1040_),
    .B_N(_1061_),
    .Y(_1062_));
 sg13g2_nand2_1 _1811_ (.Y(_1063_),
    .A(_1055_),
    .B(_1062_));
 sg13g2_and2_2 _1812_ (.A(_1036_),
    .B(_1051_),
    .X(_1064_));
 sg13g2_nand2_2 _1813_ (.Y(_1065_),
    .A(_1062_),
    .B(_1064_));
 sg13g2_nor2_1 _1814_ (.A(_1036_),
    .B(_1053_),
    .Y(_1066_));
 sg13g2_a21o_1 _1815_ (.A2(_1062_),
    .A1(_1051_),
    .B1(_1066_),
    .X(_1067_));
 sg13g2_nand2_1 _1816_ (.Y(_1068_),
    .A(_1040_),
    .B(_1061_));
 sg13g2_inv_1 _1817_ (.Y(_1069_),
    .A(_1068_));
 sg13g2_nand2_1 _1818_ (.Y(_1070_),
    .A(_1049_),
    .B(_1069_));
 sg13g2_and3_1 _1819_ (.X(_1071_),
    .A(net226),
    .B(net224),
    .C(_1070_));
 sg13g2_nor2_2 _1820_ (.A(_1040_),
    .B(_1061_),
    .Y(_1072_));
 sg13g2_nand2_1 _1821_ (.Y(_1073_),
    .A(_1055_),
    .B(_1072_));
 sg13g2_or2_1 _1822_ (.X(_1074_),
    .B(_1068_),
    .A(_1049_));
 sg13g2_nor2_1 _1823_ (.A(_1036_),
    .B(_1074_),
    .Y(_1075_));
 sg13g2_a21oi_2 _1824_ (.B1(_1075_),
    .Y(_1076_),
    .A2(_1072_),
    .A1(_1055_));
 sg13g2_and4_1 _1825_ (.A(_1053_),
    .B(_1063_),
    .C(_1065_),
    .D(_1076_),
    .X(_1077_));
 sg13g2_a22oi_1 _1826_ (.Y(_0109_),
    .B1(_1071_),
    .B2(_1077_),
    .A2(net231),
    .A1(_0594_));
 sg13g2_nand3b_1 _1827_ (.B(_1035_),
    .C(_1032_),
    .Y(_1078_),
    .A_N(_1074_));
 sg13g2_inv_1 _1828_ (.Y(_1079_),
    .A(_1078_));
 sg13g2_and2_1 _1829_ (.A(_1055_),
    .B(_1069_),
    .X(_1080_));
 sg13g2_nor3_2 _1830_ (.A(net230),
    .B(_1079_),
    .C(_1080_),
    .Y(_1081_));
 sg13g2_nand3_1 _1831_ (.B(_1076_),
    .C(_1081_),
    .A(net224),
    .Y(_1082_));
 sg13g2_o21ai_1 _1832_ (.B1(_1082_),
    .Y(_1083_),
    .A1(net172),
    .A2(net225));
 sg13g2_inv_1 _1833_ (.Y(_0110_),
    .A(_1083_));
 sg13g2_nor2_1 _1834_ (.A(net230),
    .B(_1056_),
    .Y(_1084_));
 sg13g2_a21oi_1 _1835_ (.A1(_1064_),
    .A2(_1069_),
    .Y(_1085_),
    .B1(_1056_));
 sg13g2_and2_1 _1836_ (.A(net225),
    .B(_1085_),
    .X(_1086_));
 sg13g2_nand3_1 _1837_ (.B(_1076_),
    .C(_1086_),
    .A(_1053_),
    .Y(_1087_));
 sg13g2_o21ai_1 _1838_ (.B1(_1087_),
    .Y(_0111_),
    .A1(_0558_),
    .A2(net225));
 sg13g2_nor2_1 _1839_ (.A(net230),
    .B(_1054_),
    .Y(_1088_));
 sg13g2_and2_1 _1840_ (.A(net224),
    .B(_1063_),
    .X(_1089_));
 sg13g2_nand3_1 _1841_ (.B(_1088_),
    .C(_1089_),
    .A(_1073_),
    .Y(_1090_));
 sg13g2_o21ai_1 _1842_ (.B1(_1090_),
    .Y(_1091_),
    .A1(net168),
    .A2(net225));
 sg13g2_inv_1 _1843_ (.Y(_0112_),
    .A(_1091_));
 sg13g2_nand2_1 _1844_ (.Y(_1092_),
    .A(_1064_),
    .B(_1072_));
 sg13g2_nand2_1 _1845_ (.Y(_1093_),
    .A(_1088_),
    .B(_1092_));
 sg13g2_nand2_1 _1846_ (.Y(_1094_),
    .A(net69),
    .B(net230));
 sg13g2_o21ai_1 _1847_ (.B1(_1094_),
    .Y(_0113_),
    .A1(_1056_),
    .A2(_1093_));
 sg13g2_nor2_1 _1848_ (.A(net230),
    .B(_1062_),
    .Y(_1095_));
 sg13g2_a22oi_1 _1849_ (.Y(_0114_),
    .B1(_1073_),
    .B2(_1095_),
    .A2(net231),
    .A1(_0597_));
 sg13g2_nand4_1 _1850_ (.B(_1065_),
    .C(_1074_),
    .A(_1058_),
    .Y(_1096_),
    .D(_1088_));
 sg13g2_o21ai_1 _1851_ (.B1(_1096_),
    .Y(_1097_),
    .A1(net173),
    .A2(net226));
 sg13g2_inv_1 _1852_ (.Y(_0115_),
    .A(_1097_));
 sg13g2_nand2_1 _1853_ (.Y(_1098_),
    .A(net77),
    .B(net231));
 sg13g2_nand3_1 _1854_ (.B(_1076_),
    .C(_1084_),
    .A(net224),
    .Y(_1099_));
 sg13g2_o21ai_1 _1855_ (.B1(_1098_),
    .Y(_0116_),
    .A1(_1080_),
    .A2(_1099_));
 sg13g2_a21oi_2 _1856_ (.B1(_1054_),
    .Y(_1100_),
    .A2(_1072_),
    .A1(_1051_));
 sg13g2_nand2_1 _1857_ (.Y(_1101_),
    .A(net224),
    .B(_1084_));
 sg13g2_nand3_1 _1858_ (.B(_1089_),
    .C(_1100_),
    .A(_1084_),
    .Y(_1102_));
 sg13g2_o21ai_1 _1859_ (.B1(_1102_),
    .Y(_0117_),
    .A1(_0557_),
    .A2(net225));
 sg13g2_nand2_1 _1860_ (.Y(_1103_),
    .A(net78),
    .B(_0820_));
 sg13g2_o21ai_1 _1861_ (.B1(_1103_),
    .Y(_0118_),
    .A1(_1067_),
    .A2(_1101_));
 sg13g2_nand2_2 _1862_ (.Y(_1104_),
    .A(net224),
    .B(_1085_));
 sg13g2_nand2_1 _1863_ (.Y(_1105_),
    .A(_1081_),
    .B(_1104_));
 sg13g2_a21oi_1 _1864_ (.A1(_1064_),
    .A2(_1069_),
    .Y(_1106_),
    .B1(_1105_));
 sg13g2_a21oi_1 _1865_ (.A1(_0600_),
    .A2(net229),
    .Y(_0119_),
    .B1(_1106_));
 sg13g2_nand2_1 _1866_ (.Y(_1107_),
    .A(net246),
    .B(net306));
 sg13g2_xnor2_1 _1867_ (.Y(_1108_),
    .A(_0065_),
    .B(_0834_));
 sg13g2_o21ai_1 _1868_ (.B1(_1107_),
    .Y(_1109_),
    .A1(net246),
    .A2(_1108_));
 sg13g2_o21ai_1 _1869_ (.B1(net248),
    .Y(_1110_),
    .A1(net213),
    .A2(_1109_));
 sg13g2_a21oi_1 _1870_ (.A1(_0569_),
    .A2(net213),
    .Y(_0120_),
    .B1(_1110_));
 sg13g2_xor2_1 _1871_ (.B(_0752_),
    .A(net247),
    .X(_1111_));
 sg13g2_nand2_1 _1872_ (.Y(_1112_),
    .A(net248),
    .B(_1111_));
 sg13g2_a22oi_1 _1873_ (.Y(_0121_),
    .B1(_0703_),
    .B2(_1112_),
    .A2(net214),
    .A1(_0570_));
 sg13g2_xnor2_1 _1874_ (.Y(_1113_),
    .A(_0064_),
    .B(_0834_));
 sg13g2_xnor2_1 _1875_ (.Y(_1114_),
    .A(_0063_),
    .B(_0834_));
 sg13g2_a21o_1 _1876_ (.A2(_1113_),
    .A1(_1108_),
    .B1(_1114_),
    .X(_1115_));
 sg13g2_nand3_1 _1877_ (.B(_1113_),
    .C(_1114_),
    .A(_1108_),
    .Y(_1116_));
 sg13g2_xor2_1 _1878_ (.B(_0733_),
    .A(net291),
    .X(_1117_));
 sg13g2_a21oi_1 _1879_ (.A1(_1115_),
    .A2(_1116_),
    .Y(_1118_),
    .B1(net246));
 sg13g2_a21oi_1 _1880_ (.A1(net246),
    .A2(_1117_),
    .Y(_1119_),
    .B1(_1118_));
 sg13g2_o21ai_1 _1881_ (.B1(net248),
    .Y(_1120_),
    .A1(net213),
    .A2(_1119_));
 sg13g2_a21oi_1 _1882_ (.A1(_0571_),
    .A2(net213),
    .Y(_0122_),
    .B1(_1120_));
 sg13g2_xnor2_1 _1883_ (.Y(_1121_),
    .A(_0062_),
    .B(_0834_));
 sg13g2_nand2b_1 _1884_ (.Y(_1122_),
    .B(_1121_),
    .A_N(_1116_));
 sg13g2_xnor2_1 _1885_ (.Y(_1123_),
    .A(_1116_),
    .B(_1121_));
 sg13g2_o21ai_1 _1886_ (.B1(net247),
    .Y(_1124_),
    .A1(net176),
    .A2(_0735_));
 sg13g2_a21oi_1 _1887_ (.A1(net176),
    .A2(_0735_),
    .Y(_1125_),
    .B1(_1124_));
 sg13g2_nor2b_1 _1888_ (.A(_1125_),
    .B_N(net248),
    .Y(_1126_));
 sg13g2_o21ai_1 _1889_ (.B1(_1126_),
    .Y(_1127_),
    .A1(net247),
    .A2(_1123_));
 sg13g2_nand3_1 _1890_ (.B(net248),
    .C(net214),
    .A(net123),
    .Y(_1128_));
 sg13g2_o21ai_1 _1891_ (.B1(_1128_),
    .Y(_0123_),
    .A1(net214),
    .A2(net177));
 sg13g2_xnor2_1 _1892_ (.Y(_1129_),
    .A(_0061_),
    .B(_0834_));
 sg13g2_nand2b_1 _1893_ (.Y(_1130_),
    .B(_1129_),
    .A_N(_1122_));
 sg13g2_xnor2_1 _1894_ (.Y(_1131_),
    .A(_1122_),
    .B(_1129_));
 sg13g2_xnor2_1 _1895_ (.Y(_1132_),
    .A(_0061_),
    .B(_0737_));
 sg13g2_nand2_1 _1896_ (.Y(_1133_),
    .A(net246),
    .B(_1132_));
 sg13g2_o21ai_1 _1897_ (.B1(_1133_),
    .Y(_1134_),
    .A1(net246),
    .A2(_1131_));
 sg13g2_nand2_1 _1898_ (.Y(_1135_),
    .A(net169),
    .B(net213));
 sg13g2_o21ai_1 _1899_ (.B1(_1135_),
    .Y(_1136_),
    .A1(net213),
    .A2(_1134_));
 sg13g2_and2_1 _1900_ (.A(net248),
    .B(_1136_),
    .X(_0124_));
 sg13g2_nand3_1 _1901_ (.B(net248),
    .C(net213),
    .A(net244),
    .Y(_1137_));
 sg13g2_xnor2_1 _1902_ (.Y(_1138_),
    .A(_0060_),
    .B(_0834_));
 sg13g2_xnor2_1 _1903_ (.Y(_1139_),
    .A(_1130_),
    .B(_1138_));
 sg13g2_o21ai_1 _1904_ (.B1(net246),
    .Y(_1140_),
    .A1(net302),
    .A2(_0738_));
 sg13g2_a21oi_1 _1905_ (.A1(net302),
    .A2(_0738_),
    .Y(_1141_),
    .B1(_1140_));
 sg13g2_nor2b_1 _1906_ (.A(_1141_),
    .B_N(net248),
    .Y(_1142_));
 sg13g2_o21ai_1 _1907_ (.B1(_1142_),
    .Y(_1143_),
    .A1(net246),
    .A2(_1139_));
 sg13g2_o21ai_1 _1908_ (.B1(_1137_),
    .Y(_0125_),
    .A1(net213),
    .A2(net303));
 sg13g2_and2_1 _1909_ (.A(_1071_),
    .B(_1078_),
    .X(_1144_));
 sg13g2_a22oi_1 _1910_ (.Y(_0126_),
    .B1(_1100_),
    .B2(_1144_),
    .A2(net231),
    .A1(_0593_));
 sg13g2_nor2_1 _1911_ (.A(net230),
    .B(_1066_),
    .Y(_1145_));
 sg13g2_nand4_1 _1912_ (.B(_1065_),
    .C(_1100_),
    .A(_1059_),
    .Y(_1146_),
    .D(_1145_));
 sg13g2_o21ai_1 _1913_ (.B1(_1146_),
    .Y(_1147_),
    .A1(net142),
    .A2(net225));
 sg13g2_inv_1 _1914_ (.Y(_0127_),
    .A(_1147_));
 sg13g2_nand2_1 _1915_ (.Y(_1148_),
    .A(net70),
    .B(net231));
 sg13g2_nand2_1 _1916_ (.Y(_1149_),
    .A(_1065_),
    .B(_1100_));
 sg13g2_o21ai_1 _1917_ (.B1(_1148_),
    .Y(_0128_),
    .A1(_1101_),
    .A2(_1149_));
 sg13g2_a22oi_1 _1918_ (.Y(_1150_),
    .B1(_1077_),
    .B2(_1086_),
    .A2(net231),
    .A1(net76));
 sg13g2_inv_1 _1919_ (.Y(_0129_),
    .A(_1150_));
 sg13g2_and2_1 _1920_ (.A(_1092_),
    .B(_1145_),
    .X(_1151_));
 sg13g2_a22oi_1 _1921_ (.Y(_0130_),
    .B1(_1089_),
    .B2(_1151_),
    .A2(net230),
    .A1(_0598_));
 sg13g2_a21oi_1 _1922_ (.A1(_1051_),
    .A2(_1072_),
    .Y(_1152_),
    .B1(_1075_));
 sg13g2_a22oi_1 _1923_ (.Y(_0131_),
    .B1(_1144_),
    .B2(_1152_),
    .A2(net231),
    .A1(_0596_));
 sg13g2_nand3_1 _1924_ (.B(_1068_),
    .C(_1151_),
    .A(net224),
    .Y(_1153_));
 sg13g2_o21ai_1 _1925_ (.B1(_1153_),
    .Y(_1154_),
    .A1(net167),
    .A2(net226));
 sg13g2_inv_1 _1926_ (.Y(_0132_),
    .A(_1154_));
 sg13g2_and4_1 _1927_ (.A(net225),
    .B(_1053_),
    .C(_1065_),
    .D(_1092_),
    .X(_1155_));
 sg13g2_a22oi_1 _1928_ (.Y(_0133_),
    .B1(_1070_),
    .B2(_1155_),
    .A2(net230),
    .A1(_0595_));
 sg13g2_nand2_1 _1929_ (.Y(_1156_),
    .A(net75),
    .B(net229));
 sg13g2_nand2_1 _1930_ (.Y(_1157_),
    .A(_1145_),
    .B(_1152_));
 sg13g2_o21ai_1 _1931_ (.B1(_1156_),
    .Y(_0134_),
    .A1(_1104_),
    .A2(_1157_));
 sg13g2_nand2_1 _1932_ (.Y(_1158_),
    .A(net71),
    .B(net229));
 sg13g2_o21ai_1 _1933_ (.B1(net225),
    .Y(_1159_),
    .A1(_1040_),
    .A2(_1064_));
 sg13g2_o21ai_1 _1934_ (.B1(_1158_),
    .Y(_0135_),
    .A1(_1104_),
    .A2(_1159_));
 sg13g2_nor3_1 _1935_ (.A(net229),
    .B(_1062_),
    .C(_1104_),
    .Y(_0184_));
 sg13g2_a21o_1 _1936_ (.A2(net229),
    .A1(net96),
    .B1(_0184_),
    .X(_0136_));
 sg13g2_a22oi_1 _1937_ (.Y(_0137_),
    .B1(_1081_),
    .B2(_1104_),
    .A2(net229),
    .A1(_0599_));
 sg13g2_and2_1 _1938_ (.A(net102),
    .B(net229),
    .X(_0138_));
 sg13g2_o21ai_1 _1939_ (.B1(_0841_),
    .Y(_0185_),
    .A1(_0814_),
    .A2(_0839_));
 sg13g2_or2_2 _1940_ (.X(_0186_),
    .B(_0185_),
    .A(_0986_));
 sg13g2_nor2_2 _1941_ (.A(_0819_),
    .B(net234),
    .Y(_0187_));
 sg13g2_nor2b_2 _1942_ (.A(_0186_),
    .B_N(_0187_),
    .Y(_0188_));
 sg13g2_inv_1 _1943_ (.Y(_0189_),
    .A(net223));
 sg13g2_nor2_1 _1944_ (.A(_0186_),
    .B(_0187_),
    .Y(_0190_));
 sg13g2_nand2_1 _1945_ (.Y(_0191_),
    .A(_0980_),
    .B(_0190_));
 sg13g2_nand2_1 _1946_ (.Y(_0192_),
    .A(net196),
    .B(net221));
 sg13g2_o21ai_1 _1947_ (.B1(_0192_),
    .Y(_0139_),
    .A1(net196),
    .A2(net217));
 sg13g2_nand2_1 _1948_ (.Y(_0193_),
    .A(net203),
    .B(net221));
 sg13g2_nand2_1 _1949_ (.Y(_0194_),
    .A(\sm_i.adsr_i.scnt_step[0] ),
    .B(\sm_i.adsr_i.scnt_step[1] ));
 sg13g2_xnor2_1 _1950_ (.Y(_0195_),
    .A(net196),
    .B(net203));
 sg13g2_o21ai_1 _1951_ (.B1(_0193_),
    .Y(_0140_),
    .A1(net217),
    .A2(_0195_));
 sg13g2_nand2_1 _1952_ (.Y(_0196_),
    .A(net79),
    .B(net221));
 sg13g2_nor2_1 _1953_ (.A(_0058_),
    .B(_0194_),
    .Y(_0197_));
 sg13g2_xnor2_1 _1954_ (.Y(_0198_),
    .A(_0058_),
    .B(_0194_));
 sg13g2_o21ai_1 _1955_ (.B1(_0196_),
    .Y(_0141_),
    .A1(net217),
    .A2(_0198_));
 sg13g2_nand2_1 _1956_ (.Y(_0199_),
    .A(net94),
    .B(net221));
 sg13g2_xor2_1 _1957_ (.B(_0197_),
    .A(_0057_),
    .X(_0200_));
 sg13g2_o21ai_1 _1958_ (.B1(_0199_),
    .Y(_0142_),
    .A1(net217),
    .A2(_0200_));
 sg13g2_nand2_1 _1959_ (.Y(_0201_),
    .A(net92),
    .B(net222));
 sg13g2_nand4_1 _1960_ (.B(\sm_i.adsr_i.scnt_step[1] ),
    .C(\sm_i.adsr_i.scnt_step[3] ),
    .A(\sm_i.adsr_i.scnt_step[0] ),
    .Y(_0202_),
    .D(net79));
 sg13g2_nor2_1 _1961_ (.A(_0056_),
    .B(_0202_),
    .Y(_0203_));
 sg13g2_xnor2_1 _1962_ (.Y(_0204_),
    .A(_0056_),
    .B(_0202_));
 sg13g2_o21ai_1 _1963_ (.B1(_0201_),
    .Y(_0143_),
    .A1(net218),
    .A2(_0204_));
 sg13g2_nand2_1 _1964_ (.Y(_0205_),
    .A(net100),
    .B(net222));
 sg13g2_xor2_1 _1965_ (.B(_0203_),
    .A(_0055_),
    .X(_0206_));
 sg13g2_o21ai_1 _1966_ (.B1(_0205_),
    .Y(_0144_),
    .A1(net218),
    .A2(_0206_));
 sg13g2_nand2_1 _1967_ (.Y(_0207_),
    .A(net115),
    .B(net220));
 sg13g2_nand2_1 _1968_ (.Y(_0208_),
    .A(net100),
    .B(net92));
 sg13g2_nor2_1 _1969_ (.A(_0202_),
    .B(_0208_),
    .Y(_0209_));
 sg13g2_nor3_1 _1970_ (.A(_0054_),
    .B(_0202_),
    .C(_0208_),
    .Y(_0210_));
 sg13g2_xor2_1 _1971_ (.B(_0209_),
    .A(_0054_),
    .X(_0211_));
 sg13g2_o21ai_1 _1972_ (.B1(_0207_),
    .Y(_0145_),
    .A1(net216),
    .A2(_0211_));
 sg13g2_nand2_1 _1973_ (.Y(_0212_),
    .A(net118),
    .B(net220));
 sg13g2_xnor2_1 _1974_ (.Y(_0213_),
    .A(_0583_),
    .B(_0210_));
 sg13g2_o21ai_1 _1975_ (.B1(_0212_),
    .Y(_0146_),
    .A1(net216),
    .A2(_0213_));
 sg13g2_nand2_1 _1976_ (.Y(_0214_),
    .A(net90),
    .B(net220));
 sg13g2_nand3_1 _1977_ (.B(net115),
    .C(_0209_),
    .A(net118),
    .Y(_0215_));
 sg13g2_nor2_1 _1978_ (.A(_0052_),
    .B(_0215_),
    .Y(_0216_));
 sg13g2_nand3_1 _1979_ (.B(\sm_i.adsr_i.scnt_step[6] ),
    .C(_0209_),
    .A(\sm_i.adsr_i.scnt_step[7] ),
    .Y(_0217_));
 sg13g2_xnor2_1 _1980_ (.Y(_0218_),
    .A(_0052_),
    .B(_0217_));
 sg13g2_o21ai_1 _1981_ (.B1(_0214_),
    .Y(_0147_),
    .A1(net216),
    .A2(_0218_));
 sg13g2_nand2_1 _1982_ (.Y(_0219_),
    .A(net97),
    .B(net220));
 sg13g2_xor2_1 _1983_ (.B(_0216_),
    .A(_0051_),
    .X(_0220_));
 sg13g2_o21ai_1 _1984_ (.B1(_0219_),
    .Y(_0148_),
    .A1(net216),
    .A2(_0220_));
 sg13g2_nand2_1 _1985_ (.Y(_0221_),
    .A(net127),
    .B(net220));
 sg13g2_or3_1 _1986_ (.A(_0584_),
    .B(_0585_),
    .C(_0217_),
    .X(_0222_));
 sg13g2_nor4_2 _1987_ (.A(_0584_),
    .B(_0585_),
    .C(_0586_),
    .Y(_0223_),
    .D(_0215_));
 sg13g2_nor2_1 _1988_ (.A(_0586_),
    .B(_0222_),
    .Y(_0224_));
 sg13g2_xnor2_1 _1989_ (.Y(_0225_),
    .A(_0586_),
    .B(_0222_));
 sg13g2_o21ai_1 _1990_ (.B1(_0221_),
    .Y(_0149_),
    .A1(net216),
    .A2(_0225_));
 sg13g2_nand2_1 _1991_ (.Y(_0226_),
    .A(net133),
    .B(net220));
 sg13g2_xor2_1 _1992_ (.B(_0223_),
    .A(_0050_),
    .X(_0227_));
 sg13g2_o21ai_1 _1993_ (.B1(_0226_),
    .Y(_0150_),
    .A1(net216),
    .A2(_0227_));
 sg13g2_nand2_1 _1994_ (.Y(_0228_),
    .A(net103),
    .B(net220));
 sg13g2_nand2_1 _1995_ (.Y(_0229_),
    .A(\sm_i.adsr_i.scnt_step[11] ),
    .B(_0224_));
 sg13g2_nor2_1 _1996_ (.A(_0049_),
    .B(_0229_),
    .Y(_0230_));
 sg13g2_xnor2_1 _1997_ (.Y(_0231_),
    .A(_0049_),
    .B(_0229_));
 sg13g2_o21ai_1 _1998_ (.B1(_0228_),
    .Y(_0151_),
    .A1(net216),
    .A2(_0231_));
 sg13g2_nand2_1 _1999_ (.Y(_0232_),
    .A(net108),
    .B(net221));
 sg13g2_xor2_1 _2000_ (.B(_0230_),
    .A(_0048_),
    .X(_0233_));
 sg13g2_o21ai_1 _2001_ (.B1(_0232_),
    .Y(_0152_),
    .A1(net217),
    .A2(_0233_));
 sg13g2_nand2_1 _2002_ (.Y(_0234_),
    .A(net121),
    .B(net222));
 sg13g2_and4_1 _2003_ (.A(net103),
    .B(net108),
    .C(\sm_i.adsr_i.scnt_step[11] ),
    .D(_0223_),
    .X(_0235_));
 sg13g2_nand4_1 _2004_ (.B(net108),
    .C(\sm_i.adsr_i.scnt_step[11] ),
    .A(net103),
    .Y(_0236_),
    .D(_0224_));
 sg13g2_nor2_1 _2005_ (.A(_0047_),
    .B(_0236_),
    .Y(_0237_));
 sg13g2_xor2_1 _2006_ (.B(_0235_),
    .A(_0047_),
    .X(_0238_));
 sg13g2_o21ai_1 _2007_ (.B1(_0234_),
    .Y(_0153_),
    .A1(net218),
    .A2(_0238_));
 sg13g2_nand2_1 _2008_ (.Y(_0239_),
    .A(net110),
    .B(net220));
 sg13g2_xor2_1 _2009_ (.B(_0237_),
    .A(_0046_),
    .X(_0240_));
 sg13g2_o21ai_1 _2010_ (.B1(_0239_),
    .Y(_0154_),
    .A1(net216),
    .A2(_0240_));
 sg13g2_nand2_1 _2011_ (.Y(_0241_),
    .A(net199),
    .B(net222));
 sg13g2_nand2_1 _2012_ (.Y(_0242_),
    .A(net121),
    .B(net110));
 sg13g2_nor2_1 _2013_ (.A(_0236_),
    .B(_0242_),
    .Y(_0243_));
 sg13g2_and4_1 _2014_ (.A(\sm_i.adsr_i.scnt_step[14] ),
    .B(\sm_i.adsr_i.scnt_step[15] ),
    .C(\sm_i.adsr_i.scnt_step[16] ),
    .D(_0235_),
    .X(_0244_));
 sg13g2_xnor2_1 _2015_ (.Y(_0245_),
    .A(net199),
    .B(_0243_));
 sg13g2_o21ai_1 _2016_ (.B1(_0241_),
    .Y(_0155_),
    .A1(net218),
    .A2(_0245_));
 sg13g2_xnor2_1 _2017_ (.Y(_0246_),
    .A(_0045_),
    .B(_0244_));
 sg13g2_nand3_1 _2018_ (.B(_0190_),
    .C(_0246_),
    .A(_0980_),
    .Y(_0247_));
 sg13g2_o21ai_1 _2019_ (.B1(_0247_),
    .Y(_0156_),
    .A1(_0559_),
    .A2(_0189_));
 sg13g2_nand2_1 _2020_ (.Y(_0248_),
    .A(net201),
    .B(net223));
 sg13g2_and2_1 _2021_ (.A(net165),
    .B(_0244_),
    .X(_0249_));
 sg13g2_and2_1 _2022_ (.A(net309),
    .B(_0249_),
    .X(_0250_));
 sg13g2_xnor2_1 _2023_ (.Y(_0251_),
    .A(net201),
    .B(_0249_));
 sg13g2_o21ai_1 _2024_ (.B1(_0248_),
    .Y(_0157_),
    .A1(net219),
    .A2(_0251_));
 sg13g2_nand2_1 _2025_ (.Y(_0252_),
    .A(net193),
    .B(net222));
 sg13g2_nand4_1 _2026_ (.B(net165),
    .C(\sm_i.adsr_i.scnt_step[18] ),
    .A(\sm_i.adsr_i.scnt_step[16] ),
    .Y(_0253_),
    .D(_0243_));
 sg13g2_and2_1 _2027_ (.A(\sm_i.adsr_i.scnt_step[19] ),
    .B(_0250_),
    .X(_0254_));
 sg13g2_xnor2_1 _2028_ (.Y(_0255_),
    .A(net193),
    .B(_0250_));
 sg13g2_o21ai_1 _2029_ (.B1(_0252_),
    .Y(_0158_),
    .A1(net218),
    .A2(_0255_));
 sg13g2_nand2_1 _2030_ (.Y(_0256_),
    .A(net144),
    .B(net222));
 sg13g2_xnor2_1 _2031_ (.Y(_0257_),
    .A(net144),
    .B(_0254_));
 sg13g2_o21ai_1 _2032_ (.B1(_0256_),
    .Y(_0159_),
    .A1(net218),
    .A2(_0257_));
 sg13g2_nor3_2 _2033_ (.A(_0560_),
    .B(_0561_),
    .C(_0253_),
    .Y(_0258_));
 sg13g2_nand2_1 _2034_ (.Y(_0259_),
    .A(net194),
    .B(net222));
 sg13g2_and3_1 _2035_ (.X(_0260_),
    .A(net144),
    .B(net310),
    .C(_0254_));
 sg13g2_xnor2_1 _2036_ (.Y(_0261_),
    .A(net194),
    .B(_0258_));
 sg13g2_o21ai_1 _2037_ (.B1(_0259_),
    .Y(_0160_),
    .A1(net218),
    .A2(_0261_));
 sg13g2_nand2_1 _2038_ (.Y(_0262_),
    .A(net190),
    .B(net222));
 sg13g2_and2_1 _2039_ (.A(\sm_i.adsr_i.scnt_step[22] ),
    .B(_0260_),
    .X(_0263_));
 sg13g2_xnor2_1 _2040_ (.Y(_0264_),
    .A(net190),
    .B(_0260_));
 sg13g2_o21ai_1 _2041_ (.B1(_0262_),
    .Y(_0161_),
    .A1(net218),
    .A2(_0264_));
 sg13g2_nand2_1 _2042_ (.Y(_0265_),
    .A(net183),
    .B(net223));
 sg13g2_and2_1 _2043_ (.A(\sm_i.adsr_i.scnt_step[23] ),
    .B(_0263_),
    .X(_0266_));
 sg13g2_xnor2_1 _2044_ (.Y(_0267_),
    .A(net183),
    .B(_0263_));
 sg13g2_nand4_1 _2045_ (.B(net307),
    .C(net183),
    .A(\sm_i.adsr_i.scnt_step[21] ),
    .Y(_0268_),
    .D(_0258_));
 sg13g2_o21ai_1 _2046_ (.B1(_0265_),
    .Y(_0162_),
    .A1(net219),
    .A2(_0267_));
 sg13g2_a21oi_1 _2047_ (.A1(_0189_),
    .A2(_0266_),
    .Y(_0269_),
    .B1(net140));
 sg13g2_nor3_2 _2048_ (.A(_0562_),
    .B(net223),
    .C(net308),
    .Y(_0270_));
 sg13g2_nor3_1 _2049_ (.A(_0186_),
    .B(net141),
    .C(_0270_),
    .Y(_0163_));
 sg13g2_xnor2_1 _2050_ (.Y(_0271_),
    .A(net188),
    .B(_0270_));
 sg13g2_nor2_1 _2051_ (.A(_0186_),
    .B(net189),
    .Y(_0164_));
 sg13g2_a21oi_1 _2052_ (.A1(\sm_i.adsr_i.scnt_step[25] ),
    .A2(_0270_),
    .Y(_0272_),
    .B1(net105));
 sg13g2_nand4_1 _2053_ (.B(net140),
    .C(net105),
    .A(\sm_i.adsr_i.scnt_step[25] ),
    .Y(_0273_),
    .D(_0266_));
 sg13g2_nor2_1 _2054_ (.A(_0187_),
    .B(_0273_),
    .Y(_0274_));
 sg13g2_nor3_1 _2055_ (.A(_0186_),
    .B(net106),
    .C(_0274_),
    .Y(_0165_));
 sg13g2_xnor2_1 _2056_ (.Y(_0275_),
    .A(net151),
    .B(_0274_));
 sg13g2_nor2_1 _2057_ (.A(_0186_),
    .B(net152),
    .Y(_0166_));
 sg13g2_nand2_2 _2058_ (.Y(_0276_),
    .A(_0811_),
    .B(\sm_i.scnt_pwm_on_en ));
 sg13g2_inv_1 _2059_ (.Y(_0277_),
    .A(_0276_));
 sg13g2_nand2_1 _2060_ (.Y(_0278_),
    .A(net63),
    .B(_0277_));
 sg13g2_o21ai_1 _2061_ (.B1(\sm_i.wav_gen_1.rom_ampl_sin_i.data_out[2] ),
    .Y(_0279_),
    .A1(\sm_i.wav_gen_1.rom_ampl_sin_i.data_out[0] ),
    .A2(\sm_i.wav_gen_1.rom_ampl_sin_i.data_out[1] ));
 sg13g2_or3_1 _2062_ (.A(\sm_i.wav_gen_1.rom_ampl_sin_i.data_out[2] ),
    .B(\sm_i.wav_gen_1.rom_ampl_sin_i.data_out[0] ),
    .C(\sm_i.wav_gen_1.rom_ampl_sin_i.data_out[1] ),
    .X(_0280_));
 sg13g2_nand3_1 _2063_ (.B(_0279_),
    .C(_0280_),
    .A(\sm_i.wav_gen_1.smem_rom_ampl_sin_val_is_neg ),
    .Y(_0281_));
 sg13g2_nor2_1 _2064_ (.A(\sm_i.wav_gen_1.smem_rom_ampl_sin_val_is_neg ),
    .B(_0067_),
    .Y(_0282_));
 sg13g2_and2_1 _2065_ (.A(net240),
    .B(\sm_i.ssw_reg[2][1] ),
    .X(_0283_));
 sg13g2_nand2_1 _2066_ (.Y(_0284_),
    .A(net240),
    .B(\sm_i.ssw_reg[2][1] ));
 sg13g2_nor2_1 _2067_ (.A(_0282_),
    .B(_0284_),
    .Y(_0285_));
 sg13g2_nor2b_1 _2068_ (.A(\sm_i.ssw_reg[2][1] ),
    .B_N(net240),
    .Y(_0286_));
 sg13g2_nand3b_1 _2069_ (.B(_0071_),
    .C(net241),
    .Y(_0287_),
    .A_N(\sm_i.ssw_reg[2][1] ));
 sg13g2_o21ai_1 _2070_ (.B1(_0287_),
    .Y(_0288_),
    .A1(net240),
    .A2(\sm_i.wav_gen_1.swave_saw[2] ));
 sg13g2_a21o_2 _2071_ (.A2(_0285_),
    .A1(_0281_),
    .B1(_0288_),
    .X(_0289_));
 sg13g2_nor2_1 _2072_ (.A(_0042_),
    .B(_0289_),
    .Y(_0290_));
 sg13g2_nand2_1 _2073_ (.Y(_0291_),
    .A(\sm_i.wav_gen_1.smem_rom_ampl_sin_val_is_neg ),
    .B(\sm_i.wav_gen_1.rom_ampl_sin_i.data_out[0] ));
 sg13g2_xor2_1 _2074_ (.B(_0291_),
    .A(\sm_i.wav_gen_1.rom_ampl_sin_i.data_out[1] ),
    .X(_0292_));
 sg13g2_o21ai_1 _2075_ (.B1(_0287_),
    .Y(_0293_),
    .A1(net240),
    .A2(\sm_i.wav_gen_1.swave_saw[1] ));
 sg13g2_a21oi_2 _2076_ (.B1(_0293_),
    .Y(_0294_),
    .A2(_0292_),
    .A1(_0283_));
 sg13g2_nand2_1 _2077_ (.Y(_0295_),
    .A(\sm_i.adsr_i.dout[2] ),
    .B(_0294_));
 sg13g2_nor3_1 _2078_ (.A(_0042_),
    .B(_0289_),
    .C(_0295_),
    .Y(_0296_));
 sg13g2_or2_1 _2079_ (.X(_0297_),
    .B(\sm_i.wav_gen_1.swave_saw[0] ),
    .A(net240));
 sg13g2_o21ai_1 _2080_ (.B1(_0297_),
    .Y(_0298_),
    .A1(\sm_i.wav_gen_1.rom_ampl_sin_i.data_out[0] ),
    .A2(_0284_));
 sg13g2_a21oi_2 _2081_ (.B1(_0298_),
    .Y(_0299_),
    .A2(_0286_),
    .A1(_0070_));
 sg13g2_nand2b_1 _2082_ (.Y(_0300_),
    .B(_0299_),
    .A_N(_0040_));
 sg13g2_xor2_1 _2083_ (.B(_0295_),
    .A(_0290_),
    .X(_0301_));
 sg13g2_nor2_1 _2084_ (.A(_0300_),
    .B(_0301_),
    .Y(_0302_));
 sg13g2_nor2_1 _2085_ (.A(_0296_),
    .B(_0302_),
    .Y(_0303_));
 sg13g2_xor2_1 _2086_ (.B(_0301_),
    .A(_0300_),
    .X(_0304_));
 sg13g2_nand2_1 _2087_ (.Y(_0305_),
    .A(\sm_i.wav_gen_1.rom_ampl_sin_i.data_out[3] ),
    .B(_0280_));
 sg13g2_or4_2 _2088_ (.A(\sm_i.wav_gen_1.rom_ampl_sin_i.data_out[3] ),
    .B(\sm_i.wav_gen_1.rom_ampl_sin_i.data_out[2] ),
    .C(\sm_i.wav_gen_1.rom_ampl_sin_i.data_out[0] ),
    .D(\sm_i.wav_gen_1.rom_ampl_sin_i.data_out[1] ),
    .X(_0306_));
 sg13g2_and2_1 _2089_ (.A(\sm_i.wav_gen_1.smem_rom_ampl_sin_val_is_neg ),
    .B(_0306_),
    .X(_0307_));
 sg13g2_o21ai_1 _2090_ (.B1(_0283_),
    .Y(_0308_),
    .A1(\sm_i.wav_gen_1.smem_rom_ampl_sin_val_is_neg ),
    .A2(_0068_));
 sg13g2_a21oi_2 _2091_ (.B1(_0308_),
    .Y(_0309_),
    .A2(_0307_),
    .A1(_0305_));
 sg13g2_o21ai_1 _2092_ (.B1(_0287_),
    .Y(_0310_),
    .A1(net241),
    .A2(\sm_i.wav_gen_1.swave_saw[3] ));
 sg13g2_nor2_1 _2093_ (.A(_0309_),
    .B(_0310_),
    .Y(_0311_));
 sg13g2_or2_2 _2094_ (.X(_0312_),
    .B(_0310_),
    .A(_0309_));
 sg13g2_nor2_1 _2095_ (.A(_0043_),
    .B(_0312_),
    .Y(_0313_));
 sg13g2_nand2_1 _2096_ (.Y(_0314_),
    .A(_0304_),
    .B(_0313_));
 sg13g2_a21oi_1 _2097_ (.A1(\sm_i.wav_gen_1.smem_rom_ampl_sin_val_is_neg ),
    .A2(_0306_),
    .Y(_0315_),
    .B1(_0069_));
 sg13g2_and3_1 _2098_ (.X(_0316_),
    .A(\sm_i.wav_gen_1.smem_rom_ampl_sin_val_is_neg ),
    .B(_0069_),
    .C(_0306_));
 sg13g2_nor3_2 _2099_ (.A(_0284_),
    .B(_0315_),
    .C(_0316_),
    .Y(_0317_));
 sg13g2_o21ai_1 _2100_ (.B1(_0287_),
    .Y(_0318_),
    .A1(net241),
    .A2(\sm_i.wav_gen_1.swave_saw[4] ));
 sg13g2_or2_2 _2101_ (.X(_0319_),
    .B(_0318_),
    .A(_0317_));
 sg13g2_nor2_1 _2102_ (.A(_0043_),
    .B(_0319_),
    .Y(_0320_));
 sg13g2_nor2_1 _2103_ (.A(_0042_),
    .B(_0312_),
    .Y(_0321_));
 sg13g2_or4_1 _2104_ (.A(_0043_),
    .B(_0042_),
    .C(_0312_),
    .D(_0319_),
    .X(_0322_));
 sg13g2_xnor2_1 _2105_ (.Y(_0323_),
    .A(_0320_),
    .B(_0321_));
 sg13g2_nand2_1 _2106_ (.Y(_0324_),
    .A(\sm_i.adsr_i.dout[4] ),
    .B(_0299_));
 sg13g2_inv_1 _2107_ (.Y(_0325_),
    .A(_0324_));
 sg13g2_nor2_1 _2108_ (.A(_0041_),
    .B(_0289_),
    .Y(_0326_));
 sg13g2_nand2_1 _2109_ (.Y(_0327_),
    .A(\sm_i.adsr_i.dout[3] ),
    .B(_0294_));
 sg13g2_nor3_1 _2110_ (.A(_0041_),
    .B(_0289_),
    .C(_0327_),
    .Y(_0328_));
 sg13g2_xnor2_1 _2111_ (.Y(_0329_),
    .A(_0326_),
    .B(_0327_));
 sg13g2_xnor2_1 _2112_ (.Y(_0330_),
    .A(_0324_),
    .B(_0329_));
 sg13g2_nand2b_1 _2113_ (.Y(_0331_),
    .B(_0330_),
    .A_N(_0323_));
 sg13g2_xnor2_1 _2114_ (.Y(_0332_),
    .A(_0323_),
    .B(_0330_));
 sg13g2_nand2b_1 _2115_ (.Y(_0333_),
    .B(_0332_),
    .A_N(_0314_));
 sg13g2_xor2_1 _2116_ (.B(_0332_),
    .A(_0314_),
    .X(_0334_));
 sg13g2_xor2_1 _2117_ (.B(_0334_),
    .A(_0303_),
    .X(_0335_));
 sg13g2_xnor2_1 _2118_ (.Y(_0336_),
    .A(_0304_),
    .B(_0313_));
 sg13g2_nor2b_1 _2119_ (.A(_0042_),
    .B_N(_0294_),
    .Y(_0337_));
 sg13g2_and2_1 _2120_ (.A(_0299_),
    .B(_0337_),
    .X(_0338_));
 sg13g2_a21oi_1 _2121_ (.A1(\sm_i.adsr_i.dout[2] ),
    .A2(_0299_),
    .Y(_0339_),
    .B1(_0337_));
 sg13g2_nor3_1 _2122_ (.A(_0043_),
    .B(_0289_),
    .C(_0339_),
    .Y(_0340_));
 sg13g2_a21oi_1 _2123_ (.A1(\sm_i.adsr_i.dout[2] ),
    .A2(_0338_),
    .Y(_0341_),
    .B1(_0340_));
 sg13g2_nor2_1 _2124_ (.A(_0336_),
    .B(_0341_),
    .Y(_0342_));
 sg13g2_nor2b_1 _2125_ (.A(_0043_),
    .B_N(_0301_),
    .Y(_0343_));
 sg13g2_xor2_1 _2126_ (.B(_0341_),
    .A(_0336_),
    .X(_0344_));
 sg13g2_nand3_1 _2127_ (.B(_0343_),
    .C(_0344_),
    .A(_0338_),
    .Y(_0345_));
 sg13g2_nor2b_1 _2128_ (.A(_0342_),
    .B_N(_0345_),
    .Y(_0346_));
 sg13g2_xnor2_1 _2129_ (.Y(_0347_),
    .A(_0335_),
    .B(_0346_));
 sg13g2_o21ai_1 _2130_ (.B1(_0278_),
    .Y(_0167_),
    .A1(_0811_),
    .A2(_0347_));
 sg13g2_nand4_1 _2131_ (.B(_0338_),
    .C(_0343_),
    .A(_0335_),
    .Y(_0348_),
    .D(_0344_));
 sg13g2_inv_1 _2132_ (.Y(_0349_),
    .A(_0348_));
 sg13g2_nand2_1 _2133_ (.Y(_0350_),
    .A(_0335_),
    .B(_0342_));
 sg13g2_nand2_1 _2134_ (.Y(_0351_),
    .A(\sm_i.adsr_i.dout[5] ),
    .B(_0299_));
 sg13g2_o21ai_1 _2135_ (.B1(_0333_),
    .Y(_0352_),
    .A1(_0303_),
    .A2(_0334_));
 sg13g2_a21oi_1 _2136_ (.A1(_0325_),
    .A2(_0329_),
    .Y(_0353_),
    .B1(_0328_));
 sg13g2_nand2_1 _2137_ (.Y(_0354_),
    .A(\sm_i.adsr_i.dout[4] ),
    .B(_0294_));
 sg13g2_nor3_1 _2138_ (.A(net243),
    .B(_0309_),
    .C(_0310_),
    .Y(_0355_));
 sg13g2_or2_1 _2139_ (.X(_0356_),
    .B(_0289_),
    .A(_0565_));
 sg13g2_or3_1 _2140_ (.A(net243),
    .B(_0312_),
    .C(_0356_),
    .X(_0357_));
 sg13g2_xor2_1 _2141_ (.B(_0356_),
    .A(_0355_),
    .X(_0358_));
 sg13g2_xor2_1 _2142_ (.B(_0358_),
    .A(_0354_),
    .X(_0359_));
 sg13g2_or3_1 _2143_ (.A(_0563_),
    .B(_0317_),
    .C(_0318_),
    .X(_0360_));
 sg13g2_o21ai_1 _2144_ (.B1(_0589_),
    .Y(_0361_),
    .A1(_0588_),
    .A2(_0306_));
 sg13g2_nor2_1 _2145_ (.A(net240),
    .B(\sm_i.wav_gen_1.swave_saw[5] ),
    .Y(_0362_));
 sg13g2_a221oi_1 _2146_ (.B2(_0283_),
    .C1(_0362_),
    .B1(_0361_),
    .A1(_0072_),
    .Y(_0363_),
    .A2(_0286_));
 sg13g2_inv_1 _2147_ (.Y(_0364_),
    .A(net233));
 sg13g2_nand2_1 _2148_ (.Y(_0365_),
    .A(\sm_i.adsr_i.dout[0] ),
    .B(net233));
 sg13g2_xor2_1 _2149_ (.B(_0365_),
    .A(_0360_),
    .X(_0366_));
 sg13g2_nand2b_1 _2150_ (.Y(_0367_),
    .B(_0366_),
    .A_N(_0322_));
 sg13g2_xnor2_1 _2151_ (.Y(_0368_),
    .A(_0322_),
    .B(_0366_));
 sg13g2_nand2_1 _2152_ (.Y(_0369_),
    .A(_0359_),
    .B(_0368_));
 sg13g2_xnor2_1 _2153_ (.Y(_0370_),
    .A(_0359_),
    .B(_0368_));
 sg13g2_nor2_1 _2154_ (.A(_0331_),
    .B(_0370_),
    .Y(_0371_));
 sg13g2_xor2_1 _2155_ (.B(_0370_),
    .A(_0331_),
    .X(_0372_));
 sg13g2_nor2b_1 _2156_ (.A(_0353_),
    .B_N(_0372_),
    .Y(_0373_));
 sg13g2_xnor2_1 _2157_ (.Y(_0374_),
    .A(_0353_),
    .B(_0372_));
 sg13g2_nand2_1 _2158_ (.Y(_0375_),
    .A(_0352_),
    .B(_0374_));
 sg13g2_nor2_1 _2159_ (.A(_0352_),
    .B(_0374_),
    .Y(_0376_));
 sg13g2_xor2_1 _2160_ (.B(_0374_),
    .A(_0352_),
    .X(_0377_));
 sg13g2_xnor2_1 _2161_ (.Y(_0378_),
    .A(_0351_),
    .B(_0377_));
 sg13g2_nor2b_1 _2162_ (.A(_0350_),
    .B_N(_0378_),
    .Y(_0379_));
 sg13g2_xnor2_1 _2163_ (.Y(_0380_),
    .A(_0350_),
    .B(_0378_));
 sg13g2_xnor2_1 _2164_ (.Y(_0381_),
    .A(_0348_),
    .B(_0380_));
 sg13g2_nor2_2 _2165_ (.A(_0347_),
    .B(_0381_),
    .Y(_0382_));
 sg13g2_and2_1 _2166_ (.A(_0347_),
    .B(_0378_),
    .X(_0383_));
 sg13g2_o21ai_1 _2167_ (.B1(_0810_),
    .Y(_0384_),
    .A1(_0382_),
    .A2(_0383_));
 sg13g2_a21oi_1 _2168_ (.A1(net185),
    .A2(\sm_i.scnt_pwm_on[1] ),
    .Y(_0385_),
    .B1(_0810_));
 sg13g2_a22oi_1 _2169_ (.Y(_0168_),
    .B1(net186),
    .B2(_0821_),
    .A2(_0384_),
    .A1(_0276_));
 sg13g2_xor2_1 _2170_ (.B(_0821_),
    .A(net292),
    .X(_0386_));
 sg13g2_nor2_1 _2171_ (.A(_0371_),
    .B(_0373_),
    .Y(_0387_));
 sg13g2_o21ai_1 _2172_ (.B1(_0357_),
    .Y(_0388_),
    .A1(_0354_),
    .A2(_0358_));
 sg13g2_and2_1 _2173_ (.A(_0367_),
    .B(_0369_),
    .X(_0389_));
 sg13g2_nor2_1 _2174_ (.A(_0039_),
    .B(_0289_),
    .Y(_0390_));
 sg13g2_nor2b_1 _2175_ (.A(_0038_),
    .B_N(_0294_),
    .Y(_0391_));
 sg13g2_and2_1 _2176_ (.A(_0390_),
    .B(_0391_),
    .X(_0392_));
 sg13g2_xnor2_1 _2177_ (.Y(_0393_),
    .A(_0390_),
    .B(_0391_));
 sg13g2_a21oi_1 _2178_ (.A1(\sm_i.adsr_i.dout[0] ),
    .A2(_0360_),
    .Y(_0394_),
    .B1(_0364_));
 sg13g2_nor2_1 _2179_ (.A(_0040_),
    .B(_0312_),
    .Y(_0395_));
 sg13g2_nor3_1 _2180_ (.A(net243),
    .B(_0317_),
    .C(_0318_),
    .Y(_0396_));
 sg13g2_nand2_1 _2181_ (.Y(_0397_),
    .A(_0042_),
    .B(net233));
 sg13g2_nor3_1 _2182_ (.A(net243),
    .B(_0319_),
    .C(_0397_),
    .Y(_0398_));
 sg13g2_nand2b_1 _2183_ (.Y(_0399_),
    .B(_0397_),
    .A_N(_0396_));
 sg13g2_xor2_1 _2184_ (.B(_0397_),
    .A(_0396_),
    .X(_0400_));
 sg13g2_xnor2_1 _2185_ (.Y(_0401_),
    .A(_0395_),
    .B(_0400_));
 sg13g2_nand2_1 _2186_ (.Y(_0402_),
    .A(_0394_),
    .B(_0401_));
 sg13g2_xnor2_1 _2187_ (.Y(_0403_),
    .A(_0394_),
    .B(_0401_));
 sg13g2_xor2_1 _2188_ (.B(_0403_),
    .A(_0393_),
    .X(_0404_));
 sg13g2_nor2b_1 _2189_ (.A(_0389_),
    .B_N(_0404_),
    .Y(_0405_));
 sg13g2_xnor2_1 _2190_ (.Y(_0406_),
    .A(_0389_),
    .B(_0404_));
 sg13g2_xnor2_1 _2191_ (.Y(_0407_),
    .A(_0388_),
    .B(_0406_));
 sg13g2_nor2_1 _2192_ (.A(_0387_),
    .B(_0407_),
    .Y(_0408_));
 sg13g2_xnor2_1 _2193_ (.Y(_0409_),
    .A(_0387_),
    .B(_0407_));
 sg13g2_o21ai_1 _2194_ (.B1(_0375_),
    .Y(_0410_),
    .A1(_0351_),
    .A2(_0376_));
 sg13g2_nand2b_1 _2195_ (.Y(_0411_),
    .B(_0410_),
    .A_N(_0409_));
 sg13g2_xor2_1 _2196_ (.B(_0410_),
    .A(_0409_),
    .X(_0412_));
 sg13g2_inv_1 _2197_ (.Y(_0413_),
    .A(_0412_));
 sg13g2_a21oi_1 _2198_ (.A1(_0349_),
    .A2(_0380_),
    .Y(_0414_),
    .B1(_0379_));
 sg13g2_a21o_1 _2199_ (.A2(_0380_),
    .A1(_0349_),
    .B1(_0379_),
    .X(_0415_));
 sg13g2_xnor2_1 _2200_ (.Y(_0416_),
    .A(_0412_),
    .B(_0414_));
 sg13g2_xnor2_1 _2201_ (.Y(_0417_),
    .A(_0382_),
    .B(_0416_));
 sg13g2_nand2_1 _2202_ (.Y(_0418_),
    .A(_0810_),
    .B(_0417_));
 sg13g2_o21ai_1 _2203_ (.B1(_0418_),
    .Y(_0169_),
    .A1(_0276_),
    .A2(net293));
 sg13g2_o21ai_1 _2204_ (.B1(net155),
    .Y(_0419_),
    .A1(\sm_i.scnt_pwm_on[2] ),
    .A2(_0821_));
 sg13g2_a21oi_1 _2205_ (.A1(_0822_),
    .A2(\sm_i.scnt_pwm_on_en ),
    .Y(_0420_),
    .B1(_0810_));
 sg13g2_a21oi_1 _2206_ (.A1(_0388_),
    .A2(_0406_),
    .Y(_0421_),
    .B1(_0405_));
 sg13g2_o21ai_1 _2207_ (.B1(_0402_),
    .Y(_0422_),
    .A1(_0393_),
    .A2(_0403_));
 sg13g2_or2_1 _2208_ (.X(_0423_),
    .B(_0289_),
    .A(_0567_));
 sg13g2_a21oi_1 _2209_ (.A1(_0395_),
    .A2(_0399_),
    .Y(_0424_),
    .B1(_0398_));
 sg13g2_nand2_1 _2210_ (.Y(_0425_),
    .A(\sm_i.adsr_i.dout[4] ),
    .B(_0311_));
 sg13g2_nor3_1 _2211_ (.A(_0040_),
    .B(_0317_),
    .C(_0318_),
    .Y(_0426_));
 sg13g2_nand2_1 _2212_ (.Y(_0427_),
    .A(net243),
    .B(_0363_));
 sg13g2_nand3_1 _2213_ (.B(net233),
    .C(_0426_),
    .A(net243),
    .Y(_0428_));
 sg13g2_xor2_1 _2214_ (.B(_0427_),
    .A(_0426_),
    .X(_0429_));
 sg13g2_xor2_1 _2215_ (.B(_0429_),
    .A(_0425_),
    .X(_0430_));
 sg13g2_nand2b_1 _2216_ (.Y(_0431_),
    .B(_0430_),
    .A_N(_0424_));
 sg13g2_xnor2_1 _2217_ (.Y(_0432_),
    .A(_0424_),
    .B(_0430_));
 sg13g2_nand2b_1 _2218_ (.Y(_0433_),
    .B(_0432_),
    .A_N(_0423_));
 sg13g2_xnor2_1 _2219_ (.Y(_0434_),
    .A(_0423_),
    .B(_0432_));
 sg13g2_nand2_1 _2220_ (.Y(_0435_),
    .A(_0422_),
    .B(_0434_));
 sg13g2_xor2_1 _2221_ (.B(_0434_),
    .A(_0422_),
    .X(_0436_));
 sg13g2_nand2_1 _2222_ (.Y(_0437_),
    .A(_0392_),
    .B(_0436_));
 sg13g2_xnor2_1 _2223_ (.Y(_0438_),
    .A(_0392_),
    .B(_0436_));
 sg13g2_nor2_1 _2224_ (.A(_0421_),
    .B(_0438_),
    .Y(_0439_));
 sg13g2_inv_1 _2225_ (.Y(_0440_),
    .A(_0439_));
 sg13g2_xor2_1 _2226_ (.B(_0438_),
    .A(_0421_),
    .X(_0441_));
 sg13g2_nand2_1 _2227_ (.Y(_0442_),
    .A(_0408_),
    .B(_0441_));
 sg13g2_inv_1 _2228_ (.Y(_0443_),
    .A(_0442_));
 sg13g2_nor2_1 _2229_ (.A(_0408_),
    .B(_0441_),
    .Y(_0444_));
 sg13g2_nor2_1 _2230_ (.A(_0443_),
    .B(_0444_),
    .Y(_0445_));
 sg13g2_o21ai_1 _2231_ (.B1(_0411_),
    .Y(_0446_),
    .A1(_0412_),
    .A2(_0414_));
 sg13g2_xnor2_1 _2232_ (.Y(_0447_),
    .A(_0445_),
    .B(_0446_));
 sg13g2_and3_1 _2233_ (.X(_0448_),
    .A(_0382_),
    .B(_0416_),
    .C(_0447_));
 sg13g2_a21oi_1 _2234_ (.A1(_0382_),
    .A2(_0416_),
    .Y(_0449_),
    .B1(_0447_));
 sg13g2_nor3_1 _2235_ (.A(_0811_),
    .B(_0448_),
    .C(_0449_),
    .Y(_0450_));
 sg13g2_a21oi_1 _2236_ (.A1(net156),
    .A2(_0420_),
    .Y(_0170_),
    .B1(_0450_));
 sg13g2_nand2_1 _2237_ (.Y(_0451_),
    .A(_0411_),
    .B(_0442_));
 sg13g2_a21oi_1 _2238_ (.A1(_0413_),
    .A2(_0415_),
    .Y(_0452_),
    .B1(_0451_));
 sg13g2_o21ai_1 _2239_ (.B1(_0428_),
    .Y(_0453_),
    .A1(_0425_),
    .A2(_0429_));
 sg13g2_nand2_1 _2240_ (.Y(_0454_),
    .A(\sm_i.adsr_i.dout[5] ),
    .B(_0311_));
 sg13g2_nand2_1 _2241_ (.Y(_0455_),
    .A(_0040_),
    .B(net233));
 sg13g2_or3_1 _2242_ (.A(_0039_),
    .B(_0319_),
    .C(_0455_),
    .X(_0456_));
 sg13g2_o21ai_1 _2243_ (.B1(_0455_),
    .Y(_0457_),
    .A1(_0039_),
    .A2(_0319_));
 sg13g2_nand2_1 _2244_ (.Y(_0458_),
    .A(_0456_),
    .B(_0457_));
 sg13g2_xor2_1 _2245_ (.B(_0458_),
    .A(_0454_),
    .X(_0459_));
 sg13g2_nand2_1 _2246_ (.Y(_0460_),
    .A(_0453_),
    .B(_0459_));
 sg13g2_xnor2_1 _2247_ (.Y(_0461_),
    .A(_0453_),
    .B(_0459_));
 sg13g2_a21o_1 _2248_ (.A2(_0433_),
    .A1(_0431_),
    .B1(_0461_),
    .X(_0462_));
 sg13g2_nand3_1 _2249_ (.B(_0433_),
    .C(_0461_),
    .A(_0431_),
    .Y(_0463_));
 sg13g2_nand2_1 _2250_ (.Y(_0464_),
    .A(_0462_),
    .B(_0463_));
 sg13g2_nand2_1 _2251_ (.Y(_0465_),
    .A(_0435_),
    .B(_0437_));
 sg13g2_a21oi_1 _2252_ (.A1(_0435_),
    .A2(_0437_),
    .Y(_0466_),
    .B1(_0464_));
 sg13g2_xor2_1 _2253_ (.B(_0465_),
    .A(_0464_),
    .X(_0467_));
 sg13g2_nor2_1 _2254_ (.A(_0440_),
    .B(_0467_),
    .Y(_0468_));
 sg13g2_xnor2_1 _2255_ (.Y(_0469_),
    .A(_0440_),
    .B(_0467_));
 sg13g2_nor3_1 _2256_ (.A(_0444_),
    .B(_0452_),
    .C(_0469_),
    .Y(_0470_));
 sg13g2_o21ai_1 _2257_ (.B1(_0469_),
    .Y(_0471_),
    .A1(_0444_),
    .A2(_0452_));
 sg13g2_nand2b_1 _2258_ (.Y(_0472_),
    .B(_0471_),
    .A_N(_0470_));
 sg13g2_xnor2_1 _2259_ (.Y(_0473_),
    .A(_0448_),
    .B(_0472_));
 sg13g2_a22oi_1 _2260_ (.Y(_0474_),
    .B1(_0473_),
    .B2(_0810_),
    .A2(_0420_),
    .A1(net153));
 sg13g2_o21ai_1 _2261_ (.B1(_0474_),
    .Y(_0171_),
    .A1(_0823_),
    .A2(_0276_));
 sg13g2_nand2_1 _2262_ (.Y(_0475_),
    .A(net174),
    .B(_0823_));
 sg13g2_a21oi_1 _2263_ (.A1(_0824_),
    .A2(\sm_i.scnt_pwm_on_en ),
    .Y(_0476_),
    .B1(_0810_));
 sg13g2_nand2_1 _2264_ (.Y(_0477_),
    .A(_0460_),
    .B(_0462_));
 sg13g2_o21ai_1 _2265_ (.B1(_0456_),
    .Y(_0478_),
    .A1(_0454_),
    .A2(_0458_));
 sg13g2_or2_1 _2266_ (.X(_0479_),
    .B(_0319_),
    .A(_0567_));
 sg13g2_nand2_1 _2267_ (.Y(_0480_),
    .A(_0039_),
    .B(net233));
 sg13g2_nor2_1 _2268_ (.A(_0479_),
    .B(_0480_),
    .Y(_0481_));
 sg13g2_xor2_1 _2269_ (.B(_0480_),
    .A(_0479_),
    .X(_0482_));
 sg13g2_nand2_1 _2270_ (.Y(_0483_),
    .A(_0478_),
    .B(_0482_));
 sg13g2_xnor2_1 _2271_ (.Y(_0484_),
    .A(_0478_),
    .B(_0482_));
 sg13g2_xor2_1 _2272_ (.B(_0484_),
    .A(_0477_),
    .X(_0485_));
 sg13g2_inv_1 _2273_ (.Y(_0486_),
    .A(_0485_));
 sg13g2_nand2_1 _2274_ (.Y(_0487_),
    .A(_0466_),
    .B(_0486_));
 sg13g2_xnor2_1 _2275_ (.Y(_0488_),
    .A(_0466_),
    .B(_0485_));
 sg13g2_nor3_1 _2276_ (.A(_0468_),
    .B(_0470_),
    .C(_0488_),
    .Y(_0489_));
 sg13g2_o21ai_1 _2277_ (.B1(_0488_),
    .Y(_0490_),
    .A1(_0468_),
    .A2(_0470_));
 sg13g2_nand2b_1 _2278_ (.Y(_0491_),
    .B(_0490_),
    .A_N(_0489_));
 sg13g2_a21oi_1 _2279_ (.A1(_0448_),
    .A2(_0472_),
    .Y(_0492_),
    .B1(_0491_));
 sg13g2_nand3_1 _2280_ (.B(_0472_),
    .C(_0491_),
    .A(_0448_),
    .Y(_0493_));
 sg13g2_nor2_1 _2281_ (.A(_0811_),
    .B(_0492_),
    .Y(_0494_));
 sg13g2_a22oi_1 _2282_ (.Y(_0172_),
    .B1(_0493_),
    .B2(_0494_),
    .A2(_0476_),
    .A1(_0475_));
 sg13g2_nor2_1 _2283_ (.A(_0462_),
    .B(_0484_),
    .Y(_0495_));
 sg13g2_a21oi_1 _2284_ (.A1(_0038_),
    .A2(net233),
    .Y(_0496_),
    .B1(_0481_));
 sg13g2_a21o_1 _2285_ (.A2(_0481_),
    .A1(_0038_),
    .B1(_0496_),
    .X(_0497_));
 sg13g2_inv_1 _2286_ (.Y(_0498_),
    .A(_0497_));
 sg13g2_o21ai_1 _2287_ (.B1(_0483_),
    .Y(_0499_),
    .A1(_0460_),
    .A2(_0484_));
 sg13g2_xnor2_1 _2288_ (.Y(_0500_),
    .A(_0498_),
    .B(_0499_));
 sg13g2_or3_1 _2289_ (.A(_0462_),
    .B(_0484_),
    .C(_0500_),
    .X(_0501_));
 sg13g2_xor2_1 _2290_ (.B(_0500_),
    .A(_0495_),
    .X(_0502_));
 sg13g2_a21oi_1 _2291_ (.A1(_0487_),
    .A2(_0490_),
    .Y(_0503_),
    .B1(_0502_));
 sg13g2_nand3_1 _2292_ (.B(_0490_),
    .C(_0502_),
    .A(_0487_),
    .Y(_0504_));
 sg13g2_nor2b_1 _2293_ (.A(_0503_),
    .B_N(_0504_),
    .Y(_0505_));
 sg13g2_nor2_1 _2294_ (.A(_0493_),
    .B(_0505_),
    .Y(_0506_));
 sg13g2_xor2_1 _2295_ (.B(_0505_),
    .A(_0493_),
    .X(_0507_));
 sg13g2_nor2b_1 _2296_ (.A(_0824_),
    .B_N(net204),
    .Y(_0508_));
 sg13g2_o21ai_1 _2297_ (.B1(_0277_),
    .Y(_0509_),
    .A1(_0825_),
    .A2(_0508_));
 sg13g2_o21ai_1 _2298_ (.B1(_0509_),
    .Y(_0173_),
    .A1(_0811_),
    .A2(_0507_));
 sg13g2_nand3b_1 _2299_ (.B(net85),
    .C(_0811_),
    .Y(_0510_),
    .A_N(_0825_));
 sg13g2_a22oi_1 _2300_ (.Y(_0511_),
    .B1(_0498_),
    .B2(_0499_),
    .A2(_0481_),
    .A1(_0038_));
 sg13g2_nand3_1 _2301_ (.B(_0501_),
    .C(_0511_),
    .A(net233),
    .Y(_0512_));
 sg13g2_o21ai_1 _2302_ (.B1(_0810_),
    .Y(_0513_),
    .A1(_0503_),
    .A2(_0512_));
 sg13g2_o21ai_1 _2303_ (.B1(net86),
    .Y(_0174_),
    .A1(_0506_),
    .A2(_0513_));
 sg13g2_o21ai_1 _2304_ (.B1(_0814_),
    .Y(_0514_),
    .A1(\sm_i.adsr_i.sstate[2] ),
    .A2(_0816_));
 sg13g2_nand2b_1 _2305_ (.Y(_0515_),
    .B(_0514_),
    .A_N(_0185_));
 sg13g2_nand2_1 _2306_ (.Y(_0516_),
    .A(_0852_),
    .B(_0515_));
 sg13g2_or2_1 _2307_ (.X(_0517_),
    .B(_0514_),
    .A(_0840_));
 sg13g2_o21ai_1 _2308_ (.B1(_0517_),
    .Y(_0518_),
    .A1(_0837_),
    .A2(_0515_));
 sg13g2_a221oi_1 _2309_ (.B2(_0516_),
    .C1(_0518_),
    .B1(_0980_),
    .A1(_0846_),
    .Y(_0519_),
    .A2(net234));
 sg13g2_nor2_1 _2310_ (.A(net304),
    .B(_0185_),
    .Y(_0520_));
 sg13g2_nand2_1 _2311_ (.Y(_0521_),
    .A(_0519_),
    .B(_0520_));
 sg13g2_o21ai_1 _2312_ (.B1(_0521_),
    .Y(_0175_),
    .A1(_0564_),
    .A2(net215));
 sg13g2_nor2_1 _2313_ (.A(_0563_),
    .B(net235),
    .Y(_0522_));
 sg13g2_xnor2_1 _2314_ (.Y(_0523_),
    .A(\sm_i.adsr_i.dout[1] ),
    .B(net235));
 sg13g2_xnor2_1 _2315_ (.Y(_0524_),
    .A(\sm_i.adsr_i.dout[0] ),
    .B(_0523_));
 sg13g2_nor2_1 _2316_ (.A(_0185_),
    .B(_0524_),
    .Y(_0525_));
 sg13g2_mux2_1 _2317_ (.A0(net163),
    .A1(_0525_),
    .S(net215),
    .X(_0176_));
 sg13g2_a21oi_1 _2318_ (.A1(net311),
    .A2(_0523_),
    .Y(_0526_),
    .B1(_0522_));
 sg13g2_xnor2_1 _2319_ (.Y(_0527_),
    .A(_0566_),
    .B(net235));
 sg13g2_or2_1 _2320_ (.X(_0528_),
    .B(_0527_),
    .A(_0526_));
 sg13g2_a21oi_1 _2321_ (.A1(_0526_),
    .A2(_0527_),
    .Y(_0529_),
    .B1(_0185_));
 sg13g2_nand3_1 _2322_ (.B(_0528_),
    .C(_0529_),
    .A(net215),
    .Y(_0530_));
 sg13g2_o21ai_1 _2323_ (.B1(_0530_),
    .Y(_0177_),
    .A1(_0566_),
    .A2(_0519_));
 sg13g2_o21ai_1 _2324_ (.B1(_0528_),
    .Y(_0531_),
    .A1(net243),
    .A2(net235));
 sg13g2_xnor2_1 _2325_ (.Y(_0532_),
    .A(\sm_i.adsr_i.dout[3] ),
    .B(net235));
 sg13g2_nand2_1 _2326_ (.Y(_0533_),
    .A(_0531_),
    .B(_0532_));
 sg13g2_nor2_1 _2327_ (.A(_0531_),
    .B(_0532_),
    .Y(_0534_));
 sg13g2_nor2_1 _2328_ (.A(_0185_),
    .B(_0534_),
    .Y(_0535_));
 sg13g2_nand3_1 _2329_ (.B(_0533_),
    .C(_0535_),
    .A(net215),
    .Y(_0536_));
 sg13g2_o21ai_1 _2330_ (.B1(_0536_),
    .Y(_0178_),
    .A1(_0565_),
    .A2(_0519_));
 sg13g2_xor2_1 _2331_ (.B(net234),
    .A(_0039_),
    .X(_0537_));
 sg13g2_o21ai_1 _2332_ (.B1(_0533_),
    .Y(_0538_),
    .A1(_0040_),
    .A2(net234));
 sg13g2_nand2_1 _2333_ (.Y(_0539_),
    .A(_0537_),
    .B(_0538_));
 sg13g2_nor2_1 _2334_ (.A(_0537_),
    .B(_0538_),
    .Y(_0540_));
 sg13g2_nor2_1 _2335_ (.A(_0185_),
    .B(_0540_),
    .Y(_0541_));
 sg13g2_nand3_1 _2336_ (.B(_0539_),
    .C(_0541_),
    .A(net215),
    .Y(_0542_));
 sg13g2_o21ai_1 _2337_ (.B1(_0542_),
    .Y(_0179_),
    .A1(_0568_),
    .A2(net215));
 sg13g2_o21ai_1 _2338_ (.B1(_0539_),
    .Y(_0543_),
    .A1(_0039_),
    .A2(net234));
 sg13g2_xnor2_1 _2339_ (.Y(_0544_),
    .A(_0038_),
    .B(net234));
 sg13g2_xnor2_1 _2340_ (.Y(_0545_),
    .A(_0543_),
    .B(_0544_));
 sg13g2_nand3b_1 _2341_ (.B(net215),
    .C(_0545_),
    .Y(_0546_),
    .A_N(_0185_));
 sg13g2_o21ai_1 _2342_ (.B1(_0546_),
    .Y(_0180_),
    .A1(_0567_),
    .A2(net215));
 sg13g2_nor2_1 _2343_ (.A(_0981_),
    .B(_0187_),
    .Y(_0547_));
 sg13g2_or2_1 _2344_ (.X(_0548_),
    .B(_0547_),
    .A(_0186_));
 sg13g2_inv_1 _2345_ (.Y(_0549_),
    .A(_0548_));
 sg13g2_nand2b_1 _2346_ (.Y(_0550_),
    .B(_0855_),
    .A_N(_0186_));
 sg13g2_o21ai_1 _2347_ (.B1(_0548_),
    .Y(_0551_),
    .A1(net279),
    .A2(_0550_));
 sg13g2_o21ai_1 _2348_ (.B1(_0551_),
    .Y(_0552_),
    .A1(net279),
    .A2(_0547_));
 sg13g2_inv_1 _2349_ (.Y(_0181_),
    .A(_0552_));
 sg13g2_nand2_1 _2350_ (.Y(_0553_),
    .A(net280),
    .B(_0549_));
 sg13g2_a21oi_1 _2351_ (.A1(_0582_),
    .A2(_0854_),
    .Y(_0554_),
    .B1(_0861_));
 sg13g2_nand2b_1 _2352_ (.Y(_0555_),
    .B(_0190_),
    .A_N(_0554_));
 sg13g2_o21ai_1 _2353_ (.B1(_0553_),
    .Y(_0182_),
    .A1(_0981_),
    .A2(_0555_));
 sg13g2_nand3_1 _2354_ (.B(net242),
    .C(_0548_),
    .A(net280),
    .Y(_0556_));
 sg13g2_a22oi_1 _2355_ (.Y(_0183_),
    .B1(_0556_),
    .B2(_0582_),
    .A2(_0550_),
    .A1(_0548_));
 sg13g2_dfrbp_1 _2356_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net272),
    .D(net55),
    .Q_N(_1204_),
    .Q(pwm_out_right));
 sg13g2_dfrbp_1 _2357_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net255),
    .D(_0032_),
    .Q_N(_1205_),
    .Q(\sm_i.wav_gen_1.rom_ampl_sin_i.data_out[0] ));
 sg13g2_dfrbp_1 _2358_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net255),
    .D(_0033_),
    .Q_N(_1206_),
    .Q(\sm_i.wav_gen_1.rom_ampl_sin_i.data_out[1] ));
 sg13g2_dfrbp_1 _2359_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net254),
    .D(_0034_),
    .Q_N(_0067_),
    .Q(\sm_i.wav_gen_1.rom_ampl_sin_i.data_out[2] ));
 sg13g2_dfrbp_1 _2360_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net254),
    .D(_0035_),
    .Q_N(_0068_),
    .Q(\sm_i.wav_gen_1.rom_ampl_sin_i.data_out[3] ));
 sg13g2_dfrbp_1 _2361_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net255),
    .D(_0036_),
    .Q_N(_0069_),
    .Q(\sm_i.wav_gen_1.rom_ampl_sin_i.data_out[4] ));
 sg13g2_dfrbp_1 _2362_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net249),
    .D(net65),
    .Q_N(_1203_),
    .Q(\sm_i.wav_gen_1.rom_ampl_sin_i.en ));
 sg13g2_dfrbp_1 _2363_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net249),
    .D(net132),
    .Q_N(_1207_),
    .Q(\sm_i.wav_gen_1.swave_squ_sel ));
 sg13g2_dfrbp_1 _2364_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net264),
    .D(net226),
    .Q_N(_1208_),
    .Q(\sm_i.wav_gen_1.snote_enable ));
 sg13g2_dfrbp_1 _2365_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net258),
    .D(net66),
    .Q_N(_0070_),
    .Q(\sm_i.wav_gen_1.swave_squ[0] ));
 sg13g2_dfrbp_1 _2366_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net258),
    .D(_0030_),
    .Q_N(_0071_),
    .Q(\sm_i.wav_gen_1.swave_squ[1] ));
 sg13g2_dfrbp_1 _2367_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net254),
    .D(_0031_),
    .Q_N(_0072_),
    .Q(\sm_i.wav_gen_1.swave_squ[5] ));
 sg13g2_dfrbp_1 _2368_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net268),
    .D(_0008_),
    .Q_N(_1209_),
    .Q(\sm_i.wav_gen_1.sstep_cnt[0] ));
 sg13g2_dfrbp_1 _2369_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net265),
    .D(_0015_),
    .Q_N(_1210_),
    .Q(\sm_i.wav_gen_1.sstep_cnt[1] ));
 sg13g2_dfrbp_1 _2370_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net265),
    .D(_0016_),
    .Q_N(_0073_),
    .Q(\sm_i.wav_gen_1.sstep_cnt[2] ));
 sg13g2_dfrbp_1 _2371_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net265),
    .D(net139),
    .Q_N(_1211_),
    .Q(\sm_i.wav_gen_1.sstep_cnt[3] ));
 sg13g2_dfrbp_1 _2372_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net265),
    .D(_0018_),
    .Q_N(_0074_),
    .Q(\sm_i.wav_gen_1.sstep_cnt[4] ));
 sg13g2_dfrbp_1 _2373_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net265),
    .D(_0019_),
    .Q_N(_0075_),
    .Q(\sm_i.wav_gen_1.sstep_cnt[5] ));
 sg13g2_dfrbp_1 _2374_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net265),
    .D(_0020_),
    .Q_N(_0076_),
    .Q(\sm_i.wav_gen_1.sstep_cnt[6] ));
 sg13g2_dfrbp_1 _2375_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net265),
    .D(net161),
    .Q_N(_1212_),
    .Q(\sm_i.wav_gen_1.sstep_cnt[7] ));
 sg13g2_dfrbp_1 _2376_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net265),
    .D(_0022_),
    .Q_N(_0077_),
    .Q(\sm_i.wav_gen_1.sstep_cnt[8] ));
 sg13g2_dfrbp_1 _2377_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net261),
    .D(_0023_),
    .Q_N(_0078_),
    .Q(\sm_i.wav_gen_1.sstep_cnt[9] ));
 sg13g2_dfrbp_1 _2378_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net262),
    .D(_0009_),
    .Q_N(_0079_),
    .Q(\sm_i.wav_gen_1.sstep_cnt[10] ));
 sg13g2_dfrbp_1 _2379_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net261),
    .D(net297),
    .Q_N(_1213_),
    .Q(\sm_i.wav_gen_1.sstep_cnt[11] ));
 sg13g2_dfrbp_1 _2380_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net262),
    .D(net208),
    .Q_N(_0080_),
    .Q(\sm_i.wav_gen_1.sstep_cnt[12] ));
 sg13g2_dfrbp_1 _2381_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net262),
    .D(_0012_),
    .Q_N(_0081_),
    .Q(\sm_i.wav_gen_1.sstep_cnt[13] ));
 sg13g2_dfrbp_1 _2382_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net262),
    .D(_0013_),
    .Q_N(_0082_),
    .Q(\sm_i.wav_gen_1.sstep_cnt[14] ));
 sg13g2_dfrbp_1 _2383_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net264),
    .D(_0014_),
    .Q_N(_1202_),
    .Q(\sm_i.wav_gen_1.sstep_cnt[15] ));
 sg13g2_dfrbp_1 _2384_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net253),
    .D(net288),
    .Q_N(_0083_),
    .Q(\sm_i.wav_gen_1.swave_cnt_tri_down_up_n ));
 sg13g2_dfrbp_1 _2385_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net254),
    .D(net245),
    .Q_N(_0066_),
    .Q(\sm_i.wav_gen_1.smem_rom_ampl_sin_val_is_neg ));
 sg13g2_dfrbp_1 _2386_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net263),
    .D(net286),
    .Q_N(_1201_),
    .Q(\sm_i.adsr_i.sstate[0] ));
 sg13g2_dfrbp_1 _2387_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net263),
    .D(net290),
    .Q_N(_1200_),
    .Q(\sm_i.adsr_i.sstate[1] ));
 sg13g2_dfrbp_1 _2388_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net263),
    .D(net198),
    .Q_N(_0084_),
    .Q(\sm_i.adsr_i.sstate[2] ));
 sg13g2_dfrbp_1 _2389_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net254),
    .D(_0024_),
    .Q_N(_1214_),
    .Q(\sm_i.wav_gen_1.swave_saw[0] ));
 sg13g2_dfrbp_1 _2390_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net257),
    .D(_0025_),
    .Q_N(_1215_),
    .Q(\sm_i.wav_gen_1.swave_saw[1] ));
 sg13g2_dfrbp_1 _2391_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net254),
    .D(_0026_),
    .Q_N(_1216_),
    .Q(\sm_i.wav_gen_1.swave_saw[2] ));
 sg13g2_dfrbp_1 _2392_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net258),
    .D(_0027_),
    .Q_N(_1217_),
    .Q(\sm_i.wav_gen_1.swave_saw[3] ));
 sg13g2_dfrbp_1 _2393_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net258),
    .D(_0028_),
    .Q_N(_1218_),
    .Q(\sm_i.wav_gen_1.swave_saw[4] ));
 sg13g2_dfrbp_1 _2394_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net257),
    .D(_0029_),
    .Q_N(_1199_),
    .Q(\sm_i.wav_gen_1.swave_saw[5] ));
 sg13g2_dfrbp_1 _2395_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net267),
    .D(_0109_),
    .Q_N(_1198_),
    .Q(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[0] ));
 sg13g2_dfrbp_1 _2396_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net266),
    .D(_0110_),
    .Q_N(_1197_),
    .Q(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[1] ));
 sg13g2_dfrbp_1 _2397_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net267),
    .D(_0111_),
    .Q_N(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[2] ),
    .Q(_0088_));
 sg13g2_dfrbp_1 _2398_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net267),
    .D(_0112_),
    .Q_N(_1196_),
    .Q(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[3] ));
 sg13g2_dfrbp_1 _2399_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net276),
    .D(_0113_),
    .Q_N(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[4] ),
    .Q(_0089_));
 sg13g2_dfrbp_1 _2400_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net276),
    .D(_0114_),
    .Q_N(_1195_),
    .Q(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[5] ));
 sg13g2_dfrbp_1 _2401_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net276),
    .D(_0115_),
    .Q_N(_1194_),
    .Q(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[6] ));
 sg13g2_dfrbp_1 _2402_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net266),
    .D(_0116_),
    .Q_N(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[7] ),
    .Q(_0090_));
 sg13g2_dfrbp_1 _2403_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net266),
    .D(_0117_),
    .Q_N(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[8] ),
    .Q(_0091_));
 sg13g2_dfrbp_1 _2404_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net263),
    .D(_0118_),
    .Q_N(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[9] ),
    .Q(_0092_));
 sg13g2_dfrbp_1 _2405_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net269),
    .D(_0119_),
    .Q_N(_1193_),
    .Q(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[10] ));
 sg13g2_dfrbp_1 _2406_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net254),
    .D(_0120_),
    .Q_N(_0065_),
    .Q(\sm_i.wav_gen_1.rom_ampl_sin_i.addr[0] ));
 sg13g2_dfrbp_1 _2407_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net253),
    .D(net283),
    .Q_N(_0064_),
    .Q(\sm_i.wav_gen_1.swave_cnt_tri[1] ));
 sg13g2_dfrbp_1 _2408_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net254),
    .D(_0122_),
    .Q_N(_0063_),
    .Q(\sm_i.wav_gen_1.swave_cnt_tri[2] ));
 sg13g2_dfrbp_1 _2409_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net249),
    .D(_0123_),
    .Q_N(_0062_),
    .Q(\sm_i.wav_gen_1.swave_cnt_tri[3] ));
 sg13g2_dfrbp_1 _2410_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net249),
    .D(_0124_),
    .Q_N(_0061_),
    .Q(\sm_i.wav_gen_1.swave_cnt_tri[4] ));
 sg13g2_dfrbp_1 _2411_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net249),
    .D(_0125_),
    .Q_N(_0060_),
    .Q(\sm_i.wav_gen_1.swave_cnt_tri[5] ));
 sg13g2_dfrbp_1 _2412_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net266),
    .D(_0126_),
    .Q_N(_1192_),
    .Q(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[0] ));
 sg13g2_dfrbp_1 _2413_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net267),
    .D(_0127_),
    .Q_N(_1191_),
    .Q(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[1] ));
 sg13g2_dfrbp_1 _2414_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net266),
    .D(_0128_),
    .Q_N(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[2] ),
    .Q(_0093_));
 sg13g2_dfrbp_1 _2415_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net266),
    .D(_0129_),
    .Q_N(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[3] ),
    .Q(_0094_));
 sg13g2_dfrbp_1 _2416_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net276),
    .D(_0130_),
    .Q_N(_1190_),
    .Q(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[4] ));
 sg13g2_dfrbp_1 _2417_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net267),
    .D(_0131_),
    .Q_N(_1189_),
    .Q(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[5] ));
 sg13g2_dfrbp_1 _2418_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net276),
    .D(_0132_),
    .Q_N(_1188_),
    .Q(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[6] ));
 sg13g2_dfrbp_1 _2419_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net276),
    .D(_0133_),
    .Q_N(_1187_),
    .Q(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[7] ));
 sg13g2_dfrbp_1 _2420_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net266),
    .D(_0134_),
    .Q_N(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[8] ),
    .Q(_0095_));
 sg13g2_dfrbp_1 _2421_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net263),
    .D(_0135_),
    .Q_N(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[9] ),
    .Q(_0096_));
 sg13g2_dfrbp_1 _2422_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net269),
    .D(_0136_),
    .Q_N(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[10] ),
    .Q(_0097_));
 sg13g2_dfrbp_1 _2423_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net266),
    .D(_0137_),
    .Q_N(_1186_),
    .Q(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[11] ));
 sg13g2_dfrbp_1 _2424_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net264),
    .D(_0138_),
    .Q_N(_0059_),
    .Q(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[12] ));
 sg13g2_dfrbp_1 _2425_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net249),
    .D(_0139_),
    .Q_N(_1185_),
    .Q(\sm_i.adsr_i.scnt_step[0] ));
 sg13g2_dfrbp_1 _2426_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net250),
    .D(_0140_),
    .Q_N(_1184_),
    .Q(\sm_i.adsr_i.scnt_step[1] ));
 sg13g2_dfrbp_1 _2427_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net249),
    .D(net80),
    .Q_N(_0058_),
    .Q(\sm_i.adsr_i.scnt_step[2] ));
 sg13g2_dfrbp_1 _2428_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net249),
    .D(net95),
    .Q_N(_0057_),
    .Q(\sm_i.adsr_i.scnt_step[3] ));
 sg13g2_dfrbp_1 _2429_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net251),
    .D(net93),
    .Q_N(_0056_),
    .Q(\sm_i.adsr_i.scnt_step[4] ));
 sg13g2_dfrbp_1 _2430_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net251),
    .D(net101),
    .Q_N(_0055_),
    .Q(\sm_i.adsr_i.scnt_step[5] ));
 sg13g2_dfrbp_1 _2431_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net250),
    .D(net116),
    .Q_N(_0054_),
    .Q(\sm_i.adsr_i.scnt_step[6] ));
 sg13g2_dfrbp_1 _2432_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net251),
    .D(net119),
    .Q_N(_0053_),
    .Q(\sm_i.adsr_i.scnt_step[7] ));
 sg13g2_dfrbp_1 _2433_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net250),
    .D(net91),
    .Q_N(_0052_),
    .Q(\sm_i.adsr_i.scnt_step[8] ));
 sg13g2_dfrbp_1 _2434_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net250),
    .D(net98),
    .Q_N(_0051_),
    .Q(\sm_i.adsr_i.scnt_step[9] ));
 sg13g2_dfrbp_1 _2435_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net251),
    .D(_0149_),
    .Q_N(_1183_),
    .Q(\sm_i.adsr_i.scnt_step[10] ));
 sg13g2_dfrbp_1 _2436_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net250),
    .D(net134),
    .Q_N(_0050_),
    .Q(\sm_i.adsr_i.scnt_step[11] ));
 sg13g2_dfrbp_1 _2437_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net250),
    .D(net104),
    .Q_N(_0049_),
    .Q(\sm_i.adsr_i.scnt_step[12] ));
 sg13g2_dfrbp_1 _2438_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net250),
    .D(net109),
    .Q_N(_0048_),
    .Q(\sm_i.adsr_i.scnt_step[13] ));
 sg13g2_dfrbp_1 _2439_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net251),
    .D(net122),
    .Q_N(_0047_),
    .Q(\sm_i.adsr_i.scnt_step[14] ));
 sg13g2_dfrbp_1 _2440_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net251),
    .D(net111),
    .Q_N(_0046_),
    .Q(\sm_i.adsr_i.scnt_step[15] ));
 sg13g2_dfrbp_1 _2441_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net251),
    .D(net200),
    .Q_N(_1182_),
    .Q(\sm_i.adsr_i.scnt_step[16] ));
 sg13g2_dfrbp_1 _2442_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net252),
    .D(net166),
    .Q_N(_0045_),
    .Q(\sm_i.adsr_i.scnt_step[17] ));
 sg13g2_dfrbp_1 _2443_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net251),
    .D(_0157_),
    .Q_N(_1181_),
    .Q(\sm_i.adsr_i.scnt_step[18] ));
 sg13g2_dfrbp_1 _2444_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net261),
    .D(_0158_),
    .Q_N(_1180_),
    .Q(\sm_i.adsr_i.scnt_step[19] ));
 sg13g2_dfrbp_1 _2445_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net261),
    .D(net145),
    .Q_N(_1179_),
    .Q(\sm_i.adsr_i.scnt_step[20] ));
 sg13g2_dfrbp_1 _2446_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net261),
    .D(net195),
    .Q_N(_1178_),
    .Q(\sm_i.adsr_i.scnt_step[21] ));
 sg13g2_dfrbp_1 _2447_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net261),
    .D(_0161_),
    .Q_N(_1177_),
    .Q(\sm_i.adsr_i.scnt_step[22] ));
 sg13g2_dfrbp_1 _2448_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net261),
    .D(net184),
    .Q_N(_1176_),
    .Q(\sm_i.adsr_i.scnt_step[23] ));
 sg13g2_dfrbp_1 _2449_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net261),
    .D(_0163_),
    .Q_N(_1175_),
    .Q(\sm_i.adsr_i.scnt_step[24] ));
 sg13g2_dfrbp_1 _2450_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net263),
    .D(_0164_),
    .Q_N(_1174_),
    .Q(\sm_i.adsr_i.scnt_step[25] ));
 sg13g2_dfrbp_1 _2451_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net263),
    .D(net107),
    .Q_N(_1173_),
    .Q(\sm_i.adsr_i.scnt_step[26] ));
 sg13g2_dfrbp_1 _2452_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net263),
    .D(_0166_),
    .Q_N(_1172_),
    .Q(\sm_i.adsr_i.scnt_step[27] ));
 sg13g2_dfrbp_1 _2453_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net259),
    .D(net64),
    .Q_N(_0044_),
    .Q(\sm_i.scnt_pwm_on[0] ));
 sg13g2_dfrbp_1 _2454_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net259),
    .D(net187),
    .Q_N(_1171_),
    .Q(\sm_i.scnt_pwm_on[1] ));
 sg13g2_dfrbp_1 _2455_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net259),
    .D(_0169_),
    .Q_N(_1170_),
    .Q(\sm_i.scnt_pwm_on[2] ));
 sg13g2_dfrbp_1 _2456_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net259),
    .D(net157),
    .Q_N(_1169_),
    .Q(\sm_i.scnt_pwm_on[3] ));
 sg13g2_dfrbp_1 _2457_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net258),
    .D(net154),
    .Q_N(_1168_),
    .Q(\sm_i.scnt_pwm_on[4] ));
 sg13g2_dfrbp_1 _2458_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net256),
    .D(_0172_),
    .Q_N(_1167_),
    .Q(\sm_i.scnt_pwm_on[5] ));
 sg13g2_dfrbp_1 _2459_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net256),
    .D(_0173_),
    .Q_N(_1166_),
    .Q(\sm_i.scnt_pwm_on[6] ));
 sg13g2_dfrbp_1 _2460_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net256),
    .D(net87),
    .Q_N(_1165_),
    .Q(\sm_i.scnt_pwm_on[7] ));
 sg13g2_dfrbp_1 _2461_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net269),
    .D(_0175_),
    .Q_N(_0043_),
    .Q(\sm_i.adsr_i.dout[0] ));
 sg13g2_dfrbp_1 _2462_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net269),
    .D(net164),
    .Q_N(_0042_),
    .Q(\sm_i.adsr_i.dout[1] ));
 sg13g2_dfrbp_1 _2463_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net269),
    .D(_0177_),
    .Q_N(_0041_),
    .Q(\sm_i.adsr_i.dout[2] ));
 sg13g2_dfrbp_1 _2464_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net258),
    .D(_0178_),
    .Q_N(_0040_),
    .Q(\sm_i.adsr_i.dout[3] ));
 sg13g2_dfrbp_1 _2465_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net258),
    .D(_0179_),
    .Q_N(_0039_),
    .Q(\sm_i.adsr_i.dout[4] ));
 sg13g2_dfrbp_1 _2466_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net258),
    .D(_0180_),
    .Q_N(_0038_),
    .Q(\sm_i.adsr_i.dout[5] ));
 sg13g2_dfrbp_1 _2467_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net252),
    .D(_0181_),
    .Q_N(_1164_),
    .Q(\sm_i.adsr_i.scnt_pwl[0] ));
 sg13g2_dfrbp_1 _2468_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net252),
    .D(_0182_),
    .Q_N(_0037_),
    .Q(\sm_i.adsr_i.scnt_pwl[1] ));
 sg13g2_dfrbp_1 _2469_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net252),
    .D(net300),
    .Q_N(_0085_),
    .Q(\sm_i.adsr_i.scnt_pwl[2] ));
 sg13g2_dfrbp_1 _2470_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net276),
    .D(net6),
    .Q_N(_1219_),
    .Q(\sm_i.ssw_reg[0][0] ));
 sg13g2_dfrbp_1 _2471_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net270),
    .D(net7),
    .Q_N(_1220_),
    .Q(\sm_i.ssw_reg[0][1] ));
 sg13g2_dfrbp_1 _2472_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net271),
    .D(net8),
    .Q_N(_1221_),
    .Q(\sm_i.ssw_reg[0][2] ));
 sg13g2_dfrbp_1 _2473_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net270),
    .D(net9),
    .Q_N(_1222_),
    .Q(\sm_i.ssw_reg[0][3] ));
 sg13g2_dfrbp_1 _2474_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net270),
    .D(net10),
    .Q_N(_1223_),
    .Q(\sm_i.ssw_reg[0][4] ));
 sg13g2_dfrbp_1 _2475_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net270),
    .D(net11),
    .Q_N(_1224_),
    .Q(\sm_i.ssw_reg[0][5] ));
 sg13g2_dfrbp_1 _2476_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net270),
    .D(net12),
    .Q_N(_1225_),
    .Q(\sm_i.ssw_reg[0][6] ));
 sg13g2_dfrbp_1 _2477_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net270),
    .D(net13),
    .Q_N(_1226_),
    .Q(\sm_i.ssw_reg[0][7] ));
 sg13g2_dfrbp_1 _2478_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net269),
    .D(net57),
    .Q_N(_1227_),
    .Q(\sm_i.ssw_reg[2][0] ));
 sg13g2_dfrbp_1 _2479_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net272),
    .D(net44),
    .Q_N(_1228_),
    .Q(\sm_i.ssw_reg[2][1] ));
 sg13g2_dfrbp_1 _2480_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net272),
    .D(net62),
    .Q_N(_1229_),
    .Q(\sm_i.sadsr_sel[0] ));
 sg13g2_dfrbp_1 _2481_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net271),
    .D(net51),
    .Q_N(_1230_),
    .Q(\sm_i.sadsr_sel[1] ));
 sg13g2_dfrbp_1 _2482_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net273),
    .D(net49),
    .Q_N(_1231_),
    .Q(\sm_i.snotes_sel[0] ));
 sg13g2_dfrbp_1 _2483_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net273),
    .D(net42),
    .Q_N(_1232_),
    .Q(\sm_i.snotes_sel[1] ));
 sg13g2_dfrbp_1 _2484_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net273),
    .D(net43),
    .Q_N(_1233_),
    .Q(\sm_i.snotes_sel[2] ));
 sg13g2_dfrbp_1 _2485_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net273),
    .D(net41),
    .Q_N(_1234_),
    .Q(\sm_i.snotes_sel[3] ));
 sg13g2_dfrbp_1 _2486_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net255),
    .D(_0000_),
    .Q_N(_1235_),
    .Q(\sm_i.scnt_pwm[0] ));
 sg13g2_dfrbp_1 _2487_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net255),
    .D(_0001_),
    .Q_N(_1236_),
    .Q(\sm_i.scnt_pwm[1] ));
 sg13g2_dfrbp_1 _2488_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net255),
    .D(_0002_),
    .Q_N(_1237_),
    .Q(\sm_i.scnt_pwm[2] ));
 sg13g2_dfrbp_1 _2489_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net256),
    .D(net89),
    .Q_N(_1238_),
    .Q(\sm_i.scnt_pwm[3] ));
 sg13g2_dfrbp_1 _2490_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net256),
    .D(net82),
    .Q_N(_1239_),
    .Q(\sm_i.scnt_pwm[4] ));
 sg13g2_dfrbp_1 _2491_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net255),
    .D(_0005_),
    .Q_N(_1240_),
    .Q(\sm_i.scnt_pwm[5] ));
 sg13g2_dfrbp_1 _2492_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net255),
    .D(net74),
    .Q_N(_1241_),
    .Q(\sm_i.scnt_pwm[6] ));
 sg13g2_dfrbp_1 _2493_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net256),
    .D(_0007_),
    .Q_N(_1163_),
    .Q(\sm_i.scnt_pwm[7] ));
 sg13g2_dfrbp_1 _2494_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net275),
    .D(_0101_),
    .Q_N(\sm_i.snote_synch[0][0] ),
    .Q(_0098_));
 sg13g2_dfrbp_1 _2495_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net274),
    .D(net2),
    .Q_N(_1242_),
    .Q(\sm_i.snote_synch[0][1] ));
 sg13g2_dfrbp_1 _2496_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net274),
    .D(net3),
    .Q_N(_1243_),
    .Q(\sm_i.snote_synch[0][2] ));
 sg13g2_dfrbp_1 _2497_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net273),
    .D(net4),
    .Q_N(_1244_),
    .Q(\sm_i.snote_synch[0][3] ));
 sg13g2_dfrbp_1 _2498_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net273),
    .D(net5),
    .Q_N(_1245_),
    .Q(\sm_i.snote_synch[0][4] ));
 sg13g2_dfrbp_1 _2499_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net272),
    .D(\sm_i.scnt_pwm_on_en ),
    .Q_N(_1162_),
    .Q(pwm_out_i));
 sg13g2_dfrbp_1 _2500_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net274),
    .D(_0102_),
    .Q_N(\sm_i.snote_synch[1][0] ),
    .Q(_0099_));
 sg13g2_dfrbp_1 _2501_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net274),
    .D(net53),
    .Q_N(_1246_),
    .Q(\sm_i.snote_synch[1][1] ));
 sg13g2_dfrbp_1 _2502_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net274),
    .D(net59),
    .Q_N(_1247_),
    .Q(\sm_i.snote_synch[1][2] ));
 sg13g2_dfrbp_1 _2503_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net274),
    .D(net36),
    .Q_N(_1248_),
    .Q(\sm_i.snote_synch[1][3] ));
 sg13g2_dfrbp_1 _2504_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net274),
    .D(net37),
    .Q_N(_1249_),
    .Q(\sm_i.snote_synch[1][4] ));
 sg13g2_dfrbp_1 _2505_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net271),
    .D(net54),
    .Q_N(_1250_),
    .Q(\sm_i.ssw_reg[1][0] ));
 sg13g2_dfrbp_1 _2506_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net269),
    .D(net52),
    .Q_N(_1251_),
    .Q(\sm_i.ssw_reg[1][1] ));
 sg13g2_dfrbp_1 _2507_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net269),
    .D(net47),
    .Q_N(_1252_),
    .Q(\sm_i.ssw_reg[1][2] ));
 sg13g2_dfrbp_1 _2508_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net270),
    .D(net45),
    .Q_N(_1253_),
    .Q(\sm_i.ssw_reg[1][3] ));
 sg13g2_dfrbp_1 _2509_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net273),
    .D(net40),
    .Q_N(_1254_),
    .Q(\sm_i.ssw_reg[1][4] ));
 sg13g2_dfrbp_1 _2510_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net273),
    .D(net48),
    .Q_N(_1255_),
    .Q(\sm_i.ssw_reg[1][5] ));
 sg13g2_dfrbp_1 _2511_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net270),
    .D(net39),
    .Q_N(_1256_),
    .Q(\sm_i.ssw_reg[1][6] ));
 sg13g2_dfrbp_1 _2512_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net271),
    .D(net38),
    .Q_N(_1161_),
    .Q(\sm_i.ssw_reg[1][7] ));
 sg13g2_dfrbp_1 _2513_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net275),
    .D(_0103_),
    .Q_N(\sm_i.snote_synch[2][0] ),
    .Q(_0100_));
 sg13g2_dfrbp_1 _2514_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net274),
    .D(net50),
    .Q_N(_1257_),
    .Q(\sm_i.snote_synch[2][1] ));
 sg13g2_dfrbp_1 _2515_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net275),
    .D(net56),
    .Q_N(_0086_),
    .Q(\sm_i.snote_synch[2][2] ));
 sg13g2_dfrbp_1 _2516_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net275),
    .D(net61),
    .Q_N(_0087_),
    .Q(\sm_i.snote_synch[2][3] ));
 sg13g2_dfrbp_1 _2517_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net275),
    .D(net60),
    .Q_N(_1160_),
    .Q(\sm_i.snote_synch[2][4] ));
 sg13g2_tielo tt_um_synth_simple_mm_15 (.L_LO(net15));
 sg13g2_tielo tt_um_synth_simple_mm_16 (.L_LO(net16));
 sg13g2_tielo tt_um_synth_simple_mm_17 (.L_LO(net17));
 sg13g2_tielo tt_um_synth_simple_mm_18 (.L_LO(net18));
 sg13g2_tielo tt_um_synth_simple_mm_19 (.L_LO(net19));
 sg13g2_tielo tt_um_synth_simple_mm_20 (.L_LO(net20));
 sg13g2_tielo tt_um_synth_simple_mm_21 (.L_LO(net21));
 sg13g2_tielo tt_um_synth_simple_mm_22 (.L_LO(net22));
 sg13g2_tielo tt_um_synth_simple_mm_23 (.L_LO(net23));
 sg13g2_tielo tt_um_synth_simple_mm_24 (.L_LO(net24));
 sg13g2_tielo tt_um_synth_simple_mm_25 (.L_LO(net25));
 sg13g2_tielo tt_um_synth_simple_mm_26 (.L_LO(net26));
 sg13g2_tielo tt_um_synth_simple_mm_27 (.L_LO(net27));
 sg13g2_tielo tt_um_synth_simple_mm_28 (.L_LO(net28));
 sg13g2_tielo tt_um_synth_simple_mm_29 (.L_LO(net29));
 sg13g2_tielo tt_um_synth_simple_mm_30 (.L_LO(net30));
 sg13g2_tielo tt_um_synth_simple_mm_31 (.L_LO(net31));
 sg13g2_tielo tt_um_synth_simple_mm_32 (.L_LO(net32));
 sg13g2_tielo tt_um_synth_simple_mm_33 (.L_LO(net33));
 sg13g2_tielo tt_um_synth_simple_mm_34 (.L_LO(net34));
 sg13g2_tielo tt_um_synth_simple_mm_35 (.L_LO(net35));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _2540_ (.A(pwm_out_i),
    .X(uo_out[0]));
 sg13g2_buf_1 _2541_ (.A(pwm_out_right),
    .X(uo_out[1]));
 sg13g2_buf_2 fanout211 (.A(_0703_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_0703_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(net214),
    .X(net213));
 sg13g2_buf_1 fanout214 (.A(_0702_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_0519_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(net219),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(net219),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(net219),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_0191_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_0188_),
    .X(net220));
 sg13g2_buf_1 fanout221 (.A(_0188_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(net223),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_0188_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_1058_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(net226),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(\sm_i.adsr_i.vout ),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_0896_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_0895_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_0820_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(net231),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_0820_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_0740_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_0363_),
    .X(net233));
 sg13g2_buf_4 fanout234 (.X(net234),
    .A(_0851_));
 sg13g2_buf_2 fanout235 (.A(_0851_),
    .X(net235));
 sg13g2_buf_4 fanout236 (.X(net236),
    .A(_0604_));
 sg13g2_buf_2 fanout237 (.A(_0604_),
    .X(net237));
 sg13g2_buf_4 fanout238 (.X(net238),
    .A(_0603_));
 sg13g2_buf_2 fanout239 (.A(_0572_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(net241),
    .X(net240));
 sg13g2_buf_1 fanout241 (.A(\sm_i.ssw_reg[2][0] ),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(net279),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_0041_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(net245),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(net126),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(net247),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(net287),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(net65),
    .X(net248));
 sg13g2_buf_4 fanout249 (.X(net249),
    .A(net250));
 sg13g2_buf_4 fanout250 (.X(net250),
    .A(net253));
 sg13g2_buf_4 fanout251 (.X(net251),
    .A(net252));
 sg13g2_buf_2 fanout252 (.A(net253),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(net260),
    .X(net253));
 sg13g2_buf_4 fanout254 (.X(net254),
    .A(net257));
 sg13g2_buf_4 fanout255 (.X(net255),
    .A(net256));
 sg13g2_buf_4 fanout256 (.X(net256),
    .A(net257));
 sg13g2_buf_2 fanout257 (.A(net260),
    .X(net257));
 sg13g2_buf_4 fanout258 (.X(net258),
    .A(net260));
 sg13g2_buf_2 fanout259 (.A(net260),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(rst_n),
    .X(net260));
 sg13g2_buf_4 fanout261 (.X(net261),
    .A(net264));
 sg13g2_buf_2 fanout262 (.A(net264),
    .X(net262));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(net264));
 sg13g2_buf_2 fanout264 (.A(net277),
    .X(net264));
 sg13g2_buf_4 fanout265 (.X(net265),
    .A(net268));
 sg13g2_buf_4 fanout266 (.X(net266),
    .A(net268));
 sg13g2_buf_2 fanout267 (.A(net268),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(net277),
    .X(net268));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(net272));
 sg13g2_buf_4 fanout270 (.X(net270),
    .A(net271));
 sg13g2_buf_2 fanout271 (.A(net272),
    .X(net271));
 sg13g2_buf_4 fanout272 (.X(net272),
    .A(net277));
 sg13g2_buf_4 fanout273 (.X(net273),
    .A(net277));
 sg13g2_buf_4 fanout274 (.X(net274),
    .A(net275));
 sg13g2_buf_4 fanout275 (.X(net275),
    .A(net276));
 sg13g2_buf_4 fanout276 (.X(net276),
    .A(net277));
 sg13g2_buf_2 fanout277 (.A(rst_n),
    .X(net277));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[0]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[1]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[2]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[3]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[4]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[5]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[6]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[7]),
    .X(net13));
 sg13g2_tielo tt_um_synth_simple_mm_14 (.L_LO(net14));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_17__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\sm_i.snote_synch[0][3] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold2 (.A(\sm_i.snote_synch[0][4] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold3 (.A(\sm_i.ssw_reg[0][7] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold4 (.A(\sm_i.ssw_reg[0][6] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold5 (.A(\sm_i.ssw_reg[0][4] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold6 (.A(\sm_i.ssw_reg[1][7] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold7 (.A(\sm_i.ssw_reg[1][5] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold8 (.A(\sm_i.ssw_reg[1][6] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold9 (.A(\sm_i.ssw_reg[1][1] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold10 (.A(\sm_i.ssw_reg[0][3] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold11 (.A(\sm_i.snote_synch[0][0] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold12 (.A(\sm_i.ssw_reg[0][2] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold13 (.A(\sm_i.ssw_reg[0][5] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold14 (.A(\sm_i.ssw_reg[1][4] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold15 (.A(\sm_i.snote_synch[1][1] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold16 (.A(\sm_i.ssw_reg[1][3] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold17 (.A(\sm_i.ssw_reg[0][1] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold18 (.A(\sm_i.snote_synch[0][1] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold19 (.A(\sm_i.ssw_reg[0][0] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold20 (.A(pwm_out_i),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold21 (.A(\sm_i.snote_synch[1][2] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold22 (.A(\sm_i.ssw_reg[1][0] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold23 (.A(\sm_i.snote_synch[1][0] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold24 (.A(\sm_i.snote_synch[0][2] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold25 (.A(\sm_i.snote_synch[1][4] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold26 (.A(\sm_i.snote_synch[1][3] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold27 (.A(\sm_i.ssw_reg[1][2] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0044_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0167_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold30 (.A(\sm_i.wav_gen_1.snote_enable ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold31 (.A(\sm_i.wav_gen_1.rom_ampl_sin_i.en ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold32 (.A(\sm_i.wav_gen_1.swave_squ_sel ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold33 (.A(\sm_i.scnt_pwm[0] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0089_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0093_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0096_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold37 (.A(\sm_i.scnt_pwm[6] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0809_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0006_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0095_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0094_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0090_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0092_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold44 (.A(\sm_i.adsr_i.scnt_step[2] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0141_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold46 (.A(\sm_i.scnt_pwm[4] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0004_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0088_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0091_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold50 (.A(\sm_i.scnt_pwm_on[7] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0510_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0174_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold53 (.A(\sm_i.scnt_pwm[3] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0003_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold55 (.A(\sm_i.adsr_i.scnt_step[8] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0147_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold57 (.A(\sm_i.adsr_i.scnt_step[4] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0143_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold59 (.A(\sm_i.adsr_i.scnt_step[3] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0142_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0097_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold62 (.A(\sm_i.adsr_i.scnt_step[9] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0148_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold64 (.A(\sm_i.scnt_pwm[1] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold65 (.A(\sm_i.adsr_i.scnt_step[5] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0144_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold67 (.A(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[12] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold68 (.A(\sm_i.adsr_i.scnt_step[12] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0151_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold70 (.A(\sm_i.adsr_i.scnt_step[26] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0272_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0165_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold73 (.A(\sm_i.adsr_i.scnt_step[13] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0152_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold75 (.A(\sm_i.adsr_i.scnt_step[15] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0154_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold77 (.A(\sm_i.scnt_pwm[5] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold78 (.A(\sm_i.wav_gen_1.sstep_cnt[0] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold79 (.A(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[0] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold80 (.A(\sm_i.adsr_i.scnt_step[6] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0145_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold82 (.A(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[10] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold83 (.A(\sm_i.adsr_i.scnt_step[7] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0146_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold85 (.A(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[5] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold86 (.A(\sm_i.adsr_i.scnt_step[14] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0153_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold88 (.A(\sm_i.wav_gen_1.swave_cnt_tri[3] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold89 (.A(\sm_i.scnt_pwm[7] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold90 (.A(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[11] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold91 (.A(\sm_i.wav_gen_1.swave_cnt_tri[5] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold92 (.A(\sm_i.adsr_i.scnt_step[10] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0082_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0729_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0083_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0829_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0104_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold98 (.A(\sm_i.adsr_i.scnt_step[11] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0150_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0075_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0711_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold102 (.A(\sm_i.wav_gen_1.sstep_cnt[3] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0707_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0017_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold105 (.A(\sm_i.adsr_i.scnt_step[24] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0269_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold107 (.A(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[1] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold108 (.A(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[0] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold109 (.A(\sm_i.adsr_i.scnt_step[20] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0159_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0081_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0727_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold113 (.A(\sm_i.wav_gen_1.sstep_cnt[1] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0079_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0720_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold116 (.A(\sm_i.adsr_i.scnt_step[27] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0275_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold118 (.A(\sm_i.scnt_pwm_on[4] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0171_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold120 (.A(\sm_i.scnt_pwm_on[3] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0419_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0170_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold123 (.A(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[5] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold124 (.A(\sm_i.wav_gen_1.sstep_cnt[7] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0714_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0021_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold127 (.A(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[4] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold128 (.A(\sm_i.adsr_i.dout[1] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0176_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold130 (.A(\sm_i.adsr_i.scnt_step[17] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0156_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold132 (.A(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[6] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold133 (.A(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[3] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold134 (.A(\sm_i.wav_gen_1.swave_cnt_tri[4] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0076_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0713_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold137 (.A(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[1] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold138 (.A(\sm_i.wav_gen_1.rom_freq_tri_squ_sin_i.data_out[6] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold139 (.A(\sm_i.scnt_pwm_on[5] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold140 (.A(\sm_i.wav_gen_1.rom_freq_saw_i.data_out[7] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0062_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold142 (.A(_1127_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0073_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0078_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0718_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold146 (.A(\sm_i.wav_gen_1.sstep_cnt[15] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0731_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold148 (.A(\sm_i.adsr_i.scnt_step[23] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0162_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold150 (.A(\sm_i.scnt_pwm_on[0] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0385_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0168_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold153 (.A(\sm_i.adsr_i.scnt_step[25] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0271_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold155 (.A(\sm_i.adsr_i.scnt_step[22] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0074_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0710_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold158 (.A(\sm_i.adsr_i.scnt_step[19] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold159 (.A(\sm_i.adsr_i.scnt_step[21] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0160_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold161 (.A(\sm_i.adsr_i.scnt_step[0] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold162 (.A(\sm_i.adsr_i.sstate[2] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0108_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold164 (.A(\sm_i.adsr_i.scnt_step[16] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0155_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold166 (.A(\sm_i.adsr_i.scnt_step[18] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold167 (.A(\sm_i.wav_gen_1.swave_cnt_tri[2] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold168 (.A(\sm_i.adsr_i.scnt_step[1] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold169 (.A(\sm_i.scnt_pwm_on[6] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold170 (.A(\sm_i.adsr_i.dout[3] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0080_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0725_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0011_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold174 (.A(\sm_i.adsr_i.dout[4] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0077_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0716_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold177 (.A(\sm_i.adsr_i.scnt_pwl[0] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold178 (.A(\sm_i.adsr_i.scnt_pwl[1] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold179 (.A(\sm_i.scnt_pwm[2] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold180 (.A(\sm_i.wav_gen_1.swave_cnt_tri[1] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0121_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold182 (.A(\sm_i.adsr_i.dout[2] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold183 (.A(\sm_i.adsr_i.sstate[0] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0106_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold185 (.A(\sm_i.wav_gen_1.swave_cnt_tri_down_up_n ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0105_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold187 (.A(\sm_i.adsr_i.sstate[1] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0107_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0063_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold190 (.A(\sm_i.scnt_pwm_on[2] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0386_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold192 (.A(\sm_i.wav_gen_1.sstep_cnt[8] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0722_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0723_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0010_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold196 (.A(\sm_i.scnt_pwm_on[2] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold197 (.A(\sm_i.adsr_i.scnt_pwl[2] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0183_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold199 (.A(\sm_i.adsr_i.dout[5] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0060_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold201 (.A(_1143_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold202 (.A(\sm_i.adsr_i.dout[0] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold203 (.A(\sm_i.wav_gen_1.rom_ampl_sin_i.addr[0] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0065_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold205 (.A(\sm_i.adsr_i.scnt_step[22] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0268_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold207 (.A(\sm_i.adsr_i.scnt_step[18] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold208 (.A(\sm_i.adsr_i.scnt_step[21] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold209 (.A(\sm_i.adsr_i.dout[0] ),
    .X(net311));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_4 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_131 ();
 sg13g2_decap_8 FILLER_0_138 ();
 sg13g2_decap_8 FILLER_0_145 ();
 sg13g2_decap_8 FILLER_0_152 ();
 sg13g2_decap_8 FILLER_0_159 ();
 sg13g2_decap_8 FILLER_0_166 ();
 sg13g2_decap_8 FILLER_0_173 ();
 sg13g2_decap_8 FILLER_0_180 ();
 sg13g2_decap_8 FILLER_0_187 ();
 sg13g2_decap_8 FILLER_0_194 ();
 sg13g2_decap_8 FILLER_0_201 ();
 sg13g2_decap_8 FILLER_0_208 ();
 sg13g2_decap_8 FILLER_0_215 ();
 sg13g2_decap_8 FILLER_0_222 ();
 sg13g2_decap_8 FILLER_0_229 ();
 sg13g2_decap_8 FILLER_0_236 ();
 sg13g2_decap_8 FILLER_0_243 ();
 sg13g2_decap_8 FILLER_0_250 ();
 sg13g2_decap_8 FILLER_0_257 ();
 sg13g2_decap_8 FILLER_0_264 ();
 sg13g2_decap_8 FILLER_0_271 ();
 sg13g2_decap_8 FILLER_0_278 ();
 sg13g2_decap_8 FILLER_0_285 ();
 sg13g2_decap_8 FILLER_0_292 ();
 sg13g2_decap_8 FILLER_0_299 ();
 sg13g2_decap_8 FILLER_0_306 ();
 sg13g2_decap_4 FILLER_0_313 ();
 sg13g2_fill_1 FILLER_0_347 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_4 FILLER_1_35 ();
 sg13g2_fill_1 FILLER_1_39 ();
 sg13g2_decap_8 FILLER_1_44 ();
 sg13g2_decap_8 FILLER_1_51 ();
 sg13g2_fill_2 FILLER_1_58 ();
 sg13g2_fill_1 FILLER_1_60 ();
 sg13g2_fill_2 FILLER_1_71 ();
 sg13g2_fill_1 FILLER_1_73 ();
 sg13g2_decap_8 FILLER_1_79 ();
 sg13g2_decap_8 FILLER_1_86 ();
 sg13g2_decap_8 FILLER_1_93 ();
 sg13g2_decap_8 FILLER_1_100 ();
 sg13g2_fill_2 FILLER_1_107 ();
 sg13g2_fill_1 FILLER_1_121 ();
 sg13g2_decap_8 FILLER_1_139 ();
 sg13g2_decap_8 FILLER_1_146 ();
 sg13g2_decap_8 FILLER_1_153 ();
 sg13g2_fill_2 FILLER_1_160 ();
 sg13g2_fill_2 FILLER_1_166 ();
 sg13g2_decap_8 FILLER_1_171 ();
 sg13g2_decap_8 FILLER_1_178 ();
 sg13g2_decap_8 FILLER_1_185 ();
 sg13g2_decap_8 FILLER_1_192 ();
 sg13g2_decap_8 FILLER_1_199 ();
 sg13g2_decap_8 FILLER_1_206 ();
 sg13g2_decap_8 FILLER_1_213 ();
 sg13g2_decap_8 FILLER_1_220 ();
 sg13g2_decap_8 FILLER_1_227 ();
 sg13g2_decap_8 FILLER_1_234 ();
 sg13g2_decap_8 FILLER_1_241 ();
 sg13g2_decap_8 FILLER_1_248 ();
 sg13g2_decap_8 FILLER_1_255 ();
 sg13g2_decap_8 FILLER_1_262 ();
 sg13g2_decap_8 FILLER_1_269 ();
 sg13g2_decap_8 FILLER_1_276 ();
 sg13g2_decap_8 FILLER_1_283 ();
 sg13g2_fill_1 FILLER_1_290 ();
 sg13g2_decap_8 FILLER_1_295 ();
 sg13g2_fill_1 FILLER_1_307 ();
 sg13g2_fill_1 FILLER_1_317 ();
 sg13g2_decap_4 FILLER_1_405 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_4 FILLER_2_21 ();
 sg13g2_fill_1 FILLER_2_25 ();
 sg13g2_fill_1 FILLER_2_49 ();
 sg13g2_fill_2 FILLER_2_63 ();
 sg13g2_fill_1 FILLER_2_65 ();
 sg13g2_fill_2 FILLER_2_74 ();
 sg13g2_fill_1 FILLER_2_76 ();
 sg13g2_fill_2 FILLER_2_94 ();
 sg13g2_fill_2 FILLER_2_147 ();
 sg13g2_fill_2 FILLER_2_162 ();
 sg13g2_decap_4 FILLER_2_198 ();
 sg13g2_fill_1 FILLER_2_202 ();
 sg13g2_decap_8 FILLER_2_212 ();
 sg13g2_decap_8 FILLER_2_219 ();
 sg13g2_decap_4 FILLER_2_226 ();
 sg13g2_fill_2 FILLER_2_263 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_fill_2 FILLER_3_101 ();
 sg13g2_fill_2 FILLER_3_126 ();
 sg13g2_fill_1 FILLER_3_159 ();
 sg13g2_fill_1 FILLER_3_174 ();
 sg13g2_decap_8 FILLER_3_215 ();
 sg13g2_fill_2 FILLER_3_222 ();
 sg13g2_fill_1 FILLER_3_224 ();
 sg13g2_fill_2 FILLER_3_239 ();
 sg13g2_fill_1 FILLER_3_241 ();
 sg13g2_fill_1 FILLER_3_321 ();
 sg13g2_fill_1 FILLER_3_377 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_fill_2 FILLER_4_28 ();
 sg13g2_fill_1 FILLER_4_30 ();
 sg13g2_fill_2 FILLER_4_84 ();
 sg13g2_fill_1 FILLER_4_86 ();
 sg13g2_fill_1 FILLER_4_167 ();
 sg13g2_fill_1 FILLER_4_220 ();
 sg13g2_fill_2 FILLER_4_266 ();
 sg13g2_fill_2 FILLER_4_283 ();
 sg13g2_fill_1 FILLER_4_325 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_4 FILLER_5_21 ();
 sg13g2_fill_1 FILLER_5_25 ();
 sg13g2_fill_1 FILLER_5_40 ();
 sg13g2_fill_2 FILLER_5_110 ();
 sg13g2_fill_1 FILLER_5_124 ();
 sg13g2_fill_2 FILLER_5_160 ();
 sg13g2_fill_2 FILLER_5_187 ();
 sg13g2_fill_1 FILLER_5_221 ();
 sg13g2_fill_1 FILLER_5_231 ();
 sg13g2_fill_1 FILLER_5_246 ();
 sg13g2_fill_1 FILLER_5_256 ();
 sg13g2_fill_2 FILLER_5_338 ();
 sg13g2_fill_1 FILLER_5_340 ();
 sg13g2_fill_1 FILLER_5_365 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_fill_1 FILLER_6_14 ();
 sg13g2_fill_2 FILLER_6_95 ();
 sg13g2_fill_1 FILLER_6_127 ();
 sg13g2_fill_2 FILLER_6_215 ();
 sg13g2_fill_1 FILLER_6_247 ();
 sg13g2_fill_1 FILLER_6_266 ();
 sg13g2_fill_1 FILLER_6_345 ();
 sg13g2_decap_8 FILLER_6_382 ();
 sg13g2_fill_2 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_4 FILLER_7_14 ();
 sg13g2_fill_2 FILLER_7_18 ();
 sg13g2_fill_2 FILLER_7_46 ();
 sg13g2_fill_1 FILLER_7_48 ();
 sg13g2_fill_2 FILLER_7_109 ();
 sg13g2_fill_1 FILLER_7_111 ();
 sg13g2_fill_1 FILLER_7_147 ();
 sg13g2_fill_2 FILLER_7_241 ();
 sg13g2_fill_2 FILLER_7_255 ();
 sg13g2_fill_1 FILLER_7_277 ();
 sg13g2_decap_8 FILLER_7_296 ();
 sg13g2_decap_8 FILLER_7_303 ();
 sg13g2_decap_4 FILLER_7_310 ();
 sg13g2_decap_4 FILLER_7_319 ();
 sg13g2_fill_2 FILLER_7_337 ();
 sg13g2_fill_1 FILLER_7_339 ();
 sg13g2_fill_1 FILLER_7_344 ();
 sg13g2_decap_8 FILLER_7_353 ();
 sg13g2_fill_1 FILLER_7_360 ();
 sg13g2_fill_2 FILLER_7_366 ();
 sg13g2_fill_2 FILLER_7_389 ();
 sg13g2_decap_4 FILLER_7_405 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_4 FILLER_8_7 ();
 sg13g2_fill_1 FILLER_8_11 ();
 sg13g2_fill_1 FILLER_8_38 ();
 sg13g2_fill_2 FILLER_8_48 ();
 sg13g2_fill_1 FILLER_8_64 ();
 sg13g2_fill_2 FILLER_8_78 ();
 sg13g2_fill_1 FILLER_8_80 ();
 sg13g2_fill_1 FILLER_8_100 ();
 sg13g2_fill_1 FILLER_8_132 ();
 sg13g2_fill_2 FILLER_8_167 ();
 sg13g2_fill_2 FILLER_8_273 ();
 sg13g2_fill_1 FILLER_8_275 ();
 sg13g2_decap_4 FILLER_8_297 ();
 sg13g2_fill_1 FILLER_8_313 ();
 sg13g2_decap_4 FILLER_8_357 ();
 sg13g2_fill_2 FILLER_8_361 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_fill_2 FILLER_9_28 ();
 sg13g2_fill_2 FILLER_9_86 ();
 sg13g2_fill_1 FILLER_9_88 ();
 sg13g2_decap_4 FILLER_9_105 ();
 sg13g2_decap_4 FILLER_9_114 ();
 sg13g2_decap_4 FILLER_9_127 ();
 sg13g2_fill_1 FILLER_9_141 ();
 sg13g2_fill_1 FILLER_9_178 ();
 sg13g2_fill_2 FILLER_9_220 ();
 sg13g2_fill_2 FILLER_9_261 ();
 sg13g2_decap_4 FILLER_9_287 ();
 sg13g2_fill_2 FILLER_9_303 ();
 sg13g2_fill_1 FILLER_9_305 ();
 sg13g2_fill_2 FILLER_9_315 ();
 sg13g2_fill_1 FILLER_9_317 ();
 sg13g2_decap_4 FILLER_9_323 ();
 sg13g2_fill_1 FILLER_9_327 ();
 sg13g2_decap_8 FILLER_9_361 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_4 FILLER_10_14 ();
 sg13g2_fill_2 FILLER_10_18 ();
 sg13g2_fill_2 FILLER_10_46 ();
 sg13g2_fill_1 FILLER_10_48 ();
 sg13g2_decap_4 FILLER_10_80 ();
 sg13g2_fill_1 FILLER_10_84 ();
 sg13g2_fill_1 FILLER_10_93 ();
 sg13g2_decap_8 FILLER_10_100 ();
 sg13g2_fill_1 FILLER_10_107 ();
 sg13g2_fill_1 FILLER_10_124 ();
 sg13g2_fill_1 FILLER_10_135 ();
 sg13g2_fill_1 FILLER_10_174 ();
 sg13g2_decap_4 FILLER_10_291 ();
 sg13g2_fill_1 FILLER_10_295 ();
 sg13g2_fill_1 FILLER_10_311 ();
 sg13g2_fill_1 FILLER_10_347 ();
 sg13g2_fill_2 FILLER_10_374 ();
 sg13g2_fill_1 FILLER_10_376 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_4 FILLER_11_21 ();
 sg13g2_fill_2 FILLER_11_25 ();
 sg13g2_fill_2 FILLER_11_52 ();
 sg13g2_fill_1 FILLER_11_54 ();
 sg13g2_fill_1 FILLER_11_77 ();
 sg13g2_fill_1 FILLER_11_88 ();
 sg13g2_decap_4 FILLER_11_99 ();
 sg13g2_fill_2 FILLER_11_117 ();
 sg13g2_fill_1 FILLER_11_119 ();
 sg13g2_fill_2 FILLER_11_130 ();
 sg13g2_fill_1 FILLER_11_146 ();
 sg13g2_decap_8 FILLER_11_236 ();
 sg13g2_fill_1 FILLER_11_243 ();
 sg13g2_decap_8 FILLER_11_269 ();
 sg13g2_fill_1 FILLER_11_276 ();
 sg13g2_fill_2 FILLER_11_281 ();
 sg13g2_fill_1 FILLER_11_283 ();
 sg13g2_fill_2 FILLER_11_310 ();
 sg13g2_decap_8 FILLER_11_324 ();
 sg13g2_fill_2 FILLER_11_331 ();
 sg13g2_fill_2 FILLER_11_360 ();
 sg13g2_fill_1 FILLER_11_387 ();
 sg13g2_decap_4 FILLER_11_405 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_7 ();
 sg13g2_fill_1 FILLER_12_9 ();
 sg13g2_fill_1 FILLER_12_41 ();
 sg13g2_fill_2 FILLER_12_95 ();
 sg13g2_fill_2 FILLER_12_111 ();
 sg13g2_fill_1 FILLER_12_117 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_fill_2 FILLER_12_133 ();
 sg13g2_fill_1 FILLER_12_152 ();
 sg13g2_fill_2 FILLER_12_162 ();
 sg13g2_fill_1 FILLER_12_171 ();
 sg13g2_fill_2 FILLER_12_231 ();
 sg13g2_fill_1 FILLER_12_233 ();
 sg13g2_decap_8 FILLER_12_260 ();
 sg13g2_decap_8 FILLER_12_267 ();
 sg13g2_fill_2 FILLER_12_274 ();
 sg13g2_fill_2 FILLER_12_315 ();
 sg13g2_fill_2 FILLER_12_348 ();
 sg13g2_fill_1 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_fill_1 FILLER_13_21 ();
 sg13g2_fill_2 FILLER_13_40 ();
 sg13g2_fill_2 FILLER_13_51 ();
 sg13g2_fill_2 FILLER_13_65 ();
 sg13g2_decap_4 FILLER_13_87 ();
 sg13g2_fill_1 FILLER_13_103 ();
 sg13g2_fill_1 FILLER_13_113 ();
 sg13g2_fill_2 FILLER_13_163 ();
 sg13g2_fill_2 FILLER_13_171 ();
 sg13g2_decap_4 FILLER_13_177 ();
 sg13g2_fill_2 FILLER_13_340 ();
 sg13g2_fill_1 FILLER_13_342 ();
 sg13g2_fill_1 FILLER_13_372 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_fill_1 FILLER_14_21 ();
 sg13g2_decap_4 FILLER_14_83 ();
 sg13g2_fill_1 FILLER_14_87 ();
 sg13g2_fill_2 FILLER_14_101 ();
 sg13g2_decap_4 FILLER_14_108 ();
 sg13g2_fill_1 FILLER_14_116 ();
 sg13g2_decap_4 FILLER_14_131 ();
 sg13g2_fill_1 FILLER_14_135 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_fill_2 FILLER_14_215 ();
 sg13g2_fill_2 FILLER_14_247 ();
 sg13g2_fill_1 FILLER_14_249 ();
 sg13g2_decap_4 FILLER_14_260 ();
 sg13g2_fill_2 FILLER_14_313 ();
 sg13g2_fill_1 FILLER_14_315 ();
 sg13g2_fill_1 FILLER_14_326 ();
 sg13g2_fill_2 FILLER_14_341 ();
 sg13g2_fill_1 FILLER_14_343 ();
 sg13g2_fill_2 FILLER_14_350 ();
 sg13g2_fill_1 FILLER_14_352 ();
 sg13g2_fill_2 FILLER_14_365 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_4 FILLER_15_35 ();
 sg13g2_fill_1 FILLER_15_39 ();
 sg13g2_decap_8 FILLER_15_44 ();
 sg13g2_decap_8 FILLER_15_69 ();
 sg13g2_decap_8 FILLER_15_76 ();
 sg13g2_decap_4 FILLER_15_83 ();
 sg13g2_fill_1 FILLER_15_87 ();
 sg13g2_fill_2 FILLER_15_93 ();
 sg13g2_fill_1 FILLER_15_95 ();
 sg13g2_fill_2 FILLER_15_112 ();
 sg13g2_fill_1 FILLER_15_157 ();
 sg13g2_fill_2 FILLER_15_231 ();
 sg13g2_fill_1 FILLER_15_370 ();
 sg13g2_fill_1 FILLER_15_376 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_4 FILLER_16_21 ();
 sg13g2_fill_2 FILLER_16_25 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_fill_1 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_65 ();
 sg13g2_decap_8 FILLER_16_72 ();
 sg13g2_decap_8 FILLER_16_79 ();
 sg13g2_decap_4 FILLER_16_86 ();
 sg13g2_fill_2 FILLER_16_90 ();
 sg13g2_fill_2 FILLER_16_100 ();
 sg13g2_fill_1 FILLER_16_102 ();
 sg13g2_fill_2 FILLER_16_132 ();
 sg13g2_fill_2 FILLER_16_180 ();
 sg13g2_fill_2 FILLER_16_223 ();
 sg13g2_decap_8 FILLER_16_263 ();
 sg13g2_fill_2 FILLER_16_270 ();
 sg13g2_fill_1 FILLER_16_303 ();
 sg13g2_fill_1 FILLER_16_309 ();
 sg13g2_fill_1 FILLER_16_315 ();
 sg13g2_fill_2 FILLER_16_365 ();
 sg13g2_fill_1 FILLER_16_367 ();
 sg13g2_fill_1 FILLER_16_374 ();
 sg13g2_decap_4 FILLER_16_387 ();
 sg13g2_fill_2 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_fill_2 FILLER_17_105 ();
 sg13g2_fill_1 FILLER_17_107 ();
 sg13g2_fill_2 FILLER_17_121 ();
 sg13g2_fill_1 FILLER_17_123 ();
 sg13g2_fill_2 FILLER_17_164 ();
 sg13g2_fill_1 FILLER_17_207 ();
 sg13g2_fill_2 FILLER_17_291 ();
 sg13g2_fill_1 FILLER_17_293 ();
 sg13g2_fill_1 FILLER_17_306 ();
 sg13g2_fill_1 FILLER_17_342 ();
 sg13g2_fill_1 FILLER_17_359 ();
 sg13g2_fill_2 FILLER_17_375 ();
 sg13g2_fill_1 FILLER_17_377 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_4 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_78 ();
 sg13g2_decap_4 FILLER_18_85 ();
 sg13g2_fill_1 FILLER_18_89 ();
 sg13g2_decap_8 FILLER_18_95 ();
 sg13g2_decap_8 FILLER_18_102 ();
 sg13g2_fill_2 FILLER_18_109 ();
 sg13g2_decap_8 FILLER_18_115 ();
 sg13g2_decap_8 FILLER_18_122 ();
 sg13g2_decap_8 FILLER_18_129 ();
 sg13g2_decap_4 FILLER_18_136 ();
 sg13g2_fill_2 FILLER_18_140 ();
 sg13g2_fill_1 FILLER_18_155 ();
 sg13g2_fill_1 FILLER_18_165 ();
 sg13g2_fill_1 FILLER_18_192 ();
 sg13g2_fill_1 FILLER_18_219 ();
 sg13g2_decap_4 FILLER_18_249 ();
 sg13g2_fill_1 FILLER_18_253 ();
 sg13g2_decap_8 FILLER_18_257 ();
 sg13g2_decap_4 FILLER_18_264 ();
 sg13g2_fill_1 FILLER_18_294 ();
 sg13g2_fill_2 FILLER_18_312 ();
 sg13g2_fill_1 FILLER_18_314 ();
 sg13g2_decap_8 FILLER_18_325 ();
 sg13g2_decap_4 FILLER_18_332 ();
 sg13g2_fill_2 FILLER_18_360 ();
 sg13g2_fill_1 FILLER_18_380 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_4 ();
 sg13g2_fill_1 FILLER_19_89 ();
 sg13g2_fill_1 FILLER_19_95 ();
 sg13g2_decap_8 FILLER_19_122 ();
 sg13g2_fill_2 FILLER_19_129 ();
 sg13g2_fill_1 FILLER_19_131 ();
 sg13g2_fill_2 FILLER_19_157 ();
 sg13g2_fill_1 FILLER_19_159 ();
 sg13g2_fill_2 FILLER_19_190 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_fill_1 FILLER_19_215 ();
 sg13g2_fill_2 FILLER_19_226 ();
 sg13g2_fill_2 FILLER_19_236 ();
 sg13g2_fill_1 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_265 ();
 sg13g2_decap_8 FILLER_19_272 ();
 sg13g2_fill_2 FILLER_19_279 ();
 sg13g2_fill_2 FILLER_19_289 ();
 sg13g2_fill_1 FILLER_19_291 ();
 sg13g2_fill_2 FILLER_19_340 ();
 sg13g2_fill_2 FILLER_19_347 ();
 sg13g2_fill_1 FILLER_19_349 ();
 sg13g2_fill_1 FILLER_19_368 ();
 sg13g2_fill_1 FILLER_19_396 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_67 ();
 sg13g2_fill_2 FILLER_20_100 ();
 sg13g2_fill_1 FILLER_20_102 ();
 sg13g2_decap_4 FILLER_20_129 ();
 sg13g2_fill_1 FILLER_20_163 ();
 sg13g2_fill_1 FILLER_20_189 ();
 sg13g2_fill_2 FILLER_20_221 ();
 sg13g2_fill_1 FILLER_20_223 ();
 sg13g2_decap_8 FILLER_20_237 ();
 sg13g2_decap_8 FILLER_20_244 ();
 sg13g2_fill_2 FILLER_20_251 ();
 sg13g2_decap_8 FILLER_20_305 ();
 sg13g2_fill_1 FILLER_20_312 ();
 sg13g2_decap_8 FILLER_20_370 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_4 ();
 sg13g2_decap_4 FILLER_21_14 ();
 sg13g2_fill_2 FILLER_21_50 ();
 sg13g2_fill_1 FILLER_21_61 ();
 sg13g2_fill_1 FILLER_21_79 ();
 sg13g2_fill_1 FILLER_21_92 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_4 FILLER_21_154 ();
 sg13g2_fill_2 FILLER_21_158 ();
 sg13g2_fill_2 FILLER_21_168 ();
 sg13g2_fill_1 FILLER_21_170 ();
 sg13g2_decap_8 FILLER_21_177 ();
 sg13g2_decap_4 FILLER_21_184 ();
 sg13g2_fill_2 FILLER_21_188 ();
 sg13g2_decap_8 FILLER_21_193 ();
 sg13g2_fill_1 FILLER_21_200 ();
 sg13g2_fill_1 FILLER_21_205 ();
 sg13g2_fill_2 FILLER_21_213 ();
 sg13g2_fill_1 FILLER_21_215 ();
 sg13g2_decap_8 FILLER_21_269 ();
 sg13g2_decap_8 FILLER_21_276 ();
 sg13g2_decap_8 FILLER_21_283 ();
 sg13g2_fill_1 FILLER_21_290 ();
 sg13g2_fill_2 FILLER_21_325 ();
 sg13g2_decap_4 FILLER_21_335 ();
 sg13g2_decap_8 FILLER_21_360 ();
 sg13g2_fill_2 FILLER_21_367 ();
 sg13g2_decap_4 FILLER_21_374 ();
 sg13g2_fill_1 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_384 ();
 sg13g2_fill_2 FILLER_21_391 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_15 ();
 sg13g2_fill_2 FILLER_22_22 ();
 sg13g2_fill_2 FILLER_22_38 ();
 sg13g2_fill_2 FILLER_22_58 ();
 sg13g2_decap_8 FILLER_22_135 ();
 sg13g2_decap_8 FILLER_22_142 ();
 sg13g2_decap_8 FILLER_22_149 ();
 sg13g2_fill_1 FILLER_22_156 ();
 sg13g2_fill_2 FILLER_22_182 ();
 sg13g2_fill_2 FILLER_22_198 ();
 sg13g2_fill_1 FILLER_22_255 ();
 sg13g2_decap_8 FILLER_22_282 ();
 sg13g2_fill_2 FILLER_22_289 ();
 sg13g2_fill_2 FILLER_22_343 ();
 sg13g2_fill_2 FILLER_22_380 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_fill_2 FILLER_22_389 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_2 ();
 sg13g2_fill_1 FILLER_23_16 ();
 sg13g2_fill_2 FILLER_23_45 ();
 sg13g2_decap_4 FILLER_23_52 ();
 sg13g2_fill_2 FILLER_23_72 ();
 sg13g2_fill_2 FILLER_23_83 ();
 sg13g2_fill_1 FILLER_23_85 ();
 sg13g2_fill_1 FILLER_23_93 ();
 sg13g2_fill_2 FILLER_23_122 ();
 sg13g2_fill_1 FILLER_23_154 ();
 sg13g2_fill_1 FILLER_23_170 ();
 sg13g2_fill_2 FILLER_23_185 ();
 sg13g2_fill_1 FILLER_23_187 ();
 sg13g2_fill_1 FILLER_23_206 ();
 sg13g2_fill_2 FILLER_23_221 ();
 sg13g2_fill_1 FILLER_23_235 ();
 sg13g2_fill_2 FILLER_23_272 ();
 sg13g2_decap_4 FILLER_23_310 ();
 sg13g2_fill_1 FILLER_23_314 ();
 sg13g2_fill_1 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_338 ();
 sg13g2_fill_2 FILLER_23_345 ();
 sg13g2_fill_1 FILLER_23_361 ();
 sg13g2_fill_1 FILLER_23_366 ();
 sg13g2_fill_2 FILLER_23_381 ();
 sg13g2_fill_1 FILLER_23_383 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_2 ();
 sg13g2_fill_1 FILLER_24_23 ();
 sg13g2_fill_2 FILLER_24_29 ();
 sg13g2_fill_2 FILLER_24_54 ();
 sg13g2_fill_1 FILLER_24_56 ();
 sg13g2_fill_2 FILLER_24_96 ();
 sg13g2_fill_1 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_134 ();
 sg13g2_decap_4 FILLER_24_153 ();
 sg13g2_fill_2 FILLER_24_186 ();
 sg13g2_fill_1 FILLER_24_219 ();
 sg13g2_fill_2 FILLER_24_231 ();
 sg13g2_fill_2 FILLER_24_247 ();
 sg13g2_decap_8 FILLER_24_275 ();
 sg13g2_fill_1 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_335 ();
 sg13g2_decap_4 FILLER_24_342 ();
 sg13g2_fill_2 FILLER_24_354 ();
 sg13g2_fill_1 FILLER_24_356 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_fill_1 FILLER_25_18 ();
 sg13g2_fill_1 FILLER_25_33 ();
 sg13g2_fill_1 FILLER_25_81 ();
 sg13g2_fill_2 FILLER_25_87 ();
 sg13g2_fill_1 FILLER_25_98 ();
 sg13g2_fill_1 FILLER_25_116 ();
 sg13g2_decap_4 FILLER_25_153 ();
 sg13g2_fill_1 FILLER_25_157 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_4 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_4 FILLER_25_203 ();
 sg13g2_decap_4 FILLER_25_259 ();
 sg13g2_fill_2 FILLER_25_298 ();
 sg13g2_fill_2 FILLER_25_324 ();
 sg13g2_fill_2 FILLER_25_344 ();
 sg13g2_fill_1 FILLER_25_353 ();
 sg13g2_fill_1 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_25_375 ();
 sg13g2_fill_1 FILLER_25_382 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_28 ();
 sg13g2_fill_1 FILLER_26_30 ();
 sg13g2_fill_2 FILLER_26_79 ();
 sg13g2_decap_8 FILLER_26_125 ();
 sg13g2_fill_2 FILLER_26_132 ();
 sg13g2_fill_1 FILLER_26_134 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_4 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_198 ();
 sg13g2_fill_2 FILLER_26_205 ();
 sg13g2_fill_1 FILLER_26_212 ();
 sg13g2_fill_2 FILLER_26_237 ();
 sg13g2_fill_1 FILLER_26_256 ();
 sg13g2_fill_2 FILLER_26_271 ();
 sg13g2_fill_1 FILLER_26_273 ();
 sg13g2_fill_2 FILLER_26_380 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_4 ();
 sg13g2_fill_2 FILLER_27_37 ();
 sg13g2_fill_1 FILLER_27_39 ();
 sg13g2_fill_2 FILLER_27_52 ();
 sg13g2_fill_2 FILLER_27_116 ();
 sg13g2_fill_1 FILLER_27_118 ();
 sg13g2_fill_2 FILLER_27_145 ();
 sg13g2_fill_1 FILLER_27_155 ();
 sg13g2_fill_2 FILLER_27_166 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_fill_2 FILLER_27_182 ();
 sg13g2_fill_1 FILLER_27_184 ();
 sg13g2_decap_8 FILLER_27_209 ();
 sg13g2_decap_4 FILLER_27_233 ();
 sg13g2_fill_2 FILLER_27_237 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_fill_1 FILLER_27_245 ();
 sg13g2_fill_2 FILLER_27_264 ();
 sg13g2_fill_1 FILLER_27_266 ();
 sg13g2_fill_2 FILLER_27_272 ();
 sg13g2_fill_2 FILLER_27_361 ();
 sg13g2_fill_2 FILLER_27_368 ();
 sg13g2_decap_4 FILLER_27_380 ();
 sg13g2_fill_1 FILLER_27_388 ();
 sg13g2_fill_1 FILLER_27_393 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_4 ();
 sg13g2_fill_2 FILLER_28_36 ();
 sg13g2_fill_1 FILLER_28_38 ();
 sg13g2_fill_2 FILLER_28_48 ();
 sg13g2_decap_4 FILLER_28_55 ();
 sg13g2_fill_1 FILLER_28_59 ();
 sg13g2_decap_8 FILLER_28_68 ();
 sg13g2_fill_1 FILLER_28_75 ();
 sg13g2_fill_2 FILLER_28_84 ();
 sg13g2_fill_2 FILLER_28_112 ();
 sg13g2_fill_2 FILLER_28_123 ();
 sg13g2_fill_1 FILLER_28_125 ();
 sg13g2_decap_8 FILLER_28_139 ();
 sg13g2_decap_4 FILLER_28_156 ();
 sg13g2_fill_1 FILLER_28_160 ();
 sg13g2_fill_1 FILLER_28_199 ();
 sg13g2_decap_4 FILLER_28_204 ();
 sg13g2_fill_1 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_234 ();
 sg13g2_fill_1 FILLER_28_257 ();
 sg13g2_fill_1 FILLER_28_263 ();
 sg13g2_decap_8 FILLER_28_285 ();
 sg13g2_decap_8 FILLER_28_292 ();
 sg13g2_fill_1 FILLER_28_299 ();
 sg13g2_decap_8 FILLER_28_309 ();
 sg13g2_decap_4 FILLER_28_316 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_39 ();
 sg13g2_fill_2 FILLER_29_60 ();
 sg13g2_fill_2 FILLER_29_93 ();
 sg13g2_fill_2 FILLER_29_131 ();
 sg13g2_fill_1 FILLER_29_133 ();
 sg13g2_fill_1 FILLER_29_157 ();
 sg13g2_fill_1 FILLER_29_188 ();
 sg13g2_decap_8 FILLER_29_215 ();
 sg13g2_fill_1 FILLER_29_235 ();
 sg13g2_fill_2 FILLER_29_257 ();
 sg13g2_fill_1 FILLER_29_259 ();
 sg13g2_fill_2 FILLER_29_291 ();
 sg13g2_decap_8 FILLER_29_319 ();
 sg13g2_fill_2 FILLER_29_344 ();
 sg13g2_fill_1 FILLER_29_346 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_32 ();
 sg13g2_decap_8 FILLER_30_64 ();
 sg13g2_decap_8 FILLER_30_71 ();
 sg13g2_fill_1 FILLER_30_78 ();
 sg13g2_fill_2 FILLER_30_105 ();
 sg13g2_decap_4 FILLER_30_118 ();
 sg13g2_fill_2 FILLER_30_122 ();
 sg13g2_decap_8 FILLER_30_137 ();
 sg13g2_decap_4 FILLER_30_161 ();
 sg13g2_fill_2 FILLER_30_165 ();
 sg13g2_decap_4 FILLER_30_172 ();
 sg13g2_fill_2 FILLER_30_176 ();
 sg13g2_decap_8 FILLER_30_194 ();
 sg13g2_fill_2 FILLER_30_201 ();
 sg13g2_decap_8 FILLER_30_208 ();
 sg13g2_decap_4 FILLER_30_215 ();
 sg13g2_fill_2 FILLER_30_219 ();
 sg13g2_decap_8 FILLER_30_233 ();
 sg13g2_fill_1 FILLER_30_240 ();
 sg13g2_decap_4 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_262 ();
 sg13g2_fill_1 FILLER_30_271 ();
 sg13g2_fill_2 FILLER_30_373 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_4 ();
 sg13g2_fill_2 FILLER_31_19 ();
 sg13g2_fill_1 FILLER_31_21 ();
 sg13g2_fill_1 FILLER_31_40 ();
 sg13g2_decap_4 FILLER_31_53 ();
 sg13g2_fill_1 FILLER_31_57 ();
 sg13g2_decap_4 FILLER_31_63 ();
 sg13g2_fill_2 FILLER_31_67 ();
 sg13g2_decap_8 FILLER_31_95 ();
 sg13g2_fill_2 FILLER_31_102 ();
 sg13g2_fill_1 FILLER_31_104 ();
 sg13g2_fill_2 FILLER_31_121 ();
 sg13g2_fill_2 FILLER_31_136 ();
 sg13g2_fill_1 FILLER_31_138 ();
 sg13g2_fill_2 FILLER_31_156 ();
 sg13g2_fill_2 FILLER_31_176 ();
 sg13g2_fill_2 FILLER_31_199 ();
 sg13g2_fill_2 FILLER_31_239 ();
 sg13g2_decap_8 FILLER_31_262 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_9 ();
 sg13g2_fill_2 FILLER_32_34 ();
 sg13g2_fill_1 FILLER_32_36 ();
 sg13g2_decap_4 FILLER_32_62 ();
 sg13g2_fill_1 FILLER_32_66 ();
 sg13g2_decap_8 FILLER_32_93 ();
 sg13g2_fill_2 FILLER_32_100 ();
 sg13g2_fill_1 FILLER_32_102 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_fill_2 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_159 ();
 sg13g2_fill_2 FILLER_32_166 ();
 sg13g2_fill_2 FILLER_32_185 ();
 sg13g2_fill_1 FILLER_32_187 ();
 sg13g2_decap_8 FILLER_32_198 ();
 sg13g2_decap_8 FILLER_32_205 ();
 sg13g2_decap_8 FILLER_32_212 ();
 sg13g2_decap_4 FILLER_32_219 ();
 sg13g2_fill_2 FILLER_32_223 ();
 sg13g2_decap_4 FILLER_32_237 ();
 sg13g2_decap_8 FILLER_32_253 ();
 sg13g2_fill_2 FILLER_32_290 ();
 sg13g2_fill_1 FILLER_32_292 ();
 sg13g2_fill_1 FILLER_32_352 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_14 ();
 sg13g2_fill_2 FILLER_33_19 ();
 sg13g2_fill_1 FILLER_33_36 ();
 sg13g2_fill_1 FILLER_33_78 ();
 sg13g2_decap_4 FILLER_33_84 ();
 sg13g2_fill_2 FILLER_33_88 ();
 sg13g2_fill_2 FILLER_33_111 ();
 sg13g2_fill_2 FILLER_33_121 ();
 sg13g2_fill_1 FILLER_33_123 ();
 sg13g2_decap_8 FILLER_33_132 ();
 sg13g2_fill_1 FILLER_33_148 ();
 sg13g2_fill_2 FILLER_33_165 ();
 sg13g2_fill_1 FILLER_33_179 ();
 sg13g2_decap_4 FILLER_33_204 ();
 sg13g2_fill_1 FILLER_33_208 ();
 sg13g2_decap_4 FILLER_33_224 ();
 sg13g2_fill_1 FILLER_33_228 ();
 sg13g2_fill_1 FILLER_33_237 ();
 sg13g2_fill_1 FILLER_33_242 ();
 sg13g2_fill_1 FILLER_33_264 ();
 sg13g2_fill_2 FILLER_33_277 ();
 sg13g2_fill_1 FILLER_33_279 ();
 sg13g2_fill_1 FILLER_33_368 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_4 FILLER_34_21 ();
 sg13g2_fill_1 FILLER_34_25 ();
 sg13g2_decap_8 FILLER_34_30 ();
 sg13g2_decap_8 FILLER_34_37 ();
 sg13g2_decap_8 FILLER_34_44 ();
 sg13g2_fill_1 FILLER_34_56 ();
 sg13g2_fill_1 FILLER_34_109 ();
 sg13g2_fill_1 FILLER_34_135 ();
 sg13g2_decap_4 FILLER_34_183 ();
 sg13g2_fill_2 FILLER_34_187 ();
 sg13g2_decap_8 FILLER_34_206 ();
 sg13g2_fill_1 FILLER_34_213 ();
 sg13g2_fill_1 FILLER_34_258 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_4 FILLER_35_56 ();
 sg13g2_fill_2 FILLER_35_69 ();
 sg13g2_fill_1 FILLER_35_71 ();
 sg13g2_decap_4 FILLER_35_79 ();
 sg13g2_fill_2 FILLER_35_152 ();
 sg13g2_fill_1 FILLER_35_154 ();
 sg13g2_fill_1 FILLER_35_199 ();
 sg13g2_decap_4 FILLER_35_210 ();
 sg13g2_fill_2 FILLER_35_214 ();
 sg13g2_fill_1 FILLER_35_237 ();
 sg13g2_fill_1 FILLER_35_283 ();
 sg13g2_fill_1 FILLER_35_363 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_4 FILLER_36_42 ();
 sg13g2_fill_1 FILLER_36_75 ();
 sg13g2_decap_8 FILLER_36_165 ();
 sg13g2_fill_1 FILLER_36_172 ();
 sg13g2_decap_8 FILLER_36_177 ();
 sg13g2_decap_8 FILLER_36_184 ();
 sg13g2_fill_1 FILLER_36_194 ();
 sg13g2_fill_1 FILLER_36_215 ();
 sg13g2_fill_1 FILLER_36_224 ();
 sg13g2_fill_2 FILLER_36_256 ();
 sg13g2_fill_2 FILLER_36_277 ();
 sg13g2_fill_1 FILLER_36_360 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_4 FILLER_37_49 ();
 sg13g2_fill_1 FILLER_37_53 ();
 sg13g2_fill_2 FILLER_37_62 ();
 sg13g2_decap_8 FILLER_37_90 ();
 sg13g2_fill_1 FILLER_37_97 ();
 sg13g2_fill_1 FILLER_37_142 ();
 sg13g2_fill_1 FILLER_37_173 ();
 sg13g2_fill_1 FILLER_37_223 ();
 sg13g2_fill_2 FILLER_37_233 ();
 sg13g2_fill_1 FILLER_37_268 ();
 sg13g2_fill_1 FILLER_37_278 ();
 sg13g2_fill_2 FILLER_37_288 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_fill_1 FILLER_38_49 ();
 sg13g2_fill_1 FILLER_38_80 ();
 sg13g2_fill_2 FILLER_38_137 ();
 sg13g2_fill_1 FILLER_38_139 ();
 sg13g2_fill_2 FILLER_38_149 ();
 sg13g2_fill_2 FILLER_38_172 ();
 sg13g2_fill_1 FILLER_38_174 ();
 sg13g2_fill_2 FILLER_38_200 ();
 sg13g2_fill_1 FILLER_38_202 ();
 sg13g2_fill_2 FILLER_38_242 ();
 sg13g2_fill_2 FILLER_38_305 ();
 sg13g2_fill_1 FILLER_38_307 ();
 sg13g2_fill_1 FILLER_38_354 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net14;
 assign uio_oe[1] = net15;
 assign uio_oe[2] = net16;
 assign uio_oe[3] = net17;
 assign uio_oe[4] = net18;
 assign uio_oe[5] = net19;
 assign uio_oe[6] = net20;
 assign uio_oe[7] = net21;
 assign uio_out[0] = net22;
 assign uio_out[1] = net23;
 assign uio_out[2] = net24;
 assign uio_out[3] = net25;
 assign uio_out[4] = net26;
 assign uio_out[5] = net27;
 assign uio_out[6] = net28;
 assign uio_out[7] = net29;
 assign uo_out[2] = net30;
 assign uo_out[3] = net31;
 assign uo_out[4] = net32;
 assign uo_out[5] = net33;
 assign uo_out[6] = net34;
 assign uo_out[7] = net35;
endmodule

module tt_um_favoritohjs_scroller (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire clknet_0_clk;
 wire \bd[0] ;
 wire \bd[1] ;
 wire \bd[2] ;
 wire \color_ditherer.dither ;
 wire \color_ditherer.gin[0] ;
 wire \color_ditherer.gin[1] ;
 wire \color_ditherer.gin[2] ;
 wire \count1[0] ;
 wire \count1[1] ;
 wire \count1[2] ;
 wire \count1b[0] ;
 wire \count1b[1] ;
 wire \count1b[2] ;
 wire \count2[0] ;
 wire \count2[1] ;
 wire \count2b[0] ;
 wire \count2b[1] ;
 wire count2low;
 wire \cutoff1[0] ;
 wire \cutoff1[1] ;
 wire \cutoff1[2] ;
 wire \cutoff1[3] ;
 wire \cutoff1[4] ;
 wire \cutoff2[0] ;
 wire \cutoff2[1] ;
 wire \cutoff2[2] ;
 wire \cutoff2[3] ;
 wire \cutoff2[4] ;
 wire \hcount[0] ;
 wire \hcount[1] ;
 wire \hcount[2] ;
 wire \hcount[3] ;
 wire \hcount[4] ;
 wire \hcount[5] ;
 wire \hcount[6] ;
 wire \hcount[7] ;
 wire \hcount[8] ;
 wire \hcount[9] ;
 wire hsync;
 wire \l1[0] ;
 wire \l1[1] ;
 wire \l1[2] ;
 wire \l1[3] ;
 wire \l2[0] ;
 wire \l2[1] ;
 wire \l2[2] ;
 wire \l2[3] ;
 wire \lfsr1[4] ;
 wire \lfsr1[5] ;
 wire \lfsr1[6] ;
 wire \lfsr1[7] ;
 wire \lfsr1[8] ;
 wire \lfsr1[9] ;
 wire \lfsr1b[0] ;
 wire \lfsr1b[1] ;
 wire \lfsr1b[2] ;
 wire \lfsr1b[3] ;
 wire \lfsr1b[4] ;
 wire \lfsr1b[5] ;
 wire \lfsr1b[6] ;
 wire \lfsr1b[7] ;
 wire \lfsr1b[8] ;
 wire \lfsr1b[9] ;
 wire \lfsr2[4] ;
 wire \lfsr2[5] ;
 wire \lfsr2[6] ;
 wire \lfsr2[7] ;
 wire \lfsr2[8] ;
 wire \lfsr2[9] ;
 wire \lfsr2b[0] ;
 wire \lfsr2b[1] ;
 wire \lfsr2b[2] ;
 wire \lfsr2b[3] ;
 wire \lfsr2b[4] ;
 wire \lfsr2b[5] ;
 wire \lfsr2b[6] ;
 wire \lfsr2b[7] ;
 wire \lfsr2b[8] ;
 wire \lfsr2b[9] ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire vborder1;
 wire vborder2;
 wire \vcount[0] ;
 wire \vcount[1] ;
 wire \vcount[2] ;
 wire \vcount[3] ;
 wire \vcount[4] ;
 wire \vcount[5] ;
 wire \vcount[6] ;
 wire \vcount[7] ;
 wire \vcount[8] ;
 wire \vcount[9] ;
 wire \vga_sync.vga_vsync ;
 wire \vga_sync.xvisible ;
 wire \vga_sync.yvisible ;
 wire \vscheudler1.blockline[0] ;
 wire \vscheudler1.blockline[1] ;
 wire \vscheudler1.blockline[2] ;
 wire \vscheudler1.blockline[3] ;
 wire \vscheudler1.blockline[4] ;
 wire \vscheudler1.started ;
 wire \vscheudler2.blockline[0] ;
 wire \vscheudler2.blockline[1] ;
 wire \vscheudler2.blockline[2] ;
 wire \vscheudler2.blockline[3] ;
 wire \vscheudler2.blockline[4] ;
 wire \vscheudler2.started ;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net1;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;

 sg13g2_inv_1 _0659_ (.Y(_0120_),
    .A(\l2[2] ));
 sg13g2_inv_1 _0660_ (.Y(_0121_),
    .A(\l2[1] ));
 sg13g2_inv_1 _0661_ (.Y(_0122_),
    .A(net281));
 sg13g2_inv_1 _0662_ (.Y(_0123_),
    .A(net270));
 sg13g2_inv_1 _0663_ (.Y(_0124_),
    .A(net203));
 sg13g2_inv_1 _0664_ (.Y(_0125_),
    .A(net210));
 sg13g2_inv_1 _0665_ (.Y(_0126_),
    .A(net217));
 sg13g2_inv_1 _0666_ (.Y(_0127_),
    .A(\vscheudler2.blockline[3] ));
 sg13g2_inv_1 _0667_ (.Y(_0128_),
    .A(net266));
 sg13g2_inv_1 _0668_ (.Y(_0129_),
    .A(\cutoff2[3] ));
 sg13g2_inv_1 _0669_ (.Y(_0130_),
    .A(net316));
 sg13g2_inv_1 _0670_ (.Y(_0131_),
    .A(net301));
 sg13g2_inv_1 _0671_ (.Y(_0132_),
    .A(net340));
 sg13g2_inv_1 _0672_ (.Y(_0133_),
    .A(net248));
 sg13g2_inv_1 _0673_ (.Y(_0134_),
    .A(\vcount[6] ));
 sg13g2_inv_1 _0674_ (.Y(_0135_),
    .A(net198));
 sg13g2_inv_1 _0675_ (.Y(_0136_),
    .A(net275));
 sg13g2_inv_1 _0676_ (.Y(_0137_),
    .A(\color_ditherer.dither ));
 sg13g2_inv_1 _0677_ (.Y(_0138_),
    .A(net220));
 sg13g2_inv_1 _0678_ (.Y(_0139_),
    .A(net235));
 sg13g2_inv_1 _0679_ (.Y(_0140_),
    .A(net277));
 sg13g2_inv_1 _0680_ (.Y(_0141_),
    .A(net231));
 sg13g2_inv_1 _0681_ (.Y(_0142_),
    .A(net271));
 sg13g2_inv_1 _0682_ (.Y(_0143_),
    .A(net132));
 sg13g2_nor2_1 _0683_ (.A(\vcount[3] ),
    .B(\vcount[2] ),
    .Y(_0144_));
 sg13g2_or2_2 _0684_ (.X(_0145_),
    .B(\vcount[2] ),
    .A(\vcount[3] ));
 sg13g2_nand4_1 _0685_ (.B(\vcount[7] ),
    .C(\vcount[6] ),
    .A(\vcount[8] ),
    .Y(_0146_),
    .D(\vcount[5] ));
 sg13g2_nor3_1 _0686_ (.A(\vcount[9] ),
    .B(\vcount[4] ),
    .C(_0146_),
    .Y(_0147_));
 sg13g2_nand2b_1 _0687_ (.Y(_0148_),
    .B(net120),
    .A_N(\vcount[0] ));
 sg13g2_or4_2 _0688_ (.A(\vcount[9] ),
    .B(\vcount[4] ),
    .C(_0146_),
    .D(_0148_),
    .X(_0149_));
 sg13g2_nand3b_1 _0689_ (.B(\hcount[9] ),
    .C(\hcount[7] ),
    .Y(_0150_),
    .A_N(\hcount[8] ));
 sg13g2_or2_1 _0690_ (.X(_0151_),
    .B(net200),
    .A(\hcount[3] ));
 sg13g2_or4_2 _0691_ (.A(\hcount[0] ),
    .B(\hcount[1] ),
    .C(\hcount[3] ),
    .D(\hcount[2] ),
    .X(_0152_));
 sg13g2_nand2b_1 _0692_ (.Y(_0153_),
    .B(\hcount[4] ),
    .A_N(\hcount[5] ));
 sg13g2_nor4_2 _0693_ (.A(\hcount[6] ),
    .B(_0150_),
    .C(_0152_),
    .Y(_0154_),
    .D(_0153_));
 sg13g2_nor2_1 _0694_ (.A(\hcount[6] ),
    .B(_0150_),
    .Y(_0155_));
 sg13g2_nor4_2 _0695_ (.A(\hcount[6] ),
    .B(_0150_),
    .C(_0152_),
    .Y(_0156_),
    .D(_0153_));
 sg13g2_or4_1 _0696_ (.A(\hcount[6] ),
    .B(_0150_),
    .C(_0152_),
    .D(_0153_),
    .X(_0157_));
 sg13g2_nor3_2 _0697_ (.A(_0145_),
    .B(_0149_),
    .C(net110),
    .Y(_0158_));
 sg13g2_or3_1 _0698_ (.A(net185),
    .B(\count2b[1] ),
    .C(\count2b[0] ),
    .X(_0159_));
 sg13g2_nor4_2 _0699_ (.A(_0145_),
    .B(_0149_),
    .C(net109),
    .Y(_0160_),
    .D(_0159_));
 sg13g2_or4_1 _0700_ (.A(_0145_),
    .B(_0149_),
    .C(net109),
    .D(_0159_),
    .X(_0161_));
 sg13g2_xnor2_1 _0701_ (.Y(_0162_),
    .A(net235),
    .B(net255));
 sg13g2_a21oi_1 _0702_ (.A1(net264),
    .A2(net106),
    .Y(_0163_),
    .B1(net121));
 sg13g2_o21ai_1 _0703_ (.B1(_0163_),
    .Y(_0010_),
    .A1(net106),
    .A2(_0162_));
 sg13g2_a21oi_1 _0704_ (.A1(net280),
    .A2(net105),
    .Y(_0164_),
    .B1(net122));
 sg13g2_xnor2_1 _0705_ (.Y(_0165_),
    .A(net277),
    .B(net287));
 sg13g2_o21ai_1 _0706_ (.B1(_0164_),
    .Y(_0011_),
    .A1(net105),
    .A2(_0165_));
 sg13g2_nand2_1 _0707_ (.Y(_0166_),
    .A(net271),
    .B(_0160_));
 sg13g2_o21ai_1 _0708_ (.B1(net127),
    .Y(_0167_),
    .A1(net231),
    .A2(_0166_));
 sg13g2_a21o_1 _0709_ (.A2(_0166_),
    .A1(net231),
    .B1(_0167_),
    .X(_0012_));
 sg13g2_o21ai_1 _0710_ (.B1(net128),
    .Y(_0168_),
    .A1(net257),
    .A2(net106));
 sg13g2_a21oi_1 _0711_ (.A1(_0140_),
    .A2(net105),
    .Y(_0013_),
    .B1(_0168_));
 sg13g2_o21ai_1 _0712_ (.B1(net128),
    .Y(_0169_),
    .A1(net264),
    .A2(net106));
 sg13g2_a21oi_1 _0713_ (.A1(_0139_),
    .A2(_0161_),
    .Y(_0014_),
    .B1(_0169_));
 sg13g2_o21ai_1 _0714_ (.B1(net127),
    .Y(_0170_),
    .A1(net280),
    .A2(net105));
 sg13g2_a21oi_1 _0715_ (.A1(_0142_),
    .A2(net105),
    .Y(_0015_),
    .B1(_0170_));
 sg13g2_o21ai_1 _0716_ (.B1(net127),
    .Y(_0171_),
    .A1(\lfsr2b[7] ),
    .A2(_0160_));
 sg13g2_a21oi_1 _0717_ (.A1(_0141_),
    .A2(_0160_),
    .Y(_0016_),
    .B1(_0171_));
 sg13g2_o21ai_1 _0718_ (.B1(net128),
    .Y(_0172_),
    .A1(_0140_),
    .A2(net106));
 sg13g2_a21o_1 _0719_ (.A2(net105),
    .A1(net255),
    .B1(_0172_),
    .X(_0017_));
 sg13g2_o21ai_1 _0720_ (.B1(net128),
    .Y(_0173_),
    .A1(\lfsr2b[5] ),
    .A2(net106));
 sg13g2_a21oi_1 _0721_ (.A1(_0138_),
    .A2(net106),
    .Y(_0018_),
    .B1(_0173_));
 sg13g2_and2_2 _0722_ (.A(net243),
    .B(net191),
    .X(_0174_));
 sg13g2_nand2_2 _0723_ (.Y(_0175_),
    .A(\vga_sync.xvisible ),
    .B(net191));
 sg13g2_nor2_2 _0724_ (.A(_0154_),
    .B(_0174_),
    .Y(_0176_));
 sg13g2_nand3_1 _0725_ (.B(net111),
    .C(_0174_),
    .A(net171),
    .Y(_0177_));
 sg13g2_a22oi_1 _0726_ (.Y(_0178_),
    .B1(_0176_),
    .B2(\count2[0] ),
    .A2(_0156_),
    .A1(\count2b[0] ));
 sg13g2_nand3_1 _0727_ (.B(_0177_),
    .C(_0178_),
    .A(net129),
    .Y(_0019_));
 sg13g2_nand2_1 _0728_ (.Y(_0179_),
    .A(\count2[0] ),
    .B(_0174_));
 sg13g2_xor2_1 _0729_ (.B(_0179_),
    .A(net331),
    .X(_0180_));
 sg13g2_a21oi_1 _0730_ (.A1(net187),
    .A2(net114),
    .Y(_0181_),
    .B1(net122));
 sg13g2_o21ai_1 _0731_ (.B1(_0181_),
    .Y(_0020_),
    .A1(net114),
    .A2(net332));
 sg13g2_a21oi_1 _0732_ (.A1(net272),
    .A2(_0158_),
    .Y(_0182_),
    .B1(\count2b[0] ));
 sg13g2_nand3_1 _0733_ (.B(\count2b[0] ),
    .C(_0158_),
    .A(net272),
    .Y(_0183_));
 sg13g2_inv_1 _0734_ (.Y(_0184_),
    .A(_0183_));
 sg13g2_o21ai_1 _0735_ (.B1(net127),
    .Y(_0021_),
    .A1(net273),
    .A2(_0184_));
 sg13g2_a21oi_1 _0736_ (.A1(net187),
    .A2(_0183_),
    .Y(_0185_),
    .B1(net122));
 sg13g2_o21ai_1 _0737_ (.B1(_0185_),
    .Y(_0022_),
    .A1(net187),
    .A2(_0183_));
 sg13g2_nand2b_1 _0738_ (.Y(_0186_),
    .B(count2low),
    .A_N(_0158_));
 sg13g2_nand2_1 _0739_ (.Y(_0187_),
    .A(net185),
    .B(_0158_));
 sg13g2_nand3_1 _0740_ (.B(_0186_),
    .C(_0187_),
    .A(net127),
    .Y(_0023_));
 sg13g2_o21ai_1 _0741_ (.B1(net130),
    .Y(_0188_),
    .A1(net180),
    .A2(_0176_));
 sg13g2_a21oi_1 _0742_ (.A1(_0137_),
    .A2(_0176_),
    .Y(_0024_),
    .B1(_0188_));
 sg13g2_or2_1 _0743_ (.X(_0189_),
    .B(\hcount[7] ),
    .A(\hcount[6] ));
 sg13g2_nand2b_1 _0744_ (.Y(_0190_),
    .B(\hcount[5] ),
    .A_N(\hcount[4] ));
 sg13g2_nand2_1 _0745_ (.Y(_0191_),
    .A(net329),
    .B(\hcount[9] ));
 sg13g2_nor4_2 _0746_ (.A(_0152_),
    .B(_0189_),
    .C(_0190_),
    .Y(_0192_),
    .D(_0191_));
 sg13g2_nor2_2 _0747_ (.A(net123),
    .B(_0192_),
    .Y(_0193_));
 sg13g2_nand2b_2 _0748_ (.Y(_0194_),
    .B(net130),
    .A_N(_0192_));
 sg13g2_nand2b_1 _0749_ (.Y(_0025_),
    .B(_0193_),
    .A_N(net159));
 sg13g2_xnor2_1 _0750_ (.Y(_0195_),
    .A(\hcount[0] ),
    .B(net320));
 sg13g2_nor2_1 _0751_ (.A(_0194_),
    .B(net321),
    .Y(_0026_));
 sg13g2_and3_1 _0752_ (.X(_0196_),
    .A(\hcount[0] ),
    .B(\hcount[1] ),
    .C(net200));
 sg13g2_a21oi_1 _0753_ (.A1(\hcount[0] ),
    .A2(\hcount[1] ),
    .Y(_0197_),
    .B1(net200));
 sg13g2_nor3_1 _0754_ (.A(_0194_),
    .B(_0196_),
    .C(net201),
    .Y(_0027_));
 sg13g2_and4_2 _0755_ (.A(\hcount[0] ),
    .B(net320),
    .C(net251),
    .D(net200),
    .X(_0198_));
 sg13g2_nor2_1 _0756_ (.A(net251),
    .B(_0196_),
    .Y(_0199_));
 sg13g2_nor3_1 _0757_ (.A(_0194_),
    .B(_0198_),
    .C(net252),
    .Y(_0028_));
 sg13g2_xnor2_1 _0758_ (.Y(_0200_),
    .A(net352),
    .B(_0198_));
 sg13g2_nor2_1 _0759_ (.A(_0194_),
    .B(net353),
    .Y(_0029_));
 sg13g2_a21oi_1 _0760_ (.A1(\hcount[4] ),
    .A2(_0198_),
    .Y(_0201_),
    .B1(net322));
 sg13g2_and3_1 _0761_ (.X(_0202_),
    .A(net322),
    .B(net362),
    .C(_0198_));
 sg13g2_nor3_1 _0762_ (.A(_0194_),
    .B(net323),
    .C(_0202_),
    .Y(_0030_));
 sg13g2_nor2_1 _0763_ (.A(net346),
    .B(_0202_),
    .Y(_0203_));
 sg13g2_nand3_1 _0764_ (.B(\hcount[4] ),
    .C(\hcount[6] ),
    .A(net364),
    .Y(_0204_));
 sg13g2_and4_1 _0765_ (.A(net351),
    .B(\hcount[4] ),
    .C(\hcount[6] ),
    .D(_0198_),
    .X(_0205_));
 sg13g2_nor3_1 _0766_ (.A(_0194_),
    .B(_0203_),
    .C(_0205_),
    .Y(_0031_));
 sg13g2_nor2_1 _0767_ (.A(net253),
    .B(_0205_),
    .Y(_0206_));
 sg13g2_and2_1 _0768_ (.A(net253),
    .B(_0205_),
    .X(_0207_));
 sg13g2_nor3_1 _0769_ (.A(_0194_),
    .B(net254),
    .C(_0207_),
    .Y(_0032_));
 sg13g2_and2_1 _0770_ (.A(net329),
    .B(_0207_),
    .X(_0208_));
 sg13g2_o21ai_1 _0771_ (.B1(_0193_),
    .Y(_0209_),
    .A1(net329),
    .A2(_0207_));
 sg13g2_nor2_1 _0772_ (.A(_0208_),
    .B(_0209_),
    .Y(_0033_));
 sg13g2_nor2_1 _0773_ (.A(net284),
    .B(_0208_),
    .Y(_0210_));
 sg13g2_a21oi_1 _0774_ (.A1(net284),
    .A2(_0208_),
    .Y(_0211_),
    .B1(_0194_));
 sg13g2_nor2b_1 _0775_ (.A(net285),
    .B_N(_0211_),
    .Y(_0034_));
 sg13g2_nand2_2 _0776_ (.Y(_0212_),
    .A(net129),
    .B(_0174_));
 sg13g2_nor2b_1 _0777_ (.A(\l2[0] ),
    .B_N(\cutoff2[0] ),
    .Y(_0213_));
 sg13g2_o21ai_1 _0778_ (.B1(_0213_),
    .Y(_0214_),
    .A1(_0121_),
    .A2(\cutoff2[1] ));
 sg13g2_a22oi_1 _0779_ (.Y(_0215_),
    .B1(\cutoff2[1] ),
    .B2(_0121_),
    .A2(\cutoff2[2] ),
    .A1(_0120_));
 sg13g2_nor2_1 _0780_ (.A(_0120_),
    .B(\cutoff2[2] ),
    .Y(_0216_));
 sg13g2_a221oi_1 _0781_ (.B2(_0215_),
    .C1(_0216_),
    .B1(_0214_),
    .A1(\l2[3] ),
    .Y(_0217_),
    .A2(_0129_));
 sg13g2_nor2_1 _0782_ (.A(\l2[3] ),
    .B(_0129_),
    .Y(_0218_));
 sg13g2_or3_1 _0783_ (.A(\cutoff2[4] ),
    .B(_0217_),
    .C(_0218_),
    .X(_0219_));
 sg13g2_nand2b_1 _0784_ (.Y(_0220_),
    .B(\l1[3] ),
    .A_N(\cutoff1[3] ));
 sg13g2_nor2_1 _0785_ (.A(\l1[2] ),
    .B(_0132_),
    .Y(_0221_));
 sg13g2_nand2b_1 _0786_ (.Y(_0222_),
    .B(\cutoff1[0] ),
    .A_N(\l1[0] ));
 sg13g2_nand2b_1 _0787_ (.Y(_0223_),
    .B(\cutoff1[1] ),
    .A_N(\l1[1] ));
 sg13g2_nor2b_1 _0788_ (.A(\cutoff1[1] ),
    .B_N(\l1[1] ),
    .Y(_0224_));
 sg13g2_a221oi_1 _0789_ (.B2(_0223_),
    .C1(_0224_),
    .B1(_0222_),
    .A1(\l1[2] ),
    .Y(_0225_),
    .A2(_0132_));
 sg13g2_o21ai_1 _0790_ (.B1(_0220_),
    .Y(_0226_),
    .A1(_0221_),
    .A2(_0225_));
 sg13g2_nand2b_1 _0791_ (.Y(_0227_),
    .B(\cutoff1[3] ),
    .A_N(\l1[3] ));
 sg13g2_nand3_1 _0792_ (.B(_0226_),
    .C(_0227_),
    .A(_0131_),
    .Y(_0228_));
 sg13g2_nor2b_1 _0793_ (.A(net344),
    .B_N(net331),
    .Y(_0229_));
 sg13g2_nand2b_1 _0794_ (.Y(_0230_),
    .B(net331),
    .A_N(net344));
 sg13g2_nand3b_1 _0795_ (.B(_0229_),
    .C(_0219_),
    .Y(_0231_),
    .A_N(_0228_));
 sg13g2_nor2b_1 _0796_ (.A(_0212_),
    .B_N(_0231_),
    .Y(_0035_));
 sg13g2_o21ai_1 _0797_ (.B1(_0133_),
    .Y(_0232_),
    .A1(net361),
    .A2(\count1[1] ));
 sg13g2_nand2b_1 _0798_ (.Y(_0233_),
    .B(_0228_),
    .A_N(_0232_));
 sg13g2_a21oi_1 _0799_ (.A1(_0231_),
    .A2(_0233_),
    .Y(_0036_),
    .B1(_0212_));
 sg13g2_nand4_1 _0800_ (.B(_0174_),
    .C(_0228_),
    .A(net129),
    .Y(_0234_),
    .D(_0232_));
 sg13g2_inv_1 _0801_ (.Y(_0037_),
    .A(_0234_));
 sg13g2_nor2_1 _0802_ (.A(net347),
    .B(_0192_),
    .Y(_0235_));
 sg13g2_and2_2 _0803_ (.A(net363),
    .B(_0192_),
    .X(_0236_));
 sg13g2_nor4_1 _0804_ (.A(\vcount[7] ),
    .B(\vcount[6] ),
    .C(\vcount[5] ),
    .D(\vcount[4] ),
    .Y(_0237_));
 sg13g2_and2_1 _0805_ (.A(\vcount[3] ),
    .B(\vcount[2] ),
    .X(_0238_));
 sg13g2_nor2b_1 _0806_ (.A(net120),
    .B_N(\vcount[0] ),
    .Y(_0239_));
 sg13g2_nor2b_1 _0807_ (.A(\vcount[8] ),
    .B_N(\vcount[9] ),
    .Y(_0240_));
 sg13g2_nand4_1 _0808_ (.B(_0238_),
    .C(_0239_),
    .A(_0237_),
    .Y(_0241_),
    .D(_0240_));
 sg13g2_a21oi_1 _0809_ (.A1(net130),
    .A2(_0241_),
    .Y(_0242_),
    .B1(_0193_));
 sg13g2_a21o_1 _0810_ (.A2(_0241_),
    .A1(net130),
    .B1(_0193_),
    .X(_0243_));
 sg13g2_o21ai_1 _0811_ (.B1(_0243_),
    .Y(_0038_),
    .A1(net348),
    .A2(_0236_));
 sg13g2_a21oi_1 _0812_ (.A1(_0236_),
    .A2(_0241_),
    .Y(_0244_),
    .B1(net120));
 sg13g2_nand2b_1 _0813_ (.Y(_0245_),
    .B(net130),
    .A_N(_0244_));
 sg13g2_a21oi_1 _0814_ (.A1(net120),
    .A2(_0236_),
    .Y(_0039_),
    .B1(_0245_));
 sg13g2_and3_1 _0815_ (.X(_0246_),
    .A(net275),
    .B(net120),
    .C(_0236_));
 sg13g2_a21oi_1 _0816_ (.A1(net120),
    .A2(_0236_),
    .Y(_0247_),
    .B1(net275));
 sg13g2_nor3_1 _0817_ (.A(_0242_),
    .B(_0246_),
    .C(net276),
    .Y(_0040_));
 sg13g2_o21ai_1 _0818_ (.B1(_0243_),
    .Y(_0248_),
    .A1(net308),
    .A2(_0246_));
 sg13g2_and2_1 _0819_ (.A(net120),
    .B(_0238_),
    .X(_0249_));
 sg13g2_a21oi_1 _0820_ (.A1(net308),
    .A2(_0246_),
    .Y(_0041_),
    .B1(_0248_));
 sg13g2_a21oi_1 _0821_ (.A1(_0236_),
    .A2(_0249_),
    .Y(_0250_),
    .B1(net259));
 sg13g2_nand4_1 _0822_ (.B(net120),
    .C(_0236_),
    .A(net259),
    .Y(_0251_),
    .D(_0238_));
 sg13g2_nand2_1 _0823_ (.Y(_0252_),
    .A(net130),
    .B(_0251_));
 sg13g2_nor2_1 _0824_ (.A(_0250_),
    .B(_0252_),
    .Y(_0042_));
 sg13g2_and2_1 _0825_ (.A(net198),
    .B(net259),
    .X(_0253_));
 sg13g2_and4_2 _0826_ (.A(\vcount[0] ),
    .B(_0192_),
    .C(_0249_),
    .D(_0253_),
    .X(_0254_));
 sg13g2_nand2b_1 _0827_ (.Y(_0255_),
    .B(net127),
    .A_N(_0254_));
 sg13g2_a21oi_1 _0828_ (.A1(_0135_),
    .A2(_0251_),
    .Y(_0043_),
    .B1(_0255_));
 sg13g2_xnor2_1 _0829_ (.Y(_0256_),
    .A(net342),
    .B(_0254_));
 sg13g2_nor2_1 _0830_ (.A(net122),
    .B(net343),
    .Y(_0044_));
 sg13g2_a21o_1 _0831_ (.A2(_0254_),
    .A1(net342),
    .B1(net360),
    .X(_0257_));
 sg13g2_nand3_1 _0832_ (.B(net342),
    .C(_0254_),
    .A(net360),
    .Y(_0258_));
 sg13g2_and3_1 _0833_ (.X(_0045_),
    .A(net127),
    .B(_0257_),
    .C(_0258_));
 sg13g2_nand2b_1 _0834_ (.Y(_0259_),
    .B(_0258_),
    .A_N(net356));
 sg13g2_nand4_1 _0835_ (.B(\vcount[7] ),
    .C(\vcount[6] ),
    .A(net356),
    .Y(_0260_),
    .D(_0254_));
 sg13g2_and3_1 _0836_ (.X(_0046_),
    .A(net127),
    .B(net357),
    .C(_0260_));
 sg13g2_xor2_1 _0837_ (.B(_0260_),
    .A(net333),
    .X(_0261_));
 sg13g2_nor2_1 _0838_ (.A(_0242_),
    .B(net334),
    .Y(_0047_));
 sg13g2_a21oi_1 _0839_ (.A1(\color_ditherer.dither ),
    .A2(\bd[0] ),
    .Y(_0262_),
    .B1(net182));
 sg13g2_and3_1 _0840_ (.X(_0263_),
    .A(\color_ditherer.dither ),
    .B(\bd[0] ),
    .C(net182));
 sg13g2_nor3_1 _0841_ (.A(net123),
    .B(net183),
    .C(_0263_),
    .Y(_0048_));
 sg13g2_o21ai_1 _0842_ (.B1(net129),
    .Y(_0264_),
    .A1(net164),
    .A2(_0263_));
 sg13g2_a21oi_1 _0843_ (.A1(net164),
    .A2(_0263_),
    .Y(_0049_),
    .B1(_0264_));
 sg13g2_nand3_1 _0844_ (.B(_0147_),
    .C(_0239_),
    .A(_0144_),
    .Y(_0265_));
 sg13g2_nand2_1 _0845_ (.Y(_0266_),
    .A(net191),
    .B(_0265_));
 sg13g2_nor2_1 _0846_ (.A(\vcount[9] ),
    .B(\vcount[8] ),
    .Y(_0267_));
 sg13g2_nand4_1 _0847_ (.B(_0237_),
    .C(_0239_),
    .A(_0144_),
    .Y(_0268_),
    .D(_0267_));
 sg13g2_a21oi_1 _0848_ (.A1(_0266_),
    .A2(_0268_),
    .Y(_0050_),
    .B1(net123));
 sg13g2_nand2b_1 _0849_ (.Y(_0269_),
    .B(\hcount[0] ),
    .A_N(\hcount[1] ));
 sg13g2_nor4_2 _0850_ (.A(\hcount[5] ),
    .B(\hcount[4] ),
    .C(_0151_),
    .Y(_0270_),
    .D(_0269_));
 sg13g2_nand2_1 _0851_ (.Y(_0271_),
    .A(_0155_),
    .B(_0270_));
 sg13g2_nor3_1 _0852_ (.A(\hcount[8] ),
    .B(\hcount[9] ),
    .C(_0189_),
    .Y(_0272_));
 sg13g2_a22oi_1 _0853_ (.Y(_0273_),
    .B1(_0272_),
    .B2(_0270_),
    .A2(_0271_),
    .A1(net243));
 sg13g2_nor2_1 _0854_ (.A(net123),
    .B(net244),
    .Y(_0051_));
 sg13g2_nor3_1 _0855_ (.A(_0150_),
    .B(_0152_),
    .C(_0204_),
    .Y(_0274_));
 sg13g2_o21ai_1 _0856_ (.B1(net111),
    .Y(_0275_),
    .A1(net325),
    .A2(_0274_));
 sg13g2_nand2_1 _0857_ (.Y(_0052_),
    .A(net129),
    .B(_0275_));
 sg13g2_nand2_1 _0858_ (.Y(_0276_),
    .A(\vcount[3] ),
    .B(_0136_));
 sg13g2_nor2_1 _0859_ (.A(_0149_),
    .B(_0276_),
    .Y(_0277_));
 sg13g2_nor2_1 _0860_ (.A(\vcount[1] ),
    .B(\vcount[0] ),
    .Y(_0278_));
 sg13g2_nand3_1 _0861_ (.B(_0238_),
    .C(_0278_),
    .A(_0147_),
    .Y(_0279_));
 sg13g2_nor2b_1 _0862_ (.A(net291),
    .B_N(_0279_),
    .Y(_0280_));
 sg13g2_o21ai_1 _0863_ (.B1(net129),
    .Y(_0053_),
    .A1(_0277_),
    .A2(net292));
 sg13g2_a21oi_1 _0864_ (.A1(\color_ditherer.dither ),
    .A2(\color_ditherer.gin[0] ),
    .Y(_0281_),
    .B1(net175));
 sg13g2_and3_1 _0865_ (.X(_0282_),
    .A(\color_ditherer.dither ),
    .B(\color_ditherer.gin[0] ),
    .C(net175));
 sg13g2_nor3_1 _0866_ (.A(net123),
    .B(net176),
    .C(_0282_),
    .Y(_0054_));
 sg13g2_o21ai_1 _0867_ (.B1(net132),
    .Y(_0283_),
    .A1(net162),
    .A2(_0282_));
 sg13g2_a21oi_1 _0868_ (.A1(net162),
    .A2(_0282_),
    .Y(_0055_),
    .B1(_0283_));
 sg13g2_nor3_1 _0869_ (.A(net193),
    .B(net212),
    .C(\vscheudler1.blockline[1] ),
    .Y(_0284_));
 sg13g2_and3_1 _0870_ (.X(_0285_),
    .A(net316),
    .B(_0000_),
    .C(_0154_));
 sg13g2_and3_2 _0871_ (.X(_0286_),
    .A(\vscheudler1.started ),
    .B(_0000_),
    .C(net116));
 sg13g2_nand2_1 _0872_ (.Y(_0287_),
    .A(_0284_),
    .B(_0286_));
 sg13g2_and2_1 _0873_ (.A(net291),
    .B(net131),
    .X(_0288_));
 sg13g2_nand2_1 _0874_ (.Y(_0289_),
    .A(net291),
    .B(net130));
 sg13g2_and4_1 _0875_ (.A(net193),
    .B(net212),
    .C(\vscheudler1.blockline[1] ),
    .D(\vscheudler1.blockline[0] ),
    .X(_0290_));
 sg13g2_a221oi_1 _0876_ (.B2(_0286_),
    .C1(net118),
    .B1(_0290_),
    .A1(_0133_),
    .Y(_0056_),
    .A2(_0287_));
 sg13g2_nor2b_2 _0877_ (.A(net328),
    .B_N(_0284_),
    .Y(_0291_));
 sg13g2_nor4_1 _0878_ (.A(_0131_),
    .B(\cutoff1[3] ),
    .C(\cutoff1[2] ),
    .D(\cutoff1[0] ),
    .Y(_0292_));
 sg13g2_nand2b_1 _0879_ (.Y(_0293_),
    .B(_0292_),
    .A_N(\cutoff1[1] ));
 sg13g2_nand3_1 _0880_ (.B(_0291_),
    .C(_0293_),
    .A(_0286_),
    .Y(_0294_));
 sg13g2_nor2b_1 _0881_ (.A(\cutoff1[0] ),
    .B_N(_0294_),
    .Y(_0295_));
 sg13g2_nor2_1 _0882_ (.A(net166),
    .B(_0294_),
    .Y(_0296_));
 sg13g2_nor3_1 _0883_ (.A(net118),
    .B(_0295_),
    .C(_0296_),
    .Y(_0057_));
 sg13g2_nand3_1 _0884_ (.B(_0286_),
    .C(_0291_),
    .A(\cutoff1[0] ),
    .Y(_0297_));
 sg13g2_nor2b_1 _0885_ (.A(net303),
    .B_N(_0297_),
    .Y(_0298_));
 sg13g2_nand4_1 _0886_ (.B(\cutoff1[0] ),
    .C(_0285_),
    .A(net303),
    .Y(_0299_),
    .D(_0291_));
 sg13g2_and4_1 _0887_ (.A(net303),
    .B(\cutoff1[0] ),
    .C(_0286_),
    .D(_0291_),
    .X(_0300_));
 sg13g2_nor3_1 _0888_ (.A(net118),
    .B(net304),
    .C(_0300_),
    .Y(_0058_));
 sg13g2_o21ai_1 _0889_ (.B1(_0288_),
    .Y(_0301_),
    .A1(_0132_),
    .A2(_0299_));
 sg13g2_a21oi_1 _0890_ (.A1(_0132_),
    .A2(_0299_),
    .Y(_0059_),
    .B1(_0301_));
 sg13g2_a21o_1 _0891_ (.A2(_0300_),
    .A1(net340),
    .B1(net359),
    .X(_0302_));
 sg13g2_nand3_1 _0892_ (.B(net340),
    .C(_0300_),
    .A(net359),
    .Y(_0303_));
 sg13g2_and3_1 _0893_ (.X(_0060_),
    .A(_0288_),
    .B(_0302_),
    .C(_0303_));
 sg13g2_a21o_1 _0894_ (.A2(\cutoff1[3] ),
    .A1(net301),
    .B1(net117),
    .X(_0304_));
 sg13g2_a22oi_1 _0895_ (.Y(_0061_),
    .B1(_0304_),
    .B2(_0301_),
    .A2(_0303_),
    .A1(_0131_));
 sg13g2_o21ai_1 _0896_ (.B1(net328),
    .Y(_0305_),
    .A1(_0130_),
    .A2(net111));
 sg13g2_nand3b_1 _0897_ (.B(net116),
    .C(net316),
    .Y(_0306_),
    .A_N(net328));
 sg13g2_nand3_1 _0898_ (.B(_0305_),
    .C(_0306_),
    .A(net119),
    .Y(_0062_));
 sg13g2_or2_1 _0899_ (.X(_0307_),
    .B(_0306_),
    .A(net306));
 sg13g2_a21oi_1 _0900_ (.A1(net306),
    .A2(_0306_),
    .Y(_0308_),
    .B1(net117));
 sg13g2_nand2_1 _0901_ (.Y(_0063_),
    .A(_0307_),
    .B(net307));
 sg13g2_a21oi_1 _0902_ (.A1(net212),
    .A2(_0307_),
    .Y(_0309_),
    .B1(net117));
 sg13g2_o21ai_1 _0903_ (.B1(_0309_),
    .Y(_0064_),
    .A1(net212),
    .A2(_0307_));
 sg13g2_o21ai_1 _0904_ (.B1(net193),
    .Y(_0310_),
    .A1(\vscheudler1.blockline[2] ),
    .A2(_0307_));
 sg13g2_nand3_1 _0905_ (.B(net116),
    .C(_0291_),
    .A(\vscheudler1.started ),
    .Y(_0311_));
 sg13g2_nand2_1 _0906_ (.Y(_0312_),
    .A(net119),
    .B(_0311_));
 sg13g2_nand2b_1 _0907_ (.Y(_0065_),
    .B(net194),
    .A_N(_0312_));
 sg13g2_a21oi_1 _0908_ (.A1(\vscheudler1.started ),
    .A2(net116),
    .Y(_0313_),
    .B1(net168));
 sg13g2_nor3_1 _0909_ (.A(_0286_),
    .B(_0312_),
    .C(net169),
    .Y(_0066_));
 sg13g2_nor4_1 _0910_ (.A(\vcount[7] ),
    .B(_0134_),
    .C(net308),
    .D(_0136_),
    .Y(_0314_));
 sg13g2_nand4_1 _0911_ (.B(_0267_),
    .C(_0278_),
    .A(_0253_),
    .Y(_0315_),
    .D(_0314_));
 sg13g2_a21oi_1 _0912_ (.A1(_0130_),
    .A2(_0315_),
    .Y(_0067_),
    .B1(net117));
 sg13g2_nor4_2 _0913_ (.A(net225),
    .B(net208),
    .C(\vscheudler2.blockline[1] ),
    .Y(_0316_),
    .D(\vscheudler2.blockline[0] ));
 sg13g2_nand2_1 _0914_ (.Y(_0317_),
    .A(_0001_),
    .B(_0316_));
 sg13g2_xnor2_1 _0915_ (.Y(_0318_),
    .A(\vscheudler2.blockline[2] ),
    .B(\vscheudler2.blockline[1] ));
 sg13g2_nand4_1 _0916_ (.B(\vscheudler2.blockline[0] ),
    .C(_0001_),
    .A(_0127_),
    .Y(_0319_),
    .D(_0318_));
 sg13g2_nor2_2 _0917_ (.A(_0126_),
    .B(net111),
    .Y(_0320_));
 sg13g2_nand2_2 _0918_ (.Y(_0321_),
    .A(net217),
    .B(net114));
 sg13g2_a21oi_1 _0919_ (.A1(_0317_),
    .A2(_0319_),
    .Y(_0322_),
    .B1(_0321_));
 sg13g2_o21ai_1 _0920_ (.B1(net119),
    .Y(_0323_),
    .A1(vborder2),
    .A2(_0322_));
 sg13g2_a21oi_1 _0921_ (.A1(net208),
    .A2(_0322_),
    .Y(_0068_),
    .B1(_0323_));
 sg13g2_nand2b_1 _0922_ (.Y(_0324_),
    .B(\cutoff2[4] ),
    .A_N(\cutoff2[3] ));
 sg13g2_nor4_1 _0923_ (.A(\cutoff2[2] ),
    .B(\cutoff2[1] ),
    .C(\cutoff2[0] ),
    .D(_0324_),
    .Y(_0325_));
 sg13g2_nor4_2 _0924_ (.A(_0126_),
    .B(net111),
    .C(_0317_),
    .Y(_0326_),
    .D(_0325_));
 sg13g2_nor2_1 _0925_ (.A(\cutoff2[0] ),
    .B(_0326_),
    .Y(_0327_));
 sg13g2_nor2b_1 _0926_ (.A(net160),
    .B_N(_0326_),
    .Y(_0328_));
 sg13g2_nor3_1 _0927_ (.A(net117),
    .B(_0327_),
    .C(_0328_),
    .Y(_0069_));
 sg13g2_a21oi_1 _0928_ (.A1(\cutoff2[0] ),
    .A2(_0326_),
    .Y(_0329_),
    .B1(net282));
 sg13g2_and3_1 _0929_ (.X(_0330_),
    .A(net282),
    .B(\cutoff2[0] ),
    .C(_0326_));
 sg13g2_nor3_1 _0930_ (.A(net117),
    .B(net283),
    .C(_0330_),
    .Y(_0070_));
 sg13g2_nor2_1 _0931_ (.A(net338),
    .B(_0330_),
    .Y(_0331_));
 sg13g2_and2_1 _0932_ (.A(net338),
    .B(_0330_),
    .X(_0332_));
 sg13g2_nor3_1 _0933_ (.A(net118),
    .B(net339),
    .C(_0332_),
    .Y(_0071_));
 sg13g2_a21o_1 _0934_ (.A2(_0330_),
    .A1(net338),
    .B1(net350),
    .X(_0333_));
 sg13g2_nand3_1 _0935_ (.B(net338),
    .C(_0330_),
    .A(net350),
    .Y(_0334_));
 sg13g2_and3_1 _0936_ (.X(_0072_),
    .A(net119),
    .B(_0333_),
    .C(_0334_));
 sg13g2_nor2_1 _0937_ (.A(_0128_),
    .B(_0129_),
    .Y(_0335_));
 sg13g2_a221oi_1 _0938_ (.B2(_0332_),
    .C1(net118),
    .B1(_0335_),
    .A1(_0128_),
    .Y(_0073_),
    .A2(_0334_));
 sg13g2_nand2b_2 _0939_ (.Y(_0336_),
    .B(_0320_),
    .A_N(net330));
 sg13g2_a21oi_1 _0940_ (.A1(net330),
    .A2(_0321_),
    .Y(_0337_),
    .B1(net117));
 sg13g2_nand2_1 _0941_ (.Y(_0074_),
    .A(_0336_),
    .B(_0337_));
 sg13g2_a21oi_1 _0942_ (.A1(net314),
    .A2(_0336_),
    .Y(_0338_),
    .B1(net117));
 sg13g2_o21ai_1 _0943_ (.B1(_0338_),
    .Y(_0075_),
    .A1(net314),
    .A2(_0336_));
 sg13g2_or4_1 _0944_ (.A(net208),
    .B(net314),
    .C(net330),
    .D(_0321_),
    .X(_0339_));
 sg13g2_o21ai_1 _0945_ (.B1(net208),
    .Y(_0340_),
    .A1(net314),
    .A2(_0336_));
 sg13g2_nand3_1 _0946_ (.B(_0339_),
    .C(_0340_),
    .A(net119),
    .Y(_0076_));
 sg13g2_nand3_1 _0947_ (.B(net119),
    .C(_0339_),
    .A(net225),
    .Y(_0341_));
 sg13g2_nand3b_1 _0948_ (.B(net119),
    .C(_0316_),
    .Y(_0342_),
    .A_N(_0001_));
 sg13g2_o21ai_1 _0949_ (.B1(_0341_),
    .Y(_0077_),
    .A1(_0321_),
    .A2(_0342_));
 sg13g2_o21ai_1 _0950_ (.B1(_0320_),
    .Y(_0343_),
    .A1(_0001_),
    .A2(_0316_));
 sg13g2_o21ai_1 _0951_ (.B1(net119),
    .Y(_0344_),
    .A1(net214),
    .A2(_0320_));
 sg13g2_nor2b_1 _0952_ (.A(net215),
    .B_N(_0343_),
    .Y(_0078_));
 sg13g2_nor3_1 _0953_ (.A(\vcount[1] ),
    .B(\vcount[0] ),
    .C(_0276_),
    .Y(_0345_));
 sg13g2_and4_1 _0954_ (.A(\vcount[7] ),
    .B(_0134_),
    .C(_0253_),
    .D(_0267_),
    .X(_0346_));
 sg13g2_a21oi_1 _0955_ (.A1(_0345_),
    .A2(_0346_),
    .Y(_0347_),
    .B1(net217));
 sg13g2_nor2_1 _0956_ (.A(net118),
    .B(net218),
    .Y(_0079_));
 sg13g2_or2_1 _0957_ (.X(_0348_),
    .B(_0228_),
    .A(_0219_));
 sg13g2_mux2_1 _0958_ (.A0(_0230_),
    .A1(_0232_),
    .S(_0228_),
    .X(_0349_));
 sg13g2_a21oi_1 _0959_ (.A1(_0348_),
    .A2(_0349_),
    .Y(_0080_),
    .B1(_0212_));
 sg13g2_o21ai_1 _0960_ (.B1(_0234_),
    .Y(_0081_),
    .A1(_0212_),
    .A2(_0348_));
 sg13g2_nor2b_1 _0961_ (.A(_0212_),
    .B_N(_0348_),
    .Y(_0082_));
 sg13g2_nor4_2 _0962_ (.A(\count1[2] ),
    .B(\count1[1] ),
    .C(\count1[0] ),
    .Y(_0350_),
    .D(_0175_));
 sg13g2_nor2b_2 _0963_ (.A(_0154_),
    .B_N(_0350_),
    .Y(_0351_));
 sg13g2_nand3b_1 _0964_ (.B(net288),
    .C(net104),
    .Y(_0352_),
    .A_N(net205));
 sg13g2_nor2b_1 _0965_ (.A(net288),
    .B_N(_0351_),
    .Y(_0353_));
 sg13g2_nor2_1 _0966_ (.A(_0154_),
    .B(_0350_),
    .Y(_0354_));
 sg13g2_a21oi_1 _0967_ (.A1(net227),
    .A2(net116),
    .Y(_0355_),
    .B1(net124));
 sg13g2_a22oi_1 _0968_ (.Y(_0356_),
    .B1(_0354_),
    .B2(net245),
    .A2(_0353_),
    .A1(net205));
 sg13g2_nand3_1 _0969_ (.B(_0355_),
    .C(_0356_),
    .A(_0352_),
    .Y(_0083_));
 sg13g2_xor2_1 _0970_ (.B(net260),
    .A(net240),
    .X(_0357_));
 sg13g2_a21oi_1 _0971_ (.A1(net262),
    .A2(net115),
    .Y(_0358_),
    .B1(net126));
 sg13g2_a22oi_1 _0972_ (.Y(_0359_),
    .B1(_0357_),
    .B2(net104),
    .A2(net103),
    .A1(net324));
 sg13g2_nand2_1 _0973_ (.Y(_0084_),
    .A(_0358_),
    .B(_0359_));
 sg13g2_xor2_1 _0974_ (.B(\lfsr1[4] ),
    .A(net222),
    .X(_0360_));
 sg13g2_a21oi_1 _0975_ (.A1(net210),
    .A2(net115),
    .Y(_0361_),
    .B1(net124));
 sg13g2_a22oi_1 _0976_ (.Y(_0362_),
    .B1(_0360_),
    .B2(_0351_),
    .A2(net103),
    .A1(net299));
 sg13g2_nand2_1 _0977_ (.Y(_0085_),
    .A(_0361_),
    .B(net300));
 sg13g2_o21ai_1 _0978_ (.B1(net312),
    .Y(_0363_),
    .A1(_0353_),
    .A2(_0354_));
 sg13g2_a21oi_1 _0979_ (.A1(net203),
    .A2(net115),
    .Y(_0364_),
    .B1(net126));
 sg13g2_nand3b_1 _0980_ (.B(_0351_),
    .C(net288),
    .Y(_0365_),
    .A_N(net312));
 sg13g2_nand3_1 _0981_ (.B(_0364_),
    .C(_0365_),
    .A(_0363_),
    .Y(_0086_));
 sg13g2_a21oi_1 _0982_ (.A1(\lfsr1b[4] ),
    .A2(net115),
    .Y(_0366_),
    .B1(net125));
 sg13g2_a22oi_1 _0983_ (.Y(_0367_),
    .B1(net103),
    .B2(\lfsr1[4] ),
    .A2(net104),
    .A1(net245));
 sg13g2_nand2_1 _0984_ (.Y(_0087_),
    .A(_0366_),
    .B(net246));
 sg13g2_a21oi_1 _0985_ (.A1(net260),
    .A2(net103),
    .Y(_0368_),
    .B1(net126));
 sg13g2_a22oi_1 _0986_ (.Y(_0369_),
    .B1(net104),
    .B2(\l1[1] ),
    .A2(net115),
    .A1(\lfsr1b[5] ));
 sg13g2_nand2_1 _0987_ (.Y(_0088_),
    .A(_0368_),
    .B(_0369_));
 sg13g2_a21oi_1 _0988_ (.A1(\lfsr1b[6] ),
    .A2(net115),
    .Y(_0370_),
    .B1(net125));
 sg13g2_a22oi_1 _0989_ (.Y(_0371_),
    .B1(net103),
    .B2(net288),
    .A2(net104),
    .A1(\l1[2] ));
 sg13g2_nand2_1 _0990_ (.Y(_0089_),
    .A(_0370_),
    .B(net289));
 sg13g2_a21oi_1 _0991_ (.A1(\lfsr1b[7] ),
    .A2(net116),
    .Y(_0372_),
    .B1(net124));
 sg13g2_a22oi_1 _0992_ (.Y(_0373_),
    .B1(net103),
    .B2(net222),
    .A2(net104),
    .A1(\l1[3] ));
 sg13g2_nand2_1 _0993_ (.Y(_0090_),
    .A(_0372_),
    .B(net223));
 sg13g2_a21oi_1 _0994_ (.A1(\lfsr1b[8] ),
    .A2(net115),
    .Y(_0374_),
    .B1(net125));
 sg13g2_a22oi_1 _0995_ (.Y(_0375_),
    .B1(net103),
    .B2(net240),
    .A2(net104),
    .A1(\lfsr1[4] ));
 sg13g2_nand2_1 _0996_ (.Y(_0091_),
    .A(_0374_),
    .B(net241));
 sg13g2_a21oi_1 _0997_ (.A1(\lfsr1b[9] ),
    .A2(net115),
    .Y(_0376_),
    .B1(net125));
 sg13g2_a22oi_1 _0998_ (.Y(_0377_),
    .B1(net103),
    .B2(net205),
    .A2(net104),
    .A1(\lfsr1[5] ));
 sg13g2_nand2_1 _0999_ (.Y(_0092_),
    .A(_0376_),
    .B(net206));
 sg13g2_or3_1 _1000_ (.A(\count1b[2] ),
    .B(\count1b[1] ),
    .C(\count1b[0] ),
    .X(_0378_));
 sg13g2_nor4_2 _1001_ (.A(_0145_),
    .B(_0149_),
    .C(net109),
    .Y(_0379_),
    .D(_0378_));
 sg13g2_or4_2 _1002_ (.A(_0145_),
    .B(_0149_),
    .C(net108),
    .D(_0378_),
    .X(_0380_));
 sg13g2_a21oi_1 _1003_ (.A1(net227),
    .A2(net102),
    .Y(_0381_),
    .B1(net124));
 sg13g2_xnor2_1 _1004_ (.Y(_0382_),
    .A(net278),
    .B(\lfsr1b[6] ));
 sg13g2_o21ai_1 _1005_ (.B1(_0381_),
    .Y(_0093_),
    .A1(net102),
    .A2(net279));
 sg13g2_a21oi_1 _1006_ (.A1(net262),
    .A2(net101),
    .Y(_0383_),
    .B1(net126));
 sg13g2_xnor2_1 _1007_ (.Y(_0384_),
    .A(net281),
    .B(net295));
 sg13g2_o21ai_1 _1008_ (.B1(_0383_),
    .Y(_0094_),
    .A1(net101),
    .A2(_0384_));
 sg13g2_a21oi_1 _1009_ (.A1(net210),
    .A2(net102),
    .Y(_0385_),
    .B1(net124));
 sg13g2_xnor2_1 _1010_ (.Y(_0386_),
    .A(net270),
    .B(net250));
 sg13g2_o21ai_1 _1011_ (.B1(_0385_),
    .Y(_0095_),
    .A1(net102),
    .A2(_0386_));
 sg13g2_nand2_1 _1012_ (.Y(_0387_),
    .A(\lfsr1b[6] ),
    .B(_0379_));
 sg13g2_a21oi_1 _1013_ (.A1(net203),
    .A2(_0387_),
    .Y(_0388_),
    .B1(net124));
 sg13g2_o21ai_1 _1014_ (.B1(_0388_),
    .Y(_0096_),
    .A1(net203),
    .A2(_0387_));
 sg13g2_o21ai_1 _1015_ (.B1(net132),
    .Y(_0389_),
    .A1(_0123_),
    .A2(_0379_));
 sg13g2_a21o_1 _1016_ (.A2(_0379_),
    .A1(net227),
    .B1(_0389_),
    .X(_0097_));
 sg13g2_o21ai_1 _1017_ (.B1(net132),
    .Y(_0390_),
    .A1(_0122_),
    .A2(_0379_));
 sg13g2_a21o_1 _1018_ (.A2(_0379_),
    .A1(net262),
    .B1(_0390_),
    .X(_0098_));
 sg13g2_a21oi_1 _1019_ (.A1(\lfsr1b[6] ),
    .A2(net101),
    .Y(_0391_),
    .B1(net124));
 sg13g2_o21ai_1 _1020_ (.B1(_0391_),
    .Y(_0099_),
    .A1(_0125_),
    .A2(net102));
 sg13g2_a21oi_1 _1021_ (.A1(net250),
    .A2(net101),
    .Y(_0392_),
    .B1(net124));
 sg13g2_o21ai_1 _1022_ (.B1(_0392_),
    .Y(_0100_),
    .A1(_0124_),
    .A2(net102));
 sg13g2_a21oi_1 _1023_ (.A1(net295),
    .A2(net101),
    .Y(_0393_),
    .B1(net125));
 sg13g2_o21ai_1 _1024_ (.B1(_0393_),
    .Y(_0101_),
    .A1(_0123_),
    .A2(net101));
 sg13g2_a21oi_1 _1025_ (.A1(net278),
    .A2(net101),
    .Y(_0394_),
    .B1(net125));
 sg13g2_o21ai_1 _1026_ (.B1(_0394_),
    .Y(_0102_),
    .A1(_0122_),
    .A2(net101));
 sg13g2_nand3_1 _1027_ (.B(net111),
    .C(_0174_),
    .A(net178),
    .Y(_0395_));
 sg13g2_a22oi_1 _1028_ (.Y(_0396_),
    .B1(_0176_),
    .B2(\count1[0] ),
    .A2(net114),
    .A1(\count1b[0] ));
 sg13g2_nand3_1 _1029_ (.B(_0395_),
    .C(_0396_),
    .A(net129),
    .Y(_0103_));
 sg13g2_a21oi_1 _1030_ (.A1(\count1[1] ),
    .A2(\count1[0] ),
    .Y(_0397_),
    .B1(_0175_));
 sg13g2_o21ai_1 _1031_ (.B1(_0397_),
    .Y(_0398_),
    .A1(\count1[1] ),
    .A2(\count1[0] ));
 sg13g2_o21ai_1 _1032_ (.B1(net129),
    .Y(_0399_),
    .A1(net114),
    .A2(_0398_));
 sg13g2_a221oi_1 _1033_ (.B2(net345),
    .C1(_0399_),
    .B1(_0176_),
    .A1(net309),
    .Y(_0400_),
    .A2(net114));
 sg13g2_inv_1 _1034_ (.Y(_0104_),
    .A(_0400_));
 sg13g2_nand3_1 _1035_ (.B(net318),
    .C(_0174_),
    .A(\count1[1] ),
    .Y(_0401_));
 sg13g2_xor2_1 _1036_ (.B(net319),
    .A(net313),
    .X(_0402_));
 sg13g2_a21oi_1 _1037_ (.A1(net189),
    .A2(_0154_),
    .Y(_0403_),
    .B1(net123));
 sg13g2_o21ai_1 _1038_ (.B1(_0403_),
    .Y(_0105_),
    .A1(net114),
    .A2(_0402_));
 sg13g2_nand2b_1 _1039_ (.Y(_0404_),
    .B(\count1b[0] ),
    .A_N(_0158_));
 sg13g2_nand2_1 _1040_ (.Y(_0405_),
    .A(net173),
    .B(_0158_));
 sg13g2_nand3_1 _1041_ (.B(_0404_),
    .C(_0405_),
    .A(net128),
    .Y(_0106_));
 sg13g2_a21oi_1 _1042_ (.A1(\count1b[0] ),
    .A2(_0158_),
    .Y(_0406_),
    .B1(net309));
 sg13g2_nand3_1 _1043_ (.B(\count1b[0] ),
    .C(_0158_),
    .A(net309),
    .Y(_0407_));
 sg13g2_inv_1 _1044_ (.Y(_0408_),
    .A(_0407_));
 sg13g2_o21ai_1 _1045_ (.B1(net128),
    .Y(_0107_),
    .A1(net310),
    .A2(_0408_));
 sg13g2_a21oi_1 _1046_ (.A1(net189),
    .A2(_0407_),
    .Y(_0409_),
    .B1(net122));
 sg13g2_o21ai_1 _1047_ (.B1(_0409_),
    .Y(_0108_),
    .A1(net189),
    .A2(_0407_));
 sg13g2_and2_1 _1048_ (.A(\lfsr2[6] ),
    .B(net108),
    .X(_0410_));
 sg13g2_nand2_1 _1049_ (.Y(_0411_),
    .A(\lfsr2[6] ),
    .B(net108));
 sg13g2_nor3_2 _1050_ (.A(\count2[1] ),
    .B(\count2[0] ),
    .C(_0175_),
    .Y(_0412_));
 sg13g2_or3_2 _1051_ (.A(\count2[1] ),
    .B(\count2[0] ),
    .C(_0175_),
    .X(_0413_));
 sg13g2_nor2_1 _1052_ (.A(_0154_),
    .B(_0412_),
    .Y(_0414_));
 sg13g2_nand2_1 _1053_ (.Y(_0415_),
    .A(net108),
    .B(_0413_));
 sg13g2_nor2_1 _1054_ (.A(\lfsr2[6] ),
    .B(net113),
    .Y(_0416_));
 sg13g2_o21ai_1 _1055_ (.B1(_0415_),
    .Y(_0417_),
    .A1(net296),
    .A2(_0416_));
 sg13g2_a21oi_1 _1056_ (.A1(net296),
    .A2(_0411_),
    .Y(_0418_),
    .B1(_0417_));
 sg13g2_nand2b_1 _1057_ (.Y(_0419_),
    .B(net112),
    .A_N(net257));
 sg13g2_o21ai_1 _1058_ (.B1(_0419_),
    .Y(_0420_),
    .A1(\l2[0] ),
    .A2(_0415_));
 sg13g2_o21ai_1 _1059_ (.B1(net132),
    .Y(_0109_),
    .A1(net297),
    .A2(_0420_));
 sg13g2_nor2_1 _1060_ (.A(net268),
    .B(_0415_),
    .Y(_0421_));
 sg13g2_xnor2_1 _1061_ (.Y(_0422_),
    .A(\lfsr2[8] ),
    .B(\lfsr2[5] ));
 sg13g2_nand3_1 _1062_ (.B(net107),
    .C(_0422_),
    .A(net108),
    .Y(_0423_));
 sg13g2_o21ai_1 _1063_ (.B1(_0423_),
    .Y(_0424_),
    .A1(net264),
    .A2(net108));
 sg13g2_o21ai_1 _1064_ (.B1(net132),
    .Y(_0110_),
    .A1(_0421_),
    .A2(_0424_));
 sg13g2_nor2_1 _1065_ (.A(net196),
    .B(_0415_),
    .Y(_0425_));
 sg13g2_xnor2_1 _1066_ (.Y(_0426_),
    .A(\lfsr2[7] ),
    .B(net326));
 sg13g2_nand3_1 _1067_ (.B(net107),
    .C(net327),
    .A(net109),
    .Y(_0427_));
 sg13g2_o21ai_1 _1068_ (.B1(_0427_),
    .Y(_0428_),
    .A1(net280),
    .A2(net109));
 sg13g2_o21ai_1 _1069_ (.B1(net128),
    .Y(_0111_),
    .A1(_0425_),
    .A2(_0428_));
 sg13g2_a21oi_1 _1070_ (.A1(\lfsr2[6] ),
    .A2(net107),
    .Y(_0429_),
    .B1(net113));
 sg13g2_nor2b_1 _1071_ (.A(net335),
    .B_N(_0429_),
    .Y(_0430_));
 sg13g2_nand3_1 _1072_ (.B(net109),
    .C(_0412_),
    .A(\l2[3] ),
    .Y(_0431_));
 sg13g2_nand4_1 _1073_ (.B(net335),
    .C(net110),
    .A(\lfsr2[6] ),
    .Y(_0432_),
    .D(net107));
 sg13g2_o21ai_1 _1074_ (.B1(_0432_),
    .Y(_0433_),
    .A1(net231),
    .A2(net108));
 sg13g2_o21ai_1 _1075_ (.B1(net128),
    .Y(_0112_),
    .A1(net336),
    .A2(_0433_));
 sg13g2_nand2_1 _1076_ (.Y(_0434_),
    .A(net229),
    .B(_0413_));
 sg13g2_a21oi_1 _1077_ (.A1(\l2[0] ),
    .A2(net107),
    .Y(_0435_),
    .B1(net112));
 sg13g2_a221oi_1 _1078_ (.B2(_0435_),
    .C1(net121),
    .B1(_0434_),
    .A1(_0140_),
    .Y(_0113_),
    .A2(net112));
 sg13g2_nand3_1 _1079_ (.B(net110),
    .C(_0413_),
    .A(net233),
    .Y(_0436_));
 sg13g2_nor3_1 _1080_ (.A(_0121_),
    .B(net113),
    .C(_0413_),
    .Y(_0437_));
 sg13g2_a21oi_1 _1081_ (.A1(net235),
    .A2(net113),
    .Y(_0438_),
    .B1(_0437_));
 sg13g2_a21oi_1 _1082_ (.A1(_0436_),
    .A2(net236),
    .Y(_0114_),
    .B1(net121));
 sg13g2_nand3_1 _1083_ (.B(net109),
    .C(net107),
    .A(net196),
    .Y(_0439_));
 sg13g2_a22oi_1 _1084_ (.Y(_0440_),
    .B1(_0410_),
    .B2(_0413_),
    .A2(net112),
    .A1(\lfsr2b[6] ));
 sg13g2_a21oi_1 _1085_ (.A1(_0439_),
    .A2(_0440_),
    .Y(_0115_),
    .B1(net121));
 sg13g2_a22oi_1 _1086_ (.Y(_0441_),
    .B1(_0414_),
    .B2(net237),
    .A2(net112),
    .A1(\lfsr2b[7] ));
 sg13g2_a21oi_1 _1087_ (.A1(_0431_),
    .A2(net238),
    .Y(_0116_),
    .B1(net121));
 sg13g2_and2_1 _1088_ (.A(net294),
    .B(_0413_),
    .X(_0442_));
 sg13g2_a21oi_1 _1089_ (.A1(net229),
    .A2(net107),
    .Y(_0443_),
    .B1(_0442_));
 sg13g2_a21oi_1 _1090_ (.A1(net255),
    .A2(net112),
    .Y(_0444_),
    .B1(net121));
 sg13g2_o21ai_1 _1091_ (.B1(_0444_),
    .Y(_0117_),
    .A1(net112),
    .A2(_0443_));
 sg13g2_nand3_1 _1092_ (.B(net108),
    .C(net107),
    .A(net233),
    .Y(_0445_));
 sg13g2_a22oi_1 _1093_ (.Y(_0446_),
    .B1(_0414_),
    .B2(\lfsr2[9] ),
    .A2(net112),
    .A1(net220));
 sg13g2_a21oi_1 _1094_ (.A1(_0445_),
    .A2(_0446_),
    .Y(_0118_),
    .B1(net121));
 sg13g2_a21oi_1 _1095_ (.A1(net257),
    .A2(net105),
    .Y(_0447_),
    .B1(net121));
 sg13g2_xnor2_1 _1096_ (.Y(_0448_),
    .A(net220),
    .B(\lfsr2b[6] ));
 sg13g2_o21ai_1 _1097_ (.B1(_0447_),
    .Y(_0119_),
    .A1(net105),
    .A2(_0448_));
 sg13g2_dfrbp_1 _1098_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net38),
    .D(_0010_),
    .Q_N(_0548_),
    .Q(\lfsr2b[1] ));
 sg13g2_dfrbp_1 _1099_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net136),
    .D(_0011_),
    .Q_N(_0547_),
    .Q(\lfsr2b[2] ));
 sg13g2_dfrbp_1 _1100_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net134),
    .D(_0012_),
    .Q_N(_0546_),
    .Q(\lfsr2b[3] ));
 sg13g2_dfrbp_1 _1101_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net100),
    .D(_0013_),
    .Q_N(_0545_),
    .Q(\lfsr2b[4] ));
 sg13g2_dfrbp_1 _1102_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net98),
    .D(net265),
    .Q_N(_0544_),
    .Q(\lfsr2b[5] ));
 sg13g2_dfrbp_1 _1103_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net96),
    .D(_0015_),
    .Q_N(_0543_),
    .Q(\lfsr2b[6] ));
 sg13g2_dfrbp_1 _1104_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net94),
    .D(net232),
    .Q_N(_0542_),
    .Q(\lfsr2b[7] ));
 sg13g2_dfrbp_1 _1105_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net92),
    .D(net256),
    .Q_N(_0541_),
    .Q(\lfsr2b[8] ));
 sg13g2_dfrbp_1 _1106_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net90),
    .D(net221),
    .Q_N(_0540_),
    .Q(\lfsr2b[9] ));
 sg13g2_dfrbp_1 _1107_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net88),
    .D(net172),
    .Q_N(_0002_),
    .Q(\count2[0] ));
 sg13g2_dfrbp_1 _1108_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net86),
    .D(_0020_),
    .Q_N(_0539_),
    .Q(\count2[1] ));
 sg13g2_dfrbp_1 _1109_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net84),
    .D(net274),
    .Q_N(_0538_),
    .Q(\count2b[0] ));
 sg13g2_dfrbp_1 _1110_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net82),
    .D(net188),
    .Q_N(_0537_),
    .Q(\count2b[1] ));
 sg13g2_dfrbp_1 _1111_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net80),
    .D(net186),
    .Q_N(_0009_),
    .Q(count2low));
 sg13g2_dfrbp_1 _1112_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net78),
    .D(net181),
    .Q_N(_0004_),
    .Q(\color_ditherer.dither ));
 sg13g2_dfrbp_1 _1113_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net76),
    .D(_0025_),
    .Q_N(_0008_),
    .Q(\hcount[0] ));
 sg13g2_dfrbp_1 _1114_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net75),
    .D(_0026_),
    .Q_N(_0536_),
    .Q(\hcount[1] ));
 sg13g2_dfrbp_1 _1115_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net74),
    .D(net202),
    .Q_N(_0535_),
    .Q(\hcount[2] ));
 sg13g2_dfrbp_1 _1116_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net73),
    .D(_0028_),
    .Q_N(_0534_),
    .Q(\hcount[3] ));
 sg13g2_dfrbp_1 _1117_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net72),
    .D(_0029_),
    .Q_N(_0533_),
    .Q(\hcount[4] ));
 sg13g2_dfrbp_1 _1118_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net71),
    .D(_0030_),
    .Q_N(_0532_),
    .Q(\hcount[5] ));
 sg13g2_dfrbp_1 _1119_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net70),
    .D(_0031_),
    .Q_N(_0531_),
    .Q(\hcount[6] ));
 sg13g2_dfrbp_1 _1120_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net69),
    .D(_0032_),
    .Q_N(_0530_),
    .Q(\hcount[7] ));
 sg13g2_dfrbp_1 _1121_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net68),
    .D(_0033_),
    .Q_N(_0529_),
    .Q(\hcount[8] ));
 sg13g2_dfrbp_1 _1122_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net67),
    .D(net286),
    .Q_N(_0528_),
    .Q(\hcount[9] ));
 sg13g2_dfrbp_1 _1123_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net66),
    .D(_0035_),
    .Q_N(_0527_),
    .Q(\color_ditherer.gin[1] ));
 sg13g2_dfrbp_1 _1124_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net65),
    .D(_0036_),
    .Q_N(_0526_),
    .Q(\color_ditherer.gin[2] ));
 sg13g2_dfrbp_1 _1125_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net64),
    .D(_0037_),
    .Q_N(_0525_),
    .Q(\color_ditherer.gin[0] ));
 sg13g2_dfrbp_1 _1126_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net63),
    .D(net349),
    .Q_N(_0524_),
    .Q(\vcount[0] ));
 sg13g2_dfrbp_1 _1127_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net61),
    .D(net355),
    .Q_N(_0523_),
    .Q(\vcount[1] ));
 sg13g2_dfrbp_1 _1128_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net59),
    .D(_0040_),
    .Q_N(_0522_),
    .Q(\vcount[2] ));
 sg13g2_dfrbp_1 _1129_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net57),
    .D(_0041_),
    .Q_N(_0521_),
    .Q(\vcount[3] ));
 sg13g2_dfrbp_1 _1130_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net55),
    .D(_0042_),
    .Q_N(_0520_),
    .Q(\vcount[4] ));
 sg13g2_dfrbp_1 _1131_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net53),
    .D(net199),
    .Q_N(_0519_),
    .Q(\vcount[5] ));
 sg13g2_dfrbp_1 _1132_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net51),
    .D(_0044_),
    .Q_N(_0518_),
    .Q(\vcount[6] ));
 sg13g2_dfrbp_1 _1133_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net49),
    .D(_0045_),
    .Q_N(_0517_),
    .Q(\vcount[7] ));
 sg13g2_dfrbp_1 _1134_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net47),
    .D(net358),
    .Q_N(_0516_),
    .Q(\vcount[8] ));
 sg13g2_dfrbp_1 _1135_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net45),
    .D(_0047_),
    .Q_N(_0515_),
    .Q(\vcount[9] ));
 sg13g2_dfrbp_1 _1136_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net43),
    .D(net184),
    .Q_N(_0514_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _1137_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net42),
    .D(net165),
    .Q_N(_0513_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _1138_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net41),
    .D(net192),
    .Q_N(_0512_),
    .Q(\vga_sync.yvisible ));
 sg13g2_dfrbp_1 _1139_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net39),
    .D(_0051_),
    .Q_N(_0511_),
    .Q(\vga_sync.xvisible ));
 sg13g2_dfrbp_1 _1140_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net37),
    .D(_0052_),
    .Q_N(_0510_),
    .Q(hsync));
 sg13g2_dfrbp_1 _1141_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net35),
    .D(net293),
    .Q_N(_0509_),
    .Q(\vga_sync.vga_vsync ));
 sg13g2_dfrbp_1 _1142_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net33),
    .D(net177),
    .Q_N(_0508_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _1143_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net32),
    .D(net163),
    .Q_N(_0507_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _1144_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net31),
    .D(net249),
    .Q_N(_0506_),
    .Q(vborder1));
 sg13g2_dfrbp_1 _1145_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net29),
    .D(net167),
    .Q_N(_0007_),
    .Q(\cutoff1[0] ));
 sg13g2_dfrbp_1 _1146_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net27),
    .D(net305),
    .Q_N(_0505_),
    .Q(\cutoff1[1] ));
 sg13g2_dfrbp_1 _1147_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net25),
    .D(net341),
    .Q_N(_0504_),
    .Q(\cutoff1[2] ));
 sg13g2_dfrbp_1 _1148_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net23),
    .D(_0060_),
    .Q_N(_0503_),
    .Q(\cutoff1[3] ));
 sg13g2_dfrbp_1 _1149_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net21),
    .D(net302),
    .Q_N(_0502_),
    .Q(\cutoff1[4] ));
 sg13g2_dfrbp_1 _1150_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net19),
    .D(_0062_),
    .Q_N(_0501_),
    .Q(\vscheudler1.blockline[0] ));
 sg13g2_dfrbp_1 _1151_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net17),
    .D(_0063_),
    .Q_N(_0500_),
    .Q(\vscheudler1.blockline[1] ));
 sg13g2_dfrbp_1 _1152_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net157),
    .D(net213),
    .Q_N(_0499_),
    .Q(\vscheudler1.blockline[2] ));
 sg13g2_dfrbp_1 _1153_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net155),
    .D(net195),
    .Q_N(_0498_),
    .Q(\vscheudler1.blockline[3] ));
 sg13g2_dfrbp_1 _1154_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net153),
    .D(net170),
    .Q_N(_0000_),
    .Q(\vscheudler1.blockline[4] ));
 sg13g2_dfrbp_1 _1155_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net151),
    .D(net317),
    .Q_N(_0497_),
    .Q(\vscheudler1.started ));
 sg13g2_dfrbp_1 _1156_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net149),
    .D(net209),
    .Q_N(_0496_),
    .Q(vborder2));
 sg13g2_dfrbp_1 _1157_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net147),
    .D(net161),
    .Q_N(_0006_),
    .Q(\cutoff2[0] ));
 sg13g2_dfrbp_1 _1158_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net145),
    .D(_0070_),
    .Q_N(_0495_),
    .Q(\cutoff2[1] ));
 sg13g2_dfrbp_1 _1159_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net143),
    .D(_0071_),
    .Q_N(_0494_),
    .Q(\cutoff2[2] ));
 sg13g2_dfrbp_1 _1160_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net141),
    .D(_0072_),
    .Q_N(_0493_),
    .Q(\cutoff2[3] ));
 sg13g2_dfrbp_1 _1161_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net139),
    .D(net267),
    .Q_N(_0492_),
    .Q(\cutoff2[4] ));
 sg13g2_dfrbp_1 _1162_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net137),
    .D(_0074_),
    .Q_N(_0491_),
    .Q(\vscheudler2.blockline[0] ));
 sg13g2_dfrbp_1 _1163_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net133),
    .D(net315),
    .Q_N(_0490_),
    .Q(\vscheudler2.blockline[1] ));
 sg13g2_dfrbp_1 _1164_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net97),
    .D(_0076_),
    .Q_N(_0489_),
    .Q(\vscheudler2.blockline[2] ));
 sg13g2_dfrbp_1 _1165_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net93),
    .D(net226),
    .Q_N(_0488_),
    .Q(\vscheudler2.blockline[3] ));
 sg13g2_dfrbp_1 _1166_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net89),
    .D(net216),
    .Q_N(_0001_),
    .Q(\vscheudler2.blockline[4] ));
 sg13g2_dfrbp_1 _1167_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net85),
    .D(net219),
    .Q_N(_0487_),
    .Q(\vscheudler2.started ));
 sg13g2_dfrbp_1 _1168_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net81),
    .D(_0080_),
    .Q_N(_0486_),
    .Q(\bd[0] ));
 sg13g2_dfrbp_1 _1169_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net79),
    .D(_0081_),
    .Q_N(_0485_),
    .Q(\bd[1] ));
 sg13g2_dfrbp_1 _1170_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net77),
    .D(_0082_),
    .Q_N(_0484_),
    .Q(\bd[2] ));
 sg13g2_dfrbp_1 _1171_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net62),
    .D(_0083_),
    .Q_N(_0483_),
    .Q(\l1[0] ));
 sg13g2_dfrbp_1 _1172_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net58),
    .D(_0084_),
    .Q_N(_0482_),
    .Q(\l1[1] ));
 sg13g2_dfrbp_1 _1173_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net54),
    .D(_0085_),
    .Q_N(_0481_),
    .Q(\l1[2] ));
 sg13g2_dfrbp_1 _1174_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net50),
    .D(_0086_),
    .Q_N(_0480_),
    .Q(\l1[3] ));
 sg13g2_dfrbp_1 _1175_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net46),
    .D(net247),
    .Q_N(_0479_),
    .Q(\lfsr1[4] ));
 sg13g2_dfrbp_1 _1176_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net40),
    .D(net261),
    .Q_N(_0478_),
    .Q(\lfsr1[5] ));
 sg13g2_dfrbp_1 _1177_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net36),
    .D(net290),
    .Q_N(_0477_),
    .Q(\lfsr1[6] ));
 sg13g2_dfrbp_1 _1178_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net30),
    .D(net224),
    .Q_N(_0476_),
    .Q(\lfsr1[7] ));
 sg13g2_dfrbp_1 _1179_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net26),
    .D(net242),
    .Q_N(_0475_),
    .Q(\lfsr1[8] ));
 sg13g2_dfrbp_1 _1180_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net22),
    .D(net207),
    .Q_N(_0474_),
    .Q(\lfsr1[9] ));
 sg13g2_dfrbp_1 _1181_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net18),
    .D(_0093_),
    .Q_N(_0473_),
    .Q(\lfsr1b[0] ));
 sg13g2_dfrbp_1 _1182_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net156),
    .D(_0094_),
    .Q_N(_0472_),
    .Q(\lfsr1b[1] ));
 sg13g2_dfrbp_1 _1183_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net152),
    .D(_0095_),
    .Q_N(_0471_),
    .Q(\lfsr1b[2] ));
 sg13g2_dfrbp_1 _1184_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net148),
    .D(net204),
    .Q_N(_0470_),
    .Q(\lfsr1b[3] ));
 sg13g2_dfrbp_1 _1185_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net144),
    .D(net228),
    .Q_N(_0469_),
    .Q(\lfsr1b[4] ));
 sg13g2_dfrbp_1 _1186_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net140),
    .D(net263),
    .Q_N(_0468_),
    .Q(\lfsr1b[5] ));
 sg13g2_dfrbp_1 _1187_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net135),
    .D(net211),
    .Q_N(_0467_),
    .Q(\lfsr1b[6] ));
 sg13g2_dfrbp_1 _1188_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net95),
    .D(_0100_),
    .Q_N(_0466_),
    .Q(\lfsr1b[7] ));
 sg13g2_dfrbp_1 _1189_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net87),
    .D(_0101_),
    .Q_N(_0465_),
    .Q(\lfsr1b[8] ));
 sg13g2_dfrbp_1 _1190_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net60),
    .D(_0102_),
    .Q_N(_0464_),
    .Q(\lfsr1b[9] ));
 sg13g2_dfrbp_1 _1191_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net52),
    .D(net179),
    .Q_N(_0003_),
    .Q(\count1[0] ));
 sg13g2_dfrbp_1 _1192_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net44),
    .D(_0104_),
    .Q_N(_0463_),
    .Q(\count1[1] ));
 sg13g2_dfrbp_1 _1193_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net34),
    .D(_0105_),
    .Q_N(_0462_),
    .Q(\count1[2] ));
 sg13g2_dfrbp_1 _1194_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net24),
    .D(net174),
    .Q_N(_0005_),
    .Q(\count1b[0] ));
 sg13g2_dfrbp_1 _1195_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net158),
    .D(net311),
    .Q_N(_0461_),
    .Q(\count1b[1] ));
 sg13g2_dfrbp_1 _1196_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net150),
    .D(net190),
    .Q_N(_0460_),
    .Q(\count1b[2] ));
 sg13g2_dfrbp_1 _1197_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net142),
    .D(net298),
    .Q_N(_0459_),
    .Q(\l2[0] ));
 sg13g2_dfrbp_1 _1198_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net99),
    .D(net269),
    .Q_N(_0458_),
    .Q(\l2[1] ));
 sg13g2_dfrbp_1 _1199_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net83),
    .D(_0111_),
    .Q_N(_0457_),
    .Q(\l2[2] ));
 sg13g2_dfrbp_1 _1200_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net48),
    .D(net337),
    .Q_N(_0456_),
    .Q(\l2[3] ));
 sg13g2_dfrbp_1 _1201_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net28),
    .D(net230),
    .Q_N(_0455_),
    .Q(\lfsr2[4] ));
 sg13g2_dfrbp_1 _1202_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net154),
    .D(_0114_),
    .Q_N(_0454_),
    .Q(\lfsr2[5] ));
 sg13g2_dfrbp_1 _1203_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net138),
    .D(net197),
    .Q_N(_0453_),
    .Q(\lfsr2[6] ));
 sg13g2_dfrbp_1 _1204_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net56),
    .D(net239),
    .Q_N(_0452_),
    .Q(\lfsr2[7] ));
 sg13g2_dfrbp_1 _1205_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net20),
    .D(_0117_),
    .Q_N(_0451_),
    .Q(\lfsr2[8] ));
 sg13g2_dfrbp_1 _1206_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net91),
    .D(net234),
    .Q_N(_0450_),
    .Q(\lfsr2[9] ));
 sg13g2_dfrbp_1 _1207_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net146),
    .D(net258),
    .Q_N(_0449_),
    .Q(\lfsr2b[0] ));
 sg13g2_tiehi _1181__18 (.L_HI(net18));
 sg13g2_tiehi _1150__19 (.L_HI(net19));
 sg13g2_tiehi _1205__20 (.L_HI(net20));
 sg13g2_tiehi _1149__21 (.L_HI(net21));
 sg13g2_tiehi _1180__22 (.L_HI(net22));
 sg13g2_tiehi _1148__23 (.L_HI(net23));
 sg13g2_tiehi _1194__24 (.L_HI(net24));
 sg13g2_tiehi _1147__25 (.L_HI(net25));
 sg13g2_tiehi _1179__26 (.L_HI(net26));
 sg13g2_tiehi _1146__27 (.L_HI(net27));
 sg13g2_tiehi _1201__28 (.L_HI(net28));
 sg13g2_tiehi _1145__29 (.L_HI(net29));
 sg13g2_tiehi _1178__30 (.L_HI(net30));
 sg13g2_tiehi _1144__31 (.L_HI(net31));
 sg13g2_tiehi _1143__32 (.L_HI(net32));
 sg13g2_tiehi _1142__33 (.L_HI(net33));
 sg13g2_tiehi _1193__34 (.L_HI(net34));
 sg13g2_tiehi _1141__35 (.L_HI(net35));
 sg13g2_tiehi _1177__36 (.L_HI(net36));
 sg13g2_tiehi _1140__37 (.L_HI(net37));
 sg13g2_tiehi _1098__38 (.L_HI(net38));
 sg13g2_tiehi _1139__39 (.L_HI(net39));
 sg13g2_tiehi _1176__40 (.L_HI(net40));
 sg13g2_tiehi _1138__41 (.L_HI(net41));
 sg13g2_tiehi _1137__42 (.L_HI(net42));
 sg13g2_tiehi _1136__43 (.L_HI(net43));
 sg13g2_tiehi _1192__44 (.L_HI(net44));
 sg13g2_tiehi _1135__45 (.L_HI(net45));
 sg13g2_tiehi _1175__46 (.L_HI(net46));
 sg13g2_tiehi _1134__47 (.L_HI(net47));
 sg13g2_tiehi _1200__48 (.L_HI(net48));
 sg13g2_tiehi _1133__49 (.L_HI(net49));
 sg13g2_tiehi _1174__50 (.L_HI(net50));
 sg13g2_tiehi _1132__51 (.L_HI(net51));
 sg13g2_tiehi _1191__52 (.L_HI(net52));
 sg13g2_tiehi _1131__53 (.L_HI(net53));
 sg13g2_tiehi _1173__54 (.L_HI(net54));
 sg13g2_tiehi _1130__55 (.L_HI(net55));
 sg13g2_tiehi _1204__56 (.L_HI(net56));
 sg13g2_tiehi _1129__57 (.L_HI(net57));
 sg13g2_tiehi _1172__58 (.L_HI(net58));
 sg13g2_tiehi _1128__59 (.L_HI(net59));
 sg13g2_tiehi _1190__60 (.L_HI(net60));
 sg13g2_tiehi _1127__61 (.L_HI(net61));
 sg13g2_tiehi _1171__62 (.L_HI(net62));
 sg13g2_tiehi _1126__63 (.L_HI(net63));
 sg13g2_tiehi _1125__64 (.L_HI(net64));
 sg13g2_tiehi _1124__65 (.L_HI(net65));
 sg13g2_tiehi _1123__66 (.L_HI(net66));
 sg13g2_tiehi _1122__67 (.L_HI(net67));
 sg13g2_tiehi _1121__68 (.L_HI(net68));
 sg13g2_tiehi _1120__69 (.L_HI(net69));
 sg13g2_tiehi _1119__70 (.L_HI(net70));
 sg13g2_tiehi _1118__71 (.L_HI(net71));
 sg13g2_tiehi _1117__72 (.L_HI(net72));
 sg13g2_tiehi _1116__73 (.L_HI(net73));
 sg13g2_tiehi _1115__74 (.L_HI(net74));
 sg13g2_tiehi _1114__75 (.L_HI(net75));
 sg13g2_tiehi _1113__76 (.L_HI(net76));
 sg13g2_tiehi _1170__77 (.L_HI(net77));
 sg13g2_tiehi _1112__78 (.L_HI(net78));
 sg13g2_tiehi _1169__79 (.L_HI(net79));
 sg13g2_tiehi _1111__80 (.L_HI(net80));
 sg13g2_tiehi _1168__81 (.L_HI(net81));
 sg13g2_tiehi _1110__82 (.L_HI(net82));
 sg13g2_tiehi _1199__83 (.L_HI(net83));
 sg13g2_tiehi _1109__84 (.L_HI(net84));
 sg13g2_tiehi _1167__85 (.L_HI(net85));
 sg13g2_tiehi _1108__86 (.L_HI(net86));
 sg13g2_tiehi _1189__87 (.L_HI(net87));
 sg13g2_tiehi _1107__88 (.L_HI(net88));
 sg13g2_tiehi _1166__89 (.L_HI(net89));
 sg13g2_tiehi _1106__90 (.L_HI(net90));
 sg13g2_tiehi _1206__91 (.L_HI(net91));
 sg13g2_tiehi _1105__92 (.L_HI(net92));
 sg13g2_tiehi _1165__93 (.L_HI(net93));
 sg13g2_tiehi _1104__94 (.L_HI(net94));
 sg13g2_tiehi _1188__95 (.L_HI(net95));
 sg13g2_tiehi _1103__96 (.L_HI(net96));
 sg13g2_tiehi _1164__97 (.L_HI(net97));
 sg13g2_tiehi _1102__98 (.L_HI(net98));
 sg13g2_tiehi _1198__99 (.L_HI(net99));
 sg13g2_tiehi _1101__100 (.L_HI(net100));
 sg13g2_tiehi _1163__101 (.L_HI(net133));
 sg13g2_tiehi _1100__102 (.L_HI(net134));
 sg13g2_tiehi _1187__103 (.L_HI(net135));
 sg13g2_tiehi _1099__104 (.L_HI(net136));
 sg13g2_tiehi _1162__105 (.L_HI(net137));
 sg13g2_tiehi _1203__106 (.L_HI(net138));
 sg13g2_tiehi _1161__107 (.L_HI(net139));
 sg13g2_tiehi _1186__108 (.L_HI(net140));
 sg13g2_tiehi _1160__109 (.L_HI(net141));
 sg13g2_tiehi _1197__110 (.L_HI(net142));
 sg13g2_tiehi _1159__111 (.L_HI(net143));
 sg13g2_tiehi _1185__112 (.L_HI(net144));
 sg13g2_tiehi _1158__113 (.L_HI(net145));
 sg13g2_tiehi _1207__114 (.L_HI(net146));
 sg13g2_tiehi _1157__115 (.L_HI(net147));
 sg13g2_tiehi _1184__116 (.L_HI(net148));
 sg13g2_tiehi _1156__117 (.L_HI(net149));
 sg13g2_tiehi _1196__118 (.L_HI(net150));
 sg13g2_tiehi _1155__119 (.L_HI(net151));
 sg13g2_tiehi _1183__120 (.L_HI(net152));
 sg13g2_tiehi _1154__121 (.L_HI(net153));
 sg13g2_tiehi _1202__122 (.L_HI(net154));
 sg13g2_tiehi _1153__123 (.L_HI(net155));
 sg13g2_tiehi _1182__124 (.L_HI(net156));
 sg13g2_tiehi _1152__125 (.L_HI(net157));
 sg13g2_tiehi _1195__126 (.L_HI(net158));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_favoritohjs_scroller_2 (.L_LO(net2));
 sg13g2_tielo tt_um_favoritohjs_scroller_3 (.L_LO(net3));
 sg13g2_tielo tt_um_favoritohjs_scroller_4 (.L_LO(net4));
 sg13g2_tielo tt_um_favoritohjs_scroller_5 (.L_LO(net5));
 sg13g2_tielo tt_um_favoritohjs_scroller_6 (.L_LO(net6));
 sg13g2_tielo tt_um_favoritohjs_scroller_7 (.L_LO(net7));
 sg13g2_tielo tt_um_favoritohjs_scroller_8 (.L_LO(net8));
 sg13g2_tielo tt_um_favoritohjs_scroller_9 (.L_LO(net9));
 sg13g2_tielo tt_um_favoritohjs_scroller_10 (.L_LO(net10));
 sg13g2_tielo tt_um_favoritohjs_scroller_11 (.L_LO(net11));
 sg13g2_tielo tt_um_favoritohjs_scroller_12 (.L_LO(net12));
 sg13g2_tielo tt_um_favoritohjs_scroller_13 (.L_LO(net13));
 sg13g2_tielo tt_um_favoritohjs_scroller_14 (.L_LO(net14));
 sg13g2_tielo tt_um_favoritohjs_scroller_15 (.L_LO(net15));
 sg13g2_tielo tt_um_favoritohjs_scroller_16 (.L_LO(net16));
 sg13g2_tiehi _1151__17 (.L_HI(net17));
 sg13g2_buf_1 _1334_ (.A(uo_out[1]),
    .X(uo_out[0]));
 sg13g2_buf_1 _1335_ (.A(\vga_sync.vga_vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _1336_ (.A(uo_out[5]),
    .X(uo_out[4]));
 sg13g2_buf_1 _1337_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout101 (.A(_0380_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_0380_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_0354_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_0351_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(net106),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_0161_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_0412_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(net109),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(net110),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(net111),
    .X(net110));
 sg13g2_buf_4 fanout111 (.X(net111),
    .A(_0157_));
 sg13g2_buf_2 fanout112 (.A(net113),
    .X(net112));
 sg13g2_buf_1 fanout113 (.A(net114),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_0156_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(net116),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_0156_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(net118),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_0289_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_0288_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(net354),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(net122),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(net123),
    .X(net122));
 sg13g2_buf_4 fanout123 (.X(net123),
    .A(_0143_));
 sg13g2_buf_2 fanout124 (.A(net125),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(net126),
    .X(net125));
 sg13g2_buf_1 fanout126 (.A(_0143_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(net131),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(net131),
    .X(net128));
 sg13g2_buf_4 fanout129 (.X(net129),
    .A(net130));
 sg13g2_buf_4 fanout130 (.X(net130),
    .A(net131));
 sg13g2_buf_2 fanout131 (.A(net132),
    .X(net131));
 sg13g2_buf_4 fanout132 (.X(net132),
    .A(rst_n));
 sg13g2_tielo tt_um_favoritohjs_scroller_1 (.L_LO(net1));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0008_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0006_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0069_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold4 (.A(\color_ditherer.gin[2] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0055_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold6 (.A(\bd[2] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0049_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0007_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0057_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold10 (.A(\vscheudler1.blockline[4] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0313_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0066_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0002_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0019_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0005_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0106_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold17 (.A(\color_ditherer.gin[1] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0281_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0054_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0003_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0103_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0004_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0024_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold24 (.A(\bd[1] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0262_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0048_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0009_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0023_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold29 (.A(\count2b[1] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0022_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold31 (.A(\count1b[2] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0108_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold33 (.A(\vga_sync.yvisible ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0050_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold35 (.A(\vscheudler1.blockline[3] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0310_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0065_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold38 (.A(\l2[2] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0115_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold40 (.A(\vcount[5] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0043_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold42 (.A(\hcount[2] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0197_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0027_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold45 (.A(\lfsr1b[3] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0096_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold47 (.A(\lfsr1[9] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0377_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0092_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold50 (.A(\vscheudler2.blockline[2] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0068_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold52 (.A(\lfsr1b[2] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0099_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold54 (.A(\vscheudler1.blockline[2] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0064_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold56 (.A(\vscheudler2.blockline[4] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0344_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0078_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold59 (.A(\vscheudler2.started ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0347_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0079_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold62 (.A(\lfsr2b[9] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0018_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold64 (.A(\lfsr1[7] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0373_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0090_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold67 (.A(\vscheudler2.blockline[3] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0077_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold69 (.A(\lfsr1b[0] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0097_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold71 (.A(\lfsr2[4] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0113_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold73 (.A(\lfsr2b[3] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0016_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold75 (.A(\lfsr2[5] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0118_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold77 (.A(\lfsr2b[5] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0438_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold79 (.A(\lfsr2[7] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0441_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0116_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold82 (.A(\lfsr1[8] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0375_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0091_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold85 (.A(\vga_sync.xvisible ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0273_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold87 (.A(\l1[0] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0367_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0087_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold90 (.A(vborder1),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0056_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold92 (.A(\lfsr1b[7] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold93 (.A(\hcount[3] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0199_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold95 (.A(\hcount[7] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0206_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold97 (.A(\lfsr2b[8] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0017_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold99 (.A(\lfsr2b[0] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0119_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold101 (.A(\vcount[4] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold102 (.A(\lfsr1[5] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0088_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold104 (.A(\lfsr1b[1] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0098_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold106 (.A(\lfsr2b[1] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0014_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold108 (.A(\cutoff2[4] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0073_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold110 (.A(\l2[1] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0110_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold112 (.A(\lfsr1b[4] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold113 (.A(\lfsr2b[6] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold114 (.A(count2low),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0182_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0021_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold117 (.A(\vcount[2] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0247_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold119 (.A(\lfsr2b[4] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold120 (.A(\lfsr1b[9] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0382_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold122 (.A(\lfsr2b[2] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold123 (.A(\lfsr1b[5] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold124 (.A(\cutoff2[1] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0329_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold126 (.A(\hcount[9] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0210_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0034_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold129 (.A(\lfsr2b[7] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold130 (.A(\lfsr1[6] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0371_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0089_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold133 (.A(\vga_sync.vga_vsync ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0280_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0053_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold136 (.A(\lfsr2[8] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold137 (.A(\lfsr1b[8] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold138 (.A(\lfsr2[9] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0418_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0109_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold141 (.A(\l1[2] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0362_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold143 (.A(\cutoff1[4] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0061_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold145 (.A(\cutoff1[1] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0298_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0058_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold148 (.A(\vscheudler1.blockline[1] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0308_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold150 (.A(\vcount[3] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold151 (.A(\count1b[1] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0406_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0107_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold154 (.A(\l1[3] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold155 (.A(\count1[2] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold156 (.A(\vscheudler2.blockline[1] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0075_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold158 (.A(\vscheudler1.started ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0067_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold160 (.A(\count1[0] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0401_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold162 (.A(\hcount[1] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0195_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold164 (.A(\hcount[5] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0201_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold166 (.A(\l1[1] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold167 (.A(hsync),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold168 (.A(\lfsr2[4] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0426_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold170 (.A(\vscheudler1.blockline[0] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold171 (.A(\hcount[8] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold172 (.A(\vscheudler2.blockline[0] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold173 (.A(\count2[1] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0180_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold175 (.A(\vcount[9] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0261_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold177 (.A(\l2[3] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0430_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0112_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold180 (.A(\cutoff2[2] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0331_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold182 (.A(\cutoff1[2] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0059_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold184 (.A(\vcount[6] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0256_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold186 (.A(vborder2),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold187 (.A(\count1[1] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold188 (.A(\hcount[6] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold189 (.A(\vcount[0] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0235_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0038_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold192 (.A(\cutoff2[3] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold193 (.A(\hcount[5] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold194 (.A(\hcount[4] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0200_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold196 (.A(\vcount[1] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0039_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold198 (.A(\vcount[8] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0259_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0046_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold201 (.A(\cutoff1[3] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold202 (.A(\vcount[7] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold203 (.A(\count1[2] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold204 (.A(\hcount[4] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold205 (.A(\vcount[0] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold206 (.A(\hcount[5] ),
    .X(net364));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_4 FILLER_12_105 ();
 sg13g2_fill_2 FILLER_12_109 ();
 sg13g2_decap_8 FILLER_12_116 ();
 sg13g2_decap_8 FILLER_12_123 ();
 sg13g2_decap_8 FILLER_12_130 ();
 sg13g2_decap_8 FILLER_12_137 ();
 sg13g2_decap_8 FILLER_12_144 ();
 sg13g2_decap_8 FILLER_12_151 ();
 sg13g2_decap_8 FILLER_12_158 ();
 sg13g2_decap_8 FILLER_12_165 ();
 sg13g2_decap_8 FILLER_12_172 ();
 sg13g2_decap_8 FILLER_12_179 ();
 sg13g2_decap_8 FILLER_12_186 ();
 sg13g2_decap_8 FILLER_12_193 ();
 sg13g2_decap_8 FILLER_12_200 ();
 sg13g2_decap_8 FILLER_12_207 ();
 sg13g2_decap_8 FILLER_12_214 ();
 sg13g2_decap_8 FILLER_12_221 ();
 sg13g2_decap_8 FILLER_12_228 ();
 sg13g2_decap_8 FILLER_12_235 ();
 sg13g2_decap_8 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_249 ();
 sg13g2_decap_8 FILLER_12_256 ();
 sg13g2_decap_8 FILLER_12_263 ();
 sg13g2_decap_8 FILLER_12_270 ();
 sg13g2_decap_8 FILLER_12_277 ();
 sg13g2_decap_8 FILLER_12_284 ();
 sg13g2_decap_8 FILLER_12_291 ();
 sg13g2_decap_8 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_305 ();
 sg13g2_decap_8 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_decap_8 FILLER_12_326 ();
 sg13g2_decap_8 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_decap_8 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_4 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_4 FILLER_13_98 ();
 sg13g2_fill_1 FILLER_13_117 ();
 sg13g2_fill_2 FILLER_13_123 ();
 sg13g2_fill_1 FILLER_13_125 ();
 sg13g2_fill_1 FILLER_13_130 ();
 sg13g2_fill_1 FILLER_13_145 ();
 sg13g2_fill_2 FILLER_13_153 ();
 sg13g2_fill_1 FILLER_13_169 ();
 sg13g2_fill_1 FILLER_13_184 ();
 sg13g2_decap_8 FILLER_13_190 ();
 sg13g2_fill_2 FILLER_13_197 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_4 FILLER_13_294 ();
 sg13g2_fill_1 FILLER_13_298 ();
 sg13g2_decap_8 FILLER_13_303 ();
 sg13g2_fill_2 FILLER_13_310 ();
 sg13g2_fill_1 FILLER_13_312 ();
 sg13g2_decap_8 FILLER_13_316 ();
 sg13g2_decap_8 FILLER_13_323 ();
 sg13g2_fill_1 FILLER_13_330 ();
 sg13g2_decap_8 FILLER_13_335 ();
 sg13g2_fill_2 FILLER_13_342 ();
 sg13g2_decap_4 FILLER_13_347 ();
 sg13g2_fill_1 FILLER_13_351 ();
 sg13g2_decap_8 FILLER_13_361 ();
 sg13g2_decap_8 FILLER_13_368 ();
 sg13g2_decap_8 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_4 FILLER_13_403 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_fill_1 FILLER_14_91 ();
 sg13g2_fill_2 FILLER_14_101 ();
 sg13g2_fill_1 FILLER_14_103 ();
 sg13g2_fill_1 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_218 ();
 sg13g2_decap_8 FILLER_14_225 ();
 sg13g2_decap_8 FILLER_14_232 ();
 sg13g2_decap_8 FILLER_14_239 ();
 sg13g2_decap_8 FILLER_14_246 ();
 sg13g2_decap_8 FILLER_14_253 ();
 sg13g2_decap_8 FILLER_14_260 ();
 sg13g2_decap_8 FILLER_14_267 ();
 sg13g2_decap_4 FILLER_14_274 ();
 sg13g2_fill_2 FILLER_14_282 ();
 sg13g2_fill_2 FILLER_14_314 ();
 sg13g2_fill_1 FILLER_14_342 ();
 sg13g2_decap_4 FILLER_14_369 ();
 sg13g2_fill_2 FILLER_14_373 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_fill_2 FILLER_15_77 ();
 sg13g2_fill_1 FILLER_15_79 ();
 sg13g2_fill_1 FILLER_15_84 ();
 sg13g2_fill_2 FILLER_15_111 ();
 sg13g2_fill_1 FILLER_15_113 ();
 sg13g2_fill_1 FILLER_15_211 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_fill_1 FILLER_15_266 ();
 sg13g2_fill_1 FILLER_15_346 ();
 sg13g2_fill_1 FILLER_15_352 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_4 FILLER_16_63 ();
 sg13g2_fill_2 FILLER_16_67 ();
 sg13g2_fill_1 FILLER_16_102 ();
 sg13g2_fill_2 FILLER_16_163 ();
 sg13g2_fill_1 FILLER_16_174 ();
 sg13g2_fill_2 FILLER_16_180 ();
 sg13g2_fill_1 FILLER_16_182 ();
 sg13g2_fill_1 FILLER_16_225 ();
 sg13g2_fill_1 FILLER_16_242 ();
 sg13g2_decap_8 FILLER_16_251 ();
 sg13g2_fill_2 FILLER_16_258 ();
 sg13g2_fill_2 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_fill_1 FILLER_17_70 ();
 sg13g2_fill_1 FILLER_17_94 ();
 sg13g2_fill_1 FILLER_17_136 ();
 sg13g2_fill_1 FILLER_17_174 ();
 sg13g2_fill_1 FILLER_17_195 ();
 sg13g2_fill_2 FILLER_17_206 ();
 sg13g2_fill_1 FILLER_17_243 ();
 sg13g2_fill_1 FILLER_17_283 ();
 sg13g2_fill_2 FILLER_17_308 ();
 sg13g2_fill_2 FILLER_17_344 ();
 sg13g2_fill_2 FILLER_17_367 ();
 sg13g2_fill_1 FILLER_17_369 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_fill_2 FILLER_18_63 ();
 sg13g2_fill_1 FILLER_18_65 ();
 sg13g2_fill_1 FILLER_18_112 ();
 sg13g2_fill_2 FILLER_18_139 ();
 sg13g2_fill_2 FILLER_18_176 ();
 sg13g2_fill_1 FILLER_18_178 ();
 sg13g2_decap_4 FILLER_18_221 ();
 sg13g2_fill_2 FILLER_18_225 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_fill_2 FILLER_18_238 ();
 sg13g2_fill_2 FILLER_18_271 ();
 sg13g2_fill_1 FILLER_18_273 ();
 sg13g2_fill_2 FILLER_18_327 ();
 sg13g2_fill_1 FILLER_18_339 ();
 sg13g2_fill_1 FILLER_18_345 ();
 sg13g2_fill_1 FILLER_18_351 ();
 sg13g2_fill_1 FILLER_18_361 ();
 sg13g2_fill_1 FILLER_18_372 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_fill_1 FILLER_19_63 ();
 sg13g2_fill_1 FILLER_19_90 ();
 sg13g2_fill_2 FILLER_19_99 ();
 sg13g2_fill_1 FILLER_19_106 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_fill_1 FILLER_19_140 ();
 sg13g2_fill_1 FILLER_19_242 ();
 sg13g2_decap_8 FILLER_19_247 ();
 sg13g2_fill_1 FILLER_19_254 ();
 sg13g2_fill_1 FILLER_19_305 ();
 sg13g2_fill_2 FILLER_19_336 ();
 sg13g2_fill_1 FILLER_19_338 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_fill_2 FILLER_20_63 ();
 sg13g2_fill_1 FILLER_20_127 ();
 sg13g2_fill_2 FILLER_20_133 ();
 sg13g2_fill_1 FILLER_20_135 ();
 sg13g2_fill_1 FILLER_20_162 ();
 sg13g2_fill_2 FILLER_20_192 ();
 sg13g2_decap_8 FILLER_20_220 ();
 sg13g2_fill_2 FILLER_20_231 ();
 sg13g2_fill_1 FILLER_20_233 ();
 sg13g2_decap_8 FILLER_20_253 ();
 sg13g2_decap_4 FILLER_20_260 ();
 sg13g2_fill_1 FILLER_20_264 ();
 sg13g2_fill_1 FILLER_20_274 ();
 sg13g2_fill_2 FILLER_20_303 ();
 sg13g2_fill_1 FILLER_20_305 ();
 sg13g2_fill_1 FILLER_20_337 ();
 sg13g2_fill_2 FILLER_20_370 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_fill_2 FILLER_21_63 ();
 sg13g2_fill_1 FILLER_21_65 ();
 sg13g2_fill_2 FILLER_21_141 ();
 sg13g2_fill_2 FILLER_21_166 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_4 FILLER_21_238 ();
 sg13g2_decap_4 FILLER_21_257 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_fill_2 FILLER_21_321 ();
 sg13g2_fill_1 FILLER_21_323 ();
 sg13g2_fill_2 FILLER_21_342 ();
 sg13g2_fill_2 FILLER_21_351 ();
 sg13g2_fill_1 FILLER_21_353 ();
 sg13g2_fill_2 FILLER_21_369 ();
 sg13g2_fill_1 FILLER_21_371 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_fill_1 FILLER_22_89 ();
 sg13g2_fill_1 FILLER_22_130 ();
 sg13g2_fill_2 FILLER_22_139 ();
 sg13g2_fill_1 FILLER_22_141 ();
 sg13g2_decap_4 FILLER_22_173 ();
 sg13g2_fill_2 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_221 ();
 sg13g2_decap_4 FILLER_22_228 ();
 sg13g2_fill_2 FILLER_22_255 ();
 sg13g2_decap_8 FILLER_22_317 ();
 sg13g2_fill_1 FILLER_22_349 ();
 sg13g2_fill_1 FILLER_22_376 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_108 ();
 sg13g2_decap_4 FILLER_23_115 ();
 sg13g2_fill_1 FILLER_23_119 ();
 sg13g2_fill_2 FILLER_23_134 ();
 sg13g2_fill_1 FILLER_23_136 ();
 sg13g2_fill_1 FILLER_23_161 ();
 sg13g2_fill_2 FILLER_23_166 ();
 sg13g2_fill_2 FILLER_23_275 ();
 sg13g2_fill_2 FILLER_23_299 ();
 sg13g2_fill_1 FILLER_23_301 ();
 sg13g2_fill_2 FILLER_23_306 ();
 sg13g2_fill_1 FILLER_23_308 ();
 sg13g2_fill_1 FILLER_23_350 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_fill_2 FILLER_24_49 ();
 sg13g2_fill_1 FILLER_24_51 ();
 sg13g2_fill_2 FILLER_24_142 ();
 sg13g2_fill_2 FILLER_24_149 ();
 sg13g2_fill_1 FILLER_24_177 ();
 sg13g2_decap_8 FILLER_24_230 ();
 sg13g2_fill_2 FILLER_24_237 ();
 sg13g2_fill_1 FILLER_24_264 ();
 sg13g2_fill_2 FILLER_24_307 ();
 sg13g2_fill_1 FILLER_24_318 ();
 sg13g2_fill_2 FILLER_24_345 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_4 FILLER_25_14 ();
 sg13g2_fill_1 FILLER_25_18 ();
 sg13g2_decap_4 FILLER_25_99 ();
 sg13g2_decap_4 FILLER_25_116 ();
 sg13g2_fill_1 FILLER_25_169 ();
 sg13g2_fill_1 FILLER_25_264 ();
 sg13g2_fill_1 FILLER_25_270 ();
 sg13g2_fill_1 FILLER_25_298 ();
 sg13g2_fill_1 FILLER_25_325 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_4 FILLER_26_21 ();
 sg13g2_fill_1 FILLER_26_55 ();
 sg13g2_fill_2 FILLER_26_79 ();
 sg13g2_fill_2 FILLER_26_128 ();
 sg13g2_fill_2 FILLER_26_176 ();
 sg13g2_fill_1 FILLER_26_178 ();
 sg13g2_fill_2 FILLER_26_188 ();
 sg13g2_fill_1 FILLER_26_190 ();
 sg13g2_fill_2 FILLER_26_214 ();
 sg13g2_fill_1 FILLER_26_239 ();
 sg13g2_decap_8 FILLER_26_253 ();
 sg13g2_fill_2 FILLER_26_260 ();
 sg13g2_fill_1 FILLER_26_293 ();
 sg13g2_fill_1 FILLER_26_332 ();
 sg13g2_fill_2 FILLER_26_338 ();
 sg13g2_fill_1 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_4 FILLER_27_21 ();
 sg13g2_fill_1 FILLER_27_25 ();
 sg13g2_fill_2 FILLER_27_60 ();
 sg13g2_fill_1 FILLER_27_62 ();
 sg13g2_fill_2 FILLER_27_83 ();
 sg13g2_fill_2 FILLER_27_91 ();
 sg13g2_fill_1 FILLER_27_93 ();
 sg13g2_fill_2 FILLER_27_108 ();
 sg13g2_fill_2 FILLER_27_130 ();
 sg13g2_fill_2 FILLER_27_171 ();
 sg13g2_fill_1 FILLER_27_262 ();
 sg13g2_fill_1 FILLER_27_358 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_14 ();
 sg13g2_fill_1 FILLER_28_62 ();
 sg13g2_fill_1 FILLER_28_73 ();
 sg13g2_fill_1 FILLER_28_100 ();
 sg13g2_fill_2 FILLER_28_112 ();
 sg13g2_fill_1 FILLER_28_136 ();
 sg13g2_fill_2 FILLER_28_159 ();
 sg13g2_fill_1 FILLER_28_161 ();
 sg13g2_decap_4 FILLER_28_167 ();
 sg13g2_fill_1 FILLER_28_171 ();
 sg13g2_fill_1 FILLER_28_185 ();
 sg13g2_fill_2 FILLER_28_249 ();
 sg13g2_fill_2 FILLER_28_264 ();
 sg13g2_fill_2 FILLER_28_277 ();
 sg13g2_fill_1 FILLER_28_317 ();
 sg13g2_fill_1 FILLER_28_341 ();
 sg13g2_fill_1 FILLER_28_380 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_4 FILLER_29_21 ();
 sg13g2_fill_2 FILLER_29_48 ();
 sg13g2_fill_2 FILLER_29_71 ();
 sg13g2_fill_1 FILLER_29_73 ();
 sg13g2_fill_2 FILLER_29_98 ();
 sg13g2_fill_1 FILLER_29_100 ();
 sg13g2_fill_1 FILLER_29_124 ();
 sg13g2_fill_1 FILLER_29_168 ();
 sg13g2_fill_2 FILLER_29_173 ();
 sg13g2_decap_4 FILLER_29_181 ();
 sg13g2_fill_2 FILLER_29_193 ();
 sg13g2_fill_2 FILLER_29_247 ();
 sg13g2_fill_1 FILLER_29_281 ();
 sg13g2_fill_1 FILLER_29_320 ();
 sg13g2_fill_2 FILLER_29_328 ();
 sg13g2_fill_2 FILLER_29_348 ();
 sg13g2_fill_1 FILLER_29_358 ();
 sg13g2_decap_8 FILLER_29_396 ();
 sg13g2_decap_4 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_fill_1 FILLER_30_21 ();
 sg13g2_fill_1 FILLER_30_48 ();
 sg13g2_fill_2 FILLER_30_63 ();
 sg13g2_fill_1 FILLER_30_65 ();
 sg13g2_fill_1 FILLER_30_75 ();
 sg13g2_fill_1 FILLER_30_82 ();
 sg13g2_fill_1 FILLER_30_109 ();
 sg13g2_fill_1 FILLER_30_136 ();
 sg13g2_fill_2 FILLER_30_146 ();
 sg13g2_fill_1 FILLER_30_148 ();
 sg13g2_fill_1 FILLER_30_184 ();
 sg13g2_fill_2 FILLER_30_216 ();
 sg13g2_fill_2 FILLER_30_257 ();
 sg13g2_fill_2 FILLER_30_279 ();
 sg13g2_fill_2 FILLER_30_321 ();
 sg13g2_fill_1 FILLER_30_366 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_fill_1 FILLER_31_106 ();
 sg13g2_fill_1 FILLER_31_120 ();
 sg13g2_fill_2 FILLER_31_134 ();
 sg13g2_fill_1 FILLER_31_156 ();
 sg13g2_fill_1 FILLER_31_194 ();
 sg13g2_fill_1 FILLER_31_227 ();
 sg13g2_fill_2 FILLER_31_336 ();
 sg13g2_fill_2 FILLER_31_355 ();
 sg13g2_decap_8 FILLER_31_398 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_fill_2 FILLER_32_28 ();
 sg13g2_fill_1 FILLER_32_30 ();
 sg13g2_fill_2 FILLER_32_66 ();
 sg13g2_fill_2 FILLER_32_112 ();
 sg13g2_fill_1 FILLER_32_114 ();
 sg13g2_fill_2 FILLER_32_141 ();
 sg13g2_fill_2 FILLER_32_178 ();
 sg13g2_fill_1 FILLER_32_180 ();
 sg13g2_fill_1 FILLER_32_207 ();
 sg13g2_decap_4 FILLER_32_232 ();
 sg13g2_fill_2 FILLER_32_259 ();
 sg13g2_fill_1 FILLER_32_286 ();
 sg13g2_fill_2 FILLER_32_304 ();
 sg13g2_fill_1 FILLER_32_306 ();
 sg13g2_fill_2 FILLER_32_333 ();
 sg13g2_fill_1 FILLER_32_354 ();
 sg13g2_decap_8 FILLER_32_386 ();
 sg13g2_decap_8 FILLER_32_393 ();
 sg13g2_decap_8 FILLER_32_400 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_4 FILLER_33_35 ();
 sg13g2_fill_2 FILLER_33_69 ();
 sg13g2_fill_2 FILLER_33_89 ();
 sg13g2_fill_1 FILLER_33_105 ();
 sg13g2_fill_2 FILLER_33_118 ();
 sg13g2_fill_1 FILLER_33_129 ();
 sg13g2_fill_2 FILLER_33_139 ();
 sg13g2_fill_2 FILLER_33_145 ();
 sg13g2_fill_1 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_211 ();
 sg13g2_fill_2 FILLER_33_218 ();
 sg13g2_fill_1 FILLER_33_220 ();
 sg13g2_decap_4 FILLER_33_227 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_fill_2 FILLER_33_267 ();
 sg13g2_fill_1 FILLER_33_269 ();
 sg13g2_fill_2 FILLER_33_301 ();
 sg13g2_fill_1 FILLER_33_303 ();
 sg13g2_fill_2 FILLER_33_334 ();
 sg13g2_decap_8 FILLER_33_384 ();
 sg13g2_decap_8 FILLER_33_391 ();
 sg13g2_decap_8 FILLER_33_398 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_4 FILLER_34_28 ();
 sg13g2_fill_2 FILLER_34_78 ();
 sg13g2_fill_1 FILLER_34_106 ();
 sg13g2_fill_1 FILLER_34_117 ();
 sg13g2_fill_1 FILLER_34_124 ();
 sg13g2_fill_1 FILLER_34_156 ();
 sg13g2_fill_1 FILLER_34_188 ();
 sg13g2_fill_2 FILLER_34_219 ();
 sg13g2_fill_1 FILLER_34_221 ();
 sg13g2_fill_2 FILLER_34_243 ();
 sg13g2_fill_1 FILLER_34_245 ();
 sg13g2_fill_2 FILLER_34_272 ();
 sg13g2_fill_1 FILLER_34_274 ();
 sg13g2_fill_2 FILLER_34_284 ();
 sg13g2_fill_2 FILLER_34_291 ();
 sg13g2_fill_1 FILLER_34_293 ();
 sg13g2_decap_8 FILLER_34_325 ();
 sg13g2_fill_2 FILLER_34_332 ();
 sg13g2_fill_1 FILLER_34_338 ();
 sg13g2_decap_8 FILLER_34_366 ();
 sg13g2_decap_8 FILLER_34_373 ();
 sg13g2_decap_8 FILLER_34_380 ();
 sg13g2_decap_8 FILLER_34_387 ();
 sg13g2_decap_8 FILLER_34_394 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_4 FILLER_35_35 ();
 sg13g2_fill_2 FILLER_35_39 ();
 sg13g2_fill_1 FILLER_35_71 ();
 sg13g2_fill_2 FILLER_35_125 ();
 sg13g2_fill_1 FILLER_35_127 ();
 sg13g2_fill_1 FILLER_35_135 ();
 sg13g2_fill_2 FILLER_35_171 ();
 sg13g2_fill_2 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_222 ();
 sg13g2_fill_1 FILLER_35_229 ();
 sg13g2_fill_1 FILLER_35_263 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_decap_8 FILLER_35_322 ();
 sg13g2_decap_8 FILLER_35_329 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_4 FILLER_36_28 ();
 sg13g2_fill_2 FILLER_36_82 ();
 sg13g2_fill_2 FILLER_36_109 ();
 sg13g2_fill_1 FILLER_36_111 ();
 sg13g2_fill_2 FILLER_36_173 ();
 sg13g2_fill_2 FILLER_36_206 ();
 sg13g2_fill_2 FILLER_36_235 ();
 sg13g2_fill_1 FILLER_36_237 ();
 sg13g2_fill_2 FILLER_36_264 ();
 sg13g2_fill_1 FILLER_36_266 ();
 sg13g2_fill_1 FILLER_36_299 ();
 sg13g2_decap_8 FILLER_36_305 ();
 sg13g2_decap_8 FILLER_36_312 ();
 sg13g2_decap_8 FILLER_36_319 ();
 sg13g2_decap_8 FILLER_36_326 ();
 sg13g2_decap_8 FILLER_36_333 ();
 sg13g2_decap_8 FILLER_36_340 ();
 sg13g2_decap_8 FILLER_36_347 ();
 sg13g2_decap_8 FILLER_36_354 ();
 sg13g2_decap_8 FILLER_36_361 ();
 sg13g2_decap_8 FILLER_36_368 ();
 sg13g2_decap_8 FILLER_36_375 ();
 sg13g2_decap_8 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_36_389 ();
 sg13g2_decap_8 FILLER_36_396 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_4 FILLER_37_28 ();
 sg13g2_fill_2 FILLER_37_32 ();
 sg13g2_fill_2 FILLER_37_90 ();
 sg13g2_fill_2 FILLER_37_115 ();
 sg13g2_fill_2 FILLER_37_126 ();
 sg13g2_fill_2 FILLER_37_136 ();
 sg13g2_fill_1 FILLER_37_138 ();
 sg13g2_fill_2 FILLER_37_182 ();
 sg13g2_fill_1 FILLER_37_184 ();
 sg13g2_fill_2 FILLER_37_211 ();
 sg13g2_decap_8 FILLER_37_239 ();
 sg13g2_fill_2 FILLER_37_246 ();
 sg13g2_fill_1 FILLER_37_248 ();
 sg13g2_decap_8 FILLER_37_253 ();
 sg13g2_decap_4 FILLER_37_260 ();
 sg13g2_fill_2 FILLER_37_264 ();
 sg13g2_decap_8 FILLER_37_305 ();
 sg13g2_decap_8 FILLER_37_312 ();
 sg13g2_decap_8 FILLER_37_319 ();
 sg13g2_decap_8 FILLER_37_326 ();
 sg13g2_decap_8 FILLER_37_333 ();
 sg13g2_decap_8 FILLER_37_340 ();
 sg13g2_decap_8 FILLER_37_347 ();
 sg13g2_decap_8 FILLER_37_354 ();
 sg13g2_decap_8 FILLER_37_361 ();
 sg13g2_decap_8 FILLER_37_368 ();
 sg13g2_decap_8 FILLER_37_375 ();
 sg13g2_decap_8 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_396 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_fill_2 FILLER_38_95 ();
 sg13g2_fill_1 FILLER_38_97 ();
 sg13g2_fill_2 FILLER_38_133 ();
 sg13g2_fill_2 FILLER_38_144 ();
 sg13g2_fill_1 FILLER_38_146 ();
 sg13g2_fill_1 FILLER_38_188 ();
 sg13g2_fill_1 FILLER_38_224 ();
 sg13g2_decap_8 FILLER_38_234 ();
 sg13g2_decap_8 FILLER_38_241 ();
 sg13g2_decap_8 FILLER_38_248 ();
 sg13g2_decap_8 FILLER_38_255 ();
 sg13g2_decap_8 FILLER_38_262 ();
 sg13g2_fill_2 FILLER_38_269 ();
 sg13g2_fill_2 FILLER_38_280 ();
 sg13g2_decap_8 FILLER_38_286 ();
 sg13g2_decap_8 FILLER_38_293 ();
 sg13g2_decap_8 FILLER_38_300 ();
 sg13g2_decap_8 FILLER_38_307 ();
 sg13g2_decap_8 FILLER_38_314 ();
 sg13g2_decap_8 FILLER_38_321 ();
 sg13g2_decap_8 FILLER_38_328 ();
 sg13g2_decap_8 FILLER_38_335 ();
 sg13g2_decap_8 FILLER_38_342 ();
 sg13g2_decap_8 FILLER_38_349 ();
 sg13g2_decap_8 FILLER_38_356 ();
 sg13g2_decap_8 FILLER_38_363 ();
 sg13g2_decap_8 FILLER_38_370 ();
 sg13g2_decap_8 FILLER_38_377 ();
 sg13g2_decap_8 FILLER_38_384 ();
 sg13g2_decap_8 FILLER_38_391 ();
 sg13g2_decap_8 FILLER_38_398 ();
 sg13g2_decap_4 FILLER_38_405 ();
 assign uio_oe[0] = net1;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net3;
 assign uio_oe[3] = net4;
 assign uio_oe[4] = net5;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net8;
 assign uio_out[0] = net9;
 assign uio_out[1] = net10;
 assign uio_out[2] = net11;
 assign uio_out[3] = net12;
 assign uio_out[4] = net13;
 assign uio_out[5] = net14;
 assign uio_out[6] = net15;
 assign uio_out[7] = net16;
endmodule

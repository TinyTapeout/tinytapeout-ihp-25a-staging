module tt_um_tinytapeout_logo_screensaver (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire clknet_0_clk;
 wire \color_index[0] ;
 wire \color_index[1] ;
 wire \color_index[2] ;
 wire dir_x;
 wire dir_y;
 wire \gamepad.decoder.data_reg[0] ;
 wire \gamepad.decoder.data_reg[10] ;
 wire \gamepad.decoder.data_reg[11] ;
 wire \gamepad.decoder.data_reg[1] ;
 wire \gamepad.decoder.data_reg[2] ;
 wire \gamepad.decoder.data_reg[3] ;
 wire \gamepad.decoder.data_reg[4] ;
 wire \gamepad.decoder.data_reg[5] ;
 wire \gamepad.decoder.data_reg[6] ;
 wire \gamepad.decoder.data_reg[7] ;
 wire \gamepad.decoder.data_reg[8] ;
 wire \gamepad.decoder.data_reg[9] ;
 wire \gamepad.driver.pmod_clk_prev ;
 wire \gamepad.driver.pmod_clk_sync[0] ;
 wire \gamepad.driver.pmod_clk_sync[1] ;
 wire \gamepad.driver.pmod_data_sync[0] ;
 wire \gamepad.driver.pmod_data_sync[1] ;
 wire \gamepad.driver.pmod_latch_prev ;
 wire \gamepad.driver.pmod_latch_sync[0] ;
 wire \gamepad.driver.pmod_latch_sync[1] ;
 wire \gamepad.driver.shift_reg[0] ;
 wire \gamepad.driver.shift_reg[10] ;
 wire \gamepad.driver.shift_reg[11] ;
 wire \gamepad.driver.shift_reg[1] ;
 wire \gamepad.driver.shift_reg[2] ;
 wire \gamepad.driver.shift_reg[3] ;
 wire \gamepad.driver.shift_reg[4] ;
 wire \gamepad.driver.shift_reg[5] ;
 wire \gamepad.driver.shift_reg[6] ;
 wire \gamepad.driver.shift_reg[7] ;
 wire \gamepad.driver.shift_reg[8] ;
 wire \gamepad.driver.shift_reg[9] ;
 wire gamepad_start_prev;
 wire hsync;
 wire \logo_left[0] ;
 wire \logo_left[1] ;
 wire \logo_left[2] ;
 wire \logo_left[3] ;
 wire \logo_left[4] ;
 wire \logo_left[5] ;
 wire \logo_left[6] ;
 wire \logo_left[7] ;
 wire \logo_left[8] ;
 wire \logo_left[9] ;
 wire \logo_top[0] ;
 wire \logo_top[1] ;
 wire \logo_top[2] ;
 wire \logo_top[3] ;
 wire \logo_top[4] ;
 wire \logo_top[5] ;
 wire \logo_top[6] ;
 wire \logo_top[7] ;
 wire \logo_top[8] ;
 wire \logo_top[9] ;
 wire manual_mode;
 wire \palette_inst.rrggbb[0] ;
 wire \palette_inst.rrggbb[1] ;
 wire \palette_inst.rrggbb[2] ;
 wire \palette_inst.rrggbb[3] ;
 wire \palette_inst.rrggbb[4] ;
 wire \palette_inst.rrggbb[5] ;
 wire \pix_x[0] ;
 wire \pix_x[1] ;
 wire \pix_x[2] ;
 wire \pix_x[3] ;
 wire \pix_x[4] ;
 wire \pix_x[5] ;
 wire \pix_x[6] ;
 wire \pix_x[7] ;
 wire \pix_x[8] ;
 wire \pix_x[9] ;
 wire \pix_y[0] ;
 wire \pix_y[1] ;
 wire \pix_y[2] ;
 wire \pix_y[3] ;
 wire \pix_y[4] ;
 wire \pix_y[5] ;
 wire \pix_y[6] ;
 wire \pix_y[7] ;
 wire \pix_y[8] ;
 wire \pix_y[9] ;
 wire \prev_y[0] ;
 wire \prev_y[1] ;
 wire \prev_y[2] ;
 wire \prev_y[3] ;
 wire \prev_y[4] ;
 wire \prev_y[5] ;
 wire \prev_y[6] ;
 wire \prev_y[7] ;
 wire \prev_y[8] ;
 wire \prev_y[9] ;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire \vga_sync_gen.vsync ;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;

 sg13g2_inv_1 _1676_ (.Y(_0712_),
    .A(net201));
 sg13g2_inv_1 _1677_ (.Y(_0713_),
    .A(net205));
 sg13g2_inv_1 _1678_ (.Y(_0714_),
    .A(net197));
 sg13g2_inv_1 _1679_ (.Y(_0715_),
    .A(net193));
 sg13g2_inv_1 _1680_ (.Y(_0716_),
    .A(net198));
 sg13g2_inv_1 _1681_ (.Y(_0717_),
    .A(net203));
 sg13g2_inv_1 _1682_ (.Y(_0718_),
    .A(net210));
 sg13g2_inv_2 _1683_ (.Y(_0719_),
    .A(net189));
 sg13g2_inv_1 _1684_ (.Y(_0720_),
    .A(net211));
 sg13g2_inv_1 _1685_ (.Y(_0721_),
    .A(net191));
 sg13g2_inv_1 _1686_ (.Y(_0722_),
    .A(net183));
 sg13g2_inv_2 _1687_ (.Y(_0723_),
    .A(\gamepad.driver.pmod_data_sync[1] ));
 sg13g2_inv_1 _1688_ (.Y(_0724_),
    .A(net784));
 sg13g2_inv_1 _1689_ (.Y(_0725_),
    .A(net787));
 sg13g2_inv_2 _1690_ (.Y(_0726_),
    .A(net790));
 sg13g2_inv_1 _1691_ (.Y(_0727_),
    .A(net244));
 sg13g2_inv_1 _1692_ (.Y(_0728_),
    .A(net792));
 sg13g2_inv_1 _1693_ (.Y(_0729_),
    .A(net793));
 sg13g2_inv_1 _1694_ (.Y(_0730_),
    .A(\logo_top[3] ));
 sg13g2_inv_1 _1695_ (.Y(_0731_),
    .A(net795));
 sg13g2_inv_1 _1696_ (.Y(_0732_),
    .A(net797));
 sg13g2_inv_2 _1697_ (.Y(_0733_),
    .A(\logo_left[6] ));
 sg13g2_inv_2 _1698_ (.Y(_0734_),
    .A(\logo_left[5] ));
 sg13g2_inv_1 _1699_ (.Y(_0735_),
    .A(net800));
 sg13g2_inv_1 _1700_ (.Y(_0736_),
    .A(\logo_left[2] ));
 sg13g2_inv_1 _1701_ (.Y(_0737_),
    .A(net132));
 sg13g2_inv_1 _1702_ (.Y(_0738_),
    .A(net161));
 sg13g2_inv_1 _1703_ (.Y(_0739_),
    .A(\pix_y[0] ));
 sg13g2_inv_1 _1704_ (.Y(_0740_),
    .A(net778));
 sg13g2_inv_2 _1705_ (.Y(_0741_),
    .A(\pix_y[5] ));
 sg13g2_inv_1 _1706_ (.Y(_0742_),
    .A(\pix_y[6] ));
 sg13g2_inv_1 _1707_ (.Y(_0743_),
    .A(net807));
 sg13g2_inv_1 _1708_ (.Y(_0744_),
    .A(net245));
 sg13g2_inv_1 _1709_ (.Y(_0745_),
    .A(\prev_y[4] ));
 sg13g2_inv_1 _1710_ (.Y(_0746_),
    .A(\prev_y[5] ));
 sg13g2_inv_1 _1711_ (.Y(_0747_),
    .A(\prev_y[6] ));
 sg13g2_inv_1 _1712_ (.Y(_0748_),
    .A(net187));
 sg13g2_inv_1 _1713_ (.Y(_0749_),
    .A(net152));
 sg13g2_inv_1 _1714_ (.Y(_0750_),
    .A(net148));
 sg13g2_inv_1 _1715_ (.Y(_0751_),
    .A(net150));
 sg13g2_inv_1 _1716_ (.Y(_0752_),
    .A(net144));
 sg13g2_inv_1 _1717_ (.Y(_0753_),
    .A(net206));
 sg13g2_inv_1 _1718_ (.Y(_0754_),
    .A(net208));
 sg13g2_inv_1 _1719_ (.Y(_0755_),
    .A(net200));
 sg13g2_inv_1 _1720_ (.Y(_0756_),
    .A(net163));
 sg13g2_inv_1 _1721_ (.Y(_0757_),
    .A(net154));
 sg13g2_inv_1 _1722_ (.Y(_0758_),
    .A(net165));
 sg13g2_inv_1 _1723_ (.Y(_0759_),
    .A(net169));
 sg13g2_inv_1 _1724_ (.Y(_0760_),
    .A(net142));
 sg13g2_inv_1 _1725_ (.Y(_0761_),
    .A(_0010_));
 sg13g2_inv_1 _1726_ (.Y(_0762_),
    .A(net2));
 sg13g2_nor2_2 _1727_ (.A(_0741_),
    .B(_0742_),
    .Y(_0763_));
 sg13g2_nand3_1 _1728_ (.B(net185),
    .C(_0763_),
    .A(\pix_y[8] ),
    .Y(_0764_));
 sg13g2_or2_1 _1729_ (.X(_0765_),
    .B(net246),
    .A(net239));
 sg13g2_nand3b_1 _1730_ (.B(net779),
    .C(net781),
    .Y(_0766_),
    .A_N(net780));
 sg13g2_nor3_2 _1731_ (.A(net778),
    .B(_0765_),
    .C(_0766_),
    .Y(_0006_));
 sg13g2_and3_1 _1732_ (.X(_0767_),
    .A(\pix_x[4] ),
    .B(net803),
    .C(\pix_x[6] ));
 sg13g2_nand3b_1 _1733_ (.B(\pix_x[7] ),
    .C(net221),
    .Y(_0768_),
    .A_N(net216));
 sg13g2_nor3_1 _1734_ (.A(\pix_x[4] ),
    .B(\pix_x[5] ),
    .C(\pix_x[6] ),
    .Y(_0769_));
 sg13g2_nor3_2 _1735_ (.A(_0767_),
    .B(net222),
    .C(_0769_),
    .Y(_0005_));
 sg13g2_xnor2_1 _1736_ (.Y(_0770_),
    .A(\pix_y[9] ),
    .B(\prev_y[9] ));
 sg13g2_xnor2_1 _1737_ (.Y(_0771_),
    .A(\pix_y[8] ),
    .B(\prev_y[8] ));
 sg13g2_xnor2_1 _1738_ (.Y(_0772_),
    .A(net781),
    .B(\prev_y[1] ));
 sg13g2_a22oi_1 _1739_ (.Y(_0773_),
    .B1(\prev_y[6] ),
    .B2(_0742_),
    .A2(_0745_),
    .A1(net778));
 sg13g2_nand4_1 _1740_ (.B(_0771_),
    .C(_0772_),
    .A(_0770_),
    .Y(_0774_),
    .D(_0773_));
 sg13g2_xnor2_1 _1741_ (.Y(_0775_),
    .A(\pix_y[0] ),
    .B(\prev_y[0] ));
 sg13g2_xnor2_1 _1742_ (.Y(_0776_),
    .A(net777),
    .B(\prev_y[7] ));
 sg13g2_xor2_1 _1743_ (.B(\prev_y[2] ),
    .A(net780),
    .X(_0777_));
 sg13g2_a221oi_1 _1744_ (.B2(\pix_y[6] ),
    .C1(_0777_),
    .B1(_0747_),
    .A1(\pix_y[5] ),
    .Y(_0778_),
    .A2(_0746_));
 sg13g2_xor2_1 _1745_ (.B(\prev_y[3] ),
    .A(net779),
    .X(_0779_));
 sg13g2_a221oi_1 _1746_ (.B2(_0741_),
    .C1(_0779_),
    .B1(\prev_y[5] ),
    .A1(_0740_),
    .Y(_0780_),
    .A2(\prev_y[4] ));
 sg13g2_nand4_1 _1747_ (.B(_0776_),
    .C(_0778_),
    .A(_0775_),
    .Y(_0781_),
    .D(_0780_));
 sg13g2_nor4_1 _1748_ (.A(\pix_y[2] ),
    .B(net779),
    .C(\pix_y[8] ),
    .D(\pix_y[9] ),
    .Y(_0782_));
 sg13g2_or4_1 _1749_ (.A(net778),
    .B(\pix_y[5] ),
    .C(\pix_y[6] ),
    .D(net777),
    .X(_0783_));
 sg13g2_nor3_1 _1750_ (.A(\pix_y[0] ),
    .B(net781),
    .C(_0783_),
    .Y(_0784_));
 sg13g2_and2_1 _1751_ (.A(_0782_),
    .B(_0784_),
    .X(_0785_));
 sg13g2_o21ai_1 _1752_ (.B1(_0785_),
    .Y(_0786_),
    .A1(_0774_),
    .A2(_0781_));
 sg13g2_inv_1 _1753_ (.Y(_0787_),
    .A(_0786_));
 sg13g2_nor2_2 _1754_ (.A(net785),
    .B(_0786_),
    .Y(_0788_));
 sg13g2_inv_1 _1755_ (.Y(_0789_),
    .A(_0788_));
 sg13g2_and2_1 _1756_ (.A(net796),
    .B(net797),
    .X(_0790_));
 sg13g2_nand2_1 _1757_ (.Y(_0791_),
    .A(net796),
    .B(net797));
 sg13g2_and4_1 _1758_ (.A(\logo_top[3] ),
    .B(net795),
    .C(net796),
    .D(net797),
    .X(_0792_));
 sg13g2_nand3_1 _1759_ (.B(net794),
    .C(_0792_),
    .A(net793),
    .Y(_0793_));
 sg13g2_inv_1 _1760_ (.Y(_0794_),
    .A(_0793_));
 sg13g2_nor2_1 _1761_ (.A(_0013_),
    .B(_0793_),
    .Y(_0795_));
 sg13g2_xor2_1 _1762_ (.B(_0793_),
    .A(_0013_),
    .X(_0796_));
 sg13g2_xnor2_1 _1763_ (.Y(_0797_),
    .A(net792),
    .B(_0795_));
 sg13g2_nor2b_1 _1764_ (.A(_0796_),
    .B_N(_0797_),
    .Y(_0798_));
 sg13g2_and3_1 _1765_ (.X(_0799_),
    .A(net792),
    .B(\logo_top[6] ),
    .C(_0794_));
 sg13g2_nand2b_1 _1766_ (.Y(_0800_),
    .B(_0014_),
    .A_N(_0799_));
 sg13g2_nand3b_1 _1767_ (.B(_0799_),
    .C(net791),
    .Y(_0801_),
    .A_N(_0014_));
 sg13g2_o21ai_1 _1768_ (.B1(_0801_),
    .Y(_0802_),
    .A1(net791),
    .A2(_0800_));
 sg13g2_nor2_2 _1769_ (.A(net796),
    .B(net797),
    .Y(_0803_));
 sg13g2_nand2_1 _1770_ (.Y(_0804_),
    .A(_0011_),
    .B(_0803_));
 sg13g2_xnor2_1 _1771_ (.Y(_0805_),
    .A(\logo_top[3] ),
    .B(_0804_));
 sg13g2_nand4_1 _1772_ (.B(net797),
    .C(_0011_),
    .A(_0729_),
    .Y(_0806_),
    .D(_0012_));
 sg13g2_nor4_1 _1773_ (.A(net786),
    .B(net796),
    .C(_0805_),
    .D(_0806_),
    .Y(_0807_));
 sg13g2_nand3_1 _1774_ (.B(_0802_),
    .C(_0807_),
    .A(_0798_),
    .Y(_0808_));
 sg13g2_xnor2_1 _1775_ (.Y(_0809_),
    .A(_0014_),
    .B(_0799_));
 sg13g2_nor2b_1 _1776_ (.A(net791),
    .B_N(_0809_),
    .Y(_0810_));
 sg13g2_and2_1 _1777_ (.A(_0728_),
    .B(_0796_),
    .X(_0811_));
 sg13g2_a21oi_1 _1778_ (.A1(net794),
    .A2(_0792_),
    .Y(_0812_),
    .B1(net793));
 sg13g2_nor2_1 _1779_ (.A(_0794_),
    .B(_0812_),
    .Y(_0813_));
 sg13g2_xnor2_1 _1780_ (.Y(_0814_),
    .A(_0012_),
    .B(_0792_));
 sg13g2_nor2_1 _1781_ (.A(_0011_),
    .B(_0791_),
    .Y(_0815_));
 sg13g2_xnor2_1 _1782_ (.Y(_0816_),
    .A(_0730_),
    .B(_0815_));
 sg13g2_inv_1 _1783_ (.Y(_0817_),
    .A(_0816_));
 sg13g2_nor4_1 _1784_ (.A(_0731_),
    .B(_0791_),
    .C(_0814_),
    .D(_0816_),
    .Y(_0818_));
 sg13g2_and4_1 _1785_ (.A(_0810_),
    .B(_0811_),
    .C(_0813_),
    .D(_0818_),
    .X(_0819_));
 sg13g2_nand2_1 _1786_ (.Y(_0820_),
    .A(net787),
    .B(_0819_));
 sg13g2_and2_1 _1787_ (.A(_0808_),
    .B(_0820_),
    .X(_0821_));
 sg13g2_nor2_2 _1788_ (.A(\logo_left[1] ),
    .B(net802),
    .Y(_0822_));
 sg13g2_nand2_1 _1789_ (.Y(_0823_),
    .A(_0735_),
    .B(_0736_));
 sg13g2_nor3_2 _1790_ (.A(net801),
    .B(net802),
    .C(_0823_),
    .Y(_0824_));
 sg13g2_nand2_1 _1791_ (.Y(_0825_),
    .A(_0008_),
    .B(_0824_));
 sg13g2_xnor2_1 _1792_ (.Y(_0826_),
    .A(_0008_),
    .B(_0824_));
 sg13g2_nand2_1 _1793_ (.Y(_0827_),
    .A(_0007_),
    .B(_0822_));
 sg13g2_xnor2_1 _1794_ (.Y(_0828_),
    .A(_0735_),
    .B(_0827_));
 sg13g2_nand2_1 _1795_ (.Y(_0829_),
    .A(net802),
    .B(_0007_));
 sg13g2_nor4_1 _1796_ (.A(dir_x),
    .B(\logo_left[9] ),
    .C(net801),
    .D(_0829_),
    .Y(_0830_));
 sg13g2_nand2_1 _1797_ (.Y(_0831_),
    .A(_0828_),
    .B(_0830_));
 sg13g2_nor2_2 _1798_ (.A(\logo_left[5] ),
    .B(net799),
    .Y(_0832_));
 sg13g2_nand2_1 _1799_ (.Y(_0833_),
    .A(_0824_),
    .B(_0832_));
 sg13g2_nand3_1 _1800_ (.B(_0824_),
    .C(_0832_),
    .A(_0009_),
    .Y(_0834_));
 sg13g2_xnor2_1 _1801_ (.Y(_0835_),
    .A(_0009_),
    .B(_0833_));
 sg13g2_xnor2_1 _1802_ (.Y(_0836_),
    .A(_0734_),
    .B(_0825_));
 sg13g2_nand2_1 _1803_ (.Y(_0837_),
    .A(_0835_),
    .B(_0836_));
 sg13g2_or3_1 _1804_ (.A(net798),
    .B(\logo_left[6] ),
    .C(_0833_),
    .X(_0838_));
 sg13g2_nor2_1 _1805_ (.A(_0761_),
    .B(_0838_),
    .Y(_0839_));
 sg13g2_xnor2_1 _1806_ (.Y(_0840_),
    .A(_0761_),
    .B(_0838_));
 sg13g2_xor2_1 _1807_ (.B(_0834_),
    .A(net798),
    .X(_0841_));
 sg13g2_nand2b_1 _1808_ (.Y(_0842_),
    .B(_0841_),
    .A_N(_0840_));
 sg13g2_nor4_2 _1809_ (.A(_0826_),
    .B(_0831_),
    .C(_0837_),
    .Y(_0843_),
    .D(_0842_));
 sg13g2_nand2_2 _1810_ (.Y(_0844_),
    .A(net801),
    .B(net802));
 sg13g2_nand4_1 _1811_ (.B(\logo_left[2] ),
    .C(net801),
    .A(net800),
    .Y(_0845_),
    .D(net802));
 sg13g2_nand2_1 _1812_ (.Y(_0846_),
    .A(\logo_left[5] ),
    .B(net799));
 sg13g2_nor2_1 _1813_ (.A(_0845_),
    .B(_0846_),
    .Y(_0847_));
 sg13g2_and3_1 _1814_ (.X(_0848_),
    .A(net798),
    .B(\logo_left[6] ),
    .C(_0847_));
 sg13g2_and2_1 _1815_ (.A(_0761_),
    .B(_0848_),
    .X(_0849_));
 sg13g2_xnor2_1 _1816_ (.Y(_0850_),
    .A(\logo_left[9] ),
    .B(_0849_));
 sg13g2_xnor2_1 _1817_ (.Y(_0851_),
    .A(_0733_),
    .B(_0847_));
 sg13g2_nor2_1 _1818_ (.A(_0008_),
    .B(_0845_),
    .Y(_0852_));
 sg13g2_xnor2_1 _1819_ (.Y(_0853_),
    .A(_0734_),
    .B(_0852_));
 sg13g2_xor2_1 _1820_ (.B(_0845_),
    .A(net799),
    .X(_0854_));
 sg13g2_nor2_1 _1821_ (.A(_0007_),
    .B(_0844_),
    .Y(_0855_));
 sg13g2_xnor2_1 _1822_ (.Y(_0856_),
    .A(net800),
    .B(_0855_));
 sg13g2_nor3_1 _1823_ (.A(_0726_),
    .B(_0736_),
    .C(_0844_),
    .Y(_0857_));
 sg13g2_nand3_1 _1824_ (.B(_0856_),
    .C(_0857_),
    .A(_0854_),
    .Y(_0858_));
 sg13g2_nor3_1 _1825_ (.A(_0009_),
    .B(_0845_),
    .C(_0846_),
    .Y(_0859_));
 sg13g2_xnor2_1 _1826_ (.Y(_0860_),
    .A(net798),
    .B(_0859_));
 sg13g2_xor2_1 _1827_ (.B(_0848_),
    .A(\logo_left[8] ),
    .X(_0861_));
 sg13g2_nand3_1 _1828_ (.B(\logo_left[8] ),
    .C(_0848_),
    .A(\logo_left[9] ),
    .Y(_0862_));
 sg13g2_nor4_1 _1829_ (.A(_0850_),
    .B(_0851_),
    .C(_0853_),
    .D(_0858_),
    .Y(_0863_));
 sg13g2_and2_1 _1830_ (.A(_0860_),
    .B(_0862_),
    .X(_0864_));
 sg13g2_nand3b_1 _1831_ (.B(_0863_),
    .C(_0864_),
    .Y(_0865_),
    .A_N(_0861_));
 sg13g2_nor2b_1 _1832_ (.A(_0843_),
    .B_N(_0865_),
    .Y(_0866_));
 sg13g2_a21oi_2 _1833_ (.B1(_0789_),
    .Y(_0867_),
    .A2(_0866_),
    .A1(_0821_));
 sg13g2_xnor2_1 _1834_ (.Y(_0868_),
    .A(net136),
    .B(net612));
 sg13g2_and2_1 _1835_ (.A(net810),
    .B(_0868_),
    .X(_0869_));
 sg13g2_nand2_1 _1836_ (.Y(_0870_),
    .A(net213),
    .B(\color_index[0] ));
 sg13g2_xor2_1 _1837_ (.B(_0870_),
    .A(_0015_),
    .X(_0871_));
 sg13g2_nand2_1 _1838_ (.Y(_0872_),
    .A(net612),
    .B(_0871_));
 sg13g2_o21ai_1 _1839_ (.B1(_0872_),
    .Y(_0873_),
    .A1(net226),
    .A2(net612));
 sg13g2_or2_1 _1840_ (.X(_0874_),
    .B(_0867_),
    .A(net251));
 sg13g2_nor2_1 _1841_ (.A(\color_index[1] ),
    .B(\color_index[0] ),
    .Y(_0875_));
 sg13g2_nand2_1 _1842_ (.Y(_0876_),
    .A(net612),
    .B(_0870_));
 sg13g2_o21ai_1 _1843_ (.B1(_0874_),
    .Y(_0877_),
    .A1(_0875_),
    .A2(_0876_));
 sg13g2_nand2_1 _1844_ (.Y(_0878_),
    .A(_0873_),
    .B(_0877_));
 sg13g2_nand2_1 _1845_ (.Y(_0000_),
    .A(_0869_),
    .B(_0878_));
 sg13g2_nand2_1 _1846_ (.Y(_0879_),
    .A(_0869_),
    .B(_0873_));
 sg13g2_nand2_1 _1847_ (.Y(_0880_),
    .A(net810),
    .B(_0877_));
 sg13g2_mux2_1 _1848_ (.A0(_0877_),
    .A1(_0880_),
    .S(_0879_),
    .X(_0001_));
 sg13g2_nor2_1 _1849_ (.A(_0873_),
    .B(_0880_),
    .Y(_0881_));
 sg13g2_nor2_1 _1850_ (.A(_0869_),
    .B(_0881_),
    .Y(_0882_));
 sg13g2_a21oi_1 _1851_ (.A1(_0868_),
    .A2(_0881_),
    .Y(_0002_),
    .B1(_0882_));
 sg13g2_a21o_1 _1852_ (.A2(_0873_),
    .A1(net810),
    .B1(_0869_),
    .X(_0115_));
 sg13g2_nand2_1 _1853_ (.Y(_0883_),
    .A(_0879_),
    .B(_0115_));
 sg13g2_or2_1 _1854_ (.X(_0003_),
    .B(_0883_),
    .A(_0881_));
 sg13g2_nand2b_1 _1855_ (.Y(_0884_),
    .B(net802),
    .A_N(\pix_x[0] ));
 sg13g2_nor2b_1 _1856_ (.A(net801),
    .B_N(\pix_x[1] ),
    .Y(_0885_));
 sg13g2_xnor2_1 _1857_ (.Y(_0886_),
    .A(net801),
    .B(\pix_x[1] ));
 sg13g2_xor2_1 _1858_ (.B(_0886_),
    .A(_0884_),
    .X(_0887_));
 sg13g2_xor2_1 _1859_ (.B(\pix_y[6] ),
    .A(\logo_top[6] ),
    .X(_0888_));
 sg13g2_nand2_1 _1860_ (.Y(_0889_),
    .A(\logo_top[5] ),
    .B(_0741_));
 sg13g2_nor2_1 _1861_ (.A(net793),
    .B(_0741_),
    .Y(_0890_));
 sg13g2_nand2b_1 _1862_ (.Y(_0891_),
    .B(net778),
    .A_N(\logo_top[4] ));
 sg13g2_xor2_1 _1863_ (.B(net779),
    .A(\logo_top[3] ),
    .X(_0892_));
 sg13g2_nor2b_1 _1864_ (.A(\logo_top[2] ),
    .B_N(net780),
    .Y(_0893_));
 sg13g2_nand2b_1 _1865_ (.Y(_0894_),
    .B(net781),
    .A_N(\logo_top[1] ));
 sg13g2_nor2b_2 _1866_ (.A(\pix_y[0] ),
    .B_N(\logo_top[0] ),
    .Y(_0895_));
 sg13g2_nor2b_1 _1867_ (.A(net781),
    .B_N(net796),
    .Y(_0896_));
 sg13g2_xnor2_1 _1868_ (.Y(_0897_),
    .A(\logo_top[1] ),
    .B(net781));
 sg13g2_o21ai_1 _1869_ (.B1(_0894_),
    .Y(_0898_),
    .A1(_0895_),
    .A2(_0896_));
 sg13g2_xnor2_1 _1870_ (.Y(_0899_),
    .A(net795),
    .B(net780));
 sg13g2_a21oi_2 _1871_ (.B1(_0893_),
    .Y(_0900_),
    .A2(_0899_),
    .A1(_0898_));
 sg13g2_nor2_1 _1872_ (.A(_0892_),
    .B(_0900_),
    .Y(_0901_));
 sg13g2_a21oi_2 _1873_ (.B1(_0901_),
    .Y(_0902_),
    .A2(net779),
    .A1(_0730_));
 sg13g2_nor2b_1 _1874_ (.A(net778),
    .B_N(net794),
    .Y(_0903_));
 sg13g2_xnor2_1 _1875_ (.Y(_0904_),
    .A(net794),
    .B(net778));
 sg13g2_o21ai_1 _1876_ (.B1(_0891_),
    .Y(_0905_),
    .A1(_0902_),
    .A2(_0903_));
 sg13g2_a21o_1 _1877_ (.A2(_0905_),
    .A1(_0889_),
    .B1(_0890_),
    .X(_0906_));
 sg13g2_nand2b_1 _1878_ (.Y(_0907_),
    .B(_0906_),
    .A_N(_0888_));
 sg13g2_xnor2_1 _1879_ (.Y(_0908_),
    .A(_0888_),
    .B(_0906_));
 sg13g2_xor2_1 _1880_ (.B(_0906_),
    .A(_0888_),
    .X(_0909_));
 sg13g2_xnor2_1 _1881_ (.Y(_0910_),
    .A(_0902_),
    .B(_0904_));
 sg13g2_xor2_1 _1882_ (.B(_0904_),
    .A(_0902_),
    .X(_0911_));
 sg13g2_xor2_1 _1883_ (.B(_0900_),
    .A(_0892_),
    .X(_0912_));
 sg13g2_xnor2_1 _1884_ (.Y(_0913_),
    .A(_0892_),
    .B(_0900_));
 sg13g2_xnor2_1 _1885_ (.Y(_0914_),
    .A(_0895_),
    .B(_0897_));
 sg13g2_xor2_1 _1886_ (.B(_0897_),
    .A(_0895_),
    .X(_0915_));
 sg13g2_nand2b_1 _1887_ (.Y(_0916_),
    .B(\logo_left[6] ),
    .A_N(\pix_x[6] ));
 sg13g2_nand2_1 _1888_ (.Y(_0917_),
    .A(_0733_),
    .B(\pix_x[6] ));
 sg13g2_and2_1 _1889_ (.A(_0916_),
    .B(_0917_),
    .X(_0918_));
 sg13g2_nand2_1 _1890_ (.Y(_0919_),
    .A(_0916_),
    .B(_0917_));
 sg13g2_nor2_2 _1891_ (.A(_0734_),
    .B(net803),
    .Y(_0920_));
 sg13g2_nand2b_1 _1892_ (.Y(_0921_),
    .B(\logo_left[5] ),
    .A_N(net803));
 sg13g2_nor2b_1 _1893_ (.A(\logo_left[5] ),
    .B_N(net803),
    .Y(_0922_));
 sg13g2_nor2b_1 _1894_ (.A(\logo_left[4] ),
    .B_N(\pix_x[4] ),
    .Y(_0923_));
 sg13g2_a21oi_2 _1895_ (.B1(_0885_),
    .Y(_0924_),
    .A2(_0886_),
    .A1(_0884_));
 sg13g2_a21o_1 _1896_ (.A2(_0886_),
    .A1(_0884_),
    .B1(_0885_),
    .X(_0925_));
 sg13g2_nor2b_1 _1897_ (.A(\logo_left[2] ),
    .B_N(\pix_x[2] ),
    .Y(_0926_));
 sg13g2_xnor2_1 _1898_ (.Y(_0927_),
    .A(\logo_left[2] ),
    .B(\pix_x[2] ));
 sg13g2_nor2b_1 _1899_ (.A(net800),
    .B_N(\pix_x[3] ),
    .Y(_0928_));
 sg13g2_nand2b_1 _1900_ (.Y(_0929_),
    .B(net800),
    .A_N(\pix_x[3] ));
 sg13g2_xnor2_1 _1901_ (.Y(_0930_),
    .A(net800),
    .B(\pix_x[3] ));
 sg13g2_nand2_1 _1902_ (.Y(_0931_),
    .A(_0927_),
    .B(_0930_));
 sg13g2_a21oi_1 _1903_ (.A1(_0926_),
    .A2(_0929_),
    .Y(_0932_),
    .B1(_0928_));
 sg13g2_o21ai_1 _1904_ (.B1(_0932_),
    .Y(_0933_),
    .A1(_0924_),
    .A2(_0931_));
 sg13g2_xnor2_1 _1905_ (.Y(_0934_),
    .A(net799),
    .B(\pix_x[4] ));
 sg13g2_a21o_1 _1906_ (.A2(_0934_),
    .A1(_0933_),
    .B1(_0923_),
    .X(_0935_));
 sg13g2_a221oi_1 _1907_ (.B2(_0934_),
    .C1(_0923_),
    .B1(_0933_),
    .A1(_0734_),
    .Y(_0936_),
    .A2(net803));
 sg13g2_nor3_2 _1908_ (.A(_0919_),
    .B(_0920_),
    .C(_0936_),
    .Y(_0937_));
 sg13g2_nand3b_1 _1909_ (.B(_0918_),
    .C(_0921_),
    .Y(_0938_),
    .A_N(_0936_));
 sg13g2_a221oi_1 _1910_ (.B2(_0935_),
    .C1(_0922_),
    .B1(_0921_),
    .A1(_0916_),
    .Y(_0939_),
    .A2(_0917_));
 sg13g2_o21ai_1 _1911_ (.B1(_0919_),
    .Y(_0940_),
    .A1(_0920_),
    .A2(_0936_));
 sg13g2_or3_1 _1912_ (.A(_0918_),
    .B(_0920_),
    .C(_0936_),
    .X(_0941_));
 sg13g2_o21ai_1 _1913_ (.B1(_0918_),
    .Y(_0942_),
    .A1(_0920_),
    .A2(_0936_));
 sg13g2_nor2_1 _1914_ (.A(_0937_),
    .B(_0939_),
    .Y(_0943_));
 sg13g2_nand2_1 _1915_ (.Y(_0944_),
    .A(net695),
    .B(net694));
 sg13g2_xor2_1 _1916_ (.B(_0934_),
    .A(_0933_),
    .X(_0945_));
 sg13g2_xnor2_1 _1917_ (.Y(_0946_),
    .A(_0933_),
    .B(_0934_));
 sg13g2_a21oi_1 _1918_ (.A1(_0925_),
    .A2(_0927_),
    .Y(_0947_),
    .B1(_0926_));
 sg13g2_xnor2_1 _1919_ (.Y(_0948_),
    .A(_0930_),
    .B(_0947_));
 sg13g2_xor2_1 _1920_ (.B(_0947_),
    .A(_0930_),
    .X(_0949_));
 sg13g2_nor2_1 _1921_ (.A(net710),
    .B(_0949_),
    .Y(_0950_));
 sg13g2_nand2_2 _1922_ (.Y(_0951_),
    .A(net707),
    .B(_0948_));
 sg13g2_nor2_2 _1923_ (.A(net707),
    .B(_0948_),
    .Y(_0952_));
 sg13g2_nand2_2 _1924_ (.Y(_0953_),
    .A(net709),
    .B(_0949_));
 sg13g2_nor2_1 _1925_ (.A(_0920_),
    .B(_0922_),
    .Y(_0954_));
 sg13g2_xnor2_1 _1926_ (.Y(_0955_),
    .A(_0935_),
    .B(_0954_));
 sg13g2_xor2_1 _1927_ (.B(_0954_),
    .A(_0935_),
    .X(_0956_));
 sg13g2_nand2_1 _1928_ (.Y(_0957_),
    .A(net709),
    .B(net680));
 sg13g2_nor2_2 _1929_ (.A(net711),
    .B(_0948_),
    .Y(_0958_));
 sg13g2_nand2_2 _1930_ (.Y(_0959_),
    .A(net708),
    .B(_0949_));
 sg13g2_nor2_2 _1931_ (.A(net708),
    .B(_0949_),
    .Y(_0960_));
 sg13g2_nand2_2 _1932_ (.Y(_0961_),
    .A(net711),
    .B(_0948_));
 sg13g2_xnor2_1 _1933_ (.Y(_0962_),
    .A(net708),
    .B(_0948_));
 sg13g2_xnor2_1 _1934_ (.Y(_0963_),
    .A(net709),
    .B(_0948_));
 sg13g2_a221oi_1 _1935_ (.B2(net681),
    .C1(_0950_),
    .B1(_0952_),
    .A1(net696),
    .Y(_0964_),
    .A2(net693));
 sg13g2_inv_1 _1936_ (.Y(_0965_),
    .A(_0964_));
 sg13g2_a22oi_1 _1937_ (.Y(_0966_),
    .B1(net710),
    .B2(net680),
    .A2(net689),
    .A1(net691));
 sg13g2_nand2_2 _1938_ (.Y(_0967_),
    .A(net687),
    .B(_0961_));
 sg13g2_nand2_1 _1939_ (.Y(_0968_),
    .A(net686),
    .B(_0962_));
 sg13g2_nand2_1 _1940_ (.Y(_0969_),
    .A(net652),
    .B(net651));
 sg13g2_a21oi_2 _1941_ (.B1(_0964_),
    .Y(_0970_),
    .A2(net651),
    .A1(net654));
 sg13g2_nor2_1 _1942_ (.A(net710),
    .B(net681),
    .Y(_0971_));
 sg13g2_nand2_1 _1943_ (.Y(_0972_),
    .A(net707),
    .B(net685));
 sg13g2_nand2_1 _1944_ (.Y(_0973_),
    .A(net688),
    .B(net685));
 sg13g2_nor2_2 _1945_ (.A(net710),
    .B(net685),
    .Y(_0974_));
 sg13g2_o21ai_1 _1946_ (.B1(net661),
    .Y(_0975_),
    .A1(net677),
    .A2(_0974_));
 sg13g2_xnor2_1 _1947_ (.Y(_0976_),
    .A(net797),
    .B(\pix_y[0] ));
 sg13g2_xor2_1 _1948_ (.B(\pix_y[0] ),
    .A(net797),
    .X(_0977_));
 sg13g2_nand2_2 _1949_ (.Y(_0978_),
    .A(net757),
    .B(net774));
 sg13g2_nor2_1 _1950_ (.A(_0964_),
    .B(_0978_),
    .Y(_0979_));
 sg13g2_nor2_1 _1951_ (.A(net751),
    .B(net773),
    .Y(_0980_));
 sg13g2_nand2_2 _1952_ (.Y(_0981_),
    .A(net753),
    .B(net765));
 sg13g2_nor2_1 _1953_ (.A(net659),
    .B(net707),
    .Y(_0982_));
 sg13g2_nand3_1 _1954_ (.B(net693),
    .C(_0952_),
    .A(net696),
    .Y(_0983_));
 sg13g2_nand2_1 _1955_ (.Y(_0984_),
    .A(net646),
    .B(_0983_));
 sg13g2_a21oi_1 _1956_ (.A1(net646),
    .A2(_0983_),
    .Y(_0985_),
    .B1(net742));
 sg13g2_a221oi_1 _1957_ (.B2(_0979_),
    .C1(_0985_),
    .B1(_0975_),
    .A1(net749),
    .Y(_0986_),
    .A2(_0970_));
 sg13g2_xor2_1 _1958_ (.B(_0899_),
    .A(_0898_),
    .X(_0987_));
 sg13g2_xnor2_1 _1959_ (.Y(_0988_),
    .A(_0898_),
    .B(_0899_));
 sg13g2_nor2_2 _1960_ (.A(net756),
    .B(net774),
    .Y(_0989_));
 sg13g2_nand2_2 _1961_ (.Y(_0990_),
    .A(net748),
    .B(net765));
 sg13g2_o21ai_1 _1962_ (.B1(net741),
    .Y(_0991_),
    .A1(_0975_),
    .A2(_0990_));
 sg13g2_nor2_2 _1963_ (.A(net748),
    .B(net737),
    .Y(_0992_));
 sg13g2_nand2_2 _1964_ (.Y(_0993_),
    .A(net752),
    .B(net728));
 sg13g2_nand2_1 _1965_ (.Y(_0994_),
    .A(_0970_),
    .B(net706));
 sg13g2_o21ai_1 _1966_ (.B1(_0994_),
    .Y(_0995_),
    .A1(_0986_),
    .A2(_0991_));
 sg13g2_a22oi_1 _1967_ (.Y(_0996_),
    .B1(net686),
    .B2(_0962_),
    .A2(net693),
    .A1(net696));
 sg13g2_nand2_2 _1968_ (.Y(_0997_),
    .A(net659),
    .B(net650));
 sg13g2_a21oi_1 _1969_ (.A1(net659),
    .A2(net681),
    .Y(_0998_),
    .B1(net677));
 sg13g2_o21ai_1 _1970_ (.B1(_0962_),
    .Y(_0999_),
    .A1(net661),
    .A2(net685));
 sg13g2_nand2_1 _1971_ (.Y(_1000_),
    .A(net651),
    .B(_0983_));
 sg13g2_nor2_1 _1972_ (.A(net767),
    .B(_1000_),
    .Y(_1001_));
 sg13g2_a21oi_1 _1973_ (.A1(net767),
    .A2(_0999_),
    .Y(_1002_),
    .B1(_1001_));
 sg13g2_nor2_2 _1974_ (.A(net752),
    .B(net730),
    .Y(_1003_));
 sg13g2_nand2_2 _1975_ (.Y(_1004_),
    .A(net748),
    .B(net737));
 sg13g2_nor2_1 _1976_ (.A(net715),
    .B(_1004_),
    .Y(_1005_));
 sg13g2_nor2_2 _1977_ (.A(net683),
    .B(_0958_),
    .Y(_1006_));
 sg13g2_nand2_1 _1978_ (.Y(_1007_),
    .A(net678),
    .B(_0959_));
 sg13g2_nand2_2 _1979_ (.Y(_1008_),
    .A(net681),
    .B(_0962_));
 sg13g2_a22oi_1 _1980_ (.Y(_1009_),
    .B1(net681),
    .B2(_0962_),
    .A2(net693),
    .A1(net696));
 sg13g2_nand2_2 _1981_ (.Y(_1010_),
    .A(net648),
    .B(net645));
 sg13g2_a22oi_1 _1982_ (.Y(_1011_),
    .B1(net649),
    .B2(net645),
    .A2(net651),
    .A1(net654));
 sg13g2_nor2_2 _1983_ (.A(net753),
    .B(net737),
    .Y(_1012_));
 sg13g2_nand2_1 _1984_ (.Y(_1013_),
    .A(net751),
    .B(net733));
 sg13g2_nor2_2 _1985_ (.A(net723),
    .B(net701),
    .Y(_1014_));
 sg13g2_nand2_1 _1986_ (.Y(_1015_),
    .A(_1011_),
    .B(_1014_));
 sg13g2_nor2_2 _1987_ (.A(net713),
    .B(net737),
    .Y(_1016_));
 sg13g2_nand2_2 _1988_ (.Y(_1017_),
    .A(net723),
    .B(net733));
 sg13g2_nor2_1 _1989_ (.A(net748),
    .B(net728),
    .Y(_1018_));
 sg13g2_nand2_2 _1990_ (.Y(_1019_),
    .A(net757),
    .B(net741));
 sg13g2_nor2_1 _1991_ (.A(net718),
    .B(net732),
    .Y(_1020_));
 sg13g2_nand2_2 _1992_ (.Y(_1021_),
    .A(net723),
    .B(net741));
 sg13g2_nor2_2 _1993_ (.A(net715),
    .B(_1019_),
    .Y(_1022_));
 sg13g2_nand2_2 _1994_ (.Y(_1023_),
    .A(net725),
    .B(net699));
 sg13g2_a22oi_1 _1995_ (.Y(_1024_),
    .B1(_1022_),
    .B2(_0998_),
    .A2(_1016_),
    .A1(_0984_));
 sg13g2_nand2_1 _1996_ (.Y(_1025_),
    .A(_1015_),
    .B(_1024_));
 sg13g2_a221oi_1 _1997_ (.B2(_1005_),
    .C1(_1025_),
    .B1(_1002_),
    .A1(net715),
    .Y(_1026_),
    .A2(_0995_));
 sg13g2_xnor2_1 _1998_ (.Y(_1027_),
    .A(net793),
    .B(\pix_y[5] ));
 sg13g2_xnor2_1 _1999_ (.Y(_1028_),
    .A(_0905_),
    .B(_1027_));
 sg13g2_xor2_1 _2000_ (.B(_1027_),
    .A(_0905_),
    .X(_1029_));
 sg13g2_nand2_2 _2001_ (.Y(_1030_),
    .A(net678),
    .B(_0958_));
 sg13g2_inv_1 _2002_ (.Y(_1031_),
    .A(_1030_));
 sg13g2_mux2_2 _2003_ (.A0(net708),
    .A1(_0959_),
    .S(net678),
    .X(_1032_));
 sg13g2_mux2_2 _2004_ (.A0(net711),
    .A1(_0958_),
    .S(net678),
    .X(_1033_));
 sg13g2_nand2_2 _2005_ (.Y(_1034_),
    .A(net657),
    .B(_1032_));
 sg13g2_a22oi_1 _2006_ (.Y(_1035_),
    .B1(net680),
    .B2(_0962_),
    .A2(net689),
    .A1(net691));
 sg13g2_nor3_2 _2007_ (.A(_0937_),
    .B(_0939_),
    .C(net683),
    .Y(_1036_));
 sg13g2_nand3_1 _2008_ (.B(net694),
    .C(net679),
    .A(net695),
    .Y(_1037_));
 sg13g2_nor4_2 _2009_ (.A(_0937_),
    .B(_0939_),
    .C(net685),
    .Y(_1038_),
    .D(net677));
 sg13g2_nand4_1 _2010_ (.B(net693),
    .C(net681),
    .A(net697),
    .Y(_1039_),
    .D(_0962_));
 sg13g2_a22oi_1 _2011_ (.Y(_1040_),
    .B1(net679),
    .B2(_0959_),
    .A2(net694),
    .A1(net695));
 sg13g2_a21oi_2 _2012_ (.B1(_1038_),
    .Y(_1041_),
    .A2(net642),
    .A1(net648));
 sg13g2_nor2_1 _2013_ (.A(net722),
    .B(net705),
    .Y(_1042_));
 sg13g2_nand2_1 _2014_ (.Y(_1043_),
    .A(net683),
    .B(_0958_));
 sg13g2_inv_1 _2015_ (.Y(_1044_),
    .A(net639));
 sg13g2_a21o_1 _2016_ (.A2(net639),
    .A1(net642),
    .B1(_1038_),
    .X(_1045_));
 sg13g2_a21oi_1 _2017_ (.A1(net705),
    .A2(_1045_),
    .Y(_1046_),
    .B1(net722));
 sg13g2_a22oi_1 _2018_ (.Y(_1047_),
    .B1(net688),
    .B2(_0956_),
    .A2(net689),
    .A1(net691));
 sg13g2_o21ai_1 _2019_ (.B1(net661),
    .Y(_1048_),
    .A1(_0951_),
    .A2(net685));
 sg13g2_a221oi_1 _2020_ (.B2(_1034_),
    .C1(_1017_),
    .B1(_1048_),
    .A1(net750),
    .Y(_1049_),
    .A2(_1038_));
 sg13g2_a221oi_1 _2021_ (.B2(_1046_),
    .C1(_1049_),
    .B1(_1041_),
    .A1(_1011_),
    .Y(_1050_),
    .A2(net675));
 sg13g2_mux2_1 _2022_ (.A0(_1026_),
    .A1(_1050_),
    .S(net664),
    .X(_1051_));
 sg13g2_a22oi_1 _2023_ (.Y(_1052_),
    .B1(net710),
    .B2(net686),
    .A2(net693),
    .A1(net696));
 sg13g2_a22oi_1 _2024_ (.Y(_1053_),
    .B1(net708),
    .B2(net680),
    .A2(net689),
    .A1(net691));
 sg13g2_nand2b_1 _2025_ (.Y(_1054_),
    .B(net661),
    .A_N(_0974_));
 sg13g2_nand2_1 _2026_ (.Y(_1055_),
    .A(net650),
    .B(net635));
 sg13g2_a21o_1 _2027_ (.A2(net635),
    .A1(net650),
    .B1(net637),
    .X(_1056_));
 sg13g2_a21oi_2 _2028_ (.B1(net679),
    .Y(_1057_),
    .A2(net694),
    .A1(net695));
 sg13g2_o21ai_1 _2029_ (.B1(net683),
    .Y(_1058_),
    .A1(_0937_),
    .A2(_0939_));
 sg13g2_nor2_1 _2030_ (.A(_0953_),
    .B(net680),
    .Y(_1059_));
 sg13g2_a22oi_1 _2031_ (.Y(_1060_),
    .B1(_0952_),
    .B2(net686),
    .A2(_0940_),
    .A1(net696));
 sg13g2_a21oi_1 _2032_ (.A1(net660),
    .A2(net688),
    .Y(_1061_),
    .B1(_1059_));
 sg13g2_a221oi_1 _2033_ (.B2(net709),
    .C1(_1059_),
    .B1(_1057_),
    .A1(net660),
    .Y(_1062_),
    .A2(net688));
 sg13g2_mux2_1 _2034_ (.A0(_1056_),
    .A1(_1062_),
    .S(net771),
    .X(_1063_));
 sg13g2_nor2_1 _2035_ (.A(net676),
    .B(net638),
    .Y(_1064_));
 sg13g2_nor2_2 _2036_ (.A(net752),
    .B(net763),
    .Y(_1065_));
 sg13g2_nand2_2 _2037_ (.Y(_1066_),
    .A(_0897_),
    .B(net773));
 sg13g2_o21ai_1 _2038_ (.B1(net738),
    .Y(_1067_),
    .A1(_1064_),
    .A2(_1066_));
 sg13g2_a221oi_1 _2039_ (.B2(net754),
    .C1(_1067_),
    .B1(_1063_),
    .A1(_0989_),
    .Y(_1068_),
    .A2(_1061_));
 sg13g2_a221oi_1 _2040_ (.B2(net755),
    .C1(net676),
    .B1(net638),
    .A1(net657),
    .Y(_1069_),
    .A2(net680));
 sg13g2_nand2_1 _2041_ (.Y(_1070_),
    .A(net731),
    .B(_1069_));
 sg13g2_nand2_2 _2042_ (.Y(_1071_),
    .A(net774),
    .B(net733));
 sg13g2_o21ai_1 _2043_ (.B1(_1070_),
    .Y(_1072_),
    .A1(_0999_),
    .A2(_1071_));
 sg13g2_o21ai_1 _2044_ (.B1(net715),
    .Y(_1073_),
    .A1(_1068_),
    .A2(_1072_));
 sg13g2_mux2_1 _2045_ (.A0(_0959_),
    .A1(_0961_),
    .S(net683),
    .X(_1074_));
 sg13g2_and3_1 _2046_ (.X(_1075_),
    .A(net655),
    .B(net763),
    .C(net630));
 sg13g2_nand3_1 _2047_ (.B(net766),
    .C(net631),
    .A(net657),
    .Y(_1076_));
 sg13g2_a22oi_1 _2048_ (.Y(_1077_),
    .B1(net635),
    .B2(net650),
    .A2(_1032_),
    .A1(net657));
 sg13g2_a21oi_1 _2049_ (.A1(_1076_),
    .A2(_1077_),
    .Y(_1078_),
    .B1(_1004_));
 sg13g2_and2_1 _2050_ (.A(net731),
    .B(_1056_),
    .X(_1079_));
 sg13g2_nand4_1 _2051_ (.B(net693),
    .C(net687),
    .A(net696),
    .Y(_1080_),
    .D(net676));
 sg13g2_a21oi_1 _2052_ (.A1(net656),
    .A2(net630),
    .Y(_1081_),
    .B1(_1006_));
 sg13g2_o21ai_1 _2053_ (.B1(_1007_),
    .Y(_1082_),
    .A1(net660),
    .A2(_0967_));
 sg13g2_a21oi_1 _2054_ (.A1(_1080_),
    .A2(_1081_),
    .Y(_1083_),
    .B1(_1019_));
 sg13g2_nor4_1 _2055_ (.A(net713),
    .B(_1078_),
    .C(_1079_),
    .D(_1083_),
    .Y(_1084_));
 sg13g2_nor2_1 _2056_ (.A(net667),
    .B(_1084_),
    .Y(_1085_));
 sg13g2_mux2_2 _2057_ (.A0(net711),
    .A1(_0961_),
    .S(net683),
    .X(_1086_));
 sg13g2_and2_1 _2058_ (.A(net655),
    .B(_1086_),
    .X(_1087_));
 sg13g2_nand2_1 _2059_ (.Y(_1088_),
    .A(net656),
    .B(_1086_));
 sg13g2_nand4_1 _2060_ (.B(net694),
    .C(net679),
    .A(net695),
    .Y(_1089_),
    .D(_0959_));
 sg13g2_mux2_1 _2061_ (.A0(_1006_),
    .A1(_1086_),
    .S(net656),
    .X(_1090_));
 sg13g2_nand2_1 _2062_ (.Y(_1091_),
    .A(_1080_),
    .B(_1089_));
 sg13g2_nor2_2 _2063_ (.A(net743),
    .B(net736),
    .Y(_1092_));
 sg13g2_o21ai_1 _2064_ (.B1(_1092_),
    .Y(_1093_),
    .A1(_1087_),
    .A2(_1091_));
 sg13g2_a22oi_1 _2065_ (.Y(_1094_),
    .B1(net683),
    .B2(_0961_),
    .A2(net690),
    .A1(net692));
 sg13g2_or2_2 _2066_ (.X(_1095_),
    .B(_1094_),
    .A(_1057_));
 sg13g2_nand2_1 _2067_ (.Y(_1096_),
    .A(net736),
    .B(_1095_));
 sg13g2_nand2_1 _2068_ (.Y(_1097_),
    .A(net682),
    .B(_0960_));
 sg13g2_xnor2_1 _2069_ (.Y(_1098_),
    .A(net678),
    .B(_0960_));
 sg13g2_and2_2 _2070_ (.A(net655),
    .B(_1098_),
    .X(_1099_));
 sg13g2_o21ai_1 _2071_ (.B1(net728),
    .Y(_1100_),
    .A1(_1091_),
    .A2(_1099_));
 sg13g2_nand4_1 _2072_ (.B(_1093_),
    .C(_1096_),
    .A(net714),
    .Y(_1101_),
    .D(_1100_));
 sg13g2_nor2_2 _2073_ (.A(_1036_),
    .B(_1057_),
    .Y(_1102_));
 sg13g2_and2_1 _2074_ (.A(net630),
    .B(_1102_),
    .X(_1103_));
 sg13g2_nand3_1 _2075_ (.B(net632),
    .C(net630),
    .A(net643),
    .Y(_1104_));
 sg13g2_a22oi_1 _2076_ (.Y(_1105_),
    .B1(net707),
    .B2(net684),
    .A2(net690),
    .A1(net692));
 sg13g2_a22oi_1 _2077_ (.Y(_1106_),
    .B1(net711),
    .B2(net679),
    .A2(net694),
    .A1(net695));
 sg13g2_or2_1 _2078_ (.X(_1107_),
    .B(_1106_),
    .A(net628));
 sg13g2_a22oi_1 _2079_ (.Y(_1108_),
    .B1(net682),
    .B2(_0960_),
    .A2(net694),
    .A1(net695));
 sg13g2_or3_1 _2080_ (.A(_0977_),
    .B(net628),
    .C(_1108_),
    .X(_1109_));
 sg13g2_nor3_2 _2081_ (.A(_0937_),
    .B(_0939_),
    .C(_0949_),
    .Y(_1110_));
 sg13g2_or4_1 _2082_ (.A(net764),
    .B(net628),
    .C(_1108_),
    .D(net627),
    .X(_1111_));
 sg13g2_a22oi_1 _2083_ (.Y(_1112_),
    .B1(_1111_),
    .B2(net699),
    .A2(_1107_),
    .A1(net739));
 sg13g2_nand3_1 _2084_ (.B(_1103_),
    .C(_1112_),
    .A(net720),
    .Y(_1113_));
 sg13g2_and3_1 _2085_ (.X(_1114_),
    .A(net668),
    .B(_1101_),
    .C(_1113_));
 sg13g2_a21o_1 _2086_ (.A2(_1085_),
    .A1(_1073_),
    .B1(_1114_),
    .X(_1115_));
 sg13g2_mux2_1 _2087_ (.A0(_1051_),
    .A1(_1115_),
    .S(_1029_),
    .X(_1116_));
 sg13g2_xnor2_1 _2088_ (.Y(_1117_),
    .A(\logo_left[0] ),
    .B(\pix_x[0] ));
 sg13g2_xor2_1 _2089_ (.B(\pix_x[0] ),
    .A(net802),
    .X(_1118_));
 sg13g2_nor2_1 _2090_ (.A(net770),
    .B(net628),
    .Y(_1119_));
 sg13g2_or3_1 _2091_ (.A(net773),
    .B(net629),
    .C(_1108_),
    .X(_1120_));
 sg13g2_or4_1 _2092_ (.A(net773),
    .B(net629),
    .C(_1108_),
    .D(net627),
    .X(_1121_));
 sg13g2_nand2_1 _2093_ (.Y(_1122_),
    .A(net704),
    .B(_1121_));
 sg13g2_a22oi_1 _2094_ (.Y(_1123_),
    .B1(_1121_),
    .B2(net704),
    .A2(_1107_),
    .A1(net732));
 sg13g2_nand2_1 _2095_ (.Y(_1124_),
    .A(_0981_),
    .B(_1104_));
 sg13g2_nor2_1 _2096_ (.A(_1036_),
    .B(net641),
    .Y(_1125_));
 sg13g2_or2_1 _2097_ (.X(_1126_),
    .B(net641),
    .A(_1036_));
 sg13g2_nand4_1 _2098_ (.B(_1123_),
    .C(_1124_),
    .A(net716),
    .Y(_1127_),
    .D(_1125_));
 sg13g2_nand2_1 _2099_ (.Y(_1128_),
    .A(net732),
    .B(_1102_));
 sg13g2_and2_1 _2100_ (.A(net662),
    .B(net630),
    .X(_1129_));
 sg13g2_nand2_1 _2101_ (.Y(_1130_),
    .A(net660),
    .B(net631));
 sg13g2_nor2_1 _2102_ (.A(net658),
    .B(_1033_),
    .Y(_1131_));
 sg13g2_mux2_2 _2103_ (.A0(_1032_),
    .A1(_1086_),
    .S(net655),
    .X(_1132_));
 sg13g2_a221oi_1 _2104_ (.B2(net752),
    .C1(net728),
    .B1(_1132_),
    .A1(net743),
    .Y(_1133_),
    .A2(_1129_));
 sg13g2_a21oi_2 _2105_ (.B1(net655),
    .Y(_1134_),
    .A2(_0959_),
    .A1(net683));
 sg13g2_a221oi_1 _2106_ (.B2(_1030_),
    .C1(_1099_),
    .B1(_1134_),
    .A1(net763),
    .Y(_1135_),
    .A2(_1132_));
 sg13g2_a22oi_1 _2107_ (.Y(_1136_),
    .B1(_1133_),
    .B2(_1135_),
    .A2(_1102_),
    .A1(net729));
 sg13g2_o21ai_1 _2108_ (.B1(_1127_),
    .Y(_1137_),
    .A1(net715),
    .A2(_1136_));
 sg13g2_and4_1 _2109_ (.A(net691),
    .B(net689),
    .C(net707),
    .D(net685),
    .X(_1138_));
 sg13g2_a21o_2 _2110_ (.A2(net629),
    .A1(_1008_),
    .B1(_1138_),
    .X(_1139_));
 sg13g2_and2_1 _2111_ (.A(net738),
    .B(_1139_),
    .X(_1140_));
 sg13g2_o21ai_1 _2112_ (.B1(_1140_),
    .Y(_1141_),
    .A1(net646),
    .A2(net727));
 sg13g2_or2_2 _2113_ (.X(_1142_),
    .B(net634),
    .A(net637));
 sg13g2_nor2_1 _2114_ (.A(net716),
    .B(net750),
    .Y(_1143_));
 sg13g2_nand2_2 _2115_ (.Y(_1144_),
    .A(net722),
    .B(net701));
 sg13g2_a21oi_1 _2116_ (.A1(net702),
    .A2(_1142_),
    .Y(_1145_),
    .B1(net714));
 sg13g2_nor2_2 _2117_ (.A(_0978_),
    .B(net739),
    .Y(_1146_));
 sg13g2_nor4_2 _2118_ (.A(_0937_),
    .B(_0939_),
    .C(_0951_),
    .Y(_1147_),
    .D(net685));
 sg13g2_or2_1 _2119_ (.X(_1148_),
    .B(net638),
    .A(_1047_));
 sg13g2_a22oi_1 _2120_ (.Y(_1149_),
    .B1(_1146_),
    .B2(_1148_),
    .A2(_1139_),
    .A1(net706));
 sg13g2_nand3_1 _2121_ (.B(_1145_),
    .C(_1149_),
    .A(_1141_),
    .Y(_1150_));
 sg13g2_a221oi_1 _2122_ (.B2(net738),
    .C1(net721),
    .B1(_1142_),
    .A1(net702),
    .Y(_1151_),
    .A2(net631));
 sg13g2_or2_1 _2123_ (.X(_1152_),
    .B(net641),
    .A(net652));
 sg13g2_o21ai_1 _2124_ (.B1(_0967_),
    .Y(_1153_),
    .A1(net654),
    .A2(net641));
 sg13g2_nor2_2 _2125_ (.A(net742),
    .B(net736),
    .Y(_1154_));
 sg13g2_nand2_2 _2126_ (.Y(_1155_),
    .A(net743),
    .B(net728));
 sg13g2_nand2_1 _2127_ (.Y(_1156_),
    .A(_1034_),
    .B(_1054_));
 sg13g2_a22oi_1 _2128_ (.Y(_1157_),
    .B1(_1154_),
    .B2(_1156_),
    .A2(_1153_),
    .A1(_1146_));
 sg13g2_a21oi_1 _2129_ (.A1(_1151_),
    .A2(_1157_),
    .Y(_1158_),
    .B1(net664));
 sg13g2_a21oi_1 _2130_ (.A1(_1150_),
    .A2(_1158_),
    .Y(_1159_),
    .B1(net622));
 sg13g2_o21ai_1 _2131_ (.B1(_1159_),
    .Y(_1160_),
    .A1(net667),
    .A2(_1137_));
 sg13g2_nand3_1 _2132_ (.B(net646),
    .C(_1139_),
    .A(net750),
    .Y(_1161_));
 sg13g2_and4_2 _2133_ (.A(net691),
    .B(net689),
    .C(net684),
    .D(_0958_),
    .X(_1162_));
 sg13g2_nand2b_2 _2134_ (.Y(_1163_),
    .B(net658),
    .A_N(net640));
 sg13g2_a22oi_1 _2135_ (.Y(_1164_),
    .B1(_0952_),
    .B2(net681),
    .A2(net689),
    .A1(net691));
 sg13g2_nor2_1 _2136_ (.A(net653),
    .B(_1110_),
    .Y(_1165_));
 sg13g2_nand2_1 _2137_ (.Y(_1166_),
    .A(net648),
    .B(_1164_));
 sg13g2_a21oi_1 _2138_ (.A1(net648),
    .A2(_1164_),
    .Y(_1167_),
    .B1(_1162_));
 sg13g2_a21o_1 _2139_ (.A2(_1164_),
    .A1(net647),
    .B1(_1162_),
    .X(_1168_));
 sg13g2_o21ai_1 _2140_ (.B1(_1092_),
    .Y(_1169_),
    .A1(net688),
    .A2(net705));
 sg13g2_a21oi_1 _2141_ (.A1(_1168_),
    .A2(_1169_),
    .Y(_1170_),
    .B1(net724));
 sg13g2_nor2_2 _2142_ (.A(net730),
    .B(net727),
    .Y(_1171_));
 sg13g2_nor2_1 _2143_ (.A(net653),
    .B(net644),
    .Y(_1172_));
 sg13g2_or2_1 _2144_ (.X(_1173_),
    .B(net645),
    .A(net652));
 sg13g2_a21oi_1 _2145_ (.A1(_1171_),
    .A2(_1173_),
    .Y(_1174_),
    .B1(net717));
 sg13g2_a21o_2 _2146_ (.A2(net648),
    .A1(net652),
    .B1(_1162_),
    .X(_1175_));
 sg13g2_inv_1 _2147_ (.Y(_1176_),
    .A(_1175_));
 sg13g2_nand2_1 _2148_ (.Y(_1177_),
    .A(_1092_),
    .B(_1168_));
 sg13g2_a221oi_1 _2149_ (.B2(_1071_),
    .C1(net719),
    .B1(_1175_),
    .A1(_1171_),
    .Y(_1178_),
    .A2(_1173_));
 sg13g2_a221oi_1 _2150_ (.B2(_1178_),
    .C1(net669),
    .B1(_1177_),
    .A1(_1161_),
    .Y(_1179_),
    .A2(_1170_));
 sg13g2_and2_1 _2151_ (.A(net722),
    .B(_1041_),
    .X(_1180_));
 sg13g2_a22oi_1 _2152_ (.Y(_1181_),
    .B1(net682),
    .B2(_0960_),
    .A2(net689),
    .A1(net691));
 sg13g2_a21oi_1 _2153_ (.A1(net648),
    .A2(net644),
    .Y(_1182_),
    .B1(_1181_));
 sg13g2_o21ai_1 _2154_ (.B1(_1180_),
    .Y(_1183_),
    .A1(net701),
    .A2(_1182_));
 sg13g2_nor2_1 _2155_ (.A(_1004_),
    .B(_1041_),
    .Y(_1184_));
 sg13g2_a221oi_1 _2156_ (.B2(net673),
    .C1(_1184_),
    .B1(_1183_),
    .A1(_1045_),
    .Y(_1185_),
    .A2(_1171_));
 sg13g2_a21oi_1 _2157_ (.A1(net644),
    .A2(net705),
    .Y(_1186_),
    .B1(net653));
 sg13g2_and3_1 _2158_ (.X(_1187_),
    .A(net717),
    .B(_1010_),
    .C(_1186_));
 sg13g2_nand2_1 _2159_ (.Y(_1188_),
    .A(net699),
    .B(net626));
 sg13g2_a21oi_1 _2160_ (.A1(_1187_),
    .A2(_1188_),
    .Y(_1189_),
    .B1(net665));
 sg13g2_nand2b_1 _2161_ (.Y(_1190_),
    .B(_1189_),
    .A_N(_1185_));
 sg13g2_nor2_1 _2162_ (.A(net624),
    .B(_1179_),
    .Y(_1191_));
 sg13g2_a21oi_1 _2163_ (.A1(_1190_),
    .A2(_1191_),
    .Y(_1192_),
    .B1(net620));
 sg13g2_a221oi_1 _2164_ (.B2(_1192_),
    .C1(_1117_),
    .B1(_1160_),
    .A1(net620),
    .Y(_1193_),
    .A2(_1116_));
 sg13g2_nand2_1 _2165_ (.Y(_1194_),
    .A(_0989_),
    .B(_1132_));
 sg13g2_o21ai_1 _2166_ (.B1(net748),
    .Y(_1195_),
    .A1(net769),
    .A2(_1132_));
 sg13g2_a22oi_1 _2167_ (.Y(_1196_),
    .B1(net679),
    .B2(_0961_),
    .A2(net694),
    .A1(net695));
 sg13g2_a221oi_1 _2168_ (.B2(_1030_),
    .C1(_1196_),
    .B1(_1134_),
    .A1(net763),
    .Y(_1197_),
    .A2(_1132_));
 sg13g2_o21ai_1 _2169_ (.B1(_1133_),
    .Y(_1198_),
    .A1(_1195_),
    .A2(_1197_));
 sg13g2_nand2_1 _2170_ (.Y(_1199_),
    .A(net633),
    .B(_1089_));
 sg13g2_nor2_1 _2171_ (.A(net740),
    .B(_1199_),
    .Y(_1200_));
 sg13g2_o21ai_1 _2172_ (.B1(_1200_),
    .Y(_1201_),
    .A1(net743),
    .A2(_1102_));
 sg13g2_or2_1 _2173_ (.X(_1202_),
    .B(_1106_),
    .A(_1094_));
 sg13g2_a221oi_1 _2174_ (.B2(_1065_),
    .C1(_1126_),
    .B1(_1202_),
    .A1(_0989_),
    .Y(_1203_),
    .A2(_1104_));
 sg13g2_nand2_1 _2175_ (.Y(_1204_),
    .A(net773),
    .B(_1104_));
 sg13g2_nand4_1 _2176_ (.B(_1123_),
    .C(_1203_),
    .A(net716),
    .Y(_1205_),
    .D(_1204_));
 sg13g2_a21o_1 _2177_ (.A2(_1201_),
    .A1(_1198_),
    .B1(net716),
    .X(_1206_));
 sg13g2_nand3_1 _2178_ (.B(_1205_),
    .C(_1206_),
    .A(net666),
    .Y(_1207_));
 sg13g2_or2_1 _2179_ (.X(_1208_),
    .B(_1052_),
    .A(_1035_));
 sg13g2_a221oi_1 _2180_ (.B2(_1208_),
    .C1(net714),
    .B1(_1146_),
    .A1(net706),
    .Y(_1209_),
    .A2(_1139_));
 sg13g2_nand3_1 _2181_ (.B(net688),
    .C(net687),
    .A(net754),
    .Y(_1210_));
 sg13g2_nand3_1 _2182_ (.B(_1139_),
    .C(_1210_),
    .A(net738),
    .Y(_1211_));
 sg13g2_nor2_2 _2183_ (.A(net739),
    .B(_1066_),
    .Y(_1212_));
 sg13g2_nand2_2 _2184_ (.Y(_1213_),
    .A(net733),
    .B(net727));
 sg13g2_nor2_2 _2185_ (.A(net738),
    .B(_0990_),
    .Y(_1214_));
 sg13g2_a22oi_1 _2186_ (.Y(_1215_),
    .B1(_1214_),
    .B2(_1148_),
    .A2(_1212_),
    .A1(_1142_));
 sg13g2_nand3_1 _2187_ (.B(_1211_),
    .C(_1215_),
    .A(_1209_),
    .Y(_1216_));
 sg13g2_and2_1 _2188_ (.A(net769),
    .B(net631),
    .X(_1217_));
 sg13g2_a21o_1 _2189_ (.A2(_1153_),
    .A1(net765),
    .B1(_1217_),
    .X(_1218_));
 sg13g2_and2_1 _2190_ (.A(_1142_),
    .B(_1171_),
    .X(_1219_));
 sg13g2_a21oi_1 _2191_ (.A1(net657),
    .A2(net631),
    .Y(_1220_),
    .B1(net634));
 sg13g2_a21o_1 _2192_ (.A2(net631),
    .A1(net657),
    .B1(net634),
    .X(_1221_));
 sg13g2_nand2_1 _2193_ (.Y(_1222_),
    .A(_1154_),
    .B(_1221_));
 sg13g2_a221oi_1 _2194_ (.B2(_1142_),
    .C1(net721),
    .B1(_1171_),
    .A1(net738),
    .Y(_1223_),
    .A2(_1156_));
 sg13g2_a22oi_1 _2195_ (.Y(_1224_),
    .B1(_1218_),
    .B2(net702),
    .A2(_1153_),
    .A1(_1146_));
 sg13g2_nand3_1 _2196_ (.B(_1223_),
    .C(_1224_),
    .A(_1222_),
    .Y(_1225_));
 sg13g2_and2_1 _2197_ (.A(net667),
    .B(_1216_),
    .X(_1226_));
 sg13g2_a21oi_1 _2198_ (.A1(_1225_),
    .A2(_1226_),
    .Y(_1227_),
    .B1(net622));
 sg13g2_o21ai_1 _2199_ (.B1(_1168_),
    .Y(_1228_),
    .A1(_0951_),
    .A2(_1213_));
 sg13g2_a22oi_1 _2200_ (.Y(_1229_),
    .B1(_1228_),
    .B2(net719),
    .A2(_1176_),
    .A1(_1174_));
 sg13g2_nand2_1 _2201_ (.Y(_1230_),
    .A(net665),
    .B(_1229_));
 sg13g2_a221oi_1 _2202_ (.B2(_1042_),
    .C1(net666),
    .B1(_1182_),
    .A1(_1014_),
    .Y(_1231_),
    .A2(_1172_));
 sg13g2_a21oi_1 _2203_ (.A1(_1183_),
    .A2(_1231_),
    .Y(_1232_),
    .B1(net625));
 sg13g2_a221oi_1 _2204_ (.B2(_1232_),
    .C1(net620),
    .B1(_1230_),
    .A1(_1207_),
    .Y(_1233_),
    .A2(_1227_));
 sg13g2_nand3b_1 _2205_ (.B(_1089_),
    .C(_1080_),
    .Y(_1234_),
    .A_N(_1196_));
 sg13g2_nand2_1 _2206_ (.Y(_1235_),
    .A(_1154_),
    .B(_1234_));
 sg13g2_nand3_1 _2207_ (.B(net632),
    .C(net727),
    .A(_0958_),
    .Y(_1236_));
 sg13g2_nand3_1 _2208_ (.B(_1095_),
    .C(_1236_),
    .A(net736),
    .Y(_1237_));
 sg13g2_nand4_1 _2209_ (.B(_1093_),
    .C(_1235_),
    .A(net712),
    .Y(_1238_),
    .D(_1237_));
 sg13g2_nand2_1 _2210_ (.Y(_1239_),
    .A(net743),
    .B(_1202_));
 sg13g2_nand3_1 _2211_ (.B(_1103_),
    .C(_1239_),
    .A(net720),
    .Y(_1240_));
 sg13g2_nand2b_1 _2212_ (.Y(_1241_),
    .B(_1239_),
    .A_N(_1113_));
 sg13g2_nand3_1 _2213_ (.B(_1238_),
    .C(_1241_),
    .A(net668),
    .Y(_1242_));
 sg13g2_a21oi_2 _2214_ (.B1(net638),
    .Y(_1243_),
    .A2(net676),
    .A1(net660));
 sg13g2_a21oi_1 _2215_ (.A1(net676),
    .A2(net772),
    .Y(_1244_),
    .B1(_1004_));
 sg13g2_a22oi_1 _2216_ (.Y(_1245_),
    .B1(_1243_),
    .B2(_1244_),
    .A2(_1069_),
    .A1(net730));
 sg13g2_o21ai_1 _2217_ (.B1(_1245_),
    .Y(_1246_),
    .A1(_1019_),
    .A2(_1063_));
 sg13g2_nor2_1 _2218_ (.A(net737),
    .B(_1077_),
    .Y(_1247_));
 sg13g2_and2_1 _2219_ (.A(_1056_),
    .B(_1092_),
    .X(_1248_));
 sg13g2_nor2_2 _2220_ (.A(net742),
    .B(net730),
    .Y(_1249_));
 sg13g2_nand2_1 _2221_ (.Y(_1250_),
    .A(_0980_),
    .B(net740));
 sg13g2_nand2_1 _2222_ (.Y(_1251_),
    .A(net742),
    .B(net737));
 sg13g2_a22oi_1 _2223_ (.Y(_1252_),
    .B1(net631),
    .B2(net657),
    .A2(net635),
    .A1(net650));
 sg13g2_o21ai_1 _2224_ (.B1(net721),
    .Y(_1253_),
    .A1(_1251_),
    .A2(_1252_));
 sg13g2_a21oi_1 _2225_ (.A1(net766),
    .A2(_1083_),
    .Y(_1254_),
    .B1(_1247_));
 sg13g2_nor2_1 _2226_ (.A(_1248_),
    .B(_1253_),
    .Y(_1255_));
 sg13g2_a22oi_1 _2227_ (.Y(_1256_),
    .B1(_1254_),
    .B2(_1255_),
    .A2(_1246_),
    .A1(net713));
 sg13g2_a21oi_1 _2228_ (.A1(net664),
    .A2(_1256_),
    .Y(_1257_),
    .B1(net623));
 sg13g2_nor2_1 _2229_ (.A(_0978_),
    .B(_1011_),
    .Y(_1258_));
 sg13g2_nand2_1 _2230_ (.Y(_1259_),
    .A(net650),
    .B(net626));
 sg13g2_a21oi_1 _2231_ (.A1(_1010_),
    .A2(_1259_),
    .Y(_1260_),
    .B1(net757));
 sg13g2_nor2_1 _2232_ (.A(_0970_),
    .B(net742),
    .Y(_1261_));
 sg13g2_nor4_1 _2233_ (.A(net673),
    .B(_1258_),
    .C(_1260_),
    .D(_1261_),
    .Y(_1262_));
 sg13g2_a21oi_1 _2234_ (.A1(net673),
    .A2(_1041_),
    .Y(_1263_),
    .B1(_1262_));
 sg13g2_nand2_1 _2235_ (.Y(_1264_),
    .A(net664),
    .B(_1263_));
 sg13g2_nand3_1 _2236_ (.B(net646),
    .C(_1249_),
    .A(net658),
    .Y(_1265_));
 sg13g2_a21oi_1 _2237_ (.A1(_0970_),
    .A2(_1265_),
    .Y(_1266_),
    .B1(net720));
 sg13g2_a21oi_1 _2238_ (.A1(net646),
    .A2(_0983_),
    .Y(_1267_),
    .B1(net755));
 sg13g2_a21oi_1 _2239_ (.A1(net755),
    .A2(_1000_),
    .Y(_1268_),
    .B1(_1267_));
 sg13g2_a221oi_1 _2240_ (.B2(_1268_),
    .C1(_1266_),
    .B1(_1016_),
    .A1(_0974_),
    .Y(_1269_),
    .A2(_1005_));
 sg13g2_o21ai_1 _2241_ (.B1(_1269_),
    .Y(_1270_),
    .A1(_1002_),
    .A2(net673));
 sg13g2_a21oi_1 _2242_ (.A1(net668),
    .A2(_1270_),
    .Y(_1271_),
    .B1(net622));
 sg13g2_a221oi_1 _2243_ (.B2(_1271_),
    .C1(net619),
    .B1(_1264_),
    .A1(_1242_),
    .Y(_1272_),
    .A2(_1257_));
 sg13g2_nor3_1 _2244_ (.A(_1118_),
    .B(_1233_),
    .C(_1272_),
    .Y(_1273_));
 sg13g2_o21ai_1 _2245_ (.B1(_0887_),
    .Y(_1274_),
    .A1(_1193_),
    .A2(_1273_));
 sg13g2_xnor2_1 _2246_ (.Y(_1275_),
    .A(_0924_),
    .B(_0927_));
 sg13g2_inv_1 _2247_ (.Y(_1276_),
    .A(_1275_));
 sg13g2_nand4_1 _2248_ (.B(net643),
    .C(net633),
    .A(net763),
    .Y(_1277_),
    .D(_1086_));
 sg13g2_nand3_1 _2249_ (.B(_1109_),
    .C(_1277_),
    .A(net729),
    .Y(_1278_));
 sg13g2_and2_1 _2250_ (.A(_1203_),
    .B(_1278_),
    .X(_1279_));
 sg13g2_a21oi_1 _2251_ (.A1(_1122_),
    .A2(_1279_),
    .Y(_1280_),
    .B1(net725));
 sg13g2_nor3_2 _2252_ (.A(net769),
    .B(_1036_),
    .C(_1057_),
    .Y(_1281_));
 sg13g2_a21oi_1 _2253_ (.A1(net773),
    .A2(_1125_),
    .Y(_1282_),
    .B1(_1281_));
 sg13g2_a21o_1 _2254_ (.A2(_1125_),
    .A1(net773),
    .B1(_1281_),
    .X(_1283_));
 sg13g2_o21ai_1 _2255_ (.B1(_1200_),
    .Y(_1284_),
    .A1(net756),
    .A2(_1283_));
 sg13g2_o21ai_1 _2256_ (.B1(net750),
    .Y(_1285_),
    .A1(_1131_),
    .A2(_1196_));
 sg13g2_a21oi_1 _2257_ (.A1(_1133_),
    .A2(_1285_),
    .Y(_1286_),
    .B1(net716));
 sg13g2_a21o_1 _2258_ (.A2(_1153_),
    .A1(net765),
    .B1(_1086_),
    .X(_1287_));
 sg13g2_o21ai_1 _2259_ (.B1(net712),
    .Y(_1288_),
    .A1(_0993_),
    .A2(_1220_));
 sg13g2_a21oi_1 _2260_ (.A1(net702),
    .A2(_1287_),
    .Y(_1289_),
    .B1(_1288_));
 sg13g2_nor2_1 _2261_ (.A(net731),
    .B(_1066_),
    .Y(_1290_));
 sg13g2_nand2_1 _2262_ (.Y(_1291_),
    .A(net736),
    .B(net727));
 sg13g2_a21oi_1 _2263_ (.A1(_1221_),
    .A2(_1290_),
    .Y(_1292_),
    .B1(_1219_));
 sg13g2_nand2_1 _2264_ (.Y(_1293_),
    .A(_1289_),
    .B(_1292_));
 sg13g2_o21ai_1 _2265_ (.B1(net765),
    .Y(_1294_),
    .A1(_1035_),
    .A2(net637));
 sg13g2_nand2_1 _2266_ (.Y(_1295_),
    .A(net772),
    .B(_1148_));
 sg13g2_a21o_1 _2267_ (.A2(_1295_),
    .A1(_1294_),
    .B1(net700),
    .X(_1296_));
 sg13g2_nand3b_1 _2268_ (.B(_1209_),
    .C(_1296_),
    .Y(_1297_),
    .A_N(_1140_));
 sg13g2_a21oi_1 _2269_ (.A1(_1293_),
    .A2(_1297_),
    .Y(_1298_),
    .B1(net664));
 sg13g2_a21o_1 _2270_ (.A2(_1286_),
    .A1(_1284_),
    .B1(net671),
    .X(_1299_));
 sg13g2_o21ai_1 _2271_ (.B1(net624),
    .Y(_1300_),
    .A1(_1280_),
    .A2(_1299_));
 sg13g2_nand3_1 _2272_ (.B(net732),
    .C(_1110_),
    .A(net682),
    .Y(_1301_));
 sg13g2_o21ai_1 _2273_ (.B1(_1301_),
    .Y(_1302_),
    .A1(net757),
    .A2(_1167_));
 sg13g2_a22oi_1 _2274_ (.Y(_1303_),
    .B1(net626),
    .B2(net743),
    .A2(_1152_),
    .A1(_1066_));
 sg13g2_or2_1 _2275_ (.X(_1304_),
    .B(net626),
    .A(net642));
 sg13g2_o21ai_1 _2276_ (.B1(net705),
    .Y(_1305_),
    .A1(net642),
    .A2(_1181_));
 sg13g2_and2_1 _2277_ (.A(net718),
    .B(_1305_),
    .X(_1306_));
 sg13g2_a221oi_1 _2278_ (.B2(net681),
    .C1(net688),
    .B1(net710),
    .A1(net696),
    .Y(_1307_),
    .A2(net693));
 sg13g2_inv_1 _2279_ (.Y(_1308_),
    .A(_1307_));
 sg13g2_nor2_1 _2280_ (.A(net626),
    .B(_1307_),
    .Y(_1309_));
 sg13g2_nor2_1 _2281_ (.A(_1249_),
    .B(_1309_),
    .Y(_1310_));
 sg13g2_o21ai_1 _2282_ (.B1(net768),
    .Y(_1311_),
    .A1(_1033_),
    .A2(net626));
 sg13g2_nand3_1 _2283_ (.B(_1305_),
    .C(_1311_),
    .A(net717),
    .Y(_1312_));
 sg13g2_o21ai_1 _2284_ (.B1(net704),
    .Y(_1313_),
    .A1(_1033_),
    .A2(net626));
 sg13g2_nand3_1 _2285_ (.B(_1041_),
    .C(_1313_),
    .A(net722),
    .Y(_1314_));
 sg13g2_a21oi_1 _2286_ (.A1(_1023_),
    .A2(_1175_),
    .Y(_1315_),
    .B1(net670));
 sg13g2_o21ai_1 _2287_ (.B1(_1315_),
    .Y(_1316_),
    .A1(_1021_),
    .A2(_1303_));
 sg13g2_a21o_1 _2288_ (.A2(_1302_),
    .A1(net718),
    .B1(_1316_),
    .X(_1317_));
 sg13g2_o21ai_1 _2289_ (.B1(_1314_),
    .Y(_1318_),
    .A1(_1310_),
    .A2(_1312_));
 sg13g2_a21oi_1 _2290_ (.A1(net669),
    .A2(_1318_),
    .Y(_1319_),
    .B1(net625));
 sg13g2_a21oi_1 _2291_ (.A1(_1317_),
    .A2(_1319_),
    .Y(_1320_),
    .B1(net620));
 sg13g2_o21ai_1 _2292_ (.B1(_1320_),
    .Y(_1321_),
    .A1(_1298_),
    .A2(_1300_));
 sg13g2_nand4_1 _2293_ (.B(net643),
    .C(net632),
    .A(net763),
    .Y(_1322_),
    .D(net630));
 sg13g2_nand3b_1 _2294_ (.B(net770),
    .C(net633),
    .Y(_1323_),
    .A_N(_1094_));
 sg13g2_nand2_1 _2295_ (.Y(_1324_),
    .A(_1322_),
    .B(_1323_));
 sg13g2_nand3_1 _2296_ (.B(_1322_),
    .C(_1323_),
    .A(net698),
    .Y(_1325_));
 sg13g2_nand2_1 _2297_ (.Y(_1326_),
    .A(net749),
    .B(_1095_));
 sg13g2_a21oi_1 _2298_ (.A1(_0958_),
    .A2(net632),
    .Y(_1327_),
    .B1(_1004_));
 sg13g2_o21ai_1 _2299_ (.B1(net712),
    .Y(_1328_),
    .A1(net640),
    .A2(_1291_));
 sg13g2_a221oi_1 _2300_ (.B2(_1095_),
    .C1(_1328_),
    .B1(_1327_),
    .A1(net706),
    .Y(_1329_),
    .A2(_1234_));
 sg13g2_o21ai_1 _2301_ (.B1(net703),
    .Y(_1330_),
    .A1(_1087_),
    .A2(_1091_));
 sg13g2_nand3_1 _2302_ (.B(_1329_),
    .C(_1330_),
    .A(_1325_),
    .Y(_1331_));
 sg13g2_a21oi_1 _2303_ (.A1(_1022_),
    .A2(_1109_),
    .Y(_1332_),
    .B1(net663));
 sg13g2_nor2_1 _2304_ (.A(net764),
    .B(_1202_),
    .Y(_1333_));
 sg13g2_nand2_1 _2305_ (.Y(_1334_),
    .A(net674),
    .B(_1120_));
 sg13g2_o21ai_1 _2306_ (.B1(_1332_),
    .Y(_1335_),
    .A1(_1333_),
    .A2(_1334_));
 sg13g2_a221oi_1 _2307_ (.B2(_1331_),
    .C1(_1335_),
    .B1(_1240_),
    .A1(_1022_),
    .Y(_1336_),
    .A2(net627));
 sg13g2_a21oi_1 _2308_ (.A1(_1055_),
    .A2(_1088_),
    .Y(_1337_),
    .B1(net730));
 sg13g2_nor2_1 _2309_ (.A(_1155_),
    .B(_1252_),
    .Y(_1338_));
 sg13g2_or4_1 _2310_ (.A(_1248_),
    .B(_1253_),
    .C(_1337_),
    .D(_1338_),
    .X(_1339_));
 sg13g2_and2_1 _2311_ (.A(_1062_),
    .B(_1249_),
    .X(_1340_));
 sg13g2_nor2_1 _2312_ (.A(net702),
    .B(_1249_),
    .Y(_1341_));
 sg13g2_nor2b_1 _2313_ (.A(_1243_),
    .B_N(_1341_),
    .Y(_1342_));
 sg13g2_nor2b_1 _2314_ (.A(_1064_),
    .B_N(_1092_),
    .Y(_1343_));
 sg13g2_or4_1 _2315_ (.A(net721),
    .B(_1340_),
    .C(_1342_),
    .D(_1343_),
    .X(_1344_));
 sg13g2_a21oi_1 _2316_ (.A1(_1339_),
    .A2(_1344_),
    .Y(_1345_),
    .B1(net667));
 sg13g2_or3_1 _2317_ (.A(net623),
    .B(_1336_),
    .C(_1345_),
    .X(_1346_));
 sg13g2_a21oi_1 _2318_ (.A1(net650),
    .A2(net626),
    .Y(_1347_),
    .B1(_1307_));
 sg13g2_a21oi_1 _2319_ (.A1(_0969_),
    .A2(_1308_),
    .Y(_1348_),
    .B1(_1212_));
 sg13g2_o21ai_1 _2320_ (.B1(_1265_),
    .Y(_1349_),
    .A1(_1213_),
    .A2(_1347_));
 sg13g2_o21ai_1 _2321_ (.B1(net717),
    .Y(_1350_),
    .A1(_1348_),
    .A2(_1349_));
 sg13g2_nor2_1 _2322_ (.A(_1000_),
    .B(_1144_),
    .Y(_1351_));
 sg13g2_a21oi_1 _2323_ (.A1(_0969_),
    .A2(_0997_),
    .Y(_1352_),
    .B1(_1017_));
 sg13g2_nor3_1 _2324_ (.A(net665),
    .B(_1351_),
    .C(_1352_),
    .Y(_1353_));
 sg13g2_nand2b_1 _2325_ (.Y(_1354_),
    .B(net674),
    .A_N(_1347_));
 sg13g2_nor2_1 _2326_ (.A(net719),
    .B(_1065_),
    .Y(_1355_));
 sg13g2_o21ai_1 _2327_ (.B1(_1355_),
    .Y(_1356_),
    .A1(_1038_),
    .A2(_1307_));
 sg13g2_or2_1 _2328_ (.X(_1357_),
    .B(_1143_),
    .A(_1041_));
 sg13g2_nand4_1 _2329_ (.B(_1354_),
    .C(_1356_),
    .A(net665),
    .Y(_1358_),
    .D(_1357_));
 sg13g2_a21oi_1 _2330_ (.A1(_1350_),
    .A2(_1353_),
    .Y(_1359_),
    .B1(net622));
 sg13g2_a21oi_1 _2331_ (.A1(_1358_),
    .A2(_1359_),
    .Y(_1360_),
    .B1(net619));
 sg13g2_a21oi_1 _2332_ (.A1(_1346_),
    .A2(_1360_),
    .Y(_1361_),
    .B1(_1117_));
 sg13g2_a21oi_1 _2333_ (.A1(net740),
    .A2(_1175_),
    .Y(_1362_),
    .B1(net724));
 sg13g2_a21o_1 _2334_ (.A2(_1164_),
    .A1(net647),
    .B1(_1138_),
    .X(_1363_));
 sg13g2_a22oi_1 _2335_ (.Y(_1364_),
    .B1(_1363_),
    .B2(net704),
    .A2(_1168_),
    .A1(net706));
 sg13g2_nand2_1 _2336_ (.Y(_1365_),
    .A(net733),
    .B(_1175_));
 sg13g2_a21o_1 _2337_ (.A2(net628),
    .A1(_1097_),
    .B1(_1162_),
    .X(_1366_));
 sg13g2_a221oi_1 _2338_ (.B2(_1003_),
    .C1(net716),
    .B1(_1366_),
    .A1(_1171_),
    .Y(_1367_),
    .A2(_1304_));
 sg13g2_a22oi_1 _2339_ (.Y(_1368_),
    .B1(_1365_),
    .B2(_1367_),
    .A2(_1364_),
    .A1(_1362_));
 sg13g2_a21oi_2 _2340_ (.B1(_1307_),
    .Y(_1369_),
    .A2(_1036_),
    .A1(_0952_));
 sg13g2_a22oi_1 _2341_ (.Y(_1370_),
    .B1(_1369_),
    .B2(net722),
    .A2(_1309_),
    .A1(_1306_));
 sg13g2_nor2_1 _2342_ (.A(net701),
    .B(_1309_),
    .Y(_1371_));
 sg13g2_nand2_1 _2343_ (.Y(_1372_),
    .A(net665),
    .B(_1368_));
 sg13g2_o21ai_1 _2344_ (.B1(net669),
    .Y(_1373_),
    .A1(_1370_),
    .A2(_1371_));
 sg13g2_nand3_1 _2345_ (.B(_1372_),
    .C(_1373_),
    .A(net622),
    .Y(_1374_));
 sg13g2_a21oi_1 _2346_ (.A1(net704),
    .A2(_1120_),
    .Y(_1375_),
    .B1(net725));
 sg13g2_a22oi_1 _2347_ (.Y(_1376_),
    .B1(net627),
    .B2(net679),
    .A2(_1057_),
    .A1(_0959_));
 sg13g2_or2_1 _2348_ (.X(_1377_),
    .B(_1376_),
    .A(_0978_));
 sg13g2_a21o_1 _2349_ (.A2(_1377_),
    .A1(_1285_),
    .B1(net732),
    .X(_1378_));
 sg13g2_a21oi_1 _2350_ (.A1(net698),
    .A2(_1086_),
    .Y(_1379_),
    .B1(net714));
 sg13g2_o21ai_1 _2351_ (.B1(_1379_),
    .Y(_1380_),
    .A1(net640),
    .A2(_1155_));
 sg13g2_a221oi_1 _2352_ (.B2(net704),
    .C1(_1380_),
    .B1(_1282_),
    .A1(_0992_),
    .Y(_1381_),
    .A2(_1199_));
 sg13g2_a221oi_1 _2353_ (.B2(_1381_),
    .C1(net671),
    .B1(_1378_),
    .A1(_1279_),
    .Y(_1382_),
    .A2(_1375_));
 sg13g2_o21ai_1 _2354_ (.B1(net771),
    .Y(_1383_),
    .A1(net637),
    .A2(net634));
 sg13g2_nand3_1 _2355_ (.B(_1294_),
    .C(_1383_),
    .A(net754),
    .Y(_1384_));
 sg13g2_a21oi_1 _2356_ (.A1(net749),
    .A2(_1220_),
    .Y(_1385_),
    .B1(net730));
 sg13g2_a221oi_1 _2357_ (.B2(_1385_),
    .C1(_1288_),
    .B1(_1384_),
    .A1(net702),
    .Y(_1386_),
    .A2(_1287_));
 sg13g2_nand2b_1 _2358_ (.Y(_1387_),
    .B(_1139_),
    .A_N(_1251_));
 sg13g2_a22oi_1 _2359_ (.Y(_1388_),
    .B1(_1249_),
    .B2(_1363_),
    .A2(_1208_),
    .A1(net702));
 sg13g2_nand3_1 _2360_ (.B(_1387_),
    .C(_1388_),
    .A(_1209_),
    .Y(_1389_));
 sg13g2_nand3b_1 _2361_ (.B(_1389_),
    .C(net667),
    .Y(_1390_),
    .A_N(_1386_));
 sg13g2_nand3b_1 _2362_ (.B(_1390_),
    .C(net623),
    .Y(_1391_),
    .A_N(_1382_));
 sg13g2_a21oi_1 _2363_ (.A1(_1374_),
    .A2(_1391_),
    .Y(_1392_),
    .B1(net620));
 sg13g2_a21o_1 _2364_ (.A2(_1088_),
    .A1(_1055_),
    .B1(net700),
    .X(_1393_));
 sg13g2_nand2b_1 _2365_ (.Y(_1394_),
    .B(_1214_),
    .A_N(_1376_));
 sg13g2_nand4_1 _2366_ (.B(_1329_),
    .C(_1393_),
    .A(_1325_),
    .Y(_1395_),
    .D(_1394_));
 sg13g2_a21oi_1 _2367_ (.A1(_1240_),
    .A2(_1395_),
    .Y(_1396_),
    .B1(_1335_));
 sg13g2_nand2b_1 _2368_ (.Y(_1397_),
    .B(net771),
    .A_N(_1243_));
 sg13g2_a21oi_1 _2369_ (.A1(net765),
    .A2(_1056_),
    .Y(_1398_),
    .B1(net753));
 sg13g2_a221oi_1 _2370_ (.B2(_1398_),
    .C1(net737),
    .B1(_1397_),
    .A1(net753),
    .Y(_1399_),
    .A2(_1252_));
 sg13g2_nor3_1 _2371_ (.A(_1253_),
    .B(_1337_),
    .C(_1399_),
    .Y(_1400_));
 sg13g2_nor2_1 _2372_ (.A(net771),
    .B(net638),
    .Y(_1401_));
 sg13g2_nand2_1 _2373_ (.Y(_1402_),
    .A(net765),
    .B(_1064_));
 sg13g2_nor4_1 _2374_ (.A(net676),
    .B(_0974_),
    .C(net767),
    .D(_1060_),
    .Y(_1403_));
 sg13g2_nor2_1 _2375_ (.A(net700),
    .B(_1403_),
    .Y(_1404_));
 sg13g2_o21ai_1 _2376_ (.B1(net713),
    .Y(_1405_),
    .A1(net702),
    .A2(_1243_));
 sg13g2_a21oi_1 _2377_ (.A1(_1402_),
    .A2(_1404_),
    .Y(_1406_),
    .B1(_1405_));
 sg13g2_o21ai_1 _2378_ (.B1(net664),
    .Y(_1407_),
    .A1(_1400_),
    .A2(_1406_));
 sg13g2_nor2_1 _2379_ (.A(net623),
    .B(_1396_),
    .Y(_1408_));
 sg13g2_or2_1 _2380_ (.X(_1409_),
    .B(_1347_),
    .A(net741));
 sg13g2_a21o_1 _2381_ (.A2(_1308_),
    .A1(_0969_),
    .B1(_1004_),
    .X(_1410_));
 sg13g2_a21oi_1 _2382_ (.A1(_1409_),
    .A2(_1410_),
    .Y(_1411_),
    .B1(net723));
 sg13g2_o21ai_1 _2383_ (.B1(net668),
    .Y(_1412_),
    .A1(net673),
    .A2(_1069_));
 sg13g2_o21ai_1 _2384_ (.B1(net699),
    .Y(_1413_),
    .A1(net768),
    .A2(_1152_));
 sg13g2_a22oi_1 _2385_ (.Y(_1414_),
    .B1(_1413_),
    .B2(net717),
    .A2(_0997_),
    .A1(_0969_));
 sg13g2_nor3_1 _2386_ (.A(_1411_),
    .B(_1412_),
    .C(_1414_),
    .Y(_1415_));
 sg13g2_nand3_1 _2387_ (.B(_1354_),
    .C(_1369_),
    .A(net665),
    .Y(_1416_));
 sg13g2_nand2_1 _2388_ (.Y(_1417_),
    .A(net625),
    .B(_1416_));
 sg13g2_o21ai_1 _2389_ (.B1(net620),
    .Y(_1418_),
    .A1(_1415_),
    .A2(_1417_));
 sg13g2_a21oi_1 _2390_ (.A1(_1407_),
    .A2(_1408_),
    .Y(_1419_),
    .B1(_1418_));
 sg13g2_or3_1 _2391_ (.A(_1118_),
    .B(_1392_),
    .C(_1419_),
    .X(_1420_));
 sg13g2_a21oi_1 _2392_ (.A1(_1321_),
    .A2(_1361_),
    .Y(_1421_),
    .B1(_0887_));
 sg13g2_a21oi_1 _2393_ (.A1(_1420_),
    .A2(_1421_),
    .Y(_1422_),
    .B1(_1275_));
 sg13g2_o21ai_1 _2394_ (.B1(net752),
    .Y(_1423_),
    .A1(_1075_),
    .A2(_1132_));
 sg13g2_nand3_1 _2395_ (.B(_1135_),
    .C(_1423_),
    .A(net739),
    .Y(_1424_));
 sg13g2_a21oi_1 _2396_ (.A1(_1128_),
    .A2(_1424_),
    .Y(_1425_),
    .B1(net716));
 sg13g2_a21oi_1 _2397_ (.A1(net768),
    .A2(_1095_),
    .Y(_1426_),
    .B1(net720));
 sg13g2_and3_1 _2398_ (.X(_1427_),
    .A(_1123_),
    .B(_1124_),
    .C(_1426_));
 sg13g2_o21ai_1 _2399_ (.B1(net624),
    .Y(_1428_),
    .A1(_1425_),
    .A2(_1427_));
 sg13g2_a22oi_1 _2400_ (.Y(_1429_),
    .B1(net684),
    .B2(_0958_),
    .A2(net690),
    .A1(net692));
 sg13g2_nand2_1 _2401_ (.Y(_1430_),
    .A(_1008_),
    .B(_1429_));
 sg13g2_a21oi_2 _2402_ (.B1(_1162_),
    .Y(_1431_),
    .A2(_1429_),
    .A1(_1008_));
 sg13g2_or2_1 _2403_ (.X(_1432_),
    .B(_1431_),
    .A(net740));
 sg13g2_o21ai_1 _2404_ (.B1(net740),
    .Y(_1433_),
    .A1(net627),
    .A2(_1175_));
 sg13g2_a21oi_1 _2405_ (.A1(_1432_),
    .A2(_1433_),
    .Y(_1434_),
    .B1(net725));
 sg13g2_or2_1 _2406_ (.X(_1435_),
    .B(_1164_),
    .A(net644));
 sg13g2_a22oi_1 _2407_ (.Y(_1436_),
    .B1(_1435_),
    .B2(_0989_),
    .A2(_1173_),
    .A1(net756));
 sg13g2_a21o_2 _2408_ (.A2(net648),
    .A1(net652),
    .B1(net627),
    .X(_1437_));
 sg13g2_a21oi_1 _2409_ (.A1(net751),
    .A2(_1437_),
    .Y(_1438_),
    .B1(net732));
 sg13g2_a21oi_1 _2410_ (.A1(_0981_),
    .A2(_1162_),
    .Y(_1439_),
    .B1(_1437_));
 sg13g2_a221oi_1 _2411_ (.B2(net732),
    .C1(net718),
    .B1(_1439_),
    .A1(_1436_),
    .Y(_1440_),
    .A2(_1438_));
 sg13g2_nor3_1 _2412_ (.A(net625),
    .B(_1434_),
    .C(_1440_),
    .Y(_1441_));
 sg13g2_nor2_1 _2413_ (.A(net670),
    .B(_1441_),
    .Y(_1442_));
 sg13g2_o21ai_1 _2414_ (.B1(_1146_),
    .Y(_1443_),
    .A1(_1047_),
    .A2(_1060_));
 sg13g2_and2_1 _2415_ (.A(_1145_),
    .B(_1443_),
    .X(_1444_));
 sg13g2_nor2_1 _2416_ (.A(net729),
    .B(_1431_),
    .Y(_1445_));
 sg13g2_a21oi_2 _2417_ (.B1(_1162_),
    .Y(_1446_),
    .A2(_1047_),
    .A1(net640));
 sg13g2_a21oi_1 _2418_ (.A1(_1155_),
    .A2(_1291_),
    .Y(_1447_),
    .B1(_1446_));
 sg13g2_nor2_1 _2419_ (.A(_1445_),
    .B(_1447_),
    .Y(_1448_));
 sg13g2_nand2_1 _2420_ (.Y(_1449_),
    .A(net653),
    .B(_0967_));
 sg13g2_a22oi_1 _2421_ (.Y(_1450_),
    .B1(_1057_),
    .B2(net709),
    .A2(_0967_),
    .A1(net654));
 sg13g2_nand2_1 _2422_ (.Y(_1451_),
    .A(_1034_),
    .B(_1130_));
 sg13g2_a22oi_1 _2423_ (.Y(_1452_),
    .B1(_1451_),
    .B2(_1146_),
    .A2(_1450_),
    .A1(_1154_));
 sg13g2_a221oi_1 _2424_ (.B2(_1151_),
    .C1(net622),
    .B1(_1452_),
    .A1(_1444_),
    .Y(_1453_),
    .A2(_1448_));
 sg13g2_a21oi_1 _2425_ (.A1(net642),
    .A2(net639),
    .Y(_1454_),
    .B1(_1147_));
 sg13g2_a21o_1 _2426_ (.A2(net639),
    .A1(net642),
    .B1(_1147_),
    .X(_1455_));
 sg13g2_nand2_2 _2427_ (.Y(_1456_),
    .A(net644),
    .B(net639));
 sg13g2_a21o_1 _2428_ (.A2(net639),
    .A1(net644),
    .B1(net652),
    .X(_1457_));
 sg13g2_a21oi_1 _2429_ (.A1(net704),
    .A2(_1457_),
    .Y(_1458_),
    .B1(_1455_));
 sg13g2_a21oi_1 _2430_ (.A1(_1045_),
    .A2(_1249_),
    .Y(_1459_),
    .B1(net717));
 sg13g2_o21ai_1 _2431_ (.B1(_1187_),
    .Y(_1460_),
    .A1(_1019_),
    .A2(_1456_));
 sg13g2_a21oi_1 _2432_ (.A1(_1458_),
    .A2(_1459_),
    .Y(_1461_),
    .B1(net625));
 sg13g2_a21o_1 _2433_ (.A2(_1461_),
    .A1(_1460_),
    .B1(_1453_),
    .X(_1462_));
 sg13g2_a221oi_1 _2434_ (.B2(net670),
    .C1(_0908_),
    .B1(_1462_),
    .A1(_1428_),
    .Y(_1463_),
    .A2(_1442_));
 sg13g2_nand3_1 _2435_ (.B(_1112_),
    .C(_1324_),
    .A(net720),
    .Y(_1464_));
 sg13g2_a21oi_1 _2436_ (.A1(net752),
    .A2(_1104_),
    .Y(_1465_),
    .B1(_1464_));
 sg13g2_a221oi_1 _2437_ (.B2(net769),
    .C1(_1099_),
    .B1(_1087_),
    .A1(net662),
    .Y(_1466_),
    .A2(_1006_));
 sg13g2_nor2_1 _2438_ (.A(net736),
    .B(_1466_),
    .Y(_1467_));
 sg13g2_a22oi_1 _2439_ (.Y(_1468_),
    .B1(_1214_),
    .B2(_1090_),
    .A2(_1212_),
    .A1(_1082_));
 sg13g2_nand2_1 _2440_ (.Y(_1469_),
    .A(net712),
    .B(_1468_));
 sg13g2_a21oi_1 _2441_ (.A1(net643),
    .A2(net632),
    .Y(_1470_),
    .B1(net728));
 sg13g2_nor3_1 _2442_ (.A(_1467_),
    .B(_1469_),
    .C(_1470_),
    .Y(_1471_));
 sg13g2_o21ai_1 _2443_ (.B1(net668),
    .Y(_1472_),
    .A1(_1465_),
    .A2(_1471_));
 sg13g2_a21oi_2 _2444_ (.B1(net657),
    .Y(_1473_),
    .A2(_0961_),
    .A1(_0957_));
 sg13g2_nor2_1 _2445_ (.A(net637),
    .B(_1473_),
    .Y(_1474_));
 sg13g2_o21ai_1 _2446_ (.B1(net766),
    .Y(_1475_),
    .A1(net660),
    .A2(net709));
 sg13g2_o21ai_1 _2447_ (.B1(_1475_),
    .Y(_1476_),
    .A1(net766),
    .A2(_0996_));
 sg13g2_a21oi_2 _2448_ (.B1(net688),
    .Y(_1477_),
    .A2(net687),
    .A1(_0949_));
 sg13g2_nor2_1 _2449_ (.A(net753),
    .B(_1477_),
    .Y(_1478_));
 sg13g2_a221oi_1 _2450_ (.B2(_1478_),
    .C1(net730),
    .B1(_1476_),
    .A1(net753),
    .Y(_1479_),
    .A2(_1474_));
 sg13g2_a21oi_2 _2451_ (.B1(_0996_),
    .Y(_1480_),
    .A2(net647),
    .A1(net677));
 sg13g2_nand2_1 _2452_ (.Y(_1481_),
    .A(net753),
    .B(_1477_));
 sg13g2_a21o_1 _2453_ (.A2(_1481_),
    .A1(_1480_),
    .B1(net737),
    .X(_1482_));
 sg13g2_and2_1 _2454_ (.A(net771),
    .B(_1480_),
    .X(_1483_));
 sg13g2_o21ai_1 _2455_ (.B1(net713),
    .Y(_1484_),
    .A1(_1482_),
    .A2(_1483_));
 sg13g2_or2_1 _2456_ (.X(_1485_),
    .B(_1138_),
    .A(_1006_));
 sg13g2_o21ai_1 _2457_ (.B1(_0957_),
    .Y(_0117_),
    .A1(net661),
    .A2(net709));
 sg13g2_a22oi_1 _2458_ (.Y(_0118_),
    .B1(_0117_),
    .B2(net727),
    .A2(_1082_),
    .A1(net753));
 sg13g2_a21oi_1 _2459_ (.A1(_0989_),
    .A2(_1485_),
    .Y(_0119_),
    .B1(net673));
 sg13g2_a22oi_1 _2460_ (.Y(_0120_),
    .B1(_0118_),
    .B2(_0119_),
    .A2(_1474_),
    .A1(_1016_));
 sg13g2_o21ai_1 _2461_ (.B1(_0120_),
    .Y(_0121_),
    .A1(_1479_),
    .A2(_1484_));
 sg13g2_a21oi_1 _2462_ (.A1(net664),
    .A2(_0121_),
    .Y(_0122_),
    .B1(net623));
 sg13g2_a221oi_1 _2463_ (.B2(net750),
    .C1(_1017_),
    .B1(_1455_),
    .A1(_1034_),
    .Y(_0123_),
    .A2(_1048_));
 sg13g2_a22oi_1 _2464_ (.Y(_0124_),
    .B1(net649),
    .B2(net645),
    .A2(_0967_),
    .A1(net653));
 sg13g2_a221oi_1 _2465_ (.B2(net674),
    .C1(_0123_),
    .B1(_0124_),
    .A1(_1046_),
    .Y(_0125_),
    .A2(_1454_));
 sg13g2_nand2_2 _2466_ (.Y(_0126_),
    .A(_0953_),
    .B(net629));
 sg13g2_nand3_1 _2467_ (.B(_0953_),
    .C(net629),
    .A(net757),
    .Y(_0127_));
 sg13g2_a22oi_1 _2468_ (.Y(_0128_),
    .B1(_0127_),
    .B2(_0965_),
    .A2(_0990_),
    .A1(_0978_));
 sg13g2_a21oi_1 _2469_ (.A1(_1010_),
    .A2(_0126_),
    .Y(_0129_),
    .B1(net757));
 sg13g2_a22oi_1 _2470_ (.Y(_0130_),
    .B1(net646),
    .B2(net658),
    .A2(net647),
    .A1(_0953_));
 sg13g2_o21ai_1 _2471_ (.B1(net741),
    .Y(_0131_),
    .A1(_0981_),
    .A2(_0130_));
 sg13g2_or3_1 _2472_ (.A(_0128_),
    .B(_0129_),
    .C(_0131_),
    .X(_0132_));
 sg13g2_nand3_1 _2473_ (.B(_0124_),
    .C(_0127_),
    .A(net733),
    .Y(_0133_));
 sg13g2_and2_1 _2474_ (.A(net716),
    .B(_0133_),
    .X(_0134_));
 sg13g2_a221oi_1 _2475_ (.B2(net676),
    .C1(net774),
    .B1(net647),
    .A1(net658),
    .Y(_0135_),
    .A2(net650));
 sg13g2_a22oi_1 _2476_ (.Y(_0136_),
    .B1(net646),
    .B2(net658),
    .A2(net647),
    .A1(net676));
 sg13g2_inv_1 _2477_ (.Y(_0137_),
    .A(_0136_));
 sg13g2_a21oi_1 _2478_ (.A1(net774),
    .A2(_0136_),
    .Y(_0138_),
    .B1(_0135_));
 sg13g2_a21o_1 _2479_ (.A2(_0136_),
    .A1(net774),
    .B1(_0135_),
    .X(_0139_));
 sg13g2_o21ai_1 _2480_ (.B1(net669),
    .Y(_0140_),
    .A1(_1017_),
    .A2(_0130_));
 sg13g2_nand2_1 _2481_ (.Y(_0141_),
    .A(net758),
    .B(_1480_));
 sg13g2_a21oi_1 _2482_ (.A1(net750),
    .A2(_0139_),
    .Y(_0142_),
    .B1(net673));
 sg13g2_a221oi_1 _2483_ (.B2(_0142_),
    .C1(_0140_),
    .B1(_0141_),
    .A1(_0132_),
    .Y(_0143_),
    .A2(_0134_));
 sg13g2_o21ai_1 _2484_ (.B1(net623),
    .Y(_0144_),
    .A1(net669),
    .A2(_0125_));
 sg13g2_o21ai_1 _2485_ (.B1(net620),
    .Y(_0145_),
    .A1(_0143_),
    .A2(_0144_));
 sg13g2_a21oi_1 _2486_ (.A1(_1472_),
    .A2(_0122_),
    .Y(_0146_),
    .B1(_0145_));
 sg13g2_or3_1 _2487_ (.A(_1118_),
    .B(_1463_),
    .C(_0146_),
    .X(_0147_));
 sg13g2_nand4_1 _2488_ (.B(_1037_),
    .C(net633),
    .A(net769),
    .Y(_0148_),
    .D(net630));
 sg13g2_or2_1 _2489_ (.X(_0149_),
    .B(net628),
    .A(net641));
 sg13g2_nor3_2 _2490_ (.A(net770),
    .B(net641),
    .C(net628),
    .Y(_0150_));
 sg13g2_nand2_1 _2491_ (.Y(_0151_),
    .A(net758),
    .B(_0148_));
 sg13g2_nor2_1 _2492_ (.A(_0150_),
    .B(_0151_),
    .Y(_0152_));
 sg13g2_nand3b_1 _2493_ (.B(net752),
    .C(_0148_),
    .Y(_0153_),
    .A_N(_0150_));
 sg13g2_nand4_1 _2494_ (.B(_1112_),
    .C(_1324_),
    .A(net720),
    .Y(_0154_),
    .D(_0153_));
 sg13g2_o21ai_1 _2495_ (.B1(net768),
    .Y(_0155_),
    .A1(_1036_),
    .A2(_1099_));
 sg13g2_mux4_1 _2496_ (.S0(net769),
    .A0(net678),
    .A1(_1006_),
    .A2(_1098_),
    .A3(_1086_),
    .S1(net655),
    .X(_0156_));
 sg13g2_a22oi_1 _2497_ (.Y(_0157_),
    .B1(_0156_),
    .B2(net706),
    .A2(_1470_),
    .A1(net763));
 sg13g2_nand3_1 _2498_ (.B(net643),
    .C(net632),
    .A(net752),
    .Y(_0158_));
 sg13g2_a22oi_1 _2499_ (.Y(_0159_),
    .B1(net643),
    .B2(net632),
    .A2(_0960_),
    .A1(net655));
 sg13g2_inv_1 _2500_ (.Y(_0160_),
    .A(_0159_));
 sg13g2_a221oi_1 _2501_ (.B2(net632),
    .C1(net728),
    .B1(net643),
    .A1(net655),
    .Y(_0161_),
    .A2(_0960_));
 sg13g2_nor2_1 _2502_ (.A(net698),
    .B(_0161_),
    .Y(_0162_));
 sg13g2_o21ai_1 _2503_ (.B1(_0158_),
    .Y(_0163_),
    .A1(net698),
    .A2(_0161_));
 sg13g2_nand4_1 _2504_ (.B(_1468_),
    .C(_0157_),
    .A(net712),
    .Y(_0164_),
    .D(_0163_));
 sg13g2_a21oi_1 _2505_ (.A1(_0154_),
    .A2(_0164_),
    .Y(_0165_),
    .B1(net663));
 sg13g2_mux2_1 _2506_ (.A0(net637),
    .A1(_1060_),
    .S(net771),
    .X(_0166_));
 sg13g2_o21ai_1 _2507_ (.B1(net698),
    .Y(_0167_),
    .A1(_1473_),
    .A2(_0166_));
 sg13g2_nand2_1 _2508_ (.Y(_0168_),
    .A(_1290_),
    .B(_1477_));
 sg13g2_o21ai_1 _2509_ (.B1(_1003_),
    .Y(_0169_),
    .A1(_0996_),
    .A2(_1473_));
 sg13g2_nand4_1 _2510_ (.B(_0167_),
    .C(_0168_),
    .A(_1482_),
    .Y(_0170_),
    .D(_0169_));
 sg13g2_nand3_1 _2511_ (.B(_1066_),
    .C(_1485_),
    .A(net742),
    .Y(_0171_));
 sg13g2_o21ai_1 _2512_ (.B1(_1007_),
    .Y(_0172_),
    .A1(net660),
    .A2(net709));
 sg13g2_a22oi_1 _2513_ (.Y(_0173_),
    .B1(_0172_),
    .B2(net727),
    .A2(_1082_),
    .A1(net743));
 sg13g2_nand2_1 _2514_ (.Y(_0174_),
    .A(_0171_),
    .B(_0173_));
 sg13g2_o21ai_1 _2515_ (.B1(_1092_),
    .Y(_0175_),
    .A1(net638),
    .A2(_1473_));
 sg13g2_a21oi_1 _2516_ (.A1(_1016_),
    .A2(_0117_),
    .Y(_0176_),
    .B1(net667));
 sg13g2_o21ai_1 _2517_ (.B1(_0176_),
    .Y(_0177_),
    .A1(net713),
    .A2(_0175_));
 sg13g2_a221oi_1 _2518_ (.B2(net675),
    .C1(_0177_),
    .B1(_0174_),
    .A1(net713),
    .Y(_0178_),
    .A2(_0170_));
 sg13g2_or3_1 _2519_ (.A(net619),
    .B(_0165_),
    .C(_0178_),
    .X(_0179_));
 sg13g2_a22oi_1 _2520_ (.Y(_0180_),
    .B1(_1437_),
    .B2(_1019_),
    .A2(_1435_),
    .A1(_1171_));
 sg13g2_o21ai_1 _2521_ (.B1(net666),
    .Y(_0181_),
    .A1(net718),
    .A2(_0180_));
 sg13g2_and3_1 _2522_ (.X(_0182_),
    .A(net751),
    .B(_1008_),
    .C(_1429_));
 sg13g2_a21oi_1 _2523_ (.A1(net756),
    .A2(_1437_),
    .Y(_0183_),
    .B1(_0182_));
 sg13g2_a221oi_1 _2524_ (.B2(net756),
    .C1(_0182_),
    .B1(_1437_),
    .A1(net658),
    .Y(_0184_),
    .A2(_1044_));
 sg13g2_o21ai_1 _2525_ (.B1(_1432_),
    .Y(_0185_),
    .A1(net734),
    .A2(_0184_));
 sg13g2_a21o_1 _2526_ (.A2(_0185_),
    .A1(net718),
    .B1(_0181_),
    .X(_0186_));
 sg13g2_a221oi_1 _2527_ (.B2(net639),
    .C1(net652),
    .B1(net644),
    .A1(net750),
    .Y(_0187_),
    .A2(net733));
 sg13g2_nor2_1 _2528_ (.A(net722),
    .B(_0187_),
    .Y(_0188_));
 sg13g2_nor4_2 _2529_ (.A(_0937_),
    .B(_0939_),
    .C(_0949_),
    .Y(_0189_),
    .D(net768));
 sg13g2_nor4_1 _2530_ (.A(net652),
    .B(net644),
    .C(net700),
    .D(_0189_),
    .Y(_0190_));
 sg13g2_or3_1 _2531_ (.A(net722),
    .B(_0187_),
    .C(_0190_),
    .X(_0191_));
 sg13g2_nand3_1 _2532_ (.B(_1458_),
    .C(_0191_),
    .A(net669),
    .Y(_0192_));
 sg13g2_and2_1 _2533_ (.A(net619),
    .B(_0192_),
    .X(_0193_));
 sg13g2_a21oi_1 _2534_ (.A1(_0186_),
    .A2(_0193_),
    .Y(_0194_),
    .B1(_1028_));
 sg13g2_a22oi_1 _2535_ (.Y(_0195_),
    .B1(_0149_),
    .B2(_1065_),
    .A2(_1104_),
    .A1(_0989_));
 sg13g2_nand4_1 _2536_ (.B(_1204_),
    .C(_1426_),
    .A(_1123_),
    .Y(_0196_),
    .D(_0195_));
 sg13g2_o21ai_1 _2537_ (.B1(net727),
    .Y(_0197_),
    .A1(_1099_),
    .A2(_1134_));
 sg13g2_nand4_1 _2538_ (.B(_1194_),
    .C(_1423_),
    .A(net675),
    .Y(_0198_),
    .D(_0197_));
 sg13g2_nor2_1 _2539_ (.A(_1017_),
    .B(_0159_),
    .Y(_0199_));
 sg13g2_o21ai_1 _2540_ (.B1(_0199_),
    .Y(_0200_),
    .A1(net743),
    .A2(_1102_));
 sg13g2_and4_1 _2541_ (.A(net663),
    .B(_0196_),
    .C(_0198_),
    .D(_0200_),
    .X(_0201_));
 sg13g2_nand3_1 _2542_ (.B(net640),
    .C(_1047_),
    .A(net749),
    .Y(_0202_));
 sg13g2_a21oi_1 _2543_ (.A1(_1431_),
    .A2(_0202_),
    .Y(_0203_),
    .B1(net729));
 sg13g2_nand2_1 _2544_ (.Y(_0204_),
    .A(_0997_),
    .B(_1054_));
 sg13g2_a21oi_1 _2545_ (.A1(_0997_),
    .A2(_1054_),
    .Y(_0205_),
    .B1(_1071_));
 sg13g2_o21ai_1 _2546_ (.B1(_1146_),
    .Y(_0206_),
    .A1(_0996_),
    .A2(net636));
 sg13g2_o21ai_1 _2547_ (.B1(_0206_),
    .Y(_0207_),
    .A1(_1155_),
    .A2(_1446_));
 sg13g2_or2_1 _2548_ (.X(_0208_),
    .B(_1060_),
    .A(net634));
 sg13g2_nor3_1 _2549_ (.A(net712),
    .B(_0203_),
    .C(_0207_),
    .Y(_0209_));
 sg13g2_a22oi_1 _2550_ (.Y(_0210_),
    .B1(_1214_),
    .B2(_0208_),
    .A2(_1212_),
    .A1(_1142_));
 sg13g2_a21oi_1 _2551_ (.A1(_1034_),
    .A2(_1130_),
    .Y(_0211_),
    .B1(net769));
 sg13g2_o21ai_1 _2552_ (.B1(net703),
    .Y(_0212_),
    .A1(_1217_),
    .A2(_0211_));
 sg13g2_and2_1 _2553_ (.A(net736),
    .B(_1450_),
    .X(_0213_));
 sg13g2_a21oi_2 _2554_ (.B1(net637),
    .Y(_0214_),
    .A2(net630),
    .A1(net660));
 sg13g2_o21ai_1 _2555_ (.B1(net706),
    .Y(_0215_),
    .A1(net764),
    .A2(_1030_));
 sg13g2_nor2_1 _2556_ (.A(_0214_),
    .B(_0215_),
    .Y(_0216_));
 sg13g2_nor4_1 _2557_ (.A(net721),
    .B(_1219_),
    .C(_0213_),
    .D(_0216_),
    .Y(_0217_));
 sg13g2_a221oi_1 _2558_ (.B2(_0217_),
    .C1(net663),
    .B1(_0212_),
    .A1(_0209_),
    .Y(_0218_),
    .A2(_0210_));
 sg13g2_o21ai_1 _2559_ (.B1(net619),
    .Y(_0219_),
    .A1(_0201_),
    .A2(_0218_));
 sg13g2_nand3_1 _2560_ (.B(net648),
    .C(_1249_),
    .A(net659),
    .Y(_0220_));
 sg13g2_and4_1 _2561_ (.A(net717),
    .B(_1010_),
    .C(_0126_),
    .D(_0220_),
    .X(_0221_));
 sg13g2_a221oi_1 _2562_ (.B2(net674),
    .C1(_1143_),
    .B1(_0136_),
    .A1(_1016_),
    .Y(_0222_),
    .A2(_0130_));
 sg13g2_a221oi_1 _2563_ (.B2(net699),
    .C1(_0222_),
    .B1(_0138_),
    .A1(net706),
    .Y(_0223_),
    .A2(_0137_));
 sg13g2_o21ai_1 _2564_ (.B1(net669),
    .Y(_0224_),
    .A1(_0221_),
    .A2(_0223_));
 sg13g2_a21oi_1 _2565_ (.A1(_1449_),
    .A2(_1456_),
    .Y(_0225_),
    .B1(net757));
 sg13g2_nor2_1 _2566_ (.A(net742),
    .B(_0126_),
    .Y(_0226_));
 sg13g2_o21ai_1 _2567_ (.B1(net674),
    .Y(_0227_),
    .A1(_0225_),
    .A2(_0226_));
 sg13g2_o21ai_1 _2568_ (.B1(net665),
    .Y(_0228_),
    .A1(_1023_),
    .A2(_0124_));
 sg13g2_a21oi_1 _2569_ (.A1(net673),
    .A2(_1455_),
    .Y(_0229_),
    .B1(_0228_));
 sg13g2_a21oi_1 _2570_ (.A1(_0227_),
    .A2(_0229_),
    .Y(_0230_),
    .B1(net619));
 sg13g2_a21oi_1 _2571_ (.A1(_0224_),
    .A2(_0230_),
    .Y(_0231_),
    .B1(net622));
 sg13g2_a221oi_1 _2572_ (.B2(_0231_),
    .C1(_1117_),
    .B1(_0219_),
    .A1(_0179_),
    .Y(_0232_),
    .A2(_0194_));
 sg13g2_nor2_1 _2573_ (.A(_0887_),
    .B(_0232_),
    .Y(_0233_));
 sg13g2_nor3_1 _2574_ (.A(net764),
    .B(_1106_),
    .C(_1429_),
    .Y(_0234_));
 sg13g2_or3_1 _2575_ (.A(net739),
    .B(_0150_),
    .C(_0234_),
    .X(_0235_));
 sg13g2_a21oi_1 _2576_ (.A1(net756),
    .A2(_1095_),
    .Y(_0236_),
    .B1(net720));
 sg13g2_nand3_1 _2577_ (.B(_0235_),
    .C(_0236_),
    .A(_0195_),
    .Y(_0237_));
 sg13g2_or3_1 _2578_ (.A(net773),
    .B(_1106_),
    .C(_1429_),
    .X(_0238_));
 sg13g2_a21oi_1 _2579_ (.A1(net704),
    .A2(_0238_),
    .Y(_0239_),
    .B1(_0237_));
 sg13g2_o21ai_1 _2580_ (.B1(_1016_),
    .Y(_0240_),
    .A1(_1281_),
    .A2(_1326_));
 sg13g2_o21ai_1 _2581_ (.B1(net748),
    .Y(_0241_),
    .A1(_1087_),
    .A2(_1134_));
 sg13g2_nand2_1 _2582_ (.Y(_0242_),
    .A(net675),
    .B(_0241_));
 sg13g2_a21oi_1 _2583_ (.A1(_0155_),
    .A2(_0160_),
    .Y(_0243_),
    .B1(_0993_));
 sg13g2_o21ai_1 _2584_ (.B1(_1033_),
    .Y(_0244_),
    .A1(net764),
    .A2(_0160_));
 sg13g2_a221oi_1 _2585_ (.B2(net698),
    .C1(_0243_),
    .B1(_0244_),
    .A1(_0240_),
    .Y(_0245_),
    .A2(_0242_));
 sg13g2_o21ai_1 _2586_ (.B1(net663),
    .Y(_0246_),
    .A1(_0239_),
    .A2(_0245_));
 sg13g2_nand3_1 _2587_ (.B(net640),
    .C(_1047_),
    .A(net698),
    .Y(_0247_));
 sg13g2_nand2_1 _2588_ (.Y(_0248_),
    .A(net640),
    .B(net636));
 sg13g2_nand4_1 _2589_ (.B(_1163_),
    .C(_0247_),
    .A(net721),
    .Y(_0249_),
    .D(_0248_));
 sg13g2_a21oi_1 _2590_ (.A1(_1092_),
    .A2(_0204_),
    .Y(_0250_),
    .B1(_0249_));
 sg13g2_o21ai_1 _2591_ (.B1(_1033_),
    .Y(_0251_),
    .A1(net769),
    .A2(_1130_));
 sg13g2_o21ai_1 _2592_ (.B1(net712),
    .Y(_0252_),
    .A1(_0993_),
    .A2(_0214_));
 sg13g2_o21ai_1 _2593_ (.B1(net765),
    .Y(_0253_),
    .A1(_0996_),
    .A2(net634));
 sg13g2_nand3_1 _2594_ (.B(_1383_),
    .C(_0253_),
    .A(net754),
    .Y(_0254_));
 sg13g2_a21oi_1 _2595_ (.A1(net748),
    .A2(_0214_),
    .Y(_0255_),
    .B1(net728));
 sg13g2_a221oi_1 _2596_ (.B2(_0255_),
    .C1(_0252_),
    .B1(_0254_),
    .A1(net703),
    .Y(_0256_),
    .A2(_0251_));
 sg13g2_o21ai_1 _2597_ (.B1(_0910_),
    .Y(_0257_),
    .A1(_0250_),
    .A2(_0256_));
 sg13g2_and2_1 _2598_ (.A(net623),
    .B(_0257_),
    .X(_0258_));
 sg13g2_or2_1 _2599_ (.X(_0259_),
    .B(_1196_),
    .A(_1164_));
 sg13g2_a22oi_1 _2600_ (.Y(_0260_),
    .B1(_0259_),
    .B2(_1066_),
    .A2(_1437_),
    .A1(net751));
 sg13g2_nor2_1 _2601_ (.A(_1021_),
    .B(_0260_),
    .Y(_0261_));
 sg13g2_a221oi_1 _2602_ (.B2(_0202_),
    .C1(net725),
    .B1(_1431_),
    .A1(net740),
    .Y(_0262_),
    .A2(_1430_));
 sg13g2_o21ai_1 _2603_ (.B1(net666),
    .Y(_0263_),
    .A1(_1017_),
    .A2(_0183_));
 sg13g2_nor3_1 _2604_ (.A(_0261_),
    .B(_0262_),
    .C(_0263_),
    .Y(_0264_));
 sg13g2_a22oi_1 _2605_ (.Y(_0265_),
    .B1(_1057_),
    .B2(_0959_),
    .A2(_0960_),
    .A1(net656));
 sg13g2_nor2_1 _2606_ (.A(net715),
    .B(net700),
    .Y(_0266_));
 sg13g2_a21oi_1 _2607_ (.A1(_1165_),
    .A2(_0265_),
    .Y(_0267_),
    .B1(_1014_));
 sg13g2_o21ai_1 _2608_ (.B1(net671),
    .Y(_0268_),
    .A1(_1144_),
    .A2(_1376_));
 sg13g2_a221oi_1 _2609_ (.B2(_1144_),
    .C1(_0268_),
    .B1(_0267_),
    .A1(_1014_),
    .Y(_0269_),
    .A2(_0259_));
 sg13g2_or2_1 _2610_ (.X(_0270_),
    .B(_0269_),
    .A(net625));
 sg13g2_o21ai_1 _2611_ (.B1(net619),
    .Y(_0271_),
    .A1(_0264_),
    .A2(_0270_));
 sg13g2_a21o_1 _2612_ (.A2(_0258_),
    .A1(_0246_),
    .B1(_0271_),
    .X(_0272_));
 sg13g2_and2_1 _2613_ (.A(_0983_),
    .B(net643),
    .X(_0273_));
 sg13g2_a21oi_1 _2614_ (.A1(_1088_),
    .A2(_0273_),
    .Y(_0274_),
    .B1(net748));
 sg13g2_o21ai_1 _2615_ (.B1(net730),
    .Y(_0275_),
    .A1(_0990_),
    .A2(_0208_));
 sg13g2_nor2_1 _2616_ (.A(_0274_),
    .B(_0275_),
    .Y(_0276_));
 sg13g2_a21oi_1 _2617_ (.A1(net770),
    .A2(_0273_),
    .Y(_0277_),
    .B1(_1119_));
 sg13g2_nor3_1 _2618_ (.A(_1019_),
    .B(_1057_),
    .C(_0277_),
    .Y(_0278_));
 sg13g2_nand2_1 _2619_ (.Y(_0279_),
    .A(net678),
    .B(net764));
 sg13g2_nand2_1 _2620_ (.Y(_0280_),
    .A(_1003_),
    .B(_0273_));
 sg13g2_a21oi_1 _2621_ (.A1(_1099_),
    .A2(_0279_),
    .Y(_0281_),
    .B1(_0280_));
 sg13g2_nor4_1 _2622_ (.A(net720),
    .B(_0276_),
    .C(_0278_),
    .D(_0281_),
    .Y(_0282_));
 sg13g2_o21ai_1 _2623_ (.B1(net750),
    .Y(_0283_),
    .A1(net707),
    .A2(net682));
 sg13g2_nand2_1 _2624_ (.Y(_0284_),
    .A(_1033_),
    .B(_0283_));
 sg13g2_a21oi_1 _2625_ (.A1(_1102_),
    .A2(_0284_),
    .Y(_0285_),
    .B1(_1017_));
 sg13g2_nor3_1 _2626_ (.A(net768),
    .B(net641),
    .C(net628),
    .Y(_0286_));
 sg13g2_nor2_1 _2627_ (.A(_1021_),
    .B(_0286_),
    .Y(_0287_));
 sg13g2_nand2_1 _2628_ (.Y(_0288_),
    .A(_0983_),
    .B(_1089_));
 sg13g2_nand2b_1 _2629_ (.Y(_0289_),
    .B(_1034_),
    .A_N(_0288_));
 sg13g2_and2_1 _2630_ (.A(_1014_),
    .B(_0289_),
    .X(_0290_));
 sg13g2_a21oi_1 _2631_ (.A1(_0238_),
    .A2(_0287_),
    .Y(_0291_),
    .B1(net663));
 sg13g2_o21ai_1 _2632_ (.B1(_0291_),
    .Y(_0292_),
    .A1(_1023_),
    .A2(_0234_));
 sg13g2_nor4_1 _2633_ (.A(_0282_),
    .B(_0285_),
    .C(_0290_),
    .D(_0292_),
    .Y(_0293_));
 sg13g2_a21oi_1 _2634_ (.A1(net774),
    .A2(_0997_),
    .Y(_0294_),
    .B1(_1401_));
 sg13g2_a22oi_1 _2635_ (.Y(_0295_),
    .B1(_0973_),
    .B2(net658),
    .A2(net647),
    .A1(_0951_));
 sg13g2_a21oi_1 _2636_ (.A1(net699),
    .A2(_1031_),
    .Y(_0296_),
    .B1(_1144_));
 sg13g2_o21ai_1 _2637_ (.B1(_0296_),
    .Y(_0297_),
    .A1(net638),
    .A2(_0288_));
 sg13g2_o21ai_1 _2638_ (.B1(_0266_),
    .Y(_0298_),
    .A1(_0982_),
    .A2(_0294_));
 sg13g2_nand3b_1 _2639_ (.B(_0997_),
    .C(net700),
    .Y(_0299_),
    .A_N(_0982_));
 sg13g2_nor3_1 _2640_ (.A(net772),
    .B(_1047_),
    .C(_1060_),
    .Y(_0300_));
 sg13g2_o21ai_1 _2641_ (.B1(net703),
    .Y(_0301_),
    .A1(_0295_),
    .A2(_0300_));
 sg13g2_nand3_1 _2642_ (.B(_0299_),
    .C(_0301_),
    .A(net715),
    .Y(_0302_));
 sg13g2_nand3_1 _2643_ (.B(_0298_),
    .C(_0302_),
    .A(_0297_),
    .Y(_0303_));
 sg13g2_o21ai_1 _2644_ (.B1(_1029_),
    .Y(_0304_),
    .A1(net667),
    .A2(_0303_));
 sg13g2_nor3_1 _2645_ (.A(_0978_),
    .B(_1164_),
    .C(_1196_),
    .Y(_0305_));
 sg13g2_nand2_1 _2646_ (.Y(_0306_),
    .A(net647),
    .B(_1039_));
 sg13g2_o21ai_1 _2647_ (.B1(net740),
    .Y(_0307_),
    .A1(_0960_),
    .A2(_0283_));
 sg13g2_a221oi_1 _2648_ (.B2(_1166_),
    .C1(_0305_),
    .B1(_0307_),
    .A1(net756),
    .Y(_0308_),
    .A2(_0306_));
 sg13g2_nand2_1 _2649_ (.Y(_0309_),
    .A(_1166_),
    .B(_0265_));
 sg13g2_a21oi_1 _2650_ (.A1(net732),
    .A2(_0309_),
    .Y(_0310_),
    .B1(_0308_));
 sg13g2_o21ai_1 _2651_ (.B1(net674),
    .Y(_0311_),
    .A1(net756),
    .A2(_1039_));
 sg13g2_nor2_1 _2652_ (.A(_0295_),
    .B(_0311_),
    .Y(_0312_));
 sg13g2_o21ai_1 _2653_ (.B1(net671),
    .Y(_0313_),
    .A1(_1017_),
    .A2(_0306_));
 sg13g2_nor2_1 _2654_ (.A(_0312_),
    .B(_0313_),
    .Y(_0314_));
 sg13g2_o21ai_1 _2655_ (.B1(_0314_),
    .Y(_0315_),
    .A1(net725),
    .A2(_0310_));
 sg13g2_o21ai_1 _2656_ (.B1(net666),
    .Y(_0316_),
    .A1(net674),
    .A2(_1376_));
 sg13g2_a21oi_1 _2657_ (.A1(net674),
    .A2(_0309_),
    .Y(_0317_),
    .B1(_0316_));
 sg13g2_nor2_1 _2658_ (.A(net622),
    .B(_0317_),
    .Y(_0318_));
 sg13g2_a21oi_1 _2659_ (.A1(_0315_),
    .A2(_0318_),
    .Y(_0319_),
    .B1(net619));
 sg13g2_o21ai_1 _2660_ (.B1(_0319_),
    .Y(_0320_),
    .A1(_0293_),
    .A2(_0304_));
 sg13g2_nand3_1 _2661_ (.B(_0272_),
    .C(_0320_),
    .A(_1118_),
    .Y(_0321_));
 sg13g2_nand4_1 _2662_ (.B(_0195_),
    .C(_0235_),
    .A(_1122_),
    .Y(_0322_),
    .D(_0236_));
 sg13g2_o21ai_1 _2663_ (.B1(_0199_),
    .Y(_0323_),
    .A1(_1281_),
    .A2(_1326_));
 sg13g2_nand3_1 _2664_ (.B(_1423_),
    .C(_0241_),
    .A(net675),
    .Y(_0324_));
 sg13g2_nand4_1 _2665_ (.B(_0322_),
    .C(_0323_),
    .A(net663),
    .Y(_0325_),
    .D(_0324_));
 sg13g2_o21ai_1 _2666_ (.B1(net771),
    .Y(_0326_),
    .A1(net634),
    .A2(_1060_));
 sg13g2_a21oi_1 _2667_ (.A1(_0253_),
    .A2(_0326_),
    .Y(_0327_),
    .B1(net700));
 sg13g2_nor3_1 _2668_ (.A(net771),
    .B(net731),
    .C(_1446_),
    .Y(_0328_));
 sg13g2_nor4_1 _2669_ (.A(_0205_),
    .B(_0249_),
    .C(_0327_),
    .D(_0328_),
    .Y(_0329_));
 sg13g2_o21ai_1 _2670_ (.B1(_1066_),
    .Y(_0330_),
    .A1(net637),
    .A2(net634));
 sg13g2_o21ai_1 _2671_ (.B1(_0330_),
    .Y(_0331_),
    .A1(net764),
    .A2(_0214_));
 sg13g2_a21o_1 _2672_ (.A2(_1142_),
    .A1(net736),
    .B1(_1003_),
    .X(_0332_));
 sg13g2_a221oi_1 _2673_ (.B2(_0332_),
    .C1(_0252_),
    .B1(_0331_),
    .A1(net703),
    .Y(_0333_),
    .A2(_0251_));
 sg13g2_or2_1 _2674_ (.X(_0334_),
    .B(_0333_),
    .A(_0329_));
 sg13g2_o21ai_1 _2675_ (.B1(_0325_),
    .Y(_0335_),
    .A1(net663),
    .A2(_0334_));
 sg13g2_o21ai_1 _2676_ (.B1(_1430_),
    .Y(_0336_),
    .A1(net699),
    .A2(_1163_));
 sg13g2_a21oi_1 _2677_ (.A1(net718),
    .A2(_0336_),
    .Y(_0337_),
    .B1(_0181_));
 sg13g2_o21ai_1 _2678_ (.B1(_0188_),
    .Y(_0338_),
    .A1(net700),
    .A2(_1435_));
 sg13g2_nand3_1 _2679_ (.B(net627),
    .C(_1250_),
    .A(_1042_),
    .Y(_0339_));
 sg13g2_nand4_1 _2680_ (.B(_1458_),
    .C(_0338_),
    .A(net670),
    .Y(_0340_),
    .D(_0339_));
 sg13g2_nor2_1 _2681_ (.A(net625),
    .B(_0337_),
    .Y(_0341_));
 sg13g2_a221oi_1 _2682_ (.B2(_0341_),
    .C1(net620),
    .B1(_0340_),
    .A1(net625),
    .Y(_0342_),
    .A2(_0335_));
 sg13g2_a22oi_1 _2683_ (.Y(_0343_),
    .B1(_0158_),
    .B2(net742),
    .A2(_1095_),
    .A1(net763));
 sg13g2_nor2_1 _2684_ (.A(_0162_),
    .B(_0343_),
    .Y(_0344_));
 sg13g2_a21oi_1 _2685_ (.A1(net711),
    .A2(net678),
    .Y(_0345_),
    .B1(_0159_));
 sg13g2_o21ai_1 _2686_ (.B1(_1468_),
    .Y(_0346_),
    .A1(_0993_),
    .A2(_0345_));
 sg13g2_o21ai_1 _2687_ (.B1(net712),
    .Y(_0347_),
    .A1(_0344_),
    .A2(_0346_));
 sg13g2_o21ai_1 _2688_ (.B1(_1016_),
    .Y(_0348_),
    .A1(_1095_),
    .A2(_0152_));
 sg13g2_nand2_1 _2689_ (.Y(_0349_),
    .A(_1022_),
    .B(_1111_));
 sg13g2_nand4_1 _2690_ (.B(_0347_),
    .C(_0348_),
    .A(_0291_),
    .Y(_0350_),
    .D(_0349_));
 sg13g2_nand2_1 _2691_ (.Y(_0351_),
    .A(net698),
    .B(_1485_));
 sg13g2_o21ai_1 _2692_ (.B1(_0172_),
    .Y(_0352_),
    .A1(_1003_),
    .A2(_1154_));
 sg13g2_nand4_1 _2693_ (.B(_0175_),
    .C(_0351_),
    .A(net721),
    .Y(_0353_),
    .D(_0352_));
 sg13g2_o21ai_1 _2694_ (.B1(_1341_),
    .Y(_0354_),
    .A1(_0996_),
    .A2(_1473_));
 sg13g2_o21ai_1 _2695_ (.B1(_1249_),
    .Y(_0355_),
    .A1(_1060_),
    .A2(_1473_));
 sg13g2_o21ai_1 _2696_ (.B1(_1092_),
    .Y(_0356_),
    .A1(_0996_),
    .A2(_1477_));
 sg13g2_nand4_1 _2697_ (.B(_0354_),
    .C(_0355_),
    .A(net713),
    .Y(_0357_),
    .D(_0356_));
 sg13g2_a21oi_2 _2698_ (.B1(net667),
    .Y(_0358_),
    .A2(_0357_),
    .A1(_0353_));
 sg13g2_nor2_1 _2699_ (.A(net623),
    .B(_0358_),
    .Y(_0359_));
 sg13g2_a221oi_1 _2700_ (.B2(net682),
    .C1(net740),
    .B1(net627),
    .A1(net641),
    .Y(_0360_),
    .A2(net639));
 sg13g2_nand3_1 _2701_ (.B(_1456_),
    .C(_0126_),
    .A(net741),
    .Y(_0361_));
 sg13g2_nor3_1 _2702_ (.A(net717),
    .B(_1212_),
    .C(_0360_),
    .Y(_0362_));
 sg13g2_a22oi_1 _2703_ (.Y(_0363_),
    .B1(_0361_),
    .B2(_0362_),
    .A2(_1455_),
    .A1(_1144_));
 sg13g2_nand2_1 _2704_ (.Y(_0364_),
    .A(net665),
    .B(_0363_));
 sg13g2_nand3_1 _2705_ (.B(_0126_),
    .C(_0220_),
    .A(_1456_),
    .Y(_0365_));
 sg13g2_a21oi_1 _2706_ (.A1(_0971_),
    .A2(_1213_),
    .Y(_0366_),
    .B1(net724));
 sg13g2_a21oi_1 _2707_ (.A1(net661),
    .A2(_0962_),
    .Y(_0367_),
    .B1(_0971_));
 sg13g2_o21ai_1 _2708_ (.B1(net669),
    .Y(_0368_),
    .A1(_1144_),
    .A2(_0136_));
 sg13g2_a221oi_1 _2709_ (.B2(_1016_),
    .C1(_0368_),
    .B1(_0367_),
    .A1(_0365_),
    .Y(_0369_),
    .A2(_0366_));
 sg13g2_nor2_1 _2710_ (.A(_1029_),
    .B(_0369_),
    .Y(_0370_));
 sg13g2_a221oi_1 _2711_ (.B2(_0370_),
    .C1(_0909_),
    .B1(_0364_),
    .A1(_0350_),
    .Y(_0371_),
    .A2(_0359_));
 sg13g2_or3_1 _2712_ (.A(_1118_),
    .B(_0342_),
    .C(_0371_),
    .X(_0372_));
 sg13g2_nand3_1 _2713_ (.B(_0321_),
    .C(_0372_),
    .A(_0887_),
    .Y(_0373_));
 sg13g2_a21oi_1 _2714_ (.A1(_0147_),
    .A2(_0233_),
    .Y(_0374_),
    .B1(_1276_));
 sg13g2_nor2b_1 _2715_ (.A(net792),
    .B_N(net777),
    .Y(_0375_));
 sg13g2_o21ai_1 _2716_ (.B1(_0907_),
    .Y(_0376_),
    .A1(\logo_top[6] ),
    .A2(_0742_));
 sg13g2_nand2_1 _2717_ (.Y(_0377_),
    .A(_0375_),
    .B(_0376_));
 sg13g2_nor2b_1 _2718_ (.A(\pix_x[8] ),
    .B_N(\logo_left[8] ),
    .Y(_0378_));
 sg13g2_xor2_1 _2719_ (.B(\pix_x[8] ),
    .A(\logo_left[8] ),
    .X(_0379_));
 sg13g2_nor2b_1 _2720_ (.A(\logo_left[7] ),
    .B_N(\pix_x[7] ),
    .Y(_0380_));
 sg13g2_and2_1 _2721_ (.A(_0917_),
    .B(net697),
    .X(_0381_));
 sg13g2_nor2b_1 _2722_ (.A(\pix_x[7] ),
    .B_N(net798),
    .Y(_0382_));
 sg13g2_nor3_1 _2723_ (.A(_0380_),
    .B(_0381_),
    .C(_0382_),
    .Y(_0383_));
 sg13g2_o21ai_1 _2724_ (.B1(_0379_),
    .Y(_0384_),
    .A1(_0380_),
    .A2(_0383_));
 sg13g2_a21o_1 _2725_ (.A2(_0382_),
    .A1(_0379_),
    .B1(_0380_),
    .X(_0385_));
 sg13g2_a21oi_1 _2726_ (.A1(_0381_),
    .A2(_0385_),
    .Y(_0386_),
    .B1(_0383_));
 sg13g2_xnor2_1 _2727_ (.Y(_0387_),
    .A(net791),
    .B(\pix_y[9] ));
 sg13g2_nor2_1 _2728_ (.A(_0727_),
    .B(\pix_y[8] ),
    .Y(_0388_));
 sg13g2_xnor2_1 _2729_ (.Y(_0389_),
    .A(_0387_),
    .B(_0388_));
 sg13g2_xnor2_1 _2730_ (.Y(_0390_),
    .A(\logo_left[9] ),
    .B(\pix_x[9] ));
 sg13g2_xnor2_1 _2731_ (.Y(_0391_),
    .A(_0378_),
    .B(_0390_));
 sg13g2_nor3_1 _2732_ (.A(_0386_),
    .B(_0389_),
    .C(_0391_),
    .Y(_0392_));
 sg13g2_nand2b_1 _2733_ (.Y(_0393_),
    .B(net792),
    .A_N(net777));
 sg13g2_o21ai_1 _2734_ (.B1(_0387_),
    .Y(_0394_),
    .A1(\logo_top[8] ),
    .A2(_0744_));
 sg13g2_a21o_1 _2735_ (.A2(_0393_),
    .A1(_0376_),
    .B1(_0375_),
    .X(_0395_));
 sg13g2_nor2_1 _2736_ (.A(_0376_),
    .B(_0393_),
    .Y(_0396_));
 sg13g2_mux2_1 _2737_ (.A0(_0395_),
    .A1(_0396_),
    .S(_0394_),
    .X(_0397_));
 sg13g2_nand4_1 _2738_ (.B(_0384_),
    .C(_0392_),
    .A(_0377_),
    .Y(_0398_),
    .D(_0397_));
 sg13g2_nand2b_1 _2739_ (.Y(_0399_),
    .B(_0398_),
    .A_N(net1));
 sg13g2_nor2_1 _2740_ (.A(net805),
    .B(\pix_y[9] ),
    .Y(_0400_));
 sg13g2_o21ai_1 _2741_ (.B1(\pix_x[9] ),
    .Y(_0401_),
    .A1(\pix_x[8] ),
    .A2(\pix_x[7] ));
 sg13g2_nand4_1 _2742_ (.B(_0399_),
    .C(_0400_),
    .A(_0764_),
    .Y(_0402_),
    .D(_0401_));
 sg13g2_a221oi_1 _2743_ (.B2(_0374_),
    .C1(_0402_),
    .B1(_0373_),
    .A1(_1274_),
    .Y(_0403_),
    .A2(_1422_));
 sg13g2_nand2b_1 _2744_ (.Y(_0404_),
    .B(net668),
    .A_N(_0008_));
 sg13g2_xnor2_1 _2745_ (.Y(_0405_),
    .A(net799),
    .B(net668));
 sg13g2_o21ai_1 _2746_ (.B1(_0404_),
    .Y(_0406_),
    .A1(net711),
    .A2(_0405_));
 sg13g2_nor2_1 _2747_ (.A(_0734_),
    .B(net624),
    .Y(_0407_));
 sg13g2_xnor2_1 _2748_ (.Y(_0408_),
    .A(\logo_left[5] ),
    .B(net624));
 sg13g2_xnor2_1 _2749_ (.Y(_0409_),
    .A(net682),
    .B(_0408_));
 sg13g2_xnor2_1 _2750_ (.Y(_0410_),
    .A(net707),
    .B(_0405_));
 sg13g2_nand2_1 _2751_ (.Y(_0411_),
    .A(\logo_left[3] ),
    .B(net725));
 sg13g2_xnor2_1 _2752_ (.Y(_0412_),
    .A(\logo_left[3] ),
    .B(net725));
 sg13g2_o21ai_1 _2753_ (.B1(_0411_),
    .Y(_0413_),
    .A1(_0948_),
    .A2(_0412_));
 sg13g2_nand2_1 _2754_ (.Y(_0414_),
    .A(_0410_),
    .B(_0413_));
 sg13g2_nand2_1 _2755_ (.Y(_0415_),
    .A(_0007_),
    .B(_1275_));
 sg13g2_xnor2_1 _2756_ (.Y(_0416_),
    .A(_0949_),
    .B(_0412_));
 sg13g2_xnor2_1 _2757_ (.Y(_0417_),
    .A(\pix_x[2] ),
    .B(_0924_));
 sg13g2_nor2_1 _2758_ (.A(net734),
    .B(_0417_),
    .Y(_0418_));
 sg13g2_xnor2_1 _2759_ (.Y(_0419_),
    .A(_0415_),
    .B(_0416_));
 sg13g2_nor3_1 _2760_ (.A(net734),
    .B(_0417_),
    .C(_0419_),
    .Y(_0420_));
 sg13g2_a21oi_1 _2761_ (.A1(_0415_),
    .A2(_0416_),
    .Y(_0421_),
    .B1(_0420_));
 sg13g2_xor2_1 _2762_ (.B(_0413_),
    .A(_0410_),
    .X(_0422_));
 sg13g2_nand2b_1 _2763_ (.Y(_0423_),
    .B(_0422_),
    .A_N(_0421_));
 sg13g2_xnor2_1 _2764_ (.Y(_0424_),
    .A(_0406_),
    .B(_0409_));
 sg13g2_a21oi_2 _2765_ (.B1(_0424_),
    .Y(_0425_),
    .A2(_0423_),
    .A1(_0414_));
 sg13g2_a21oi_1 _2766_ (.A1(_0406_),
    .A2(_0409_),
    .Y(_0426_),
    .B1(_0425_));
 sg13g2_a21oi_1 _2767_ (.A1(net684),
    .A2(_0408_),
    .Y(_0427_),
    .B1(_0407_));
 sg13g2_xnor2_1 _2768_ (.Y(_0428_),
    .A(\logo_left[6] ),
    .B(net662));
 sg13g2_xnor2_1 _2769_ (.Y(_0429_),
    .A(_0908_),
    .B(_0428_));
 sg13g2_xnor2_1 _2770_ (.Y(_0430_),
    .A(_0427_),
    .B(_0429_));
 sg13g2_xnor2_1 _2771_ (.Y(_0431_),
    .A(_0426_),
    .B(_0430_));
 sg13g2_nand2_1 _2772_ (.Y(_0432_),
    .A(net2),
    .B(net232));
 sg13g2_o21ai_1 _2773_ (.B1(_0432_),
    .Y(_0433_),
    .A1(net2),
    .A2(_0431_));
 sg13g2_and2_1 _2774_ (.A(_0403_),
    .B(_0433_),
    .X(_0022_));
 sg13g2_nand2b_1 _2775_ (.Y(_0434_),
    .B(net2),
    .A_N(net227));
 sg13g2_and2_1 _2776_ (.A(_0403_),
    .B(_0434_),
    .X(_0023_));
 sg13g2_nor2b_1 _2777_ (.A(\gamepad.driver.pmod_latch_prev ),
    .B_N(\gamepad.driver.pmod_latch_sync[1] ),
    .Y(_0435_));
 sg13g2_nor2_1 _2778_ (.A(net805),
    .B(net761),
    .Y(_0436_));
 sg13g2_a22oi_1 _2779_ (.Y(_0024_),
    .B1(net747),
    .B2(_0750_),
    .A2(net762),
    .A1(_0722_));
 sg13g2_a22oi_1 _2780_ (.Y(_0025_),
    .B1(net747),
    .B2(_0749_),
    .A2(net762),
    .A1(_0721_));
 sg13g2_a22oi_1 _2781_ (.Y(_0026_),
    .B1(net747),
    .B2(_0752_),
    .A2(net762),
    .A1(_0720_));
 sg13g2_a22oi_1 _2782_ (.Y(_0027_),
    .B1(net747),
    .B2(_0751_),
    .A2(net762),
    .A1(_0719_));
 sg13g2_a22oi_1 _2783_ (.Y(_0028_),
    .B1(net746),
    .B2(_0754_),
    .A2(net761),
    .A1(_0718_));
 sg13g2_a22oi_1 _2784_ (.Y(_0029_),
    .B1(net746),
    .B2(_0753_),
    .A2(net761),
    .A1(_0717_));
 sg13g2_a22oi_1 _2785_ (.Y(_0030_),
    .B1(net746),
    .B2(_0756_),
    .A2(net761),
    .A1(_0716_));
 sg13g2_a22oi_1 _2786_ (.Y(_0031_),
    .B1(net746),
    .B2(_0755_),
    .A2(net761),
    .A1(_0715_));
 sg13g2_a22oi_1 _2787_ (.Y(_0032_),
    .B1(net746),
    .B2(_0758_),
    .A2(net761),
    .A1(_0714_));
 sg13g2_a22oi_1 _2788_ (.Y(_0033_),
    .B1(net746),
    .B2(_0757_),
    .A2(net761),
    .A1(_0713_));
 sg13g2_a22oi_1 _2789_ (.Y(_0034_),
    .B1(net746),
    .B2(_0760_),
    .A2(net761),
    .A1(_0712_));
 sg13g2_a22oi_1 _2790_ (.Y(_0035_),
    .B1(net746),
    .B2(_0759_),
    .A2(net762),
    .A1(_0738_));
 sg13g2_nand2_1 _2791_ (.Y(_0437_),
    .A(net140),
    .B(_0786_));
 sg13g2_nand4_1 _2792_ (.B(\gamepad.decoder.data_reg[8] ),
    .C(\gamepad.decoder.data_reg[11] ),
    .A(\gamepad.decoder.data_reg[9] ),
    .Y(_0438_),
    .D(\gamepad.decoder.data_reg[10] ));
 sg13g2_nand4_1 _2793_ (.B(\gamepad.decoder.data_reg[4] ),
    .C(\gamepad.decoder.data_reg[7] ),
    .A(\gamepad.decoder.data_reg[5] ),
    .Y(_0439_),
    .D(\gamepad.decoder.data_reg[6] ));
 sg13g2_nand4_1 _2794_ (.B(\gamepad.decoder.data_reg[0] ),
    .C(\gamepad.decoder.data_reg[3] ),
    .A(\gamepad.decoder.data_reg[1] ),
    .Y(_0440_),
    .D(\gamepad.decoder.data_reg[2] ));
 sg13g2_or3_2 _2795_ (.A(_0438_),
    .B(_0439_),
    .C(_0440_),
    .X(_0441_));
 sg13g2_nand3_1 _2796_ (.B(_0787_),
    .C(_0441_),
    .A(\gamepad.decoder.data_reg[8] ),
    .Y(_0442_));
 sg13g2_a21oi_1 _2797_ (.A1(_0437_),
    .A2(_0442_),
    .Y(_0036_),
    .B1(net805));
 sg13g2_and3_1 _2798_ (.X(_0443_),
    .A(\pix_x[0] ),
    .B(net218),
    .C(\pix_x[1] ));
 sg13g2_and2_1 _2799_ (.A(net233),
    .B(_0443_),
    .X(_0444_));
 sg13g2_and2_1 _2800_ (.A(net241),
    .B(_0444_),
    .X(_0445_));
 sg13g2_nor4_1 _2801_ (.A(net803),
    .B(\pix_x[6] ),
    .C(\pix_x[7] ),
    .D(_0401_),
    .Y(_0446_));
 sg13g2_and2_2 _2802_ (.A(_0445_),
    .B(_0446_),
    .X(_0447_));
 sg13g2_nor2_1 _2803_ (.A(net804),
    .B(_0447_),
    .Y(_0448_));
 sg13g2_nand2b_1 _2804_ (.Y(_0449_),
    .B(net807),
    .A_N(_0447_));
 sg13g2_and2_1 _2805_ (.A(net127),
    .B(_0448_),
    .X(_0037_));
 sg13g2_xnor2_1 _2806_ (.Y(_0450_),
    .A(\pix_x[0] ),
    .B(net224));
 sg13g2_nor2_1 _2807_ (.A(net672),
    .B(net225),
    .Y(_0038_));
 sg13g2_a21oi_1 _2808_ (.A1(\pix_x[0] ),
    .A2(\pix_x[1] ),
    .Y(_0451_),
    .B1(net218));
 sg13g2_nor3_1 _2809_ (.A(net805),
    .B(_0443_),
    .C(net219),
    .Y(_0039_));
 sg13g2_o21ai_1 _2810_ (.B1(net807),
    .Y(_0452_),
    .A1(net233),
    .A2(_0443_));
 sg13g2_nor2_1 _2811_ (.A(_0444_),
    .B(net234),
    .Y(_0040_));
 sg13g2_o21ai_1 _2812_ (.B1(net807),
    .Y(_0453_),
    .A1(net241),
    .A2(_0444_));
 sg13g2_nor2_1 _2813_ (.A(_0445_),
    .B(_0453_),
    .Y(_0041_));
 sg13g2_and2_1 _2814_ (.A(net803),
    .B(_0445_),
    .X(_0454_));
 sg13g2_nor2_1 _2815_ (.A(net803),
    .B(_0445_),
    .Y(_0455_));
 sg13g2_nor3_1 _2816_ (.A(net672),
    .B(_0454_),
    .C(_0455_),
    .Y(_0042_));
 sg13g2_nor2_1 _2817_ (.A(net230),
    .B(_0454_),
    .Y(_0456_));
 sg13g2_and2_1 _2818_ (.A(_0767_),
    .B(_0444_),
    .X(_0457_));
 sg13g2_nor3_1 _2819_ (.A(net672),
    .B(net231),
    .C(_0457_),
    .Y(_0043_));
 sg13g2_xnor2_1 _2820_ (.Y(_0458_),
    .A(net235),
    .B(_0457_));
 sg13g2_nor2_1 _2821_ (.A(net672),
    .B(_0458_),
    .Y(_0044_));
 sg13g2_a21oi_1 _2822_ (.A1(\pix_x[7] ),
    .A2(_0457_),
    .Y(_0459_),
    .B1(net216));
 sg13g2_and3_1 _2823_ (.X(_0460_),
    .A(net216),
    .B(\pix_x[7] ),
    .C(_0457_));
 sg13g2_nor3_1 _2824_ (.A(net672),
    .B(net217),
    .C(net236),
    .Y(_0045_));
 sg13g2_a21oi_1 _2825_ (.A1(net221),
    .A2(_0460_),
    .Y(_0461_),
    .B1(net672));
 sg13g2_o21ai_1 _2826_ (.B1(_0461_),
    .Y(_0462_),
    .A1(net221),
    .A2(_0460_));
 sg13g2_inv_1 _2827_ (.Y(_0046_),
    .A(_0462_));
 sg13g2_and2_1 _2828_ (.A(\gamepad.decoder.data_reg[5] ),
    .B(_0441_),
    .X(_0463_));
 sg13g2_or2_1 _2829_ (.X(_0464_),
    .B(\logo_left[8] ),
    .A(\logo_left[9] ));
 sg13g2_o21ai_1 _2830_ (.B1(_0463_),
    .Y(_0465_),
    .A1(_0838_),
    .A2(_0464_));
 sg13g2_and3_1 _2831_ (.X(_0466_),
    .A(\gamepad.decoder.data_reg[4] ),
    .B(_0850_),
    .C(_0441_));
 sg13g2_and2_2 _2832_ (.A(_0862_),
    .B(_0466_),
    .X(_0467_));
 sg13g2_nand2_1 _2833_ (.Y(_0468_),
    .A(_0862_),
    .B(_0466_));
 sg13g2_nor2_1 _2834_ (.A(net776),
    .B(_0467_),
    .Y(_0469_));
 sg13g2_a21oi_1 _2835_ (.A1(_0465_),
    .A2(_0469_),
    .Y(_0470_),
    .B1(_0786_));
 sg13g2_a21o_1 _2836_ (.A2(_0469_),
    .A1(_0465_),
    .B1(_0786_),
    .X(_0471_));
 sg13g2_o21ai_1 _2837_ (.B1(net806),
    .Y(_0472_),
    .A1(net802),
    .A2(net616));
 sg13g2_a21oi_1 _2838_ (.A1(_0737_),
    .A2(net616),
    .Y(_0047_),
    .B1(_0472_));
 sg13g2_nand2b_1 _2839_ (.Y(_0473_),
    .B(_0844_),
    .A_N(_0822_));
 sg13g2_xnor2_1 _2840_ (.Y(_0474_),
    .A(net621),
    .B(_0473_));
 sg13g2_nand2_1 _2841_ (.Y(_0475_),
    .A(net782),
    .B(_0474_));
 sg13g2_xor2_1 _2842_ (.B(net801),
    .A(net790),
    .X(_0476_));
 sg13g2_xnor2_1 _2843_ (.Y(_0477_),
    .A(_0737_),
    .B(_0476_));
 sg13g2_a21oi_1 _2844_ (.A1(net776),
    .A2(_0477_),
    .Y(_0478_),
    .B1(net615));
 sg13g2_o21ai_1 _2845_ (.B1(net806),
    .Y(_0479_),
    .A1(net801),
    .A2(net616));
 sg13g2_a21oi_1 _2846_ (.A1(_0475_),
    .A2(_0478_),
    .Y(_0048_),
    .B1(_0479_));
 sg13g2_xor2_1 _2847_ (.B(_0822_),
    .A(_0007_),
    .X(_0480_));
 sg13g2_xnor2_1 _2848_ (.Y(_0481_),
    .A(\logo_left[2] ),
    .B(_0844_));
 sg13g2_o21ai_1 _2849_ (.B1(net782),
    .Y(_0482_),
    .A1(net621),
    .A2(_0481_));
 sg13g2_a21oi_1 _2850_ (.A1(net621),
    .A2(_0480_),
    .Y(_0483_),
    .B1(_0482_));
 sg13g2_xnor2_1 _2851_ (.Y(_0484_),
    .A(net790),
    .B(\logo_left[2] ));
 sg13g2_a21oi_1 _2852_ (.A1(net790),
    .A2(_0844_),
    .Y(_0485_),
    .B1(_0822_));
 sg13g2_and2_1 _2853_ (.A(_0484_),
    .B(_0485_),
    .X(_0486_));
 sg13g2_o21ai_1 _2854_ (.B1(net776),
    .Y(_0487_),
    .A1(_0484_),
    .A2(_0485_));
 sg13g2_nor2_1 _2855_ (.A(_0486_),
    .B(_0487_),
    .Y(_0488_));
 sg13g2_nor3_1 _2856_ (.A(net615),
    .B(_0483_),
    .C(_0488_),
    .Y(_0489_));
 sg13g2_o21ai_1 _2857_ (.B1(net806),
    .Y(_0490_),
    .A1(net256),
    .A2(net616));
 sg13g2_nor2_1 _2858_ (.A(_0489_),
    .B(_0490_),
    .Y(_0049_));
 sg13g2_nor2_1 _2859_ (.A(net800),
    .B(net616),
    .Y(_0491_));
 sg13g2_nand2_1 _2860_ (.Y(_0492_),
    .A(_0856_),
    .B(_0467_));
 sg13g2_a21oi_1 _2861_ (.A1(_0828_),
    .A2(net621),
    .Y(_0493_),
    .B1(net776));
 sg13g2_nand2_1 _2862_ (.Y(_0494_),
    .A(net790),
    .B(_0735_));
 sg13g2_xnor2_1 _2863_ (.Y(_0495_),
    .A(net790),
    .B(net800));
 sg13g2_a21oi_1 _2864_ (.A1(_0726_),
    .A2(\logo_left[2] ),
    .Y(_0496_),
    .B1(_0486_));
 sg13g2_xnor2_1 _2865_ (.Y(_0497_),
    .A(_0495_),
    .B(_0496_));
 sg13g2_a221oi_1 _2866_ (.B2(net776),
    .C1(net615),
    .B1(_0497_),
    .A1(_0492_),
    .Y(_0498_),
    .A2(_0493_));
 sg13g2_o21ai_1 _2867_ (.B1(net806),
    .Y(_0050_),
    .A1(_0491_),
    .A2(_0498_));
 sg13g2_o21ai_1 _2868_ (.B1(net782),
    .Y(_0499_),
    .A1(_0826_),
    .A2(_0467_));
 sg13g2_a21oi_1 _2869_ (.A1(_0854_),
    .A2(_0467_),
    .Y(_0500_),
    .B1(_0499_));
 sg13g2_xor2_1 _2870_ (.B(net799),
    .A(net790),
    .X(_0501_));
 sg13g2_a22oi_1 _2871_ (.Y(_0502_),
    .B1(_0486_),
    .B2(_0494_),
    .A2(_0823_),
    .A1(_0726_));
 sg13g2_nor2_1 _2872_ (.A(_0501_),
    .B(_0502_),
    .Y(_0503_));
 sg13g2_a21oi_1 _2873_ (.A1(_0501_),
    .A2(_0502_),
    .Y(_0504_),
    .B1(net782));
 sg13g2_nor2b_1 _2874_ (.A(_0503_),
    .B_N(_0504_),
    .Y(_0505_));
 sg13g2_nor3_1 _2875_ (.A(net615),
    .B(_0500_),
    .C(_0505_),
    .Y(_0506_));
 sg13g2_o21ai_1 _2876_ (.B1(net806),
    .Y(_0507_),
    .A1(net799),
    .A2(net616));
 sg13g2_nor2_1 _2877_ (.A(_0506_),
    .B(_0507_),
    .Y(_0051_));
 sg13g2_nand2_1 _2878_ (.Y(_0508_),
    .A(_0836_),
    .B(_0468_));
 sg13g2_o21ai_1 _2879_ (.B1(_0508_),
    .Y(_0509_),
    .A1(_0853_),
    .A2(net621));
 sg13g2_xnor2_1 _2880_ (.Y(_0510_),
    .A(net789),
    .B(\logo_left[5] ));
 sg13g2_a21oi_1 _2881_ (.A1(_0726_),
    .A2(net799),
    .Y(_0511_),
    .B1(_0503_));
 sg13g2_xnor2_1 _2882_ (.Y(_0512_),
    .A(_0510_),
    .B(_0511_));
 sg13g2_nor2_1 _2883_ (.A(net782),
    .B(_0512_),
    .Y(_0513_));
 sg13g2_a21oi_1 _2884_ (.A1(net783),
    .A2(_0509_),
    .Y(_0514_),
    .B1(_0513_));
 sg13g2_o21ai_1 _2885_ (.B1(net806),
    .Y(_0515_),
    .A1(_0471_),
    .A2(_0514_));
 sg13g2_a21oi_1 _2886_ (.A1(_0734_),
    .A2(_0471_),
    .Y(_0052_),
    .B1(_0515_));
 sg13g2_o21ai_1 _2887_ (.B1(net783),
    .Y(_0516_),
    .A1(_0851_),
    .A2(net621));
 sg13g2_a21oi_1 _2888_ (.A1(_0835_),
    .A2(net621),
    .Y(_0517_),
    .B1(_0516_));
 sg13g2_xnor2_1 _2889_ (.Y(_0518_),
    .A(net789),
    .B(\logo_left[6] ));
 sg13g2_nand2_1 _2890_ (.Y(_0519_),
    .A(_0503_),
    .B(_0510_));
 sg13g2_nor2_1 _2891_ (.A(net789),
    .B(_0832_),
    .Y(_0520_));
 sg13g2_o21ai_1 _2892_ (.B1(_0519_),
    .Y(_0521_),
    .A1(net789),
    .A2(_0832_));
 sg13g2_nor2_1 _2893_ (.A(_0518_),
    .B(_0521_),
    .Y(_0522_));
 sg13g2_nand2_1 _2894_ (.Y(_0523_),
    .A(_0518_),
    .B(_0521_));
 sg13g2_nor2_1 _2895_ (.A(net782),
    .B(_0522_),
    .Y(_0524_));
 sg13g2_a21oi_1 _2896_ (.A1(_0523_),
    .A2(_0524_),
    .Y(_0525_),
    .B1(_0517_));
 sg13g2_o21ai_1 _2897_ (.B1(net806),
    .Y(_0526_),
    .A1(net615),
    .A2(_0525_));
 sg13g2_a21o_1 _2898_ (.A2(net615),
    .A1(net252),
    .B1(_0526_),
    .X(_0053_));
 sg13g2_a21oi_1 _2899_ (.A1(net798),
    .A2(_0471_),
    .Y(_0527_),
    .B1(net805));
 sg13g2_mux2_1 _2900_ (.A0(_0841_),
    .A1(_0860_),
    .S(_0467_),
    .X(_0528_));
 sg13g2_xnor2_1 _2901_ (.Y(_0529_),
    .A(net789),
    .B(net798));
 sg13g2_o21ai_1 _2902_ (.B1(_0523_),
    .Y(_0530_),
    .A1(net789),
    .A2(_0733_));
 sg13g2_xor2_1 _2903_ (.B(_0530_),
    .A(_0529_),
    .X(_0531_));
 sg13g2_a21oi_1 _2904_ (.A1(net782),
    .A2(_0528_),
    .Y(_0532_),
    .B1(net615));
 sg13g2_o21ai_1 _2905_ (.B1(_0532_),
    .Y(_0533_),
    .A1(net782),
    .A2(_0531_));
 sg13g2_nand2_1 _2906_ (.Y(_0054_),
    .A(_0527_),
    .B(_0533_));
 sg13g2_nand2_1 _2907_ (.Y(_0534_),
    .A(_0726_),
    .B(\logo_left[8] ));
 sg13g2_xor2_1 _2908_ (.B(\logo_left[8] ),
    .A(net789),
    .X(_0535_));
 sg13g2_nand2_1 _2909_ (.Y(_0536_),
    .A(_0518_),
    .B(_0529_));
 sg13g2_o21ai_1 _2910_ (.B1(_0726_),
    .Y(_0537_),
    .A1(net798),
    .A2(\logo_left[6] ));
 sg13g2_o21ai_1 _2911_ (.B1(_0537_),
    .Y(_0538_),
    .A1(_0519_),
    .A2(_0536_));
 sg13g2_nor2_1 _2912_ (.A(_0520_),
    .B(_0538_),
    .Y(_0539_));
 sg13g2_xor2_1 _2913_ (.B(_0539_),
    .A(_0535_),
    .X(_0540_));
 sg13g2_a22oi_1 _2914_ (.Y(_0541_),
    .B1(net621),
    .B2(_0840_),
    .A2(_0466_),
    .A1(_0861_));
 sg13g2_nand2_1 _2915_ (.Y(_0542_),
    .A(net783),
    .B(_0541_));
 sg13g2_o21ai_1 _2916_ (.B1(_0542_),
    .Y(_0543_),
    .A1(net783),
    .A2(_0540_));
 sg13g2_o21ai_1 _2917_ (.B1(net806),
    .Y(_0544_),
    .A1(net257),
    .A2(_0470_));
 sg13g2_a21oi_1 _2918_ (.A1(net616),
    .A2(_0543_),
    .Y(_0055_),
    .B1(_0544_));
 sg13g2_o21ai_1 _2919_ (.B1(_0534_),
    .Y(_0545_),
    .A1(_0535_),
    .A2(_0539_));
 sg13g2_xor2_1 _2920_ (.B(\logo_left[9] ),
    .A(net789),
    .X(_0546_));
 sg13g2_xnor2_1 _2921_ (.Y(_0547_),
    .A(_0545_),
    .B(_0546_));
 sg13g2_xor2_1 _2922_ (.B(_0839_),
    .A(\logo_left[9] ),
    .X(_0548_));
 sg13g2_a221oi_1 _2923_ (.B2(_0469_),
    .C1(net615),
    .B1(_0548_),
    .A1(net776),
    .Y(_0549_),
    .A2(_0547_));
 sg13g2_o21ai_1 _2924_ (.B1(net807),
    .Y(_0550_),
    .A1(net260),
    .A2(net616));
 sg13g2_nor2_1 _2925_ (.A(_0549_),
    .B(_0550_),
    .Y(_0056_));
 sg13g2_nand2b_1 _2926_ (.Y(_0551_),
    .B(_0811_),
    .A_N(_0813_));
 sg13g2_nand2b_1 _2927_ (.Y(_0552_),
    .B(_0551_),
    .A_N(_0798_));
 sg13g2_a21oi_1 _2928_ (.A1(_0810_),
    .A2(_0552_),
    .Y(_0553_),
    .B1(_0802_));
 sg13g2_and2_1 _2929_ (.A(net791),
    .B(\logo_top[8] ),
    .X(_0554_));
 sg13g2_nand2_1 _2930_ (.Y(_0555_),
    .A(\gamepad.decoder.data_reg[6] ),
    .B(_0441_));
 sg13g2_nor4_1 _2931_ (.A(_0819_),
    .B(_0553_),
    .C(_0554_),
    .D(_0555_),
    .Y(_0556_));
 sg13g2_and2_1 _2932_ (.A(\gamepad.decoder.data_reg[7] ),
    .B(_0441_),
    .X(_0557_));
 sg13g2_nand2_1 _2933_ (.Y(_0558_),
    .A(\gamepad.decoder.data_reg[7] ),
    .B(_0441_));
 sg13g2_nor2_1 _2934_ (.A(\logo_top[3] ),
    .B(net795),
    .Y(_0559_));
 sg13g2_and2_1 _2935_ (.A(_0803_),
    .B(_0559_),
    .X(_0560_));
 sg13g2_nor2_1 _2936_ (.A(net793),
    .B(net794),
    .Y(_0561_));
 sg13g2_nand2_1 _2937_ (.Y(_0562_),
    .A(_0560_),
    .B(_0561_));
 sg13g2_nor3_2 _2938_ (.A(net792),
    .B(\logo_top[6] ),
    .C(_0562_),
    .Y(_0563_));
 sg13g2_nor2_1 _2939_ (.A(net791),
    .B(\logo_top[8] ),
    .Y(_0564_));
 sg13g2_a21oi_1 _2940_ (.A1(_0563_),
    .A2(_0564_),
    .Y(_0565_),
    .B1(_0558_));
 sg13g2_nand2b_1 _2941_ (.Y(_0566_),
    .B(net785),
    .A_N(_0565_));
 sg13g2_nor2_1 _2942_ (.A(net618),
    .B(_0566_),
    .Y(_0567_));
 sg13g2_nor2_2 _2943_ (.A(_0786_),
    .B(_0567_),
    .Y(_0568_));
 sg13g2_o21ai_1 _2944_ (.B1(_0787_),
    .Y(_0569_),
    .A1(net618),
    .A2(_0566_));
 sg13g2_o21ai_1 _2945_ (.B1(net809),
    .Y(_0570_),
    .A1(net195),
    .A2(net613));
 sg13g2_a21oi_1 _2946_ (.A1(_0732_),
    .A2(net613),
    .Y(_0057_),
    .B1(_0570_));
 sg13g2_o21ai_1 _2947_ (.B1(net617),
    .Y(_0571_),
    .A1(_0790_),
    .A2(_0803_));
 sg13g2_nor3_1 _2948_ (.A(_0790_),
    .B(_0803_),
    .C(net617),
    .Y(_0572_));
 sg13g2_nor2_1 _2949_ (.A(net775),
    .B(_0572_),
    .Y(_0573_));
 sg13g2_xnor2_1 _2950_ (.Y(_0574_),
    .A(net786),
    .B(net796));
 sg13g2_xnor2_1 _2951_ (.Y(_0575_),
    .A(net195),
    .B(_0574_));
 sg13g2_a221oi_1 _2952_ (.B2(net775),
    .C1(net613),
    .B1(_0575_),
    .A1(_0571_),
    .Y(_0576_),
    .A2(_0573_));
 sg13g2_o21ai_1 _2953_ (.B1(net809),
    .Y(_0577_),
    .A1(net796),
    .A2(_0568_));
 sg13g2_nor2_1 _2954_ (.A(_0576_),
    .B(_0577_),
    .Y(_0058_));
 sg13g2_xnor2_1 _2955_ (.Y(_0578_),
    .A(net795),
    .B(_0790_));
 sg13g2_xnor2_1 _2956_ (.Y(_0579_),
    .A(_0011_),
    .B(_0803_));
 sg13g2_o21ai_1 _2957_ (.B1(net784),
    .Y(_0580_),
    .A1(net617),
    .A2(_0579_));
 sg13g2_a21oi_1 _2958_ (.A1(net617),
    .A2(_0578_),
    .Y(_0581_),
    .B1(_0580_));
 sg13g2_xnor2_1 _2959_ (.Y(_0582_),
    .A(net786),
    .B(net795));
 sg13g2_a21oi_1 _2960_ (.A1(net786),
    .A2(_0791_),
    .Y(_0583_),
    .B1(_0803_));
 sg13g2_and2_1 _2961_ (.A(_0582_),
    .B(_0583_),
    .X(_0584_));
 sg13g2_o21ai_1 _2962_ (.B1(net775),
    .Y(_0585_),
    .A1(_0582_),
    .A2(_0583_));
 sg13g2_nor2_1 _2963_ (.A(_0584_),
    .B(_0585_),
    .Y(_0586_));
 sg13g2_nor3_1 _2964_ (.A(net613),
    .B(_0581_),
    .C(_0586_),
    .Y(_0587_));
 sg13g2_o21ai_1 _2965_ (.B1(net809),
    .Y(_0588_),
    .A1(net795),
    .A2(_0568_));
 sg13g2_nor2_1 _2966_ (.A(_0587_),
    .B(_0588_),
    .Y(_0059_));
 sg13g2_o21ai_1 _2967_ (.B1(net784),
    .Y(_0589_),
    .A1(_0805_),
    .A2(net617));
 sg13g2_a21oi_1 _2968_ (.A1(_0817_),
    .A2(net617),
    .Y(_0590_),
    .B1(_0589_));
 sg13g2_xor2_1 _2969_ (.B(\logo_top[3] ),
    .A(net786),
    .X(_0591_));
 sg13g2_a21oi_1 _2970_ (.A1(_0725_),
    .A2(net795),
    .Y(_0592_),
    .B1(_0584_));
 sg13g2_xnor2_1 _2971_ (.Y(_0593_),
    .A(_0591_),
    .B(_0592_));
 sg13g2_nor2_1 _2972_ (.A(net784),
    .B(_0593_),
    .Y(_0594_));
 sg13g2_o21ai_1 _2973_ (.B1(_0568_),
    .Y(_0595_),
    .A1(_0590_),
    .A2(_0594_));
 sg13g2_a21oi_1 _2974_ (.A1(net250),
    .A2(net613),
    .Y(_0596_),
    .B1(net804));
 sg13g2_nand2_1 _2975_ (.Y(_0060_),
    .A(_0595_),
    .B(_0596_));
 sg13g2_nand2_1 _2976_ (.Y(_0597_),
    .A(_0012_),
    .B(_0560_));
 sg13g2_xnor2_1 _2977_ (.Y(_0598_),
    .A(_0012_),
    .B(_0560_));
 sg13g2_mux2_1 _2978_ (.A0(_0598_),
    .A1(_0814_),
    .S(net617),
    .X(_0599_));
 sg13g2_nand2_1 _2979_ (.Y(_0600_),
    .A(net785),
    .B(_0599_));
 sg13g2_nor2b_1 _2980_ (.A(net787),
    .B_N(net794),
    .Y(_0601_));
 sg13g2_xnor2_1 _2981_ (.Y(_0602_),
    .A(net787),
    .B(net794));
 sg13g2_o21ai_1 _2982_ (.B1(_0584_),
    .Y(_0603_),
    .A1(_0725_),
    .A2(\logo_top[3] ));
 sg13g2_o21ai_1 _2983_ (.B1(_0603_),
    .Y(_0604_),
    .A1(net786),
    .A2(_0559_));
 sg13g2_xor2_1 _2984_ (.B(_0604_),
    .A(_0602_),
    .X(_0605_));
 sg13g2_a21oi_1 _2985_ (.A1(net775),
    .A2(_0605_),
    .Y(_0606_),
    .B1(net613));
 sg13g2_o21ai_1 _2986_ (.B1(net809),
    .Y(_0607_),
    .A1(net794),
    .A2(_0568_));
 sg13g2_a21oi_1 _2987_ (.A1(_0600_),
    .A2(_0606_),
    .Y(_0061_),
    .B1(_0607_));
 sg13g2_xnor2_1 _2988_ (.Y(_0608_),
    .A(net793),
    .B(_0597_));
 sg13g2_nand2b_1 _2989_ (.Y(_0609_),
    .B(_0608_),
    .A_N(net617));
 sg13g2_a21oi_1 _2990_ (.A1(_0813_),
    .A2(net618),
    .Y(_0610_),
    .B1(net775));
 sg13g2_a21o_1 _2991_ (.A2(_0604_),
    .A1(_0602_),
    .B1(_0601_),
    .X(_0611_));
 sg13g2_xnor2_1 _2992_ (.Y(_0612_),
    .A(net787),
    .B(net793));
 sg13g2_xnor2_1 _2993_ (.Y(_0613_),
    .A(_0611_),
    .B(_0612_));
 sg13g2_a22oi_1 _2994_ (.Y(_0614_),
    .B1(_0613_),
    .B2(net775),
    .A2(_0610_),
    .A1(_0609_));
 sg13g2_o21ai_1 _2995_ (.B1(net809),
    .Y(_0615_),
    .A1(net613),
    .A2(_0614_));
 sg13g2_a21oi_1 _2996_ (.A1(_0729_),
    .A2(net613),
    .Y(_0062_),
    .B1(_0615_));
 sg13g2_nand3_1 _2997_ (.B(_0560_),
    .C(_0561_),
    .A(_0013_),
    .Y(_0616_));
 sg13g2_xor2_1 _2998_ (.B(_0562_),
    .A(_0013_),
    .X(_0617_));
 sg13g2_mux2_1 _2999_ (.A0(_0617_),
    .A1(_0796_),
    .S(net618),
    .X(_0618_));
 sg13g2_xor2_1 _3000_ (.B(\logo_top[6] ),
    .A(net788),
    .X(_0619_));
 sg13g2_nand3_1 _3001_ (.B(_0604_),
    .C(_0612_),
    .A(_0602_),
    .Y(_0620_));
 sg13g2_or2_1 _3002_ (.X(_0621_),
    .B(_0561_),
    .A(net788));
 sg13g2_and3_1 _3003_ (.X(_0622_),
    .A(_0619_),
    .B(_0620_),
    .C(_0621_));
 sg13g2_a21oi_1 _3004_ (.A1(_0620_),
    .A2(_0621_),
    .Y(_0623_),
    .B1(_0619_));
 sg13g2_nor3_1 _3005_ (.A(net784),
    .B(_0622_),
    .C(_0623_),
    .Y(_0624_));
 sg13g2_a21oi_1 _3006_ (.A1(net784),
    .A2(_0618_),
    .Y(_0625_),
    .B1(_0624_));
 sg13g2_a21oi_1 _3007_ (.A1(net255),
    .A2(net614),
    .Y(_0626_),
    .B1(net804));
 sg13g2_o21ai_1 _3008_ (.B1(_0626_),
    .Y(_0063_),
    .A1(net614),
    .A2(_0625_));
 sg13g2_xnor2_1 _3009_ (.Y(_0627_),
    .A(_0728_),
    .B(_0616_));
 sg13g2_nand2b_1 _3010_ (.Y(_0628_),
    .B(_0627_),
    .A_N(net618));
 sg13g2_a21oi_1 _3011_ (.A1(_0797_),
    .A2(net618),
    .Y(_0629_),
    .B1(net775));
 sg13g2_xor2_1 _3012_ (.B(\logo_top[7] ),
    .A(net788),
    .X(_0630_));
 sg13g2_a21o_1 _3013_ (.A2(\logo_top[6] ),
    .A1(_0725_),
    .B1(_0623_),
    .X(_0631_));
 sg13g2_xnor2_1 _3014_ (.Y(_0632_),
    .A(_0630_),
    .B(_0631_));
 sg13g2_a221oi_1 _3015_ (.B2(net775),
    .C1(net614),
    .B1(_0632_),
    .A1(_0628_),
    .Y(_0633_),
    .A2(_0629_));
 sg13g2_nor2_1 _3016_ (.A(net792),
    .B(_0568_),
    .Y(_0634_));
 sg13g2_o21ai_1 _3017_ (.B1(net808),
    .Y(_0064_),
    .A1(_0633_),
    .A2(_0634_));
 sg13g2_nand2_1 _3018_ (.Y(_0635_),
    .A(_0014_),
    .B(_0563_));
 sg13g2_xnor2_1 _3019_ (.Y(_0636_),
    .A(_0014_),
    .B(_0563_));
 sg13g2_mux2_1 _3020_ (.A0(_0636_),
    .A1(_0809_),
    .S(net618),
    .X(_0637_));
 sg13g2_nand2_1 _3021_ (.Y(_0638_),
    .A(net785),
    .B(_0637_));
 sg13g2_xnor2_1 _3022_ (.Y(_0639_),
    .A(net788),
    .B(\logo_top[8] ));
 sg13g2_nor3_1 _3023_ (.A(_0619_),
    .B(_0620_),
    .C(_0630_),
    .Y(_0640_));
 sg13g2_o21ai_1 _3024_ (.B1(_0725_),
    .Y(_0641_),
    .A1(net792),
    .A2(\logo_top[6] ));
 sg13g2_nand2_1 _3025_ (.Y(_0642_),
    .A(_0621_),
    .B(_0641_));
 sg13g2_o21ai_1 _3026_ (.B1(_0639_),
    .Y(_0643_),
    .A1(_0640_),
    .A2(_0642_));
 sg13g2_nor3_1 _3027_ (.A(_0639_),
    .B(_0640_),
    .C(_0642_),
    .Y(_0644_));
 sg13g2_nor2_1 _3028_ (.A(net784),
    .B(_0644_),
    .Y(_0645_));
 sg13g2_a21oi_1 _3029_ (.A1(_0643_),
    .A2(_0645_),
    .Y(_0646_),
    .B1(net614));
 sg13g2_a221oi_1 _3030_ (.B2(_0646_),
    .C1(net804),
    .B1(_0638_),
    .A1(_0727_),
    .Y(_0065_),
    .A2(net614));
 sg13g2_o21ai_1 _3031_ (.B1(_0643_),
    .Y(_0647_),
    .A1(net788),
    .A2(_0727_));
 sg13g2_xnor2_1 _3032_ (.Y(_0648_),
    .A(net788),
    .B(\logo_top[9] ));
 sg13g2_xnor2_1 _3033_ (.Y(_0649_),
    .A(_0647_),
    .B(_0648_));
 sg13g2_nor2_1 _3034_ (.A(net784),
    .B(_0649_),
    .Y(_0650_));
 sg13g2_xor2_1 _3035_ (.B(_0635_),
    .A(net791),
    .X(_0651_));
 sg13g2_nor3_1 _3036_ (.A(_0724_),
    .B(net618),
    .C(_0651_),
    .Y(_0652_));
 sg13g2_nor3_1 _3037_ (.A(net614),
    .B(_0650_),
    .C(_0652_),
    .Y(_0653_));
 sg13g2_o21ai_1 _3038_ (.B1(net808),
    .Y(_0654_),
    .A1(net791),
    .A2(_0568_));
 sg13g2_nor2_1 _3039_ (.A(_0653_),
    .B(_0654_),
    .Y(_0066_));
 sg13g2_o21ai_1 _3040_ (.B1(_0441_),
    .Y(_0655_),
    .A1(\gamepad.decoder.data_reg[5] ),
    .A2(\gamepad.decoder.data_reg[4] ));
 sg13g2_nand2_1 _3041_ (.Y(_0656_),
    .A(_0866_),
    .B(_0655_));
 sg13g2_a21o_1 _3042_ (.A2(_0656_),
    .A1(_0788_),
    .B1(_0726_),
    .X(_0657_));
 sg13g2_nand2b_1 _3043_ (.Y(_0658_),
    .B(_0463_),
    .A_N(_0843_));
 sg13g2_nand4_1 _3044_ (.B(_0865_),
    .C(_0656_),
    .A(_0788_),
    .Y(_0659_),
    .D(_0658_));
 sg13g2_nand3_1 _3045_ (.B(_0657_),
    .C(_0659_),
    .A(net807),
    .Y(_0067_));
 sg13g2_nand3_1 _3046_ (.B(_0555_),
    .C(_0558_),
    .A(_0821_),
    .Y(_0660_));
 sg13g2_nand2_1 _3047_ (.Y(_0661_),
    .A(_0788_),
    .B(_0660_));
 sg13g2_a22oi_1 _3048_ (.Y(_0662_),
    .B1(_0557_),
    .B2(_0808_),
    .A2(_0819_),
    .A1(net786));
 sg13g2_mux2_1 _3049_ (.A0(_0662_),
    .A1(net786),
    .S(_0661_),
    .X(_0663_));
 sg13g2_and2_1 _3050_ (.A(net809),
    .B(_0663_),
    .X(_0068_));
 sg13g2_or2_1 _3051_ (.X(_0664_),
    .B(_0442_),
    .A(gamepad_start_prev));
 sg13g2_o21ai_1 _3052_ (.B1(net807),
    .Y(_0665_),
    .A1(net133),
    .A2(_0664_));
 sg13g2_a21oi_1 _3053_ (.A1(net776),
    .A2(_0664_),
    .Y(_0069_),
    .B1(net134));
 sg13g2_nand2b_1 _3054_ (.Y(_0666_),
    .B(\color_index[0] ),
    .A_N(net612));
 sg13g2_nand2_1 _3055_ (.Y(_0667_),
    .A(net136),
    .B(net612));
 sg13g2_a21oi_1 _3056_ (.A1(_0666_),
    .A2(_0667_),
    .Y(_0070_),
    .B1(net804));
 sg13g2_nand2b_1 _3057_ (.Y(_0668_),
    .B(net213),
    .A_N(net612));
 sg13g2_o21ai_1 _3058_ (.B1(net810),
    .Y(_0669_),
    .A1(net213),
    .A2(\color_index[0] ));
 sg13g2_a21oi_1 _3059_ (.A1(_0876_),
    .A2(_0668_),
    .Y(_0071_),
    .B1(_0669_));
 sg13g2_nand2b_1 _3060_ (.Y(_0670_),
    .B(net138),
    .A_N(net612));
 sg13g2_a21oi_1 _3061_ (.A1(_0872_),
    .A2(_0670_),
    .Y(_0072_),
    .B1(net804));
 sg13g2_nor2_1 _3062_ (.A(net808),
    .B(net171),
    .Y(_0671_));
 sg13g2_a21oi_1 _3063_ (.A1(_0739_),
    .A2(net808),
    .Y(_0073_),
    .B1(_0671_));
 sg13g2_mux2_1 _3064_ (.A0(net186),
    .A1(net781),
    .S(net808),
    .X(_0074_));
 sg13g2_mux2_1 _3065_ (.A0(net177),
    .A1(net780),
    .S(net811),
    .X(_0075_));
 sg13g2_mux2_1 _3066_ (.A0(net173),
    .A1(net779),
    .S(net811),
    .X(_0076_));
 sg13g2_nor2_1 _3067_ (.A(net811),
    .B(net160),
    .Y(_0672_));
 sg13g2_a21oi_1 _3068_ (.A1(_0740_),
    .A2(net811),
    .Y(_0077_),
    .B1(_0672_));
 sg13g2_nor2_1 _3069_ (.A(net811),
    .B(net167),
    .Y(_0673_));
 sg13g2_a21oi_1 _3070_ (.A1(_0741_),
    .A2(net811),
    .Y(_0078_),
    .B1(_0673_));
 sg13g2_nor2_1 _3071_ (.A(net809),
    .B(net175),
    .Y(_0674_));
 sg13g2_a21oi_1 _3072_ (.A1(_0742_),
    .A2(net813),
    .Y(_0079_),
    .B1(_0674_));
 sg13g2_mux2_1 _3073_ (.A0(net179),
    .A1(net777),
    .S(net811),
    .X(_0080_));
 sg13g2_nor2_1 _3074_ (.A(net808),
    .B(net158),
    .Y(_0675_));
 sg13g2_a21oi_1 _3075_ (.A1(net808),
    .A2(_0744_),
    .Y(_0081_),
    .B1(_0675_));
 sg13g2_a21oi_1 _3076_ (.A1(net804),
    .A2(_0748_),
    .Y(_0082_),
    .B1(_0400_));
 sg13g2_xnor2_1 _3077_ (.Y(_0676_),
    .A(net733),
    .B(_0417_));
 sg13g2_nand2_1 _3078_ (.Y(_0677_),
    .A(net229),
    .B(net2));
 sg13g2_o21ai_1 _3079_ (.B1(_0677_),
    .Y(_0678_),
    .A1(net2),
    .A2(_0676_));
 sg13g2_and2_1 _3080_ (.A(_0403_),
    .B(_0678_),
    .X(_0083_));
 sg13g2_xnor2_1 _3081_ (.Y(_0679_),
    .A(_0418_),
    .B(_0419_));
 sg13g2_mux2_1 _3082_ (.A0(net240),
    .A1(_0679_),
    .S(_0762_),
    .X(_0680_));
 sg13g2_and2_1 _3083_ (.A(_0403_),
    .B(_0680_),
    .X(_0084_));
 sg13g2_xnor2_1 _3084_ (.Y(_0681_),
    .A(_0421_),
    .B(_0422_));
 sg13g2_mux2_1 _3085_ (.A0(net228),
    .A1(_0681_),
    .S(_0762_),
    .X(_0682_));
 sg13g2_and2_1 _3086_ (.A(_0403_),
    .B(_0682_),
    .X(_0085_));
 sg13g2_nand2b_1 _3087_ (.Y(_0683_),
    .B(net2),
    .A_N(net215));
 sg13g2_and3_1 _3088_ (.X(_0684_),
    .A(_0414_),
    .B(_0423_),
    .C(_0424_));
 sg13g2_o21ai_1 _3089_ (.B1(_0762_),
    .Y(_0685_),
    .A1(_0425_),
    .A2(_0684_));
 sg13g2_and3_1 _3090_ (.X(_0086_),
    .A(_0403_),
    .B(_0683_),
    .C(_0685_));
 sg13g2_nor2b_1 _3091_ (.A(\gamepad.driver.pmod_clk_prev ),
    .B_N(\gamepad.driver.pmod_clk_sync[1] ),
    .Y(_0686_));
 sg13g2_nor2_1 _3092_ (.A(net804),
    .B(net759),
    .Y(_0687_));
 sg13g2_a22oi_1 _3093_ (.Y(_0087_),
    .B1(net744),
    .B2(_0722_),
    .A2(net760),
    .A1(_0723_));
 sg13g2_a22oi_1 _3094_ (.Y(_0088_),
    .B1(net745),
    .B2(_0721_),
    .A2(net760),
    .A1(_0722_));
 sg13g2_a22oi_1 _3095_ (.Y(_0089_),
    .B1(net745),
    .B2(_0720_),
    .A2(net760),
    .A1(_0721_));
 sg13g2_a22oi_1 _3096_ (.Y(_0090_),
    .B1(net745),
    .B2(_0719_),
    .A2(net760),
    .A1(_0720_));
 sg13g2_a22oi_1 _3097_ (.Y(_0091_),
    .B1(net744),
    .B2(_0718_),
    .A2(net759),
    .A1(_0719_));
 sg13g2_a22oi_1 _3098_ (.Y(_0092_),
    .B1(net744),
    .B2(_0717_),
    .A2(net759),
    .A1(_0718_));
 sg13g2_a22oi_1 _3099_ (.Y(_0093_),
    .B1(net744),
    .B2(_0716_),
    .A2(net759),
    .A1(_0717_));
 sg13g2_a22oi_1 _3100_ (.Y(_0094_),
    .B1(net744),
    .B2(_0715_),
    .A2(net759),
    .A1(_0716_));
 sg13g2_a22oi_1 _3101_ (.Y(_0095_),
    .B1(net744),
    .B2(_0714_),
    .A2(net759),
    .A1(_0715_));
 sg13g2_a22oi_1 _3102_ (.Y(_0096_),
    .B1(net744),
    .B2(_0713_),
    .A2(net759),
    .A1(_0714_));
 sg13g2_a22oi_1 _3103_ (.Y(_0097_),
    .B1(net744),
    .B2(_0712_),
    .A2(net759),
    .A1(_0713_));
 sg13g2_a22oi_1 _3104_ (.Y(_0098_),
    .B1(net745),
    .B2(_0738_),
    .A2(net760),
    .A1(_0712_));
 sg13g2_and2_1 _3105_ (.A(net810),
    .B(net5),
    .X(_0099_));
 sg13g2_and2_1 _3106_ (.A(net812),
    .B(net131),
    .X(_0100_));
 sg13g2_and2_1 _3107_ (.A(net812),
    .B(net4),
    .X(_0101_));
 sg13g2_and2_1 _3108_ (.A(net812),
    .B(net130),
    .X(_0102_));
 sg13g2_and2_1 _3109_ (.A(net810),
    .B(net3),
    .X(_0103_));
 sg13g2_and2_1 _3110_ (.A(net810),
    .B(net157),
    .X(_0104_));
 sg13g2_and2_1 _3111_ (.A(net780),
    .B(net779),
    .X(_0688_));
 sg13g2_nand4_1 _3112_ (.B(\pix_y[9] ),
    .C(_0784_),
    .A(_0744_),
    .Y(_0689_),
    .D(_0688_));
 sg13g2_and2_2 _3113_ (.A(net808),
    .B(_0689_),
    .X(_0690_));
 sg13g2_nand3_1 _3114_ (.B(_0447_),
    .C(_0690_),
    .A(net128),
    .Y(_0691_));
 sg13g2_o21ai_1 _3115_ (.B1(_0691_),
    .Y(_0105_),
    .A1(_0739_),
    .A2(_0449_));
 sg13g2_a21oi_1 _3116_ (.A1(\pix_y[0] ),
    .A2(net672),
    .Y(_0692_),
    .B1(net146));
 sg13g2_and2_1 _3117_ (.A(\pix_y[0] ),
    .B(net781),
    .X(_0693_));
 sg13g2_and2_1 _3118_ (.A(net672),
    .B(_0693_),
    .X(_0694_));
 sg13g2_nor2_2 _3119_ (.A(_0448_),
    .B(_0690_),
    .Y(_0695_));
 sg13g2_nor3_1 _3120_ (.A(net147),
    .B(_0694_),
    .C(_0695_),
    .Y(_0106_));
 sg13g2_a21o_1 _3121_ (.A2(_0694_),
    .A1(net237),
    .B1(_0695_),
    .X(_0696_));
 sg13g2_nor2_1 _3122_ (.A(net780),
    .B(_0694_),
    .Y(_0697_));
 sg13g2_nor2_1 _3123_ (.A(_0696_),
    .B(_0697_),
    .Y(_0107_));
 sg13g2_and4_1 _3124_ (.A(net780),
    .B(_0447_),
    .C(_0690_),
    .D(_0693_),
    .X(_0698_));
 sg13g2_nor2_1 _3125_ (.A(net181),
    .B(_0698_),
    .Y(_0699_));
 sg13g2_a21oi_1 _3126_ (.A1(net779),
    .A2(_0696_),
    .Y(_0108_),
    .B1(_0699_));
 sg13g2_and3_2 _3127_ (.X(_0700_),
    .A(net156),
    .B(_0688_),
    .C(_0694_));
 sg13g2_nor2_1 _3128_ (.A(_0695_),
    .B(_0700_),
    .Y(_0701_));
 sg13g2_a21oi_1 _3129_ (.A1(_0688_),
    .A2(_0694_),
    .Y(_0702_),
    .B1(net156));
 sg13g2_nor3_1 _3130_ (.A(_0695_),
    .B(_0700_),
    .C(_0702_),
    .Y(_0109_));
 sg13g2_nand2_1 _3131_ (.Y(_0703_),
    .A(net238),
    .B(_0701_));
 sg13g2_nand2_1 _3132_ (.Y(_0704_),
    .A(_0690_),
    .B(_0700_));
 sg13g2_o21ai_1 _3133_ (.B1(_0703_),
    .Y(_0110_),
    .A1(net238),
    .A2(_0704_));
 sg13g2_a21oi_1 _3134_ (.A1(_0763_),
    .A2(_0700_),
    .Y(_0705_),
    .B1(_0695_));
 sg13g2_a21o_1 _3135_ (.A2(_0700_),
    .A1(net238),
    .B1(net247),
    .X(_0706_));
 sg13g2_and2_1 _3136_ (.A(_0705_),
    .B(_0706_),
    .X(_0111_));
 sg13g2_nand2_1 _3137_ (.Y(_0707_),
    .A(net777),
    .B(_0705_));
 sg13g2_nand4_1 _3138_ (.B(net778),
    .C(_0763_),
    .A(net181),
    .Y(_0708_),
    .D(_0698_));
 sg13g2_o21ai_1 _3139_ (.B1(_0707_),
    .Y(_0112_),
    .A1(net777),
    .A2(_0708_));
 sg13g2_a21oi_1 _3140_ (.A1(_0764_),
    .A2(_0690_),
    .Y(_0709_),
    .B1(_0701_));
 sg13g2_nand3_1 _3141_ (.B(_0763_),
    .C(_0700_),
    .A(net777),
    .Y(_0710_));
 sg13g2_a21oi_1 _3142_ (.A1(_0744_),
    .A2(_0710_),
    .Y(_0113_),
    .B1(_0709_));
 sg13g2_nand2b_1 _3143_ (.Y(_0711_),
    .B(net239),
    .A_N(_0709_));
 sg13g2_o21ai_1 _3144_ (.B1(_0711_),
    .Y(_0114_),
    .A1(_0765_),
    .A2(_0704_));
 sg13g2_a21o_1 _3145_ (.A2(_0877_),
    .A1(net810),
    .B1(_0115_),
    .X(_0116_));
 sg13g2_dfrbp_1 _3146_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net87),
    .D(_0022_),
    .Q_N(_1564_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _3147_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net40),
    .D(_0023_),
    .Q_N(_1563_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _3148_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net39),
    .D(net149),
    .Q_N(_1562_),
    .Q(\gamepad.decoder.data_reg[0] ));
 sg13g2_dfrbp_1 _3149_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net37),
    .D(net153),
    .Q_N(_1561_),
    .Q(\gamepad.decoder.data_reg[1] ));
 sg13g2_dfrbp_1 _3150_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net35),
    .D(net145),
    .Q_N(_1560_),
    .Q(\gamepad.decoder.data_reg[2] ));
 sg13g2_dfrbp_1 _3151_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net33),
    .D(net151),
    .Q_N(_1559_),
    .Q(\gamepad.decoder.data_reg[3] ));
 sg13g2_dfrbp_1 _3152_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net31),
    .D(net209),
    .Q_N(_1558_),
    .Q(\gamepad.decoder.data_reg[4] ));
 sg13g2_dfrbp_1 _3153_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net29),
    .D(net207),
    .Q_N(_1557_),
    .Q(\gamepad.decoder.data_reg[5] ));
 sg13g2_dfrbp_1 _3154_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net27),
    .D(net164),
    .Q_N(_1556_),
    .Q(\gamepad.decoder.data_reg[6] ));
 sg13g2_dfrbp_1 _3155_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net25),
    .D(_0031_),
    .Q_N(_1555_),
    .Q(\gamepad.decoder.data_reg[7] ));
 sg13g2_dfrbp_1 _3156_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net23),
    .D(net166),
    .Q_N(_1554_),
    .Q(\gamepad.decoder.data_reg[8] ));
 sg13g2_dfrbp_1 _3157_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net124),
    .D(net155),
    .Q_N(_1553_),
    .Q(\gamepad.decoder.data_reg[9] ));
 sg13g2_dfrbp_1 _3158_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net117),
    .D(net143),
    .Q_N(_1552_),
    .Q(\gamepad.decoder.data_reg[10] ));
 sg13g2_dfrbp_1 _3159_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net115),
    .D(net170),
    .Q_N(_1551_),
    .Q(\gamepad.decoder.data_reg[11] ));
 sg13g2_dfrbp_1 _3160_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net113),
    .D(net141),
    .Q_N(_1550_),
    .Q(gamepad_start_prev));
 sg13g2_dfrbp_1 _3161_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net111),
    .D(_0037_),
    .Q_N(_0021_),
    .Q(\pix_x[0] ));
 sg13g2_dfrbp_1 _3162_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net110),
    .D(_0038_),
    .Q_N(_1549_),
    .Q(\pix_x[1] ));
 sg13g2_dfrbp_1 _3163_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net109),
    .D(net220),
    .Q_N(_1548_),
    .Q(\pix_x[2] ));
 sg13g2_dfrbp_1 _3164_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net108),
    .D(_0040_),
    .Q_N(_1547_),
    .Q(\pix_x[3] ));
 sg13g2_dfrbp_1 _3165_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net106),
    .D(_0041_),
    .Q_N(_1546_),
    .Q(\pix_x[4] ));
 sg13g2_dfrbp_1 _3166_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net105),
    .D(_0042_),
    .Q_N(_1545_),
    .Q(\pix_x[5] ));
 sg13g2_dfrbp_1 _3167_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net104),
    .D(_0043_),
    .Q_N(_1544_),
    .Q(\pix_x[6] ));
 sg13g2_dfrbp_1 _3168_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net103),
    .D(_0044_),
    .Q_N(_1543_),
    .Q(\pix_x[7] ));
 sg13g2_dfrbp_1 _3169_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net102),
    .D(_0045_),
    .Q_N(_1542_),
    .Q(\pix_x[8] ));
 sg13g2_dfrbp_1 _3170_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net101),
    .D(_0046_),
    .Q_N(_1541_),
    .Q(\pix_x[9] ));
 sg13g2_dfrbp_1 _3171_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net100),
    .D(_0047_),
    .Q_N(_0020_),
    .Q(\logo_left[0] ));
 sg13g2_dfrbp_1 _3172_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net98),
    .D(_0048_),
    .Q_N(_1540_),
    .Q(\logo_left[1] ));
 sg13g2_dfrbp_1 _3173_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net96),
    .D(_0049_),
    .Q_N(_0007_),
    .Q(\logo_left[2] ));
 sg13g2_dfrbp_1 _3174_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net94),
    .D(_0050_),
    .Q_N(_1539_),
    .Q(\logo_left[3] ));
 sg13g2_dfrbp_1 _3175_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net92),
    .D(_0051_),
    .Q_N(_0008_),
    .Q(\logo_left[4] ));
 sg13g2_dfrbp_1 _3176_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net90),
    .D(_0052_),
    .Q_N(_1538_),
    .Q(\logo_left[5] ));
 sg13g2_dfrbp_1 _3177_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net86),
    .D(_0053_),
    .Q_N(_0009_),
    .Q(\logo_left[6] ));
 sg13g2_dfrbp_1 _3178_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net84),
    .D(_0054_),
    .Q_N(_1537_),
    .Q(\logo_left[7] ));
 sg13g2_dfrbp_1 _3179_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net82),
    .D(_0055_),
    .Q_N(_0010_),
    .Q(\logo_left[8] ));
 sg13g2_dfrbp_1 _3180_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net80),
    .D(_0056_),
    .Q_N(_1536_),
    .Q(\logo_left[9] ));
 sg13g2_dfrbp_1 _3181_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net78),
    .D(net196),
    .Q_N(_0019_),
    .Q(\logo_top[0] ));
 sg13g2_dfrbp_1 _3182_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net76),
    .D(_0058_),
    .Q_N(_1535_),
    .Q(\logo_top[1] ));
 sg13g2_dfrbp_1 _3183_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net74),
    .D(_0059_),
    .Q_N(_0011_),
    .Q(\logo_top[2] ));
 sg13g2_dfrbp_1 _3184_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net72),
    .D(_0060_),
    .Q_N(_1534_),
    .Q(\logo_top[3] ));
 sg13g2_dfrbp_1 _3185_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net70),
    .D(net243),
    .Q_N(_0012_),
    .Q(\logo_top[4] ));
 sg13g2_dfrbp_1 _3186_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net68),
    .D(_0062_),
    .Q_N(_1533_),
    .Q(\logo_top[5] ));
 sg13g2_dfrbp_1 _3187_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net66),
    .D(_0063_),
    .Q_N(_0013_),
    .Q(\logo_top[6] ));
 sg13g2_dfrbp_1 _3188_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net64),
    .D(_0064_),
    .Q_N(_1532_),
    .Q(\logo_top[7] ));
 sg13g2_dfrbp_1 _3189_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net62),
    .D(_0065_),
    .Q_N(_0014_),
    .Q(\logo_top[8] ));
 sg13g2_dfrbp_1 _3190_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net60),
    .D(_0066_),
    .Q_N(_1531_),
    .Q(\logo_top[9] ));
 sg13g2_dfrbp_1 _3191_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net58),
    .D(_0067_),
    .Q_N(_1530_),
    .Q(dir_x));
 sg13g2_dfrbp_1 _3192_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net56),
    .D(_0068_),
    .Q_N(_1529_),
    .Q(dir_y));
 sg13g2_dfrbp_1 _3193_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net54),
    .D(net135),
    .Q_N(_0004_),
    .Q(manual_mode));
 sg13g2_dfrbp_1 _3194_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net52),
    .D(net137),
    .Q_N(_0018_),
    .Q(\color_index[0] ));
 sg13g2_dfrbp_1 _3195_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net50),
    .D(net214),
    .Q_N(_0016_),
    .Q(\color_index[1] ));
 sg13g2_dfrbp_1 _3196_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net48),
    .D(net139),
    .Q_N(_0015_),
    .Q(\color_index[2] ));
 sg13g2_dfrbp_1 _3197_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net46),
    .D(net172),
    .Q_N(_1528_),
    .Q(\prev_y[0] ));
 sg13g2_dfrbp_1 _3198_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net45),
    .D(_0074_),
    .Q_N(_1527_),
    .Q(\prev_y[1] ));
 sg13g2_dfrbp_1 _3199_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net44),
    .D(net178),
    .Q_N(_1526_),
    .Q(\prev_y[2] ));
 sg13g2_dfrbp_1 _3200_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net43),
    .D(net174),
    .Q_N(_1525_),
    .Q(\prev_y[3] ));
 sg13g2_dfrbp_1 _3201_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net42),
    .D(_0077_),
    .Q_N(_1524_),
    .Q(\prev_y[4] ));
 sg13g2_dfrbp_1 _3202_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net41),
    .D(net168),
    .Q_N(_1523_),
    .Q(\prev_y[5] ));
 sg13g2_dfrbp_1 _3203_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net38),
    .D(net176),
    .Q_N(_1522_),
    .Q(\prev_y[6] ));
 sg13g2_dfrbp_1 _3204_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net36),
    .D(net180),
    .Q_N(_1521_),
    .Q(\prev_y[7] ));
 sg13g2_dfrbp_1 _3205_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net34),
    .D(net159),
    .Q_N(_1520_),
    .Q(\prev_y[8] ));
 sg13g2_dfrbp_1 _3206_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net32),
    .D(net188),
    .Q_N(_1519_),
    .Q(\prev_y[9] ));
 sg13g2_dfrbp_1 _3207_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net30),
    .D(_0083_),
    .Q_N(_1518_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _3208_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net28),
    .D(_0084_),
    .Q_N(_1517_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _3209_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net26),
    .D(_0085_),
    .Q_N(_1516_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _3210_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net88),
    .D(_0086_),
    .Q_N(_1565_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _3211_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net107),
    .D(net126),
    .Q_N(_1566_),
    .Q(\gamepad.driver.pmod_clk_prev ));
 sg13g2_dfrbp_1 _3212_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net24),
    .D(net125),
    .Q_N(_1515_),
    .Q(\gamepad.driver.pmod_latch_prev ));
 sg13g2_dfrbp_1 _3213_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net22),
    .D(net184),
    .Q_N(_1514_),
    .Q(\gamepad.driver.shift_reg[0] ));
 sg13g2_dfrbp_1 _3214_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net116),
    .D(net192),
    .Q_N(_1513_),
    .Q(\gamepad.driver.shift_reg[1] ));
 sg13g2_dfrbp_1 _3215_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net112),
    .D(net212),
    .Q_N(_1512_),
    .Q(\gamepad.driver.shift_reg[2] ));
 sg13g2_dfrbp_1 _3216_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net97),
    .D(net190),
    .Q_N(_1511_),
    .Q(\gamepad.driver.shift_reg[3] ));
 sg13g2_dfrbp_1 _3217_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net93),
    .D(_0091_),
    .Q_N(_1510_),
    .Q(\gamepad.driver.shift_reg[4] ));
 sg13g2_dfrbp_1 _3218_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net89),
    .D(net204),
    .Q_N(_1509_),
    .Q(\gamepad.driver.shift_reg[5] ));
 sg13g2_dfrbp_1 _3219_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net83),
    .D(net199),
    .Q_N(_1508_),
    .Q(\gamepad.driver.shift_reg[6] ));
 sg13g2_dfrbp_1 _3220_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net79),
    .D(net194),
    .Q_N(_1507_),
    .Q(\gamepad.driver.shift_reg[7] ));
 sg13g2_dfrbp_1 _3221_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net75),
    .D(_0095_),
    .Q_N(_1506_),
    .Q(\gamepad.driver.shift_reg[8] ));
 sg13g2_dfrbp_1 _3222_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net71),
    .D(_0096_),
    .Q_N(_1505_),
    .Q(\gamepad.driver.shift_reg[9] ));
 sg13g2_dfrbp_1 _3223_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net67),
    .D(net202),
    .Q_N(_1504_),
    .Q(\gamepad.driver.shift_reg[10] ));
 sg13g2_dfrbp_1 _3224_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net63),
    .D(net162),
    .Q_N(_1503_),
    .Q(\gamepad.driver.shift_reg[11] ));
 sg13g2_dfrbp_1 _3225_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net59),
    .D(_0099_),
    .Q_N(_1502_),
    .Q(\gamepad.driver.pmod_data_sync[0] ));
 sg13g2_dfrbp_1 _3226_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net57),
    .D(_0100_),
    .Q_N(_1501_),
    .Q(\gamepad.driver.pmod_data_sync[1] ));
 sg13g2_dfrbp_1 _3227_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net55),
    .D(_0101_),
    .Q_N(_1500_),
    .Q(\gamepad.driver.pmod_clk_sync[0] ));
 sg13g2_dfrbp_1 _3228_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net53),
    .D(_0102_),
    .Q_N(_1499_),
    .Q(\gamepad.driver.pmod_clk_sync[1] ));
 sg13g2_dfrbp_1 _3229_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net51),
    .D(_0103_),
    .Q_N(_1498_),
    .Q(\gamepad.driver.pmod_latch_sync[0] ));
 sg13g2_dfrbp_1 _3230_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net118),
    .D(_0104_),
    .Q_N(_1567_),
    .Q(\gamepad.driver.pmod_latch_sync[1] ));
 sg13g2_dfrbp_1 _3231_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net49),
    .D(net223),
    .Q_N(_1497_),
    .Q(hsync));
 sg13g2_dfrbp_1 _3232_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net47),
    .D(net129),
    .Q_N(_0017_),
    .Q(\pix_y[0] ));
 sg13g2_dfrbp_1 _3233_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net114),
    .D(_0106_),
    .Q_N(_1496_),
    .Q(\pix_y[1] ));
 sg13g2_dfrbp_1 _3234_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net95),
    .D(_0107_),
    .Q_N(_1495_),
    .Q(\pix_y[2] ));
 sg13g2_dfrbp_1 _3235_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net85),
    .D(net182),
    .Q_N(_1494_),
    .Q(\pix_y[3] ));
 sg13g2_dfrbp_1 _3236_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net77),
    .D(_0109_),
    .Q_N(_1493_),
    .Q(\pix_y[4] ));
 sg13g2_dfrbp_1 _3237_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net69),
    .D(_0110_),
    .Q_N(_1492_),
    .Q(\pix_y[5] ));
 sg13g2_dfrbp_1 _3238_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net61),
    .D(_0111_),
    .Q_N(_1491_),
    .Q(\pix_y[6] ));
 sg13g2_dfrbp_1 _3239_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net99),
    .D(_0112_),
    .Q_N(_1490_),
    .Q(\pix_y[7] ));
 sg13g2_dfrbp_1 _3240_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net81),
    .D(_0113_),
    .Q_N(_1489_),
    .Q(\pix_y[8] ));
 sg13g2_dfrbp_1 _3241_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net119),
    .D(_0114_),
    .Q_N(_1568_),
    .Q(\pix_y[9] ));
 sg13g2_dfrbp_1 _3242_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net120),
    .D(_0006_),
    .Q_N(_1569_),
    .Q(\vga_sync_gen.vsync ));
 sg13g2_dfrbp_1 _3243_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net121),
    .D(_0000_),
    .Q_N(_1570_),
    .Q(\palette_inst.rrggbb[0] ));
 sg13g2_dfrbp_1 _3244_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net122),
    .D(_0001_),
    .Q_N(_1571_),
    .Q(\palette_inst.rrggbb[1] ));
 sg13g2_dfrbp_1 _3245_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net123),
    .D(_0002_),
    .Q_N(_1572_),
    .Q(\palette_inst.rrggbb[2] ));
 sg13g2_dfrbp_1 _3246_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net65),
    .D(_0003_),
    .Q_N(_1488_),
    .Q(\palette_inst.rrggbb[3] ));
 sg13g2_dfrbp_1 _3247_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net91),
    .D(_0115_),
    .Q_N(_1487_),
    .Q(\palette_inst.rrggbb[4] ));
 sg13g2_dfrbp_1 _3248_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net73),
    .D(_0116_),
    .Q_N(_1486_),
    .Q(\palette_inst.rrggbb[5] ));
 sg13g2_tiehi _3156__23 (.L_HI(net23));
 sg13g2_tiehi _3212__24 (.L_HI(net24));
 sg13g2_tiehi _3155__25 (.L_HI(net25));
 sg13g2_tiehi _3209__26 (.L_HI(net26));
 sg13g2_tiehi _3154__27 (.L_HI(net27));
 sg13g2_tiehi _3208__28 (.L_HI(net28));
 sg13g2_tiehi _3153__29 (.L_HI(net29));
 sg13g2_tiehi _3207__30 (.L_HI(net30));
 sg13g2_tiehi _3152__31 (.L_HI(net31));
 sg13g2_tiehi _3206__32 (.L_HI(net32));
 sg13g2_tiehi _3151__33 (.L_HI(net33));
 sg13g2_tiehi _3205__34 (.L_HI(net34));
 sg13g2_tiehi _3150__35 (.L_HI(net35));
 sg13g2_tiehi _3204__36 (.L_HI(net36));
 sg13g2_tiehi _3149__37 (.L_HI(net37));
 sg13g2_tiehi _3203__38 (.L_HI(net38));
 sg13g2_tiehi _3148__39 (.L_HI(net39));
 sg13g2_tiehi _3147__40 (.L_HI(net40));
 sg13g2_tiehi _3202__41 (.L_HI(net41));
 sg13g2_tiehi _3201__42 (.L_HI(net42));
 sg13g2_tiehi _3200__43 (.L_HI(net43));
 sg13g2_tiehi _3199__44 (.L_HI(net44));
 sg13g2_tiehi _3198__45 (.L_HI(net45));
 sg13g2_tiehi _3197__46 (.L_HI(net46));
 sg13g2_tiehi _3232__47 (.L_HI(net47));
 sg13g2_tiehi _3196__48 (.L_HI(net48));
 sg13g2_tiehi _3231__49 (.L_HI(net49));
 sg13g2_tiehi _3195__50 (.L_HI(net50));
 sg13g2_tiehi _3229__51 (.L_HI(net51));
 sg13g2_tiehi _3194__52 (.L_HI(net52));
 sg13g2_tiehi _3228__53 (.L_HI(net53));
 sg13g2_tiehi _3193__54 (.L_HI(net54));
 sg13g2_tiehi _3227__55 (.L_HI(net55));
 sg13g2_tiehi _3192__56 (.L_HI(net56));
 sg13g2_tiehi _3226__57 (.L_HI(net57));
 sg13g2_tiehi _3191__58 (.L_HI(net58));
 sg13g2_tiehi _3225__59 (.L_HI(net59));
 sg13g2_tiehi _3190__60 (.L_HI(net60));
 sg13g2_tiehi _3238__61 (.L_HI(net61));
 sg13g2_tiehi _3189__62 (.L_HI(net62));
 sg13g2_tiehi _3224__63 (.L_HI(net63));
 sg13g2_tiehi _3188__64 (.L_HI(net64));
 sg13g2_tiehi _3246__65 (.L_HI(net65));
 sg13g2_tiehi _3187__66 (.L_HI(net66));
 sg13g2_tiehi _3223__67 (.L_HI(net67));
 sg13g2_tiehi _3186__68 (.L_HI(net68));
 sg13g2_tiehi _3237__69 (.L_HI(net69));
 sg13g2_tiehi _3185__70 (.L_HI(net70));
 sg13g2_tiehi _3222__71 (.L_HI(net71));
 sg13g2_tiehi _3184__72 (.L_HI(net72));
 sg13g2_tiehi _3248__73 (.L_HI(net73));
 sg13g2_tiehi _3183__74 (.L_HI(net74));
 sg13g2_tiehi _3221__75 (.L_HI(net75));
 sg13g2_tiehi _3182__76 (.L_HI(net76));
 sg13g2_tiehi _3236__77 (.L_HI(net77));
 sg13g2_tiehi _3181__78 (.L_HI(net78));
 sg13g2_tiehi _3220__79 (.L_HI(net79));
 sg13g2_tiehi _3180__80 (.L_HI(net80));
 sg13g2_tiehi _3240__81 (.L_HI(net81));
 sg13g2_tiehi _3179__82 (.L_HI(net82));
 sg13g2_tiehi _3219__83 (.L_HI(net83));
 sg13g2_tiehi _3178__84 (.L_HI(net84));
 sg13g2_tiehi _3235__85 (.L_HI(net85));
 sg13g2_tiehi _3177__86 (.L_HI(net86));
 sg13g2_tiehi _3146__87 (.L_HI(net87));
 sg13g2_tiehi _3210__88 (.L_HI(net88));
 sg13g2_tiehi _3218__89 (.L_HI(net89));
 sg13g2_tiehi _3176__90 (.L_HI(net90));
 sg13g2_tiehi _3247__91 (.L_HI(net91));
 sg13g2_tiehi _3175__92 (.L_HI(net92));
 sg13g2_tiehi _3217__93 (.L_HI(net93));
 sg13g2_tiehi _3174__94 (.L_HI(net94));
 sg13g2_tiehi _3234__95 (.L_HI(net95));
 sg13g2_tiehi _3173__96 (.L_HI(net96));
 sg13g2_tiehi _3216__97 (.L_HI(net97));
 sg13g2_tiehi _3172__98 (.L_HI(net98));
 sg13g2_tiehi _3239__99 (.L_HI(net99));
 sg13g2_tiehi _3171__100 (.L_HI(net100));
 sg13g2_tiehi _3170__101 (.L_HI(net101));
 sg13g2_tiehi _3169__102 (.L_HI(net102));
 sg13g2_tiehi _3168__103 (.L_HI(net103));
 sg13g2_tiehi _3167__104 (.L_HI(net104));
 sg13g2_tiehi _3166__105 (.L_HI(net105));
 sg13g2_tiehi _3165__106 (.L_HI(net106));
 sg13g2_tiehi _3211__107 (.L_HI(net107));
 sg13g2_tiehi _3164__108 (.L_HI(net108));
 sg13g2_tiehi _3163__109 (.L_HI(net109));
 sg13g2_tiehi _3162__110 (.L_HI(net110));
 sg13g2_tiehi _3161__111 (.L_HI(net111));
 sg13g2_tiehi _3215__112 (.L_HI(net112));
 sg13g2_tiehi _3160__113 (.L_HI(net113));
 sg13g2_tiehi _3233__114 (.L_HI(net114));
 sg13g2_tiehi _3159__115 (.L_HI(net115));
 sg13g2_tiehi _3214__116 (.L_HI(net116));
 sg13g2_tiehi _3158__117 (.L_HI(net117));
 sg13g2_tiehi _3230__118 (.L_HI(net118));
 sg13g2_tiehi _3241__119 (.L_HI(net119));
 sg13g2_tiehi _3242__120 (.L_HI(net120));
 sg13g2_tiehi _3243__121 (.L_HI(net121));
 sg13g2_tiehi _3244__122 (.L_HI(net122));
 sg13g2_tiehi _3245__123 (.L_HI(net123));
 sg13g2_tiehi _3157__124 (.L_HI(net124));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_7 (.L_LO(net7));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_8 (.L_LO(net8));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_9 (.L_LO(net9));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_10 (.L_LO(net10));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_11 (.L_LO(net11));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_12 (.L_LO(net12));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_13 (.L_LO(net13));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_14 (.L_LO(net14));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_15 (.L_LO(net15));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_16 (.L_LO(net16));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_17 (.L_LO(net17));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_18 (.L_LO(net18));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_19 (.L_LO(net19));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_20 (.L_LO(net20));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_21 (.L_LO(net21));
 sg13g2_tiehi _3213__22 (.L_HI(net22));
 sg13g2_buf_1 _3368_ (.A(\vga_sync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _3369_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout612 (.A(_0867_),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(_0569_),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(_0569_),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(_0471_),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(_0470_),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(_0556_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_0556_),
    .X(net618));
 sg13g2_buf_4 fanout619 (.X(net619),
    .A(_0909_));
 sg13g2_buf_2 fanout620 (.A(_0908_),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(_0468_),
    .X(net621));
 sg13g2_buf_4 fanout622 (.X(net622),
    .A(_1029_));
 sg13g2_buf_2 fanout623 (.A(net624),
    .X(net623));
 sg13g2_buf_4 fanout624 (.X(net624),
    .A(_1028_));
 sg13g2_buf_2 fanout625 (.A(_1028_),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(_1181_),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(_1110_),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(net629),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(_1105_),
    .X(net629));
 sg13g2_buf_4 fanout630 (.X(net630),
    .A(_1074_));
 sg13g2_buf_2 fanout631 (.A(_1074_),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(net633),
    .X(net632));
 sg13g2_buf_1 fanout633 (.A(_1058_),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(net636),
    .X(net634));
 sg13g2_buf_1 fanout635 (.A(net636),
    .X(net635));
 sg13g2_buf_1 fanout636 (.A(_1053_),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(net638),
    .X(net637));
 sg13g2_buf_4 fanout638 (.X(net638),
    .A(_1052_));
 sg13g2_buf_4 fanout639 (.X(net639),
    .A(net640));
 sg13g2_buf_4 fanout640 (.X(net640),
    .A(_1043_));
 sg13g2_buf_4 fanout641 (.X(net641),
    .A(_1040_));
 sg13g2_buf_2 fanout642 (.A(_1040_),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(_1037_),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(net645),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(_1009_),
    .X(net645));
 sg13g2_buf_4 fanout646 (.X(net646),
    .A(_0973_));
 sg13g2_buf_2 fanout647 (.A(net649),
    .X(net647));
 sg13g2_buf_4 fanout648 (.X(net648),
    .A(net649));
 sg13g2_buf_2 fanout649 (.A(_0972_),
    .X(net649));
 sg13g2_buf_4 fanout650 (.X(net650),
    .A(_0968_));
 sg13g2_buf_2 fanout651 (.A(_0968_),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(net653),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(net654),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(_0966_),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(net656),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(net659),
    .X(net656));
 sg13g2_buf_4 fanout657 (.X(net657),
    .A(net659));
 sg13g2_buf_4 fanout658 (.X(net658),
    .A(net659));
 sg13g2_buf_4 fanout659 (.X(net659),
    .A(_0944_));
 sg13g2_buf_4 fanout660 (.X(net660),
    .A(net661));
 sg13g2_buf_4 fanout661 (.X(net661),
    .A(net662));
 sg13g2_buf_2 fanout662 (.A(_0943_),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(_0911_),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(_0911_),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(net666),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(_0911_),
    .X(net666));
 sg13g2_buf_4 fanout667 (.X(net667),
    .A(net668));
 sg13g2_buf_4 fanout668 (.X(net668),
    .A(_0910_));
 sg13g2_buf_4 fanout669 (.X(net669),
    .A(net671));
 sg13g2_buf_1 fanout670 (.A(net671),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(_0910_),
    .X(net671));
 sg13g2_buf_4 fanout672 (.X(net672),
    .A(_0449_));
 sg13g2_buf_4 fanout673 (.X(net673),
    .A(_1021_));
 sg13g2_buf_4 fanout674 (.X(net674),
    .A(net675));
 sg13g2_buf_4 fanout675 (.X(net675),
    .A(_1020_));
 sg13g2_buf_2 fanout676 (.A(_0963_),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(_0963_),
    .X(net677));
 sg13g2_buf_4 fanout678 (.X(net678),
    .A(net680));
 sg13g2_buf_2 fanout679 (.A(net680),
    .X(net679));
 sg13g2_buf_4 fanout680 (.X(net680),
    .A(_0956_));
 sg13g2_buf_2 fanout681 (.A(net682),
    .X(net681));
 sg13g2_buf_4 fanout682 (.X(net682),
    .A(_0956_));
 sg13g2_buf_4 fanout683 (.X(net683),
    .A(_0955_));
 sg13g2_buf_2 fanout684 (.A(_0955_),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(net687),
    .X(net685));
 sg13g2_buf_1 fanout686 (.A(net687),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(_0955_),
    .X(net687));
 sg13g2_buf_4 fanout688 (.X(net688),
    .A(_0950_));
 sg13g2_buf_2 fanout689 (.A(net690),
    .X(net689));
 sg13g2_buf_1 fanout690 (.A(_0942_),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(net692),
    .X(net691));
 sg13g2_buf_1 fanout692 (.A(_0941_),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(_0940_),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(_0940_),
    .X(net694));
 sg13g2_buf_2 fanout695 (.A(net697),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(net697),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(_0938_),
    .X(net697));
 sg13g2_buf_4 fanout698 (.X(net698),
    .A(net699));
 sg13g2_buf_4 fanout699 (.X(net699),
    .A(_1018_));
 sg13g2_buf_4 fanout700 (.X(net700),
    .A(_1013_));
 sg13g2_buf_2 fanout701 (.A(_1013_),
    .X(net701));
 sg13g2_buf_2 fanout702 (.A(net703),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(_1012_),
    .X(net703));
 sg13g2_buf_4 fanout704 (.X(net704),
    .A(_1012_));
 sg13g2_buf_2 fanout705 (.A(_1012_),
    .X(net705));
 sg13g2_buf_4 fanout706 (.X(net706),
    .A(_0992_));
 sg13g2_buf_4 fanout707 (.X(net707),
    .A(net708));
 sg13g2_buf_4 fanout708 (.X(net708),
    .A(_0946_));
 sg13g2_buf_4 fanout709 (.X(net709),
    .A(_0945_));
 sg13g2_buf_2 fanout710 (.A(net711),
    .X(net710));
 sg13g2_buf_4 fanout711 (.X(net711),
    .A(_0945_));
 sg13g2_buf_2 fanout712 (.A(net714),
    .X(net712));
 sg13g2_buf_2 fanout713 (.A(net714),
    .X(net713));
 sg13g2_buf_2 fanout714 (.A(net715),
    .X(net714));
 sg13g2_buf_4 fanout715 (.X(net715),
    .A(_0913_));
 sg13g2_buf_2 fanout716 (.A(net719),
    .X(net716));
 sg13g2_buf_2 fanout717 (.A(net718),
    .X(net717));
 sg13g2_buf_2 fanout718 (.A(net719),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(_0913_),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(net726),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(net726),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(net724),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(net724),
    .X(net723));
 sg13g2_buf_2 fanout724 (.A(net726),
    .X(net724));
 sg13g2_buf_4 fanout725 (.X(net725),
    .A(net726));
 sg13g2_buf_2 fanout726 (.A(_0912_),
    .X(net726));
 sg13g2_buf_4 fanout727 (.X(net727),
    .A(_1065_));
 sg13g2_buf_2 fanout728 (.A(net735),
    .X(net728));
 sg13g2_buf_1 fanout729 (.A(net735),
    .X(net729));
 sg13g2_buf_4 fanout730 (.X(net730),
    .A(net731));
 sg13g2_buf_2 fanout731 (.A(net735),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(net734),
    .X(net732));
 sg13g2_buf_4 fanout733 (.X(net733),
    .A(net734));
 sg13g2_buf_2 fanout734 (.A(net735),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(_0988_),
    .X(net735));
 sg13g2_buf_2 fanout736 (.A(net739),
    .X(net736));
 sg13g2_buf_4 fanout737 (.X(net737),
    .A(net738));
 sg13g2_buf_2 fanout738 (.A(net739),
    .X(net738));
 sg13g2_buf_4 fanout739 (.X(net739),
    .A(_0987_));
 sg13g2_buf_2 fanout740 (.A(_0987_),
    .X(net740));
 sg13g2_buf_2 fanout741 (.A(_0987_),
    .X(net741));
 sg13g2_buf_4 fanout742 (.X(net742),
    .A(_0981_));
 sg13g2_buf_4 fanout743 (.X(net743),
    .A(_0980_));
 sg13g2_buf_4 fanout744 (.X(net744),
    .A(_0687_));
 sg13g2_buf_2 fanout745 (.A(_0687_),
    .X(net745));
 sg13g2_buf_4 fanout746 (.X(net746),
    .A(_0436_));
 sg13g2_buf_1 fanout747 (.A(_0436_),
    .X(net747));
 sg13g2_buf_4 fanout748 (.X(net748),
    .A(net749));
 sg13g2_buf_4 fanout749 (.X(net749),
    .A(_0915_));
 sg13g2_buf_4 fanout750 (.X(net750),
    .A(_0915_));
 sg13g2_buf_2 fanout751 (.A(_0915_),
    .X(net751));
 sg13g2_buf_4 fanout752 (.X(net752),
    .A(net758));
 sg13g2_buf_2 fanout753 (.A(net754),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(net755),
    .X(net754));
 sg13g2_buf_1 fanout755 (.A(net758),
    .X(net755));
 sg13g2_buf_4 fanout756 (.X(net756),
    .A(net757));
 sg13g2_buf_4 fanout757 (.X(net757),
    .A(net758));
 sg13g2_buf_2 fanout758 (.A(_0914_),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(_0686_),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(_0686_),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(_0435_),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(_0435_),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(net764),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(net768),
    .X(net764));
 sg13g2_buf_4 fanout765 (.X(net765),
    .A(net767));
 sg13g2_buf_1 fanout766 (.A(net767),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(net768),
    .X(net767));
 sg13g2_buf_4 fanout768 (.X(net768),
    .A(_0977_));
 sg13g2_buf_4 fanout769 (.X(net769),
    .A(net772));
 sg13g2_buf_2 fanout770 (.A(net772),
    .X(net770));
 sg13g2_buf_4 fanout771 (.X(net771),
    .A(net772));
 sg13g2_buf_4 fanout772 (.X(net772),
    .A(_0976_));
 sg13g2_buf_2 fanout773 (.A(net774),
    .X(net773));
 sg13g2_buf_4 fanout774 (.X(net774),
    .A(_0976_));
 sg13g2_buf_2 fanout775 (.A(net776),
    .X(net775));
 sg13g2_buf_4 fanout776 (.X(net776),
    .A(_0724_));
 sg13g2_buf_2 fanout777 (.A(net185),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(net156),
    .X(net778));
 sg13g2_buf_4 fanout779 (.X(net779),
    .A(net181));
 sg13g2_buf_2 fanout780 (.A(net237),
    .X(net780));
 sg13g2_buf_4 fanout781 (.X(net781),
    .A(net146));
 sg13g2_buf_2 fanout782 (.A(net785),
    .X(net782));
 sg13g2_buf_1 fanout783 (.A(net785),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(net785),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(net242),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(net788),
    .X(net786));
 sg13g2_buf_2 fanout787 (.A(net788),
    .X(net787));
 sg13g2_buf_4 fanout788 (.X(net788),
    .A(dir_y));
 sg13g2_buf_4 fanout789 (.X(net789),
    .A(net790));
 sg13g2_buf_4 fanout790 (.X(net790),
    .A(dir_x));
 sg13g2_buf_2 fanout791 (.A(net262),
    .X(net791));
 sg13g2_buf_2 fanout792 (.A(net261),
    .X(net792));
 sg13g2_buf_4 fanout793 (.X(net793),
    .A(net248));
 sg13g2_buf_2 fanout794 (.A(\logo_top[4] ),
    .X(net794));
 sg13g2_buf_4 fanout795 (.X(net795),
    .A(net254));
 sg13g2_buf_2 fanout796 (.A(\logo_top[1] ),
    .X(net796));
 sg13g2_buf_2 fanout797 (.A(\logo_top[0] ),
    .X(net797));
 sg13g2_buf_2 fanout798 (.A(net259),
    .X(net798));
 sg13g2_buf_4 fanout799 (.X(net799),
    .A(net258));
 sg13g2_buf_2 fanout800 (.A(\logo_left[3] ),
    .X(net800));
 sg13g2_buf_4 fanout801 (.X(net801),
    .A(net253));
 sg13g2_buf_4 fanout802 (.X(net802),
    .A(\logo_left[0] ));
 sg13g2_buf_2 fanout803 (.A(net249),
    .X(net803));
 sg13g2_buf_4 fanout804 (.X(net804),
    .A(net805));
 sg13g2_buf_4 fanout805 (.X(net805),
    .A(_0743_));
 sg13g2_buf_4 fanout806 (.X(net806),
    .A(net807));
 sg13g2_buf_4 fanout807 (.X(net807),
    .A(net813));
 sg13g2_buf_2 fanout808 (.A(net809),
    .X(net808));
 sg13g2_buf_4 fanout809 (.X(net809),
    .A(net813));
 sg13g2_buf_2 fanout810 (.A(net811),
    .X(net810));
 sg13g2_buf_2 fanout811 (.A(net812),
    .X(net811));
 sg13g2_buf_1 fanout812 (.A(net813),
    .X(net812));
 sg13g2_buf_2 fanout813 (.A(rst_n),
    .X(net813));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[4]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[5]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[6]),
    .X(net5));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_6 (.L_LO(net6));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\gamepad.driver.pmod_latch_sync[1] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold2 (.A(\gamepad.driver.pmod_clk_sync[1] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0021_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0017_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0105_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold6 (.A(\gamepad.driver.pmod_clk_sync[0] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold7 (.A(\gamepad.driver.pmod_data_sync[0] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0020_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0004_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0665_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0069_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0018_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0070_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold14 (.A(\color_index[2] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0072_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold16 (.A(gamepad_start_prev),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0036_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold18 (.A(\gamepad.decoder.data_reg[10] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0034_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold20 (.A(\gamepad.decoder.data_reg[2] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0026_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold22 (.A(\pix_y[1] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0692_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold24 (.A(\gamepad.decoder.data_reg[0] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0024_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold26 (.A(\gamepad.decoder.data_reg[3] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0027_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold28 (.A(\gamepad.decoder.data_reg[1] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0025_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold30 (.A(\gamepad.decoder.data_reg[9] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0033_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold32 (.A(\pix_y[4] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold33 (.A(\gamepad.driver.pmod_latch_sync[0] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold34 (.A(\prev_y[8] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0081_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold36 (.A(\prev_y[4] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold37 (.A(\gamepad.driver.shift_reg[11] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0098_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold39 (.A(\gamepad.decoder.data_reg[6] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0030_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold41 (.A(\gamepad.decoder.data_reg[8] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0032_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold43 (.A(\prev_y[5] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0078_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold45 (.A(\gamepad.decoder.data_reg[11] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0035_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold47 (.A(\prev_y[0] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0073_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold49 (.A(\prev_y[3] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0076_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold51 (.A(\prev_y[6] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0079_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold53 (.A(\prev_y[2] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0075_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold55 (.A(\prev_y[7] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0080_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold57 (.A(\pix_y[3] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0108_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold59 (.A(\gamepad.driver.shift_reg[0] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0087_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold61 (.A(\pix_y[7] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold62 (.A(\prev_y[1] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold63 (.A(\prev_y[9] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0082_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold65 (.A(\gamepad.driver.shift_reg[3] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0090_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold67 (.A(\gamepad.driver.shift_reg[1] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0088_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold69 (.A(\gamepad.driver.shift_reg[7] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0094_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0019_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0057_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold73 (.A(\gamepad.driver.shift_reg[8] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold74 (.A(\gamepad.driver.shift_reg[6] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0093_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold76 (.A(\gamepad.decoder.data_reg[7] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold77 (.A(\gamepad.driver.shift_reg[10] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0097_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold79 (.A(\gamepad.driver.shift_reg[5] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0092_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold81 (.A(\gamepad.driver.shift_reg[9] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold82 (.A(\gamepad.decoder.data_reg[5] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0029_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold84 (.A(\gamepad.decoder.data_reg[4] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0028_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold86 (.A(\gamepad.driver.shift_reg[4] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold87 (.A(\gamepad.driver.shift_reg[2] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0089_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold89 (.A(\color_index[1] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0071_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold91 (.A(\palette_inst.rrggbb[3] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold92 (.A(\pix_x[8] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0459_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold94 (.A(\pix_x[2] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0451_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0039_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold97 (.A(\pix_x[9] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0768_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0005_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold100 (.A(\pix_x[1] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0450_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0015_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold103 (.A(\palette_inst.rrggbb[5] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold104 (.A(\palette_inst.rrggbb[2] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold105 (.A(\palette_inst.rrggbb[0] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold106 (.A(\pix_x[6] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0456_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold108 (.A(\palette_inst.rrggbb[4] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold109 (.A(\pix_x[3] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0452_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold111 (.A(\pix_x[7] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0460_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold113 (.A(\pix_y[2] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold114 (.A(\pix_y[5] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold115 (.A(\pix_y[9] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold116 (.A(\palette_inst.rrggbb[1] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold117 (.A(\pix_x[4] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold118 (.A(manual_mode),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0061_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold120 (.A(\logo_top[8] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold121 (.A(\pix_y[8] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0764_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold123 (.A(\pix_y[6] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold124 (.A(\logo_top[5] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold125 (.A(\pix_x[5] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold126 (.A(\logo_top[3] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0016_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold128 (.A(\logo_left[6] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold129 (.A(\logo_left[1] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold130 (.A(\logo_top[2] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold131 (.A(\logo_top[6] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold132 (.A(\logo_left[2] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold133 (.A(\logo_left[8] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold134 (.A(\logo_left[4] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold135 (.A(\logo_left[7] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold136 (.A(\logo_left[9] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold137 (.A(\logo_top[7] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold138 (.A(\logo_top[9] ),
    .X(net262));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_fill_2 FILLER_0_14 ();
 sg13g2_decap_4 FILLER_0_30 ();
 sg13g2_fill_1 FILLER_0_34 ();
 sg13g2_fill_2 FILLER_0_38 ();
 sg13g2_fill_1 FILLER_0_40 ();
 sg13g2_fill_2 FILLER_0_71 ();
 sg13g2_fill_2 FILLER_0_82 ();
 sg13g2_fill_1 FILLER_0_161 ();
 sg13g2_fill_1 FILLER_0_184 ();
 sg13g2_fill_2 FILLER_0_245 ();
 sg13g2_fill_2 FILLER_0_271 ();
 sg13g2_fill_2 FILLER_0_327 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_fill_2 FILLER_1_7 ();
 sg13g2_fill_2 FILLER_1_52 ();
 sg13g2_fill_1 FILLER_1_72 ();
 sg13g2_fill_2 FILLER_1_106 ();
 sg13g2_fill_1 FILLER_1_108 ();
 sg13g2_fill_2 FILLER_1_134 ();
 sg13g2_fill_1 FILLER_1_310 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_fill_2 FILLER_2_14 ();
 sg13g2_fill_1 FILLER_2_37 ();
 sg13g2_fill_2 FILLER_2_58 ();
 sg13g2_fill_2 FILLER_2_90 ();
 sg13g2_fill_2 FILLER_2_100 ();
 sg13g2_fill_1 FILLER_2_102 ();
 sg13g2_fill_2 FILLER_2_142 ();
 sg13g2_fill_1 FILLER_2_170 ();
 sg13g2_fill_1 FILLER_2_184 ();
 sg13g2_fill_1 FILLER_2_228 ();
 sg13g2_fill_1 FILLER_2_257 ();
 sg13g2_fill_2 FILLER_2_267 ();
 sg13g2_fill_2 FILLER_2_287 ();
 sg13g2_fill_1 FILLER_2_315 ();
 sg13g2_fill_1 FILLER_3_44 ();
 sg13g2_fill_2 FILLER_3_50 ();
 sg13g2_decap_8 FILLER_3_83 ();
 sg13g2_fill_2 FILLER_3_95 ();
 sg13g2_fill_1 FILLER_3_97 ();
 sg13g2_fill_2 FILLER_3_117 ();
 sg13g2_fill_1 FILLER_3_124 ();
 sg13g2_fill_1 FILLER_3_143 ();
 sg13g2_fill_2 FILLER_3_304 ();
 sg13g2_fill_2 FILLER_3_315 ();
 sg13g2_fill_2 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_95 ();
 sg13g2_decap_8 FILLER_4_103 ();
 sg13g2_fill_2 FILLER_4_110 ();
 sg13g2_fill_1 FILLER_4_131 ();
 sg13g2_fill_2 FILLER_4_176 ();
 sg13g2_fill_1 FILLER_4_207 ();
 sg13g2_fill_2 FILLER_4_217 ();
 sg13g2_fill_1 FILLER_4_246 ();
 sg13g2_fill_1 FILLER_4_303 ();
 sg13g2_fill_2 FILLER_4_312 ();
 sg13g2_fill_2 FILLER_4_328 ();
 sg13g2_fill_2 FILLER_4_362 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_4 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_16 ();
 sg13g2_fill_2 FILLER_5_23 ();
 sg13g2_fill_1 FILLER_5_25 ();
 sg13g2_decap_4 FILLER_5_58 ();
 sg13g2_fill_1 FILLER_5_62 ();
 sg13g2_fill_2 FILLER_5_67 ();
 sg13g2_fill_1 FILLER_5_91 ();
 sg13g2_fill_2 FILLER_5_104 ();
 sg13g2_fill_2 FILLER_5_125 ();
 sg13g2_fill_1 FILLER_5_140 ();
 sg13g2_fill_2 FILLER_5_167 ();
 sg13g2_fill_1 FILLER_5_225 ();
 sg13g2_fill_2 FILLER_5_251 ();
 sg13g2_fill_1 FILLER_5_279 ();
 sg13g2_fill_1 FILLER_5_314 ();
 sg13g2_fill_2 FILLER_5_350 ();
 sg13g2_fill_2 FILLER_5_361 ();
 sg13g2_decap_4 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_4 ();
 sg13g2_fill_2 FILLER_6_28 ();
 sg13g2_fill_2 FILLER_6_56 ();
 sg13g2_fill_2 FILLER_6_63 ();
 sg13g2_fill_2 FILLER_6_86 ();
 sg13g2_fill_1 FILLER_6_88 ();
 sg13g2_fill_2 FILLER_6_125 ();
 sg13g2_fill_1 FILLER_6_127 ();
 sg13g2_fill_1 FILLER_6_211 ();
 sg13g2_fill_2 FILLER_6_238 ();
 sg13g2_fill_1 FILLER_6_298 ();
 sg13g2_fill_1 FILLER_6_324 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_20 ();
 sg13g2_fill_1 FILLER_7_22 ();
 sg13g2_fill_2 FILLER_7_39 ();
 sg13g2_fill_1 FILLER_7_41 ();
 sg13g2_fill_1 FILLER_7_51 ();
 sg13g2_fill_1 FILLER_7_60 ();
 sg13g2_fill_1 FILLER_7_73 ();
 sg13g2_fill_2 FILLER_7_86 ();
 sg13g2_fill_1 FILLER_7_88 ();
 sg13g2_fill_2 FILLER_7_104 ();
 sg13g2_fill_1 FILLER_7_106 ();
 sg13g2_decap_8 FILLER_7_121 ();
 sg13g2_decap_8 FILLER_7_128 ();
 sg13g2_fill_2 FILLER_7_135 ();
 sg13g2_fill_1 FILLER_7_149 ();
 sg13g2_fill_2 FILLER_7_203 ();
 sg13g2_fill_1 FILLER_7_226 ();
 sg13g2_fill_1 FILLER_7_246 ();
 sg13g2_fill_1 FILLER_7_268 ();
 sg13g2_fill_1 FILLER_7_283 ();
 sg13g2_fill_1 FILLER_7_288 ();
 sg13g2_fill_1 FILLER_7_313 ();
 sg13g2_fill_1 FILLER_7_357 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_4 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_4 ();
 sg13g2_fill_2 FILLER_8_72 ();
 sg13g2_fill_1 FILLER_8_98 ();
 sg13g2_fill_1 FILLER_8_108 ();
 sg13g2_fill_1 FILLER_8_145 ();
 sg13g2_fill_2 FILLER_8_225 ();
 sg13g2_fill_2 FILLER_8_241 ();
 sg13g2_fill_1 FILLER_8_264 ();
 sg13g2_fill_2 FILLER_8_353 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_7 ();
 sg13g2_fill_1 FILLER_9_40 ();
 sg13g2_fill_1 FILLER_9_46 ();
 sg13g2_fill_1 FILLER_9_64 ();
 sg13g2_fill_1 FILLER_9_73 ();
 sg13g2_fill_2 FILLER_9_95 ();
 sg13g2_fill_1 FILLER_9_97 ();
 sg13g2_fill_1 FILLER_9_131 ();
 sg13g2_fill_2 FILLER_9_167 ();
 sg13g2_fill_1 FILLER_9_169 ();
 sg13g2_fill_1 FILLER_9_282 ();
 sg13g2_fill_1 FILLER_9_337 ();
 sg13g2_fill_2 FILLER_9_369 ();
 sg13g2_fill_2 FILLER_10_111 ();
 sg13g2_fill_1 FILLER_10_136 ();
 sg13g2_decap_4 FILLER_10_153 ();
 sg13g2_fill_1 FILLER_10_157 ();
 sg13g2_fill_2 FILLER_10_171 ();
 sg13g2_fill_2 FILLER_10_178 ();
 sg13g2_fill_1 FILLER_10_180 ();
 sg13g2_fill_1 FILLER_10_191 ();
 sg13g2_fill_2 FILLER_10_210 ();
 sg13g2_fill_2 FILLER_10_228 ();
 sg13g2_fill_2 FILLER_10_263 ();
 sg13g2_fill_2 FILLER_10_328 ();
 sg13g2_fill_2 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_7 ();
 sg13g2_fill_1 FILLER_11_122 ();
 sg13g2_fill_2 FILLER_11_158 ();
 sg13g2_fill_1 FILLER_11_160 ();
 sg13g2_fill_1 FILLER_11_182 ();
 sg13g2_fill_1 FILLER_11_188 ();
 sg13g2_fill_1 FILLER_11_194 ();
 sg13g2_fill_2 FILLER_11_199 ();
 sg13g2_fill_2 FILLER_11_322 ();
 sg13g2_fill_2 FILLER_11_360 ();
 sg13g2_fill_1 FILLER_11_390 ();
 sg13g2_fill_1 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_41 ();
 sg13g2_fill_1 FILLER_12_58 ();
 sg13g2_fill_1 FILLER_12_100 ();
 sg13g2_decap_8 FILLER_12_136 ();
 sg13g2_decap_8 FILLER_12_153 ();
 sg13g2_decap_4 FILLER_12_160 ();
 sg13g2_fill_2 FILLER_12_186 ();
 sg13g2_fill_1 FILLER_12_220 ();
 sg13g2_fill_2 FILLER_12_242 ();
 sg13g2_fill_1 FILLER_12_275 ();
 sg13g2_fill_2 FILLER_12_319 ();
 sg13g2_fill_1 FILLER_12_376 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_fill_2 FILLER_13_26 ();
 sg13g2_fill_1 FILLER_13_28 ();
 sg13g2_fill_1 FILLER_13_52 ();
 sg13g2_fill_2 FILLER_13_79 ();
 sg13g2_fill_1 FILLER_13_95 ();
 sg13g2_fill_1 FILLER_13_105 ();
 sg13g2_fill_2 FILLER_13_124 ();
 sg13g2_fill_2 FILLER_13_168 ();
 sg13g2_fill_2 FILLER_13_175 ();
 sg13g2_fill_2 FILLER_13_182 ();
 sg13g2_decap_4 FILLER_13_197 ();
 sg13g2_fill_2 FILLER_13_201 ();
 sg13g2_fill_1 FILLER_13_212 ();
 sg13g2_fill_1 FILLER_13_227 ();
 sg13g2_fill_1 FILLER_13_263 ();
 sg13g2_fill_1 FILLER_13_269 ();
 sg13g2_fill_2 FILLER_13_305 ();
 sg13g2_fill_1 FILLER_13_325 ();
 sg13g2_fill_2 FILLER_13_331 ();
 sg13g2_fill_1 FILLER_13_352 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_25 ();
 sg13g2_fill_1 FILLER_14_33 ();
 sg13g2_fill_2 FILLER_14_42 ();
 sg13g2_fill_1 FILLER_14_44 ();
 sg13g2_fill_1 FILLER_14_112 ();
 sg13g2_fill_1 FILLER_14_125 ();
 sg13g2_decap_4 FILLER_14_138 ();
 sg13g2_fill_2 FILLER_14_142 ();
 sg13g2_fill_2 FILLER_14_147 ();
 sg13g2_fill_1 FILLER_14_149 ();
 sg13g2_fill_1 FILLER_14_186 ();
 sg13g2_fill_2 FILLER_14_213 ();
 sg13g2_fill_2 FILLER_14_223 ();
 sg13g2_fill_1 FILLER_14_256 ();
 sg13g2_fill_2 FILLER_14_263 ();
 sg13g2_fill_1 FILLER_14_355 ();
 sg13g2_fill_1 FILLER_14_378 ();
 sg13g2_fill_2 FILLER_14_384 ();
 sg13g2_fill_2 FILLER_15_34 ();
 sg13g2_fill_1 FILLER_15_36 ();
 sg13g2_fill_1 FILLER_15_52 ();
 sg13g2_fill_2 FILLER_15_94 ();
 sg13g2_fill_2 FILLER_15_110 ();
 sg13g2_fill_2 FILLER_15_117 ();
 sg13g2_fill_1 FILLER_15_119 ();
 sg13g2_fill_1 FILLER_15_136 ();
 sg13g2_decap_4 FILLER_15_147 ();
 sg13g2_fill_2 FILLER_15_196 ();
 sg13g2_fill_2 FILLER_15_202 ();
 sg13g2_fill_1 FILLER_15_204 ();
 sg13g2_fill_1 FILLER_15_240 ();
 sg13g2_fill_1 FILLER_15_245 ();
 sg13g2_fill_2 FILLER_15_312 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_35 ();
 sg13g2_fill_1 FILLER_16_49 ();
 sg13g2_fill_1 FILLER_16_60 ();
 sg13g2_fill_1 FILLER_16_85 ();
 sg13g2_fill_1 FILLER_16_101 ();
 sg13g2_fill_1 FILLER_16_120 ();
 sg13g2_decap_4 FILLER_16_142 ();
 sg13g2_fill_2 FILLER_16_146 ();
 sg13g2_fill_1 FILLER_16_160 ();
 sg13g2_fill_2 FILLER_16_169 ();
 sg13g2_decap_8 FILLER_16_176 ();
 sg13g2_fill_1 FILLER_16_183 ();
 sg13g2_decap_4 FILLER_16_200 ();
 sg13g2_decap_8 FILLER_16_208 ();
 sg13g2_decap_4 FILLER_16_220 ();
 sg13g2_fill_2 FILLER_16_354 ();
 sg13g2_fill_2 FILLER_16_370 ();
 sg13g2_fill_2 FILLER_16_381 ();
 sg13g2_fill_2 FILLER_17_26 ();
 sg13g2_fill_1 FILLER_17_54 ();
 sg13g2_fill_1 FILLER_17_78 ();
 sg13g2_decap_8 FILLER_17_115 ();
 sg13g2_fill_2 FILLER_17_122 ();
 sg13g2_fill_1 FILLER_17_124 ();
 sg13g2_fill_2 FILLER_17_143 ();
 sg13g2_fill_1 FILLER_17_150 ();
 sg13g2_fill_2 FILLER_17_191 ();
 sg13g2_decap_8 FILLER_17_218 ();
 sg13g2_fill_2 FILLER_17_225 ();
 sg13g2_fill_2 FILLER_17_232 ();
 sg13g2_fill_1 FILLER_17_234 ();
 sg13g2_fill_2 FILLER_17_248 ();
 sg13g2_fill_1 FILLER_17_250 ();
 sg13g2_fill_1 FILLER_17_263 ();
 sg13g2_fill_2 FILLER_17_279 ();
 sg13g2_fill_2 FILLER_17_306 ();
 sg13g2_fill_2 FILLER_17_312 ();
 sg13g2_fill_1 FILLER_17_370 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_7 ();
 sg13g2_fill_1 FILLER_18_26 ();
 sg13g2_decap_8 FILLER_18_47 ();
 sg13g2_fill_2 FILLER_18_54 ();
 sg13g2_fill_1 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_81 ();
 sg13g2_fill_2 FILLER_18_88 ();
 sg13g2_fill_1 FILLER_18_90 ();
 sg13g2_fill_2 FILLER_18_104 ();
 sg13g2_decap_8 FILLER_18_116 ();
 sg13g2_fill_1 FILLER_18_123 ();
 sg13g2_fill_1 FILLER_18_149 ();
 sg13g2_fill_2 FILLER_18_163 ();
 sg13g2_decap_8 FILLER_18_170 ();
 sg13g2_decap_4 FILLER_18_177 ();
 sg13g2_decap_8 FILLER_18_191 ();
 sg13g2_fill_1 FILLER_18_198 ();
 sg13g2_fill_1 FILLER_18_220 ();
 sg13g2_fill_1 FILLER_18_250 ();
 sg13g2_fill_1 FILLER_18_292 ();
 sg13g2_fill_2 FILLER_18_319 ();
 sg13g2_fill_2 FILLER_18_333 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_4 ();
 sg13g2_fill_2 FILLER_19_23 ();
 sg13g2_decap_4 FILLER_19_39 ();
 sg13g2_decap_8 FILLER_19_61 ();
 sg13g2_decap_8 FILLER_19_68 ();
 sg13g2_decap_8 FILLER_19_75 ();
 sg13g2_fill_1 FILLER_19_102 ();
 sg13g2_fill_1 FILLER_19_124 ();
 sg13g2_fill_1 FILLER_19_131 ();
 sg13g2_fill_2 FILLER_19_141 ();
 sg13g2_decap_4 FILLER_19_153 ();
 sg13g2_fill_2 FILLER_19_163 ();
 sg13g2_fill_1 FILLER_19_165 ();
 sg13g2_fill_2 FILLER_19_202 ();
 sg13g2_fill_2 FILLER_19_209 ();
 sg13g2_decap_4 FILLER_19_227 ();
 sg13g2_fill_1 FILLER_19_252 ();
 sg13g2_decap_4 FILLER_19_258 ();
 sg13g2_fill_2 FILLER_19_262 ();
 sg13g2_fill_2 FILLER_19_280 ();
 sg13g2_fill_1 FILLER_19_365 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_9 ();
 sg13g2_fill_1 FILLER_20_25 ();
 sg13g2_decap_4 FILLER_20_77 ();
 sg13g2_fill_2 FILLER_20_81 ();
 sg13g2_decap_8 FILLER_20_92 ();
 sg13g2_decap_8 FILLER_20_99 ();
 sg13g2_fill_2 FILLER_20_106 ();
 sg13g2_fill_2 FILLER_20_117 ();
 sg13g2_fill_1 FILLER_20_124 ();
 sg13g2_fill_2 FILLER_20_136 ();
 sg13g2_fill_1 FILLER_20_170 ();
 sg13g2_decap_4 FILLER_20_175 ();
 sg13g2_fill_2 FILLER_20_179 ();
 sg13g2_decap_4 FILLER_20_188 ();
 sg13g2_fill_2 FILLER_20_192 ();
 sg13g2_fill_2 FILLER_20_199 ();
 sg13g2_fill_1 FILLER_20_201 ();
 sg13g2_fill_2 FILLER_20_208 ();
 sg13g2_fill_1 FILLER_20_210 ();
 sg13g2_fill_2 FILLER_20_216 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_fill_2 FILLER_20_231 ();
 sg13g2_fill_1 FILLER_20_233 ();
 sg13g2_decap_8 FILLER_20_263 ();
 sg13g2_fill_2 FILLER_20_270 ();
 sg13g2_fill_2 FILLER_20_280 ();
 sg13g2_fill_2 FILLER_20_302 ();
 sg13g2_fill_2 FILLER_20_352 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_4 ();
 sg13g2_fill_1 FILLER_21_31 ();
 sg13g2_decap_8 FILLER_21_43 ();
 sg13g2_decap_8 FILLER_21_50 ();
 sg13g2_fill_1 FILLER_21_57 ();
 sg13g2_decap_4 FILLER_21_99 ();
 sg13g2_fill_2 FILLER_21_114 ();
 sg13g2_fill_1 FILLER_21_116 ();
 sg13g2_fill_2 FILLER_21_124 ();
 sg13g2_fill_1 FILLER_21_126 ();
 sg13g2_fill_1 FILLER_21_144 ();
 sg13g2_fill_1 FILLER_21_166 ();
 sg13g2_fill_2 FILLER_21_178 ();
 sg13g2_fill_1 FILLER_21_198 ();
 sg13g2_fill_2 FILLER_21_217 ();
 sg13g2_decap_4 FILLER_21_232 ();
 sg13g2_fill_1 FILLER_21_236 ();
 sg13g2_fill_2 FILLER_21_249 ();
 sg13g2_decap_4 FILLER_21_255 ();
 sg13g2_fill_1 FILLER_21_259 ();
 sg13g2_fill_1 FILLER_21_270 ();
 sg13g2_decap_4 FILLER_21_276 ();
 sg13g2_fill_1 FILLER_21_280 ();
 sg13g2_fill_1 FILLER_21_286 ();
 sg13g2_decap_4 FILLER_21_291 ();
 sg13g2_fill_1 FILLER_21_295 ();
 sg13g2_fill_2 FILLER_21_311 ();
 sg13g2_fill_1 FILLER_21_352 ();
 sg13g2_fill_2 FILLER_21_367 ();
 sg13g2_fill_2 FILLER_21_378 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_4 ();
 sg13g2_fill_2 FILLER_22_24 ();
 sg13g2_fill_2 FILLER_22_70 ();
 sg13g2_fill_1 FILLER_22_77 ();
 sg13g2_fill_1 FILLER_22_89 ();
 sg13g2_fill_2 FILLER_22_95 ();
 sg13g2_decap_4 FILLER_22_102 ();
 sg13g2_fill_1 FILLER_22_106 ();
 sg13g2_fill_2 FILLER_22_127 ();
 sg13g2_fill_1 FILLER_22_129 ();
 sg13g2_decap_8 FILLER_22_137 ();
 sg13g2_decap_8 FILLER_22_144 ();
 sg13g2_fill_2 FILLER_22_151 ();
 sg13g2_fill_1 FILLER_22_153 ();
 sg13g2_fill_1 FILLER_22_158 ();
 sg13g2_decap_4 FILLER_22_163 ();
 sg13g2_fill_1 FILLER_22_167 ();
 sg13g2_fill_1 FILLER_22_178 ();
 sg13g2_fill_1 FILLER_22_186 ();
 sg13g2_fill_1 FILLER_22_213 ();
 sg13g2_fill_1 FILLER_22_231 ();
 sg13g2_fill_2 FILLER_22_264 ();
 sg13g2_fill_2 FILLER_22_276 ();
 sg13g2_fill_1 FILLER_22_297 ();
 sg13g2_fill_1 FILLER_22_323 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_7 ();
 sg13g2_fill_2 FILLER_23_11 ();
 sg13g2_decap_8 FILLER_23_65 ();
 sg13g2_fill_2 FILLER_23_77 ();
 sg13g2_fill_2 FILLER_23_84 ();
 sg13g2_fill_2 FILLER_23_124 ();
 sg13g2_fill_1 FILLER_23_126 ();
 sg13g2_decap_4 FILLER_23_143 ();
 sg13g2_decap_8 FILLER_23_160 ();
 sg13g2_fill_2 FILLER_23_178 ();
 sg13g2_fill_1 FILLER_23_180 ();
 sg13g2_decap_8 FILLER_23_202 ();
 sg13g2_fill_2 FILLER_23_209 ();
 sg13g2_fill_1 FILLER_23_234 ();
 sg13g2_fill_2 FILLER_23_244 ();
 sg13g2_decap_8 FILLER_23_251 ();
 sg13g2_decap_4 FILLER_23_258 ();
 sg13g2_decap_8 FILLER_23_279 ();
 sg13g2_fill_2 FILLER_23_294 ();
 sg13g2_fill_1 FILLER_23_296 ();
 sg13g2_fill_2 FILLER_23_309 ();
 sg13g2_fill_1 FILLER_23_357 ();
 sg13g2_fill_1 FILLER_23_363 ();
 sg13g2_fill_1 FILLER_23_368 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_decap_4 FILLER_24_23 ();
 sg13g2_fill_2 FILLER_24_27 ();
 sg13g2_fill_2 FILLER_24_44 ();
 sg13g2_fill_2 FILLER_24_50 ();
 sg13g2_fill_1 FILLER_24_52 ();
 sg13g2_fill_1 FILLER_24_62 ();
 sg13g2_fill_2 FILLER_24_68 ();
 sg13g2_fill_1 FILLER_24_78 ();
 sg13g2_decap_4 FILLER_24_101 ();
 sg13g2_fill_1 FILLER_24_105 ();
 sg13g2_decap_4 FILLER_24_111 ();
 sg13g2_fill_2 FILLER_24_128 ();
 sg13g2_fill_1 FILLER_24_130 ();
 sg13g2_fill_1 FILLER_24_141 ();
 sg13g2_fill_1 FILLER_24_152 ();
 sg13g2_fill_1 FILLER_24_159 ();
 sg13g2_fill_2 FILLER_24_178 ();
 sg13g2_fill_1 FILLER_24_180 ();
 sg13g2_decap_8 FILLER_24_204 ();
 sg13g2_fill_1 FILLER_24_211 ();
 sg13g2_fill_2 FILLER_24_219 ();
 sg13g2_fill_1 FILLER_24_221 ();
 sg13g2_decap_4 FILLER_24_235 ();
 sg13g2_fill_2 FILLER_24_255 ();
 sg13g2_fill_2 FILLER_24_268 ();
 sg13g2_fill_2 FILLER_24_292 ();
 sg13g2_fill_1 FILLER_24_312 ();
 sg13g2_fill_1 FILLER_24_329 ();
 sg13g2_fill_2 FILLER_24_338 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_9 ();
 sg13g2_decap_8 FILLER_25_20 ();
 sg13g2_fill_2 FILLER_25_27 ();
 sg13g2_fill_2 FILLER_25_50 ();
 sg13g2_fill_1 FILLER_25_52 ();
 sg13g2_fill_2 FILLER_25_80 ();
 sg13g2_fill_2 FILLER_25_110 ();
 sg13g2_fill_1 FILLER_25_112 ();
 sg13g2_decap_4 FILLER_25_125 ();
 sg13g2_fill_2 FILLER_25_134 ();
 sg13g2_fill_1 FILLER_25_136 ();
 sg13g2_fill_2 FILLER_25_147 ();
 sg13g2_fill_1 FILLER_25_149 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_4 FILLER_25_201 ();
 sg13g2_fill_1 FILLER_25_205 ();
 sg13g2_fill_1 FILLER_25_215 ();
 sg13g2_decap_8 FILLER_25_220 ();
 sg13g2_fill_2 FILLER_25_227 ();
 sg13g2_decap_8 FILLER_25_244 ();
 sg13g2_fill_2 FILLER_25_251 ();
 sg13g2_fill_2 FILLER_25_262 ();
 sg13g2_decap_8 FILLER_25_278 ();
 sg13g2_decap_4 FILLER_25_304 ();
 sg13g2_decap_4 FILLER_25_326 ();
 sg13g2_fill_2 FILLER_25_334 ();
 sg13g2_fill_2 FILLER_25_392 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_30 ();
 sg13g2_fill_2 FILLER_26_59 ();
 sg13g2_fill_1 FILLER_26_88 ();
 sg13g2_fill_1 FILLER_26_99 ();
 sg13g2_fill_2 FILLER_26_116 ();
 sg13g2_decap_8 FILLER_26_134 ();
 sg13g2_decap_4 FILLER_26_141 ();
 sg13g2_fill_1 FILLER_26_145 ();
 sg13g2_fill_1 FILLER_26_155 ();
 sg13g2_fill_1 FILLER_26_169 ();
 sg13g2_fill_2 FILLER_26_179 ();
 sg13g2_fill_1 FILLER_26_181 ();
 sg13g2_fill_2 FILLER_26_200 ();
 sg13g2_fill_1 FILLER_26_202 ();
 sg13g2_fill_2 FILLER_26_212 ();
 sg13g2_fill_2 FILLER_26_258 ();
 sg13g2_fill_1 FILLER_26_281 ();
 sg13g2_decap_4 FILLER_26_302 ();
 sg13g2_fill_1 FILLER_26_306 ();
 sg13g2_fill_2 FILLER_26_333 ();
 sg13g2_fill_1 FILLER_26_343 ();
 sg13g2_fill_1 FILLER_26_362 ();
 sg13g2_fill_2 FILLER_26_368 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_2 ();
 sg13g2_fill_2 FILLER_27_54 ();
 sg13g2_fill_2 FILLER_27_65 ();
 sg13g2_fill_2 FILLER_27_77 ();
 sg13g2_fill_1 FILLER_27_79 ();
 sg13g2_fill_2 FILLER_27_112 ();
 sg13g2_fill_2 FILLER_27_135 ();
 sg13g2_fill_1 FILLER_27_137 ();
 sg13g2_fill_1 FILLER_27_172 ();
 sg13g2_fill_2 FILLER_27_183 ();
 sg13g2_fill_1 FILLER_27_185 ();
 sg13g2_decap_8 FILLER_27_206 ();
 sg13g2_fill_2 FILLER_27_218 ();
 sg13g2_fill_2 FILLER_27_229 ();
 sg13g2_fill_1 FILLER_27_236 ();
 sg13g2_fill_1 FILLER_27_262 ();
 sg13g2_fill_2 FILLER_27_294 ();
 sg13g2_decap_4 FILLER_27_329 ();
 sg13g2_fill_1 FILLER_27_399 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_7 ();
 sg13g2_decap_4 FILLER_28_23 ();
 sg13g2_fill_2 FILLER_28_27 ();
 sg13g2_fill_2 FILLER_28_33 ();
 sg13g2_fill_1 FILLER_28_40 ();
 sg13g2_decap_8 FILLER_28_45 ();
 sg13g2_decap_4 FILLER_28_52 ();
 sg13g2_fill_1 FILLER_28_72 ();
 sg13g2_fill_2 FILLER_28_88 ();
 sg13g2_fill_2 FILLER_28_118 ();
 sg13g2_fill_1 FILLER_28_120 ();
 sg13g2_fill_2 FILLER_28_141 ();
 sg13g2_fill_1 FILLER_28_143 ();
 sg13g2_fill_2 FILLER_28_149 ();
 sg13g2_fill_2 FILLER_28_163 ();
 sg13g2_fill_1 FILLER_28_165 ();
 sg13g2_fill_2 FILLER_28_176 ();
 sg13g2_fill_1 FILLER_28_178 ();
 sg13g2_fill_2 FILLER_28_184 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_fill_2 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_227 ();
 sg13g2_fill_1 FILLER_28_242 ();
 sg13g2_decap_4 FILLER_28_250 ();
 sg13g2_decap_4 FILLER_28_270 ();
 sg13g2_fill_2 FILLER_28_282 ();
 sg13g2_fill_1 FILLER_28_284 ();
 sg13g2_decap_8 FILLER_28_297 ();
 sg13g2_fill_2 FILLER_28_304 ();
 sg13g2_fill_2 FILLER_28_314 ();
 sg13g2_fill_1 FILLER_28_316 ();
 sg13g2_fill_2 FILLER_28_355 ();
 sg13g2_fill_1 FILLER_28_366 ();
 sg13g2_fill_1 FILLER_28_384 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_fill_1 FILLER_29_30 ();
 sg13g2_fill_1 FILLER_29_48 ();
 sg13g2_decap_4 FILLER_29_87 ();
 sg13g2_decap_4 FILLER_29_97 ();
 sg13g2_fill_2 FILLER_29_111 ();
 sg13g2_fill_1 FILLER_29_113 ();
 sg13g2_fill_2 FILLER_29_120 ();
 sg13g2_fill_2 FILLER_29_127 ();
 sg13g2_fill_2 FILLER_29_143 ();
 sg13g2_fill_1 FILLER_29_145 ();
 sg13g2_fill_2 FILLER_29_198 ();
 sg13g2_fill_1 FILLER_29_200 ();
 sg13g2_fill_1 FILLER_29_213 ();
 sg13g2_decap_4 FILLER_29_234 ();
 sg13g2_fill_2 FILLER_29_243 ();
 sg13g2_decap_4 FILLER_29_260 ();
 sg13g2_fill_2 FILLER_29_297 ();
 sg13g2_fill_1 FILLER_29_299 ();
 sg13g2_fill_1 FILLER_29_312 ();
 sg13g2_fill_2 FILLER_29_340 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_4 FILLER_30_31 ();
 sg13g2_fill_1 FILLER_30_35 ();
 sg13g2_decap_4 FILLER_30_51 ();
 sg13g2_fill_1 FILLER_30_55 ();
 sg13g2_decap_4 FILLER_30_69 ();
 sg13g2_decap_8 FILLER_30_78 ();
 sg13g2_fill_1 FILLER_30_85 ();
 sg13g2_decap_4 FILLER_30_101 ();
 sg13g2_decap_4 FILLER_30_115 ();
 sg13g2_fill_1 FILLER_30_126 ();
 sg13g2_decap_4 FILLER_30_155 ();
 sg13g2_fill_1 FILLER_30_163 ();
 sg13g2_fill_2 FILLER_30_170 ();
 sg13g2_fill_1 FILLER_30_172 ();
 sg13g2_fill_2 FILLER_30_179 ();
 sg13g2_fill_1 FILLER_30_181 ();
 sg13g2_decap_4 FILLER_30_198 ();
 sg13g2_fill_2 FILLER_30_202 ();
 sg13g2_decap_4 FILLER_30_212 ();
 sg13g2_fill_1 FILLER_30_216 ();
 sg13g2_fill_2 FILLER_30_222 ();
 sg13g2_fill_2 FILLER_30_238 ();
 sg13g2_fill_1 FILLER_30_258 ();
 sg13g2_fill_2 FILLER_30_264 ();
 sg13g2_fill_1 FILLER_30_266 ();
 sg13g2_decap_8 FILLER_30_277 ();
 sg13g2_fill_1 FILLER_30_284 ();
 sg13g2_fill_1 FILLER_30_300 ();
 sg13g2_fill_1 FILLER_30_306 ();
 sg13g2_fill_1 FILLER_30_360 ();
 sg13g2_fill_1 FILLER_30_371 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_4 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_11 ();
 sg13g2_fill_2 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_58 ();
 sg13g2_fill_2 FILLER_31_69 ();
 sg13g2_fill_1 FILLER_31_71 ();
 sg13g2_fill_2 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_79 ();
 sg13g2_decap_4 FILLER_31_87 ();
 sg13g2_fill_2 FILLER_31_113 ();
 sg13g2_fill_1 FILLER_31_134 ();
 sg13g2_decap_4 FILLER_31_146 ();
 sg13g2_fill_1 FILLER_31_162 ();
 sg13g2_fill_2 FILLER_31_176 ();
 sg13g2_fill_1 FILLER_31_178 ();
 sg13g2_decap_4 FILLER_31_187 ();
 sg13g2_fill_1 FILLER_31_191 ();
 sg13g2_fill_1 FILLER_31_200 ();
 sg13g2_fill_2 FILLER_31_237 ();
 sg13g2_fill_1 FILLER_31_239 ();
 sg13g2_fill_1 FILLER_31_286 ();
 sg13g2_fill_2 FILLER_31_317 ();
 sg13g2_fill_1 FILLER_31_337 ();
 sg13g2_fill_1 FILLER_31_399 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_26 ();
 sg13g2_fill_1 FILLER_32_33 ();
 sg13g2_decap_4 FILLER_32_52 ();
 sg13g2_fill_1 FILLER_32_56 ();
 sg13g2_fill_1 FILLER_32_70 ();
 sg13g2_fill_2 FILLER_32_88 ();
 sg13g2_fill_1 FILLER_32_100 ();
 sg13g2_fill_1 FILLER_32_111 ();
 sg13g2_decap_8 FILLER_32_117 ();
 sg13g2_fill_1 FILLER_32_124 ();
 sg13g2_decap_4 FILLER_32_139 ();
 sg13g2_fill_1 FILLER_32_143 ();
 sg13g2_fill_2 FILLER_32_155 ();
 sg13g2_fill_1 FILLER_32_157 ();
 sg13g2_decap_4 FILLER_32_168 ();
 sg13g2_fill_2 FILLER_32_172 ();
 sg13g2_fill_1 FILLER_32_190 ();
 sg13g2_fill_2 FILLER_32_214 ();
 sg13g2_fill_1 FILLER_32_216 ();
 sg13g2_fill_2 FILLER_32_222 ();
 sg13g2_fill_2 FILLER_32_234 ();
 sg13g2_decap_4 FILLER_32_242 ();
 sg13g2_decap_4 FILLER_32_251 ();
 sg13g2_fill_1 FILLER_32_255 ();
 sg13g2_decap_8 FILLER_32_269 ();
 sg13g2_fill_2 FILLER_32_276 ();
 sg13g2_fill_1 FILLER_32_278 ();
 sg13g2_fill_1 FILLER_32_293 ();
 sg13g2_fill_2 FILLER_32_298 ();
 sg13g2_fill_2 FILLER_32_310 ();
 sg13g2_decap_4 FILLER_32_343 ();
 sg13g2_fill_2 FILLER_32_367 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_4 ();
 sg13g2_fill_1 FILLER_33_16 ();
 sg13g2_fill_2 FILLER_33_70 ();
 sg13g2_fill_2 FILLER_33_96 ();
 sg13g2_fill_2 FILLER_33_103 ();
 sg13g2_fill_1 FILLER_33_105 ();
 sg13g2_fill_2 FILLER_33_126 ();
 sg13g2_fill_1 FILLER_33_138 ();
 sg13g2_fill_2 FILLER_33_151 ();
 sg13g2_fill_1 FILLER_33_153 ();
 sg13g2_decap_8 FILLER_33_165 ();
 sg13g2_decap_4 FILLER_33_184 ();
 sg13g2_fill_2 FILLER_33_188 ();
 sg13g2_decap_8 FILLER_33_195 ();
 sg13g2_fill_2 FILLER_33_202 ();
 sg13g2_fill_1 FILLER_33_217 ();
 sg13g2_decap_4 FILLER_33_248 ();
 sg13g2_fill_2 FILLER_33_262 ();
 sg13g2_decap_8 FILLER_33_281 ();
 sg13g2_fill_2 FILLER_33_306 ();
 sg13g2_decap_8 FILLER_33_336 ();
 sg13g2_fill_2 FILLER_33_343 ();
 sg13g2_fill_1 FILLER_33_345 ();
 sg13g2_fill_2 FILLER_33_354 ();
 sg13g2_fill_1 FILLER_33_356 ();
 sg13g2_fill_1 FILLER_33_364 ();
 sg13g2_fill_1 FILLER_33_377 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_2 ();
 sg13g2_fill_2 FILLER_34_25 ();
 sg13g2_fill_1 FILLER_34_27 ();
 sg13g2_fill_2 FILLER_34_34 ();
 sg13g2_fill_1 FILLER_34_36 ();
 sg13g2_fill_2 FILLER_34_51 ();
 sg13g2_fill_2 FILLER_34_116 ();
 sg13g2_fill_1 FILLER_34_122 ();
 sg13g2_fill_2 FILLER_34_128 ();
 sg13g2_fill_1 FILLER_34_135 ();
 sg13g2_fill_2 FILLER_34_145 ();
 sg13g2_fill_1 FILLER_34_187 ();
 sg13g2_fill_2 FILLER_34_203 ();
 sg13g2_fill_1 FILLER_34_205 ();
 sg13g2_decap_8 FILLER_34_223 ();
 sg13g2_fill_1 FILLER_34_236 ();
 sg13g2_fill_2 FILLER_34_265 ();
 sg13g2_fill_1 FILLER_34_286 ();
 sg13g2_fill_2 FILLER_34_291 ();
 sg13g2_fill_2 FILLER_34_297 ();
 sg13g2_fill_1 FILLER_34_299 ();
 sg13g2_decap_4 FILLER_34_309 ();
 sg13g2_fill_2 FILLER_34_313 ();
 sg13g2_fill_1 FILLER_34_391 ();
 sg13g2_fill_2 FILLER_34_397 ();
 sg13g2_fill_1 FILLER_34_399 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_15 ();
 sg13g2_fill_1 FILLER_35_17 ();
 sg13g2_fill_1 FILLER_35_27 ();
 sg13g2_fill_2 FILLER_35_37 ();
 sg13g2_fill_1 FILLER_35_39 ();
 sg13g2_fill_2 FILLER_35_50 ();
 sg13g2_fill_1 FILLER_35_52 ();
 sg13g2_fill_1 FILLER_35_58 ();
 sg13g2_fill_2 FILLER_35_65 ();
 sg13g2_fill_1 FILLER_35_67 ();
 sg13g2_fill_1 FILLER_35_81 ();
 sg13g2_fill_2 FILLER_35_88 ();
 sg13g2_fill_1 FILLER_35_96 ();
 sg13g2_fill_2 FILLER_35_113 ();
 sg13g2_decap_4 FILLER_35_130 ();
 sg13g2_fill_2 FILLER_35_147 ();
 sg13g2_fill_1 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_fill_2 FILLER_35_210 ();
 sg13g2_fill_2 FILLER_35_228 ();
 sg13g2_fill_2 FILLER_35_246 ();
 sg13g2_fill_2 FILLER_35_285 ();
 sg13g2_fill_1 FILLER_35_287 ();
 sg13g2_fill_1 FILLER_35_321 ();
 sg13g2_fill_2 FILLER_35_327 ();
 sg13g2_fill_2 FILLER_35_356 ();
 sg13g2_fill_2 FILLER_35_372 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_7 ();
 sg13g2_decap_4 FILLER_36_24 ();
 sg13g2_fill_2 FILLER_36_47 ();
 sg13g2_fill_2 FILLER_36_64 ();
 sg13g2_fill_1 FILLER_36_79 ();
 sg13g2_fill_2 FILLER_36_124 ();
 sg13g2_fill_1 FILLER_36_126 ();
 sg13g2_fill_2 FILLER_36_140 ();
 sg13g2_fill_1 FILLER_36_142 ();
 sg13g2_fill_2 FILLER_36_156 ();
 sg13g2_fill_2 FILLER_36_172 ();
 sg13g2_fill_1 FILLER_36_174 ();
 sg13g2_fill_2 FILLER_36_179 ();
 sg13g2_fill_1 FILLER_36_181 ();
 sg13g2_fill_2 FILLER_36_203 ();
 sg13g2_fill_1 FILLER_36_205 ();
 sg13g2_decap_4 FILLER_36_223 ();
 sg13g2_fill_1 FILLER_36_227 ();
 sg13g2_fill_1 FILLER_36_233 ();
 sg13g2_fill_2 FILLER_36_239 ();
 sg13g2_fill_1 FILLER_36_241 ();
 sg13g2_fill_1 FILLER_36_253 ();
 sg13g2_decap_4 FILLER_36_271 ();
 sg13g2_fill_1 FILLER_36_280 ();
 sg13g2_decap_4 FILLER_36_301 ();
 sg13g2_decap_4 FILLER_36_310 ();
 sg13g2_fill_2 FILLER_36_314 ();
 sg13g2_fill_2 FILLER_36_356 ();
 sg13g2_fill_1 FILLER_36_358 ();
 sg13g2_fill_2 FILLER_36_398 ();
 sg13g2_fill_1 FILLER_36_400 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_fill_2 FILLER_37_26 ();
 sg13g2_decap_4 FILLER_37_33 ();
 sg13g2_fill_1 FILLER_37_67 ();
 sg13g2_fill_1 FILLER_37_79 ();
 sg13g2_fill_2 FILLER_37_92 ();
 sg13g2_fill_1 FILLER_37_94 ();
 sg13g2_fill_1 FILLER_37_100 ();
 sg13g2_fill_1 FILLER_37_114 ();
 sg13g2_fill_2 FILLER_37_123 ();
 sg13g2_fill_1 FILLER_37_125 ();
 sg13g2_fill_2 FILLER_37_220 ();
 sg13g2_fill_1 FILLER_37_263 ();
 sg13g2_fill_1 FILLER_37_309 ();
 sg13g2_fill_1 FILLER_37_375 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_fill_2 FILLER_38_28 ();
 sg13g2_fill_1 FILLER_38_30 ();
 sg13g2_fill_1 FILLER_38_81 ();
 sg13g2_fill_2 FILLER_38_102 ();
 sg13g2_fill_1 FILLER_38_104 ();
 sg13g2_fill_2 FILLER_38_133 ();
 sg13g2_fill_1 FILLER_38_135 ();
 sg13g2_fill_2 FILLER_38_152 ();
 sg13g2_fill_2 FILLER_38_175 ();
 sg13g2_fill_2 FILLER_38_189 ();
 sg13g2_fill_1 FILLER_38_191 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_fill_2 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_218 ();
 sg13g2_fill_2 FILLER_38_225 ();
 sg13g2_fill_1 FILLER_38_247 ();
 sg13g2_decap_8 FILLER_38_256 ();
 sg13g2_decap_8 FILLER_38_263 ();
 sg13g2_decap_4 FILLER_38_270 ();
 sg13g2_fill_2 FILLER_38_278 ();
 sg13g2_fill_1 FILLER_38_280 ();
 sg13g2_fill_1 FILLER_38_291 ();
 sg13g2_decap_8 FILLER_38_303 ();
 sg13g2_fill_1 FILLER_38_310 ();
 sg13g2_fill_2 FILLER_38_353 ();
 sg13g2_fill_1 FILLER_38_393 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net6;
 assign uio_oe[1] = net7;
 assign uio_oe[2] = net8;
 assign uio_oe[3] = net9;
 assign uio_oe[4] = net10;
 assign uio_oe[5] = net11;
 assign uio_oe[6] = net12;
 assign uio_oe[7] = net13;
 assign uio_out[0] = net14;
 assign uio_out[1] = net15;
 assign uio_out[2] = net16;
 assign uio_out[3] = net17;
 assign uio_out[4] = net18;
 assign uio_out[5] = net19;
 assign uio_out[6] = net20;
 assign uio_out[7] = net21;
endmodule

module tt_um_iitbbs (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \C1.Program[0] ;
 wire \C1.Program[1] ;
 wire \C1.counter1[0] ;
 wire \C1.counter1[10] ;
 wire \C1.counter1[11] ;
 wire \C1.counter1[1] ;
 wire \C1.counter1[2] ;
 wire \C1.counter1[3] ;
 wire \C1.counter1[4] ;
 wire \C1.counter1[5] ;
 wire \C1.counter1[6] ;
 wire \C1.counter1[7] ;
 wire \C1.counter1[8] ;
 wire \C1.counter1[9] ;
 wire \C1.counter2[0] ;
 wire \C1.counter2[10] ;
 wire \C1.counter2[11] ;
 wire \C1.counter2[12] ;
 wire \C1.counter2[13] ;
 wire \C1.counter2[14] ;
 wire \C1.counter2[15] ;
 wire \C1.counter2[16] ;
 wire \C1.counter2[17] ;
 wire \C1.counter2[18] ;
 wire \C1.counter2[19] ;
 wire \C1.counter2[1] ;
 wire \C1.counter2[20] ;
 wire \C1.counter2[21] ;
 wire \C1.counter2[22] ;
 wire \C1.counter2[23] ;
 wire \C1.counter2[24] ;
 wire \C1.counter2[25] ;
 wire \C1.counter2[26] ;
 wire \C1.counter2[27] ;
 wire \C1.counter2[28] ;
 wire \C1.counter2[29] ;
 wire \C1.counter2[2] ;
 wire \C1.counter2[30] ;
 wire \C1.counter2[31] ;
 wire \C1.counter2[3] ;
 wire \C1.counter2[4] ;
 wire \C1.counter2[5] ;
 wire \C1.counter2[6] ;
 wire \C1.counter2[7] ;
 wire \C1.counter2[8] ;
 wire \C1.counter2[9] ;
 wire \C1.counter_status[0] ;
 wire \C1.counter_status[1] ;
 wire \C1.counter_status[2] ;
 wire \C1.dry_status ;
 wire \C1.dura_op ;
 wire \C1.heating ;
 wire \C1.level[0] ;
 wire \C1.level[1] ;
 wire \C1.level_op ;
 wire \C1.max_count[10] ;
 wire \C1.max_count[11] ;
 wire \C1.max_count[1] ;
 wire \C1.max_count[2] ;
 wire \C1.max_count[3] ;
 wire \C1.max_count[4] ;
 wire \C1.max_count[5] ;
 wire \C1.max_count[6] ;
 wire \C1.max_count[7] ;
 wire \C1.max_count[8] ;
 wire \C1.max_count[9] ;
 wire \C1.next_state_var[0] ;
 wire \C1.next_state_var[1] ;
 wire \C1.next_state_var[2] ;
 wire \C1.next_state_var[3] ;
 wire \C1.next_state_var[4] ;
 wire \C1.next_state_var[5] ;
 wire \C1.next_state_var[6] ;
 wire \C1.next_state_var[7] ;
 wire \C1.pouring ;
 wire \C1.prog_op ;
 wire \C1.rinse_status ;
 wire \C1.spinning ;
 wire \C1.temp[0] ;
 wire \C1.temp[1] ;
 wire \C1.temp_op ;
 wire \C1.timer[0] ;
 wire \C1.timer[1] ;
 wire \C1.waiting ;
 wire \FpgaPins_Fpga_FSM_data_a1[0] ;
 wire \FpgaPins_Fpga_FSM_data_a1[1] ;
 wire \FpgaPins_Fpga_FSM_data_a1[2] ;
 wire \FpgaPins_Fpga_FSM_data_a1[3] ;
 wire \FpgaPins_Fpga_FSM_data_a1[4] ;
 wire \FpgaPins_Fpga_FSM_data_a1[5] ;
 wire \FpgaPins_Fpga_FSM_data_a1[6] ;
 wire \FpgaPins_Fpga_FSM_data_a1[7] ;
 wire \FpgaPins_Fpga_FSM_idata_rd_addr_a1[0] ;
 wire \FpgaPins_Fpga_FSM_idata_rd_addr_a1[1] ;
 wire \FpgaPins_Fpga_FSM_idata_rd_addr_a1[2] ;
 wire \FpgaPins_Fpga_FSM_idata_rd_addr_a1[3] ;
 wire \FpgaPins_Fpga_FSM_imem_rd_addr_a1[0] ;
 wire \FpgaPins_Fpga_FSM_imem_rd_addr_a1[1] ;
 wire \FpgaPins_Fpga_FSM_imem_rd_addr_a1[2] ;
 wire \FpgaPins_Fpga_FSM_imem_rd_addr_a1[3] ;
 wire \FpgaPins_Fpga_FSM_imem_wr_addr_a1[0] ;
 wire \FpgaPins_Fpga_FSM_imem_wr_addr_a1[1] ;
 wire \FpgaPins_Fpga_FSM_imem_wr_addr_a1[2] ;
 wire \FpgaPins_Fpga_FSM_imem_wr_addr_a1[3] ;
 wire \FpgaPins_Fpga_FSM_instr_a1[0] ;
 wire \FpgaPins_Fpga_FSM_instr_a1[1] ;
 wire \FpgaPins_Fpga_FSM_instr_a1[2] ;
 wire \FpgaPins_Fpga_FSM_instr_a1[3] ;
 wire \FpgaPins_Fpga_FSM_instr_a1[4] ;
 wire \FpgaPins_Fpga_FSM_instr_a1[5] ;
 wire \FpgaPins_Fpga_FSM_instr_a1[6] ;
 wire \FpgaPins_Fpga_FSM_instr_a1[7] ;
 wire \FpgaPins_Fpga_FSM_instr_wr_a1[0] ;
 wire \FpgaPins_Fpga_FSM_instr_wr_a1[1] ;
 wire \FpgaPins_Fpga_FSM_instr_wr_a1[2] ;
 wire \FpgaPins_Fpga_FSM_instr_wr_a1[3] ;
 wire \FpgaPins_Fpga_FSM_instr_wr_a1[4] ;
 wire \FpgaPins_Fpga_FSM_instr_wr_a1[5] ;
 wire \FpgaPins_Fpga_FSM_instr_wr_a1[6] ;
 wire \FpgaPins_Fpga_FSM_instr_wr_a1[7] ;
 wire FpgaPins_Fpga_GAME_clk_pulse1_a1;
 wire FpgaPins_Fpga_GAME_clk_pulse1_a2;
 wire FpgaPins_Fpga_GAME_clk_pulse2_a1;
 wire FpgaPins_Fpga_GAME_clk_pulse2_a2;
 wire FpgaPins_Fpga_GAME_clk_pulse3_a1;
 wire FpgaPins_Fpga_GAME_clk_pulse3_a2;
 wire FpgaPins_Fpga_GAME_clk_pulse4_a1;
 wire FpgaPins_Fpga_GAME_clk_pulse4_a2;
 wire FpgaPins_Fpga_GAME_clk_pulse_a1;
 wire FpgaPins_Fpga_GAME_clk_pulse_a2;
 wire FpgaPins_Fpga_GAME_clk_pulse_a3;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[0] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[10] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[11] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[12] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[13] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[14] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[15] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[16] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[17] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[18] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[19] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[1] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[20] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[21] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[22] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[23] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[2] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[3] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[4] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[5] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[6] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[7] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[8] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a1[9] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[0] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[10] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[11] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[12] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[13] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[14] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[15] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[16] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[17] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[18] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[19] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[1] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[20] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[21] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[22] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[23] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[2] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[3] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[4] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[5] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[6] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[7] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[8] ;
 wire \FpgaPins_Fpga_GAME_count_speed1_a2[9] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[0] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[10] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[11] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[12] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[13] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[14] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[15] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[16] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[17] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[18] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[19] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[1] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[20] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[2] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[3] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[4] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[5] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[6] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[7] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[8] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a1[9] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[0] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[10] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[11] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[12] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[13] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[14] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[15] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[16] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[17] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[18] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[19] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[1] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[20] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[2] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[3] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[4] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[5] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[6] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[7] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[8] ;
 wire \FpgaPins_Fpga_GAME_count_speed2_a2[9] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a1[0] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a1[10] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a1[11] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a1[12] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a1[13] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a1[14] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a1[15] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a1[16] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a1[17] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a1[18] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a1[19] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a1[1] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a1[2] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a1[3] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a1[4] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a1[5] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a1[6] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a1[7] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a1[8] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a1[9] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a2[0] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a2[10] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a2[11] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a2[12] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a2[13] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a2[14] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a2[15] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a2[16] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a2[17] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a2[18] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a2[19] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a2[1] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a2[2] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a2[3] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a2[4] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a2[5] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a2[6] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a2[7] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a2[8] ;
 wire \FpgaPins_Fpga_GAME_count_speed3_a2[9] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a1[0] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a1[10] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a1[11] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a1[12] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a1[13] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a1[14] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a1[15] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a1[16] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a1[17] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a1[18] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a1[1] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a1[2] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a1[3] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a1[4] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a1[5] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a1[6] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a1[7] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a1[8] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a1[9] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a2[0] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a2[10] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a2[11] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a2[12] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a2[13] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a2[14] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a2[15] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a2[16] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a2[17] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a2[18] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a2[1] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a2[2] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a2[3] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a2[4] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a2[5] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a2[6] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a2[7] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a2[8] ;
 wire \FpgaPins_Fpga_GAME_count_speed4_a2[9] ;
 wire FpgaPins_Fpga_GAME_forward_a2;
 wire \FpgaPins_Fpga_GAME_led_output_a1[0] ;
 wire \FpgaPins_Fpga_GAME_led_output_a1[1] ;
 wire \FpgaPins_Fpga_GAME_led_output_a1[2] ;
 wire \FpgaPins_Fpga_GAME_led_output_a1[3] ;
 wire \FpgaPins_Fpga_GAME_led_output_a1[4] ;
 wire \FpgaPins_Fpga_GAME_led_output_a1[5] ;
 wire \FpgaPins_Fpga_GAME_led_output_a1[6] ;
 wire \FpgaPins_Fpga_GAME_led_output_a1[7] ;
 wire \FpgaPins_Fpga_GAME_led_output_a2[0] ;
 wire \FpgaPins_Fpga_GAME_led_output_a2[1] ;
 wire \FpgaPins_Fpga_GAME_led_output_a2[2] ;
 wire \FpgaPins_Fpga_GAME_led_output_a2[3] ;
 wire \FpgaPins_Fpga_GAME_led_output_a2[4] ;
 wire \FpgaPins_Fpga_GAME_led_output_a2[5] ;
 wire \FpgaPins_Fpga_GAME_led_output_a2[6] ;
 wire \FpgaPins_Fpga_GAME_led_output_a2[7] ;
 wire \FpgaPins_Fpga_GAME_led_output_a3[0] ;
 wire \FpgaPins_Fpga_GAME_led_output_a3[1] ;
 wire \FpgaPins_Fpga_GAME_led_output_a3[2] ;
 wire \FpgaPins_Fpga_GAME_led_output_a3[3] ;
 wire \FpgaPins_Fpga_GAME_led_output_a3[4] ;
 wire \FpgaPins_Fpga_GAME_led_output_a3[5] ;
 wire \FpgaPins_Fpga_GAME_led_output_a3[6] ;
 wire \FpgaPins_Fpga_GAME_led_output_a3[7] ;
 wire FpgaPins_Fpga_GAME_left_btn_a2;
 wire FpgaPins_Fpga_GAME_reset_a1;
 wire FpgaPins_Fpga_GAME_reset_a2;
 wire FpgaPins_Fpga_GAME_right_btn_a2;
 wire \FpgaPins_Fpga_GAME_score_a2[0] ;
 wire \FpgaPins_Fpga_GAME_score_a2[1] ;
 wire \FpgaPins_Fpga_GAME_score_a2[2] ;
 wire \FpgaPins_Fpga_GAME_score_a2[3] ;
 wire \FpgaPins_Fpga_GAME_score_a2[4] ;
 wire \FpgaPins_Fpga_GAME_score_a2[5] ;
 wire \FpgaPins_Fpga_GAME_score_a2[6] ;
 wire \FpgaPins_Fpga_GAME_score_a2[7] ;
 wire \FpgaPins_Fpga_GAME_score_a3[0] ;
 wire \FpgaPins_Fpga_GAME_score_a3[1] ;
 wire \FpgaPins_Fpga_GAME_score_a3[2] ;
 wire \FpgaPins_Fpga_GAME_score_a3[3] ;
 wire \FpgaPins_Fpga_GAME_score_a3[4] ;
 wire \FpgaPins_Fpga_GAME_score_a3[5] ;
 wire \FpgaPins_Fpga_GAME_score_a3[6] ;
 wire \FpgaPins_Fpga_GAME_score_a3[7] ;
 wire \FpgaPins_Fpga_GAME_score_a4[0] ;
 wire \FpgaPins_Fpga_GAME_score_a4[1] ;
 wire \FpgaPins_Fpga_GAME_score_a4[2] ;
 wire \FpgaPins_Fpga_GAME_score_a4[3] ;
 wire \FpgaPins_Fpga_GAME_score_a4[4] ;
 wire \FpgaPins_Fpga_GAME_score_a4[5] ;
 wire \FpgaPins_Fpga_GAME_score_a4[6] ;
 wire \FpgaPins_Fpga_GAME_score_a4[7] ;
 wire \FpgaPins_Fpga_GAME_speed_level_a2[1] ;
 wire \FpgaPins_Fpga_GAME_speed_level_a2[2] ;
 wire \FpgaPins_Fpga_GAME_speed_level_a2[3] ;
 wire \FpgaPins_Fpga_GAME_state_a2[0] ;
 wire \FpgaPins_Fpga_GAME_state_a2[1] ;
 wire \FpgaPins_Fpga_GAME_state_a3[0] ;
 wire \FpgaPins_Fpga_GAME_state_a3[1] ;
 wire \FpgaPins_Fpga_GAME_state_a4[0] ;
 wire \FpgaPins_Fpga_GAME_state_a4[1] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[0] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[10] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[11] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[12] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[13] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[14] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[15] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[16] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[17] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[18] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[19] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[1] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[20] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[21] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[22] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[23] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[24] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[2] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[3] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[4] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[5] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[6] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[7] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[8] ;
 wire \FpgaPins_Fpga_GAME_wait_counter_a2[9] ;
 wire \FpgaPins_Fpga_GAME_win_a1[0] ;
 wire \FpgaPins_Fpga_GAME_win_a1[1] ;
 wire \FpgaPins_Fpga_GAME_win_a2[1] ;
 wire \FpgaPins_Fpga_GAME_win_a2[2] ;
 wire \FpgaPins_Fpga_LIPSI_acc_a1[0] ;
 wire \FpgaPins_Fpga_LIPSI_acc_a1[1] ;
 wire \FpgaPins_Fpga_LIPSI_acc_a1[2] ;
 wire \FpgaPins_Fpga_LIPSI_acc_a1[3] ;
 wire \FpgaPins_Fpga_LIPSI_acc_a1[4] ;
 wire \FpgaPins_Fpga_LIPSI_acc_a1[5] ;
 wire \FpgaPins_Fpga_LIPSI_acc_a1[6] ;
 wire \FpgaPins_Fpga_LIPSI_acc_a1[7] ;
 wire \FpgaPins_Fpga_LIPSI_acc_a2[0] ;
 wire \FpgaPins_Fpga_LIPSI_acc_a2[1] ;
 wire \FpgaPins_Fpga_LIPSI_acc_a2[2] ;
 wire \FpgaPins_Fpga_LIPSI_acc_a2[3] ;
 wire \FpgaPins_Fpga_LIPSI_acc_a2[4] ;
 wire \FpgaPins_Fpga_LIPSI_acc_a2[5] ;
 wire \FpgaPins_Fpga_LIPSI_acc_a2[6] ;
 wire \FpgaPins_Fpga_LIPSI_acc_a2[7] ;
 wire FpgaPins_Fpga_LIPSI_c_a2;
 wire \FpgaPins_Fpga_LIPSI_data_a2[0] ;
 wire \FpgaPins_Fpga_LIPSI_data_a2[1] ;
 wire \FpgaPins_Fpga_LIPSI_data_a2[2] ;
 wire \FpgaPins_Fpga_LIPSI_data_a2[3] ;
 wire \FpgaPins_Fpga_LIPSI_data_a2[4] ;
 wire \FpgaPins_Fpga_LIPSI_data_a2[5] ;
 wire \FpgaPins_Fpga_LIPSI_data_a2[6] ;
 wire \FpgaPins_Fpga_LIPSI_data_a2[7] ;
 wire \FpgaPins_Fpga_LIPSI_data_wr_a1[0] ;
 wire \FpgaPins_Fpga_LIPSI_data_wr_a1[1] ;
 wire \FpgaPins_Fpga_LIPSI_data_wr_a1[2] ;
 wire \FpgaPins_Fpga_LIPSI_data_wr_a1[3] ;
 wire \FpgaPins_Fpga_LIPSI_data_wr_a1[4] ;
 wire \FpgaPins_Fpga_LIPSI_data_wr_a1[5] ;
 wire \FpgaPins_Fpga_LIPSI_data_wr_a1[6] ;
 wire \FpgaPins_Fpga_LIPSI_data_wr_a1[7] ;
 wire \FpgaPins_Fpga_LIPSI_data_wr_a2[0] ;
 wire \FpgaPins_Fpga_LIPSI_data_wr_a2[1] ;
 wire \FpgaPins_Fpga_LIPSI_data_wr_a2[2] ;
 wire \FpgaPins_Fpga_LIPSI_data_wr_a2[3] ;
 wire \FpgaPins_Fpga_LIPSI_data_wr_a2[4] ;
 wire \FpgaPins_Fpga_LIPSI_data_wr_a2[5] ;
 wire \FpgaPins_Fpga_LIPSI_data_wr_a2[6] ;
 wire \FpgaPins_Fpga_LIPSI_data_wr_a2[7] ;
 wire \FpgaPins_Fpga_LIPSI_dptr_a2[0] ;
 wire \FpgaPins_Fpga_LIPSI_dptr_a2[1] ;
 wire \FpgaPins_Fpga_LIPSI_dptr_a2[2] ;
 wire \FpgaPins_Fpga_LIPSI_dptr_a2[3] ;
 wire FpgaPins_Fpga_LIPSI_exit_a1;
 wire FpgaPins_Fpga_LIPSI_exit_a2;
 wire \FpgaPins_Fpga_LIPSI_instr_a2[0] ;
 wire \FpgaPins_Fpga_LIPSI_instr_a2[1] ;
 wire \FpgaPins_Fpga_LIPSI_instr_a2[2] ;
 wire \FpgaPins_Fpga_LIPSI_instr_a2[3] ;
 wire \FpgaPins_Fpga_LIPSI_instr_a2[4] ;
 wire \FpgaPins_Fpga_LIPSI_instr_a2[5] ;
 wire \FpgaPins_Fpga_LIPSI_instr_a2[6] ;
 wire \FpgaPins_Fpga_LIPSI_instr_a2[7] ;
 wire FpgaPins_Fpga_LIPSI_is_2cyc_a1;
 wire FpgaPins_Fpga_LIPSI_is_2cyc_a2;
 wire FpgaPins_Fpga_LIPSI_is_ALU_imm_a1;
 wire FpgaPins_Fpga_LIPSI_is_ALU_imm_a2;
 wire FpgaPins_Fpga_LIPSI_is_br_a1;
 wire FpgaPins_Fpga_LIPSI_is_br_a2;
 wire FpgaPins_Fpga_LIPSI_is_br_a3;
 wire FpgaPins_Fpga_LIPSI_is_brl_a1;
 wire FpgaPins_Fpga_LIPSI_is_brl_a2;
 wire FpgaPins_Fpga_LIPSI_is_brnz_a1;
 wire FpgaPins_Fpga_LIPSI_is_brnz_a2;
 wire FpgaPins_Fpga_LIPSI_is_brnz_a3;
 wire FpgaPins_Fpga_LIPSI_is_brz_a1;
 wire FpgaPins_Fpga_LIPSI_is_brz_a2;
 wire FpgaPins_Fpga_LIPSI_is_brz_a3;
 wire FpgaPins_Fpga_LIPSI_is_ld_ind_a1;
 wire FpgaPins_Fpga_LIPSI_is_ld_ind_a2;
 wire FpgaPins_Fpga_LIPSI_is_ret_a1;
 wire FpgaPins_Fpga_LIPSI_is_ret_a2;
 wire FpgaPins_Fpga_LIPSI_is_st_ind_a1;
 wire FpgaPins_Fpga_LIPSI_is_st_ind_a2;
 wire \FpgaPins_Fpga_LIPSI_pc_a1[4] ;
 wire \FpgaPins_Fpga_LIPSI_pc_a1[5] ;
 wire \FpgaPins_Fpga_LIPSI_pc_a1[6] ;
 wire \FpgaPins_Fpga_LIPSI_pc_a1[7] ;
 wire \FpgaPins_Fpga_LIPSI_pc_a2[0] ;
 wire \FpgaPins_Fpga_LIPSI_pc_a2[1] ;
 wire \FpgaPins_Fpga_LIPSI_pc_a2[2] ;
 wire \FpgaPins_Fpga_LIPSI_pc_a2[3] ;
 wire \FpgaPins_Fpga_LIPSI_pc_a2[4] ;
 wire \FpgaPins_Fpga_LIPSI_pc_a2[5] ;
 wire \FpgaPins_Fpga_LIPSI_pc_a2[6] ;
 wire \FpgaPins_Fpga_LIPSI_pc_a2[7] ;
 wire FpgaPins_Fpga_LIPSI_reset_a1;
 wire FpgaPins_Fpga_LIPSI_reset_a2;
 wire FpgaPins_Fpga_LIPSI_z_a1;
 wire FpgaPins_Fpga_LIPSI_z_a2;
 wire FpgaPins_Fpga_UART_comment_a1;
 wire FpgaPins_Fpga_UART_comment_a2;
 wire \FpgaPins_Fpga_UART_data_a2[0] ;
 wire \FpgaPins_Fpga_UART_data_a2[1] ;
 wire \FpgaPins_Fpga_UART_data_a2[2] ;
 wire \FpgaPins_Fpga_UART_data_a2[3] ;
 wire \FpgaPins_Fpga_UART_data_a2[4] ;
 wire \FpgaPins_Fpga_UART_data_a2[5] ;
 wire \FpgaPins_Fpga_UART_data_a2[6] ;
 wire \FpgaPins_Fpga_UART_data_a2[7] ;
 wire \FpgaPins_Fpga_UART_dptr_a2[0] ;
 wire \FpgaPins_Fpga_UART_dptr_a2[1] ;
 wire \FpgaPins_Fpga_UART_dptr_a2[2] ;
 wire \FpgaPins_Fpga_UART_dptr_a2[3] ;
 wire FpgaPins_Fpga_UART_first_byte_a2;
 wire FpgaPins_Fpga_UART_is_enter_a1;
 wire FpgaPins_Fpga_UART_is_enter_a2;
 wire \L1_Digit[0].L2_Leds[7].L2_viz_lit_a0 ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire clknet_leaf_0_clk;
 wire \datam[0][0] ;
 wire \datam[0][1] ;
 wire \datam[0][2] ;
 wire \datam[0][3] ;
 wire \datam[0][4] ;
 wire \datam[0][5] ;
 wire \datam[0][6] ;
 wire \datam[0][7] ;
 wire \datam[10][0] ;
 wire \datam[10][1] ;
 wire \datam[10][2] ;
 wire \datam[10][3] ;
 wire \datam[10][4] ;
 wire \datam[10][5] ;
 wire \datam[10][6] ;
 wire \datam[10][7] ;
 wire \datam[11][0] ;
 wire \datam[11][1] ;
 wire \datam[11][2] ;
 wire \datam[11][3] ;
 wire \datam[11][4] ;
 wire \datam[11][5] ;
 wire \datam[11][6] ;
 wire \datam[11][7] ;
 wire \datam[12][0] ;
 wire \datam[12][1] ;
 wire \datam[12][2] ;
 wire \datam[12][3] ;
 wire \datam[12][4] ;
 wire \datam[12][5] ;
 wire \datam[12][6] ;
 wire \datam[12][7] ;
 wire \datam[13][0] ;
 wire \datam[13][1] ;
 wire \datam[13][2] ;
 wire \datam[13][3] ;
 wire \datam[13][4] ;
 wire \datam[13][5] ;
 wire \datam[13][6] ;
 wire \datam[13][7] ;
 wire \datam[14][0] ;
 wire \datam[14][1] ;
 wire \datam[14][2] ;
 wire \datam[14][3] ;
 wire \datam[14][4] ;
 wire \datam[14][5] ;
 wire \datam[14][6] ;
 wire \datam[14][7] ;
 wire \datam[15][0] ;
 wire \datam[15][1] ;
 wire \datam[15][2] ;
 wire \datam[15][3] ;
 wire \datam[15][4] ;
 wire \datam[15][5] ;
 wire \datam[15][6] ;
 wire \datam[15][7] ;
 wire \datam[1][0] ;
 wire \datam[1][1] ;
 wire \datam[1][2] ;
 wire \datam[1][3] ;
 wire \datam[1][4] ;
 wire \datam[1][5] ;
 wire \datam[1][6] ;
 wire \datam[1][7] ;
 wire \datam[2][0] ;
 wire \datam[2][1] ;
 wire \datam[2][2] ;
 wire \datam[2][3] ;
 wire \datam[2][4] ;
 wire \datam[2][5] ;
 wire \datam[2][6] ;
 wire \datam[2][7] ;
 wire \datam[3][0] ;
 wire \datam[3][1] ;
 wire \datam[3][2] ;
 wire \datam[3][3] ;
 wire \datam[3][4] ;
 wire \datam[3][5] ;
 wire \datam[3][6] ;
 wire \datam[3][7] ;
 wire \datam[4][0] ;
 wire \datam[4][1] ;
 wire \datam[4][2] ;
 wire \datam[4][3] ;
 wire \datam[4][4] ;
 wire \datam[4][5] ;
 wire \datam[4][6] ;
 wire \datam[4][7] ;
 wire \datam[5][0] ;
 wire \datam[5][1] ;
 wire \datam[5][2] ;
 wire \datam[5][3] ;
 wire \datam[5][4] ;
 wire \datam[5][5] ;
 wire \datam[5][6] ;
 wire \datam[5][7] ;
 wire \datam[6][0] ;
 wire \datam[6][1] ;
 wire \datam[6][2] ;
 wire \datam[6][3] ;
 wire \datam[6][4] ;
 wire \datam[6][5] ;
 wire \datam[6][6] ;
 wire \datam[6][7] ;
 wire \datam[7][0] ;
 wire \datam[7][1] ;
 wire \datam[7][2] ;
 wire \datam[7][3] ;
 wire \datam[7][4] ;
 wire \datam[7][5] ;
 wire \datam[7][6] ;
 wire \datam[7][7] ;
 wire \datam[8][0] ;
 wire \datam[8][1] ;
 wire \datam[8][2] ;
 wire \datam[8][3] ;
 wire \datam[8][4] ;
 wire \datam[8][5] ;
 wire \datam[8][6] ;
 wire \datam[8][7] ;
 wire \datam[9][0] ;
 wire \datam[9][1] ;
 wire \datam[9][2] ;
 wire \datam[9][3] ;
 wire \datam[9][4] ;
 wire \datam[9][5] ;
 wire \datam[9][6] ;
 wire \datam[9][7] ;
 wire \instrs[0][0] ;
 wire \instrs[0][1] ;
 wire \instrs[0][2] ;
 wire \instrs[0][3] ;
 wire \instrs[0][4] ;
 wire \instrs[0][5] ;
 wire \instrs[0][6] ;
 wire \instrs[0][7] ;
 wire \instrs[10][0] ;
 wire \instrs[10][1] ;
 wire \instrs[10][2] ;
 wire \instrs[10][3] ;
 wire \instrs[10][4] ;
 wire \instrs[10][5] ;
 wire \instrs[10][6] ;
 wire \instrs[10][7] ;
 wire \instrs[11][0] ;
 wire \instrs[11][1] ;
 wire \instrs[11][2] ;
 wire \instrs[11][3] ;
 wire \instrs[11][4] ;
 wire \instrs[11][5] ;
 wire \instrs[11][6] ;
 wire \instrs[11][7] ;
 wire \instrs[12][0] ;
 wire \instrs[12][1] ;
 wire \instrs[12][2] ;
 wire \instrs[12][3] ;
 wire \instrs[12][4] ;
 wire \instrs[12][5] ;
 wire \instrs[12][6] ;
 wire \instrs[12][7] ;
 wire \instrs[13][0] ;
 wire \instrs[13][1] ;
 wire \instrs[13][2] ;
 wire \instrs[13][3] ;
 wire \instrs[13][4] ;
 wire \instrs[13][5] ;
 wire \instrs[13][6] ;
 wire \instrs[13][7] ;
 wire \instrs[14][0] ;
 wire \instrs[14][1] ;
 wire \instrs[14][2] ;
 wire \instrs[14][3] ;
 wire \instrs[14][4] ;
 wire \instrs[14][5] ;
 wire \instrs[14][6] ;
 wire \instrs[14][7] ;
 wire \instrs[15][0] ;
 wire \instrs[15][1] ;
 wire \instrs[15][2] ;
 wire \instrs[15][3] ;
 wire \instrs[15][4] ;
 wire \instrs[15][5] ;
 wire \instrs[15][6] ;
 wire \instrs[15][7] ;
 wire \instrs[1][0] ;
 wire \instrs[1][1] ;
 wire \instrs[1][2] ;
 wire \instrs[1][3] ;
 wire \instrs[1][4] ;
 wire \instrs[1][5] ;
 wire \instrs[1][6] ;
 wire \instrs[1][7] ;
 wire \instrs[2][0] ;
 wire \instrs[2][1] ;
 wire \instrs[2][2] ;
 wire \instrs[2][3] ;
 wire \instrs[2][4] ;
 wire \instrs[2][5] ;
 wire \instrs[2][6] ;
 wire \instrs[2][7] ;
 wire \instrs[3][0] ;
 wire \instrs[3][1] ;
 wire \instrs[3][2] ;
 wire \instrs[3][3] ;
 wire \instrs[3][4] ;
 wire \instrs[3][5] ;
 wire \instrs[3][6] ;
 wire \instrs[3][7] ;
 wire \instrs[4][0] ;
 wire \instrs[4][1] ;
 wire \instrs[4][2] ;
 wire \instrs[4][3] ;
 wire \instrs[4][4] ;
 wire \instrs[4][5] ;
 wire \instrs[4][6] ;
 wire \instrs[4][7] ;
 wire \instrs[5][0] ;
 wire \instrs[5][1] ;
 wire \instrs[5][2] ;
 wire \instrs[5][3] ;
 wire \instrs[5][4] ;
 wire \instrs[5][5] ;
 wire \instrs[5][6] ;
 wire \instrs[5][7] ;
 wire \instrs[6][0] ;
 wire \instrs[6][1] ;
 wire \instrs[6][2] ;
 wire \instrs[6][3] ;
 wire \instrs[6][4] ;
 wire \instrs[6][5] ;
 wire \instrs[6][6] ;
 wire \instrs[6][7] ;
 wire \instrs[7][0] ;
 wire \instrs[7][1] ;
 wire \instrs[7][2] ;
 wire \instrs[7][3] ;
 wire \instrs[7][4] ;
 wire \instrs[7][5] ;
 wire \instrs[7][6] ;
 wire \instrs[7][7] ;
 wire \instrs[8][0] ;
 wire \instrs[8][1] ;
 wire \instrs[8][2] ;
 wire \instrs[8][3] ;
 wire \instrs[8][4] ;
 wire \instrs[8][5] ;
 wire \instrs[8][6] ;
 wire \instrs[8][7] ;
 wire \instrs[9][0] ;
 wire \instrs[9][1] ;
 wire \instrs[9][2] ;
 wire \instrs[9][3] ;
 wire \instrs[9][4] ;
 wire \instrs[9][5] ;
 wire \instrs[9][6] ;
 wire \instrs[9][7] ;
 wire \uart_rx_1.r_Bit_Index[0] ;
 wire \uart_rx_1.r_Bit_Index[10] ;
 wire \uart_rx_1.r_Bit_Index[11] ;
 wire \uart_rx_1.r_Bit_Index[12] ;
 wire \uart_rx_1.r_Bit_Index[13] ;
 wire \uart_rx_1.r_Bit_Index[14] ;
 wire \uart_rx_1.r_Bit_Index[15] ;
 wire \uart_rx_1.r_Bit_Index[16] ;
 wire \uart_rx_1.r_Bit_Index[17] ;
 wire \uart_rx_1.r_Bit_Index[18] ;
 wire \uart_rx_1.r_Bit_Index[19] ;
 wire \uart_rx_1.r_Bit_Index[1] ;
 wire \uart_rx_1.r_Bit_Index[20] ;
 wire \uart_rx_1.r_Bit_Index[21] ;
 wire \uart_rx_1.r_Bit_Index[22] ;
 wire \uart_rx_1.r_Bit_Index[23] ;
 wire \uart_rx_1.r_Bit_Index[24] ;
 wire \uart_rx_1.r_Bit_Index[25] ;
 wire \uart_rx_1.r_Bit_Index[26] ;
 wire \uart_rx_1.r_Bit_Index[27] ;
 wire \uart_rx_1.r_Bit_Index[28] ;
 wire \uart_rx_1.r_Bit_Index[29] ;
 wire \uart_rx_1.r_Bit_Index[2] ;
 wire \uart_rx_1.r_Bit_Index[30] ;
 wire \uart_rx_1.r_Bit_Index[31] ;
 wire \uart_rx_1.r_Bit_Index[3] ;
 wire \uart_rx_1.r_Bit_Index[4] ;
 wire \uart_rx_1.r_Bit_Index[5] ;
 wire \uart_rx_1.r_Bit_Index[6] ;
 wire \uart_rx_1.r_Bit_Index[7] ;
 wire \uart_rx_1.r_Bit_Index[8] ;
 wire \uart_rx_1.r_Bit_Index[9] ;
 wire \uart_rx_1.r_Clock_Count[0] ;
 wire \uart_rx_1.r_Clock_Count[10] ;
 wire \uart_rx_1.r_Clock_Count[11] ;
 wire \uart_rx_1.r_Clock_Count[12] ;
 wire \uart_rx_1.r_Clock_Count[13] ;
 wire \uart_rx_1.r_Clock_Count[14] ;
 wire \uart_rx_1.r_Clock_Count[15] ;
 wire \uart_rx_1.r_Clock_Count[16] ;
 wire \uart_rx_1.r_Clock_Count[17] ;
 wire \uart_rx_1.r_Clock_Count[18] ;
 wire \uart_rx_1.r_Clock_Count[19] ;
 wire \uart_rx_1.r_Clock_Count[1] ;
 wire \uart_rx_1.r_Clock_Count[20] ;
 wire \uart_rx_1.r_Clock_Count[21] ;
 wire \uart_rx_1.r_Clock_Count[22] ;
 wire \uart_rx_1.r_Clock_Count[23] ;
 wire \uart_rx_1.r_Clock_Count[24] ;
 wire \uart_rx_1.r_Clock_Count[25] ;
 wire \uart_rx_1.r_Clock_Count[26] ;
 wire \uart_rx_1.r_Clock_Count[27] ;
 wire \uart_rx_1.r_Clock_Count[28] ;
 wire \uart_rx_1.r_Clock_Count[29] ;
 wire \uart_rx_1.r_Clock_Count[2] ;
 wire \uart_rx_1.r_Clock_Count[30] ;
 wire \uart_rx_1.r_Clock_Count[31] ;
 wire \uart_rx_1.r_Clock_Count[3] ;
 wire \uart_rx_1.r_Clock_Count[4] ;
 wire \uart_rx_1.r_Clock_Count[5] ;
 wire \uart_rx_1.r_Clock_Count[6] ;
 wire \uart_rx_1.r_Clock_Count[7] ;
 wire \uart_rx_1.r_Clock_Count[8] ;
 wire \uart_rx_1.r_Clock_Count[9] ;
 wire \uart_rx_1.r_Rx_Byte[0] ;
 wire \uart_rx_1.r_Rx_Byte[1] ;
 wire \uart_rx_1.r_Rx_Byte[2] ;
 wire \uart_rx_1.r_Rx_Byte[3] ;
 wire \uart_rx_1.r_Rx_Byte[4] ;
 wire \uart_rx_1.r_Rx_Byte[5] ;
 wire \uart_rx_1.r_Rx_Byte[6] ;
 wire \uart_rx_1.r_Rx_Byte[7] ;
 wire \uart_rx_1.r_Rx_DV ;
 wire \uart_rx_1.r_Rx_Data ;
 wire \uart_rx_1.r_Rx_Data_R ;
 wire \uart_rx_1.r_SM_Main[0] ;
 wire \uart_rx_1.r_SM_Main[1] ;
 wire \uart_rx_1.r_SM_Main[2] ;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;

 sg13g2_inv_1 _4042_ (.Y(_0660_),
    .A(\uart_rx_1.r_Clock_Count[7] ));
 sg13g2_inv_1 _4043_ (.Y(_0661_),
    .A(net1519));
 sg13g2_inv_1 _4044_ (.Y(_0662_),
    .A(net1400));
 sg13g2_inv_1 _4045_ (.Y(_0663_),
    .A(net1262));
 sg13g2_inv_1 _4046_ (.Y(_0664_),
    .A(\uart_rx_1.r_Bit_Index[1] ));
 sg13g2_inv_1 _4047_ (.Y(_0665_),
    .A(net1515));
 sg13g2_inv_1 _4048_ (.Y(_0666_),
    .A(\uart_rx_1.r_Rx_Byte[3] ));
 sg13g2_inv_1 _4049_ (.Y(_0667_),
    .A(\uart_rx_1.r_Rx_Byte[2] ));
 sg13g2_inv_1 _4050_ (.Y(_0668_),
    .A(net1659));
 sg13g2_inv_2 _4051_ (.Y(_0669_),
    .A(net1744));
 sg13g2_inv_4 _4052_ (.A(net1750),
    .Y(_0670_));
 sg13g2_inv_1 _4053_ (.Y(_0671_),
    .A(net1742));
 sg13g2_inv_2 _4054_ (.Y(_0672_),
    .A(net1741));
 sg13g2_inv_1 _4055_ (.Y(_0673_),
    .A(net1359));
 sg13g2_inv_1 _4056_ (.Y(_0674_),
    .A(net1424));
 sg13g2_inv_1 _4057_ (.Y(_0675_),
    .A(net1654));
 sg13g2_inv_2 _4058_ (.Y(_0676_),
    .A(net1736));
 sg13g2_inv_1 _4059_ (.Y(_0677_),
    .A(net1014));
 sg13g2_inv_1 _4060_ (.Y(_0678_),
    .A(net1123));
 sg13g2_inv_1 _4061_ (.Y(_0679_),
    .A(net1109));
 sg13g2_inv_1 _4062_ (.Y(_0680_),
    .A(net1235));
 sg13g2_inv_1 _4063_ (.Y(_0681_),
    .A(\FpgaPins_Fpga_GAME_score_a2[3] ));
 sg13g2_inv_1 _4064_ (.Y(_0682_),
    .A(net713));
 sg13g2_inv_1 _4065_ (.Y(_0683_),
    .A(net712));
 sg13g2_inv_1 _4066_ (.Y(_0684_),
    .A(net704));
 sg13g2_inv_1 _4067_ (.Y(_0685_),
    .A(net726));
 sg13g2_inv_2 _4068_ (.Y(_0686_),
    .A(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[3] ));
 sg13g2_inv_1 _4069_ (.Y(_0687_),
    .A(net991));
 sg13g2_inv_1 _4070_ (.Y(_0688_),
    .A(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[0] ));
 sg13g2_inv_1 _4071_ (.Y(_0689_),
    .A(\C1.max_count[9] ));
 sg13g2_inv_1 _4072_ (.Y(_0690_),
    .A(\C1.max_count[3] ));
 sg13g2_inv_1 _4073_ (.Y(_0691_),
    .A(\FpgaPins_Fpga_GAME_count_speed1_a2[6] ));
 sg13g2_inv_1 _4074_ (.Y(_0692_),
    .A(\FpgaPins_Fpga_GAME_count_speed1_a2[10] ));
 sg13g2_inv_2 _4075_ (.Y(_0693_),
    .A(net1492));
 sg13g2_inv_1 _4076_ (.Y(_0694_),
    .A(\FpgaPins_Fpga_GAME_score_a4[7] ));
 sg13g2_inv_1 _4077_ (.Y(_0695_),
    .A(net1527));
 sg13g2_inv_1 _4078_ (.Y(_0696_),
    .A(\FpgaPins_Fpga_GAME_win_a2[1] ));
 sg13g2_inv_1 _4079_ (.Y(_0697_),
    .A(_0022_));
 sg13g2_inv_1 _4080_ (.Y(_0698_),
    .A(net987));
 sg13g2_inv_2 _4081_ (.Y(_0699_),
    .A(net988));
 sg13g2_inv_1 _4082_ (.Y(_0700_),
    .A(FpgaPins_Fpga_LIPSI_reset_a2));
 sg13g2_inv_1 _4083_ (.Y(_0701_),
    .A(\FpgaPins_Fpga_LIPSI_acc_a2[1] ));
 sg13g2_inv_1 _4084_ (.Y(_0702_),
    .A(_0024_));
 sg13g2_inv_2 _4085_ (.Y(_0703_),
    .A(_0028_));
 sg13g2_inv_1 _4086_ (.Y(_0704_),
    .A(_0031_));
 sg13g2_inv_1 _4087_ (.Y(_0705_),
    .A(\FpgaPins_Fpga_GAME_count_speed4_a2[13] ));
 sg13g2_inv_1 _4088_ (.Y(_0706_),
    .A(\FpgaPins_Fpga_GAME_count_speed4_a2[8] ));
 sg13g2_inv_1 _4089_ (.Y(_0707_),
    .A(\FpgaPins_Fpga_GAME_count_speed3_a2[10] ));
 sg13g2_inv_1 _4090_ (.Y(_0708_),
    .A(net1710));
 sg13g2_inv_1 _4091_ (.Y(_0709_),
    .A(net992));
 sg13g2_inv_2 _4092_ (.Y(_0710_),
    .A(net995));
 sg13g2_inv_1 _4093_ (.Y(_0711_),
    .A(\C1.spinning ));
 sg13g2_inv_1 _4094_ (.Y(_0712_),
    .A(\C1.counter1[2] ));
 sg13g2_inv_1 _4095_ (.Y(_0713_),
    .A(net1745));
 sg13g2_inv_1 _4096_ (.Y(_0714_),
    .A(\C1.counter1[6] ));
 sg13g2_inv_1 _4097_ (.Y(_0715_),
    .A(net1751));
 sg13g2_inv_1 _4098_ (.Y(_0716_),
    .A(\C1.counter2[6] ));
 sg13g2_inv_1 _4099_ (.Y(_0717_),
    .A(net753));
 sg13g2_inv_1 _4100_ (.Y(_0718_),
    .A(\FpgaPins_Fpga_GAME_led_output_a2[2] ));
 sg13g2_inv_1 _4101_ (.Y(_0719_),
    .A(\FpgaPins_Fpga_GAME_score_a4[6] ));
 sg13g2_inv_1 _4102_ (.Y(_0720_),
    .A(\FpgaPins_Fpga_GAME_led_output_a2[4] ));
 sg13g2_inv_1 _4103_ (.Y(_0721_),
    .A(\FpgaPins_Fpga_GAME_led_output_a2[3] ));
 sg13g2_inv_1 _4104_ (.Y(_0722_),
    .A(net999));
 sg13g2_inv_1 _4105_ (.Y(_0723_),
    .A(net3));
 sg13g2_inv_1 _4106_ (.Y(_0724_),
    .A(net1546));
 sg13g2_inv_1 _4107_ (.Y(_0725_),
    .A(net1495));
 sg13g2_inv_1 _4108_ (.Y(_0726_),
    .A(\FpgaPins_Fpga_GAME_wait_counter_a2[19] ));
 sg13g2_inv_1 _4109_ (.Y(_0727_),
    .A(_0099_));
 sg13g2_inv_1 _4110_ (.Y(_0728_),
    .A(FpgaPins_Fpga_LIPSI_is_ALU_imm_a2));
 sg13g2_inv_1 _4111_ (.Y(_0729_),
    .A(_0110_));
 sg13g2_inv_1 _4112_ (.Y(_0730_),
    .A(_0119_));
 sg13g2_inv_1 _4113_ (.Y(_0731_),
    .A(\FpgaPins_Fpga_LIPSI_acc_a2[7] ));
 sg13g2_inv_1 _4114_ (.Y(_0732_),
    .A(_0128_));
 sg13g2_inv_1 _4115_ (.Y(_0733_),
    .A(_0137_));
 sg13g2_inv_1 _4116_ (.Y(_0734_),
    .A(_0144_));
 sg13g2_inv_1 _4117_ (.Y(_0735_),
    .A(_0148_));
 sg13g2_inv_1 _4118_ (.Y(_0736_),
    .A(_0152_));
 sg13g2_inv_1 _4119_ (.Y(_0737_),
    .A(_0160_));
 sg13g2_inv_1 _4120_ (.Y(_0738_),
    .A(_0169_));
 sg13g2_inv_1 _4121_ (.Y(_0739_),
    .A(_0172_));
 sg13g2_inv_1 _4122_ (.Y(_0740_),
    .A(_0177_));
 sg13g2_inv_1 _4123_ (.Y(_0741_),
    .A(_0186_));
 sg13g2_inv_1 _4124_ (.Y(_0742_),
    .A(\FpgaPins_Fpga_LIPSI_acc_a2[5] ));
 sg13g2_inv_1 _4125_ (.Y(_0743_),
    .A(_0189_));
 sg13g2_inv_1 _4126_ (.Y(_0744_),
    .A(net1283));
 sg13g2_inv_1 _4127_ (.Y(_0745_),
    .A(net1099));
 sg13g2_inv_2 _4128_ (.Y(_0746_),
    .A(_0190_));
 sg13g2_inv_1 _4129_ (.Y(_0747_),
    .A(\datam[4][6] ));
 sg13g2_inv_1 _4130_ (.Y(_0748_),
    .A(\datam[8][6] ));
 sg13g2_inv_1 _4131_ (.Y(_0749_),
    .A(\datam[12][6] ));
 sg13g2_inv_1 _4132_ (.Y(_0750_),
    .A(\datam[4][7] ));
 sg13g2_inv_1 _4133_ (.Y(_0751_),
    .A(\datam[13][7] ));
 sg13g2_inv_1 _4134_ (.Y(_0752_),
    .A(_0191_));
 sg13g2_inv_1 _4135_ (.Y(_0753_),
    .A(\FpgaPins_Fpga_UART_data_a2[4] ));
 sg13g2_inv_1 _4136_ (.Y(_0754_),
    .A(_0197_));
 sg13g2_inv_1 _4137_ (.Y(_0755_),
    .A(_0199_));
 sg13g2_inv_1 _4138_ (.Y(_0756_),
    .A(\FpgaPins_Fpga_UART_data_a2[6] ));
 sg13g2_inv_1 _4139_ (.Y(_0757_),
    .A(_0201_));
 sg13g2_inv_1 _4140_ (.Y(_0758_),
    .A(net1478));
 sg13g2_and2_1 _4141_ (.A(net1616),
    .B(net725),
    .X(_0759_));
 sg13g2_and2_1 _4142_ (.A(net1432),
    .B(_0759_),
    .X(_0760_));
 sg13g2_and2_1 _4143_ (.A(net1446),
    .B(_0760_),
    .X(_0761_));
 sg13g2_and2_1 _4144_ (.A(net1450),
    .B(_0761_),
    .X(_0762_));
 sg13g2_and2_1 _4145_ (.A(net1494),
    .B(_0762_),
    .X(_0763_));
 sg13g2_and2_1 _4146_ (.A(net1393),
    .B(_0763_),
    .X(_0764_));
 sg13g2_and2_1 _4147_ (.A(net1721),
    .B(_0764_),
    .X(_0765_));
 sg13g2_and2_1 _4148_ (.A(net1579),
    .B(_0765_),
    .X(_0766_));
 sg13g2_and2_1 _4149_ (.A(net1556),
    .B(_0766_),
    .X(_0767_));
 sg13g2_and2_1 _4150_ (.A(net1615),
    .B(_0767_),
    .X(_0768_));
 sg13g2_nor4_1 _4151_ (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[5] ),
    .B(\FpgaPins_Fpga_GAME_count_speed1_a2[4] ),
    .C(\FpgaPins_Fpga_GAME_count_speed1_a2[3] ),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a2[2] ),
    .Y(_0769_));
 sg13g2_nor2_1 _4152_ (.A(net1616),
    .B(net725),
    .Y(_0770_));
 sg13g2_nand4_1 _4153_ (.B(_0691_),
    .C(_0769_),
    .A(\FpgaPins_Fpga_GAME_count_speed1_a2[7] ),
    .Y(_0771_),
    .D(_0770_));
 sg13g2_nor3_1 _4154_ (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[13] ),
    .B(\FpgaPins_Fpga_GAME_count_speed1_a2[12] ),
    .C(\FpgaPins_Fpga_GAME_count_speed1_a2[14] ),
    .Y(_0772_));
 sg13g2_nor4_1 _4155_ (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[9] ),
    .B(\FpgaPins_Fpga_GAME_count_speed1_a2[8] ),
    .C(_0692_),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a2[11] ),
    .Y(_0773_));
 sg13g2_nand3_1 _4156_ (.B(_0772_),
    .C(_0773_),
    .A(\FpgaPins_Fpga_GAME_count_speed1_a2[15] ),
    .Y(_0774_));
 sg13g2_nor2b_1 _4157_ (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[16] ),
    .B_N(\FpgaPins_Fpga_GAME_count_speed1_a2[17] ),
    .Y(_0775_));
 sg13g2_nand2b_1 _4158_ (.Y(_0776_),
    .B(\FpgaPins_Fpga_GAME_count_speed1_a2[20] ),
    .A_N(\FpgaPins_Fpga_GAME_count_speed1_a2[21] ));
 sg13g2_nor4_1 _4159_ (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[23] ),
    .B(\FpgaPins_Fpga_GAME_count_speed1_a2[22] ),
    .C(_0774_),
    .D(_0776_),
    .Y(_0777_));
 sg13g2_nand4_1 _4160_ (.B(\FpgaPins_Fpga_GAME_count_speed1_a2[18] ),
    .C(_0775_),
    .A(\FpgaPins_Fpga_GAME_count_speed1_a2[19] ),
    .Y(_0778_),
    .D(_0777_));
 sg13g2_o21ai_1 _4161_ (.B1(net985),
    .Y(_0779_),
    .A1(_0771_),
    .A2(_0778_));
 sg13g2_inv_1 _4162_ (.Y(_0780_),
    .A(net898));
 sg13g2_o21ai_1 _4163_ (.B1(net892),
    .Y(_0781_),
    .A1(net1615),
    .A2(_0767_));
 sg13g2_nor2_1 _4164_ (.A(_0768_),
    .B(_0781_),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[10] ));
 sg13g2_o21ai_1 _4165_ (.B1(net1687),
    .Y(_0782_),
    .A1(_0695_),
    .A2(_0696_));
 sg13g2_nor2b_2 _4166_ (.A(FpgaPins_Fpga_GAME_clk_pulse_a3),
    .B_N(FpgaPins_Fpga_GAME_clk_pulse_a2),
    .Y(_0783_));
 sg13g2_nand2b_1 _4167_ (.Y(_0784_),
    .B(FpgaPins_Fpga_GAME_clk_pulse_a2),
    .A_N(FpgaPins_Fpga_GAME_clk_pulse_a3));
 sg13g2_nor2b_1 _4168_ (.A(\FpgaPins_Fpga_GAME_state_a3[0] ),
    .B_N(\FpgaPins_Fpga_GAME_state_a3[1] ),
    .Y(_0785_));
 sg13g2_nand2b_1 _4169_ (.Y(_0786_),
    .B(\FpgaPins_Fpga_GAME_state_a3[1] ),
    .A_N(\FpgaPins_Fpga_GAME_state_a3[0] ));
 sg13g2_nand3_1 _4170_ (.B(\FpgaPins_Fpga_GAME_led_output_a2[6] ),
    .C(_0783_),
    .A(net984),
    .Y(_0787_));
 sg13g2_a21oi_1 _4171_ (.A1(\FpgaPins_Fpga_GAME_led_output_a2[7] ),
    .A2(_0784_),
    .Y(_0788_),
    .B1(net979));
 sg13g2_nor2_1 _4172_ (.A(\FpgaPins_Fpga_GAME_state_a3[1] ),
    .B(\FpgaPins_Fpga_GAME_state_a4[0] ),
    .Y(_0789_));
 sg13g2_nand3_1 _4173_ (.B(\FpgaPins_Fpga_GAME_state_a4[1] ),
    .C(_0789_),
    .A(\FpgaPins_Fpga_GAME_state_a3[0] ),
    .Y(_0790_));
 sg13g2_nand2_2 _4174_ (.Y(_0791_),
    .A(net985),
    .B(_0790_));
 sg13g2_a221oi_1 _4175_ (.B2(_0788_),
    .C1(_0791_),
    .B1(_0787_),
    .A1(_0694_),
    .Y(_0792_),
    .A2(net979));
 sg13g2_nor2_1 _4176_ (.A(net1636),
    .B(_0792_),
    .Y(_0793_));
 sg13g2_nor2_1 _4177_ (.A(_0782_),
    .B(_0793_),
    .Y(\FpgaPins_Fpga_GAME_led_output_a1[7] ));
 sg13g2_o21ai_1 _4178_ (.B1(net892),
    .Y(_0794_),
    .A1(net1721),
    .A2(_0764_));
 sg13g2_nor2_1 _4179_ (.A(_0765_),
    .B(_0794_),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[7] ));
 sg13g2_nor2b_2 _4180_ (.A(net8),
    .B_N(net1),
    .Y(_0795_));
 sg13g2_nor2b_1 _4181_ (.A(net2),
    .B_N(_0795_),
    .Y(_0796_));
 sg13g2_inv_1 _4182_ (.Y(FpgaPins_Fpga_LIPSI_reset_a1),
    .A(net975));
 sg13g2_nor2_2 _4183_ (.A(net989),
    .B(FpgaPins_Fpga_LIPSI_is_st_ind_a2),
    .Y(_0797_));
 sg13g2_nor3_1 _4184_ (.A(FpgaPins_Fpga_LIPSI_exit_a2),
    .B(net989),
    .C(FpgaPins_Fpga_LIPSI_is_st_ind_a2),
    .Y(_0798_));
 sg13g2_nand2b_1 _4185_ (.Y(_0799_),
    .B(_0797_),
    .A_N(FpgaPins_Fpga_LIPSI_exit_a2));
 sg13g2_nand2b_1 _4186_ (.Y(_0800_),
    .B(FpgaPins_Fpga_LIPSI_is_brnz_a3),
    .A_N(FpgaPins_Fpga_LIPSI_z_a2));
 sg13g2_a21oi_1 _4187_ (.A1(FpgaPins_Fpga_LIPSI_is_brz_a3),
    .A2(FpgaPins_Fpga_LIPSI_z_a2),
    .Y(_0801_),
    .B1(FpgaPins_Fpga_LIPSI_is_br_a3));
 sg13g2_nand2_1 _4188_ (.Y(_0802_),
    .A(_0800_),
    .B(_0801_));
 sg13g2_mux2_2 _4189_ (.A0(\FpgaPins_Fpga_LIPSI_pc_a2[0] ),
    .A1(\FpgaPins_Fpga_LIPSI_data_a2[0] ),
    .S(FpgaPins_Fpga_LIPSI_is_ret_a2),
    .X(_0803_));
 sg13g2_mux2_1 _4190_ (.A0(_0022_),
    .A1(_0803_),
    .S(_0698_),
    .X(_0804_));
 sg13g2_mux2_1 _4191_ (.A0(_0804_),
    .A1(_0021_),
    .S(net940),
    .X(_0805_));
 sg13g2_nand3b_1 _4192_ (.B(_0700_),
    .C(_0795_),
    .Y(_0806_),
    .A_N(net2));
 sg13g2_a21o_1 _4193_ (.A2(net943),
    .A1(_0020_),
    .B1(_0806_),
    .X(_0807_));
 sg13g2_a21o_1 _4194_ (.A2(_0805_),
    .A1(_0798_),
    .B1(_0807_),
    .X(_0808_));
 sg13g2_inv_1 _4195_ (.Y(\FpgaPins_Fpga_FSM_imem_rd_addr_a1[0] ),
    .A(net929));
 sg13g2_mux2_1 _4196_ (.A0(\FpgaPins_Fpga_LIPSI_pc_a2[1] ),
    .A1(\FpgaPins_Fpga_LIPSI_data_a2[1] ),
    .S(FpgaPins_Fpga_LIPSI_is_ret_a2),
    .X(_0809_));
 sg13g2_xor2_1 _4197_ (.B(_0809_),
    .A(_0803_),
    .X(_0810_));
 sg13g2_nand2_1 _4198_ (.Y(_0811_),
    .A(net986),
    .B(_0025_));
 sg13g2_and3_1 _4199_ (.X(_0812_),
    .A(_0800_),
    .B(_0801_),
    .C(_0811_));
 sg13g2_o21ai_1 _4200_ (.B1(_0812_),
    .Y(_0813_),
    .A1(net987),
    .A2(_0810_));
 sg13g2_a21oi_2 _4201_ (.B1(net943),
    .Y(_0814_),
    .A2(net941),
    .A1(_0702_));
 sg13g2_a21o_2 _4202_ (.A2(net943),
    .A1(_0023_),
    .B1(_0806_),
    .X(_0815_));
 sg13g2_a21oi_1 _4203_ (.A1(_0813_),
    .A2(_0814_),
    .Y(\FpgaPins_Fpga_FSM_imem_rd_addr_a1[1] ),
    .B1(_0815_));
 sg13g2_mux2_1 _4204_ (.A0(\FpgaPins_Fpga_LIPSI_pc_a2[2] ),
    .A1(\FpgaPins_Fpga_LIPSI_data_a2[2] ),
    .S(net990),
    .X(_0816_));
 sg13g2_a21oi_1 _4205_ (.A1(_0803_),
    .A2(_0809_),
    .Y(_0817_),
    .B1(_0816_));
 sg13g2_and3_1 _4206_ (.X(_0818_),
    .A(_0803_),
    .B(_0809_),
    .C(_0816_));
 sg13g2_or3_1 _4207_ (.A(net987),
    .B(_0817_),
    .C(_0818_),
    .X(_0819_));
 sg13g2_a21oi_1 _4208_ (.A1(net987),
    .A2(_0703_),
    .Y(_0820_),
    .B1(net941));
 sg13g2_a22oi_1 _4209_ (.Y(_0821_),
    .B1(_0819_),
    .B2(_0820_),
    .A2(net941),
    .A1(_0027_));
 sg13g2_a21oi_1 _4210_ (.A1(_0026_),
    .A2(net943),
    .Y(_0822_),
    .B1(_0806_));
 sg13g2_o21ai_1 _4211_ (.B1(_0822_),
    .Y(_0823_),
    .A1(net943),
    .A2(_0821_));
 sg13g2_inv_1 _4212_ (.Y(\FpgaPins_Fpga_FSM_imem_rd_addr_a1[2] ),
    .A(net906));
 sg13g2_mux4_1 _4213_ (.S0(net926),
    .A0(\instrs[9][1] ),
    .A1(\instrs[8][1] ),
    .A2(\instrs[11][1] ),
    .A3(\instrs[10][1] ),
    .S1(net920),
    .X(_0824_));
 sg13g2_and2_1 _4214_ (.A(net906),
    .B(_0824_),
    .X(_0825_));
 sg13g2_nand2_1 _4215_ (.Y(_0826_),
    .A(\instrs[13][1] ),
    .B(net913));
 sg13g2_a21oi_1 _4216_ (.A1(\instrs[12][1] ),
    .A2(net930),
    .Y(_0827_),
    .B1(net922));
 sg13g2_nand2_1 _4217_ (.Y(_0828_),
    .A(\instrs[14][1] ),
    .B(net930));
 sg13g2_a221oi_1 _4218_ (.B2(_0814_),
    .C1(_0815_),
    .B1(_0813_),
    .A1(\instrs[15][1] ),
    .Y(_0829_),
    .A2(net913));
 sg13g2_a221oi_1 _4219_ (.B2(_0829_),
    .C1(net910),
    .B1(_0828_),
    .A1(_0826_),
    .Y(_0830_),
    .A2(_0827_));
 sg13g2_nor2b_1 _4220_ (.A(net990),
    .B_N(_0029_),
    .Y(_0831_));
 sg13g2_a21oi_1 _4221_ (.A1(net990),
    .A2(_0032_),
    .Y(_0832_),
    .B1(_0831_));
 sg13g2_and2_1 _4222_ (.A(_0818_),
    .B(_0832_),
    .X(_0833_));
 sg13g2_o21ai_1 _4223_ (.B1(_0698_),
    .Y(_0834_),
    .A1(_0818_),
    .A2(_0832_));
 sg13g2_a21oi_1 _4224_ (.A1(net987),
    .A2(_0704_),
    .Y(_0835_),
    .B1(net941));
 sg13g2_o21ai_1 _4225_ (.B1(_0835_),
    .Y(_0836_),
    .A1(_0833_),
    .A2(_0834_));
 sg13g2_nand2_1 _4226_ (.Y(_0837_),
    .A(_0030_),
    .B(net941));
 sg13g2_a21oi_1 _4227_ (.A1(_0836_),
    .A2(_0837_),
    .Y(_0838_),
    .B1(net943));
 sg13g2_a21oi_1 _4228_ (.A1(net1752),
    .A2(net943),
    .Y(_0839_),
    .B1(_0806_));
 sg13g2_nand2b_2 _4229_ (.Y(_0840_),
    .B(_0839_),
    .A_N(_0838_));
 sg13g2_inv_1 _4230_ (.Y(\FpgaPins_Fpga_FSM_imem_rd_addr_a1[3] ),
    .A(net896));
 sg13g2_or3_1 _4231_ (.A(_0825_),
    .B(_0830_),
    .C(net896),
    .X(_0841_));
 sg13g2_mux4_1 _4232_ (.S0(net931),
    .A0(\instrs[1][1] ),
    .A1(\instrs[0][1] ),
    .A2(\instrs[3][1] ),
    .A3(\instrs[2][1] ),
    .S1(net923),
    .X(_0842_));
 sg13g2_and2_1 _4233_ (.A(net908),
    .B(_0842_),
    .X(_0843_));
 sg13g2_nand2_1 _4234_ (.Y(_0844_),
    .A(\instrs[5][1] ),
    .B(net914));
 sg13g2_a21oi_1 _4235_ (.A1(\instrs[4][1] ),
    .A2(net928),
    .Y(_0845_),
    .B1(net921));
 sg13g2_nand2_1 _4236_ (.Y(_0846_),
    .A(\instrs[6][1] ),
    .B(net928));
 sg13g2_a221oi_1 _4237_ (.B2(_0814_),
    .C1(_0815_),
    .B1(_0813_),
    .A1(\instrs[7][1] ),
    .Y(_0847_),
    .A2(net913));
 sg13g2_a221oi_1 _4238_ (.B2(_0847_),
    .C1(net908),
    .B1(_0846_),
    .A1(_0844_),
    .Y(_0848_),
    .A2(_0845_));
 sg13g2_or3_1 _4239_ (.A(\FpgaPins_Fpga_FSM_imem_rd_addr_a1[3] ),
    .B(_0843_),
    .C(_0848_),
    .X(_0849_));
 sg13g2_and2_2 _4240_ (.A(_0841_),
    .B(_0849_),
    .X(\FpgaPins_Fpga_FSM_instr_a1[1] ));
 sg13g2_inv_2 _4241_ (.Y(_0850_),
    .A(\FpgaPins_Fpga_FSM_instr_a1[1] ));
 sg13g2_mux4_1 _4242_ (.S0(net926),
    .A0(_0042_),
    .A1(_0041_),
    .A2(_0044_),
    .A3(_0043_),
    .S1(net920),
    .X(_0851_));
 sg13g2_nand2_1 _4243_ (.Y(_0852_),
    .A(net906),
    .B(_0851_));
 sg13g2_nand2_1 _4244_ (.Y(_0853_),
    .A(_0046_),
    .B(net912));
 sg13g2_a21oi_1 _4245_ (.A1(_0045_),
    .A2(net927),
    .Y(_0854_),
    .B1(net919));
 sg13g2_nand2_1 _4246_ (.Y(_0855_),
    .A(_0047_),
    .B(net925));
 sg13g2_a221oi_1 _4247_ (.B2(_0814_),
    .C1(_0815_),
    .B1(_0813_),
    .A1(_0048_),
    .Y(_0856_),
    .A2(net912));
 sg13g2_a221oi_1 _4248_ (.B2(_0856_),
    .C1(net907),
    .B1(_0855_),
    .A1(_0853_),
    .Y(_0857_),
    .A2(_0854_));
 sg13g2_nand3b_1 _4249_ (.B(net891),
    .C(_0852_),
    .Y(_0858_),
    .A_N(_0857_));
 sg13g2_mux4_1 _4250_ (.S0(net932),
    .A0(_0034_),
    .A1(_0033_),
    .A2(_0036_),
    .A3(_0035_),
    .S1(net924),
    .X(_0859_));
 sg13g2_and2_1 _4251_ (.A(net908),
    .B(_0859_),
    .X(_0860_));
 sg13g2_nand2_1 _4252_ (.Y(_0861_),
    .A(_0038_),
    .B(net913));
 sg13g2_a21oi_1 _4253_ (.A1(_0037_),
    .A2(net928),
    .Y(_0862_),
    .B1(net921));
 sg13g2_nand2_1 _4254_ (.Y(_0863_),
    .A(_0039_),
    .B(net930));
 sg13g2_a221oi_1 _4255_ (.B2(_0814_),
    .C1(_0815_),
    .B1(_0813_),
    .A1(_0040_),
    .Y(_0864_),
    .A2(net913));
 sg13g2_a221oi_1 _4256_ (.B2(_0864_),
    .C1(net910),
    .B1(_0863_),
    .A1(_0861_),
    .Y(_0865_),
    .A2(_0862_));
 sg13g2_or3_1 _4257_ (.A(net891),
    .B(_0860_),
    .C(_0865_),
    .X(_0866_));
 sg13g2_and2_2 _4258_ (.A(_0858_),
    .B(_0866_),
    .X(_0867_));
 sg13g2_inv_1 _4259_ (.Y(\FpgaPins_Fpga_FSM_instr_a1[0] ),
    .A(_0867_));
 sg13g2_and3_1 _4260_ (.X(_0868_),
    .A(net1164),
    .B(\FpgaPins_Fpga_GAME_count_speed4_a2[1] ),
    .C(net1207));
 sg13g2_and2_1 _4261_ (.A(net1513),
    .B(_0868_),
    .X(_0869_));
 sg13g2_and2_1 _4262_ (.A(net1366),
    .B(_0869_),
    .X(_0870_));
 sg13g2_and2_1 _4263_ (.A(net1551),
    .B(_0870_),
    .X(_0871_));
 sg13g2_and2_1 _4264_ (.A(net1389),
    .B(_0871_),
    .X(_0872_));
 sg13g2_and2_1 _4265_ (.A(net1417),
    .B(_0872_),
    .X(_0873_));
 sg13g2_and2_1 _4266_ (.A(net1607),
    .B(_0873_),
    .X(_0874_));
 sg13g2_and2_1 _4267_ (.A(net1574),
    .B(_0874_),
    .X(_0875_));
 sg13g2_and2_1 _4268_ (.A(net1621),
    .B(_0875_),
    .X(_0876_));
 sg13g2_and2_1 _4269_ (.A(net1554),
    .B(_0876_),
    .X(_0877_));
 sg13g2_and2_1 _4270_ (.A(net1565),
    .B(_0877_),
    .X(_0878_));
 sg13g2_and2_1 _4271_ (.A(net1599),
    .B(_0878_),
    .X(_0879_));
 sg13g2_nand2_1 _4272_ (.Y(_0880_),
    .A(\FpgaPins_Fpga_GAME_count_speed4_a2[13] ),
    .B(_0878_));
 sg13g2_nor2_1 _4273_ (.A(net1405),
    .B(_0880_),
    .Y(_0881_));
 sg13g2_nor4_1 _4274_ (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[11] ),
    .B(\FpgaPins_Fpga_GAME_count_speed4_a2[10] ),
    .C(_0706_),
    .D(\FpgaPins_Fpga_GAME_count_speed4_a2[9] ),
    .Y(_0882_));
 sg13g2_nand4_1 _4275_ (.B(\FpgaPins_Fpga_GAME_count_speed4_a2[16] ),
    .C(\FpgaPins_Fpga_GAME_count_speed4_a2[18] ),
    .A(\FpgaPins_Fpga_GAME_count_speed4_a2[17] ),
    .Y(_0883_),
    .D(_0882_));
 sg13g2_or4_1 _4276_ (.A(_0705_),
    .B(\FpgaPins_Fpga_GAME_count_speed4_a2[12] ),
    .C(\FpgaPins_Fpga_GAME_count_speed4_a2[7] ),
    .D(\FpgaPins_Fpga_GAME_count_speed4_a2[6] ),
    .X(_0884_));
 sg13g2_nor3_1 _4277_ (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[14] ),
    .B(\FpgaPins_Fpga_GAME_count_speed4_a2[1] ),
    .C(\FpgaPins_Fpga_GAME_count_speed4_a2[0] ),
    .Y(_0885_));
 sg13g2_nor3_1 _4278_ (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[4] ),
    .B(\FpgaPins_Fpga_GAME_count_speed4_a2[3] ),
    .C(\FpgaPins_Fpga_GAME_count_speed4_a2[2] ),
    .Y(_0886_));
 sg13g2_nand4_1 _4279_ (.B(\FpgaPins_Fpga_GAME_count_speed4_a2[15] ),
    .C(_0885_),
    .A(\FpgaPins_Fpga_GAME_count_speed4_a2[5] ),
    .Y(_0887_),
    .D(_0886_));
 sg13g2_or2_1 _4280_ (.X(_0888_),
    .B(_0887_),
    .A(_0884_));
 sg13g2_o21ai_1 _4281_ (.B1(net985),
    .Y(_0889_),
    .A1(_0883_),
    .A2(_0888_));
 sg13g2_inv_2 _4282_ (.Y(_0890_),
    .A(net916));
 sg13g2_o21ai_1 _4283_ (.B1(_0890_),
    .Y(_0891_),
    .A1(net1498),
    .A2(_0881_));
 sg13g2_a21oi_1 _4284_ (.A1(net1498),
    .A2(_0881_),
    .Y(\FpgaPins_Fpga_GAME_count_speed4_a1[15] ),
    .B1(_0891_));
 sg13g2_o21ai_1 _4285_ (.B1(_0890_),
    .Y(_0892_),
    .A1(net1599),
    .A2(_0878_));
 sg13g2_nor2_1 _4286_ (.A(_0879_),
    .B(_0892_),
    .Y(\FpgaPins_Fpga_GAME_count_speed4_a1[13] ));
 sg13g2_o21ai_1 _4287_ (.B1(_0890_),
    .Y(_0893_),
    .A1(net1607),
    .A2(_0873_));
 sg13g2_nor2_1 _4288_ (.A(_0874_),
    .B(_0893_),
    .Y(\FpgaPins_Fpga_GAME_count_speed4_a1[8] ));
 sg13g2_nor2_1 _4289_ (.A(net1551),
    .B(_0870_),
    .Y(_0894_));
 sg13g2_nor3_1 _4290_ (.A(_0871_),
    .B(net916),
    .C(_0894_),
    .Y(\FpgaPins_Fpga_GAME_count_speed4_a1[5] ));
 sg13g2_and2_1 _4291_ (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[14] ),
    .B(\FpgaPins_Fpga_GAME_count_speed4_a2[15] ),
    .X(_0895_));
 sg13g2_and3_1 _4292_ (.X(_0896_),
    .A(net1114),
    .B(_0879_),
    .C(_0895_));
 sg13g2_nor2_1 _4293_ (.A(net1503),
    .B(_0896_),
    .Y(_0897_));
 sg13g2_and2_1 _4294_ (.A(net1503),
    .B(_0896_),
    .X(_0898_));
 sg13g2_nor3_1 _4295_ (.A(net916),
    .B(_0897_),
    .C(_0898_),
    .Y(\FpgaPins_Fpga_GAME_count_speed4_a1[17] ));
 sg13g2_a21oi_1 _4296_ (.A1(_0879_),
    .A2(_0895_),
    .Y(_0899_),
    .B1(net1114));
 sg13g2_nor3_1 _4297_ (.A(net916),
    .B(_0896_),
    .C(net1115),
    .Y(\FpgaPins_Fpga_GAME_count_speed4_a1[16] ));
 sg13g2_o21ai_1 _4298_ (.B1(_0890_),
    .Y(_0900_),
    .A1(net1030),
    .A2(_0898_));
 sg13g2_a21oi_1 _4299_ (.A1(net1030),
    .A2(_0898_),
    .Y(\FpgaPins_Fpga_GAME_count_speed4_a1[18] ),
    .B1(_0900_));
 sg13g2_and3_1 _4300_ (.X(_0901_),
    .A(net1191),
    .B(net1091),
    .C(net1060));
 sg13g2_and2_1 _4301_ (.A(net1399),
    .B(_0901_),
    .X(_0902_));
 sg13g2_and2_2 _4302_ (.A(net1381),
    .B(_0902_),
    .X(_0903_));
 sg13g2_nand3_1 _4303_ (.B(\FpgaPins_Fpga_GAME_count_speed3_a2[5] ),
    .C(_0903_),
    .A(net1364),
    .Y(_0904_));
 sg13g2_nor2_1 _4304_ (.A(_0708_),
    .B(_0904_),
    .Y(_0905_));
 sg13g2_and2_1 _4305_ (.A(net1383),
    .B(_0905_),
    .X(_0906_));
 sg13g2_nand2_1 _4306_ (.Y(_0907_),
    .A(net1558),
    .B(net1383));
 sg13g2_nor3_2 _4307_ (.A(_0708_),
    .B(_0904_),
    .C(_0907_),
    .Y(_0908_));
 sg13g2_and2_1 _4308_ (.A(net1552),
    .B(_0908_),
    .X(_0909_));
 sg13g2_and2_1 _4309_ (.A(net1627),
    .B(_0909_),
    .X(_0910_));
 sg13g2_nand3_1 _4310_ (.B(net1756),
    .C(_0910_),
    .A(net1200),
    .Y(_0911_));
 sg13g2_inv_1 _4311_ (.Y(_0912_),
    .A(_0911_));
 sg13g2_nor2_1 _4312_ (.A(net1385),
    .B(_0911_),
    .Y(_0913_));
 sg13g2_nand4_1 _4313_ (.B(\FpgaPins_Fpga_GAME_count_speed3_a2[12] ),
    .C(\FpgaPins_Fpga_GAME_count_speed3_a2[11] ),
    .A(\FpgaPins_Fpga_GAME_count_speed3_a2[13] ),
    .Y(_0914_),
    .D(_0707_));
 sg13g2_nor4_1 _4314_ (.A(_0708_),
    .B(\FpgaPins_Fpga_GAME_count_speed3_a2[17] ),
    .C(_0907_),
    .D(_0914_),
    .Y(_0915_));
 sg13g2_and4_1 _4315_ (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[16] ),
    .B(\FpgaPins_Fpga_GAME_count_speed3_a2[18] ),
    .C(\FpgaPins_Fpga_GAME_count_speed3_a2[19] ),
    .D(_0915_),
    .X(_0916_));
 sg13g2_nor2_1 _4316_ (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[3] ),
    .B(\FpgaPins_Fpga_GAME_count_speed3_a2[2] ),
    .Y(_0917_));
 sg13g2_or2_1 _4317_ (.X(_0918_),
    .B(net1060),
    .A(net1091));
 sg13g2_nand2b_1 _4318_ (.Y(_0919_),
    .B(\FpgaPins_Fpga_GAME_count_speed3_a2[5] ),
    .A_N(\FpgaPins_Fpga_GAME_count_speed3_a2[4] ));
 sg13g2_nor4_1 _4319_ (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[14] ),
    .B(\FpgaPins_Fpga_GAME_count_speed3_a2[6] ),
    .C(_0918_),
    .D(_0919_),
    .Y(_0920_));
 sg13g2_nand4_1 _4320_ (.B(_0916_),
    .C(_0917_),
    .A(\FpgaPins_Fpga_GAME_count_speed3_a2[15] ),
    .Y(_0921_),
    .D(_0920_));
 sg13g2_nand2_1 _4321_ (.Y(_0922_),
    .A(net985),
    .B(_0921_));
 sg13g2_inv_2 _4322_ (.Y(_0923_),
    .A(net894));
 sg13g2_o21ai_1 _4323_ (.B1(_0923_),
    .Y(_0924_),
    .A1(net1684),
    .A2(_0913_));
 sg13g2_and2_1 _4324_ (.A(net1684),
    .B(_0913_),
    .X(_0925_));
 sg13g2_nor2_1 _4325_ (.A(_0924_),
    .B(_0925_),
    .Y(\FpgaPins_Fpga_GAME_count_speed3_a1[15] ));
 sg13g2_a21oi_1 _4326_ (.A1(\FpgaPins_Fpga_GAME_count_speed3_a2[12] ),
    .A2(_0910_),
    .Y(_0926_),
    .B1(net1200));
 sg13g2_nor3_1 _4327_ (.A(_0912_),
    .B(net895),
    .C(net1201),
    .Y(\FpgaPins_Fpga_GAME_count_speed3_a1[13] ));
 sg13g2_o21ai_1 _4328_ (.B1(_0923_),
    .Y(_0927_),
    .A1(net1395),
    .A2(_0910_));
 sg13g2_a21oi_1 _4329_ (.A1(net1395),
    .A2(_0910_),
    .Y(\FpgaPins_Fpga_GAME_count_speed3_a1[12] ),
    .B1(_0927_));
 sg13g2_o21ai_1 _4330_ (.B1(_0923_),
    .Y(_0928_),
    .A1(net1627),
    .A2(_0909_));
 sg13g2_nor2_1 _4331_ (.A(_0910_),
    .B(_0928_),
    .Y(\FpgaPins_Fpga_GAME_count_speed3_a1[11] ));
 sg13g2_o21ai_1 _4332_ (.B1(_0923_),
    .Y(_0929_),
    .A1(net1558),
    .A2(_0906_));
 sg13g2_nor2_1 _4333_ (.A(_0908_),
    .B(_0929_),
    .Y(\FpgaPins_Fpga_GAME_count_speed3_a1[9] ));
 sg13g2_nor2_1 _4334_ (.A(net1383),
    .B(_0905_),
    .Y(_0930_));
 sg13g2_nor3_1 _4335_ (.A(_0906_),
    .B(net894),
    .C(net1384),
    .Y(\FpgaPins_Fpga_GAME_count_speed3_a1[8] ));
 sg13g2_and2_1 _4336_ (.A(_0708_),
    .B(_0904_),
    .X(_0931_));
 sg13g2_nor3_1 _4337_ (.A(_0905_),
    .B(net894),
    .C(net1711),
    .Y(\FpgaPins_Fpga_GAME_count_speed3_a1[7] ));
 sg13g2_o21ai_1 _4338_ (.B1(_0923_),
    .Y(_0932_),
    .A1(net1404),
    .A2(_0903_));
 sg13g2_a21oi_1 _4339_ (.A1(net1404),
    .A2(_0903_),
    .Y(\FpgaPins_Fpga_GAME_count_speed3_a1[5] ),
    .B1(_0932_));
 sg13g2_and3_1 _4340_ (.X(_0933_),
    .A(\FpgaPins_Fpga_GAME_count_speed3_a2[14] ),
    .B(\FpgaPins_Fpga_GAME_count_speed3_a2[15] ),
    .C(_0912_));
 sg13g2_and2_1 _4341_ (.A(net1373),
    .B(_0933_),
    .X(_0934_));
 sg13g2_and2_1 _4342_ (.A(net1427),
    .B(_0934_),
    .X(_0935_));
 sg13g2_a21oi_1 _4343_ (.A1(\FpgaPins_Fpga_GAME_count_speed3_a2[18] ),
    .A2(_0935_),
    .Y(_0936_),
    .B1(net1265));
 sg13g2_and3_1 _4344_ (.X(_0937_),
    .A(\FpgaPins_Fpga_GAME_count_speed3_a2[18] ),
    .B(net1265),
    .C(_0935_));
 sg13g2_nor3_1 _4345_ (.A(net894),
    .B(net1266),
    .C(_0937_),
    .Y(\FpgaPins_Fpga_GAME_count_speed3_a1[19] ));
 sg13g2_xnor2_1 _4346_ (.Y(_0938_),
    .A(net1586),
    .B(_0935_));
 sg13g2_nor2_1 _4347_ (.A(net894),
    .B(_0938_),
    .Y(\FpgaPins_Fpga_GAME_count_speed3_a1[18] ));
 sg13g2_nor2_1 _4348_ (.A(net1373),
    .B(_0933_),
    .Y(_0939_));
 sg13g2_nor3_1 _4349_ (.A(net894),
    .B(_0934_),
    .C(net1374),
    .Y(\FpgaPins_Fpga_GAME_count_speed3_a1[16] ));
 sg13g2_and3_1 _4350_ (.X(_0940_),
    .A(net1127),
    .B(\FpgaPins_Fpga_GAME_count_speed2_a2[1] ),
    .C(net1190));
 sg13g2_and2_1 _4351_ (.A(net1452),
    .B(_0940_),
    .X(_0941_));
 sg13g2_and2_1 _4352_ (.A(net1368),
    .B(_0941_),
    .X(_0942_));
 sg13g2_inv_1 _4353_ (.Y(_0943_),
    .A(_0942_));
 sg13g2_and2_1 _4354_ (.A(net1391),
    .B(_0942_),
    .X(_0944_));
 sg13g2_and2_1 _4355_ (.A(net1521),
    .B(_0944_),
    .X(_0945_));
 sg13g2_and2_1 _4356_ (.A(net1484),
    .B(_0945_),
    .X(_0946_));
 sg13g2_and2_1 _4357_ (.A(net1500),
    .B(_0946_),
    .X(_0947_));
 sg13g2_and2_1 _4358_ (.A(net1377),
    .B(_0947_),
    .X(_0948_));
 sg13g2_and2_1 _4359_ (.A(net1441),
    .B(_0948_),
    .X(_0949_));
 sg13g2_and2_1 _4360_ (.A(net1402),
    .B(_0949_),
    .X(_0950_));
 sg13g2_and2_1 _4361_ (.A(net1564),
    .B(_0950_),
    .X(_0951_));
 sg13g2_and2_1 _4362_ (.A(net1566),
    .B(_0951_),
    .X(_0952_));
 sg13g2_nor2_1 _4363_ (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[18] ),
    .B(_0052_),
    .Y(_0953_));
 sg13g2_nand2b_1 _4364_ (.Y(_0954_),
    .B(\FpgaPins_Fpga_GAME_count_speed2_a2[7] ),
    .A_N(\FpgaPins_Fpga_GAME_count_speed2_a2[9] ));
 sg13g2_nor2_1 _4365_ (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[11] ),
    .B(\FpgaPins_Fpga_GAME_count_speed2_a2[10] ),
    .Y(_0955_));
 sg13g2_nand3_1 _4366_ (.B(\FpgaPins_Fpga_GAME_count_speed2_a2[12] ),
    .C(_0955_),
    .A(\FpgaPins_Fpga_GAME_count_speed2_a2[13] ),
    .Y(_0956_));
 sg13g2_nor4_1 _4367_ (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[8] ),
    .B(\FpgaPins_Fpga_GAME_count_speed2_a2[17] ),
    .C(_0954_),
    .D(_0956_),
    .Y(_0957_));
 sg13g2_nand4_1 _4368_ (.B(net1193),
    .C(_0953_),
    .A(\FpgaPins_Fpga_GAME_count_speed2_a2[16] ),
    .Y(_0958_),
    .D(_0957_));
 sg13g2_nor3_1 _4369_ (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[4] ),
    .B(\FpgaPins_Fpga_GAME_count_speed2_a2[3] ),
    .C(\FpgaPins_Fpga_GAME_count_speed2_a2[2] ),
    .Y(_0959_));
 sg13g2_and2_1 _4370_ (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[14] ),
    .B(\FpgaPins_Fpga_GAME_count_speed2_a2[15] ),
    .X(_0960_));
 sg13g2_nor3_1 _4371_ (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[6] ),
    .B(\FpgaPins_Fpga_GAME_count_speed2_a2[1] ),
    .C(\FpgaPins_Fpga_GAME_count_speed2_a2[0] ),
    .Y(_0961_));
 sg13g2_nand4_1 _4372_ (.B(_0959_),
    .C(_0960_),
    .A(\FpgaPins_Fpga_GAME_count_speed2_a2[5] ),
    .Y(_0962_),
    .D(_0961_));
 sg13g2_o21ai_1 _4373_ (.B1(net985),
    .Y(_0963_),
    .A1(_0958_),
    .A2(_0962_));
 sg13g2_nand3_1 _4374_ (.B(\FpgaPins_Fpga_GAME_count_speed2_a2[12] ),
    .C(_0950_),
    .A(\FpgaPins_Fpga_GAME_count_speed2_a2[13] ),
    .Y(_0964_));
 sg13g2_nor2_1 _4375_ (.A(net1346),
    .B(_0964_),
    .Y(_0965_));
 sg13g2_xnor2_1 _4376_ (.Y(_0966_),
    .A(net1540),
    .B(_0965_));
 sg13g2_nor2_1 _4377_ (.A(net905),
    .B(net1541),
    .Y(\FpgaPins_Fpga_GAME_count_speed2_a1[15] ));
 sg13g2_a21oi_1 _4378_ (.A1(net1346),
    .A2(_0964_),
    .Y(_0967_),
    .B1(net904));
 sg13g2_nor2b_1 _4379_ (.A(_0965_),
    .B_N(net1347),
    .Y(\FpgaPins_Fpga_GAME_count_speed2_a1[14] ));
 sg13g2_nor2_1 _4380_ (.A(net1566),
    .B(_0951_),
    .Y(_0968_));
 sg13g2_nor3_1 _4381_ (.A(_0952_),
    .B(net905),
    .C(_0968_),
    .Y(\FpgaPins_Fpga_GAME_count_speed2_a1[13] ));
 sg13g2_nor2_1 _4382_ (.A(net1564),
    .B(_0950_),
    .Y(_0969_));
 sg13g2_nor3_1 _4383_ (.A(_0951_),
    .B(net903),
    .C(_0969_),
    .Y(\FpgaPins_Fpga_GAME_count_speed2_a1[12] ));
 sg13g2_nor2_1 _4384_ (.A(net1484),
    .B(_0945_),
    .Y(_0970_));
 sg13g2_nor3_1 _4385_ (.A(_0946_),
    .B(net905),
    .C(net1485),
    .Y(\FpgaPins_Fpga_GAME_count_speed2_a1[7] ));
 sg13g2_nor2_1 _4386_ (.A(net1391),
    .B(_0942_),
    .Y(_0971_));
 sg13g2_nor3_1 _4387_ (.A(_0944_),
    .B(net904),
    .C(_0971_),
    .Y(\FpgaPins_Fpga_GAME_count_speed2_a1[5] ));
 sg13g2_and4_2 _4388_ (.A(net1443),
    .B(net1509),
    .C(_0952_),
    .D(_0960_),
    .X(_0972_));
 sg13g2_and4_1 _4389_ (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[13] ),
    .B(\FpgaPins_Fpga_GAME_count_speed2_a2[12] ),
    .C(_0950_),
    .D(_0960_),
    .X(_0973_));
 sg13g2_and2_1 _4390_ (.A(net1509),
    .B(_0973_),
    .X(_0974_));
 sg13g2_a21oi_1 _4391_ (.A1(\FpgaPins_Fpga_GAME_count_speed2_a2[18] ),
    .A2(_0972_),
    .Y(_0975_),
    .B1(net1193));
 sg13g2_nand3_1 _4392_ (.B(net1193),
    .C(_0972_),
    .A(\FpgaPins_Fpga_GAME_count_speed2_a2[18] ),
    .Y(_0976_));
 sg13g2_nand2b_1 _4393_ (.Y(_0977_),
    .B(_0976_),
    .A_N(net903));
 sg13g2_nor2_1 _4394_ (.A(net1194),
    .B(_0977_),
    .Y(\FpgaPins_Fpga_GAME_count_speed2_a1[19] ));
 sg13g2_nor2_1 _4395_ (.A(net1509),
    .B(_0973_),
    .Y(_0978_));
 sg13g2_nor3_1 _4396_ (.A(net903),
    .B(_0974_),
    .C(net1510),
    .Y(\FpgaPins_Fpga_GAME_count_speed2_a1[16] ));
 sg13g2_a21oi_1 _4397_ (.A1(net1422),
    .A2(_0976_),
    .Y(_0979_),
    .B1(net903));
 sg13g2_o21ai_1 _4398_ (.B1(_0979_),
    .Y(_0980_),
    .A1(net1422),
    .A2(_0976_));
 sg13g2_inv_1 _4399_ (.Y(\FpgaPins_Fpga_GAME_count_speed2_a1[20] ),
    .A(net1423));
 sg13g2_and2_1 _4400_ (.A(net1572),
    .B(_0768_),
    .X(_0981_));
 sg13g2_and2_1 _4401_ (.A(net1626),
    .B(_0981_),
    .X(_0982_));
 sg13g2_and2_1 _4402_ (.A(net1610),
    .B(_0982_),
    .X(_0983_));
 sg13g2_and2_1 _4403_ (.A(net1560),
    .B(_0983_),
    .X(_0984_));
 sg13g2_and2_1 _4404_ (.A(net1570),
    .B(_0984_),
    .X(_0985_));
 sg13g2_o21ai_1 _4405_ (.B1(net893),
    .Y(_0986_),
    .A1(net1570),
    .A2(_0984_));
 sg13g2_nor2_1 _4406_ (.A(_0985_),
    .B(_0986_),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[15] ));
 sg13g2_and2_1 _4407_ (.A(net1549),
    .B(_0985_),
    .X(_0987_));
 sg13g2_and4_1 _4408_ (.A(net1465),
    .B(net1511),
    .C(net1303),
    .D(_0987_),
    .X(_0988_));
 sg13g2_and3_1 _4409_ (.X(_0989_),
    .A(net1465),
    .B(net1303),
    .C(_0987_));
 sg13g2_nor2_1 _4410_ (.A(net1520),
    .B(_0988_),
    .Y(_0990_));
 sg13g2_and3_1 _4411_ (.X(_0991_),
    .A(net1511),
    .B(net1520),
    .C(_0989_));
 sg13g2_nor3_1 _4412_ (.A(net898),
    .B(_0990_),
    .C(_0991_),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[20] ));
 sg13g2_a21oi_1 _4413_ (.A1(\FpgaPins_Fpga_GAME_count_speed1_a2[17] ),
    .A2(_0987_),
    .Y(_0992_),
    .B1(net1303));
 sg13g2_nor3_1 _4414_ (.A(net898),
    .B(_0989_),
    .C(net1304),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[18] ));
 sg13g2_nor2_1 _4415_ (.A(net1511),
    .B(_0989_),
    .Y(_0993_));
 sg13g2_nor3_1 _4416_ (.A(net897),
    .B(_0988_),
    .C(_0993_),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[19] ));
 sg13g2_o21ai_1 _4417_ (.B1(net893),
    .Y(_0994_),
    .A1(net1465),
    .A2(_0987_));
 sg13g2_a21oi_1 _4418_ (.A1(net1465),
    .A2(_0987_),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[17] ),
    .B1(_0994_));
 sg13g2_mux4_1 _4419_ (.S0(net926),
    .A0(_0062_),
    .A1(_0061_),
    .A2(_0064_),
    .A3(_0063_),
    .S1(net920),
    .X(_0995_));
 sg13g2_nand2_1 _4420_ (.Y(_0996_),
    .A(_0066_),
    .B(net911));
 sg13g2_a21oi_1 _4421_ (.A1(_0065_),
    .A2(net925),
    .Y(_0997_),
    .B1(net918));
 sg13g2_nand2_1 _4422_ (.Y(_0998_),
    .A(_0067_),
    .B(net925));
 sg13g2_nand2_1 _4423_ (.Y(_0999_),
    .A(_0068_),
    .B(net911));
 sg13g2_nand3_1 _4424_ (.B(_0998_),
    .C(_0999_),
    .A(net918),
    .Y(_1000_));
 sg13g2_a21oi_1 _4425_ (.A1(_0996_),
    .A2(_0997_),
    .Y(_1001_),
    .B1(net907));
 sg13g2_a221oi_1 _4426_ (.B2(_1001_),
    .C1(net896),
    .B1(_1000_),
    .A1(net906),
    .Y(_1002_),
    .A2(_0995_));
 sg13g2_mux4_1 _4427_ (.S0(net931),
    .A0(_0054_),
    .A1(_0053_),
    .A2(_0056_),
    .A3(_0055_),
    .S1(net923),
    .X(_1003_));
 sg13g2_nand2_1 _4428_ (.Y(_1004_),
    .A(_0058_),
    .B(net915));
 sg13g2_a21oi_1 _4429_ (.A1(_0057_),
    .A2(net929),
    .Y(_1005_),
    .B1(net921));
 sg13g2_nand2_1 _4430_ (.Y(_1006_),
    .A(_0059_),
    .B(net930));
 sg13g2_nand2_1 _4431_ (.Y(_1007_),
    .A(_0060_),
    .B(net913));
 sg13g2_nand3_1 _4432_ (.B(_1006_),
    .C(_1007_),
    .A(net922),
    .Y(_1008_));
 sg13g2_a21oi_1 _4433_ (.A1(_1004_),
    .A2(_1005_),
    .Y(_1009_),
    .B1(net910));
 sg13g2_a221oi_1 _4434_ (.B2(_1009_),
    .C1(net891),
    .B1(_1008_),
    .A1(net910),
    .Y(_1010_),
    .A2(_1003_));
 sg13g2_or2_2 _4435_ (.X(\FpgaPins_Fpga_FSM_instr_a1[5] ),
    .B(_1010_),
    .A(_1002_));
 sg13g2_mux4_1 _4436_ (.S0(net926),
    .A0(\instrs[9][3] ),
    .A1(\instrs[8][3] ),
    .A2(\instrs[11][3] ),
    .A3(\instrs[10][3] ),
    .S1(net920),
    .X(_1011_));
 sg13g2_nand2_1 _4437_ (.Y(_1012_),
    .A(\instrs[13][3] ),
    .B(net913));
 sg13g2_a21oi_1 _4438_ (.A1(\instrs[12][3] ),
    .A2(net930),
    .Y(_1013_),
    .B1(net922));
 sg13g2_nand2_1 _4439_ (.Y(_1014_),
    .A(\instrs[14][3] ),
    .B(net930));
 sg13g2_nand2_1 _4440_ (.Y(_1015_),
    .A(\instrs[15][3] ),
    .B(net915));
 sg13g2_nand3_1 _4441_ (.B(_1014_),
    .C(_1015_),
    .A(net922),
    .Y(_1016_));
 sg13g2_a21oi_1 _4442_ (.A1(_1012_),
    .A2(_1013_),
    .Y(_1017_),
    .B1(net910));
 sg13g2_a221oi_1 _4443_ (.B2(_1017_),
    .C1(net896),
    .B1(_1016_),
    .A1(net907),
    .Y(_1018_),
    .A2(_1011_));
 sg13g2_mux4_1 _4444_ (.S0(net931),
    .A0(\instrs[1][3] ),
    .A1(\instrs[0][3] ),
    .A2(\instrs[3][3] ),
    .A3(\instrs[2][3] ),
    .S1(net923),
    .X(_1019_));
 sg13g2_nand2_1 _4445_ (.Y(_1020_),
    .A(\instrs[5][3] ),
    .B(net915));
 sg13g2_a21oi_1 _4446_ (.A1(\instrs[4][3] ),
    .A2(net929),
    .Y(_1021_),
    .B1(net923));
 sg13g2_and2_1 _4447_ (.A(\instrs[6][3] ),
    .B(net929),
    .X(_1022_));
 sg13g2_a21oi_1 _4448_ (.A1(\instrs[7][3] ),
    .A2(net914),
    .Y(_1023_),
    .B1(_1022_));
 sg13g2_a221oi_1 _4449_ (.B2(net922),
    .C1(net909),
    .B1(_1023_),
    .A1(_1020_),
    .Y(_1024_),
    .A2(_1021_));
 sg13g2_a21oi_2 _4450_ (.B1(_1024_),
    .Y(_1025_),
    .A2(_1019_),
    .A1(net909));
 sg13g2_a21o_2 _4451_ (.A2(_1025_),
    .A1(_0840_),
    .B1(_1018_),
    .X(_1026_));
 sg13g2_inv_1 _4452_ (.Y(\FpgaPins_Fpga_FSM_instr_a1[3] ),
    .A(_1026_));
 sg13g2_mux4_1 _4453_ (.S0(net926),
    .A0(\instrs[9][2] ),
    .A1(\instrs[8][2] ),
    .A2(\instrs[11][2] ),
    .A3(\instrs[10][2] ),
    .S1(net924),
    .X(_1027_));
 sg13g2_nand2_1 _4454_ (.Y(_1028_),
    .A(\instrs[13][2] ),
    .B(net911));
 sg13g2_a21oi_1 _4455_ (.A1(\instrs[12][2] ),
    .A2(net925),
    .Y(_1029_),
    .B1(net918));
 sg13g2_nand2_1 _4456_ (.Y(_1030_),
    .A(\instrs[14][2] ),
    .B(net930));
 sg13g2_nand2_1 _4457_ (.Y(_1031_),
    .A(\instrs[15][2] ),
    .B(net912));
 sg13g2_nand3_1 _4458_ (.B(_1030_),
    .C(_1031_),
    .A(net919),
    .Y(_1032_));
 sg13g2_a21oi_1 _4459_ (.A1(_1028_),
    .A2(_1029_),
    .Y(_1033_),
    .B1(net907));
 sg13g2_a221oi_1 _4460_ (.B2(_1033_),
    .C1(_0840_),
    .B1(_1032_),
    .A1(net907),
    .Y(_1034_),
    .A2(_1027_));
 sg13g2_mux4_1 _4461_ (.S0(net932),
    .A0(\instrs[1][2] ),
    .A1(\instrs[0][2] ),
    .A2(\instrs[3][2] ),
    .A3(\instrs[2][2] ),
    .S1(net924),
    .X(_1035_));
 sg13g2_nand2_1 _4462_ (.Y(_1036_),
    .A(\instrs[5][2] ),
    .B(net914));
 sg13g2_a21oi_1 _4463_ (.A1(\instrs[4][2] ),
    .A2(net928),
    .Y(_1037_),
    .B1(net921));
 sg13g2_nand2_1 _4464_ (.Y(_1038_),
    .A(\instrs[6][2] ),
    .B(net928));
 sg13g2_nand2_1 _4465_ (.Y(_1039_),
    .A(\instrs[7][2] ),
    .B(net914));
 sg13g2_nand3_1 _4466_ (.B(_1038_),
    .C(_1039_),
    .A(net921),
    .Y(_1040_));
 sg13g2_a21oi_1 _4467_ (.A1(_1036_),
    .A2(_1037_),
    .Y(_1041_),
    .B1(net908));
 sg13g2_a22oi_1 _4468_ (.Y(_1042_),
    .B1(_1040_),
    .B2(_1041_),
    .A2(_1035_),
    .A1(net908));
 sg13g2_a21o_2 _4469_ (.A2(_1042_),
    .A1(_0840_),
    .B1(_1034_),
    .X(_1043_));
 sg13g2_inv_1 _4470_ (.Y(\FpgaPins_Fpga_FSM_instr_a1[2] ),
    .A(_1043_));
 sg13g2_mux4_1 _4471_ (.S0(net926),
    .A0(\instrs[9][4] ),
    .A1(\instrs[8][4] ),
    .A2(\instrs[11][4] ),
    .A3(\instrs[10][4] ),
    .S1(net924),
    .X(_1044_));
 sg13g2_nand2_1 _4472_ (.Y(_1045_),
    .A(\instrs[13][4] ),
    .B(net912));
 sg13g2_a21oi_1 _4473_ (.A1(\instrs[12][4] ),
    .A2(net927),
    .Y(_1046_),
    .B1(net919));
 sg13g2_nand2_1 _4474_ (.Y(_1047_),
    .A(\instrs[14][4] ),
    .B(net927));
 sg13g2_nand2_1 _4475_ (.Y(_1048_),
    .A(\instrs[15][4] ),
    .B(net912));
 sg13g2_nand3_1 _4476_ (.B(_1047_),
    .C(_1048_),
    .A(net919),
    .Y(_1049_));
 sg13g2_a21oi_1 _4477_ (.A1(_1045_),
    .A2(_1046_),
    .Y(_1050_),
    .B1(net907));
 sg13g2_a221oi_1 _4478_ (.B2(_1050_),
    .C1(net896),
    .B1(_1049_),
    .A1(net907),
    .Y(_1051_),
    .A2(_1044_));
 sg13g2_mux4_1 _4479_ (.S0(net931),
    .A0(\instrs[1][4] ),
    .A1(\instrs[0][4] ),
    .A2(\instrs[3][4] ),
    .A3(\instrs[2][4] ),
    .S1(net923),
    .X(_1052_));
 sg13g2_nand2_1 _4480_ (.Y(_1053_),
    .A(\instrs[5][4] ),
    .B(net915));
 sg13g2_a21oi_1 _4481_ (.A1(\instrs[4][4] ),
    .A2(net929),
    .Y(_1054_),
    .B1(net922));
 sg13g2_nand2_1 _4482_ (.Y(_1055_),
    .A(\instrs[6][4] ),
    .B(net929));
 sg13g2_nand2_1 _4483_ (.Y(_1056_),
    .A(\instrs[7][4] ),
    .B(net914));
 sg13g2_nand3_1 _4484_ (.B(_1055_),
    .C(_1056_),
    .A(net921),
    .Y(_1057_));
 sg13g2_a21oi_1 _4485_ (.A1(_1053_),
    .A2(_1054_),
    .Y(_1058_),
    .B1(net909));
 sg13g2_a221oi_1 _4486_ (.B2(_1058_),
    .C1(net891),
    .B1(_1057_),
    .A1(net908),
    .Y(_1059_),
    .A2(_1052_));
 sg13g2_or2_2 _4487_ (.X(_1060_),
    .B(_1059_),
    .A(_1051_));
 sg13g2_inv_1 _4488_ (.Y(\FpgaPins_Fpga_FSM_instr_a1[4] ),
    .A(_1060_));
 sg13g2_mux4_1 _4489_ (.S0(net926),
    .A0(_0078_),
    .A1(_0077_),
    .A2(_0080_),
    .A3(_0079_),
    .S1(net920),
    .X(_1061_));
 sg13g2_nand2_1 _4490_ (.Y(_1062_),
    .A(net906),
    .B(_1061_));
 sg13g2_nand2_1 _4491_ (.Y(_1063_),
    .A(_0082_),
    .B(net911));
 sg13g2_a21oi_1 _4492_ (.A1(_0081_),
    .A2(net925),
    .Y(_1064_),
    .B1(net918));
 sg13g2_nand2_1 _4493_ (.Y(_1065_),
    .A(_0083_),
    .B(net925));
 sg13g2_a221oi_1 _4494_ (.B2(_0814_),
    .C1(_0815_),
    .B1(_0813_),
    .A1(_0084_),
    .Y(_1066_),
    .A2(net912));
 sg13g2_a221oi_1 _4495_ (.B2(_1066_),
    .C1(net906),
    .B1(_1065_),
    .A1(_1063_),
    .Y(_1067_),
    .A2(_1064_));
 sg13g2_nand3b_1 _4496_ (.B(net891),
    .C(_1062_),
    .Y(_1068_),
    .A_N(_1067_));
 sg13g2_mux4_1 _4497_ (.S0(net931),
    .A0(_0070_),
    .A1(_0069_),
    .A2(_0072_),
    .A3(_0071_),
    .S1(net923),
    .X(_1069_));
 sg13g2_and2_1 _4498_ (.A(net909),
    .B(_1069_),
    .X(_1070_));
 sg13g2_nand2_1 _4499_ (.Y(_1071_),
    .A(_0074_),
    .B(net914));
 sg13g2_a21oi_1 _4500_ (.A1(_0073_),
    .A2(net928),
    .Y(_1072_),
    .B1(net922));
 sg13g2_nand2_1 _4501_ (.Y(_1073_),
    .A(_0075_),
    .B(net930));
 sg13g2_a221oi_1 _4502_ (.B2(_0814_),
    .C1(_0815_),
    .B1(_0813_),
    .A1(_0076_),
    .Y(_1074_),
    .A2(net913));
 sg13g2_a221oi_1 _4503_ (.B2(_1074_),
    .C1(net910),
    .B1(_1073_),
    .A1(_1071_),
    .Y(_1075_),
    .A2(_1072_));
 sg13g2_or3_2 _4504_ (.A(net891),
    .B(_1070_),
    .C(_1075_),
    .X(_1076_));
 sg13g2_nand2_1 _4505_ (.Y(\FpgaPins_Fpga_FSM_instr_a1[7] ),
    .A(_1068_),
    .B(_1076_));
 sg13g2_mux4_1 _4506_ (.S0(net926),
    .A0(\instrs[9][6] ),
    .A1(\instrs[8][6] ),
    .A2(\instrs[11][6] ),
    .A3(\instrs[10][6] ),
    .S1(net920),
    .X(_1077_));
 sg13g2_nand2_1 _4507_ (.Y(_1078_),
    .A(\instrs[13][6] ),
    .B(net911));
 sg13g2_a21oi_1 _4508_ (.A1(\instrs[12][6] ),
    .A2(net925),
    .Y(_1079_),
    .B1(net918));
 sg13g2_nand2_1 _4509_ (.Y(_1080_),
    .A(\instrs[14][6] ),
    .B(net925));
 sg13g2_nand2_1 _4510_ (.Y(_1081_),
    .A(\instrs[15][6] ),
    .B(net911));
 sg13g2_nand3_1 _4511_ (.B(_1080_),
    .C(_1081_),
    .A(net918),
    .Y(_1082_));
 sg13g2_a21oi_1 _4512_ (.A1(_1078_),
    .A2(_1079_),
    .Y(_1083_),
    .B1(net906));
 sg13g2_a221oi_1 _4513_ (.B2(_1083_),
    .C1(net896),
    .B1(_1082_),
    .A1(net906),
    .Y(_1084_),
    .A2(_1077_));
 sg13g2_mux4_1 _4514_ (.S0(net931),
    .A0(\instrs[1][6] ),
    .A1(\instrs[0][6] ),
    .A2(\instrs[3][6] ),
    .A3(\instrs[2][6] ),
    .S1(net923),
    .X(_1085_));
 sg13g2_nand2_1 _4515_ (.Y(_1086_),
    .A(\instrs[5][6] ),
    .B(net914));
 sg13g2_a21oi_1 _4516_ (.A1(\instrs[4][6] ),
    .A2(net928),
    .Y(_1087_),
    .B1(net921));
 sg13g2_nand2_1 _4517_ (.Y(_1088_),
    .A(\instrs[6][6] ),
    .B(net928));
 sg13g2_nand2_1 _4518_ (.Y(_1089_),
    .A(\instrs[7][6] ),
    .B(net914));
 sg13g2_nand3_1 _4519_ (.B(_1088_),
    .C(_1089_),
    .A(net921),
    .Y(_1090_));
 sg13g2_a21oi_1 _4520_ (.A1(_1086_),
    .A2(_1087_),
    .Y(_1091_),
    .B1(net908));
 sg13g2_a22oi_1 _4521_ (.Y(_1092_),
    .B1(_1090_),
    .B2(_1091_),
    .A2(_1085_),
    .A1(net908));
 sg13g2_a21oi_2 _4522_ (.B1(_1084_),
    .Y(\FpgaPins_Fpga_FSM_instr_a1[6] ),
    .A2(_1092_),
    .A1(net896));
 sg13g2_nor2_1 _4523_ (.A(net1207),
    .B(net917),
    .Y(\FpgaPins_Fpga_GAME_count_speed4_a1[0] ));
 sg13g2_xnor2_1 _4524_ (.Y(_1093_),
    .A(net1612),
    .B(net1207));
 sg13g2_nor2_1 _4525_ (.A(net917),
    .B(_1093_),
    .Y(\FpgaPins_Fpga_GAME_count_speed4_a1[1] ));
 sg13g2_a21oi_1 _4526_ (.A1(\FpgaPins_Fpga_GAME_count_speed4_a2[1] ),
    .A2(\FpgaPins_Fpga_GAME_count_speed4_a2[0] ),
    .Y(_1094_),
    .B1(net1164));
 sg13g2_nor3_1 _4527_ (.A(_0868_),
    .B(net917),
    .C(net1165),
    .Y(\FpgaPins_Fpga_GAME_count_speed4_a1[2] ));
 sg13g2_nor2_1 _4528_ (.A(net1513),
    .B(_0868_),
    .Y(_1095_));
 sg13g2_nor3_1 _4529_ (.A(_0869_),
    .B(net917),
    .C(net1514),
    .Y(\FpgaPins_Fpga_GAME_count_speed4_a1[3] ));
 sg13g2_nor2_1 _4530_ (.A(net1366),
    .B(_0869_),
    .Y(_1096_));
 sg13g2_nor3_1 _4531_ (.A(_0870_),
    .B(net916),
    .C(net1367),
    .Y(\FpgaPins_Fpga_GAME_count_speed4_a1[4] ));
 sg13g2_nor2_1 _4532_ (.A(net1389),
    .B(_0871_),
    .Y(_1097_));
 sg13g2_nor3_1 _4533_ (.A(_0872_),
    .B(net916),
    .C(net1390),
    .Y(\FpgaPins_Fpga_GAME_count_speed4_a1[6] ));
 sg13g2_nor2_1 _4534_ (.A(net1417),
    .B(_0872_),
    .Y(_1098_));
 sg13g2_nor3_1 _4535_ (.A(_0873_),
    .B(net916),
    .C(_1098_),
    .Y(\FpgaPins_Fpga_GAME_count_speed4_a1[7] ));
 sg13g2_o21ai_1 _4536_ (.B1(_0890_),
    .Y(_1099_),
    .A1(net1574),
    .A2(_0874_));
 sg13g2_nor2_1 _4537_ (.A(_0875_),
    .B(net1575),
    .Y(\FpgaPins_Fpga_GAME_count_speed4_a1[9] ));
 sg13g2_o21ai_1 _4538_ (.B1(_0890_),
    .Y(_1100_),
    .A1(net1621),
    .A2(_0875_));
 sg13g2_nor2_1 _4539_ (.A(_0876_),
    .B(_1100_),
    .Y(\FpgaPins_Fpga_GAME_count_speed4_a1[10] ));
 sg13g2_o21ai_1 _4540_ (.B1(_0890_),
    .Y(_1101_),
    .A1(net1554),
    .A2(_0876_));
 sg13g2_nor2_1 _4541_ (.A(_0877_),
    .B(net1555),
    .Y(\FpgaPins_Fpga_GAME_count_speed4_a1[11] ));
 sg13g2_o21ai_1 _4542_ (.B1(_0890_),
    .Y(_1102_),
    .A1(net1565),
    .A2(_0877_));
 sg13g2_nor2_1 _4543_ (.A(_0878_),
    .B(_1102_),
    .Y(\FpgaPins_Fpga_GAME_count_speed4_a1[12] ));
 sg13g2_a21oi_1 _4544_ (.A1(net1405),
    .A2(_0880_),
    .Y(_1103_),
    .B1(net916));
 sg13g2_nand2b_1 _4545_ (.Y(_1104_),
    .B(net1406),
    .A_N(_0881_));
 sg13g2_inv_1 _4546_ (.Y(\FpgaPins_Fpga_GAME_count_speed4_a1[14] ),
    .A(_1104_));
 sg13g2_nor2_1 _4547_ (.A(net1060),
    .B(net895),
    .Y(\FpgaPins_Fpga_GAME_count_speed3_a1[0] ));
 sg13g2_nand2_1 _4548_ (.Y(_1105_),
    .A(net985),
    .B(_0918_));
 sg13g2_a21oi_1 _4549_ (.A1(net1091),
    .A2(net1060),
    .Y(\FpgaPins_Fpga_GAME_count_speed3_a1[1] ),
    .B1(_1105_));
 sg13g2_a21oi_1 _4550_ (.A1(net1091),
    .A2(net1060),
    .Y(_1106_),
    .B1(net1191));
 sg13g2_nor3_1 _4551_ (.A(_0901_),
    .B(net895),
    .C(_1106_),
    .Y(\FpgaPins_Fpga_GAME_count_speed3_a1[2] ));
 sg13g2_nor2_1 _4552_ (.A(net1399),
    .B(_0901_),
    .Y(_1107_));
 sg13g2_nor3_1 _4553_ (.A(_0902_),
    .B(net895),
    .C(_1107_),
    .Y(\FpgaPins_Fpga_GAME_count_speed3_a1[3] ));
 sg13g2_nor2_1 _4554_ (.A(net1381),
    .B(_0902_),
    .Y(_1108_));
 sg13g2_nor3_1 _4555_ (.A(_0903_),
    .B(net895),
    .C(net1382),
    .Y(\FpgaPins_Fpga_GAME_count_speed3_a1[4] ));
 sg13g2_a21oi_1 _4556_ (.A1(\FpgaPins_Fpga_GAME_count_speed3_a2[5] ),
    .A2(_0903_),
    .Y(_1109_),
    .B1(net1364));
 sg13g2_nand2_1 _4557_ (.Y(_1110_),
    .A(_0904_),
    .B(_0923_));
 sg13g2_nor2_1 _4558_ (.A(net1365),
    .B(_1110_),
    .Y(\FpgaPins_Fpga_GAME_count_speed3_a1[6] ));
 sg13g2_o21ai_1 _4559_ (.B1(_0923_),
    .Y(_1111_),
    .A1(net1552),
    .A2(_0908_));
 sg13g2_nor2_1 _4560_ (.A(_0909_),
    .B(net1553),
    .Y(\FpgaPins_Fpga_GAME_count_speed3_a1[10] ));
 sg13g2_and2_1 _4561_ (.A(net1385),
    .B(_0911_),
    .X(_1112_));
 sg13g2_nor3_1 _4562_ (.A(_0913_),
    .B(net894),
    .C(net1386),
    .Y(\FpgaPins_Fpga_GAME_count_speed3_a1[14] ));
 sg13g2_nor2_1 _4563_ (.A(net1427),
    .B(_0934_),
    .Y(_1113_));
 sg13g2_nor3_1 _4564_ (.A(net894),
    .B(_0935_),
    .C(net1428),
    .Y(\FpgaPins_Fpga_GAME_count_speed3_a1[17] ));
 sg13g2_nor2_1 _4565_ (.A(net1190),
    .B(net904),
    .Y(\FpgaPins_Fpga_GAME_count_speed2_a1[0] ));
 sg13g2_xnor2_1 _4566_ (.Y(_1114_),
    .A(net1593),
    .B(net1190));
 sg13g2_nor2_1 _4567_ (.A(net904),
    .B(_1114_),
    .Y(\FpgaPins_Fpga_GAME_count_speed2_a1[1] ));
 sg13g2_a21oi_1 _4568_ (.A1(\FpgaPins_Fpga_GAME_count_speed2_a2[1] ),
    .A2(\FpgaPins_Fpga_GAME_count_speed2_a2[0] ),
    .Y(_1115_),
    .B1(net1127));
 sg13g2_nor3_1 _4569_ (.A(_0940_),
    .B(net904),
    .C(net1128),
    .Y(\FpgaPins_Fpga_GAME_count_speed2_a1[2] ));
 sg13g2_nor2_1 _4570_ (.A(net1452),
    .B(_0940_),
    .Y(_1116_));
 sg13g2_nor3_1 _4571_ (.A(_0941_),
    .B(net904),
    .C(net1453),
    .Y(\FpgaPins_Fpga_GAME_count_speed2_a1[3] ));
 sg13g2_nor2_1 _4572_ (.A(net1368),
    .B(_0941_),
    .Y(_1117_));
 sg13g2_nor3_1 _4573_ (.A(_0942_),
    .B(net904),
    .C(net1369),
    .Y(\FpgaPins_Fpga_GAME_count_speed2_a1[4] ));
 sg13g2_nor2_1 _4574_ (.A(net1521),
    .B(_0944_),
    .Y(_1118_));
 sg13g2_nor3_1 _4575_ (.A(_0945_),
    .B(net904),
    .C(_1118_),
    .Y(\FpgaPins_Fpga_GAME_count_speed2_a1[6] ));
 sg13g2_nor2_1 _4576_ (.A(net1500),
    .B(_0946_),
    .Y(_1119_));
 sg13g2_nor3_1 _4577_ (.A(_0947_),
    .B(net903),
    .C(_1119_),
    .Y(\FpgaPins_Fpga_GAME_count_speed2_a1[8] ));
 sg13g2_nor2_1 _4578_ (.A(net1377),
    .B(_0947_),
    .Y(_1120_));
 sg13g2_nor3_1 _4579_ (.A(_0948_),
    .B(net903),
    .C(net1378),
    .Y(\FpgaPins_Fpga_GAME_count_speed2_a1[9] ));
 sg13g2_nor2_1 _4580_ (.A(net1441),
    .B(_0948_),
    .Y(_1121_));
 sg13g2_nor3_1 _4581_ (.A(_0949_),
    .B(net905),
    .C(_1121_),
    .Y(\FpgaPins_Fpga_GAME_count_speed2_a1[10] ));
 sg13g2_nor2_1 _4582_ (.A(net1402),
    .B(_0949_),
    .Y(_1122_));
 sg13g2_nor3_1 _4583_ (.A(_0950_),
    .B(net905),
    .C(net1403),
    .Y(\FpgaPins_Fpga_GAME_count_speed2_a1[11] ));
 sg13g2_nor2_1 _4584_ (.A(net1443),
    .B(_0974_),
    .Y(_1123_));
 sg13g2_nor3_1 _4585_ (.A(net903),
    .B(_0972_),
    .C(net1444),
    .Y(\FpgaPins_Fpga_GAME_count_speed2_a1[17] ));
 sg13g2_xnor2_1 _4586_ (.Y(_1124_),
    .A(net1609),
    .B(_0972_));
 sg13g2_nor2_1 _4587_ (.A(net903),
    .B(_1124_),
    .Y(\FpgaPins_Fpga_GAME_count_speed2_a1[18] ));
 sg13g2_nor2_1 _4588_ (.A(net725),
    .B(net897),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[0] ));
 sg13g2_nor3_1 _4589_ (.A(_0759_),
    .B(_0770_),
    .C(net897),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[1] ));
 sg13g2_nor2_1 _4590_ (.A(net1432),
    .B(_0759_),
    .Y(_1125_));
 sg13g2_nor3_1 _4591_ (.A(_0760_),
    .B(net897),
    .C(net1433),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[2] ));
 sg13g2_nor2_1 _4592_ (.A(net1446),
    .B(_0760_),
    .Y(_1126_));
 sg13g2_nor3_1 _4593_ (.A(_0761_),
    .B(net897),
    .C(_1126_),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[3] ));
 sg13g2_nor2_1 _4594_ (.A(net1450),
    .B(_0761_),
    .Y(_1127_));
 sg13g2_nor3_1 _4595_ (.A(_0762_),
    .B(net897),
    .C(_1127_),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[4] ));
 sg13g2_nor2_1 _4596_ (.A(net1494),
    .B(_0762_),
    .Y(_1128_));
 sg13g2_nor3_1 _4597_ (.A(_0763_),
    .B(net897),
    .C(_1128_),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[5] ));
 sg13g2_nor2_1 _4598_ (.A(net1393),
    .B(_0763_),
    .Y(_1129_));
 sg13g2_nor3_1 _4599_ (.A(_0764_),
    .B(net897),
    .C(net1394),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[6] ));
 sg13g2_o21ai_1 _4600_ (.B1(net892),
    .Y(_1130_),
    .A1(net1579),
    .A2(_0765_));
 sg13g2_nor2_1 _4601_ (.A(_0766_),
    .B(net1580),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[8] ));
 sg13g2_o21ai_1 _4602_ (.B1(net892),
    .Y(_1131_),
    .A1(net1556),
    .A2(_0766_));
 sg13g2_nor2_1 _4603_ (.A(_0767_),
    .B(net1557),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[9] ));
 sg13g2_o21ai_1 _4604_ (.B1(net892),
    .Y(_1132_),
    .A1(net1572),
    .A2(_0768_));
 sg13g2_nor2_1 _4605_ (.A(_0981_),
    .B(net1573),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[11] ));
 sg13g2_o21ai_1 _4606_ (.B1(net892),
    .Y(_1133_),
    .A1(net1626),
    .A2(_0981_));
 sg13g2_nor2_1 _4607_ (.A(_0982_),
    .B(_1133_),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[12] ));
 sg13g2_o21ai_1 _4608_ (.B1(net893),
    .Y(_1134_),
    .A1(net1610),
    .A2(_0982_));
 sg13g2_nor2_1 _4609_ (.A(_0983_),
    .B(net1611),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[13] ));
 sg13g2_o21ai_1 _4610_ (.B1(net893),
    .Y(_1135_),
    .A1(net1560),
    .A2(_0983_));
 sg13g2_nor2_1 _4611_ (.A(_0984_),
    .B(net1561),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[14] ));
 sg13g2_o21ai_1 _4612_ (.B1(net893),
    .Y(_1136_),
    .A1(net1549),
    .A2(_0985_));
 sg13g2_nor2_1 _4613_ (.A(_0987_),
    .B(net1550),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[16] ));
 sg13g2_o21ai_1 _4614_ (.B1(net892),
    .Y(_1137_),
    .A1(net1361),
    .A2(_0991_));
 sg13g2_a21oi_1 _4615_ (.A1(net1361),
    .A2(_0991_),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[21] ),
    .B1(_1137_));
 sg13g2_a21o_1 _4616_ (.A2(_0991_),
    .A1(net1361),
    .B1(net1677),
    .X(_1138_));
 sg13g2_nand3_1 _4617_ (.B(net1677),
    .C(_0991_),
    .A(net1361),
    .Y(_1139_));
 sg13g2_and3_1 _4618_ (.X(\FpgaPins_Fpga_GAME_count_speed1_a1[22] ),
    .A(net892),
    .B(_1138_),
    .C(_1139_));
 sg13g2_xor2_1 _4619_ (.B(_1139_),
    .A(net1522),
    .X(_1140_));
 sg13g2_nor2_1 _4620_ (.A(net898),
    .B(net1523),
    .Y(\FpgaPins_Fpga_GAME_count_speed1_a1[23] ));
 sg13g2_nand2b_1 _4621_ (.Y(_1141_),
    .B(net1671),
    .A_N(\FpgaPins_Fpga_GAME_win_a2[2] ));
 sg13g2_nor2_1 _4622_ (.A(_0791_),
    .B(_1141_),
    .Y(_1142_));
 sg13g2_o21ai_1 _4623_ (.B1(_0783_),
    .Y(_1143_),
    .A1(net983),
    .A2(_0718_));
 sg13g2_a21oi_1 _4624_ (.A1(net983),
    .A2(\FpgaPins_Fpga_GAME_led_output_a2[0] ),
    .Y(_1144_),
    .B1(_1143_));
 sg13g2_o21ai_1 _4625_ (.B1(_0786_),
    .Y(_1145_),
    .A1(\FpgaPins_Fpga_GAME_led_output_a2[1] ),
    .A2(_0783_));
 sg13g2_nand2_1 _4626_ (.Y(_1146_),
    .A(\FpgaPins_Fpga_GAME_score_a4[1] ),
    .B(net978));
 sg13g2_o21ai_1 _4627_ (.B1(_1146_),
    .Y(_1147_),
    .A1(_1144_),
    .A2(_1145_));
 sg13g2_and2_1 _4628_ (.A(_1142_),
    .B(_1147_),
    .X(_1148_));
 sg13g2_nand2_2 _4629_ (.Y(_1149_),
    .A(net1589),
    .B(net1669));
 sg13g2_nand2b_2 _4630_ (.Y(\FpgaPins_Fpga_GAME_led_output_a1[1] ),
    .B(_1149_),
    .A_N(_1148_));
 sg13g2_a21oi_1 _4631_ (.A1(\FpgaPins_Fpga_GAME_led_output_a2[6] ),
    .A2(net980),
    .Y(_1150_),
    .B1(net979));
 sg13g2_nand2b_1 _4632_ (.Y(_1151_),
    .B(net984),
    .A_N(\FpgaPins_Fpga_GAME_led_output_a2[5] ));
 sg13g2_o21ai_1 _4633_ (.B1(_1151_),
    .Y(_1152_),
    .A1(FpgaPins_Fpga_GAME_forward_a2),
    .A2(\FpgaPins_Fpga_GAME_led_output_a2[7] ));
 sg13g2_o21ai_1 _4634_ (.B1(_1150_),
    .Y(_1153_),
    .A1(net980),
    .A2(_1152_));
 sg13g2_a21oi_1 _4635_ (.A1(_0719_),
    .A2(net979),
    .Y(_1154_),
    .B1(_0791_));
 sg13g2_a21oi_1 _4636_ (.A1(_1153_),
    .A2(_1154_),
    .Y(_1155_),
    .B1(net1636));
 sg13g2_nor2_1 _4637_ (.A(_0782_),
    .B(_1155_),
    .Y(\FpgaPins_Fpga_GAME_led_output_a1[6] ));
 sg13g2_nand2b_1 _4638_ (.Y(_1156_),
    .B(\FpgaPins_Fpga_GAME_led_output_a2[1] ),
    .A_N(net983));
 sg13g2_o21ai_1 _4639_ (.B1(_0786_),
    .Y(_1157_),
    .A1(\FpgaPins_Fpga_GAME_led_output_a2[0] ),
    .A2(_0783_));
 sg13g2_a21oi_1 _4640_ (.A1(_0783_),
    .A2(_1156_),
    .Y(_1158_),
    .B1(_1157_));
 sg13g2_a21oi_1 _4641_ (.A1(net1725),
    .A2(net978),
    .Y(_1159_),
    .B1(_1158_));
 sg13g2_nor2b_1 _4642_ (.A(_1159_),
    .B_N(_1142_),
    .Y(_1160_));
 sg13g2_a21oi_2 _4643_ (.B1(_1160_),
    .Y(_1161_),
    .A2(net1669),
    .A1(net1589));
 sg13g2_inv_1 _4644_ (.Y(\FpgaPins_Fpga_GAME_led_output_a1[0] ),
    .A(_1161_));
 sg13g2_or2_1 _4645_ (.X(_1162_),
    .B(\FpgaPins_Fpga_GAME_led_output_a2[4] ),
    .A(net984));
 sg13g2_a21oi_1 _4646_ (.A1(net983),
    .A2(_0718_),
    .Y(_1163_),
    .B1(net980));
 sg13g2_a22oi_1 _4647_ (.Y(_1164_),
    .B1(_1162_),
    .B2(_1163_),
    .A2(net980),
    .A1(\FpgaPins_Fpga_GAME_led_output_a2[3] ));
 sg13g2_nand2_1 _4648_ (.Y(_1165_),
    .A(\FpgaPins_Fpga_GAME_score_a4[3] ),
    .B(net979));
 sg13g2_o21ai_1 _4649_ (.B1(_1165_),
    .Y(_1166_),
    .A1(net978),
    .A2(_1164_));
 sg13g2_nor2_1 _4650_ (.A(_0791_),
    .B(_1166_),
    .Y(_1167_));
 sg13g2_o21ai_1 _4651_ (.B1(_1149_),
    .Y(\FpgaPins_Fpga_GAME_led_output_a1[3] ),
    .A1(_1141_),
    .A2(_1167_));
 sg13g2_a21oi_1 _4652_ (.A1(net984),
    .A2(_0721_),
    .Y(_1168_),
    .B1(net980));
 sg13g2_o21ai_1 _4653_ (.B1(_1168_),
    .Y(_1169_),
    .A1(net983),
    .A2(\FpgaPins_Fpga_GAME_led_output_a2[5] ));
 sg13g2_a21oi_1 _4654_ (.A1(\FpgaPins_Fpga_GAME_led_output_a2[4] ),
    .A2(net980),
    .Y(_1170_),
    .B1(net978));
 sg13g2_nand2b_1 _4655_ (.Y(_1171_),
    .B(net978),
    .A_N(\FpgaPins_Fpga_GAME_score_a4[4] ));
 sg13g2_a21oi_1 _4656_ (.A1(_1169_),
    .A2(_1170_),
    .Y(_1172_),
    .B1(_0791_));
 sg13g2_a21oi_2 _4657_ (.B1(net1636),
    .Y(_1173_),
    .A2(_1172_),
    .A1(_1171_));
 sg13g2_nor2_2 _4658_ (.A(_0782_),
    .B(_1173_),
    .Y(\FpgaPins_Fpga_GAME_led_output_a1[4] ));
 sg13g2_a21oi_1 _4659_ (.A1(net983),
    .A2(_0720_),
    .Y(_1174_),
    .B1(net980));
 sg13g2_o21ai_1 _4660_ (.B1(_1174_),
    .Y(_1175_),
    .A1(net984),
    .A2(\FpgaPins_Fpga_GAME_led_output_a2[6] ));
 sg13g2_a21oi_1 _4661_ (.A1(\FpgaPins_Fpga_GAME_led_output_a2[5] ),
    .A2(net980),
    .Y(_1176_),
    .B1(net978));
 sg13g2_nand2b_1 _4662_ (.Y(_1177_),
    .B(net978),
    .A_N(net1691));
 sg13g2_a21oi_1 _4663_ (.A1(_1175_),
    .A2(_1176_),
    .Y(_1178_),
    .B1(_0791_));
 sg13g2_a21oi_2 _4664_ (.B1(net1636),
    .Y(_1179_),
    .A2(_1178_),
    .A1(_1177_));
 sg13g2_nor2_1 _4665_ (.A(_0782_),
    .B(_1179_),
    .Y(\FpgaPins_Fpga_GAME_led_output_a1[5] ));
 sg13g2_o21ai_1 _4666_ (.B1(_0783_),
    .Y(_1180_),
    .A1(net983),
    .A2(_0721_));
 sg13g2_a21oi_1 _4667_ (.A1(net983),
    .A2(\FpgaPins_Fpga_GAME_led_output_a2[1] ),
    .Y(_1181_),
    .B1(_1180_));
 sg13g2_o21ai_1 _4668_ (.B1(_0786_),
    .Y(_1182_),
    .A1(\FpgaPins_Fpga_GAME_led_output_a2[2] ),
    .A2(_0783_));
 sg13g2_nand2_1 _4669_ (.Y(_1183_),
    .A(\FpgaPins_Fpga_GAME_score_a4[2] ),
    .B(net978));
 sg13g2_o21ai_1 _4670_ (.B1(_1183_),
    .Y(_1184_),
    .A1(_1181_),
    .A2(_1182_));
 sg13g2_nand2_1 _4671_ (.Y(_1185_),
    .A(_1142_),
    .B(_1184_));
 sg13g2_nand2_2 _4672_ (.Y(\FpgaPins_Fpga_GAME_led_output_a1[2] ),
    .A(_1149_),
    .B(_1185_));
 sg13g2_and2_1 _4673_ (.A(net8),
    .B(net2),
    .X(_1186_));
 sg13g2_and2_1 _4674_ (.A(net1),
    .B(net996),
    .X(_1187_));
 sg13g2_nand2_1 _4675_ (.Y(_1188_),
    .A(net1),
    .B(net996));
 sg13g2_nor3_2 _4676_ (.A(net3),
    .B(net4),
    .C(net5),
    .Y(_1189_));
 sg13g2_or3_2 _4677_ (.A(net3),
    .B(net4),
    .C(net5),
    .X(_1190_));
 sg13g2_o21ai_1 _4678_ (.B1(_1189_),
    .Y(_1191_),
    .A1(net1359),
    .A2(net1424));
 sg13g2_nand2_1 _4679_ (.Y(_1192_),
    .A(net1457),
    .B(_1191_));
 sg13g2_nand3_1 _4680_ (.B(net1457),
    .C(_1191_),
    .A(\C1.next_state_var[4] ),
    .Y(_1193_));
 sg13g2_nand2_1 _4681_ (.Y(_1194_),
    .A(\C1.next_state_var[4] ),
    .B(_1190_));
 sg13g2_a21oi_1 _4682_ (.A1(\C1.next_state_var[4] ),
    .A2(_1190_),
    .Y(_1195_),
    .B1(net1001));
 sg13g2_a21oi_1 _4683_ (.A1(net1458),
    .A2(_1195_),
    .Y(_0007_),
    .B1(net968));
 sg13g2_nor4_2 _4684_ (.A(\FpgaPins_Fpga_GAME_led_output_a2[1] ),
    .B(\FpgaPins_Fpga_GAME_led_output_a2[5] ),
    .C(\FpgaPins_Fpga_GAME_led_output_a2[4] ),
    .Y(_1196_),
    .D(\FpgaPins_Fpga_GAME_led_output_a2[3] ));
 sg13g2_nor4_2 _4685_ (.A(\FpgaPins_Fpga_GAME_led_output_a2[6] ),
    .B(\FpgaPins_Fpga_GAME_led_output_a2[7] ),
    .C(\FpgaPins_Fpga_GAME_led_output_a2[2] ),
    .Y(_1197_),
    .D(\FpgaPins_Fpga_GAME_led_output_a2[0] ));
 sg13g2_nor2_1 _4686_ (.A(\FpgaPins_Fpga_GAME_led_output_a3[1] ),
    .B(\FpgaPins_Fpga_GAME_led_output_a3[3] ),
    .Y(_1198_));
 sg13g2_nor4_1 _4687_ (.A(\FpgaPins_Fpga_GAME_led_output_a3[2] ),
    .B(\FpgaPins_Fpga_GAME_led_output_a3[5] ),
    .C(\FpgaPins_Fpga_GAME_led_output_a3[4] ),
    .D(\FpgaPins_Fpga_GAME_led_output_a3[6] ),
    .Y(_1199_));
 sg13g2_and4_2 _4688_ (.A(_1196_),
    .B(_1197_),
    .C(_1198_),
    .D(_1199_),
    .X(_1200_));
 sg13g2_nand3b_1 _4689_ (.B(_1200_),
    .C(\FpgaPins_Fpga_GAME_led_output_a3[0] ),
    .Y(_1201_),
    .A_N(\FpgaPins_Fpga_GAME_led_output_a3[7] ));
 sg13g2_inv_1 _4690_ (.Y(_1202_),
    .A(_1201_));
 sg13g2_or4_1 _4691_ (.A(\FpgaPins_Fpga_GAME_score_a2[5] ),
    .B(\FpgaPins_Fpga_GAME_score_a2[4] ),
    .C(\FpgaPins_Fpga_GAME_score_a2[3] ),
    .D(\FpgaPins_Fpga_GAME_score_a2[2] ),
    .X(_1203_));
 sg13g2_nor4_1 _4692_ (.A(\FpgaPins_Fpga_GAME_score_a2[7] ),
    .B(\FpgaPins_Fpga_GAME_score_a2[6] ),
    .C(net1581),
    .D(_1203_),
    .Y(_1204_));
 sg13g2_nand2_1 _4693_ (.Y(_1205_),
    .A(\FpgaPins_Fpga_GAME_led_output_a3[0] ),
    .B(_1200_));
 sg13g2_nor2_1 _4694_ (.A(net1571),
    .B(_1205_),
    .Y(_1206_));
 sg13g2_and3_1 _4695_ (.X(_1207_),
    .A(net720),
    .B(_1204_),
    .C(_1206_));
 sg13g2_nor2b_1 _4696_ (.A(_1207_),
    .B_N(net1589),
    .Y(_1208_));
 sg13g2_nand3b_1 _4697_ (.B(_0683_),
    .C(net714),
    .Y(_1209_),
    .A_N(\FpgaPins_Fpga_GAME_score_a2[6] ));
 sg13g2_nand2_1 _4698_ (.Y(_1210_),
    .A(net1571),
    .B(_1200_));
 sg13g2_nor2_2 _4699_ (.A(net1562),
    .B(_1210_),
    .Y(_1211_));
 sg13g2_or2_2 _4700_ (.X(_1212_),
    .B(_1210_),
    .A(\FpgaPins_Fpga_GAME_led_output_a3[0] ));
 sg13g2_nor4_1 _4701_ (.A(net720),
    .B(_1203_),
    .C(_1209_),
    .D(_1212_),
    .Y(_1213_));
 sg13g2_nor2_1 _4702_ (.A(_1208_),
    .B(_1213_),
    .Y(_1214_));
 sg13g2_nor2_1 _4703_ (.A(net1492),
    .B(net1590),
    .Y(\FpgaPins_Fpga_GAME_win_a1[0] ));
 sg13g2_nor2_1 _4704_ (.A(net1636),
    .B(_1207_),
    .Y(_1215_));
 sg13g2_nor3_1 _4705_ (.A(net1492),
    .B(_1213_),
    .C(_1215_),
    .Y(\FpgaPins_Fpga_GAME_win_a1[1] ));
 sg13g2_nor3_1 _4706_ (.A(_0677_),
    .B(net994),
    .C(net1747),
    .Y(_1216_));
 sg13g2_nand2b_1 _4707_ (.Y(_0000_),
    .B(net970),
    .A_N(_1216_));
 sg13g2_nand2_2 _4708_ (.Y(_1217_),
    .A(_0669_),
    .B(_0670_));
 sg13g2_a21oi_1 _4709_ (.A1(_1189_),
    .A2(_1217_),
    .Y(_1218_),
    .B1(net1546));
 sg13g2_nor2_2 _4710_ (.A(net1001),
    .B(net968),
    .Y(_1219_));
 sg13g2_nand2_2 _4711_ (.Y(_1220_),
    .A(_0722_),
    .B(net971));
 sg13g2_nor2_1 _4712_ (.A(_1189_),
    .B(_1220_),
    .Y(_1221_));
 sg13g2_nand2_1 _4713_ (.Y(_1222_),
    .A(net1546),
    .B(_1221_));
 sg13g2_nor2_1 _4714_ (.A(_1190_),
    .B(_1220_),
    .Y(_1223_));
 sg13g2_nand2_1 _4715_ (.Y(_1224_),
    .A(_0675_),
    .B(_0676_));
 sg13g2_a21oi_1 _4716_ (.A1(_1189_),
    .A2(_1224_),
    .Y(_1225_),
    .B1(net995));
 sg13g2_and2_1 _4717_ (.A(net1546),
    .B(_1225_),
    .X(_1226_));
 sg13g2_o21ai_1 _4718_ (.B1(_1223_),
    .Y(_1227_),
    .A1(\C1.next_state_var[6] ),
    .A2(_1226_));
 sg13g2_o21ai_1 _4719_ (.B1(_1222_),
    .Y(_0004_),
    .A1(_1218_),
    .A2(_1227_));
 sg13g2_nand3_1 _4720_ (.B(\C1.counter_status[1] ),
    .C(_1219_),
    .A(net1179),
    .Y(_1228_));
 sg13g2_a21oi_1 _4721_ (.A1(\C1.next_state_var[0] ),
    .A2(net997),
    .Y(_1229_),
    .B1(net968));
 sg13g2_nand2_1 _4722_ (.Y(_0003_),
    .A(net1180),
    .B(_1229_));
 sg13g2_nor2_1 _4723_ (.A(net997),
    .B(net1728),
    .Y(_1230_));
 sg13g2_a21oi_1 _4724_ (.A1(_1173_),
    .A2(_1179_),
    .Y(_1231_),
    .B1(_0782_));
 sg13g2_a21oi_1 _4725_ (.A1(_0793_),
    .A2(_1155_),
    .Y(_1232_),
    .B1(_0782_));
 sg13g2_or2_1 _4726_ (.X(_1233_),
    .B(_1232_),
    .A(_1231_));
 sg13g2_nor4_1 _4727_ (.A(net997),
    .B(FpgaPins_Fpga_GAME_right_btn_a2),
    .C(\FpgaPins_Fpga_GAME_led_output_a1[3] ),
    .D(_1233_),
    .Y(_1234_));
 sg13g2_nor2b_1 _4728_ (.A(\FpgaPins_Fpga_GAME_led_output_a1[2] ),
    .B_N(_1234_),
    .Y(_1235_));
 sg13g2_nand3b_1 _4729_ (.B(_1160_),
    .C(_1235_),
    .Y(_1236_),
    .A_N(\FpgaPins_Fpga_GAME_led_output_a1[1] ));
 sg13g2_nand2b_1 _4730_ (.Y(_1237_),
    .B(_1161_),
    .A_N(_1148_));
 sg13g2_nand2b_1 _4731_ (.Y(_1238_),
    .B(_1185_),
    .A_N(_1237_));
 sg13g2_nand2b_1 _4732_ (.Y(_1239_),
    .B(net4),
    .A_N(FpgaPins_Fpga_GAME_left_btn_a2));
 sg13g2_nor3_1 _4733_ (.A(\FpgaPins_Fpga_GAME_led_output_a1[3] ),
    .B(_1238_),
    .C(_1239_),
    .Y(_1240_));
 sg13g2_nor2b_1 _4734_ (.A(_1231_),
    .B_N(_1240_),
    .Y(_1241_));
 sg13g2_nand3_1 _4735_ (.B(_1155_),
    .C(_1241_),
    .A(\FpgaPins_Fpga_GAME_led_output_a1[7] ),
    .Y(_1242_));
 sg13g2_nand2_1 _4736_ (.Y(_1243_),
    .A(_1236_),
    .B(_1242_));
 sg13g2_nor2_1 _4737_ (.A(_1185_),
    .B(_1237_),
    .Y(_1244_));
 sg13g2_nor2b_1 _4738_ (.A(_1232_),
    .B_N(_1240_),
    .Y(_1245_));
 sg13g2_and2_1 _4739_ (.A(_1173_),
    .B(\FpgaPins_Fpga_GAME_led_output_a1[5] ),
    .X(_1246_));
 sg13g2_a22oi_1 _4740_ (.Y(_1247_),
    .B1(_1245_),
    .B2(_1246_),
    .A2(_1244_),
    .A1(_1234_));
 sg13g2_nand3_1 _4741_ (.B(\FpgaPins_Fpga_GAME_led_output_a1[6] ),
    .C(_1241_),
    .A(_0793_),
    .Y(_1248_));
 sg13g2_nand3_1 _4742_ (.B(_1161_),
    .C(_1235_),
    .A(_1148_),
    .Y(_1249_));
 sg13g2_nand2_1 _4743_ (.Y(_1250_),
    .A(_1248_),
    .B(_1249_));
 sg13g2_nand3_1 _4744_ (.B(_1179_),
    .C(_1245_),
    .A(\FpgaPins_Fpga_GAME_led_output_a1[4] ),
    .Y(_1251_));
 sg13g2_nor2_1 _4745_ (.A(_1233_),
    .B(_1238_),
    .Y(_1252_));
 sg13g2_nand3_1 _4746_ (.B(_1230_),
    .C(_1252_),
    .A(\FpgaPins_Fpga_GAME_led_output_a1[3] ),
    .Y(_1253_));
 sg13g2_nand4_1 _4747_ (.B(_0790_),
    .C(_1251_),
    .A(net985),
    .Y(_1254_),
    .D(_1253_));
 sg13g2_nor3_1 _4748_ (.A(_1243_),
    .B(_1250_),
    .C(_1254_),
    .Y(_1255_));
 sg13g2_and3_1 _4749_ (.X(_1256_),
    .A(net1686),
    .B(_1247_),
    .C(_1255_));
 sg13g2_or2_1 _4750_ (.X(_0013_),
    .B(_1256_),
    .A(_1243_));
 sg13g2_inv_1 _4751_ (.Y(_1257_),
    .A(_0013_));
 sg13g2_nand2_1 _4752_ (.Y(_1258_),
    .A(net1578),
    .B(_1255_));
 sg13g2_nand2_1 _4753_ (.Y(_0012_),
    .A(_1247_),
    .B(_1258_));
 sg13g2_and3_1 _4754_ (.X(_1259_),
    .A(net1720),
    .B(_1247_),
    .C(_1255_));
 sg13g2_or2_1 _4755_ (.X(_0011_),
    .B(_1259_),
    .A(_1250_));
 sg13g2_nand2b_1 _4756_ (.Y(_1260_),
    .B(net992),
    .A_N(net1532));
 sg13g2_nand2_1 _4757_ (.Y(_1261_),
    .A(net1594),
    .B(net1532));
 sg13g2_nor2_1 _4758_ (.A(net1532),
    .B(_1220_),
    .Y(_1262_));
 sg13g2_a21oi_1 _4759_ (.A1(_1260_),
    .A2(_1261_),
    .Y(_0010_),
    .B1(_1220_));
 sg13g2_a21o_1 _4760_ (.A2(_1218_),
    .A1(net993),
    .B1(net1692),
    .X(_1263_));
 sg13g2_nor2_2 _4761_ (.A(\C1.temp[1] ),
    .B(\C1.temp[0] ),
    .Y(_1264_));
 sg13g2_nor2_1 _4762_ (.A(_1190_),
    .B(_1264_),
    .Y(_1265_));
 sg13g2_nor2_1 _4763_ (.A(net993),
    .B(_1265_),
    .Y(_1266_));
 sg13g2_a22oi_1 _4764_ (.Y(_1267_),
    .B1(_1223_),
    .B2(_1263_),
    .A2(_1221_),
    .A1(net993));
 sg13g2_nor2_1 _4765_ (.A(_1266_),
    .B(_1267_),
    .Y(_0009_));
 sg13g2_nor2_1 _4766_ (.A(_0724_),
    .B(_1190_),
    .Y(_1268_));
 sg13g2_a22oi_1 _4767_ (.Y(_1269_),
    .B1(_1268_),
    .B2(_1219_),
    .A2(_1262_),
    .A1(net995));
 sg13g2_nor2_1 _4768_ (.A(_1225_),
    .B(_1269_),
    .Y(_0008_));
 sg13g2_nand3_1 _4769_ (.B(net1532),
    .C(_1219_),
    .A(net995),
    .Y(_1270_));
 sg13g2_nand2_1 _4770_ (.Y(_1271_),
    .A(\C1.next_state_var[3] ),
    .B(_1262_));
 sg13g2_nand2_1 _4771_ (.Y(_0006_),
    .A(net1533),
    .B(_1271_));
 sg13g2_a22oi_1 _4772_ (.Y(_1272_),
    .B1(_1266_),
    .B2(net1692),
    .A2(_1192_),
    .A1(\C1.next_state_var[4] ));
 sg13g2_nor2b_1 _4773_ (.A(_1272_),
    .B_N(_1223_),
    .Y(_1273_));
 sg13g2_a21o_1 _4774_ (.A2(_1221_),
    .A1(net1692),
    .B1(_1273_),
    .X(_0005_));
 sg13g2_a22oi_1 _4775_ (.Y(_1274_),
    .B1(_0858_),
    .B2(_0866_),
    .A2(_0849_),
    .A1(_0841_));
 sg13g2_nand2_1 _4776_ (.Y(_1275_),
    .A(_0850_),
    .B(net859));
 sg13g2_nor2_2 _4777_ (.A(net1731),
    .B(net947),
    .Y(_1276_));
 sg13g2_nand2b_1 _4778_ (.Y(_1277_),
    .B(net977),
    .A_N(net1757));
 sg13g2_a221oi_1 _4779_ (.B2(net896),
    .C1(_1084_),
    .B1(_1092_),
    .A1(_1068_),
    .Y(_1278_),
    .A2(_1076_));
 sg13g2_nand2_1 _4780_ (.Y(_1279_),
    .A(_1276_),
    .B(_1278_));
 sg13g2_nor4_2 _4781_ (.A(_1002_),
    .B(_1010_),
    .C(_1051_),
    .Y(_1280_),
    .D(_1059_));
 sg13g2_nand3_1 _4782_ (.B(_1278_),
    .C(_1280_),
    .A(_1276_),
    .Y(_1281_));
 sg13g2_nand4_1 _4783_ (.B(_1276_),
    .C(_1278_),
    .A(_1274_),
    .Y(_1282_),
    .D(_1280_));
 sg13g2_inv_1 _4784_ (.Y(FpgaPins_Fpga_LIPSI_is_ret_a1),
    .A(_1282_));
 sg13g2_nor2_1 _4785_ (.A(\FpgaPins_Fpga_FSM_instr_a1[6] ),
    .B(_1277_),
    .Y(_1283_));
 sg13g2_nand2_1 _4786_ (.Y(_1284_),
    .A(\FpgaPins_Fpga_FSM_instr_a1[7] ),
    .B(_1283_));
 sg13g2_nand3_1 _4787_ (.B(_1280_),
    .C(_1283_),
    .A(\FpgaPins_Fpga_FSM_instr_a1[7] ),
    .Y(_1285_));
 sg13g2_inv_1 _4788_ (.Y(FpgaPins_Fpga_LIPSI_is_brl_a1),
    .A(net822));
 sg13g2_nand3_1 _4789_ (.B(\FpgaPins_Fpga_FSM_instr_a1[7] ),
    .C(_1283_),
    .A(\FpgaPins_Fpga_FSM_instr_a1[5] ),
    .Y(_1286_));
 sg13g2_nor2_1 _4790_ (.A(\FpgaPins_Fpga_FSM_instr_a1[4] ),
    .B(_1286_),
    .Y(FpgaPins_Fpga_LIPSI_is_ld_ind_a1));
 sg13g2_nor2_1 _4791_ (.A(_1060_),
    .B(_1286_),
    .Y(FpgaPins_Fpga_LIPSI_is_st_ind_a1));
 sg13g2_nand3_1 _4792_ (.B(_1076_),
    .C(_1276_),
    .A(_1068_),
    .Y(_1287_));
 sg13g2_nand2_1 _4793_ (.Y(_1288_),
    .A(_0024_),
    .B(_1287_));
 sg13g2_o21ai_1 _4794_ (.B1(_1288_),
    .Y(_1289_),
    .A1(net875),
    .A2(_1287_));
 sg13g2_inv_1 _4795_ (.Y(_1290_),
    .A(_1289_));
 sg13g2_nand2_1 _4796_ (.Y(_1291_),
    .A(_0021_),
    .B(_1287_));
 sg13g2_o21ai_1 _4797_ (.B1(_1291_),
    .Y(_1292_),
    .A1(\FpgaPins_Fpga_FSM_instr_a1[4] ),
    .A2(_1287_));
 sg13g2_nor2_2 _4798_ (.A(_1289_),
    .B(_1292_),
    .Y(_1293_));
 sg13g2_and2_2 _4799_ (.A(net981),
    .B(_1287_),
    .X(_1294_));
 sg13g2_nand2_1 _4800_ (.Y(_1295_),
    .A(_0027_),
    .B(_1287_));
 sg13g2_o21ai_1 _4801_ (.B1(_1295_),
    .Y(_1296_),
    .A1(\FpgaPins_Fpga_FSM_instr_a1[6] ),
    .A2(_1287_));
 sg13g2_nor2_2 _4802_ (.A(_1294_),
    .B(_1296_),
    .Y(_1297_));
 sg13g2_and2_1 _4803_ (.A(_1293_),
    .B(_1297_),
    .X(_1298_));
 sg13g2_nand2_2 _4804_ (.Y(_1299_),
    .A(_1293_),
    .B(_1297_));
 sg13g2_mux2_1 _4805_ (.A0(_0106_),
    .A1(_0107_),
    .S(_0797_),
    .X(_1300_));
 sg13g2_nand2b_2 _4806_ (.Y(_1301_),
    .B(_1276_),
    .A_N(_1278_));
 sg13g2_nor2_1 _4807_ (.A(_1277_),
    .B(_1278_),
    .Y(_1302_));
 sg13g2_mux2_1 _4808_ (.A0(_1026_),
    .A1(_1300_),
    .S(_1282_),
    .X(_1303_));
 sg13g2_o21ai_1 _4809_ (.B1(net977),
    .Y(_1304_),
    .A1(\FpgaPins_Fpga_FSM_instr_a1[1] ),
    .A2(_1301_));
 sg13g2_a21oi_2 _4810_ (.B1(_1304_),
    .Y(\FpgaPins_Fpga_FSM_idata_rd_addr_a1[1] ),
    .A2(_1303_),
    .A1(_1301_));
 sg13g2_nand2b_1 _4811_ (.Y(_1305_),
    .B(_0797_),
    .A_N(_0105_));
 sg13g2_o21ai_1 _4812_ (.B1(_1305_),
    .Y(_1306_),
    .A1(_0104_),
    .A2(_0797_));
 sg13g2_or2_1 _4813_ (.X(_1307_),
    .B(_1282_),
    .A(_1043_));
 sg13g2_a21oi_1 _4814_ (.A1(_1282_),
    .A2(_1306_),
    .Y(_1308_),
    .B1(_1302_));
 sg13g2_o21ai_1 _4815_ (.B1(net977),
    .Y(_1309_),
    .A1(net859),
    .A2(_1301_));
 sg13g2_a21o_1 _4816_ (.A2(_1308_),
    .A1(_1307_),
    .B1(_1309_),
    .X(_1310_));
 sg13g2_inv_1 _4817_ (.Y(\FpgaPins_Fpga_FSM_idata_rd_addr_a1[0] ),
    .A(net809));
 sg13g2_mux2_1 _4818_ (.A0(_0121_),
    .A1(_0120_),
    .S(net810),
    .X(_1311_));
 sg13g2_nand2b_1 _4819_ (.Y(_1312_),
    .B(_0797_),
    .A_N(\FpgaPins_Fpga_LIPSI_dptr_a2[2] ));
 sg13g2_o21ai_1 _4820_ (.B1(_1312_),
    .Y(_1313_),
    .A1(\FpgaPins_Fpga_LIPSI_data_a2[2] ),
    .A2(_0797_));
 sg13g2_nand3_1 _4821_ (.B(_1301_),
    .C(_1313_),
    .A(_1282_),
    .Y(_1314_));
 sg13g2_nand2_1 _4822_ (.Y(_1315_),
    .A(_1043_),
    .B(_1302_));
 sg13g2_nand3_1 _4823_ (.B(_1314_),
    .C(_1315_),
    .A(net977),
    .Y(_1316_));
 sg13g2_inv_1 _4824_ (.Y(\FpgaPins_Fpga_FSM_idata_rd_addr_a1[2] ),
    .A(net803));
 sg13g2_a21oi_1 _4825_ (.A1(_0730_),
    .A2(net798),
    .Y(_1317_),
    .B1(net818));
 sg13g2_o21ai_1 _4826_ (.B1(_1317_),
    .Y(_1318_),
    .A1(net1640),
    .A2(net798));
 sg13g2_a21oi_1 _4827_ (.A1(net818),
    .A2(_1311_),
    .Y(_1319_),
    .B1(_1316_));
 sg13g2_mux4_1 _4828_ (.S0(net804),
    .A0(_0115_),
    .A1(_0114_),
    .A2(_0117_),
    .A3(_0116_),
    .S1(net813),
    .X(_1320_));
 sg13g2_nand2b_1 _4829_ (.Y(_1321_),
    .B(_0797_),
    .A_N(\FpgaPins_Fpga_LIPSI_dptr_a2[3] ));
 sg13g2_o21ai_1 _4830_ (.B1(_1321_),
    .Y(_1322_),
    .A1(\FpgaPins_Fpga_LIPSI_data_a2[3] ),
    .A2(_0797_));
 sg13g2_nand3_1 _4831_ (.B(_1301_),
    .C(_1322_),
    .A(_1282_),
    .Y(_1323_));
 sg13g2_nand2_1 _4832_ (.Y(_1324_),
    .A(_1026_),
    .B(_1302_));
 sg13g2_nand3_1 _4833_ (.B(_1323_),
    .C(_1324_),
    .A(net977),
    .Y(_1325_));
 sg13g2_inv_1 _4834_ (.Y(\FpgaPins_Fpga_FSM_idata_rd_addr_a1[3] ),
    .A(_1325_));
 sg13g2_o21ai_1 _4835_ (.B1(\FpgaPins_Fpga_FSM_idata_rd_addr_a1[3] ),
    .Y(_1326_),
    .A1(net797),
    .A2(_1320_));
 sg13g2_a21oi_2 _4836_ (.B1(_1326_),
    .Y(_1327_),
    .A2(_1319_),
    .A1(net1641));
 sg13g2_a21oi_1 _4837_ (.A1(_0729_),
    .A2(net807),
    .Y(_1328_),
    .B1(net815));
 sg13g2_o21ai_1 _4838_ (.B1(_1328_),
    .Y(_1329_),
    .A1(_0111_),
    .A2(net807));
 sg13g2_mux2_1 _4839_ (.A0(_0113_),
    .A1(_0112_),
    .S(net809),
    .X(_1330_));
 sg13g2_a21oi_1 _4840_ (.A1(net816),
    .A2(_1330_),
    .Y(_1331_),
    .B1(net802));
 sg13g2_mux4_1 _4841_ (.S0(net805),
    .A0(_0103_),
    .A1(_0102_),
    .A2(_0109_),
    .A3(_0108_),
    .S1(net814),
    .X(_1332_));
 sg13g2_o21ai_1 _4842_ (.B1(_1325_),
    .Y(_1333_),
    .A1(net796),
    .A2(_1332_));
 sg13g2_a21oi_2 _4843_ (.B1(_1333_),
    .Y(_1334_),
    .A2(_1331_),
    .A1(_1329_));
 sg13g2_nor2_1 _4844_ (.A(net1642),
    .B(_1334_),
    .Y(\FpgaPins_Fpga_FSM_data_a1[0] ));
 sg13g2_nor3_1 _4845_ (.A(_0699_),
    .B(_1327_),
    .C(_1334_),
    .Y(_1335_));
 sg13g2_nor2_1 _4846_ (.A(\FpgaPins_Fpga_FSM_instr_a1[4] ),
    .B(_1279_),
    .Y(_1336_));
 sg13g2_nand2_2 _4847_ (.Y(_1337_),
    .A(\FpgaPins_Fpga_FSM_instr_a1[1] ),
    .B(\FpgaPins_Fpga_FSM_instr_a1[0] ));
 sg13g2_nand2_2 _4848_ (.Y(_1338_),
    .A(net875),
    .B(_1336_));
 sg13g2_nor2_1 _4849_ (.A(_1337_),
    .B(_1338_),
    .Y(_1339_));
 sg13g2_or2_2 _4850_ (.X(_1340_),
    .B(_1338_),
    .A(_1337_));
 sg13g2_o21ai_1 _4851_ (.B1(_1340_),
    .Y(_1341_),
    .A1(_0022_),
    .A2(net988));
 sg13g2_nor2_1 _4852_ (.A(net859),
    .B(_1338_),
    .Y(_1342_));
 sg13g2_nor3_1 _4853_ (.A(_0850_),
    .B(net859),
    .C(_1338_),
    .Y(_1343_));
 sg13g2_nor3_1 _4854_ (.A(_0850_),
    .B(net859),
    .C(_1338_),
    .Y(_1344_));
 sg13g2_a21oi_1 _4855_ (.A1(_0025_),
    .A2(net793),
    .Y(_1345_),
    .B1(net792));
 sg13g2_o21ai_1 _4856_ (.B1(_1345_),
    .Y(_1346_),
    .A1(_1335_),
    .A2(_1341_));
 sg13g2_nor2_2 _4857_ (.A(\FpgaPins_Fpga_FSM_instr_a1[1] ),
    .B(_1338_),
    .Y(_1347_));
 sg13g2_nand3_1 _4858_ (.B(net875),
    .C(_1336_),
    .A(_0850_),
    .Y(_1348_));
 sg13g2_nand2b_1 _4859_ (.Y(_1349_),
    .B(net792),
    .A_N(_0123_));
 sg13g2_nand3_1 _4860_ (.B(_1348_),
    .C(_1349_),
    .A(_1346_),
    .Y(_1350_));
 sg13g2_nor2_1 _4861_ (.A(net859),
    .B(_1348_),
    .Y(_1351_));
 sg13g2_nor2_2 _4862_ (.A(_0867_),
    .B(_1348_),
    .Y(_1352_));
 sg13g2_a22oi_1 _4863_ (.Y(_1353_),
    .B1(_1352_),
    .B2(_0025_),
    .A2(_1351_),
    .A1(_0122_));
 sg13g2_nor2_1 _4864_ (.A(_1275_),
    .B(_1338_),
    .Y(_1354_));
 sg13g2_a21oi_1 _4865_ (.A1(_1350_),
    .A2(_1353_),
    .Y(_1355_),
    .B1(net800));
 sg13g2_nor2_2 _4866_ (.A(_1290_),
    .B(_1292_),
    .Y(_1356_));
 sg13g2_and2_1 _4867_ (.A(_1297_),
    .B(_1356_),
    .X(_1357_));
 sg13g2_nor2b_2 _4868_ (.A(_1289_),
    .B_N(_1292_),
    .Y(_1358_));
 sg13g2_and2_1 _4869_ (.A(_1297_),
    .B(_1358_),
    .X(_1359_));
 sg13g2_nor2_2 _4870_ (.A(net781),
    .B(net790),
    .Y(_1360_));
 sg13g2_o21ai_1 _4871_ (.B1(net981),
    .Y(_1361_),
    .A1(_1327_),
    .A2(_1334_));
 sg13g2_nand2_1 _4872_ (.Y(_1362_),
    .A(FpgaPins_Fpga_LIPSI_is_ALU_imm_a2),
    .B(_0867_));
 sg13g2_and2_2 _4873_ (.A(_1361_),
    .B(_1362_),
    .X(_1363_));
 sg13g2_o21ai_1 _4874_ (.B1(_1360_),
    .Y(_1364_),
    .A1(_1299_),
    .A2(_1363_));
 sg13g2_and2_1 _4875_ (.A(_1289_),
    .B(_1292_),
    .X(_1365_));
 sg13g2_and2_1 _4876_ (.A(_1297_),
    .B(_1365_),
    .X(_1366_));
 sg13g2_or2_1 _4877_ (.X(_1367_),
    .B(_1363_),
    .A(\FpgaPins_Fpga_LIPSI_acc_a2[0] ));
 sg13g2_nand2_1 _4878_ (.Y(_1368_),
    .A(\FpgaPins_Fpga_LIPSI_acc_a2[0] ),
    .B(_1363_));
 sg13g2_xor2_1 _4879_ (.B(_1363_),
    .A(\FpgaPins_Fpga_LIPSI_acc_a2[0] ),
    .X(_1369_));
 sg13g2_a221oi_1 _4880_ (.B2(net790),
    .C1(net789),
    .B1(_1369_),
    .A1(net781),
    .Y(_1370_),
    .A2(_1367_));
 sg13g2_o21ai_1 _4881_ (.B1(_1370_),
    .Y(_1371_),
    .A1(_1355_),
    .A2(_1364_));
 sg13g2_nor2b_1 _4882_ (.A(_1294_),
    .B_N(_1296_),
    .Y(_1372_));
 sg13g2_and2_1 _4883_ (.A(_1293_),
    .B(net801),
    .X(_1373_));
 sg13g2_nand2_2 _4884_ (.Y(_1374_),
    .A(_1293_),
    .B(net801));
 sg13g2_a21oi_1 _4885_ (.A1(net789),
    .A2(_1368_),
    .Y(_1375_),
    .B1(net786));
 sg13g2_and2_1 _4886_ (.A(_1358_),
    .B(net801),
    .X(_1376_));
 sg13g2_nand2_2 _4887_ (.Y(_1377_),
    .A(_1358_),
    .B(net801));
 sg13g2_or2_1 _4888_ (.X(_1378_),
    .B(_1369_),
    .A(_0122_));
 sg13g2_xnor2_1 _4889_ (.Y(_1379_),
    .A(_0122_),
    .B(_1369_));
 sg13g2_a221oi_1 _4890_ (.B2(net786),
    .C1(net785),
    .B1(_1379_),
    .A1(_1371_),
    .Y(_1380_),
    .A2(_1375_));
 sg13g2_xor2_1 _4891_ (.B(_1369_),
    .A(FpgaPins_Fpga_LIPSI_c_a2),
    .X(_1381_));
 sg13g2_and2_1 _4892_ (.A(_1356_),
    .B(_1372_),
    .X(_1382_));
 sg13g2_nand2_2 _4893_ (.Y(_1383_),
    .A(_1356_),
    .B(_1372_));
 sg13g2_o21ai_1 _4894_ (.B1(_1383_),
    .Y(_1384_),
    .A1(_1377_),
    .A2(_1381_));
 sg13g2_and2_1 _4895_ (.A(_1365_),
    .B(net801),
    .X(_1385_));
 sg13g2_nand2_2 _4896_ (.Y(_1386_),
    .A(_1365_),
    .B(net801));
 sg13g2_a21oi_1 _4897_ (.A1(_1369_),
    .A2(net780),
    .Y(_1387_),
    .B1(net784));
 sg13g2_o21ai_1 _4898_ (.B1(_1387_),
    .Y(_1388_),
    .A1(_1380_),
    .A2(_1384_));
 sg13g2_o21ai_1 _4899_ (.B1(net976),
    .Y(_1389_),
    .A1(_1369_),
    .A2(_1386_));
 sg13g2_nor2b_2 _4900_ (.A(_1389_),
    .B_N(_1388_),
    .Y(\FpgaPins_Fpga_LIPSI_acc_a1[0] ));
 sg13g2_mux2_1 _4901_ (.A0(_0139_),
    .A1(_0138_),
    .S(net808),
    .X(_1390_));
 sg13g2_a21oi_1 _4902_ (.A1(_0733_),
    .A2(net798),
    .Y(_1391_),
    .B1(net819));
 sg13g2_o21ai_1 _4903_ (.B1(_1391_),
    .Y(_1392_),
    .A1(net1737),
    .A2(net798));
 sg13g2_a21oi_1 _4904_ (.A1(net819),
    .A2(_1390_),
    .Y(_1393_),
    .B1(net803));
 sg13g2_mux4_1 _4905_ (.S0(net804),
    .A0(_0133_),
    .A1(_0132_),
    .A2(_0135_),
    .A3(_0134_),
    .S1(net813),
    .X(_1394_));
 sg13g2_o21ai_1 _4906_ (.B1(\FpgaPins_Fpga_FSM_idata_rd_addr_a1[3] ),
    .Y(_1395_),
    .A1(net797),
    .A2(_1394_));
 sg13g2_a21oi_1 _4907_ (.A1(_1392_),
    .A2(_1393_),
    .Y(_1396_),
    .B1(_1395_));
 sg13g2_mux4_1 _4908_ (.S0(net804),
    .A0(_0125_),
    .A1(_0124_),
    .A2(_0127_),
    .A3(_0126_),
    .S1(net812),
    .X(_1397_));
 sg13g2_nor2_1 _4909_ (.A(net796),
    .B(_1397_),
    .Y(_1398_));
 sg13g2_mux2_1 _4910_ (.A0(_0131_),
    .A1(_0130_),
    .S(net807),
    .X(_1399_));
 sg13g2_nand2b_1 _4911_ (.Y(_1400_),
    .B(net799),
    .A_N(_0129_));
 sg13g2_a21oi_1 _4912_ (.A1(_0732_),
    .A2(net807),
    .Y(_1401_),
    .B1(net817));
 sg13g2_a221oi_1 _4913_ (.B2(_1401_),
    .C1(net803),
    .B1(_1400_),
    .A1(net817),
    .Y(_1402_),
    .A2(_1399_));
 sg13g2_nor3_2 _4914_ (.A(net794),
    .B(_1398_),
    .C(_1402_),
    .Y(_1403_));
 sg13g2_nor2_1 _4915_ (.A(_1396_),
    .B(_1403_),
    .Y(\FpgaPins_Fpga_FSM_data_a1[1] ));
 sg13g2_o21ai_1 _4916_ (.B1(net981),
    .Y(_1404_),
    .A1(_1396_),
    .A2(_1403_));
 sg13g2_nand2_2 _4917_ (.Y(_1405_),
    .A(FpgaPins_Fpga_LIPSI_is_ALU_imm_a2),
    .B(_0850_));
 sg13g2_and2_1 _4918_ (.A(_1404_),
    .B(_1405_),
    .X(_1406_));
 sg13g2_a21o_1 _4919_ (.A2(_1405_),
    .A1(_1404_),
    .B1(\FpgaPins_Fpga_LIPSI_acc_a2[1] ),
    .X(_1407_));
 sg13g2_nand3_1 _4920_ (.B(_1404_),
    .C(_1405_),
    .A(\FpgaPins_Fpga_LIPSI_acc_a2[1] ),
    .Y(_1408_));
 sg13g2_a21oi_1 _4921_ (.A1(_1404_),
    .A2(_1405_),
    .Y(_1409_),
    .B1(_0701_));
 sg13g2_nand3_1 _4922_ (.B(_1404_),
    .C(_1405_),
    .A(_0701_),
    .Y(_1410_));
 sg13g2_and2_1 _4923_ (.A(_1407_),
    .B(_1408_),
    .X(_1411_));
 sg13g2_nand3_1 _4924_ (.B(_1361_),
    .C(_1362_),
    .A(_0022_),
    .Y(_1412_));
 sg13g2_xnor2_1 _4925_ (.Y(_1413_),
    .A(_1411_),
    .B(_1412_));
 sg13g2_o21ai_1 _4926_ (.B1(net786),
    .Y(_1414_),
    .A1(_1378_),
    .A2(_1413_));
 sg13g2_a21oi_1 _4927_ (.A1(_1378_),
    .A2(_1413_),
    .Y(_1415_),
    .B1(_1414_));
 sg13g2_a21o_1 _4928_ (.A2(_1408_),
    .A1(net790),
    .B1(net781),
    .X(_1416_));
 sg13g2_nand2_1 _4929_ (.Y(_1417_),
    .A(_1407_),
    .B(_1416_));
 sg13g2_nor3_1 _4930_ (.A(_0699_),
    .B(_1396_),
    .C(_1403_),
    .Y(_1418_));
 sg13g2_o21ai_1 _4931_ (.B1(_1340_),
    .Y(_1419_),
    .A1(net988),
    .A2(_0025_));
 sg13g2_a21oi_1 _4932_ (.A1(_0028_),
    .A2(net793),
    .Y(_1420_),
    .B1(net792));
 sg13g2_o21ai_1 _4933_ (.B1(_1420_),
    .Y(_1421_),
    .A1(_1418_),
    .A2(_1419_));
 sg13g2_nand2_1 _4934_ (.Y(_1422_),
    .A(_0697_),
    .B(net792));
 sg13g2_nand3_1 _4935_ (.B(_1421_),
    .C(_1422_),
    .A(_1348_),
    .Y(_1423_));
 sg13g2_nand2_1 _4936_ (.Y(_1424_),
    .A(_1299_),
    .B(_1360_));
 sg13g2_a221oi_1 _4937_ (.B2(_0028_),
    .C1(_1424_),
    .B1(_1352_),
    .A1(_0022_),
    .Y(_1425_),
    .A2(net791));
 sg13g2_a221oi_1 _4938_ (.B2(_1425_),
    .C1(net788),
    .B1(_1423_),
    .A1(net800),
    .Y(_1426_),
    .A2(_1406_));
 sg13g2_nand2b_1 _4939_ (.Y(_1427_),
    .B(_1406_),
    .A_N(_0025_));
 sg13g2_a22oi_1 _4940_ (.Y(_1428_),
    .B1(_1427_),
    .B2(net788),
    .A2(_1426_),
    .A1(_1417_));
 sg13g2_nor2_1 _4941_ (.A(net786),
    .B(_1428_),
    .Y(_1429_));
 sg13g2_nand4_1 _4942_ (.B(_1363_),
    .C(_1407_),
    .A(\FpgaPins_Fpga_LIPSI_acc_a2[0] ),
    .Y(_1430_),
    .D(_1408_));
 sg13g2_xnor2_1 _4943_ (.Y(_1431_),
    .A(_1368_),
    .B(_1411_));
 sg13g2_a21oi_1 _4944_ (.A1(FpgaPins_Fpga_LIPSI_c_a2),
    .A2(_1369_),
    .Y(_1432_),
    .B1(_1431_));
 sg13g2_and3_1 _4945_ (.X(_1433_),
    .A(FpgaPins_Fpga_LIPSI_c_a2),
    .B(_1369_),
    .C(_1411_));
 sg13g2_o21ai_1 _4946_ (.B1(net785),
    .Y(_1434_),
    .A1(_1432_),
    .A2(_1433_));
 sg13g2_o21ai_1 _4947_ (.B1(_1377_),
    .Y(_1435_),
    .A1(_1415_),
    .A2(_1429_));
 sg13g2_nand3_1 _4948_ (.B(_1434_),
    .C(_1435_),
    .A(_1383_),
    .Y(_1436_));
 sg13g2_a21oi_1 _4949_ (.A1(net780),
    .A2(_1413_),
    .Y(_1437_),
    .B1(net784));
 sg13g2_o21ai_1 _4950_ (.B1(net976),
    .Y(_1438_),
    .A1(_1386_),
    .A2(_1431_));
 sg13g2_a21oi_2 _4951_ (.B1(_1438_),
    .Y(\FpgaPins_Fpga_LIPSI_acc_a1[1] ),
    .A2(_1437_),
    .A1(_1436_));
 sg13g2_mux2_1 _4952_ (.A0(_0151_),
    .A1(_0150_),
    .S(net806),
    .X(_1439_));
 sg13g2_a21oi_1 _4953_ (.A1(_0735_),
    .A2(net806),
    .Y(_1440_),
    .B1(net814));
 sg13g2_o21ai_1 _4954_ (.B1(_1440_),
    .Y(_1441_),
    .A1(_0149_),
    .A2(net805));
 sg13g2_a21oi_1 _4955_ (.A1(net813),
    .A2(_1439_),
    .Y(_1442_),
    .B1(net797));
 sg13g2_a21oi_1 _4956_ (.A1(_0736_),
    .A2(net808),
    .Y(_1443_),
    .B1(net819));
 sg13g2_o21ai_1 _4957_ (.B1(_1443_),
    .Y(_1444_),
    .A1(net1738),
    .A2(net808));
 sg13g2_mux2_1 _4958_ (.A0(_0155_),
    .A1(_0154_),
    .S(net808),
    .X(_1445_));
 sg13g2_a21oi_1 _4959_ (.A1(net819),
    .A2(_1445_),
    .Y(_1446_),
    .B1(net803));
 sg13g2_a221oi_1 _4960_ (.B2(_1446_),
    .C1(_1325_),
    .B1(_1444_),
    .A1(_1441_),
    .Y(_1447_),
    .A2(_1442_));
 sg13g2_mux4_1 _4961_ (.S0(net805),
    .A0(_0141_),
    .A1(_0140_),
    .A2(_0143_),
    .A3(_0142_),
    .S1(net814),
    .X(_1448_));
 sg13g2_nor2_1 _4962_ (.A(net795),
    .B(_1448_),
    .Y(_1449_));
 sg13g2_mux2_1 _4963_ (.A0(_0147_),
    .A1(_0146_),
    .S(net807),
    .X(_1450_));
 sg13g2_nand2b_1 _4964_ (.Y(_1451_),
    .B(net799),
    .A_N(_0145_));
 sg13g2_a21oi_1 _4965_ (.A1(_0734_),
    .A2(net807),
    .Y(_1452_),
    .B1(net817));
 sg13g2_a221oi_1 _4966_ (.B2(_1452_),
    .C1(net803),
    .B1(_1451_),
    .A1(net817),
    .Y(_1453_),
    .A2(_1450_));
 sg13g2_nor3_2 _4967_ (.A(net794),
    .B(_1449_),
    .C(_1453_),
    .Y(_1454_));
 sg13g2_nor2_2 _4968_ (.A(net1739),
    .B(_1454_),
    .Y(\FpgaPins_Fpga_FSM_data_a1[2] ));
 sg13g2_nor2_1 _4969_ (.A(_0728_),
    .B(_1043_),
    .Y(_1455_));
 sg13g2_a21oi_2 _4970_ (.B1(_1455_),
    .Y(_1456_),
    .A2(\FpgaPins_Fpga_FSM_data_a1[2] ),
    .A1(net981));
 sg13g2_inv_1 _4971_ (.Y(_1457_),
    .A(_1456_));
 sg13g2_nor2b_1 _4972_ (.A(_1456_),
    .B_N(\FpgaPins_Fpga_LIPSI_acc_a2[2] ),
    .Y(_1458_));
 sg13g2_nor2_1 _4973_ (.A(\FpgaPins_Fpga_LIPSI_acc_a2[2] ),
    .B(_1457_),
    .Y(_1459_));
 sg13g2_xnor2_1 _4974_ (.Y(_1460_),
    .A(\FpgaPins_Fpga_LIPSI_acc_a2[2] ),
    .B(_1456_));
 sg13g2_xor2_1 _4975_ (.B(_1456_),
    .A(\FpgaPins_Fpga_LIPSI_acc_a2[2] ),
    .X(_1461_));
 sg13g2_a21oi_1 _4976_ (.A1(_1410_),
    .A2(_1412_),
    .Y(_1462_),
    .B1(_1409_));
 sg13g2_xnor2_1 _4977_ (.Y(_1463_),
    .A(_1461_),
    .B(_1462_));
 sg13g2_o21ai_1 _4978_ (.B1(_1463_),
    .Y(_1464_),
    .A1(_1378_),
    .A2(_1413_));
 sg13g2_nor3_2 _4979_ (.A(_1378_),
    .B(_1413_),
    .C(_1463_),
    .Y(_1465_));
 sg13g2_nor2_1 _4980_ (.A(_1374_),
    .B(_1465_),
    .Y(_1466_));
 sg13g2_o21ai_1 _4981_ (.B1(_1340_),
    .Y(_1467_),
    .A1(net988),
    .A2(_0028_));
 sg13g2_a21oi_1 _4982_ (.A1(net988),
    .A2(\FpgaPins_Fpga_FSM_data_a1[2] ),
    .Y(_1468_),
    .B1(_1467_));
 sg13g2_a21oi_1 _4983_ (.A1(_0031_),
    .A2(net793),
    .Y(_1469_),
    .B1(net792));
 sg13g2_nand2b_1 _4984_ (.Y(_1470_),
    .B(_1469_),
    .A_N(_1468_));
 sg13g2_nand2b_1 _4985_ (.Y(_1471_),
    .B(net792),
    .A_N(_0025_));
 sg13g2_nand3_1 _4986_ (.B(_1470_),
    .C(_1471_),
    .A(_1348_),
    .Y(_1472_));
 sg13g2_a221oi_1 _4987_ (.B2(_0031_),
    .C1(net800),
    .B1(_1352_),
    .A1(_0025_),
    .Y(_1473_),
    .A2(net791));
 sg13g2_a22oi_1 _4988_ (.Y(_1474_),
    .B1(_1472_),
    .B2(_1473_),
    .A2(_1457_),
    .A1(net800));
 sg13g2_a21oi_1 _4989_ (.A1(net790),
    .A2(_1460_),
    .Y(_1475_),
    .B1(net781));
 sg13g2_o21ai_1 _4990_ (.B1(_1475_),
    .Y(_1476_),
    .A1(net790),
    .A2(_1474_));
 sg13g2_a21oi_1 _4991_ (.A1(net781),
    .A2(_1459_),
    .Y(_1477_),
    .B1(net788));
 sg13g2_a221oi_1 _4992_ (.B2(_1477_),
    .C1(net786),
    .B1(_1476_),
    .A1(net788),
    .Y(_1478_),
    .A2(_1458_));
 sg13g2_a221oi_1 _4993_ (.B2(_1466_),
    .C1(_1478_),
    .B1(_1464_),
    .A1(_1358_),
    .Y(_1479_),
    .A2(net801));
 sg13g2_nand2_1 _4994_ (.Y(_1480_),
    .A(_1427_),
    .B(_1430_));
 sg13g2_a21oi_1 _4995_ (.A1(_1427_),
    .A2(_1430_),
    .Y(_1481_),
    .B1(_1461_));
 sg13g2_xnor2_1 _4996_ (.Y(_1482_),
    .A(_1461_),
    .B(_1480_));
 sg13g2_xnor2_1 _4997_ (.Y(_1483_),
    .A(_1460_),
    .B(_1480_));
 sg13g2_nand2_1 _4998_ (.Y(_1484_),
    .A(_1433_),
    .B(_1482_));
 sg13g2_o21ai_1 _4999_ (.B1(net785),
    .Y(_1485_),
    .A1(_1433_),
    .A2(_1482_));
 sg13g2_nor2b_1 _5000_ (.A(_1485_),
    .B_N(_1484_),
    .Y(_1486_));
 sg13g2_o21ai_1 _5001_ (.B1(_1383_),
    .Y(_1487_),
    .A1(_1479_),
    .A2(_1486_));
 sg13g2_a21oi_1 _5002_ (.A1(net780),
    .A2(_1463_),
    .Y(_1488_),
    .B1(net784));
 sg13g2_a221oi_1 _5003_ (.B2(_1488_),
    .C1(net947),
    .B1(_1487_),
    .A1(net784),
    .Y(\FpgaPins_Fpga_LIPSI_acc_a1[2] ),
    .A2(_1483_));
 sg13g2_mux2_1 _5004_ (.A0(_0171_),
    .A1(_0170_),
    .S(net810),
    .X(_1489_));
 sg13g2_a21oi_1 _5005_ (.A1(_0738_),
    .A2(\FpgaPins_Fpga_FSM_idata_rd_addr_a1[0] ),
    .Y(_1490_),
    .B1(net819));
 sg13g2_o21ai_1 _5006_ (.B1(_1490_),
    .Y(_1491_),
    .A1(net1718),
    .A2(net798));
 sg13g2_a21oi_1 _5007_ (.A1(net819),
    .A2(_1489_),
    .Y(_1492_),
    .B1(_1316_));
 sg13g2_mux4_1 _5008_ (.S0(net804),
    .A0(_0165_),
    .A1(_0164_),
    .A2(_0167_),
    .A3(_0166_),
    .S1(net813),
    .X(_1493_));
 sg13g2_o21ai_1 _5009_ (.B1(\FpgaPins_Fpga_FSM_idata_rd_addr_a1[3] ),
    .Y(_1494_),
    .A1(net797),
    .A2(_1493_));
 sg13g2_a21oi_1 _5010_ (.A1(net1719),
    .A2(_1492_),
    .Y(_1495_),
    .B1(_1494_));
 sg13g2_mux4_1 _5011_ (.S0(net805),
    .A0(_0157_),
    .A1(_0156_),
    .A2(_0159_),
    .A3(_0158_),
    .S1(net812),
    .X(_1496_));
 sg13g2_nor2_1 _5012_ (.A(net796),
    .B(_1496_),
    .Y(_1497_));
 sg13g2_mux2_1 _5013_ (.A0(_0163_),
    .A1(_0162_),
    .S(net811),
    .X(_1498_));
 sg13g2_nand2b_1 _5014_ (.Y(_1499_),
    .B(net799),
    .A_N(_0161_));
 sg13g2_a21oi_1 _5015_ (.A1(_0737_),
    .A2(net809),
    .Y(_1500_),
    .B1(net815));
 sg13g2_a221oi_1 _5016_ (.B2(_1500_),
    .C1(net802),
    .B1(_1499_),
    .A1(net815),
    .Y(_1501_),
    .A2(_1498_));
 sg13g2_nor3_2 _5017_ (.A(net794),
    .B(_1497_),
    .C(_1501_),
    .Y(_1502_));
 sg13g2_nor2_2 _5018_ (.A(_1495_),
    .B(_1502_),
    .Y(\FpgaPins_Fpga_FSM_data_a1[3] ));
 sg13g2_mux2_2 _5019_ (.A0(\FpgaPins_Fpga_FSM_instr_a1[3] ),
    .A1(\FpgaPins_Fpga_FSM_data_a1[3] ),
    .S(net981),
    .X(_1503_));
 sg13g2_inv_1 _5020_ (.Y(_1504_),
    .A(_1503_));
 sg13g2_nor2_1 _5021_ (.A(\FpgaPins_Fpga_LIPSI_acc_a2[3] ),
    .B(_1503_),
    .Y(_1505_));
 sg13g2_nand2_2 _5022_ (.Y(_1506_),
    .A(_0704_),
    .B(_1503_));
 sg13g2_inv_1 _5023_ (.Y(_1507_),
    .A(_1506_));
 sg13g2_nand2b_1 _5024_ (.Y(_1508_),
    .B(_1506_),
    .A_N(_1505_));
 sg13g2_nand2_1 _5025_ (.Y(_1509_),
    .A(_0703_),
    .B(_1456_));
 sg13g2_o21ai_1 _5026_ (.B1(_1509_),
    .Y(_1510_),
    .A1(_1460_),
    .A2(_1462_));
 sg13g2_xnor2_1 _5027_ (.Y(_1511_),
    .A(_1508_),
    .B(_1510_));
 sg13g2_nor2_1 _5028_ (.A(_1465_),
    .B(_1511_),
    .Y(_1512_));
 sg13g2_nand2_2 _5029_ (.Y(_1513_),
    .A(_1465_),
    .B(_1511_));
 sg13g2_nor2_1 _5030_ (.A(_1374_),
    .B(_1512_),
    .Y(_1514_));
 sg13g2_o21ai_1 _5031_ (.B1(_1340_),
    .Y(_1515_),
    .A1(net988),
    .A2(_0031_));
 sg13g2_a21oi_1 _5032_ (.A1(net988),
    .A2(\FpgaPins_Fpga_FSM_data_a1[3] ),
    .Y(_1516_),
    .B1(_1515_));
 sg13g2_a21o_1 _5033_ (.A2(net793),
    .A1(_0172_),
    .B1(net792),
    .X(_1517_));
 sg13g2_a21oi_1 _5034_ (.A1(_0703_),
    .A2(_1342_),
    .Y(_1518_),
    .B1(_1347_));
 sg13g2_o21ai_1 _5035_ (.B1(_1518_),
    .Y(_1519_),
    .A1(_1516_),
    .A2(_1517_));
 sg13g2_a221oi_1 _5036_ (.B2(_0172_),
    .C1(net800),
    .B1(_1354_),
    .A1(_0028_),
    .Y(_1520_),
    .A2(net791));
 sg13g2_xor2_1 _5037_ (.B(_1503_),
    .A(\FpgaPins_Fpga_LIPSI_acc_a2[3] ),
    .X(_1521_));
 sg13g2_nand2_1 _5038_ (.Y(_1522_),
    .A(net790),
    .B(_1521_));
 sg13g2_a22oi_1 _5039_ (.Y(_1523_),
    .B1(_1519_),
    .B2(_1520_),
    .A2(_1503_),
    .A1(net800));
 sg13g2_o21ai_1 _5040_ (.B1(_1522_),
    .Y(_1524_),
    .A1(net790),
    .A2(_1523_));
 sg13g2_a21oi_1 _5041_ (.A1(net781),
    .A2(_1505_),
    .Y(_1525_),
    .B1(net788));
 sg13g2_o21ai_1 _5042_ (.B1(_1525_),
    .Y(_1526_),
    .A1(net781),
    .A2(_1524_));
 sg13g2_a21oi_1 _5043_ (.A1(net789),
    .A2(_1507_),
    .Y(_1527_),
    .B1(net786));
 sg13g2_a22oi_1 _5044_ (.Y(_1528_),
    .B1(_1526_),
    .B2(_1527_),
    .A2(_1514_),
    .A1(_1513_));
 sg13g2_o21ai_1 _5045_ (.B1(_1521_),
    .Y(_1529_),
    .A1(_1458_),
    .A2(_1481_));
 sg13g2_or3_1 _5046_ (.A(_1458_),
    .B(_1481_),
    .C(_1521_),
    .X(_1530_));
 sg13g2_nand2_2 _5047_ (.Y(_1531_),
    .A(_1529_),
    .B(_1530_));
 sg13g2_nor2_2 _5048_ (.A(_1484_),
    .B(_1531_),
    .Y(_1532_));
 sg13g2_nand2_1 _5049_ (.Y(_1533_),
    .A(_1484_),
    .B(_1531_));
 sg13g2_nor2_1 _5050_ (.A(_1377_),
    .B(_1532_),
    .Y(_1534_));
 sg13g2_a22oi_1 _5051_ (.Y(_1535_),
    .B1(_1533_),
    .B2(_1534_),
    .A2(_1528_),
    .A1(_1377_));
 sg13g2_nor2_1 _5052_ (.A(net780),
    .B(_1535_),
    .Y(_1536_));
 sg13g2_o21ai_1 _5053_ (.B1(_1386_),
    .Y(_1537_),
    .A1(_1383_),
    .A2(_1511_));
 sg13g2_o21ai_1 _5054_ (.B1(net976),
    .Y(_1538_),
    .A1(_1536_),
    .A2(_1537_));
 sg13g2_a21oi_2 _5055_ (.B1(_1538_),
    .Y(\FpgaPins_Fpga_LIPSI_acc_a1[3] ),
    .A2(_1531_),
    .A1(net784));
 sg13g2_mux4_1 _5056_ (.S0(net804),
    .A0(_0182_),
    .A1(_0181_),
    .A2(_0184_),
    .A3(_0183_),
    .S1(net813),
    .X(_1539_));
 sg13g2_nor2_1 _5057_ (.A(net797),
    .B(_1539_),
    .Y(_1540_));
 sg13g2_nand2b_1 _5058_ (.Y(_1541_),
    .B(net810),
    .A_N(_0185_));
 sg13g2_a21oi_1 _5059_ (.A1(_0741_),
    .A2(net798),
    .Y(_1542_),
    .B1(net818));
 sg13g2_mux2_1 _5060_ (.A0(_0188_),
    .A1(_0187_),
    .S(net810),
    .X(_1543_));
 sg13g2_a221oi_1 _5061_ (.B2(net818),
    .C1(net802),
    .B1(_1543_),
    .A1(_1541_),
    .Y(_1544_),
    .A2(_1542_));
 sg13g2_nor3_1 _5062_ (.A(_1325_),
    .B(_1540_),
    .C(_1544_),
    .Y(_1545_));
 sg13g2_mux4_1 _5063_ (.S0(net804),
    .A0(_0174_),
    .A1(_0173_),
    .A2(_0176_),
    .A3(_0175_),
    .S1(net812),
    .X(_1546_));
 sg13g2_nor2_1 _5064_ (.A(net795),
    .B(_1546_),
    .Y(_1547_));
 sg13g2_mux2_1 _5065_ (.A0(_0180_),
    .A1(_0179_),
    .S(net807),
    .X(_1548_));
 sg13g2_nand2b_1 _5066_ (.Y(_1549_),
    .B(net799),
    .A_N(_0178_));
 sg13g2_a21oi_1 _5067_ (.A1(_0740_),
    .A2(net807),
    .Y(_1550_),
    .B1(net817));
 sg13g2_a221oi_1 _5068_ (.B2(_1550_),
    .C1(net803),
    .B1(_1549_),
    .A1(net817),
    .Y(_1551_),
    .A2(_1548_));
 sg13g2_nor3_2 _5069_ (.A(net794),
    .B(_1547_),
    .C(_1551_),
    .Y(_1552_));
 sg13g2_nor2_2 _5070_ (.A(_1545_),
    .B(_1552_),
    .Y(\FpgaPins_Fpga_FSM_data_a1[4] ));
 sg13g2_nand2_1 _5071_ (.Y(_1553_),
    .A(net981),
    .B(\FpgaPins_Fpga_FSM_data_a1[4] ));
 sg13g2_o21ai_1 _5072_ (.B1(_1553_),
    .Y(_1554_),
    .A1(net981),
    .A2(_1060_));
 sg13g2_and2_1 _5073_ (.A(\FpgaPins_Fpga_LIPSI_acc_a2[4] ),
    .B(_1554_),
    .X(_1555_));
 sg13g2_inv_1 _5074_ (.Y(_1556_),
    .A(_1555_));
 sg13g2_xor2_1 _5075_ (.B(_1554_),
    .A(\FpgaPins_Fpga_LIPSI_acc_a2[4] ),
    .X(_1557_));
 sg13g2_inv_1 _5076_ (.Y(_1558_),
    .A(_1557_));
 sg13g2_a22oi_1 _5077_ (.Y(_1559_),
    .B1(_1508_),
    .B2(_1510_),
    .A2(_1504_),
    .A1(\FpgaPins_Fpga_LIPSI_acc_a2[3] ));
 sg13g2_xnor2_1 _5078_ (.Y(_1560_),
    .A(_1557_),
    .B(_1559_));
 sg13g2_nor2b_1 _5079_ (.A(_1513_),
    .B_N(_1560_),
    .Y(_1561_));
 sg13g2_xor2_1 _5080_ (.B(_1560_),
    .A(_1513_),
    .X(_1562_));
 sg13g2_nor2_1 _5081_ (.A(_0743_),
    .B(_1337_),
    .Y(_1563_));
 sg13g2_a21oi_1 _5082_ (.A1(_0699_),
    .A2(_0172_),
    .Y(_1564_),
    .B1(_1339_));
 sg13g2_o21ai_1 _5083_ (.B1(_1564_),
    .Y(_1565_),
    .A1(_0699_),
    .A2(\FpgaPins_Fpga_FSM_data_a1[4] ));
 sg13g2_o21ai_1 _5084_ (.B1(_1565_),
    .Y(_1566_),
    .A1(_1338_),
    .A2(_1563_));
 sg13g2_a22oi_1 _5085_ (.Y(_1567_),
    .B1(_1352_),
    .B2(_0189_),
    .A2(_1342_),
    .A1(_0031_));
 sg13g2_a21oi_1 _5086_ (.A1(_1566_),
    .A2(_1567_),
    .Y(_1568_),
    .B1(_1298_));
 sg13g2_o21ai_1 _5087_ (.B1(_1360_),
    .Y(_1569_),
    .A1(_1299_),
    .A2(_1554_));
 sg13g2_nor2_1 _5088_ (.A(_1568_),
    .B(_1569_),
    .Y(_1570_));
 sg13g2_o21ai_1 _5089_ (.B1(net781),
    .Y(_1571_),
    .A1(\FpgaPins_Fpga_LIPSI_acc_a2[4] ),
    .A2(_1554_));
 sg13g2_o21ai_1 _5090_ (.B1(_1571_),
    .Y(_1572_),
    .A1(_1360_),
    .A2(_1558_));
 sg13g2_or3_1 _5091_ (.A(net788),
    .B(_1570_),
    .C(_1572_),
    .X(_1573_));
 sg13g2_a21oi_1 _5092_ (.A1(net789),
    .A2(_1556_),
    .Y(_1574_),
    .B1(net787));
 sg13g2_a221oi_1 _5093_ (.B2(_1574_),
    .C1(net785),
    .B1(_1573_),
    .A1(net787),
    .Y(_1575_),
    .A2(_1562_));
 sg13g2_a21oi_2 _5094_ (.B1(_1558_),
    .Y(_1576_),
    .A2(_1529_),
    .A1(_1506_));
 sg13g2_nand3_1 _5095_ (.B(_1529_),
    .C(_1558_),
    .A(_1506_),
    .Y(_1577_));
 sg13g2_nor2b_2 _5096_ (.A(_1576_),
    .B_N(_1577_),
    .Y(_1578_));
 sg13g2_xnor2_1 _5097_ (.Y(_1579_),
    .A(_1532_),
    .B(_1578_));
 sg13g2_a221oi_1 _5098_ (.B2(_1579_),
    .C1(_1575_),
    .B1(net785),
    .A1(_1356_),
    .Y(_1580_),
    .A2(net801));
 sg13g2_o21ai_1 _5099_ (.B1(_1386_),
    .Y(_1581_),
    .A1(_1383_),
    .A2(_1560_));
 sg13g2_nor2_1 _5100_ (.A(_1386_),
    .B(_1578_),
    .Y(_1582_));
 sg13g2_o21ai_1 _5101_ (.B1(net975),
    .Y(_1583_),
    .A1(_1580_),
    .A2(_1581_));
 sg13g2_nor2_2 _5102_ (.A(_1582_),
    .B(_1583_),
    .Y(\FpgaPins_Fpga_LIPSI_acc_a1[4] ));
 sg13g2_mux4_1 _5103_ (.S0(net806),
    .A0(\datam[9][5] ),
    .A1(\datam[8][5] ),
    .A2(\datam[11][5] ),
    .A3(\datam[10][5] ),
    .S1(net812),
    .X(_1584_));
 sg13g2_nor2_1 _5104_ (.A(net795),
    .B(_1584_),
    .Y(_1585_));
 sg13g2_nand2b_1 _5105_ (.Y(_1586_),
    .B(net811),
    .A_N(\datam[12][5] ));
 sg13g2_a21oi_1 _5106_ (.A1(_0745_),
    .A2(net798),
    .Y(_1587_),
    .B1(net818));
 sg13g2_mux2_1 _5107_ (.A0(\datam[15][5] ),
    .A1(\datam[14][5] ),
    .S(net810),
    .X(_1588_));
 sg13g2_a221oi_1 _5108_ (.B2(net818),
    .C1(net802),
    .B1(_1588_),
    .A1(_1586_),
    .Y(_1589_),
    .A2(_1587_));
 sg13g2_nor3_1 _5109_ (.A(_1325_),
    .B(_1585_),
    .C(_1589_),
    .Y(_1590_));
 sg13g2_mux4_1 _5110_ (.S0(net804),
    .A0(\datam[1][5] ),
    .A1(\datam[0][5] ),
    .A2(\datam[3][5] ),
    .A3(\datam[2][5] ),
    .S1(net812),
    .X(_1591_));
 sg13g2_nor2_1 _5111_ (.A(net795),
    .B(_1591_),
    .Y(_1592_));
 sg13g2_mux2_1 _5112_ (.A0(\datam[7][5] ),
    .A1(\datam[6][5] ),
    .S(net811),
    .X(_1593_));
 sg13g2_nand2b_1 _5113_ (.Y(_1594_),
    .B(net799),
    .A_N(\datam[5][5] ));
 sg13g2_a21oi_1 _5114_ (.A1(_0744_),
    .A2(net808),
    .Y(_1595_),
    .B1(net815));
 sg13g2_a221oi_1 _5115_ (.B2(_1595_),
    .C1(net802),
    .B1(_1594_),
    .A1(net815),
    .Y(_1596_),
    .A2(_1593_));
 sg13g2_nor3_2 _5116_ (.A(net794),
    .B(_1592_),
    .C(_1596_),
    .Y(_1597_));
 sg13g2_nor2_2 _5117_ (.A(_1590_),
    .B(_1597_),
    .Y(_1598_));
 sg13g2_inv_1 _5118_ (.Y(\FpgaPins_Fpga_FSM_data_a1[5] ),
    .A(_1598_));
 sg13g2_nor2_1 _5119_ (.A(FpgaPins_Fpga_LIPSI_is_ALU_imm_a2),
    .B(_1598_),
    .Y(_1599_));
 sg13g2_a21oi_2 _5120_ (.B1(_1599_),
    .Y(_1600_),
    .A2(net875),
    .A1(FpgaPins_Fpga_LIPSI_is_ALU_imm_a2));
 sg13g2_nor2_1 _5121_ (.A(_0189_),
    .B(_1600_),
    .Y(_1601_));
 sg13g2_inv_1 _5122_ (.Y(_1602_),
    .A(_1601_));
 sg13g2_a21oi_1 _5123_ (.A1(_0742_),
    .A2(_1600_),
    .Y(_1603_),
    .B1(_1601_));
 sg13g2_inv_1 _5124_ (.Y(_1604_),
    .A(_1603_));
 sg13g2_nand2b_1 _5125_ (.Y(_1605_),
    .B(_0739_),
    .A_N(_1554_));
 sg13g2_o21ai_1 _5126_ (.B1(_1605_),
    .Y(_1606_),
    .A1(_1557_),
    .A2(_1559_));
 sg13g2_xnor2_1 _5127_ (.Y(_1607_),
    .A(_1604_),
    .B(_1606_));
 sg13g2_and2_1 _5128_ (.A(_1561_),
    .B(_1607_),
    .X(_1608_));
 sg13g2_o21ai_1 _5129_ (.B1(net787),
    .Y(_1609_),
    .A1(_1561_),
    .A2(_1607_));
 sg13g2_o21ai_1 _5130_ (.B1(_1347_),
    .Y(_1610_),
    .A1(_0746_),
    .A2(_0867_));
 sg13g2_a21oi_1 _5131_ (.A1(_0699_),
    .A2(_0189_),
    .Y(_1611_),
    .B1(net793));
 sg13g2_o21ai_1 _5132_ (.B1(_1611_),
    .Y(_1612_),
    .A1(_0699_),
    .A2(\FpgaPins_Fpga_FSM_data_a1[5] ));
 sg13g2_a21oi_1 _5133_ (.A1(_0746_),
    .A2(_1339_),
    .Y(_1613_),
    .B1(_1344_));
 sg13g2_a21o_1 _5134_ (.A2(net792),
    .A1(_0172_),
    .B1(_1354_),
    .X(_1614_));
 sg13g2_a21o_1 _5135_ (.A2(_1613_),
    .A1(_1612_),
    .B1(_1614_),
    .X(_1615_));
 sg13g2_a221oi_1 _5136_ (.B2(_1615_),
    .C1(_1298_),
    .B1(_1610_),
    .A1(_0172_),
    .Y(_1616_),
    .A2(net791));
 sg13g2_o21ai_1 _5137_ (.B1(_1360_),
    .Y(_1617_),
    .A1(_1299_),
    .A2(_1600_));
 sg13g2_xnor2_1 _5138_ (.Y(_1618_),
    .A(\FpgaPins_Fpga_LIPSI_acc_a2[5] ),
    .B(_1600_));
 sg13g2_inv_1 _5139_ (.Y(_1619_),
    .A(_1618_));
 sg13g2_a21oi_1 _5140_ (.A1(\FpgaPins_Fpga_LIPSI_acc_a2[5] ),
    .A2(net782),
    .Y(_1620_),
    .B1(_1360_));
 sg13g2_a21oi_1 _5141_ (.A1(_1619_),
    .A2(_1620_),
    .Y(_1621_),
    .B1(net788));
 sg13g2_o21ai_1 _5142_ (.B1(_1621_),
    .Y(_1622_),
    .A1(_1616_),
    .A2(_1617_));
 sg13g2_a21oi_1 _5143_ (.A1(net789),
    .A2(_1601_),
    .Y(_1623_),
    .B1(net786));
 sg13g2_a21oi_1 _5144_ (.A1(_1622_),
    .A2(_1623_),
    .Y(_1624_),
    .B1(net785));
 sg13g2_o21ai_1 _5145_ (.B1(_1624_),
    .Y(_1625_),
    .A1(_1608_),
    .A2(_1609_));
 sg13g2_o21ai_1 _5146_ (.B1(_1618_),
    .Y(_1626_),
    .A1(_1555_),
    .A2(_1576_));
 sg13g2_or3_1 _5147_ (.A(_1555_),
    .B(_1576_),
    .C(_1618_),
    .X(_1627_));
 sg13g2_nand2_1 _5148_ (.Y(_1628_),
    .A(_1626_),
    .B(_1627_));
 sg13g2_nand4_1 _5149_ (.B(_1578_),
    .C(_1626_),
    .A(_1532_),
    .Y(_1629_),
    .D(_1627_));
 sg13g2_a22oi_1 _5150_ (.Y(_1630_),
    .B1(_1626_),
    .B2(_1627_),
    .A2(_1578_),
    .A1(_1532_));
 sg13g2_nand3b_1 _5151_ (.B(_1376_),
    .C(_1629_),
    .Y(_1631_),
    .A_N(_1630_));
 sg13g2_a21o_1 _5152_ (.A2(_1631_),
    .A1(_1625_),
    .B1(_1382_),
    .X(_1632_));
 sg13g2_nor2_1 _5153_ (.A(_1383_),
    .B(_1607_),
    .Y(_1633_));
 sg13g2_nor2_1 _5154_ (.A(_1385_),
    .B(_1633_),
    .Y(_1634_));
 sg13g2_a221oi_1 _5155_ (.B2(_1634_),
    .C1(net944),
    .B1(_1632_),
    .A1(_1385_),
    .Y(\FpgaPins_Fpga_LIPSI_acc_a1[5] ),
    .A2(_1628_));
 sg13g2_mux2_1 _5156_ (.A0(\datam[11][6] ),
    .A1(\datam[10][6] ),
    .S(net805),
    .X(_1635_));
 sg13g2_a21oi_1 _5157_ (.A1(_0748_),
    .A2(net805),
    .Y(_1636_),
    .B1(net813));
 sg13g2_o21ai_1 _5158_ (.B1(_1636_),
    .Y(_1637_),
    .A1(\datam[9][6] ),
    .A2(net806));
 sg13g2_a21oi_1 _5159_ (.A1(net812),
    .A2(_1635_),
    .Y(_1638_),
    .B1(net795));
 sg13g2_a21oi_1 _5160_ (.A1(_0749_),
    .A2(net809),
    .Y(_1639_),
    .B1(net816));
 sg13g2_o21ai_1 _5161_ (.B1(_1639_),
    .Y(_1640_),
    .A1(\datam[13][6] ),
    .A2(net810));
 sg13g2_mux2_1 _5162_ (.A0(\datam[15][6] ),
    .A1(\datam[14][6] ),
    .S(net810),
    .X(_1641_));
 sg13g2_a21oi_1 _5163_ (.A1(net819),
    .A2(_1641_),
    .Y(_1642_),
    .B1(net803));
 sg13g2_a221oi_1 _5164_ (.B2(_1642_),
    .C1(_1325_),
    .B1(_1640_),
    .A1(_1637_),
    .Y(_1643_),
    .A2(_1638_));
 sg13g2_mux4_1 _5165_ (.S0(net805),
    .A0(\datam[1][6] ),
    .A1(\datam[0][6] ),
    .A2(\datam[3][6] ),
    .A3(\datam[2][6] ),
    .S1(net812),
    .X(_1644_));
 sg13g2_nor2_1 _5166_ (.A(net795),
    .B(_1644_),
    .Y(_1645_));
 sg13g2_mux2_1 _5167_ (.A0(\datam[7][6] ),
    .A1(\datam[6][6] ),
    .S(net809),
    .X(_1646_));
 sg13g2_nand2b_1 _5168_ (.Y(_1647_),
    .B(net799),
    .A_N(\datam[5][6] ));
 sg13g2_a21oi_1 _5169_ (.A1(_0747_),
    .A2(net809),
    .Y(_1648_),
    .B1(net815));
 sg13g2_a221oi_1 _5170_ (.B2(_1648_),
    .C1(net802),
    .B1(_1647_),
    .A1(net816),
    .Y(_1649_),
    .A2(_1646_));
 sg13g2_nor3_1 _5171_ (.A(net794),
    .B(_1645_),
    .C(_1649_),
    .Y(_1650_));
 sg13g2_or2_2 _5172_ (.X(\FpgaPins_Fpga_FSM_data_a1[6] ),
    .B(_1650_),
    .A(_1643_));
 sg13g2_nand2b_1 _5173_ (.Y(_1651_),
    .B(FpgaPins_Fpga_LIPSI_is_ALU_imm_a2),
    .A_N(\FpgaPins_Fpga_FSM_instr_a1[6] ));
 sg13g2_o21ai_1 _5174_ (.B1(_1651_),
    .Y(_1652_),
    .A1(FpgaPins_Fpga_LIPSI_is_ALU_imm_a2),
    .A2(\FpgaPins_Fpga_FSM_data_a1[6] ));
 sg13g2_nor2b_2 _5175_ (.A(_1652_),
    .B_N(\FpgaPins_Fpga_LIPSI_acc_a2[6] ),
    .Y(_1653_));
 sg13g2_nor2b_1 _5176_ (.A(\FpgaPins_Fpga_LIPSI_acc_a2[6] ),
    .B_N(_1652_),
    .Y(_1654_));
 sg13g2_nor2_2 _5177_ (.A(_1653_),
    .B(_1654_),
    .Y(_1655_));
 sg13g2_inv_1 _5178_ (.Y(_1656_),
    .A(_1655_));
 sg13g2_a22oi_1 _5179_ (.Y(_1657_),
    .B1(_1604_),
    .B2(_1606_),
    .A2(_1600_),
    .A1(_0743_));
 sg13g2_xnor2_1 _5180_ (.Y(_1658_),
    .A(_1655_),
    .B(_1657_));
 sg13g2_and2_1 _5181_ (.A(_1608_),
    .B(_1658_),
    .X(_1659_));
 sg13g2_nand2_1 _5182_ (.Y(_1660_),
    .A(_1608_),
    .B(_1658_));
 sg13g2_o21ai_1 _5183_ (.B1(net787),
    .Y(_1661_),
    .A1(_1608_),
    .A2(_1658_));
 sg13g2_o21ai_1 _5184_ (.B1(_1340_),
    .Y(_1662_),
    .A1(net989),
    .A2(_0190_));
 sg13g2_a21oi_1 _5185_ (.A1(net988),
    .A2(\FpgaPins_Fpga_FSM_data_a1[6] ),
    .Y(_1663_),
    .B1(_1662_));
 sg13g2_a21o_1 _5186_ (.A2(net793),
    .A1(_0123_),
    .B1(_1343_),
    .X(_1664_));
 sg13g2_a21oi_1 _5187_ (.A1(_0743_),
    .A2(_1342_),
    .Y(_1665_),
    .B1(_1347_));
 sg13g2_o21ai_1 _5188_ (.B1(_1665_),
    .Y(_1666_),
    .A1(_1663_),
    .A2(_1664_));
 sg13g2_a221oi_1 _5189_ (.B2(_0123_),
    .C1(net800),
    .B1(_1354_),
    .A1(_0189_),
    .Y(_1667_),
    .A2(net791));
 sg13g2_nor2_1 _5190_ (.A(_1299_),
    .B(_1652_),
    .Y(_1668_));
 sg13g2_a21oi_1 _5191_ (.A1(_1666_),
    .A2(_1667_),
    .Y(_1669_),
    .B1(_1668_));
 sg13g2_a21oi_1 _5192_ (.A1(_1359_),
    .A2(_1655_),
    .Y(_1670_),
    .B1(net782));
 sg13g2_o21ai_1 _5193_ (.B1(_1670_),
    .Y(_1671_),
    .A1(net790),
    .A2(_1669_));
 sg13g2_a21oi_1 _5194_ (.A1(net782),
    .A2(_1654_),
    .Y(_1672_),
    .B1(_1366_));
 sg13g2_a221oi_1 _5195_ (.B2(_1672_),
    .C1(net787),
    .B1(_1671_),
    .A1(net788),
    .Y(_1673_),
    .A2(_1653_));
 sg13g2_nor2_1 _5196_ (.A(net785),
    .B(_1673_),
    .Y(_1674_));
 sg13g2_o21ai_1 _5197_ (.B1(_1674_),
    .Y(_1675_),
    .A1(_1659_),
    .A2(_1661_));
 sg13g2_a21oi_2 _5198_ (.B1(_1656_),
    .Y(_1676_),
    .A2(_1626_),
    .A1(_1602_));
 sg13g2_and3_1 _5199_ (.X(_1677_),
    .A(_1602_),
    .B(_1626_),
    .C(_1656_));
 sg13g2_nor3_1 _5200_ (.A(_1629_),
    .B(_1676_),
    .C(_1677_),
    .Y(_1678_));
 sg13g2_o21ai_1 _5201_ (.B1(_1629_),
    .Y(_1679_),
    .A1(_1676_),
    .A2(_1677_));
 sg13g2_nand3b_1 _5202_ (.B(_1679_),
    .C(_1376_),
    .Y(_1680_),
    .A_N(_1678_));
 sg13g2_a21oi_1 _5203_ (.A1(_1675_),
    .A2(_1680_),
    .Y(_1681_),
    .B1(net780));
 sg13g2_o21ai_1 _5204_ (.B1(_1386_),
    .Y(_1682_),
    .A1(_1383_),
    .A2(_1658_));
 sg13g2_o21ai_1 _5205_ (.B1(net784),
    .Y(_1683_),
    .A1(_1676_),
    .A2(_1677_));
 sg13g2_and2_1 _5206_ (.A(net975),
    .B(_1683_),
    .X(_1684_));
 sg13g2_o21ai_1 _5207_ (.B1(_1684_),
    .Y(_1685_),
    .A1(_1681_),
    .A2(_1682_));
 sg13g2_inv_1 _5208_ (.Y(\FpgaPins_Fpga_LIPSI_acc_a1[6] ),
    .A(_1685_));
 sg13g2_mux4_1 _5209_ (.S0(net806),
    .A0(\datam[9][7] ),
    .A1(\datam[8][7] ),
    .A2(\datam[11][7] ),
    .A3(\datam[10][7] ),
    .S1(net813),
    .X(_1686_));
 sg13g2_a21oi_1 _5210_ (.A1(_0751_),
    .A2(net799),
    .Y(_1687_),
    .B1(net816));
 sg13g2_o21ai_1 _5211_ (.B1(_1687_),
    .Y(_1688_),
    .A1(\datam[12][7] ),
    .A2(net799));
 sg13g2_mux2_1 _5212_ (.A0(\datam[15][7] ),
    .A1(\datam[14][7] ),
    .S(net810),
    .X(_1689_));
 sg13g2_a21oi_1 _5213_ (.A1(net818),
    .A2(_1689_),
    .Y(_1690_),
    .B1(net802));
 sg13g2_a21oi_1 _5214_ (.A1(_1688_),
    .A2(_1690_),
    .Y(_1691_),
    .B1(_1325_));
 sg13g2_o21ai_1 _5215_ (.B1(_1691_),
    .Y(_1692_),
    .A1(net795),
    .A2(_1686_));
 sg13g2_mux4_1 _5216_ (.S0(net804),
    .A0(\datam[1][7] ),
    .A1(\datam[0][7] ),
    .A2(\datam[3][7] ),
    .A3(\datam[2][7] ),
    .S1(net812),
    .X(_1693_));
 sg13g2_mux2_1 _5217_ (.A0(\datam[7][7] ),
    .A1(\datam[6][7] ),
    .S(net811),
    .X(_1694_));
 sg13g2_a21oi_1 _5218_ (.A1(_0750_),
    .A2(net809),
    .Y(_1695_),
    .B1(net815));
 sg13g2_o21ai_1 _5219_ (.B1(_1695_),
    .Y(_1696_),
    .A1(\datam[5][7] ),
    .A2(net809));
 sg13g2_a21oi_1 _5220_ (.A1(net815),
    .A2(_1694_),
    .Y(_1697_),
    .B1(net802));
 sg13g2_nand2_1 _5221_ (.Y(_1698_),
    .A(_1696_),
    .B(_1697_));
 sg13g2_o21ai_1 _5222_ (.B1(_1698_),
    .Y(_1699_),
    .A1(net795),
    .A2(_1693_));
 sg13g2_o21ai_1 _5223_ (.B1(_1692_),
    .Y(\FpgaPins_Fpga_FSM_data_a1[7] ),
    .A1(net794),
    .A2(_1699_));
 sg13g2_a21oi_1 _5224_ (.A1(_1068_),
    .A2(_1076_),
    .Y(_1700_),
    .B1(_0728_));
 sg13g2_a21oi_2 _5225_ (.B1(_1700_),
    .Y(_1701_),
    .A2(\FpgaPins_Fpga_FSM_data_a1[7] ),
    .A1(net981));
 sg13g2_nor2_2 _5226_ (.A(_0731_),
    .B(_1701_),
    .Y(_1702_));
 sg13g2_xnor2_1 _5227_ (.Y(_1703_),
    .A(\FpgaPins_Fpga_LIPSI_acc_a2[7] ),
    .B(_1701_));
 sg13g2_or3_1 _5228_ (.A(_1653_),
    .B(_1676_),
    .C(_1703_),
    .X(_1704_));
 sg13g2_o21ai_1 _5229_ (.B1(_1703_),
    .Y(_1705_),
    .A1(_1653_),
    .A2(_1676_));
 sg13g2_a21oi_1 _5230_ (.A1(_1704_),
    .A2(_1705_),
    .Y(_1706_),
    .B1(_1678_));
 sg13g2_and3_1 _5231_ (.X(_1707_),
    .A(_1678_),
    .B(_1704_),
    .C(_1705_));
 sg13g2_or3_1 _5232_ (.A(_1377_),
    .B(_1706_),
    .C(_1707_),
    .X(_1708_));
 sg13g2_nand2b_1 _5233_ (.Y(_1709_),
    .B(_1702_),
    .A_N(net782));
 sg13g2_a21oi_1 _5234_ (.A1(_0731_),
    .A2(_1701_),
    .Y(_1710_),
    .B1(_1360_));
 sg13g2_or2_1 _5235_ (.X(_1711_),
    .B(\FpgaPins_Fpga_FSM_data_a1[7] ),
    .A(_0699_));
 sg13g2_a21oi_1 _5236_ (.A1(_0699_),
    .A2(_0123_),
    .Y(_1712_),
    .B1(net793));
 sg13g2_a22oi_1 _5237_ (.Y(_1713_),
    .B1(_1711_),
    .B2(_1712_),
    .A2(net793),
    .A1(_0697_));
 sg13g2_a21oi_1 _5238_ (.A1(_0746_),
    .A2(_1343_),
    .Y(_1714_),
    .B1(_1352_));
 sg13g2_o21ai_1 _5239_ (.B1(_1714_),
    .Y(_1715_),
    .A1(_1343_),
    .A2(_1713_));
 sg13g2_a21oi_1 _5240_ (.A1(_0122_),
    .A2(_1347_),
    .Y(_1716_),
    .B1(net791));
 sg13g2_a221oi_1 _5241_ (.B2(_1716_),
    .C1(net800),
    .B1(_1715_),
    .A1(_0746_),
    .Y(_1717_),
    .A2(net791));
 sg13g2_a21oi_1 _5242_ (.A1(_1298_),
    .A2(_1701_),
    .Y(_1718_),
    .B1(_1717_));
 sg13g2_a22oi_1 _5243_ (.Y(_1719_),
    .B1(_1718_),
    .B2(_1360_),
    .A2(_1710_),
    .A1(_1709_));
 sg13g2_a21oi_1 _5244_ (.A1(net789),
    .A2(_1702_),
    .Y(_1720_),
    .B1(net787));
 sg13g2_o21ai_1 _5245_ (.B1(_1720_),
    .Y(_1721_),
    .A1(net789),
    .A2(_1719_));
 sg13g2_and2_1 _5246_ (.A(_1377_),
    .B(_1721_),
    .X(_1722_));
 sg13g2_nand2_1 _5247_ (.Y(_1723_),
    .A(_0746_),
    .B(_1652_));
 sg13g2_o21ai_1 _5248_ (.B1(_1723_),
    .Y(_1724_),
    .A1(_1655_),
    .A2(_1657_));
 sg13g2_nor2b_1 _5249_ (.A(_1703_),
    .B_N(_1724_),
    .Y(_1725_));
 sg13g2_xnor2_1 _5250_ (.Y(_1726_),
    .A(_1703_),
    .B(_1724_));
 sg13g2_nor2_1 _5251_ (.A(_1660_),
    .B(_1726_),
    .Y(_1727_));
 sg13g2_o21ai_1 _5252_ (.B1(_1722_),
    .Y(_1728_),
    .A1(_1374_),
    .A2(_1727_));
 sg13g2_a21oi_1 _5253_ (.A1(_1708_),
    .A2(_1728_),
    .Y(_1729_),
    .B1(net780));
 sg13g2_a21o_1 _5254_ (.A2(_1722_),
    .A1(_1660_),
    .B1(net780),
    .X(_1730_));
 sg13g2_a21o_1 _5255_ (.A2(_1730_),
    .A1(_1726_),
    .B1(net784),
    .X(_1731_));
 sg13g2_a21oi_1 _5256_ (.A1(_1704_),
    .A2(_1705_),
    .Y(_1732_),
    .B1(_1386_));
 sg13g2_nor2_1 _5257_ (.A(net944),
    .B(_1732_),
    .Y(_1733_));
 sg13g2_o21ai_1 _5258_ (.B1(_1733_),
    .Y(_1734_),
    .A1(_1729_),
    .A2(_1731_));
 sg13g2_inv_1 _5259_ (.Y(\FpgaPins_Fpga_LIPSI_acc_a1[7] ),
    .A(_1734_));
 sg13g2_nor2_2 _5260_ (.A(net992),
    .B(\C1.next_state_var[3] ),
    .Y(_1735_));
 sg13g2_inv_1 _5261_ (.Y(_1736_),
    .A(_1735_));
 sg13g2_nor2_1 _5262_ (.A(net995),
    .B(_1736_),
    .Y(_1737_));
 sg13g2_nand2_2 _5263_ (.Y(_1738_),
    .A(_0710_),
    .B(_1735_));
 sg13g2_nand2_2 _5264_ (.Y(_1739_),
    .A(\C1.timer[0] ),
    .B(\C1.counter_status[0] ));
 sg13g2_nor2_2 _5265_ (.A(\C1.timer[1] ),
    .B(_1739_),
    .Y(_1740_));
 sg13g2_nand2b_1 _5266_ (.Y(_1741_),
    .B(_0675_),
    .A_N(_1739_));
 sg13g2_nand2_1 _5267_ (.Y(_1742_),
    .A(\C1.next_state_var[5] ),
    .B(net939));
 sg13g2_nand2_2 _5268_ (.Y(_1743_),
    .A(\C1.temp[1] ),
    .B(\C1.temp[0] ));
 sg13g2_nor2_2 _5269_ (.A(_0669_),
    .B(_1743_),
    .Y(_1744_));
 sg13g2_nand3_1 _5270_ (.B(\C1.temp[1] ),
    .C(\C1.temp[0] ),
    .A(\C1.level[1] ),
    .Y(_1745_));
 sg13g2_a21oi_2 _5271_ (.B1(_1264_),
    .Y(_1746_),
    .A2(_0670_),
    .A1(_0669_));
 sg13g2_nand2_1 _5272_ (.Y(_1747_),
    .A(_1745_),
    .B(_1746_));
 sg13g2_o21ai_1 _5273_ (.B1(net994),
    .Y(_1748_),
    .A1(net939),
    .A2(_1747_));
 sg13g2_and2_2 _5274_ (.A(\C1.timer[1] ),
    .B(\C1.counter_status[0] ),
    .X(_1749_));
 sg13g2_nand2_2 _5275_ (.Y(_1750_),
    .A(\C1.timer[1] ),
    .B(\C1.counter_status[0] ));
 sg13g2_nor3_1 _5276_ (.A(\C1.counter1[6] ),
    .B(\C1.counter1[10] ),
    .C(\C1.counter1[9] ),
    .Y(_1751_));
 sg13g2_nor4_2 _5277_ (.A(\C1.counter1[2] ),
    .B(\C1.counter1[1] ),
    .C(\C1.counter1[0] ),
    .Y(_1752_),
    .D(\C1.counter1[3] ));
 sg13g2_nor4_1 _5278_ (.A(\C1.counter1[5] ),
    .B(\C1.counter1[4] ),
    .C(\C1.counter1[7] ),
    .D(\C1.counter1[8] ),
    .Y(_1753_));
 sg13g2_nand3_1 _5279_ (.B(_1752_),
    .C(_1753_),
    .A(_1751_),
    .Y(_1754_));
 sg13g2_or2_2 _5280_ (.X(_1755_),
    .B(_1754_),
    .A(\C1.counter1[11] ));
 sg13g2_nor3_1 _5281_ (.A(net1545),
    .B(net1689),
    .C(net1734),
    .Y(_1756_));
 sg13g2_nor4_2 _5282_ (.A(net1545),
    .B(\C1.counter2[1] ),
    .C(\C1.counter2[2] ),
    .Y(_1757_),
    .D(\C1.counter2[3] ));
 sg13g2_nor2b_1 _5283_ (.A(net1604),
    .B_N(_1757_),
    .Y(_1758_));
 sg13g2_nor2b_1 _5284_ (.A(\C1.counter2[5] ),
    .B_N(_1758_),
    .Y(_1759_));
 sg13g2_nand3b_1 _5285_ (.B(_0716_),
    .C(_1758_),
    .Y(_1760_),
    .A_N(\C1.counter2[5] ));
 sg13g2_or2_1 _5286_ (.X(_1761_),
    .B(_1760_),
    .A(net1754));
 sg13g2_nor4_2 _5287_ (.A(net1685),
    .B(net1706),
    .C(net1683),
    .Y(_1762_),
    .D(_1760_));
 sg13g2_nand2b_2 _5288_ (.Y(_1763_),
    .B(_1762_),
    .A_N(\C1.counter2[10] ));
 sg13g2_nor3_2 _5289_ (.A(net1681),
    .B(net1712),
    .C(_1763_),
    .Y(_1764_));
 sg13g2_nand2b_2 _5290_ (.Y(_1765_),
    .B(_1764_),
    .A_N(\C1.counter2[13] ));
 sg13g2_nor3_2 _5291_ (.A(net1715),
    .B(net1694),
    .C(_1765_),
    .Y(_1766_));
 sg13g2_nand2b_2 _5292_ (.Y(_1767_),
    .B(_1766_),
    .A_N(\C1.counter2[16] ));
 sg13g2_nor3_2 _5293_ (.A(net1696),
    .B(net1702),
    .C(_1767_),
    .Y(_1768_));
 sg13g2_nand2b_2 _5294_ (.Y(_1769_),
    .B(_1768_),
    .A_N(net1576));
 sg13g2_nor3_2 _5295_ (.A(net1704),
    .B(net1672),
    .C(_1769_),
    .Y(_1770_));
 sg13g2_nand2b_2 _5296_ (.Y(_1771_),
    .B(_1770_),
    .A_N(net1271));
 sg13g2_nor3_2 _5297_ (.A(net1617),
    .B(net1651),
    .C(_1771_),
    .Y(_1772_));
 sg13g2_nand2b_2 _5298_ (.Y(_1773_),
    .B(_1772_),
    .A_N(net1186));
 sg13g2_nor3_2 _5299_ (.A(net1658),
    .B(net1632),
    .C(_1773_),
    .Y(_1774_));
 sg13g2_nand2b_2 _5300_ (.Y(_1775_),
    .B(_1774_),
    .A_N(net1286));
 sg13g2_nor3_1 _5301_ (.A(net1613),
    .B(net1656),
    .C(_1775_),
    .Y(_1776_));
 sg13g2_and2_1 _5302_ (.A(_0717_),
    .B(_1776_),
    .X(_1777_));
 sg13g2_and2_2 _5303_ (.A(_1755_),
    .B(_1777_),
    .X(_1778_));
 sg13g2_nand2_2 _5304_ (.Y(_1779_),
    .A(_1755_),
    .B(_1777_));
 sg13g2_nor3_1 _5305_ (.A(\C1.counter1[1] ),
    .B(\C1.counter1[0] ),
    .C(_1779_),
    .Y(_1780_));
 sg13g2_and2_1 _5306_ (.A(_0712_),
    .B(_1780_),
    .X(_1781_));
 sg13g2_nand2_1 _5307_ (.Y(_1782_),
    .A(_1752_),
    .B(_1778_));
 sg13g2_nand3_1 _5308_ (.B(_1752_),
    .C(_1778_),
    .A(_0713_),
    .Y(_1783_));
 sg13g2_nor2_1 _5309_ (.A(\C1.counter1[5] ),
    .B(_1783_),
    .Y(_1784_));
 sg13g2_nor3_1 _5310_ (.A(\C1.counter1[5] ),
    .B(\C1.counter1[6] ),
    .C(_1783_),
    .Y(_1785_));
 sg13g2_nor4_2 _5311_ (.A(\C1.counter1[5] ),
    .B(\C1.counter1[6] ),
    .C(\C1.counter1[7] ),
    .Y(_1786_),
    .D(_1783_));
 sg13g2_nor2b_1 _5312_ (.A(\C1.counter1[8] ),
    .B_N(_1786_),
    .Y(_1787_));
 sg13g2_and2_1 _5313_ (.A(_0715_),
    .B(_1787_),
    .X(_1788_));
 sg13g2_xnor2_1 _5314_ (.Y(_1789_),
    .A(_0097_),
    .B(_1788_));
 sg13g2_xnor2_1 _5315_ (.Y(_1790_),
    .A(_0676_),
    .B(_1747_));
 sg13g2_o21ai_1 _5316_ (.B1(net939),
    .Y(_1791_),
    .A1(_1750_),
    .A2(_1790_));
 sg13g2_a21oi_1 _5317_ (.A1(_1750_),
    .A2(_1789_),
    .Y(_1792_),
    .B1(_1791_));
 sg13g2_nor2_1 _5318_ (.A(\C1.rinse_status ),
    .B(_1755_),
    .Y(_1793_));
 sg13g2_o21ai_1 _5319_ (.B1(\C1.next_state_var[3] ),
    .Y(_1794_),
    .A1(\C1.rinse_status ),
    .A2(_1755_));
 sg13g2_nor2_1 _5320_ (.A(\C1.dry_status ),
    .B(_1755_),
    .Y(_1795_));
 sg13g2_o21ai_1 _5321_ (.B1(net992),
    .Y(_1796_),
    .A1(\C1.dry_status ),
    .A2(_1755_));
 sg13g2_and2_2 _5322_ (.A(_1794_),
    .B(_1796_),
    .X(_1797_));
 sg13g2_nand2_2 _5323_ (.Y(_1798_),
    .A(_1794_),
    .B(_1796_));
 sg13g2_a21oi_1 _5324_ (.A1(_1789_),
    .A2(_1798_),
    .Y(_1799_),
    .B1(net933));
 sg13g2_o21ai_1 _5325_ (.B1(_1799_),
    .Y(_1800_),
    .A1(_1748_),
    .A2(_1792_));
 sg13g2_o21ai_1 _5326_ (.B1(_1800_),
    .Y(_1801_),
    .A1(net1700),
    .A2(_1738_));
 sg13g2_xnor2_1 _5327_ (.Y(_1802_),
    .A(net1726),
    .B(_1785_));
 sg13g2_nor2_1 _5328_ (.A(_1749_),
    .B(_1802_),
    .Y(_1803_));
 sg13g2_nor2_2 _5329_ (.A(\C1.timer[0] ),
    .B(_1750_),
    .Y(_1804_));
 sg13g2_nand2_2 _5330_ (.Y(_1805_),
    .A(_0676_),
    .B(_1749_));
 sg13g2_nand2_1 _5331_ (.Y(_1806_),
    .A(\C1.level[1] ),
    .B(_0670_));
 sg13g2_nor2_2 _5332_ (.A(\C1.level[0] ),
    .B(_1745_),
    .Y(_1807_));
 sg13g2_nor2_2 _5333_ (.A(\C1.temp[1] ),
    .B(_0672_),
    .Y(_1808_));
 sg13g2_nor3_2 _5334_ (.A(_0669_),
    .B(\C1.temp[1] ),
    .C(_0672_),
    .Y(_1809_));
 sg13g2_nand2_2 _5335_ (.Y(_1810_),
    .A(\C1.level[1] ),
    .B(_1808_));
 sg13g2_nor2_2 _5336_ (.A(_0671_),
    .B(\C1.temp[0] ),
    .Y(_1811_));
 sg13g2_nor2_1 _5337_ (.A(\C1.level[1] ),
    .B(_0670_),
    .Y(_1812_));
 sg13g2_nand2_2 _5338_ (.Y(_1813_),
    .A(_1811_),
    .B(_1812_));
 sg13g2_nand2_1 _5339_ (.Y(_1814_),
    .A(_1810_),
    .B(_1813_));
 sg13g2_o21ai_1 _5340_ (.B1(_1804_),
    .Y(_1815_),
    .A1(_1807_),
    .A2(_1814_));
 sg13g2_nand2_2 _5341_ (.Y(_1816_),
    .A(\C1.timer[0] ),
    .B(_1749_));
 sg13g2_inv_1 _5342_ (.Y(_1817_),
    .A(_1816_));
 sg13g2_nand2_2 _5343_ (.Y(_1818_),
    .A(_1808_),
    .B(_1812_));
 sg13g2_nand3_1 _5344_ (.B(_1813_),
    .C(_1818_),
    .A(_1745_),
    .Y(_1819_));
 sg13g2_nand2_2 _5345_ (.Y(_1820_),
    .A(\C1.level[0] ),
    .B(_1809_));
 sg13g2_nor2b_1 _5346_ (.A(_1819_),
    .B_N(_1820_),
    .Y(_1821_));
 sg13g2_o21ai_1 _5347_ (.B1(_1815_),
    .Y(_1822_),
    .A1(_1816_),
    .A2(_1821_));
 sg13g2_o21ai_1 _5348_ (.B1(net938),
    .Y(_1823_),
    .A1(_1803_),
    .A2(_1822_));
 sg13g2_nor3_2 _5349_ (.A(_0669_),
    .B(_0670_),
    .C(_0671_),
    .Y(_1824_));
 sg13g2_nand2_2 _5350_ (.Y(_1825_),
    .A(_0672_),
    .B(_1824_));
 sg13g2_a21oi_2 _5351_ (.B1(_1807_),
    .Y(_1826_),
    .A2(_1811_),
    .A1(\C1.level[0] ));
 sg13g2_a21o_1 _5352_ (.A2(_1826_),
    .A1(_1810_),
    .B1(net938),
    .X(_1827_));
 sg13g2_nand3_1 _5353_ (.B(_1823_),
    .C(_1827_),
    .A(net994),
    .Y(_1828_));
 sg13g2_a22oi_1 _5354_ (.Y(_1829_),
    .B1(_1798_),
    .B2(_1802_),
    .A2(net934),
    .A1(\C1.counter1[7] ));
 sg13g2_nand2_1 _5355_ (.Y(_1830_),
    .A(_1828_),
    .B(_1829_));
 sg13g2_nor2_1 _5356_ (.A(_0710_),
    .B(_1749_),
    .Y(_1831_));
 sg13g2_nand2_1 _5357_ (.Y(_1832_),
    .A(_1739_),
    .B(_1831_));
 sg13g2_xor2_1 _5358_ (.B(_1787_),
    .A(_0096_),
    .X(_1833_));
 sg13g2_a21oi_1 _5359_ (.A1(_1735_),
    .A2(_1832_),
    .Y(_1834_),
    .B1(_1833_));
 sg13g2_a22oi_1 _5360_ (.Y(_1835_),
    .B1(_1795_),
    .B2(net992),
    .A2(_1793_),
    .A1(\C1.next_state_var[3] ));
 sg13g2_inv_1 _5361_ (.Y(_1836_),
    .A(_1835_));
 sg13g2_a21oi_1 _5362_ (.A1(_1739_),
    .A2(_1750_),
    .Y(_1837_),
    .B1(_0710_));
 sg13g2_nand3_1 _5363_ (.B(\C1.counter_status[0] ),
    .C(_1224_),
    .A(\C1.next_state_var[5] ),
    .Y(_1838_));
 sg13g2_a21oi_1 _5364_ (.A1(_1217_),
    .A2(_1808_),
    .Y(_1839_),
    .B1(_1744_));
 sg13g2_nand2_1 _5365_ (.Y(_1840_),
    .A(net936),
    .B(_1839_));
 sg13g2_nor3_1 _5366_ (.A(net933),
    .B(_1834_),
    .C(_1836_),
    .Y(_1841_));
 sg13g2_a22oi_1 _5367_ (.Y(_1842_),
    .B1(_1840_),
    .B2(_1841_),
    .A2(net933),
    .A1(_0715_));
 sg13g2_o21ai_1 _5368_ (.B1(_1818_),
    .Y(_1843_),
    .A1(\C1.level[0] ),
    .A2(_1810_));
 sg13g2_nand2b_1 _5369_ (.Y(_1844_),
    .B(_1813_),
    .A_N(_1843_));
 sg13g2_o21ai_1 _5370_ (.B1(_1740_),
    .Y(_1845_),
    .A1(_1824_),
    .A2(_1844_));
 sg13g2_nor3_2 _5371_ (.A(\C1.level[1] ),
    .B(_0670_),
    .C(_1743_),
    .Y(_1846_));
 sg13g2_nor3_1 _5372_ (.A(_1805_),
    .B(_1807_),
    .C(_1846_),
    .Y(_1847_));
 sg13g2_nand3_1 _5373_ (.B(_1825_),
    .C(_1847_),
    .A(_1820_),
    .Y(_1848_));
 sg13g2_and4_1 _5374_ (.A(net994),
    .B(_1816_),
    .C(_1845_),
    .D(_1848_),
    .X(_1849_));
 sg13g2_xnor2_1 _5375_ (.Y(_1850_),
    .A(_0093_),
    .B(_1784_));
 sg13g2_o21ai_1 _5376_ (.B1(_1850_),
    .Y(_1851_),
    .A1(_1798_),
    .A2(_1849_));
 sg13g2_nor3_1 _5377_ (.A(_1744_),
    .B(_1804_),
    .C(_1843_),
    .Y(_1852_));
 sg13g2_nand2_1 _5378_ (.Y(_1853_),
    .A(_1825_),
    .B(_1852_));
 sg13g2_a21oi_1 _5379_ (.A1(_1848_),
    .A2(_1853_),
    .Y(_1854_),
    .B1(_1740_));
 sg13g2_nor2_1 _5380_ (.A(_1838_),
    .B(_1854_),
    .Y(_1855_));
 sg13g2_a21oi_1 _5381_ (.A1(_1845_),
    .A2(_1855_),
    .Y(_1856_),
    .B1(net934));
 sg13g2_a22oi_1 _5382_ (.Y(_1857_),
    .B1(_1851_),
    .B2(_1856_),
    .A2(net934),
    .A1(_0714_));
 sg13g2_nand2_1 _5383_ (.Y(_1858_),
    .A(_1217_),
    .B(_1811_));
 sg13g2_and3_1 _5384_ (.X(_1859_),
    .A(_1745_),
    .B(_1804_),
    .C(_1818_));
 sg13g2_o21ai_1 _5385_ (.B1(_1858_),
    .Y(_1860_),
    .A1(_1852_),
    .A2(_1859_));
 sg13g2_a21oi_1 _5386_ (.A1(_1749_),
    .A2(_1860_),
    .Y(_1861_),
    .B1(_1742_));
 sg13g2_nor2b_2 _5387_ (.A(_1806_),
    .B_N(_1811_),
    .Y(_1862_));
 sg13g2_nor3_1 _5388_ (.A(net938),
    .B(_1819_),
    .C(_1862_),
    .Y(_1863_));
 sg13g2_a22oi_1 _5389_ (.Y(_1864_),
    .B1(_1863_),
    .B2(net994),
    .A2(net934),
    .A1(\C1.counter1[8] ));
 sg13g2_a21o_1 _5390_ (.A2(_1859_),
    .A1(_1858_),
    .B1(_1817_),
    .X(_1865_));
 sg13g2_xnor2_1 _5391_ (.Y(_1866_),
    .A(_0095_),
    .B(_1786_));
 sg13g2_o21ai_1 _5392_ (.B1(_1861_),
    .Y(_1867_),
    .A1(_1865_),
    .A2(_1866_));
 sg13g2_nand2_1 _5393_ (.Y(_1868_),
    .A(_1736_),
    .B(_1866_));
 sg13g2_nand4_1 _5394_ (.B(_1864_),
    .C(_1867_),
    .A(_1835_),
    .Y(_1869_),
    .D(_1868_));
 sg13g2_nor2_1 _5395_ (.A(_1754_),
    .B(_1779_),
    .Y(_1870_));
 sg13g2_xnor2_1 _5396_ (.Y(_1871_),
    .A(_0098_),
    .B(_1870_));
 sg13g2_a22oi_1 _5397_ (.Y(_1872_),
    .B1(_1817_),
    .B2(_1746_),
    .A2(_1804_),
    .A1(_1744_));
 sg13g2_o21ai_1 _5398_ (.B1(_1872_),
    .Y(_1873_),
    .A1(_1749_),
    .A2(_1871_));
 sg13g2_nand2_1 _5399_ (.Y(_1874_),
    .A(net938),
    .B(_1873_));
 sg13g2_o21ai_1 _5400_ (.B1(_1746_),
    .Y(_1875_),
    .A1(_1744_),
    .A2(_1805_));
 sg13g2_o21ai_1 _5401_ (.B1(_1874_),
    .Y(_1876_),
    .A1(net938),
    .A2(_1746_));
 sg13g2_a22oi_1 _5402_ (.Y(_1877_),
    .B1(_1798_),
    .B2(_1871_),
    .A2(net934),
    .A1(\C1.counter1[11] ));
 sg13g2_o21ai_1 _5403_ (.B1(_1877_),
    .Y(_1878_),
    .A1(_0710_),
    .A2(_1876_));
 sg13g2_nand2_2 _5404_ (.Y(_1879_),
    .A(\C1.level[0] ),
    .B(_1744_));
 sg13g2_nand2b_2 _5405_ (.Y(_1880_),
    .B(_1879_),
    .A_N(_1844_));
 sg13g2_o21ai_1 _5406_ (.B1(net994),
    .Y(_1881_),
    .A1(net939),
    .A2(_1880_));
 sg13g2_xnor2_1 _5407_ (.Y(_1882_),
    .A(_0676_),
    .B(_1880_));
 sg13g2_o21ai_1 _5408_ (.B1(net939),
    .Y(_1883_),
    .A1(_1750_),
    .A2(_1882_));
 sg13g2_xnor2_1 _5409_ (.Y(_1884_),
    .A(_0090_),
    .B(_1781_));
 sg13g2_a21oi_1 _5410_ (.A1(_1750_),
    .A2(_1884_),
    .Y(_1885_),
    .B1(_1883_));
 sg13g2_a21oi_1 _5411_ (.A1(_1798_),
    .A2(_1884_),
    .Y(_1886_),
    .B1(net933));
 sg13g2_o21ai_1 _5412_ (.B1(_1886_),
    .Y(_1887_),
    .A1(_1881_),
    .A2(_1885_));
 sg13g2_o21ai_1 _5413_ (.B1(_1887_),
    .Y(_1888_),
    .A1(net1740),
    .A2(_1738_));
 sg13g2_o21ai_1 _5414_ (.B1(_1826_),
    .Y(_1889_),
    .A1(\C1.level[0] ),
    .A2(_1810_));
 sg13g2_o21ai_1 _5415_ (.B1(_1831_),
    .Y(_1890_),
    .A1(net939),
    .A2(_1889_));
 sg13g2_xor2_1 _5416_ (.B(_1780_),
    .A(_0089_),
    .X(_1891_));
 sg13g2_a21oi_1 _5417_ (.A1(_1797_),
    .A2(_1890_),
    .Y(_1892_),
    .B1(_1891_));
 sg13g2_nand2_1 _5418_ (.Y(_1893_),
    .A(net936),
    .B(_1889_));
 sg13g2_nor2_1 _5419_ (.A(net933),
    .B(_1892_),
    .Y(_1894_));
 sg13g2_a22oi_1 _5420_ (.Y(_1895_),
    .B1(_1893_),
    .B2(_1894_),
    .A2(net933),
    .A1(_0712_));
 sg13g2_xnor2_1 _5421_ (.Y(_1896_),
    .A(\C1.counter1[1] ),
    .B(\C1.counter1[0] ));
 sg13g2_nor2_2 _5422_ (.A(_1264_),
    .B(_1806_),
    .Y(_1897_));
 sg13g2_o21ai_1 _5423_ (.B1(_1831_),
    .Y(_1898_),
    .A1(net939),
    .A2(_1897_));
 sg13g2_a22oi_1 _5424_ (.Y(_1899_),
    .B1(_1797_),
    .B2(_1898_),
    .A2(_1779_),
    .A1(_0088_));
 sg13g2_o21ai_1 _5425_ (.B1(_1899_),
    .Y(_1900_),
    .A1(_1779_),
    .A2(_1896_));
 sg13g2_nand2_1 _5426_ (.Y(_1901_),
    .A(net936),
    .B(_1897_));
 sg13g2_nand3_1 _5427_ (.B(_1900_),
    .C(_1901_),
    .A(_1738_),
    .Y(_1902_));
 sg13g2_o21ai_1 _5428_ (.B1(_1902_),
    .Y(_1903_),
    .A1(net1748),
    .A2(_1738_));
 sg13g2_nand2_1 _5429_ (.Y(_1904_),
    .A(_1797_),
    .B(_1832_));
 sg13g2_xnor2_1 _5430_ (.Y(_1905_),
    .A(net1665),
    .B(_1778_));
 sg13g2_a22oi_1 _5431_ (.Y(_1906_),
    .B1(_1904_),
    .B2(_1905_),
    .A2(net933),
    .A1(\C1.counter1[0] ));
 sg13g2_nor3_2 _5432_ (.A(_1809_),
    .B(_1824_),
    .C(_1846_),
    .Y(_1907_));
 sg13g2_o21ai_1 _5433_ (.B1(net994),
    .Y(_1908_),
    .A1(net938),
    .A2(_1907_));
 sg13g2_o21ai_1 _5434_ (.B1(_1797_),
    .Y(_1909_),
    .A1(_1749_),
    .A2(_1908_));
 sg13g2_xor2_1 _5435_ (.B(_1782_),
    .A(_0091_),
    .X(_1910_));
 sg13g2_nor2_1 _5436_ (.A(_1816_),
    .B(_1907_),
    .Y(_1911_));
 sg13g2_nor3_2 _5437_ (.A(_0670_),
    .B(_1264_),
    .C(_1744_),
    .Y(_1912_));
 sg13g2_o21ai_1 _5438_ (.B1(net938),
    .Y(_1913_),
    .A1(_1805_),
    .A2(_1912_));
 sg13g2_nor2_1 _5439_ (.A(_1911_),
    .B(_1913_),
    .Y(_1914_));
 sg13g2_o21ai_1 _5440_ (.B1(_1738_),
    .Y(_1915_),
    .A1(_1908_),
    .A2(_1914_));
 sg13g2_a21oi_1 _5441_ (.A1(_1909_),
    .A2(_1910_),
    .Y(_1916_),
    .B1(_1915_));
 sg13g2_a21oi_1 _5442_ (.A1(_0713_),
    .A2(net933),
    .Y(_1917_),
    .B1(_1916_));
 sg13g2_xnor2_1 _5443_ (.Y(_1918_),
    .A(net1743),
    .B(_1783_));
 sg13g2_a21oi_1 _5444_ (.A1(_1735_),
    .A2(_1832_),
    .Y(_1919_),
    .B1(_1918_));
 sg13g2_nand2_1 _5445_ (.Y(_1920_),
    .A(\C1.counter1[5] ),
    .B(net934));
 sg13g2_nand2b_1 _5446_ (.Y(_1921_),
    .B(_1217_),
    .A_N(_1743_));
 sg13g2_nand3_1 _5447_ (.B(_1813_),
    .C(_1921_),
    .A(_1810_),
    .Y(_1922_));
 sg13g2_a21oi_1 _5448_ (.A1(\C1.temp[0] ),
    .A2(_1217_),
    .Y(_1923_),
    .B1(_1805_));
 sg13g2_a221oi_1 _5449_ (.B2(_1740_),
    .C1(_1923_),
    .B1(_1922_),
    .A1(_1817_),
    .Y(_1924_),
    .A2(_1826_));
 sg13g2_o21ai_1 _5450_ (.B1(_1920_),
    .Y(_1925_),
    .A1(_0710_),
    .A2(_1924_));
 sg13g2_nor3_2 _5451_ (.A(_1836_),
    .B(_1919_),
    .C(_1925_),
    .Y(_1926_));
 sg13g2_nand3_1 _5452_ (.B(_1906_),
    .C(_1926_),
    .A(_1903_),
    .Y(_1927_));
 sg13g2_nor4_1 _5453_ (.A(_1830_),
    .B(_1869_),
    .C(_1917_),
    .D(_1927_),
    .Y(_1928_));
 sg13g2_nor4_1 _5454_ (.A(_1842_),
    .B(_1857_),
    .C(_1878_),
    .D(_1895_),
    .Y(_1929_));
 sg13g2_and4_1 _5455_ (.A(_1801_),
    .B(_1888_),
    .C(_1928_),
    .D(_1929_),
    .X(_1930_));
 sg13g2_nand2_1 _5456_ (.Y(_1931_),
    .A(net751),
    .B(_1930_));
 sg13g2_a21oi_1 _5457_ (.A1(net751),
    .A2(_1930_),
    .Y(_0002_),
    .B1(_0000_));
 sg13g2_nor2_1 _5458_ (.A(_0000_),
    .B(_1931_),
    .Y(_0001_));
 sg13g2_nor2_1 _5459_ (.A(\uart_rx_1.r_Rx_Byte[1] ),
    .B(net1674),
    .Y(_1932_));
 sg13g2_or4_1 _5460_ (.A(net1419),
    .B(net1595),
    .C(\uart_rx_1.r_Rx_Byte[3] ),
    .D(net1667),
    .X(_1933_));
 sg13g2_nor4_1 _5461_ (.A(net1352),
    .B(_0665_),
    .C(_0668_),
    .D(_1933_),
    .Y(_1934_));
 sg13g2_nand3_1 _5462_ (.B(_0667_),
    .C(_1932_),
    .A(_0666_),
    .Y(_1935_));
 sg13g2_and2_1 _5463_ (.A(net1675),
    .B(_1934_),
    .X(FpgaPins_Fpga_UART_is_enter_a1));
 sg13g2_nand2_1 _5464_ (.Y(_1936_),
    .A(\uart_rx_1.r_Rx_Byte[1] ),
    .B(\uart_rx_1.r_Rx_Byte[0] ));
 sg13g2_nand2b_1 _5465_ (.Y(_1937_),
    .B(_1936_),
    .A_N(_1932_));
 sg13g2_a21oi_1 _5466_ (.A1(_1934_),
    .A2(_1937_),
    .Y(_1938_),
    .B1(FpgaPins_Fpga_UART_comment_a2));
 sg13g2_and2_1 _5467_ (.A(net2),
    .B(_0795_),
    .X(_1939_));
 sg13g2_nand2_1 _5468_ (.Y(_1940_),
    .A(net2),
    .B(_0795_));
 sg13g2_or3_1 _5469_ (.A(net1543),
    .B(_1938_),
    .C(net950),
    .X(_1941_));
 sg13g2_inv_1 _5470_ (.Y(FpgaPins_Fpga_UART_comment_a1),
    .A(net1544));
 sg13g2_nor4_1 _5471_ (.A(\FpgaPins_Fpga_LIPSI_acc_a1[0] ),
    .B(\FpgaPins_Fpga_LIPSI_acc_a1[1] ),
    .C(\FpgaPins_Fpga_LIPSI_acc_a1[2] ),
    .D(\FpgaPins_Fpga_LIPSI_acc_a1[3] ),
    .Y(_1942_));
 sg13g2_nand2b_1 _5472_ (.Y(_1943_),
    .B(_1942_),
    .A_N(\FpgaPins_Fpga_LIPSI_acc_a1[4] ));
 sg13g2_nor4_1 _5473_ (.A(\FpgaPins_Fpga_LIPSI_acc_a1[5] ),
    .B(\FpgaPins_Fpga_LIPSI_acc_a1[6] ),
    .C(\FpgaPins_Fpga_LIPSI_acc_a1[7] ),
    .D(_1943_),
    .Y(FpgaPins_Fpga_LIPSI_z_a1));
 sg13g2_nor2b_2 _5474_ (.A(net2),
    .B_N(net998),
    .Y(_1944_));
 sg13g2_nand2_1 _5475_ (.Y(FpgaPins_Fpga_GAME_reset_a1),
    .A(net1),
    .B(_1944_));
 sg13g2_nor4_1 _5476_ (.A(_1026_),
    .B(_1043_),
    .C(_1060_),
    .D(_1279_),
    .Y(_1945_));
 sg13g2_and4_1 _5477_ (.A(\FpgaPins_Fpga_FSM_instr_a1[1] ),
    .B(\FpgaPins_Fpga_FSM_instr_a1[0] ),
    .C(\FpgaPins_Fpga_FSM_instr_a1[5] ),
    .D(_1945_),
    .X(FpgaPins_Fpga_LIPSI_exit_a1));
 sg13g2_nor3_1 _5478_ (.A(net875),
    .B(\FpgaPins_Fpga_FSM_instr_a1[4] ),
    .C(_1279_),
    .Y(FpgaPins_Fpga_LIPSI_is_ALU_imm_a1));
 sg13g2_nor3_1 _5479_ (.A(\FpgaPins_Fpga_FSM_instr_a1[1] ),
    .B(net859),
    .C(_1281_),
    .Y(FpgaPins_Fpga_LIPSI_is_br_a1));
 sg13g2_nor3_1 _5480_ (.A(_0850_),
    .B(\FpgaPins_Fpga_FSM_instr_a1[0] ),
    .C(_1281_),
    .Y(FpgaPins_Fpga_LIPSI_is_brz_a1));
 sg13g2_nor2_1 _5481_ (.A(_1281_),
    .B(_1337_),
    .Y(FpgaPins_Fpga_LIPSI_is_brnz_a1));
 sg13g2_nor2_1 _5482_ (.A(_1274_),
    .B(_1281_),
    .Y(_1946_));
 sg13g2_nor2_1 _5483_ (.A(FpgaPins_Fpga_LIPSI_is_ALU_imm_a1),
    .B(_1946_),
    .Y(_1947_));
 sg13g2_nand2_1 _5484_ (.Y(FpgaPins_Fpga_LIPSI_is_2cyc_a1),
    .A(_1286_),
    .B(_1947_));
 sg13g2_nor2_1 _5485_ (.A(net875),
    .B(_1284_),
    .Y(_1948_));
 sg13g2_nor3_1 _5486_ (.A(net875),
    .B(_1060_),
    .C(_1284_),
    .Y(_1949_));
 sg13g2_nor2_1 _5487_ (.A(FpgaPins_Fpga_LIPSI_is_brl_a1),
    .B(\FpgaPins_Fpga_LIPSI_acc_a1[0] ),
    .Y(_1950_));
 sg13g2_nor2_2 _5488_ (.A(FpgaPins_Fpga_LIPSI_is_st_ind_a2),
    .B(_1948_),
    .Y(_1951_));
 sg13g2_or2_1 _5489_ (.X(_1952_),
    .B(_1948_),
    .A(FpgaPins_Fpga_LIPSI_is_st_ind_a2));
 sg13g2_o21ai_1 _5490_ (.B1(_1952_),
    .Y(_1953_),
    .A1(net911),
    .A2(net822));
 sg13g2_nand2_1 _5491_ (.Y(_1954_),
    .A(net1105),
    .B(_1951_));
 sg13g2_o21ai_1 _5492_ (.B1(_1954_),
    .Y(\FpgaPins_Fpga_LIPSI_data_wr_a1[0] ),
    .A1(_1950_),
    .A2(_1953_));
 sg13g2_nor2_1 _5493_ (.A(_0668_),
    .B(FpgaPins_Fpga_UART_comment_a1),
    .Y(_1955_));
 sg13g2_nand2_1 _5494_ (.Y(_1956_),
    .A(\uart_rx_1.r_Rx_DV ),
    .B(_1941_));
 sg13g2_nor2_2 _5495_ (.A(_0191_),
    .B(net902),
    .Y(_1957_));
 sg13g2_nor3_1 _5496_ (.A(\uart_rx_1.r_Rx_Byte[7] ),
    .B(\uart_rx_1.r_Rx_Byte[4] ),
    .C(\uart_rx_1.r_Rx_Byte[3] ),
    .Y(_1958_));
 sg13g2_nand3_1 _5497_ (.B(\uart_rx_1.r_Rx_Byte[1] ),
    .C(\uart_rx_1.r_Rx_Byte[0] ),
    .A(\uart_rx_1.r_Rx_Byte[2] ),
    .Y(_1959_));
 sg13g2_nand4_1 _5498_ (.B(_1935_),
    .C(_1958_),
    .A(\uart_rx_1.r_Rx_Byte[6] ),
    .Y(_1960_),
    .D(_1959_));
 sg13g2_inv_1 _5499_ (.Y(_1961_),
    .A(_1960_));
 sg13g2_and3_1 _5500_ (.X(_1962_),
    .A(FpgaPins_Fpga_UART_first_byte_a2),
    .B(_1955_),
    .C(_1961_));
 sg13g2_nand3_1 _5501_ (.B(_1955_),
    .C(_1961_),
    .A(FpgaPins_Fpga_UART_first_byte_a2),
    .Y(_1963_));
 sg13g2_nor2_2 _5502_ (.A(_1957_),
    .B(_1962_),
    .Y(_1964_));
 sg13g2_mux2_1 _5503_ (.A0(_0192_),
    .A1(\uart_rx_1.r_Rx_Byte[0] ),
    .S(_1960_),
    .X(_1965_));
 sg13g2_mux2_1 _5504_ (.A0(_1965_),
    .A1(\FpgaPins_Fpga_UART_data_a2[0] ),
    .S(_1956_),
    .X(_1966_));
 sg13g2_nand2_1 _5505_ (.Y(_1967_),
    .A(_1964_),
    .B(_1966_));
 sg13g2_inv_1 _5506_ (.Y(\FpgaPins_Fpga_FSM_instr_wr_a1[0] ),
    .A(net874));
 sg13g2_nand2_1 _5507_ (.Y(_1968_),
    .A(net1116),
    .B(_1951_));
 sg13g2_nor2_1 _5508_ (.A(FpgaPins_Fpga_LIPSI_is_brl_a1),
    .B(\FpgaPins_Fpga_LIPSI_acc_a1[1] ),
    .Y(_1969_));
 sg13g2_o21ai_1 _5509_ (.B1(net783),
    .Y(_1970_),
    .A1(net918),
    .A2(net822));
 sg13g2_o21ai_1 _5510_ (.B1(_1968_),
    .Y(\FpgaPins_Fpga_LIPSI_data_wr_a1[1] ),
    .A1(_1969_),
    .A2(_1970_));
 sg13g2_nand2_1 _5511_ (.Y(_1971_),
    .A(\FpgaPins_Fpga_UART_data_a2[1] ),
    .B(net902));
 sg13g2_nor2_1 _5512_ (.A(_1937_),
    .B(_1960_),
    .Y(_1972_));
 sg13g2_a21oi_1 _5513_ (.A1(\uart_rx_1.r_Rx_Byte[1] ),
    .A2(_1960_),
    .Y(_1973_),
    .B1(_1972_));
 sg13g2_o21ai_1 _5514_ (.B1(_1971_),
    .Y(_1974_),
    .A1(net902),
    .A2(_1973_));
 sg13g2_nand2_2 _5515_ (.Y(_1975_),
    .A(_1964_),
    .B(_1974_));
 sg13g2_inv_1 _5516_ (.Y(\FpgaPins_Fpga_FSM_instr_wr_a1[1] ),
    .A(net871));
 sg13g2_nor2_1 _5517_ (.A(FpgaPins_Fpga_LIPSI_is_brl_a1),
    .B(\FpgaPins_Fpga_LIPSI_acc_a1[2] ),
    .Y(_1976_));
 sg13g2_o21ai_1 _5518_ (.B1(net783),
    .Y(_1977_),
    .A1(\FpgaPins_Fpga_FSM_imem_rd_addr_a1[2] ),
    .A2(_1285_));
 sg13g2_nand2_1 _5519_ (.Y(_1978_),
    .A(net1117),
    .B(_1951_));
 sg13g2_o21ai_1 _5520_ (.B1(_1978_),
    .Y(\FpgaPins_Fpga_LIPSI_data_wr_a1[2] ),
    .A1(_1976_),
    .A2(_1977_));
 sg13g2_nand2_1 _5521_ (.Y(_1979_),
    .A(\FpgaPins_Fpga_UART_data_a2[2] ),
    .B(net902));
 sg13g2_nor2_1 _5522_ (.A(_0193_),
    .B(_1936_),
    .Y(_1980_));
 sg13g2_xor2_1 _5523_ (.B(_1936_),
    .A(_0193_),
    .X(_1981_));
 sg13g2_nor2b_1 _5524_ (.A(_1960_),
    .B_N(_1981_),
    .Y(_1982_));
 sg13g2_a21oi_1 _5525_ (.A1(\uart_rx_1.r_Rx_Byte[2] ),
    .A2(_1960_),
    .Y(_1983_),
    .B1(_1982_));
 sg13g2_o21ai_1 _5526_ (.B1(_1979_),
    .Y(_1984_),
    .A1(net902),
    .A2(_1983_));
 sg13g2_nand2_1 _5527_ (.Y(_1985_),
    .A(_1964_),
    .B(_1984_));
 sg13g2_inv_1 _5528_ (.Y(\FpgaPins_Fpga_FSM_instr_wr_a1[2] ),
    .A(net868));
 sg13g2_nor2_1 _5529_ (.A(FpgaPins_Fpga_LIPSI_is_brl_a1),
    .B(\FpgaPins_Fpga_LIPSI_acc_a1[3] ),
    .Y(_1986_));
 sg13g2_o21ai_1 _5530_ (.B1(net783),
    .Y(_1987_),
    .A1(net891),
    .A2(_1285_));
 sg13g2_nand2_1 _5531_ (.Y(_1988_),
    .A(net1130),
    .B(_1951_));
 sg13g2_o21ai_1 _5532_ (.B1(_1988_),
    .Y(\FpgaPins_Fpga_LIPSI_data_wr_a1[3] ),
    .A1(_1986_),
    .A2(_1987_));
 sg13g2_o21ai_1 _5533_ (.B1(_0666_),
    .Y(_1989_),
    .A1(_1960_),
    .A2(_1980_));
 sg13g2_xnor2_1 _5534_ (.Y(_1990_),
    .A(\uart_rx_1.r_Rx_Byte[3] ),
    .B(_1980_));
 sg13g2_mux2_1 _5535_ (.A0(_1989_),
    .A1(\FpgaPins_Fpga_UART_data_a2[3] ),
    .S(net902),
    .X(_1991_));
 sg13g2_nand2_1 _5536_ (.Y(_1992_),
    .A(_1964_),
    .B(_1991_));
 sg13g2_inv_1 _5537_ (.Y(\FpgaPins_Fpga_FSM_instr_wr_a1[3] ),
    .A(net865));
 sg13g2_mux2_1 _5538_ (.A0(\FpgaPins_Fpga_LIPSI_pc_a2[4] ),
    .A1(\FpgaPins_Fpga_LIPSI_data_a2[4] ),
    .S(net990),
    .X(_1993_));
 sg13g2_nand2_1 _5539_ (.Y(_1994_),
    .A(_0833_),
    .B(_1993_));
 sg13g2_o21ai_1 _5540_ (.B1(_0698_),
    .Y(_1995_),
    .A1(_0833_),
    .A2(_1993_));
 sg13g2_nand2b_1 _5541_ (.Y(_1996_),
    .B(_1994_),
    .A_N(_1995_));
 sg13g2_a21oi_1 _5542_ (.A1(net986),
    .A2(_0739_),
    .Y(_1997_),
    .B1(net940));
 sg13g2_a22oi_1 _5543_ (.Y(_1998_),
    .B1(_1996_),
    .B2(_1997_),
    .A2(net940),
    .A1(_0195_));
 sg13g2_nand2_1 _5544_ (.Y(_1999_),
    .A(net1102),
    .B(net942));
 sg13g2_o21ai_1 _5545_ (.B1(_1999_),
    .Y(_2000_),
    .A1(net942),
    .A2(_1998_));
 sg13g2_nor2_1 _5546_ (.A(_0806_),
    .B(net1103),
    .Y(\FpgaPins_Fpga_LIPSI_pc_a1[4] ));
 sg13g2_nor2_1 _5547_ (.A(_1285_),
    .B(\FpgaPins_Fpga_LIPSI_pc_a1[4] ),
    .Y(_2001_));
 sg13g2_o21ai_1 _5548_ (.B1(net783),
    .Y(_2002_),
    .A1(\FpgaPins_Fpga_LIPSI_acc_a1[4] ),
    .A2(_1949_));
 sg13g2_nand2_1 _5549_ (.Y(_2003_),
    .A(net1185),
    .B(_1951_));
 sg13g2_o21ai_1 _5550_ (.B1(_2003_),
    .Y(\FpgaPins_Fpga_LIPSI_data_wr_a1[4] ),
    .A1(_2001_),
    .A2(_2002_));
 sg13g2_a21oi_1 _5551_ (.A1(\uart_rx_1.r_Rx_Byte[0] ),
    .A2(_1957_),
    .Y(_2004_),
    .B1(_1962_));
 sg13g2_o21ai_1 _5552_ (.B1(_2004_),
    .Y(_2005_),
    .A1(_0753_),
    .A2(_1957_));
 sg13g2_o21ai_1 _5553_ (.B1(_2005_),
    .Y(_2006_),
    .A1(_0192_),
    .A2(_1963_));
 sg13g2_inv_1 _5554_ (.Y(\FpgaPins_Fpga_FSM_instr_wr_a1[4] ),
    .A(net856));
 sg13g2_mux2_1 _5555_ (.A0(\FpgaPins_Fpga_LIPSI_pc_a2[5] ),
    .A1(\FpgaPins_Fpga_LIPSI_data_a2[5] ),
    .S(net990),
    .X(_2007_));
 sg13g2_nand3_1 _5556_ (.B(_1993_),
    .C(_2007_),
    .A(_0833_),
    .Y(_2008_));
 sg13g2_a21oi_1 _5557_ (.A1(_0754_),
    .A2(net940),
    .Y(_2009_),
    .B1(net942));
 sg13g2_xnor2_1 _5558_ (.Y(_2010_),
    .A(_1994_),
    .B(_2007_));
 sg13g2_a21oi_1 _5559_ (.A1(net986),
    .A2(_0189_),
    .Y(_2011_),
    .B1(net940));
 sg13g2_o21ai_1 _5560_ (.B1(_2011_),
    .Y(_2012_),
    .A1(net986),
    .A2(_2010_));
 sg13g2_a221oi_1 _5561_ (.B2(_2012_),
    .C1(_0806_),
    .B1(_2009_),
    .A1(net739),
    .Y(\FpgaPins_Fpga_LIPSI_pc_a1[5] ),
    .A2(net942));
 sg13g2_nand2_1 _5562_ (.Y(_2013_),
    .A(net1135),
    .B(_1951_));
 sg13g2_nor2_1 _5563_ (.A(FpgaPins_Fpga_LIPSI_is_brl_a1),
    .B(\FpgaPins_Fpga_LIPSI_acc_a1[5] ),
    .Y(_2014_));
 sg13g2_o21ai_1 _5564_ (.B1(net783),
    .Y(_2015_),
    .A1(net822),
    .A2(\FpgaPins_Fpga_LIPSI_pc_a1[5] ));
 sg13g2_o21ai_1 _5565_ (.B1(_2013_),
    .Y(\FpgaPins_Fpga_LIPSI_data_wr_a1[5] ),
    .A1(_2014_),
    .A2(_2015_));
 sg13g2_mux2_1 _5566_ (.A0(\FpgaPins_Fpga_UART_data_a2[5] ),
    .A1(\uart_rx_1.r_Rx_Byte[1] ),
    .S(_1957_),
    .X(_2016_));
 sg13g2_nor2_1 _5567_ (.A(_1937_),
    .B(_1963_),
    .Y(_2017_));
 sg13g2_a21oi_1 _5568_ (.A1(_1963_),
    .A2(_2016_),
    .Y(_2018_),
    .B1(_2017_));
 sg13g2_inv_1 _5569_ (.Y(\FpgaPins_Fpga_FSM_instr_wr_a1[5] ),
    .A(net862));
 sg13g2_mux2_1 _5570_ (.A0(\FpgaPins_Fpga_LIPSI_pc_a2[6] ),
    .A1(\FpgaPins_Fpga_LIPSI_data_a2[6] ),
    .S(net990),
    .X(_2019_));
 sg13g2_nor2b_1 _5571_ (.A(_2008_),
    .B_N(_2019_),
    .Y(_2020_));
 sg13g2_xnor2_1 _5572_ (.Y(_2021_),
    .A(_2008_),
    .B(_2019_));
 sg13g2_a21oi_1 _5573_ (.A1(net986),
    .A2(_0190_),
    .Y(_2022_),
    .B1(net940));
 sg13g2_o21ai_1 _5574_ (.B1(_2022_),
    .Y(_2023_),
    .A1(net986),
    .A2(_2021_));
 sg13g2_a21oi_1 _5575_ (.A1(_0755_),
    .A2(net940),
    .Y(_2024_),
    .B1(net942));
 sg13g2_a221oi_1 _5576_ (.B2(_2024_),
    .C1(_0806_),
    .B1(_2023_),
    .A1(net717),
    .Y(\FpgaPins_Fpga_LIPSI_pc_a1[6] ),
    .A2(net942));
 sg13g2_o21ai_1 _5577_ (.B1(net783),
    .Y(_2025_),
    .A1(net822),
    .A2(\FpgaPins_Fpga_LIPSI_pc_a1[6] ));
 sg13g2_a21oi_1 _5578_ (.A1(net822),
    .A2(_1685_),
    .Y(_2026_),
    .B1(_2025_));
 sg13g2_a21o_1 _5579_ (.A2(_1951_),
    .A1(net1300),
    .B1(_2026_),
    .X(\FpgaPins_Fpga_LIPSI_data_wr_a1[6] ));
 sg13g2_a21oi_1 _5580_ (.A1(\uart_rx_1.r_Rx_Byte[2] ),
    .A2(_1957_),
    .Y(_2027_),
    .B1(_1962_));
 sg13g2_o21ai_1 _5581_ (.B1(_2027_),
    .Y(_2028_),
    .A1(_0756_),
    .A2(_1957_));
 sg13g2_o21ai_1 _5582_ (.B1(_2028_),
    .Y(_2029_),
    .A1(_1963_),
    .A2(_1981_));
 sg13g2_inv_1 _5583_ (.Y(\FpgaPins_Fpga_FSM_instr_wr_a1[6] ),
    .A(net853));
 sg13g2_nor2b_1 _5584_ (.A(net990),
    .B_N(\FpgaPins_Fpga_LIPSI_pc_a2[7] ),
    .Y(_2030_));
 sg13g2_a21oi_1 _5585_ (.A1(net990),
    .A2(\FpgaPins_Fpga_LIPSI_data_a2[7] ),
    .Y(_2031_),
    .B1(_2030_));
 sg13g2_xnor2_1 _5586_ (.Y(_2032_),
    .A(_2020_),
    .B(_2031_));
 sg13g2_a21oi_1 _5587_ (.A1(net986),
    .A2(_0123_),
    .Y(_2033_),
    .B1(net940));
 sg13g2_o21ai_1 _5588_ (.B1(_2033_),
    .Y(_2034_),
    .A1(net986),
    .A2(_2032_));
 sg13g2_a21oi_1 _5589_ (.A1(_0757_),
    .A2(net941),
    .Y(_2035_),
    .B1(net942));
 sg13g2_a221oi_1 _5590_ (.B2(_2035_),
    .C1(_0806_),
    .B1(_2034_),
    .A1(net735),
    .Y(\FpgaPins_Fpga_LIPSI_pc_a1[7] ),
    .A2(net942));
 sg13g2_o21ai_1 _5591_ (.B1(net783),
    .Y(_2036_),
    .A1(net822),
    .A2(\FpgaPins_Fpga_LIPSI_pc_a1[7] ));
 sg13g2_a21oi_1 _5592_ (.A1(net822),
    .A2(_1734_),
    .Y(_2037_),
    .B1(_2036_));
 sg13g2_a21o_1 _5593_ (.A2(_1951_),
    .A1(net1282),
    .B1(_2037_),
    .X(\FpgaPins_Fpga_LIPSI_data_wr_a1[7] ));
 sg13g2_o21ai_1 _5594_ (.B1(_1963_),
    .Y(_2038_),
    .A1(\FpgaPins_Fpga_UART_data_a2[7] ),
    .A2(_1957_));
 sg13g2_a21oi_1 _5595_ (.A1(_0666_),
    .A2(_1957_),
    .Y(_2039_),
    .B1(_2038_));
 sg13g2_a21oi_1 _5596_ (.A1(_1962_),
    .A2(_1990_),
    .Y(_2040_),
    .B1(_2039_));
 sg13g2_inv_1 _5597_ (.Y(\FpgaPins_Fpga_FSM_instr_wr_a1[7] ),
    .A(net852));
 sg13g2_o21ai_1 _5598_ (.B1(net999),
    .Y(_2041_),
    .A1(_1582_),
    .A2(_1583_));
 sg13g2_a21o_1 _5599_ (.A2(net975),
    .A1(net999),
    .B1(\FpgaPins_Fpga_LIPSI_acc_a1[0] ),
    .X(_2042_));
 sg13g2_nor2_1 _5600_ (.A(net1002),
    .B(\FpgaPins_Fpga_FSM_instr_wr_a1[0] ),
    .Y(_2043_));
 sg13g2_a21oi_1 _5601_ (.A1(net1002),
    .A2(net856),
    .Y(_2044_),
    .B1(_2043_));
 sg13g2_a22oi_1 _5602_ (.Y(_2045_),
    .B1(_2044_),
    .B2(net944),
    .A2(_2042_),
    .A1(_2041_));
 sg13g2_nand2b_1 _5603_ (.Y(_2046_),
    .B(net999),
    .A_N(\FpgaPins_Fpga_LIPSI_acc_a1[5] ));
 sg13g2_a21o_1 _5604_ (.A2(net975),
    .A1(net999),
    .B1(\FpgaPins_Fpga_LIPSI_acc_a1[1] ),
    .X(_2047_));
 sg13g2_nand2_1 _5605_ (.Y(_2048_),
    .A(net1000),
    .B(net862));
 sg13g2_a21oi_1 _5606_ (.A1(net997),
    .A2(net871),
    .Y(_2049_),
    .B1(net975));
 sg13g2_a22oi_1 _5607_ (.Y(_2050_),
    .B1(_2048_),
    .B2(_2049_),
    .A2(_2047_),
    .A1(_2046_));
 sg13g2_nor2b_2 _5608_ (.A(_2045_),
    .B_N(_2050_),
    .Y(_2051_));
 sg13g2_a21oi_1 _5609_ (.A1(net999),
    .A2(net975),
    .Y(_2052_),
    .B1(\FpgaPins_Fpga_LIPSI_acc_a1[3] ));
 sg13g2_a21oi_2 _5610_ (.B1(_2052_),
    .Y(_2053_),
    .A2(_1734_),
    .A1(net1000));
 sg13g2_a21o_1 _5611_ (.A2(_1734_),
    .A1(net1000),
    .B1(_2052_),
    .X(_2054_));
 sg13g2_nor2_1 _5612_ (.A(net1002),
    .B(\FpgaPins_Fpga_FSM_instr_wr_a1[3] ),
    .Y(_2055_));
 sg13g2_a21oi_1 _5613_ (.A1(net1002),
    .A2(net852),
    .Y(_2056_),
    .B1(_2055_));
 sg13g2_and2_1 _5614_ (.A(net944),
    .B(_2056_),
    .X(_2057_));
 sg13g2_nand2_1 _5615_ (.Y(_2058_),
    .A(net944),
    .B(_2056_));
 sg13g2_nor2_1 _5616_ (.A(_2053_),
    .B(_2057_),
    .Y(_2059_));
 sg13g2_nand2_1 _5617_ (.Y(_2060_),
    .A(net999),
    .B(_1685_));
 sg13g2_a21o_1 _5618_ (.A2(net975),
    .A1(net999),
    .B1(\FpgaPins_Fpga_LIPSI_acc_a1[2] ),
    .X(_2061_));
 sg13g2_o21ai_1 _5619_ (.B1(net945),
    .Y(_2062_),
    .A1(net1002),
    .A2(\FpgaPins_Fpga_FSM_instr_wr_a1[2] ));
 sg13g2_a21oi_2 _5620_ (.B1(_2062_),
    .Y(_2063_),
    .A2(net853),
    .A1(net1002));
 sg13g2_a21oi_2 _5621_ (.B1(_2063_),
    .Y(_2064_),
    .A2(_2061_),
    .A1(_2060_));
 sg13g2_a21o_1 _5622_ (.A2(_2061_),
    .A1(_2060_),
    .B1(_2063_),
    .X(_2065_));
 sg13g2_a21oi_1 _5623_ (.A1(_2054_),
    .A2(_2058_),
    .Y(_2066_),
    .B1(_2065_));
 sg13g2_a21oi_2 _5624_ (.B1(_2064_),
    .Y(_2067_),
    .A2(_2058_),
    .A1(_2054_));
 sg13g2_nor3_2 _5625_ (.A(_2053_),
    .B(_2057_),
    .C(_2065_),
    .Y(_2068_));
 sg13g2_nand2_1 _5626_ (.Y(_2069_),
    .A(_2059_),
    .B(_2064_));
 sg13g2_or2_1 _5627_ (.X(_2070_),
    .B(_2068_),
    .A(_2067_));
 sg13g2_and2_1 _5628_ (.A(_2045_),
    .B(_2050_),
    .X(_2071_));
 sg13g2_or2_1 _5629_ (.X(_2072_),
    .B(_2050_),
    .A(_2045_));
 sg13g2_inv_1 _5630_ (.Y(_2073_),
    .A(_2072_));
 sg13g2_and3_1 _5631_ (.X(_2074_),
    .A(_2054_),
    .B(_2058_),
    .C(_2071_));
 sg13g2_a21o_1 _5632_ (.A2(_2073_),
    .A1(_2064_),
    .B1(_2074_),
    .X(_2075_));
 sg13g2_nand2_1 _5633_ (.Y(_2076_),
    .A(_2051_),
    .B(_2064_));
 sg13g2_a221oi_1 _5634_ (.B2(_2069_),
    .C1(net998),
    .B1(_2075_),
    .A1(_2051_),
    .Y(_2077_),
    .A2(_2070_));
 sg13g2_a22oi_1 _5635_ (.Y(_2078_),
    .B1(_1944_),
    .B2(\FpgaPins_Fpga_GAME_led_output_a1[0] ),
    .A2(_1186_),
    .A1(\C1.dura_op ));
 sg13g2_nand2b_2 _5636_ (.Y(uo_out[0]),
    .B(_2078_),
    .A_N(_2077_));
 sg13g2_nor4_1 _5637_ (.A(_2053_),
    .B(_2057_),
    .C(_2064_),
    .D(_2072_),
    .Y(_2079_));
 sg13g2_a21oi_1 _5638_ (.A1(_2051_),
    .A2(_2067_),
    .Y(_2080_),
    .B1(_2079_));
 sg13g2_nand2_1 _5639_ (.Y(_2081_),
    .A(_2066_),
    .B(_2072_));
 sg13g2_nor2_1 _5640_ (.A(_2068_),
    .B(_2074_),
    .Y(_2082_));
 sg13g2_and3_1 _5641_ (.X(_2083_),
    .A(_2080_),
    .B(_2081_),
    .C(_2082_));
 sg13g2_a22oi_1 _5642_ (.Y(_2084_),
    .B1(_1944_),
    .B2(\FpgaPins_Fpga_GAME_led_output_a1[1] ),
    .A2(net996),
    .A1(\C1.temp_op ));
 sg13g2_o21ai_1 _5643_ (.B1(_2084_),
    .Y(uo_out[1]),
    .A1(net998),
    .A2(_2083_));
 sg13g2_nor2b_1 _5644_ (.A(_2051_),
    .B_N(_2067_),
    .Y(_2085_));
 sg13g2_nor2b_1 _5645_ (.A(_2050_),
    .B_N(_2045_),
    .Y(_2086_));
 sg13g2_a21o_1 _5646_ (.A2(_2086_),
    .A1(_2068_),
    .B1(_2085_),
    .X(_2087_));
 sg13g2_a22oi_1 _5647_ (.Y(_2088_),
    .B1(_1944_),
    .B2(\FpgaPins_Fpga_GAME_led_output_a1[2] ),
    .A2(net996),
    .A1(\C1.level_op ));
 sg13g2_o21ai_1 _5648_ (.B1(_2088_),
    .Y(uo_out[2]),
    .A1(net998),
    .A2(_2087_));
 sg13g2_a21oi_1 _5649_ (.A1(_2051_),
    .A2(_2068_),
    .Y(_2089_),
    .B1(_1944_));
 sg13g2_nor2_1 _5650_ (.A(_2065_),
    .B(_2086_),
    .Y(_2090_));
 sg13g2_nor3_1 _5651_ (.A(_2066_),
    .B(_2073_),
    .C(_2074_),
    .Y(_2091_));
 sg13g2_o21ai_1 _5652_ (.B1(_2089_),
    .Y(_2092_),
    .A1(_2090_),
    .A2(_2091_));
 sg13g2_o21ai_1 _5653_ (.B1(net998),
    .Y(_2093_),
    .A1(net2),
    .A2(\FpgaPins_Fpga_GAME_led_output_a1[3] ));
 sg13g2_a22oi_1 _5654_ (.Y(uo_out[3]),
    .B1(_2092_),
    .B2(_2093_),
    .A2(net996),
    .A1(_0680_));
 sg13g2_nand2_1 _5655_ (.Y(_2094_),
    .A(_2045_),
    .B(_2064_));
 sg13g2_nand2_1 _5656_ (.Y(_2095_),
    .A(_2059_),
    .B(_2094_));
 sg13g2_a21oi_1 _5657_ (.A1(_2076_),
    .A2(_2095_),
    .Y(_2096_),
    .B1(_2086_));
 sg13g2_a22oi_1 _5658_ (.Y(_2097_),
    .B1(_1944_),
    .B2(\FpgaPins_Fpga_GAME_led_output_a1[4] ),
    .A2(_1186_),
    .A1(\C1.waiting ));
 sg13g2_o21ai_1 _5659_ (.B1(_2097_),
    .Y(uo_out[4]),
    .A1(net998),
    .A2(_2096_));
 sg13g2_a22oi_1 _5660_ (.Y(_2098_),
    .B1(_2080_),
    .B2(_2069_),
    .A2(_2074_),
    .A1(_2064_));
 sg13g2_a22oi_1 _5661_ (.Y(_2099_),
    .B1(_1944_),
    .B2(\FpgaPins_Fpga_GAME_led_output_a1[5] ),
    .A2(net996),
    .A1(\C1.pouring ));
 sg13g2_o21ai_1 _5662_ (.B1(_2099_),
    .Y(uo_out[5]),
    .A1(net998),
    .A2(_2098_));
 sg13g2_o21ai_1 _5663_ (.B1(_2071_),
    .Y(_2100_),
    .A1(_2067_),
    .A2(_2068_));
 sg13g2_nand3b_1 _5664_ (.B(_2089_),
    .C(_2100_),
    .Y(_2101_),
    .A_N(_2079_));
 sg13g2_o21ai_1 _5665_ (.B1(net998),
    .Y(_2102_),
    .A1(net2),
    .A2(\FpgaPins_Fpga_GAME_led_output_a1[6] ));
 sg13g2_a22oi_1 _5666_ (.Y(uo_out[6]),
    .B1(_2101_),
    .B2(_2102_),
    .A2(net996),
    .A1(_0711_));
 sg13g2_a22oi_1 _5667_ (.Y(_2103_),
    .B1(_1944_),
    .B2(\FpgaPins_Fpga_GAME_led_output_a1[7] ),
    .A2(net996),
    .A1(\C1.heating ));
 sg13g2_inv_1 _5668_ (.Y(\L1_Digit[0].L2_Leds[7].L2_viz_lit_a0 ),
    .A(_2103_));
 sg13g2_nor3_1 _5669_ (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[5] ),
    .B(_0883_),
    .C(_0884_),
    .Y(_2104_));
 sg13g2_and4_1 _5670_ (.A(\FpgaPins_Fpga_GAME_count_speed4_a1[15] ),
    .B(\FpgaPins_Fpga_GAME_count_speed4_a1[5] ),
    .C(_1104_),
    .D(_2104_),
    .X(_2105_));
 sg13g2_o21ai_1 _5671_ (.B1(net985),
    .Y(_2106_),
    .A1(net1313),
    .A2(_2105_));
 sg13g2_a21oi_2 _5672_ (.B1(_2106_),
    .Y(FpgaPins_Fpga_GAME_clk_pulse4_a1),
    .A2(_2105_),
    .A1(net1313));
 sg13g2_and2_1 _5673_ (.A(_0903_),
    .B(_0916_),
    .X(_2107_));
 sg13g2_nand3b_1 _5674_ (.B(_2107_),
    .C(\FpgaPins_Fpga_GAME_count_speed3_a1[7] ),
    .Y(_2108_),
    .A_N(\FpgaPins_Fpga_GAME_count_speed3_a1[6] ));
 sg13g2_nor4_2 _5675_ (.A(_0924_),
    .B(_0925_),
    .C(\FpgaPins_Fpga_GAME_count_speed3_a1[14] ),
    .Y(_2109_),
    .D(_2108_));
 sg13g2_o21ai_1 _5676_ (.B1(_0017_),
    .Y(_2110_),
    .A1(net1159),
    .A2(_2109_));
 sg13g2_a21oi_1 _5677_ (.A1(net1159),
    .A2(_2109_),
    .Y(FpgaPins_Fpga_GAME_clk_pulse3_a1),
    .B1(_2110_));
 sg13g2_nor3_1 _5678_ (.A(_0943_),
    .B(_0958_),
    .C(\FpgaPins_Fpga_GAME_count_speed2_a1[6] ),
    .Y(_2111_));
 sg13g2_nand4_1 _5679_ (.B(\FpgaPins_Fpga_GAME_count_speed2_a1[14] ),
    .C(\FpgaPins_Fpga_GAME_count_speed2_a1[7] ),
    .A(\FpgaPins_Fpga_GAME_count_speed2_a1[15] ),
    .Y(_2112_),
    .D(_2111_));
 sg13g2_o21ai_1 _5680_ (.B1(_0017_),
    .Y(_2113_),
    .A1(_0758_),
    .A2(_2112_));
 sg13g2_a21oi_1 _5681_ (.A1(_0758_),
    .A2(_2112_),
    .Y(FpgaPins_Fpga_GAME_clk_pulse2_a1),
    .B1(_2113_));
 sg13g2_nor3_2 _5682_ (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[7] ),
    .B(_0778_),
    .C(_0794_),
    .Y(_2114_));
 sg13g2_o21ai_1 _5683_ (.B1(_0017_),
    .Y(_2115_),
    .A1(_0695_),
    .A2(_2114_));
 sg13g2_a21oi_1 _5684_ (.A1(_0695_),
    .A2(_2114_),
    .Y(FpgaPins_Fpga_GAME_clk_pulse1_a1),
    .B1(_2115_));
 sg13g2_nand2b_1 _5685_ (.Y(_2116_),
    .B(_0012_),
    .A_N(_0011_));
 sg13g2_a21oi_1 _5686_ (.A1(_0012_),
    .A2(_0011_),
    .Y(_2117_),
    .B1(_0013_));
 sg13g2_nand2b_1 _5687_ (.Y(_2118_),
    .B(FpgaPins_Fpga_GAME_clk_pulse1_a1),
    .A_N(_0011_));
 sg13g2_a21oi_1 _5688_ (.A1(_0011_),
    .A2(FpgaPins_Fpga_GAME_clk_pulse3_a1),
    .Y(_2119_),
    .B1(_0012_));
 sg13g2_nand2_1 _5689_ (.Y(_2120_),
    .A(_2118_),
    .B(_2119_));
 sg13g2_o21ai_1 _5690_ (.B1(_2120_),
    .Y(_2121_),
    .A1(FpgaPins_Fpga_GAME_clk_pulse2_a1),
    .A2(_2116_));
 sg13g2_nor2_1 _5691_ (.A(FpgaPins_Fpga_GAME_clk_pulse4_a1),
    .B(_2117_),
    .Y(_2122_));
 sg13g2_a21oi_1 _5692_ (.A1(_1257_),
    .A2(_2121_),
    .Y(FpgaPins_Fpga_GAME_clk_pulse_a1),
    .B1(_2122_));
 sg13g2_nor2_2 _5693_ (.A(_0711_),
    .B(net1707),
    .Y(_2123_));
 sg13g2_nand2_1 _5694_ (.Y(_2124_),
    .A(net995),
    .B(_2123_));
 sg13g2_nor2_1 _5695_ (.A(_1749_),
    .B(_1778_),
    .Y(_2125_));
 sg13g2_nor2b_1 _5696_ (.A(\C1.counter1[10] ),
    .B_N(\C1.max_count[10] ),
    .Y(_2126_));
 sg13g2_nand2b_1 _5697_ (.Y(_2127_),
    .B(\C1.counter1[10] ),
    .A_N(\C1.max_count[10] ));
 sg13g2_nand2b_1 _5698_ (.Y(_2128_),
    .B(_2127_),
    .A_N(_2126_));
 sg13g2_nor2b_1 _5699_ (.A(\C1.counter1[8] ),
    .B_N(\C1.max_count[8] ),
    .Y(_2129_));
 sg13g2_nand2b_1 _5700_ (.Y(_2130_),
    .B(\C1.max_count[7] ),
    .A_N(\C1.counter1[7] ));
 sg13g2_xor2_1 _5701_ (.B(\C1.counter1[7] ),
    .A(\C1.max_count[7] ),
    .X(_2131_));
 sg13g2_nor2b_1 _5702_ (.A(\C1.counter1[6] ),
    .B_N(\C1.max_count[6] ),
    .Y(_2132_));
 sg13g2_xnor2_1 _5703_ (.Y(_2133_),
    .A(\C1.max_count[6] ),
    .B(\C1.counter1[6] ));
 sg13g2_nand2b_1 _5704_ (.Y(_2134_),
    .B(\C1.max_count[5] ),
    .A_N(\C1.counter1[5] ));
 sg13g2_xor2_1 _5705_ (.B(\C1.counter1[5] ),
    .A(\C1.max_count[5] ),
    .X(_2135_));
 sg13g2_nor2b_1 _5706_ (.A(\C1.counter1[4] ),
    .B_N(\C1.max_count[4] ),
    .Y(_2136_));
 sg13g2_xnor2_1 _5707_ (.Y(_2137_),
    .A(\C1.max_count[3] ),
    .B(\C1.counter1[3] ));
 sg13g2_nand2b_1 _5708_ (.Y(_2138_),
    .B(\C1.counter1[1] ),
    .A_N(\C1.max_count[1] ));
 sg13g2_nor2b_1 _5709_ (.A(\C1.counter1[1] ),
    .B_N(\C1.max_count[1] ),
    .Y(_2139_));
 sg13g2_o21ai_1 _5710_ (.B1(_2138_),
    .Y(_2140_),
    .A1(_0085_),
    .A2(_2139_));
 sg13g2_xnor2_1 _5711_ (.Y(_2141_),
    .A(\C1.max_count[2] ),
    .B(\C1.counter1[2] ));
 sg13g2_nor2b_1 _5712_ (.A(_2140_),
    .B_N(_2141_),
    .Y(_2142_));
 sg13g2_a21oi_1 _5713_ (.A1(\C1.max_count[2] ),
    .A2(_0712_),
    .Y(_2143_),
    .B1(_2142_));
 sg13g2_nand2b_1 _5714_ (.Y(_2144_),
    .B(_2137_),
    .A_N(_2143_));
 sg13g2_o21ai_1 _5715_ (.B1(_2144_),
    .Y(_2145_),
    .A1(_0690_),
    .A2(\C1.counter1[3] ));
 sg13g2_nand2b_1 _5716_ (.Y(_2146_),
    .B(\C1.counter1[4] ),
    .A_N(\C1.max_count[4] ));
 sg13g2_nand2b_1 _5717_ (.Y(_2147_),
    .B(_2146_),
    .A_N(_2136_));
 sg13g2_a21oi_1 _5718_ (.A1(_2145_),
    .A2(_2146_),
    .Y(_2148_),
    .B1(_2136_));
 sg13g2_o21ai_1 _5719_ (.B1(_2134_),
    .Y(_2149_),
    .A1(_2135_),
    .A2(_2148_));
 sg13g2_a21oi_1 _5720_ (.A1(_2133_),
    .A2(_2149_),
    .Y(_2150_),
    .B1(_2132_));
 sg13g2_o21ai_1 _5721_ (.B1(_2130_),
    .Y(_2151_),
    .A1(_2131_),
    .A2(_2150_));
 sg13g2_xnor2_1 _5722_ (.Y(_2152_),
    .A(\C1.max_count[8] ),
    .B(\C1.counter1[8] ));
 sg13g2_a21oi_1 _5723_ (.A1(_2151_),
    .A2(_2152_),
    .Y(_2153_),
    .B1(_2129_));
 sg13g2_xnor2_1 _5724_ (.Y(_2154_),
    .A(\C1.max_count[9] ),
    .B(\C1.counter1[9] ));
 sg13g2_nand2b_1 _5725_ (.Y(_2155_),
    .B(_2154_),
    .A_N(_2153_));
 sg13g2_o21ai_1 _5726_ (.B1(_2155_),
    .Y(_2156_),
    .A1(_0689_),
    .A2(\C1.counter1[9] ));
 sg13g2_xnor2_1 _5727_ (.Y(_2157_),
    .A(_2128_),
    .B(_2156_));
 sg13g2_a21oi_1 _5728_ (.A1(_2127_),
    .A2(_2156_),
    .Y(_2158_),
    .B1(_2126_));
 sg13g2_xor2_1 _5729_ (.B(\C1.counter1[11] ),
    .A(\C1.max_count[11] ),
    .X(_2159_));
 sg13g2_xnor2_1 _5730_ (.Y(_2160_),
    .A(_2158_),
    .B(_2159_));
 sg13g2_nor2b_2 _5731_ (.A(_2157_),
    .B_N(_2160_),
    .Y(_2161_));
 sg13g2_nand2b_1 _5732_ (.Y(_2162_),
    .B(_2160_),
    .A_N(_2157_));
 sg13g2_xnor2_1 _5733_ (.Y(_2163_),
    .A(_2131_),
    .B(_2150_));
 sg13g2_xor2_1 _5734_ (.B(_2149_),
    .A(_2133_),
    .X(_2164_));
 sg13g2_xnor2_1 _5735_ (.Y(_2165_),
    .A(_2133_),
    .B(_2149_));
 sg13g2_xnor2_1 _5736_ (.Y(_2166_),
    .A(_2135_),
    .B(_2148_));
 sg13g2_xnor2_1 _5737_ (.Y(_2167_),
    .A(_2145_),
    .B(_2147_));
 sg13g2_xor2_1 _5738_ (.B(_2147_),
    .A(_2145_),
    .X(_2168_));
 sg13g2_xnor2_1 _5739_ (.Y(_2169_),
    .A(_2140_),
    .B(_2141_));
 sg13g2_xnor2_1 _5740_ (.Y(_2170_),
    .A(_2137_),
    .B(_2143_));
 sg13g2_nor2_1 _5741_ (.A(_2169_),
    .B(_2170_),
    .Y(_2171_));
 sg13g2_xnor2_1 _5742_ (.Y(_2172_),
    .A(\C1.max_count[1] ),
    .B(\C1.counter1[1] ));
 sg13g2_nor2b_1 _5743_ (.A(\C1.counter1[0] ),
    .B_N(_2172_),
    .Y(_2173_));
 sg13g2_nand2b_1 _5744_ (.Y(_2174_),
    .B(_2172_),
    .A_N(\C1.counter1[0] ));
 sg13g2_nor3_1 _5745_ (.A(_2169_),
    .B(_2170_),
    .C(_2174_),
    .Y(_2175_));
 sg13g2_and2_1 _5746_ (.A(_2166_),
    .B(_2168_),
    .X(_2176_));
 sg13g2_o21ai_1 _5747_ (.B1(net880),
    .Y(_2177_),
    .A1(_2168_),
    .A2(_2175_));
 sg13g2_inv_1 _5748_ (.Y(_2178_),
    .A(_2177_));
 sg13g2_xnor2_1 _5749_ (.Y(_2179_),
    .A(_2153_),
    .B(_2154_));
 sg13g2_xor2_1 _5750_ (.B(_2152_),
    .A(_2151_),
    .X(_2180_));
 sg13g2_nor2_1 _5751_ (.A(_2179_),
    .B(_2180_),
    .Y(_2181_));
 sg13g2_and2_1 _5752_ (.A(_2160_),
    .B(_2181_),
    .X(_2182_));
 sg13g2_and4_1 _5753_ (.A(net849),
    .B(_2165_),
    .C(_2178_),
    .D(_2182_),
    .X(_2183_));
 sg13g2_o21ai_1 _5754_ (.B1(_1846_),
    .Y(_2184_),
    .A1(_2161_),
    .A2(_2183_));
 sg13g2_nand2_1 _5755_ (.Y(_2185_),
    .A(net880),
    .B(_2167_));
 sg13g2_nand2_1 _5756_ (.Y(_2186_),
    .A(_2169_),
    .B(_2170_));
 sg13g2_o21ai_1 _5757_ (.B1(_2170_),
    .Y(_2187_),
    .A1(_2169_),
    .A2(_2174_));
 sg13g2_nand3_1 _5758_ (.B(_2167_),
    .C(_2187_),
    .A(net880),
    .Y(_2188_));
 sg13g2_nor2_1 _5759_ (.A(_2165_),
    .B(_2176_),
    .Y(_2189_));
 sg13g2_nand3b_1 _5760_ (.B(_2188_),
    .C(_2189_),
    .Y(_2190_),
    .A_N(net849));
 sg13g2_nand3_1 _5761_ (.B(_2182_),
    .C(_2190_),
    .A(_2157_),
    .Y(_2191_));
 sg13g2_nand2_1 _5762_ (.Y(_2192_),
    .A(_2162_),
    .B(_2191_));
 sg13g2_a21oi_1 _5763_ (.A1(_2165_),
    .A2(net880),
    .Y(_2193_),
    .B1(net849));
 sg13g2_nor2_1 _5764_ (.A(net880),
    .B(_2167_),
    .Y(_2194_));
 sg13g2_nand2_1 _5765_ (.Y(_2195_),
    .A(\C1.counter1[0] ),
    .B(_2172_));
 sg13g2_nand3_1 _5766_ (.B(_2169_),
    .C(_2172_),
    .A(\C1.counter1[0] ),
    .Y(_2196_));
 sg13g2_nand3_1 _5767_ (.B(_2194_),
    .C(_2196_),
    .A(_2165_),
    .Y(_2197_));
 sg13g2_o21ai_1 _5768_ (.B1(_2193_),
    .Y(_2198_),
    .A1(_2170_),
    .A2(_2197_));
 sg13g2_a21oi_1 _5769_ (.A1(_2182_),
    .A2(_2198_),
    .Y(_2199_),
    .B1(_2161_));
 sg13g2_a21oi_1 _5770_ (.A1(_1807_),
    .A2(_2199_),
    .Y(_2200_),
    .B1(_1846_));
 sg13g2_o21ai_1 _5771_ (.B1(_2200_),
    .Y(_2201_),
    .A1(_1879_),
    .A2(_2192_));
 sg13g2_a22oi_1 _5772_ (.Y(_2202_),
    .B1(_2184_),
    .B2(_2201_),
    .A2(_1824_),
    .A1(_0672_));
 sg13g2_nor2_2 _5773_ (.A(_2162_),
    .B(_2179_),
    .Y(_2203_));
 sg13g2_nor2_1 _5774_ (.A(_2162_),
    .B(_2180_),
    .Y(_2204_));
 sg13g2_nor2_2 _5775_ (.A(_2203_),
    .B(_2204_),
    .Y(_2205_));
 sg13g2_nand3_1 _5776_ (.B(net849),
    .C(_2165_),
    .A(_2161_),
    .Y(_2206_));
 sg13g2_nand3_1 _5777_ (.B(_2176_),
    .C(_2195_),
    .A(_2171_),
    .Y(_2207_));
 sg13g2_o21ai_1 _5778_ (.B1(_2205_),
    .Y(_2208_),
    .A1(_2206_),
    .A2(_2207_));
 sg13g2_nand2_1 _5779_ (.Y(_2209_),
    .A(_1862_),
    .B(_2208_));
 sg13g2_a21o_1 _5780_ (.A2(_2174_),
    .A1(_2169_),
    .B1(_2170_),
    .X(_2210_));
 sg13g2_nor2_1 _5781_ (.A(net880),
    .B(_2168_),
    .Y(_2211_));
 sg13g2_a21o_1 _5782_ (.A2(_2211_),
    .A1(_2210_),
    .B1(_2206_),
    .X(_2212_));
 sg13g2_a21oi_1 _5783_ (.A1(_2205_),
    .A2(_2212_),
    .Y(_2213_),
    .B1(_1825_));
 sg13g2_a21o_1 _5784_ (.A2(_2208_),
    .A1(_1862_),
    .B1(_2213_),
    .X(_2214_));
 sg13g2_nor2_1 _5785_ (.A(_2202_),
    .B(_2214_),
    .Y(_2215_));
 sg13g2_o21ai_1 _5786_ (.B1(_2209_),
    .Y(_2216_),
    .A1(_1862_),
    .A2(_2215_));
 sg13g2_o21ai_1 _5787_ (.B1(_2168_),
    .Y(_2217_),
    .A1(_2173_),
    .A2(_2186_));
 sg13g2_nor2_1 _5788_ (.A(_2165_),
    .B(net880),
    .Y(_2218_));
 sg13g2_nand2_1 _5789_ (.Y(_2219_),
    .A(_2217_),
    .B(_2218_));
 sg13g2_and3_1 _5790_ (.X(_2220_),
    .A(net849),
    .B(_2179_),
    .C(_2219_));
 sg13g2_a22oi_1 _5791_ (.Y(_2221_),
    .B1(_2204_),
    .B2(_2220_),
    .A2(_2203_),
    .A1(_2180_));
 sg13g2_nor2_1 _5792_ (.A(_1813_),
    .B(_2221_),
    .Y(_2222_));
 sg13g2_nor4_1 _5793_ (.A(_2164_),
    .B(net880),
    .C(_2167_),
    .D(_2210_),
    .Y(_2223_));
 sg13g2_nand2_1 _5794_ (.Y(_2224_),
    .A(_2180_),
    .B(_2193_));
 sg13g2_o21ai_1 _5795_ (.B1(_2203_),
    .Y(_2225_),
    .A1(_2223_),
    .A2(_2224_));
 sg13g2_a21oi_1 _5796_ (.A1(_2221_),
    .A2(_2225_),
    .Y(_2226_),
    .B1(_1813_));
 sg13g2_a21o_1 _5797_ (.A2(_2216_),
    .A1(_1813_),
    .B1(_2226_),
    .X(_2227_));
 sg13g2_o21ai_1 _5798_ (.B1(_2180_),
    .Y(_2228_),
    .A1(_2164_),
    .A2(_2177_));
 sg13g2_o21ai_1 _5799_ (.B1(_2203_),
    .Y(_2229_),
    .A1(net849),
    .A2(_2228_));
 sg13g2_nand2b_1 _5800_ (.Y(_2230_),
    .B(_2229_),
    .A_N(_1820_));
 sg13g2_nor2_1 _5801_ (.A(_2186_),
    .B(_2195_),
    .Y(_2231_));
 sg13g2_o21ai_1 _5802_ (.B1(_2189_),
    .Y(_2232_),
    .A1(_2185_),
    .A2(_2231_));
 sg13g2_and2_1 _5803_ (.A(_2163_),
    .B(_2232_),
    .X(_2233_));
 sg13g2_nand4_1 _5804_ (.B(_2180_),
    .C(_2203_),
    .A(_1818_),
    .Y(_2234_),
    .D(_2233_));
 sg13g2_a21o_1 _5805_ (.A2(_2187_),
    .A1(_2176_),
    .B1(_2165_),
    .X(_2235_));
 sg13g2_or3_1 _5806_ (.A(_1818_),
    .B(net849),
    .C(_2235_),
    .X(_2236_));
 sg13g2_nand3_1 _5807_ (.B(_2181_),
    .C(_2236_),
    .A(_2161_),
    .Y(_2237_));
 sg13g2_nand3_1 _5808_ (.B(_2234_),
    .C(_2237_),
    .A(_1843_),
    .Y(_2238_));
 sg13g2_nand4_1 _5809_ (.B(_2227_),
    .C(_2230_),
    .A(_2125_),
    .Y(_2239_),
    .D(_2238_));
 sg13g2_o21ai_1 _5810_ (.B1(_2239_),
    .Y(_2240_),
    .A1(_2123_),
    .A2(_2125_));
 sg13g2_a22oi_1 _5811_ (.Y(_2241_),
    .B1(_2240_),
    .B2(_1741_),
    .A2(_2124_),
    .A1(_1742_));
 sg13g2_a21oi_1 _5812_ (.A1(_1736_),
    .A2(net1708),
    .Y(_2242_),
    .B1(_2241_));
 sg13g2_nor2_1 _5813_ (.A(net967),
    .B(net1709),
    .Y(_0209_));
 sg13g2_nand2_2 _5814_ (.Y(_2243_),
    .A(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[1] ),
    .B(_0688_));
 sg13g2_nand4_1 _5815_ (.B(net6),
    .C(net955),
    .A(_0191_),
    .Y(_2244_),
    .D(_1955_));
 sg13g2_inv_1 _5816_ (.Y(_2245_),
    .A(_2244_));
 sg13g2_nor2_1 _5817_ (.A(_0686_),
    .B(net991),
    .Y(_2246_));
 sg13g2_nand2_1 _5818_ (.Y(_2247_),
    .A(_2245_),
    .B(_2246_));
 sg13g2_nor2_1 _5819_ (.A(_2243_),
    .B(_2247_),
    .Y(_2248_));
 sg13g2_nor2_1 _5820_ (.A(net1020),
    .B(net847),
    .Y(_2249_));
 sg13g2_a21oi_1 _5821_ (.A1(net874),
    .A2(net847),
    .Y(_0210_),
    .B1(_2249_));
 sg13g2_nor2_1 _5822_ (.A(net1172),
    .B(net848),
    .Y(_2250_));
 sg13g2_a21oi_1 _5823_ (.A1(net871),
    .A2(net847),
    .Y(_0211_),
    .B1(_2250_));
 sg13g2_nor2_1 _5824_ (.A(net1161),
    .B(net848),
    .Y(_2251_));
 sg13g2_a21oi_1 _5825_ (.A1(net866),
    .A2(net848),
    .Y(_0212_),
    .B1(_2251_));
 sg13g2_nor2_1 _5826_ (.A(net1251),
    .B(net848),
    .Y(_2252_));
 sg13g2_a21oi_1 _5827_ (.A1(net863),
    .A2(net848),
    .Y(_0213_),
    .B1(_2252_));
 sg13g2_nor2_1 _5828_ (.A(net1198),
    .B(net848),
    .Y(_2253_));
 sg13g2_a21oi_1 _5829_ (.A1(net856),
    .A2(_2248_),
    .Y(_0214_),
    .B1(_2253_));
 sg13g2_nor2_1 _5830_ (.A(net1089),
    .B(net848),
    .Y(_2254_));
 sg13g2_a21oi_1 _5831_ (.A1(net860),
    .A2(net847),
    .Y(_0215_),
    .B1(_2254_));
 sg13g2_nor2_1 _5832_ (.A(net1329),
    .B(net847),
    .Y(_2255_));
 sg13g2_a21oi_1 _5833_ (.A1(net853),
    .A2(net847),
    .Y(_0216_),
    .B1(_2255_));
 sg13g2_nor2_1 _5834_ (.A(net1077),
    .B(net847),
    .Y(_2256_));
 sg13g2_a21oi_1 _5835_ (.A1(net852),
    .A2(net847),
    .Y(_0217_),
    .B1(_2256_));
 sg13g2_a21o_2 _5836_ (.A2(net947),
    .A1(\FpgaPins_Fpga_UART_dptr_a2[1] ),
    .B1(net813),
    .X(_2257_));
 sg13g2_o21ai_1 _5837_ (.B1(net805),
    .Y(_2258_),
    .A1(_0207_),
    .A2(net976));
 sg13g2_nand2b_2 _5838_ (.Y(_2259_),
    .B(_2257_),
    .A_N(_2258_));
 sg13g2_o21ai_1 _5839_ (.B1(_1325_),
    .Y(_2260_),
    .A1(_0204_),
    .A2(net977));
 sg13g2_nor4_2 _5840_ (.A(_0752_),
    .B(net6),
    .C(net950),
    .Y(_2261_),
    .D(net902));
 sg13g2_a21oi_2 _5841_ (.B1(_2261_),
    .Y(_2262_),
    .A2(net783),
    .A1(net976));
 sg13g2_o21ai_1 _5842_ (.B1(net803),
    .Y(_2263_),
    .A1(_0203_),
    .A2(net977));
 sg13g2_nor2b_1 _5843_ (.A(_2262_),
    .B_N(_2263_),
    .Y(_2264_));
 sg13g2_nand2_2 _5844_ (.Y(_2265_),
    .A(_2260_),
    .B(_2264_));
 sg13g2_or2_2 _5845_ (.X(_2266_),
    .B(_2265_),
    .A(_2259_));
 sg13g2_nor2_1 _5846_ (.A(net947),
    .B(\FpgaPins_Fpga_LIPSI_data_wr_a1[0] ),
    .Y(_2267_));
 sg13g2_a21oi_2 _5847_ (.B1(_2267_),
    .Y(_2268_),
    .A2(net874),
    .A1(net947));
 sg13g2_mux2_1 _5848_ (.A0(net777),
    .A1(net1250),
    .S(_2266_),
    .X(_0218_));
 sg13g2_nor2_1 _5849_ (.A(net946),
    .B(\FpgaPins_Fpga_LIPSI_data_wr_a1[1] ),
    .Y(_2269_));
 sg13g2_a21oi_2 _5850_ (.B1(_2269_),
    .Y(_2270_),
    .A2(net871),
    .A1(net945));
 sg13g2_mux2_1 _5851_ (.A0(net775),
    .A1(net1284),
    .S(_2266_),
    .X(_0219_));
 sg13g2_nor2_1 _5852_ (.A(net945),
    .B(\FpgaPins_Fpga_LIPSI_data_wr_a1[2] ),
    .Y(_2271_));
 sg13g2_a21oi_2 _5853_ (.B1(_2271_),
    .Y(_2272_),
    .A2(net868),
    .A1(net945));
 sg13g2_mux2_1 _5854_ (.A0(net773),
    .A1(net1311),
    .S(_2266_),
    .X(_0220_));
 sg13g2_nor2_1 _5855_ (.A(net945),
    .B(\FpgaPins_Fpga_LIPSI_data_wr_a1[3] ),
    .Y(_2273_));
 sg13g2_a21oi_2 _5856_ (.B1(_2273_),
    .Y(_2274_),
    .A2(net865),
    .A1(net945));
 sg13g2_mux2_1 _5857_ (.A0(net762),
    .A1(net1306),
    .S(_2266_),
    .X(_0221_));
 sg13g2_nor2_1 _5858_ (.A(net947),
    .B(\FpgaPins_Fpga_LIPSI_data_wr_a1[4] ),
    .Y(_2275_));
 sg13g2_a21oi_2 _5859_ (.B1(_2275_),
    .Y(_2276_),
    .A2(net856),
    .A1(net947));
 sg13g2_mux2_1 _5860_ (.A0(net767),
    .A1(net1227),
    .S(_2266_),
    .X(_0222_));
 sg13g2_nor2_1 _5861_ (.A(net945),
    .B(\FpgaPins_Fpga_LIPSI_data_wr_a1[5] ),
    .Y(_2277_));
 sg13g2_a21oi_2 _5862_ (.B1(_2277_),
    .Y(_2278_),
    .A2(net862),
    .A1(net946));
 sg13g2_mux2_1 _5863_ (.A0(net765),
    .A1(net1438),
    .S(_2266_),
    .X(_0223_));
 sg13g2_nor2_1 _5864_ (.A(net946),
    .B(\FpgaPins_Fpga_LIPSI_data_wr_a1[6] ),
    .Y(_2279_));
 sg13g2_a21oi_2 _5865_ (.B1(_2279_),
    .Y(_2280_),
    .A2(net853),
    .A1(net945));
 sg13g2_mux2_1 _5866_ (.A0(net760),
    .A1(net1426),
    .S(_2266_),
    .X(_0224_));
 sg13g2_nor2_1 _5867_ (.A(net944),
    .B(\FpgaPins_Fpga_LIPSI_data_wr_a1[7] ),
    .Y(_2281_));
 sg13g2_a21oi_2 _5868_ (.B1(_2281_),
    .Y(_2282_),
    .A2(net852),
    .A1(net944));
 sg13g2_mux2_1 _5869_ (.A0(net758),
    .A1(net1490),
    .S(_2266_),
    .X(_0225_));
 sg13g2_or2_1 _5870_ (.X(_2283_),
    .B(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[0] ),
    .A(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[1] ));
 sg13g2_nor4_1 _5871_ (.A(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[3] ),
    .B(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[2] ),
    .C(_2244_),
    .D(_2283_),
    .Y(_2284_));
 sg13g2_nor2_1 _5872_ (.A(net1039),
    .B(net878),
    .Y(_2285_));
 sg13g2_a21oi_1 _5873_ (.A1(net873),
    .A2(net878),
    .Y(_0226_),
    .B1(_2285_));
 sg13g2_nor2_1 _5874_ (.A(net1113),
    .B(net878),
    .Y(_2286_));
 sg13g2_a21oi_1 _5875_ (.A1(net870),
    .A2(net878),
    .Y(_0227_),
    .B1(_2286_));
 sg13g2_nor2_1 _5876_ (.A(net1196),
    .B(net879),
    .Y(_2287_));
 sg13g2_a21oi_1 _5877_ (.A1(net867),
    .A2(net879),
    .Y(_0228_),
    .B1(_2287_));
 sg13g2_nor2_1 _5878_ (.A(net1152),
    .B(net879),
    .Y(_2288_));
 sg13g2_a21oi_1 _5879_ (.A1(net864),
    .A2(net879),
    .Y(_0229_),
    .B1(_2288_));
 sg13g2_nor2_1 _5880_ (.A(net1222),
    .B(net879),
    .Y(_2289_));
 sg13g2_a21oi_1 _5881_ (.A1(net858),
    .A2(net879),
    .Y(_0230_),
    .B1(_2289_));
 sg13g2_nor2_1 _5882_ (.A(net1122),
    .B(net878),
    .Y(_2290_));
 sg13g2_a21oi_1 _5883_ (.A1(net861),
    .A2(net878),
    .Y(_0231_),
    .B1(_2290_));
 sg13g2_nor2_1 _5884_ (.A(net1192),
    .B(net879),
    .Y(_2291_));
 sg13g2_a21oi_1 _5885_ (.A1(net855),
    .A2(net879),
    .Y(_0232_),
    .B1(_2291_));
 sg13g2_nor2_1 _5886_ (.A(net1044),
    .B(net878),
    .Y(_2292_));
 sg13g2_a21oi_1 _5887_ (.A1(net850),
    .A2(net878),
    .Y(_0233_),
    .B1(_2292_));
 sg13g2_nor2_1 _5888_ (.A(_2247_),
    .B(_2283_),
    .Y(_2293_));
 sg13g2_nor2_1 _5889_ (.A(net1100),
    .B(net845),
    .Y(_2294_));
 sg13g2_a21oi_1 _5890_ (.A1(net874),
    .A2(net845),
    .Y(_0234_),
    .B1(_2294_));
 sg13g2_nor2_1 _5891_ (.A(net1171),
    .B(net846),
    .Y(_2295_));
 sg13g2_a21oi_1 _5892_ (.A1(net871),
    .A2(net845),
    .Y(_0235_),
    .B1(_2295_));
 sg13g2_nor2_1 _5893_ (.A(net1213),
    .B(net846),
    .Y(_2296_));
 sg13g2_a21oi_1 _5894_ (.A1(net866),
    .A2(net846),
    .Y(_0236_),
    .B1(_2296_));
 sg13g2_nor2_1 _5895_ (.A(net1392),
    .B(net846),
    .Y(_2297_));
 sg13g2_a21oi_1 _5896_ (.A1(net863),
    .A2(net846),
    .Y(_0237_),
    .B1(_2297_));
 sg13g2_nor2_1 _5897_ (.A(net1182),
    .B(net846),
    .Y(_2298_));
 sg13g2_a21oi_1 _5898_ (.A1(net856),
    .A2(_2293_),
    .Y(_0238_),
    .B1(_2298_));
 sg13g2_nor2_1 _5899_ (.A(net1093),
    .B(net846),
    .Y(_2299_));
 sg13g2_a21oi_1 _5900_ (.A1(net860),
    .A2(net845),
    .Y(_0239_),
    .B1(_2299_));
 sg13g2_nor2_1 _5901_ (.A(net1146),
    .B(net845),
    .Y(_2300_));
 sg13g2_a21oi_1 _5902_ (.A1(net853),
    .A2(net845),
    .Y(_0240_),
    .B1(_2300_));
 sg13g2_nor2_1 _5903_ (.A(net1131),
    .B(net845),
    .Y(_2301_));
 sg13g2_a21oi_1 _5904_ (.A1(net852),
    .A2(net845),
    .Y(_0241_),
    .B1(_2301_));
 sg13g2_nor2_2 _5905_ (.A(_0688_),
    .B(_2244_),
    .Y(_2302_));
 sg13g2_and2_2 _5906_ (.A(net1649),
    .B(_2302_),
    .X(_2303_));
 sg13g2_nand2_1 _5907_ (.Y(_2304_),
    .A(net991),
    .B(_2303_));
 sg13g2_nand3_1 _5908_ (.B(net991),
    .C(_2303_),
    .A(_0686_),
    .Y(_2305_));
 sg13g2_nand2_1 _5909_ (.Y(_2306_),
    .A(net737),
    .B(net843));
 sg13g2_o21ai_1 _5910_ (.B1(_2306_),
    .Y(_0242_),
    .A1(net872),
    .A2(net843));
 sg13g2_nand2_1 _5911_ (.Y(_2307_),
    .A(net1079),
    .B(net843));
 sg13g2_o21ai_1 _5912_ (.B1(_2307_),
    .Y(_0243_),
    .A1(net869),
    .A2(net843));
 sg13g2_nand2_1 _5913_ (.Y(_2308_),
    .A(net1037),
    .B(_2305_));
 sg13g2_o21ai_1 _5914_ (.B1(_2308_),
    .Y(_0244_),
    .A1(net867),
    .A2(_2305_));
 sg13g2_nand2_1 _5915_ (.Y(_2309_),
    .A(net1015),
    .B(net844));
 sg13g2_o21ai_1 _5916_ (.B1(_2309_),
    .Y(_0245_),
    .A1(net864),
    .A2(net844));
 sg13g2_nand2_1 _5917_ (.Y(_2310_),
    .A(net1040),
    .B(net844));
 sg13g2_o21ai_1 _5918_ (.B1(_2310_),
    .Y(_0246_),
    .A1(net858),
    .A2(net844));
 sg13g2_nand2_1 _5919_ (.Y(_2311_),
    .A(net1010),
    .B(net843));
 sg13g2_o21ai_1 _5920_ (.B1(_2311_),
    .Y(_0247_),
    .A1(net861),
    .A2(net844));
 sg13g2_nand2_1 _5921_ (.Y(_2312_),
    .A(net1026),
    .B(net844));
 sg13g2_o21ai_1 _5922_ (.B1(_2312_),
    .Y(_0248_),
    .A1(net854),
    .A2(net844));
 sg13g2_nand2_1 _5923_ (.Y(_2313_),
    .A(net750),
    .B(net843));
 sg13g2_o21ai_1 _5924_ (.B1(_2313_),
    .Y(_0249_),
    .A1(net851),
    .A2(net843));
 sg13g2_nand2_2 _5925_ (.Y(_2314_),
    .A(_2257_),
    .B(_2258_));
 sg13g2_nor2_1 _5926_ (.A(_2262_),
    .B(_2263_),
    .Y(_2315_));
 sg13g2_nand2b_2 _5927_ (.Y(_2316_),
    .B(_2315_),
    .A_N(_2260_));
 sg13g2_or2_2 _5928_ (.X(_2317_),
    .B(_2316_),
    .A(_2314_));
 sg13g2_mux2_1 _5929_ (.A0(net776),
    .A1(net1295),
    .S(_2317_),
    .X(_0250_));
 sg13g2_mux2_1 _5930_ (.A0(net774),
    .A1(net1252),
    .S(_2317_),
    .X(_0251_));
 sg13g2_mux2_1 _5931_ (.A0(net772),
    .A1(net1225),
    .S(_2317_),
    .X(_0252_));
 sg13g2_mux2_1 _5932_ (.A0(net761),
    .A1(net1278),
    .S(_2317_),
    .X(_0253_));
 sg13g2_mux2_1 _5933_ (.A0(net766),
    .A1(net1234),
    .S(_2317_),
    .X(_0254_));
 sg13g2_mux2_1 _5934_ (.A0(net764),
    .A1(net1416),
    .S(_2317_),
    .X(_0255_));
 sg13g2_mux2_1 _5935_ (.A0(net759),
    .A1(net1486),
    .S(_2317_),
    .X(_0256_));
 sg13g2_mux2_1 _5936_ (.A0(net757),
    .A1(net1461),
    .S(_2317_),
    .X(_0257_));
 sg13g2_or2_2 _5937_ (.X(_2318_),
    .B(_2258_),
    .A(_2257_));
 sg13g2_nand2b_1 _5938_ (.Y(_2319_),
    .B(_2264_),
    .A_N(_2260_));
 sg13g2_nor2_1 _5939_ (.A(_2318_),
    .B(_2319_),
    .Y(_2320_));
 sg13g2_mux2_1 _5940_ (.A0(net1053),
    .A1(net777),
    .S(_2320_),
    .X(_0258_));
 sg13g2_mux2_1 _5941_ (.A0(net1065),
    .A1(net775),
    .S(net779),
    .X(_0259_));
 sg13g2_mux2_1 _5942_ (.A0(net1059),
    .A1(net772),
    .S(net779),
    .X(_0260_));
 sg13g2_mux2_1 _5943_ (.A0(net1087),
    .A1(net762),
    .S(net779),
    .X(_0261_));
 sg13g2_mux2_1 _5944_ (.A0(net1056),
    .A1(net767),
    .S(net779),
    .X(_0262_));
 sg13g2_nand2_1 _5945_ (.Y(_2321_),
    .A(net765),
    .B(net779));
 sg13g2_o21ai_1 _5946_ (.B1(_2321_),
    .Y(_0263_),
    .A1(_0744_),
    .A2(net779));
 sg13g2_mux2_1 _5947_ (.A0(net1208),
    .A1(net760),
    .S(net779),
    .X(_0264_));
 sg13g2_mux2_1 _5948_ (.A0(net1217),
    .A1(net758),
    .S(net779),
    .X(_0265_));
 sg13g2_nand2_1 _5949_ (.Y(_2322_),
    .A(_2246_),
    .B(_2303_));
 sg13g2_nand2_1 _5950_ (.Y(_2323_),
    .A(net1009),
    .B(net841));
 sg13g2_o21ai_1 _5951_ (.B1(_2323_),
    .Y(_0266_),
    .A1(net874),
    .A2(net841));
 sg13g2_nand2_1 _5952_ (.Y(_2324_),
    .A(net1027),
    .B(net841));
 sg13g2_o21ai_1 _5953_ (.B1(_2324_),
    .Y(_0267_),
    .A1(net871),
    .A2(net841));
 sg13g2_nand2_1 _5954_ (.Y(_2325_),
    .A(net1018),
    .B(net842));
 sg13g2_o21ai_1 _5955_ (.B1(_2325_),
    .Y(_0268_),
    .A1(net866),
    .A2(net842));
 sg13g2_nand2_1 _5956_ (.Y(_2326_),
    .A(net1019),
    .B(net842));
 sg13g2_o21ai_1 _5957_ (.B1(_2326_),
    .Y(_0269_),
    .A1(net863),
    .A2(net842));
 sg13g2_nand2_1 _5958_ (.Y(_2327_),
    .A(net1061),
    .B(net842));
 sg13g2_o21ai_1 _5959_ (.B1(_2327_),
    .Y(_0270_),
    .A1(net856),
    .A2(_2322_));
 sg13g2_nand2_1 _5960_ (.Y(_2328_),
    .A(net728),
    .B(net842));
 sg13g2_o21ai_1 _5961_ (.B1(_2328_),
    .Y(_0271_),
    .A1(net860),
    .A2(net841));
 sg13g2_nand2_1 _5962_ (.Y(_2329_),
    .A(net1206),
    .B(net841));
 sg13g2_o21ai_1 _5963_ (.B1(_2329_),
    .Y(_0272_),
    .A1(net853),
    .A2(net842));
 sg13g2_nand2_1 _5964_ (.Y(_2330_),
    .A(net1008),
    .B(net841));
 sg13g2_o21ai_1 _5965_ (.B1(_2330_),
    .Y(_0273_),
    .A1(net852),
    .A2(net841));
 sg13g2_or2_2 _5966_ (.X(_2331_),
    .B(_2316_),
    .A(_2259_));
 sg13g2_mux2_1 _5967_ (.A0(net776),
    .A1(net1253),
    .S(_2331_),
    .X(_0274_));
 sg13g2_mux2_1 _5968_ (.A0(net774),
    .A1(net1317),
    .S(_2331_),
    .X(_0275_));
 sg13g2_mux2_1 _5969_ (.A0(net772),
    .A1(net1231),
    .S(_2331_),
    .X(_0276_));
 sg13g2_mux2_1 _5970_ (.A0(net761),
    .A1(net1310),
    .S(_2331_),
    .X(_0277_));
 sg13g2_mux2_1 _5971_ (.A0(net766),
    .A1(net1299),
    .S(_2331_),
    .X(_0278_));
 sg13g2_mux2_1 _5972_ (.A0(net764),
    .A1(net1476),
    .S(_2331_),
    .X(_0279_));
 sg13g2_mux2_1 _5973_ (.A0(net759),
    .A1(net1474),
    .S(_2331_),
    .X(_0280_));
 sg13g2_mux2_1 _5974_ (.A0(net757),
    .A1(net1477),
    .S(_2331_),
    .X(_0281_));
 sg13g2_nand2b_2 _5975_ (.Y(_2332_),
    .B(_2258_),
    .A_N(_2257_));
 sg13g2_or2_2 _5976_ (.X(_2333_),
    .B(_2332_),
    .A(_2316_));
 sg13g2_mux2_1 _5977_ (.A0(net776),
    .A1(net1259),
    .S(_2333_),
    .X(_0282_));
 sg13g2_mux2_1 _5978_ (.A0(net774),
    .A1(net1258),
    .S(_2333_),
    .X(_0283_));
 sg13g2_mux2_1 _5979_ (.A0(net772),
    .A1(net1226),
    .S(_2333_),
    .X(_0284_));
 sg13g2_mux2_1 _5980_ (.A0(net761),
    .A1(net1215),
    .S(_2333_),
    .X(_0285_));
 sg13g2_mux2_1 _5981_ (.A0(net766),
    .A1(net1320),
    .S(_2333_),
    .X(_0286_));
 sg13g2_mux2_1 _5982_ (.A0(net764),
    .A1(net1475),
    .S(_2333_),
    .X(_0287_));
 sg13g2_mux2_1 _5983_ (.A0(net759),
    .A1(net1442),
    .S(_2333_),
    .X(_0288_));
 sg13g2_mux2_1 _5984_ (.A0(net757),
    .A1(net1470),
    .S(_2333_),
    .X(_0289_));
 sg13g2_nand2_1 _5985_ (.Y(_2334_),
    .A(net1512),
    .B(_1838_));
 sg13g2_a21oi_1 _5986_ (.A1(_1901_),
    .A2(_2334_),
    .Y(_0290_),
    .B1(net966));
 sg13g2_nand2_1 _5987_ (.Y(_2335_),
    .A(net1489),
    .B(_1838_));
 sg13g2_a21oi_1 _5988_ (.A1(_1893_),
    .A2(_2335_),
    .Y(_0291_),
    .B1(net966));
 sg13g2_o21ai_1 _5989_ (.B1(net974),
    .Y(_2336_),
    .A1(net1606),
    .A2(net936));
 sg13g2_a21oi_1 _5990_ (.A1(net936),
    .A2(_1882_),
    .Y(_0292_),
    .B1(_2336_));
 sg13g2_nor2_1 _5991_ (.A(_1804_),
    .B(_1880_),
    .Y(_2337_));
 sg13g2_xnor2_1 _5992_ (.Y(_2338_),
    .A(_1740_),
    .B(_1912_));
 sg13g2_xnor2_1 _5993_ (.Y(_2339_),
    .A(_2337_),
    .B(_2338_));
 sg13g2_o21ai_1 _5994_ (.B1(net974),
    .Y(_2340_),
    .A1(net1518),
    .A2(net937));
 sg13g2_a21oi_1 _5995_ (.A1(net937),
    .A2(_2339_),
    .Y(_0293_),
    .B1(_2340_));
 sg13g2_a21oi_1 _5996_ (.A1(_1805_),
    .A2(_1826_),
    .Y(_2341_),
    .B1(_1923_));
 sg13g2_o21ai_1 _5997_ (.B1(net937),
    .Y(_2342_),
    .A1(_1740_),
    .A2(_2341_));
 sg13g2_a21oi_1 _5998_ (.A1(_1740_),
    .A2(_1922_),
    .Y(_2343_),
    .B1(_2342_));
 sg13g2_o21ai_1 _5999_ (.B1(net974),
    .Y(_2344_),
    .A1(net1646),
    .A2(net937));
 sg13g2_nor2_1 _6000_ (.A(_2343_),
    .B(_2344_),
    .Y(_0294_));
 sg13g2_a22oi_1 _6001_ (.Y(_2345_),
    .B1(_1845_),
    .B2(_1855_),
    .A2(_1838_),
    .A1(net1440));
 sg13g2_nor2_1 _6002_ (.A(net967),
    .B(_2345_),
    .Y(_0295_));
 sg13g2_o21ai_1 _6003_ (.B1(_1815_),
    .Y(_2346_),
    .A1(_1804_),
    .A2(_1821_));
 sg13g2_nand2_1 _6004_ (.Y(_2347_),
    .A(_1827_),
    .B(net937));
 sg13g2_a21oi_1 _6005_ (.A1(net938),
    .A2(_2346_),
    .Y(_2348_),
    .B1(_2347_));
 sg13g2_a21oi_1 _6006_ (.A1(net1542),
    .A2(_1838_),
    .Y(_2349_),
    .B1(_2348_));
 sg13g2_nor2_1 _6007_ (.A(net967),
    .B(_2349_),
    .Y(_0296_));
 sg13g2_nor2_1 _6008_ (.A(_1838_),
    .B(_1863_),
    .Y(_2350_));
 sg13g2_o21ai_1 _6009_ (.B1(_2350_),
    .Y(_2351_),
    .A1(_1740_),
    .A2(_1860_));
 sg13g2_o21ai_1 _6010_ (.B1(_2351_),
    .Y(_2352_),
    .A1(net1631),
    .A2(net936));
 sg13g2_nor2_1 _6011_ (.A(net967),
    .B(_2352_),
    .Y(_0297_));
 sg13g2_nand2_1 _6012_ (.Y(_2353_),
    .A(net1473),
    .B(_1838_));
 sg13g2_a21oi_1 _6013_ (.A1(_1840_),
    .A2(_2353_),
    .Y(_0298_),
    .B1(net968));
 sg13g2_o21ai_1 _6014_ (.B1(net970),
    .Y(_2354_),
    .A1(net1635),
    .A2(net936));
 sg13g2_a21oi_1 _6015_ (.A1(_1790_),
    .A2(net936),
    .Y(_0299_),
    .B1(_2354_));
 sg13g2_xnor2_1 _6016_ (.Y(_2355_),
    .A(_1740_),
    .B(_1875_));
 sg13g2_o21ai_1 _6017_ (.B1(net970),
    .Y(_2356_),
    .A1(net1563),
    .A2(net937));
 sg13g2_a21oi_1 _6018_ (.A1(net937),
    .A2(_2355_),
    .Y(_0300_),
    .B1(_2356_));
 sg13g2_or2_2 _6019_ (.X(_2357_),
    .B(_2314_),
    .A(_2265_));
 sg13g2_mux2_1 _6020_ (.A0(net777),
    .A1(net1238),
    .S(_2357_),
    .X(_0301_));
 sg13g2_mux2_1 _6021_ (.A0(net775),
    .A1(net1263),
    .S(_2357_),
    .X(_0302_));
 sg13g2_mux2_1 _6022_ (.A0(net773),
    .A1(net1323),
    .S(_2357_),
    .X(_0303_));
 sg13g2_mux2_1 _6023_ (.A0(net762),
    .A1(net1293),
    .S(_2357_),
    .X(_0304_));
 sg13g2_mux2_1 _6024_ (.A0(net767),
    .A1(net1239),
    .S(_2357_),
    .X(_0305_));
 sg13g2_mux2_1 _6025_ (.A0(net765),
    .A1(net1337),
    .S(_2357_),
    .X(_0306_));
 sg13g2_mux2_1 _6026_ (.A0(net760),
    .A1(net1431),
    .S(_2357_),
    .X(_0307_));
 sg13g2_mux2_1 _6027_ (.A0(net758),
    .A1(net1372),
    .S(_2357_),
    .X(_0308_));
 sg13g2_nand3_1 _6028_ (.B(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[2] ),
    .C(_2245_),
    .A(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[3] ),
    .Y(_2358_));
 sg13g2_nor2_1 _6029_ (.A(_2283_),
    .B(_2358_),
    .Y(_2359_));
 sg13g2_nor2_1 _6030_ (.A(net1153),
    .B(_2359_),
    .Y(_2360_));
 sg13g2_a21oi_1 _6031_ (.A1(net872),
    .A2(net840),
    .Y(_0309_),
    .B1(net1154));
 sg13g2_nor2_1 _6032_ (.A(net1148),
    .B(net840),
    .Y(_2361_));
 sg13g2_a21oi_1 _6033_ (.A1(net869),
    .A2(net840),
    .Y(_0310_),
    .B1(_2361_));
 sg13g2_nor2_1 _6034_ (.A(net1126),
    .B(net839),
    .Y(_2362_));
 sg13g2_a21oi_1 _6035_ (.A1(net866),
    .A2(net839),
    .Y(_0311_),
    .B1(_2362_));
 sg13g2_nor2_1 _6036_ (.A(net1149),
    .B(net840),
    .Y(_2363_));
 sg13g2_a21oi_1 _6037_ (.A1(net863),
    .A2(net840),
    .Y(_0312_),
    .B1(_2363_));
 sg13g2_nor2_1 _6038_ (.A(net1151),
    .B(net839),
    .Y(_2364_));
 sg13g2_a21oi_1 _6039_ (.A1(net857),
    .A2(net840),
    .Y(_0313_),
    .B1(_2364_));
 sg13g2_nor2_1 _6040_ (.A(net1096),
    .B(net840),
    .Y(_2365_));
 sg13g2_a21oi_1 _6041_ (.A1(net860),
    .A2(net839),
    .Y(_0314_),
    .B1(_2365_));
 sg13g2_nor2_1 _6042_ (.A(net1155),
    .B(net839),
    .Y(_2366_));
 sg13g2_a21oi_1 _6043_ (.A1(net854),
    .A2(net839),
    .Y(_0315_),
    .B1(_2366_));
 sg13g2_nor2_1 _6044_ (.A(net1111),
    .B(net839),
    .Y(_2367_));
 sg13g2_a21oi_1 _6045_ (.A1(net850),
    .A2(net839),
    .Y(_0316_),
    .B1(_2367_));
 sg13g2_nand2b_2 _6046_ (.Y(_2368_),
    .B(_2302_),
    .A_N(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[1] ));
 sg13g2_nor3_2 _6047_ (.A(_0686_),
    .B(_0687_),
    .C(_2368_),
    .Y(_2369_));
 sg13g2_nor2_1 _6048_ (.A(net1118),
    .B(net837),
    .Y(_2370_));
 sg13g2_a21oi_1 _6049_ (.A1(net872),
    .A2(net837),
    .Y(_0317_),
    .B1(_2370_));
 sg13g2_nor2_1 _6050_ (.A(net1341),
    .B(net837),
    .Y(_2371_));
 sg13g2_a21oi_1 _6051_ (.A1(net869),
    .A2(net837),
    .Y(_0318_),
    .B1(_2371_));
 sg13g2_nor2_1 _6052_ (.A(net1221),
    .B(net838),
    .Y(_2372_));
 sg13g2_a21oi_1 _6053_ (.A1(net866),
    .A2(_2369_),
    .Y(_0319_),
    .B1(_2372_));
 sg13g2_nor2_1 _6054_ (.A(net1150),
    .B(net837),
    .Y(_2373_));
 sg13g2_a21oi_1 _6055_ (.A1(net863),
    .A2(net837),
    .Y(_0320_),
    .B1(_2373_));
 sg13g2_nor2_1 _6056_ (.A(net1230),
    .B(net837),
    .Y(_2374_));
 sg13g2_a21oi_1 _6057_ (.A1(net857),
    .A2(net837),
    .Y(_0321_),
    .B1(_2374_));
 sg13g2_nor2_1 _6058_ (.A(net1025),
    .B(net838),
    .Y(_2375_));
 sg13g2_a21oi_1 _6059_ (.A1(net860),
    .A2(net838),
    .Y(_0322_),
    .B1(_2375_));
 sg13g2_nor2_1 _6060_ (.A(net1248),
    .B(net838),
    .Y(_2376_));
 sg13g2_a21oi_1 _6061_ (.A1(net854),
    .A2(net838),
    .Y(_0323_),
    .B1(_2376_));
 sg13g2_nor2_1 _6062_ (.A(net1069),
    .B(net838),
    .Y(_2377_));
 sg13g2_a21oi_1 _6063_ (.A1(net850),
    .A2(net838),
    .Y(_0324_),
    .B1(_2377_));
 sg13g2_o21ai_1 _6064_ (.B1(net961),
    .Y(_2378_),
    .A1(net1042),
    .A2(_2244_));
 sg13g2_a21oi_1 _6065_ (.A1(_0688_),
    .A2(_2244_),
    .Y(_0325_),
    .B1(_2378_));
 sg13g2_o21ai_1 _6066_ (.B1(net961),
    .Y(_2379_),
    .A1(net1649),
    .A2(_2302_));
 sg13g2_nor2_1 _6067_ (.A(_2303_),
    .B(net1650),
    .Y(_0326_));
 sg13g2_o21ai_1 _6068_ (.B1(net961),
    .Y(_2380_),
    .A1(net991),
    .A2(_2303_));
 sg13g2_nor2b_1 _6069_ (.A(_2380_),
    .B_N(_2304_),
    .Y(_0327_));
 sg13g2_nor2_1 _6070_ (.A(_0686_),
    .B(_2304_),
    .Y(_2381_));
 sg13g2_nand2_1 _6071_ (.Y(_2382_),
    .A(net1690),
    .B(_2304_));
 sg13g2_a21oi_1 _6072_ (.A1(net843),
    .A2(_2382_),
    .Y(_0328_),
    .B1(net952));
 sg13g2_nor2_1 _6073_ (.A(_1777_),
    .B(_1930_),
    .Y(_2383_));
 sg13g2_nand2_1 _6074_ (.Y(_2384_),
    .A(net970),
    .B(net771));
 sg13g2_nand2b_1 _6075_ (.Y(_2385_),
    .B(net1271),
    .A_N(_1770_));
 sg13g2_a21oi_1 _6076_ (.A1(_1771_),
    .A2(net1272),
    .Y(_0329_),
    .B1(net763));
 sg13g2_xor2_1 _6077_ (.B(_1771_),
    .A(net1617),
    .X(_2386_));
 sg13g2_nor2_1 _6078_ (.A(net763),
    .B(net1618),
    .Y(_0330_));
 sg13g2_o21ai_1 _6079_ (.B1(net1651),
    .Y(_2387_),
    .A1(net1617),
    .A2(_1771_));
 sg13g2_nor2b_1 _6080_ (.A(net1652),
    .B_N(_2387_),
    .Y(_2388_));
 sg13g2_nor2_1 _6081_ (.A(net763),
    .B(_2388_),
    .Y(_0331_));
 sg13g2_nand2b_1 _6082_ (.Y(_2389_),
    .B(net1186),
    .A_N(_1772_));
 sg13g2_a21oi_1 _6083_ (.A1(_1773_),
    .A2(net1187),
    .Y(_0332_),
    .B1(net763));
 sg13g2_xor2_1 _6084_ (.B(_1773_),
    .A(net1632),
    .X(_2390_));
 sg13g2_nor2_1 _6085_ (.A(net763),
    .B(net1633),
    .Y(_0333_));
 sg13g2_o21ai_1 _6086_ (.B1(net1658),
    .Y(_2391_),
    .A1(net1632),
    .A2(_1773_));
 sg13g2_nor2b_1 _6087_ (.A(_1774_),
    .B_N(_2391_),
    .Y(_2392_));
 sg13g2_nor2_1 _6088_ (.A(net763),
    .B(_2392_),
    .Y(_0334_));
 sg13g2_nand2b_1 _6089_ (.Y(_2393_),
    .B(net1286),
    .A_N(_1774_));
 sg13g2_a21oi_1 _6090_ (.A1(_1775_),
    .A2(net1287),
    .Y(_0335_),
    .B1(net763));
 sg13g2_xor2_1 _6091_ (.B(_1775_),
    .A(net1613),
    .X(_2394_));
 sg13g2_nor2_1 _6092_ (.A(net763),
    .B(net1614),
    .Y(_0336_));
 sg13g2_o21ai_1 _6093_ (.B1(net1656),
    .Y(_2395_),
    .A1(net1613),
    .A2(_1775_));
 sg13g2_nor2b_1 _6094_ (.A(net1657),
    .B_N(_2395_),
    .Y(_2396_));
 sg13g2_nor2_1 _6095_ (.A(_2384_),
    .B(_2396_),
    .Y(_0337_));
 sg13g2_nor3_1 _6096_ (.A(_0717_),
    .B(_1776_),
    .C(_2384_),
    .Y(_0338_));
 sg13g2_o21ai_1 _6097_ (.B1(net962),
    .Y(_2397_),
    .A1(\FpgaPins_Fpga_UART_dptr_a2[0] ),
    .A2(_2261_));
 sg13g2_a21oi_1 _6098_ (.A1(_0685_),
    .A2(_2261_),
    .Y(_0339_),
    .B1(_2397_));
 sg13g2_and2_1 _6099_ (.A(\FpgaPins_Fpga_UART_dptr_a2[0] ),
    .B(_2261_),
    .X(_2398_));
 sg13g2_and2_1 _6100_ (.A(net1587),
    .B(_2398_),
    .X(_2399_));
 sg13g2_o21ai_1 _6101_ (.B1(net962),
    .Y(_2400_),
    .A1(net1587),
    .A2(_2398_));
 sg13g2_nor2_1 _6102_ (.A(_2399_),
    .B(net1588),
    .Y(_0340_));
 sg13g2_o21ai_1 _6103_ (.B1(net962),
    .Y(_2401_),
    .A1(net745),
    .A2(_2399_));
 sg13g2_a21oi_1 _6104_ (.A1(net745),
    .A2(_2399_),
    .Y(_0341_),
    .B1(_2401_));
 sg13g2_nor2b_1 _6105_ (.A(_0203_),
    .B_N(_2399_),
    .Y(_2402_));
 sg13g2_o21ai_1 _6106_ (.B1(net962),
    .Y(_2403_),
    .A1(net729),
    .A2(_2402_));
 sg13g2_a21oi_1 _6107_ (.A1(net729),
    .A2(_2402_),
    .Y(_0342_),
    .B1(_2403_));
 sg13g2_a21oi_1 _6108_ (.A1(\FpgaPins_Fpga_LIPSI_acc_a2[7] ),
    .A2(_1701_),
    .Y(_2404_),
    .B1(_1725_));
 sg13g2_o21ai_1 _6109_ (.B1(net787),
    .Y(_2405_),
    .A1(_1727_),
    .A2(_2404_));
 sg13g2_a21oi_1 _6110_ (.A1(_1727_),
    .A2(_2404_),
    .Y(_2406_),
    .B1(_2405_));
 sg13g2_nor2_1 _6111_ (.A(\FpgaPins_Fpga_LIPSI_acc_a2[0] ),
    .B(_0867_),
    .Y(_2407_));
 sg13g2_or4_1 _6112_ (.A(_1297_),
    .B(_1348_),
    .C(net786),
    .D(_2407_),
    .X(_2408_));
 sg13g2_a21oi_2 _6113_ (.B1(_2408_),
    .Y(_2409_),
    .A2(net791),
    .A1(_0123_));
 sg13g2_o21ai_1 _6114_ (.B1(_1377_),
    .Y(_2410_),
    .A1(_2406_),
    .A2(_2409_));
 sg13g2_nand2b_1 _6115_ (.Y(_2411_),
    .B(_1705_),
    .A_N(_1702_));
 sg13g2_o21ai_1 _6116_ (.B1(net785),
    .Y(_2412_),
    .A1(_1707_),
    .A2(_2411_));
 sg13g2_a21oi_1 _6117_ (.A1(_1707_),
    .A2(_2411_),
    .Y(_2413_),
    .B1(_2412_));
 sg13g2_nor2_1 _6118_ (.A(net780),
    .B(_2413_),
    .Y(_2414_));
 sg13g2_o21ai_1 _6119_ (.B1(_1386_),
    .Y(_2415_),
    .A1(_1383_),
    .A2(_2404_));
 sg13g2_a21o_1 _6120_ (.A2(_2414_),
    .A1(_2410_),
    .B1(_2415_),
    .X(_2416_));
 sg13g2_a21oi_1 _6121_ (.A1(_1294_),
    .A2(_1348_),
    .Y(_2417_),
    .B1(_1297_));
 sg13g2_a221oi_1 _6122_ (.B2(_2411_),
    .C1(_1297_),
    .B1(net784),
    .A1(_1294_),
    .Y(_2418_),
    .A2(_1348_));
 sg13g2_o21ai_1 _6123_ (.B1(net976),
    .Y(_2419_),
    .A1(net1653),
    .A2(_2417_));
 sg13g2_a21oi_1 _6124_ (.A1(_2416_),
    .A2(_2418_),
    .Y(_0343_),
    .B1(_2419_));
 sg13g2_xor2_1 _6125_ (.B(net902),
    .A(net1664),
    .X(_2420_));
 sg13g2_nand2_1 _6126_ (.Y(_0344_),
    .A(net955),
    .B(_2420_));
 sg13g2_nand3_1 _6127_ (.B(_1214_),
    .C(_1215_),
    .A(_0693_),
    .Y(_2421_));
 sg13g2_nor4_1 _6128_ (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[10] ),
    .B(\FpgaPins_Fpga_GAME_wait_counter_a2[11] ),
    .C(\FpgaPins_Fpga_GAME_wait_counter_a2[13] ),
    .D(\FpgaPins_Fpga_GAME_wait_counter_a2[12] ),
    .Y(_2422_));
 sg13g2_nor2_1 _6129_ (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[6] ),
    .B(\FpgaPins_Fpga_GAME_wait_counter_a2[21] ),
    .Y(_2423_));
 sg13g2_nand3_1 _6130_ (.B(\FpgaPins_Fpga_GAME_wait_counter_a2[8] ),
    .C(net1524),
    .A(net1504),
    .Y(_2424_));
 sg13g2_nand3_1 _6131_ (.B(\FpgaPins_Fpga_GAME_wait_counter_a2[23] ),
    .C(\FpgaPins_Fpga_GAME_wait_counter_a2[24] ),
    .A(\FpgaPins_Fpga_GAME_wait_counter_a2[22] ),
    .Y(_2425_));
 sg13g2_nor2_1 _6132_ (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[17] ),
    .B(\FpgaPins_Fpga_GAME_wait_counter_a2[18] ),
    .Y(_2426_));
 sg13g2_nand2b_1 _6133_ (.Y(_2427_),
    .B(\FpgaPins_Fpga_GAME_state_a2[1] ),
    .A_N(\FpgaPins_Fpga_GAME_state_a2[0] ));
 sg13g2_nor3_1 _6134_ (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[3] ),
    .B(\FpgaPins_Fpga_GAME_wait_counter_a2[2] ),
    .C(\FpgaPins_Fpga_GAME_wait_counter_a2[5] ),
    .Y(_2428_));
 sg13g2_nand2b_1 _6135_ (.Y(_2429_),
    .B(\FpgaPins_Fpga_GAME_wait_counter_a2[20] ),
    .A_N(\FpgaPins_Fpga_GAME_wait_counter_a2[21] ));
 sg13g2_nand4_1 _6136_ (.B(\FpgaPins_Fpga_GAME_wait_counter_a2[19] ),
    .C(_2423_),
    .A(net1243),
    .Y(_2430_),
    .D(_2428_));
 sg13g2_nand4_1 _6137_ (.B(\FpgaPins_Fpga_GAME_wait_counter_a2[8] ),
    .C(\FpgaPins_Fpga_GAME_wait_counter_a2[9] ),
    .A(\FpgaPins_Fpga_GAME_wait_counter_a2[7] ),
    .Y(_2431_),
    .D(_2422_));
 sg13g2_nand4_1 _6138_ (.B(\FpgaPins_Fpga_GAME_wait_counter_a2[23] ),
    .C(\FpgaPins_Fpga_GAME_wait_counter_a2[24] ),
    .A(\FpgaPins_Fpga_GAME_wait_counter_a2[22] ),
    .Y(_2432_),
    .D(_2429_));
 sg13g2_or2_1 _6139_ (.X(_2433_),
    .B(_2432_),
    .A(_2431_));
 sg13g2_nor3_1 _6140_ (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[0] ),
    .B(\FpgaPins_Fpga_GAME_wait_counter_a2[1] ),
    .C(_2427_),
    .Y(_2434_));
 sg13g2_nand4_1 _6141_ (.B(net1678),
    .C(_2426_),
    .A(net1495),
    .Y(_2435_),
    .D(_2434_));
 sg13g2_nor4_2 _6142_ (.A(net1501),
    .B(_2430_),
    .C(_2433_),
    .Y(_2436_),
    .D(_2435_));
 sg13g2_nand4_1 _6143_ (.B(net706),
    .C(_1196_),
    .A(_0684_),
    .Y(_2437_),
    .D(_1197_));
 sg13g2_o21ai_1 _6144_ (.B1(_2437_),
    .Y(_2438_),
    .A1(net706),
    .A2(net1679));
 sg13g2_nand2b_1 _6145_ (.Y(_0345_),
    .B(net1680),
    .A_N(_2421_));
 sg13g2_o21ai_1 _6146_ (.B1(_2437_),
    .Y(_2439_),
    .A1(_0684_),
    .A2(_2436_));
 sg13g2_nor2b_1 _6147_ (.A(_2421_),
    .B_N(_2439_),
    .Y(_0346_));
 sg13g2_nor2_1 _6148_ (.A(net712),
    .B(_1201_),
    .Y(_2440_));
 sg13g2_nor2_1 _6149_ (.A(net720),
    .B(_1202_),
    .Y(_2441_));
 sg13g2_nor4_1 _6150_ (.A(net1492),
    .B(_1211_),
    .C(_2440_),
    .D(_2441_),
    .Y(_0347_));
 sg13g2_nor2_1 _6151_ (.A(_1202_),
    .B(_1211_),
    .Y(_2442_));
 sg13g2_nand2_2 _6152_ (.Y(_2443_),
    .A(_1201_),
    .B(_1212_));
 sg13g2_o21ai_1 _6153_ (.B1(_0693_),
    .Y(_2444_),
    .A1(net720),
    .A2(_1212_));
 sg13g2_a221oi_1 _6154_ (.B2(_0683_),
    .C1(_2444_),
    .B1(_2442_),
    .A1(_0682_),
    .Y(_0348_),
    .A2(_1202_));
 sg13g2_a22oi_1 _6155_ (.Y(_2445_),
    .B1(_1212_),
    .B2(_0681_),
    .A2(_1201_),
    .A1(_0683_));
 sg13g2_mux2_1 _6156_ (.A0(net713),
    .A1(_2445_),
    .S(_2443_),
    .X(_2446_));
 sg13g2_and2_1 _6157_ (.A(_0693_),
    .B(_2446_),
    .X(_0349_));
 sg13g2_nor2b_1 _6158_ (.A(net720),
    .B_N(_1204_),
    .Y(_2447_));
 sg13g2_nor3_1 _6159_ (.A(net716),
    .B(_1201_),
    .C(_2447_),
    .Y(_2448_));
 sg13g2_o21ai_1 _6160_ (.B1(_0693_),
    .Y(_2449_),
    .A1(net713),
    .A2(_1212_));
 sg13g2_nor2_1 _6161_ (.A(net715),
    .B(_2443_),
    .Y(_2450_));
 sg13g2_nor3_1 _6162_ (.A(_2448_),
    .B(_2449_),
    .C(_2450_),
    .Y(_0350_));
 sg13g2_a22oi_1 _6163_ (.Y(_2451_),
    .B1(_2442_),
    .B2(net716),
    .A2(_1202_),
    .A1(net710));
 sg13g2_o21ai_1 _6164_ (.B1(_1211_),
    .Y(_2452_),
    .A1(net715),
    .A2(_2447_));
 sg13g2_a21oi_1 _6165_ (.A1(_2451_),
    .A2(_2452_),
    .Y(_0351_),
    .B1(net1492));
 sg13g2_nor2_1 _6166_ (.A(net710),
    .B(_2443_),
    .Y(_2453_));
 sg13g2_nor2_1 _6167_ (.A(net721),
    .B(_1201_),
    .Y(_2454_));
 sg13g2_o21ai_1 _6168_ (.B1(_0693_),
    .Y(_2455_),
    .A1(net716),
    .A2(_1212_));
 sg13g2_nor3_1 _6169_ (.A(_2453_),
    .B(_2454_),
    .C(_2455_),
    .Y(_0352_));
 sg13g2_nor2_1 _6170_ (.A(net721),
    .B(_2443_),
    .Y(_2456_));
 sg13g2_o21ai_1 _6171_ (.B1(_0693_),
    .Y(_2457_),
    .A1(net714),
    .A2(_1201_));
 sg13g2_nor2_1 _6172_ (.A(net710),
    .B(_1212_),
    .Y(_2458_));
 sg13g2_nor3_1 _6173_ (.A(_2456_),
    .B(_2457_),
    .C(_2458_),
    .Y(_0353_));
 sg13g2_a22oi_1 _6174_ (.Y(_2459_),
    .B1(_2442_),
    .B2(net714),
    .A2(_1211_),
    .A1(net721));
 sg13g2_nor2_1 _6175_ (.A(net1492),
    .B(_2459_),
    .Y(_0354_));
 sg13g2_a21oi_1 _6176_ (.A1(\FpgaPins_Fpga_GAME_led_output_a1[3] ),
    .A2(_1238_),
    .Y(_2460_),
    .B1(_1233_));
 sg13g2_o21ai_1 _6177_ (.B1(_2460_),
    .Y(_2461_),
    .A1(net984),
    .A2(_1230_));
 sg13g2_a21oi_1 _6178_ (.A1(net984),
    .A2(_1239_),
    .Y(_2462_),
    .B1(_0791_));
 sg13g2_nand2_1 _6179_ (.Y(_0355_),
    .A(net1729),
    .B(_2462_));
 sg13g2_or2_1 _6180_ (.X(_2463_),
    .B(_2332_),
    .A(_2265_));
 sg13g2_mux2_1 _6181_ (.A0(net777),
    .A1(net1312),
    .S(net778),
    .X(_0356_));
 sg13g2_mux2_1 _6182_ (.A0(net775),
    .A1(net1316),
    .S(net778),
    .X(_0357_));
 sg13g2_mux2_1 _6183_ (.A0(net773),
    .A1(net1297),
    .S(net778),
    .X(_0358_));
 sg13g2_mux2_1 _6184_ (.A0(net762),
    .A1(net1246),
    .S(net778),
    .X(_0359_));
 sg13g2_mux2_1 _6185_ (.A0(net767),
    .A1(net1247),
    .S(_2463_),
    .X(_0360_));
 sg13g2_nor2_1 _6186_ (.A(net765),
    .B(net778),
    .Y(_2464_));
 sg13g2_a21oi_1 _6187_ (.A1(_0745_),
    .A2(net778),
    .Y(_0361_),
    .B1(_2464_));
 sg13g2_mux2_1 _6188_ (.A0(net760),
    .A1(net1447),
    .S(net778),
    .X(_0362_));
 sg13g2_mux2_1 _6189_ (.A0(net758),
    .A1(net1491),
    .S(net778),
    .X(_0363_));
 sg13g2_nand3_1 _6190_ (.B(net991),
    .C(_2245_),
    .A(_0686_),
    .Y(_2465_));
 sg13g2_nor2_1 _6191_ (.A(_2243_),
    .B(_2465_),
    .Y(_2466_));
 sg13g2_nor2_1 _6192_ (.A(net1049),
    .B(net835),
    .Y(_2467_));
 sg13g2_a21oi_1 _6193_ (.A1(net872),
    .A2(net835),
    .Y(_0364_),
    .B1(_2467_));
 sg13g2_nor2_1 _6194_ (.A(net1344),
    .B(net835),
    .Y(_2468_));
 sg13g2_a21oi_1 _6195_ (.A1(net869),
    .A2(net835),
    .Y(_0365_),
    .B1(_2468_));
 sg13g2_nor2_1 _6196_ (.A(net1256),
    .B(net836),
    .Y(_2469_));
 sg13g2_a21oi_1 _6197_ (.A1(net867),
    .A2(net836),
    .Y(_0366_),
    .B1(_2469_));
 sg13g2_nor2_1 _6198_ (.A(net1141),
    .B(net836),
    .Y(_2470_));
 sg13g2_a21oi_1 _6199_ (.A1(net864),
    .A2(net836),
    .Y(_0367_),
    .B1(_2470_));
 sg13g2_nor2_1 _6200_ (.A(net1331),
    .B(net836),
    .Y(_2471_));
 sg13g2_a21oi_1 _6201_ (.A1(net857),
    .A2(_2466_),
    .Y(_0368_),
    .B1(_2471_));
 sg13g2_nor2_1 _6202_ (.A(net1051),
    .B(net836),
    .Y(_2472_));
 sg13g2_a21oi_1 _6203_ (.A1(net861),
    .A2(net836),
    .Y(_0369_),
    .B1(_2472_));
 sg13g2_nor2_1 _6204_ (.A(net1132),
    .B(net835),
    .Y(_2473_));
 sg13g2_a21oi_1 _6205_ (.A1(net854),
    .A2(net835),
    .Y(_0370_),
    .B1(_2473_));
 sg13g2_nor2_1 _6206_ (.A(net1071),
    .B(net835),
    .Y(_2474_));
 sg13g2_a21oi_1 _6207_ (.A1(net851),
    .A2(net835),
    .Y(_0371_),
    .B1(_2474_));
 sg13g2_nor2_2 _6208_ (.A(_2265_),
    .B(_2318_),
    .Y(_2475_));
 sg13g2_mux2_1 _6209_ (.A0(net1074),
    .A1(net777),
    .S(_2475_),
    .X(_0372_));
 sg13g2_mux2_1 _6210_ (.A0(net1072),
    .A1(net775),
    .S(_2475_),
    .X(_0373_));
 sg13g2_mux2_1 _6211_ (.A0(net1088),
    .A1(net773),
    .S(_2475_),
    .X(_0374_));
 sg13g2_mux2_1 _6212_ (.A0(net1050),
    .A1(net762),
    .S(_2475_),
    .X(_0375_));
 sg13g2_mux2_1 _6213_ (.A0(net1045),
    .A1(net767),
    .S(_2475_),
    .X(_0376_));
 sg13g2_mux2_1 _6214_ (.A0(net1220),
    .A1(net765),
    .S(_2475_),
    .X(_0377_));
 sg13g2_mux2_1 _6215_ (.A0(net1322),
    .A1(net760),
    .S(_2475_),
    .X(_0378_));
 sg13g2_mux2_1 _6216_ (.A0(net1237),
    .A1(net758),
    .S(_2475_),
    .X(_0379_));
 sg13g2_nor3_2 _6217_ (.A(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[3] ),
    .B(_0687_),
    .C(_2368_),
    .Y(_2476_));
 sg13g2_nor2_1 _6218_ (.A(net1147),
    .B(net833),
    .Y(_2477_));
 sg13g2_a21oi_1 _6219_ (.A1(net872),
    .A2(net833),
    .Y(_0380_),
    .B1(_2477_));
 sg13g2_nor2_1 _6220_ (.A(net1158),
    .B(net833),
    .Y(_2478_));
 sg13g2_a21oi_1 _6221_ (.A1(net869),
    .A2(net833),
    .Y(_0381_),
    .B1(_2478_));
 sg13g2_nor2_1 _6222_ (.A(net1229),
    .B(net833),
    .Y(_2479_));
 sg13g2_a21oi_1 _6223_ (.A1(net867),
    .A2(net833),
    .Y(_0382_),
    .B1(_2479_));
 sg13g2_nor2_1 _6224_ (.A(net1294),
    .B(net834),
    .Y(_2480_));
 sg13g2_a21oi_1 _6225_ (.A1(net864),
    .A2(net834),
    .Y(_0383_),
    .B1(_2480_));
 sg13g2_nor2_1 _6226_ (.A(net1335),
    .B(net834),
    .Y(_2481_));
 sg13g2_a21oi_1 _6227_ (.A1(net857),
    .A2(net834),
    .Y(_0384_),
    .B1(_2481_));
 sg13g2_nor2_1 _6228_ (.A(net1106),
    .B(net834),
    .Y(_2482_));
 sg13g2_a21oi_1 _6229_ (.A1(net861),
    .A2(net834),
    .Y(_0385_),
    .B1(_2482_));
 sg13g2_nor2_1 _6230_ (.A(net1112),
    .B(net833),
    .Y(_2483_));
 sg13g2_a21oi_1 _6231_ (.A1(net854),
    .A2(net833),
    .Y(_0386_),
    .B1(_2483_));
 sg13g2_nor2_1 _6232_ (.A(net1036),
    .B(net834),
    .Y(_2484_));
 sg13g2_a21oi_1 _6233_ (.A1(net851),
    .A2(net834),
    .Y(_0387_),
    .B1(_2484_));
 sg13g2_nand2_1 _6234_ (.Y(_2485_),
    .A(_2260_),
    .B(_2315_));
 sg13g2_or2_2 _6235_ (.X(_2486_),
    .B(_2485_),
    .A(_2314_));
 sg13g2_mux2_1 _6236_ (.A0(net776),
    .A1(net1232),
    .S(_2486_),
    .X(_0388_));
 sg13g2_mux2_1 _6237_ (.A0(net774),
    .A1(net1241),
    .S(_2486_),
    .X(_0389_));
 sg13g2_mux2_1 _6238_ (.A0(net773),
    .A1(net1290),
    .S(_2486_),
    .X(_0390_));
 sg13g2_mux2_1 _6239_ (.A0(net761),
    .A1(net1261),
    .S(_2486_),
    .X(_0391_));
 sg13g2_mux2_1 _6240_ (.A0(net766),
    .A1(net1279),
    .S(_2486_),
    .X(_0392_));
 sg13g2_mux2_1 _6241_ (.A0(net764),
    .A1(net1425),
    .S(_2486_),
    .X(_0393_));
 sg13g2_mux2_1 _6242_ (.A0(net759),
    .A1(net1355),
    .S(_2486_),
    .X(_0394_));
 sg13g2_mux2_1 _6243_ (.A0(net757),
    .A1(net1439),
    .S(_2486_),
    .X(_0395_));
 sg13g2_nor2_1 _6244_ (.A(_2283_),
    .B(_2465_),
    .Y(_2487_));
 sg13g2_nor2_1 _6245_ (.A(net1035),
    .B(net831),
    .Y(_2488_));
 sg13g2_a21oi_1 _6246_ (.A1(net872),
    .A2(net831),
    .Y(_0396_),
    .B1(_2488_));
 sg13g2_nor2_1 _6247_ (.A(net1254),
    .B(net831),
    .Y(_2489_));
 sg13g2_a21oi_1 _6248_ (.A1(net869),
    .A2(net831),
    .Y(_0397_),
    .B1(_2489_));
 sg13g2_nor2_1 _6249_ (.A(net1328),
    .B(net832),
    .Y(_2490_));
 sg13g2_a21oi_1 _6250_ (.A1(net867),
    .A2(net831),
    .Y(_0398_),
    .B1(_2490_));
 sg13g2_nor2_1 _6251_ (.A(net1264),
    .B(net832),
    .Y(_2491_));
 sg13g2_a21oi_1 _6252_ (.A1(net864),
    .A2(net832),
    .Y(_0399_),
    .B1(_2491_));
 sg13g2_nor2_1 _6253_ (.A(net1360),
    .B(net832),
    .Y(_2492_));
 sg13g2_a21oi_1 _6254_ (.A1(net857),
    .A2(_2487_),
    .Y(_0400_),
    .B1(_2492_));
 sg13g2_nor2_1 _6255_ (.A(net1034),
    .B(net832),
    .Y(_2493_));
 sg13g2_a21oi_1 _6256_ (.A1(net860),
    .A2(net832),
    .Y(_0401_),
    .B1(_2493_));
 sg13g2_nor2_1 _6257_ (.A(net1133),
    .B(net831),
    .Y(_2494_));
 sg13g2_a21oi_1 _6258_ (.A1(net854),
    .A2(net832),
    .Y(_0402_),
    .B1(_2494_));
 sg13g2_nor2_1 _6259_ (.A(net1084),
    .B(net831),
    .Y(_2495_));
 sg13g2_a21oi_1 _6260_ (.A1(net851),
    .A2(net831),
    .Y(_0403_),
    .B1(_2495_));
 sg13g2_or2_2 _6261_ (.X(_2496_),
    .B(_2485_),
    .A(_2259_));
 sg13g2_mux2_1 _6262_ (.A0(net776),
    .A1(net1274),
    .S(_2496_),
    .X(_0404_));
 sg13g2_mux2_1 _6263_ (.A0(net774),
    .A1(net1276),
    .S(_2496_),
    .X(_0405_));
 sg13g2_mux2_1 _6264_ (.A0(net773),
    .A1(net1233),
    .S(_2496_),
    .X(_0406_));
 sg13g2_mux2_1 _6265_ (.A0(net761),
    .A1(net1240),
    .S(_2496_),
    .X(_0407_));
 sg13g2_mux2_1 _6266_ (.A0(net766),
    .A1(net1260),
    .S(_2496_),
    .X(_0408_));
 sg13g2_mux2_1 _6267_ (.A0(net764),
    .A1(net1460),
    .S(_2496_),
    .X(_0409_));
 sg13g2_mux2_1 _6268_ (.A0(net759),
    .A1(net1455),
    .S(_2496_),
    .X(_0410_));
 sg13g2_mux2_1 _6269_ (.A0(net757),
    .A1(net1454),
    .S(_2496_),
    .X(_0411_));
 sg13g2_nand3_1 _6270_ (.B(_0687_),
    .C(_2303_),
    .A(_0686_),
    .Y(_2497_));
 sg13g2_nand2_1 _6271_ (.Y(_2498_),
    .A(net744),
    .B(net829));
 sg13g2_o21ai_1 _6272_ (.B1(_2498_),
    .Y(_0412_),
    .A1(net873),
    .A2(net829));
 sg13g2_nand2_1 _6273_ (.Y(_2499_),
    .A(net1162),
    .B(net829));
 sg13g2_o21ai_1 _6274_ (.B1(_2499_),
    .Y(_0413_),
    .A1(net870),
    .A2(net829));
 sg13g2_nand2_1 _6275_ (.Y(_2500_),
    .A(net1021),
    .B(net830));
 sg13g2_o21ai_1 _6276_ (.B1(_2500_),
    .Y(_0414_),
    .A1(net867),
    .A2(net830));
 sg13g2_nand2_1 _6277_ (.Y(_2501_),
    .A(net1023),
    .B(net830));
 sg13g2_o21ai_1 _6278_ (.B1(_2501_),
    .Y(_0415_),
    .A1(net864),
    .A2(net830));
 sg13g2_nand2_1 _6279_ (.Y(_2502_),
    .A(net1033),
    .B(net830));
 sg13g2_o21ai_1 _6280_ (.B1(_2502_),
    .Y(_0416_),
    .A1(net857),
    .A2(net830));
 sg13g2_nand2_1 _6281_ (.Y(_2503_),
    .A(net1004),
    .B(net829));
 sg13g2_o21ai_1 _6282_ (.B1(_2503_),
    .Y(_0417_),
    .A1(net861),
    .A2(net829));
 sg13g2_nand2_1 _6283_ (.Y(_2504_),
    .A(net1022),
    .B(net830));
 sg13g2_o21ai_1 _6284_ (.B1(_2504_),
    .Y(_0418_),
    .A1(net855),
    .A2(net830));
 sg13g2_nand2_1 _6285_ (.Y(_2505_),
    .A(net749),
    .B(net829));
 sg13g2_o21ai_1 _6286_ (.B1(_2505_),
    .Y(_0419_),
    .A1(net850),
    .A2(net829));
 sg13g2_nor2_2 _6287_ (.A(_2316_),
    .B(_2318_),
    .Y(_2506_));
 sg13g2_mux2_1 _6288_ (.A0(net1078),
    .A1(net776),
    .S(_2506_),
    .X(_0420_));
 sg13g2_mux2_1 _6289_ (.A0(net1052),
    .A1(net774),
    .S(_2506_),
    .X(_0421_));
 sg13g2_mux2_1 _6290_ (.A0(net1085),
    .A1(net772),
    .S(_2506_),
    .X(_0422_));
 sg13g2_mux2_1 _6291_ (.A0(net1073),
    .A1(net761),
    .S(_2506_),
    .X(_0423_));
 sg13g2_mux2_1 _6292_ (.A0(net1057),
    .A1(net766),
    .S(_2506_),
    .X(_0424_));
 sg13g2_mux2_1 _6293_ (.A0(net1205),
    .A1(net764),
    .S(_2506_),
    .X(_0425_));
 sg13g2_mux2_1 _6294_ (.A0(net1249),
    .A1(net759),
    .S(_2506_),
    .X(_0426_));
 sg13g2_mux2_1 _6295_ (.A0(net1197),
    .A1(net757),
    .S(_2506_),
    .X(_0427_));
 sg13g2_nor2_2 _6296_ (.A(_2318_),
    .B(_2485_),
    .Y(_2507_));
 sg13g2_mux2_1 _6297_ (.A0(net1058),
    .A1(net776),
    .S(_2507_),
    .X(_0428_));
 sg13g2_mux2_1 _6298_ (.A0(net1055),
    .A1(net774),
    .S(_2507_),
    .X(_0429_));
 sg13g2_mux2_1 _6299_ (.A0(net1064),
    .A1(net773),
    .S(_2507_),
    .X(_0430_));
 sg13g2_mux2_1 _6300_ (.A0(net1038),
    .A1(net761),
    .S(_2507_),
    .X(_0431_));
 sg13g2_mux2_1 _6301_ (.A0(net1063),
    .A1(net766),
    .S(_2507_),
    .X(_0432_));
 sg13g2_mux2_1 _6302_ (.A0(net1219),
    .A1(net764),
    .S(_2507_),
    .X(_0433_));
 sg13g2_mux2_1 _6303_ (.A0(net1275),
    .A1(net759),
    .S(_2507_),
    .X(_0434_));
 sg13g2_mux2_1 _6304_ (.A0(net1342),
    .A1(net757),
    .S(_2507_),
    .X(_0435_));
 sg13g2_or2_2 _6305_ (.X(_2508_),
    .B(_2319_),
    .A(_2314_));
 sg13g2_mux2_1 _6306_ (.A0(net777),
    .A1(net1326),
    .S(_2508_),
    .X(_0436_));
 sg13g2_mux2_1 _6307_ (.A0(net775),
    .A1(net1307),
    .S(_2508_),
    .X(_0437_));
 sg13g2_mux2_1 _6308_ (.A0(net772),
    .A1(net1296),
    .S(_2508_),
    .X(_0438_));
 sg13g2_mux2_1 _6309_ (.A0(net762),
    .A1(net1345),
    .S(_2508_),
    .X(_0439_));
 sg13g2_mux2_1 _6310_ (.A0(net767),
    .A1(net1324),
    .S(_2508_),
    .X(_0440_));
 sg13g2_mux2_1 _6311_ (.A0(net765),
    .A1(net1327),
    .S(_2508_),
    .X(_0441_));
 sg13g2_mux2_1 _6312_ (.A0(net760),
    .A1(net1363),
    .S(_2508_),
    .X(_0442_));
 sg13g2_mux2_1 _6313_ (.A0(net758),
    .A1(net1343),
    .S(_2508_),
    .X(_0443_));
 sg13g2_or2_2 _6314_ (.X(_2509_),
    .B(_2319_),
    .A(_2259_));
 sg13g2_mux2_1 _6315_ (.A0(net777),
    .A1(net1318),
    .S(_2509_),
    .X(_0444_));
 sg13g2_mux2_1 _6316_ (.A0(net775),
    .A1(net1308),
    .S(_2509_),
    .X(_0445_));
 sg13g2_mux2_1 _6317_ (.A0(net772),
    .A1(net1270),
    .S(_2509_),
    .X(_0446_));
 sg13g2_mux2_1 _6318_ (.A0(net762),
    .A1(net1289),
    .S(_2509_),
    .X(_0447_));
 sg13g2_mux2_1 _6319_ (.A0(net767),
    .A1(net1319),
    .S(_2509_),
    .X(_0448_));
 sg13g2_mux2_1 _6320_ (.A0(net765),
    .A1(net1488),
    .S(_2509_),
    .X(_0449_));
 sg13g2_mux2_1 _6321_ (.A0(net760),
    .A1(net1464),
    .S(_2509_),
    .X(_0450_));
 sg13g2_mux2_1 _6322_ (.A0(net758),
    .A1(net1502),
    .S(_2509_),
    .X(_0451_));
 sg13g2_nor4_2 _6323_ (.A(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[3] ),
    .B(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[2] ),
    .C(_2243_),
    .Y(_2510_),
    .D(_2244_));
 sg13g2_nor2_1 _6324_ (.A(net1136),
    .B(net876),
    .Y(_2511_));
 sg13g2_a21oi_1 _6325_ (.A1(net873),
    .A2(net876),
    .Y(_0452_),
    .B1(_2511_));
 sg13g2_nor2_1 _6326_ (.A(net1212),
    .B(net877),
    .Y(_2512_));
 sg13g2_a21oi_1 _6327_ (.A1(net870),
    .A2(net877),
    .Y(_0453_),
    .B1(_2512_));
 sg13g2_nor2_1 _6328_ (.A(net1210),
    .B(_2510_),
    .Y(_2513_));
 sg13g2_a21oi_1 _6329_ (.A1(net867),
    .A2(net876),
    .Y(_0454_),
    .B1(net1211));
 sg13g2_nor2_1 _6330_ (.A(net1280),
    .B(net876),
    .Y(_2514_));
 sg13g2_a21oi_1 _6331_ (.A1(net864),
    .A2(net876),
    .Y(_0455_),
    .B1(_2514_));
 sg13g2_nor2_1 _6332_ (.A(net1336),
    .B(net876),
    .Y(_2515_));
 sg13g2_a21oi_1 _6333_ (.A1(net857),
    .A2(net877),
    .Y(_0456_),
    .B1(_2515_));
 sg13g2_nor2_1 _6334_ (.A(net1134),
    .B(net877),
    .Y(_2516_));
 sg13g2_a21oi_1 _6335_ (.A1(net861),
    .A2(net877),
    .Y(_0457_),
    .B1(_2516_));
 sg13g2_nor2_1 _6336_ (.A(net1255),
    .B(net876),
    .Y(_2517_));
 sg13g2_a21oi_1 _6337_ (.A1(net855),
    .A2(net876),
    .Y(_0458_),
    .B1(_2517_));
 sg13g2_nor2_1 _6338_ (.A(net1163),
    .B(net877),
    .Y(_2518_));
 sg13g2_a21oi_1 _6339_ (.A1(net850),
    .A2(net877),
    .Y(_0459_),
    .B1(_2518_));
 sg13g2_nor3_1 _6340_ (.A(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[3] ),
    .B(net991),
    .C(_2368_),
    .Y(_2519_));
 sg13g2_nor2_1 _6341_ (.A(net1086),
    .B(net827),
    .Y(_2520_));
 sg13g2_a21oi_1 _6342_ (.A1(net873),
    .A2(net827),
    .Y(_0460_),
    .B1(_2520_));
 sg13g2_nor2_1 _6343_ (.A(net1145),
    .B(net828),
    .Y(_2521_));
 sg13g2_a21oi_1 _6344_ (.A1(net870),
    .A2(net828),
    .Y(_0461_),
    .B1(_2521_));
 sg13g2_nor2_1 _6345_ (.A(net1349),
    .B(_2519_),
    .Y(_2522_));
 sg13g2_a21oi_1 _6346_ (.A1(net867),
    .A2(net827),
    .Y(_0462_),
    .B1(net1350));
 sg13g2_nor2_1 _6347_ (.A(net1125),
    .B(net827),
    .Y(_2523_));
 sg13g2_a21oi_1 _6348_ (.A1(net864),
    .A2(net827),
    .Y(_0463_),
    .B1(_2523_));
 sg13g2_nor2_1 _6349_ (.A(net1137),
    .B(net827),
    .Y(_2524_));
 sg13g2_a21oi_1 _6350_ (.A1(net857),
    .A2(net828),
    .Y(_0464_),
    .B1(_2524_));
 sg13g2_nor2_1 _6351_ (.A(net1066),
    .B(net828),
    .Y(_2525_));
 sg13g2_a21oi_1 _6352_ (.A1(net861),
    .A2(net828),
    .Y(_0465_),
    .B1(_2525_));
 sg13g2_nor2_1 _6353_ (.A(net1298),
    .B(net827),
    .Y(_2526_));
 sg13g2_a21oi_1 _6354_ (.A1(net855),
    .A2(net827),
    .Y(_0466_),
    .B1(_2526_));
 sg13g2_nor2_1 _6355_ (.A(net1024),
    .B(net828),
    .Y(_2527_));
 sg13g2_a21oi_1 _6356_ (.A1(net850),
    .A2(net828),
    .Y(_0467_),
    .B1(_2527_));
 sg13g2_nor2_1 _6357_ (.A(net1046),
    .B(net821),
    .Y(_2528_));
 sg13g2_a21oi_1 _6358_ (.A1(net872),
    .A2(net821),
    .Y(_0468_),
    .B1(_2528_));
 sg13g2_nor2_1 _6359_ (.A(net1301),
    .B(net821),
    .Y(_2529_));
 sg13g2_a21oi_1 _6360_ (.A1(net869),
    .A2(net821),
    .Y(_0469_),
    .B1(_2529_));
 sg13g2_nor2_1 _6361_ (.A(net1202),
    .B(net821),
    .Y(_2530_));
 sg13g2_a21oi_1 _6362_ (.A1(net866),
    .A2(net821),
    .Y(_0470_),
    .B1(_2530_));
 sg13g2_nor2_1 _6363_ (.A(net1189),
    .B(net821),
    .Y(_2531_));
 sg13g2_a21oi_1 _6364_ (.A1(net863),
    .A2(net821),
    .Y(_0471_),
    .B1(_2531_));
 sg13g2_nor2_1 _6365_ (.A(net1370),
    .B(net820),
    .Y(_2532_));
 sg13g2_a21oi_1 _6366_ (.A1(net858),
    .A2(net820),
    .Y(_0472_),
    .B1(_2532_));
 sg13g2_nor2_1 _6367_ (.A(net1032),
    .B(net820),
    .Y(_2533_));
 sg13g2_a21oi_1 _6368_ (.A1(net860),
    .A2(net820),
    .Y(_0473_),
    .B1(_2533_));
 sg13g2_nor2_1 _6369_ (.A(net1203),
    .B(net820),
    .Y(_2534_));
 sg13g2_a21oi_1 _6370_ (.A1(net854),
    .A2(net820),
    .Y(_0474_),
    .B1(_2534_));
 sg13g2_nor2_1 _6371_ (.A(net1138),
    .B(net820),
    .Y(_2535_));
 sg13g2_a21oi_1 _6372_ (.A1(net850),
    .A2(net820),
    .Y(_0475_),
    .B1(_2535_));
 sg13g2_or2_2 _6373_ (.X(_2536_),
    .B(_2332_),
    .A(_2319_));
 sg13g2_mux2_1 _6374_ (.A0(net777),
    .A1(net1321),
    .S(_2536_),
    .X(_0476_));
 sg13g2_mux2_1 _6375_ (.A0(net775),
    .A1(net1269),
    .S(_2536_),
    .X(_0477_));
 sg13g2_mux2_1 _6376_ (.A0(net772),
    .A1(net1325),
    .S(_2536_),
    .X(_0478_));
 sg13g2_mux2_1 _6377_ (.A0(net762),
    .A1(net1315),
    .S(_2536_),
    .X(_0479_));
 sg13g2_mux2_1 _6378_ (.A0(net767),
    .A1(net1291),
    .S(_2536_),
    .X(_0480_));
 sg13g2_mux2_1 _6379_ (.A0(net765),
    .A1(net1401),
    .S(_2536_),
    .X(_0481_));
 sg13g2_mux2_1 _6380_ (.A0(net760),
    .A1(net1410),
    .S(_2536_),
    .X(_0482_));
 sg13g2_mux2_1 _6381_ (.A0(net758),
    .A1(net1467),
    .S(_2536_),
    .X(_0483_));
 sg13g2_or2_2 _6382_ (.X(_2537_),
    .B(_2485_),
    .A(_2332_));
 sg13g2_mux2_1 _6383_ (.A0(net776),
    .A1(net1281),
    .S(_2537_),
    .X(_0484_));
 sg13g2_mux2_1 _6384_ (.A0(net774),
    .A1(net1285),
    .S(_2537_),
    .X(_0485_));
 sg13g2_mux2_1 _6385_ (.A0(net773),
    .A1(net1228),
    .S(_2537_),
    .X(_0486_));
 sg13g2_mux2_1 _6386_ (.A0(net761),
    .A1(net1242),
    .S(_2537_),
    .X(_0487_));
 sg13g2_mux2_1 _6387_ (.A0(net766),
    .A1(net1292),
    .S(_2537_),
    .X(_0488_));
 sg13g2_mux2_1 _6388_ (.A0(net764),
    .A1(net1469),
    .S(_2537_),
    .X(_0489_));
 sg13g2_mux2_1 _6389_ (.A0(net759),
    .A1(net1456),
    .S(_2537_),
    .X(_0490_));
 sg13g2_mux2_1 _6390_ (.A0(net757),
    .A1(net1468),
    .S(_2537_),
    .X(_0491_));
 sg13g2_a21oi_1 _6391_ (.A1(net1545),
    .A2(net768),
    .Y(_0492_),
    .B1(net963));
 sg13g2_xor2_1 _6392_ (.B(net1689),
    .A(net1545),
    .X(_2538_));
 sg13g2_a21oi_1 _6393_ (.A1(net768),
    .A2(_2538_),
    .Y(_0493_),
    .B1(net963));
 sg13g2_o21ai_1 _6394_ (.B1(net1734),
    .Y(_2539_),
    .A1(\C1.counter2[0] ),
    .A2(\C1.counter2[1] ));
 sg13g2_nor2b_1 _6395_ (.A(_1756_),
    .B_N(_2539_),
    .Y(_2540_));
 sg13g2_a21oi_1 _6396_ (.A1(net768),
    .A2(net1735),
    .Y(_0494_),
    .B1(net964));
 sg13g2_xnor2_1 _6397_ (.Y(_2541_),
    .A(net1647),
    .B(_1756_));
 sg13g2_a21oi_1 _6398_ (.A1(net768),
    .A2(net1648),
    .Y(_0495_),
    .B1(net963));
 sg13g2_xnor2_1 _6399_ (.Y(_2542_),
    .A(net1604),
    .B(_1757_));
 sg13g2_a21oi_1 _6400_ (.A1(net770),
    .A2(net1605),
    .Y(_0496_),
    .B1(net963));
 sg13g2_xnor2_1 _6401_ (.Y(_2543_),
    .A(net1634),
    .B(_1758_));
 sg13g2_a21oi_1 _6402_ (.A1(net770),
    .A2(_2543_),
    .Y(_0497_),
    .B1(net964));
 sg13g2_xnor2_1 _6403_ (.Y(_2544_),
    .A(net1600),
    .B(_1759_));
 sg13g2_a21oi_1 _6404_ (.A1(net771),
    .A2(net1601),
    .Y(_0498_),
    .B1(net964));
 sg13g2_xor2_1 _6405_ (.B(_1760_),
    .A(net1685),
    .X(_2545_));
 sg13g2_a21oi_1 _6406_ (.A1(net768),
    .A2(_2545_),
    .Y(_0499_),
    .B1(net964));
 sg13g2_xor2_1 _6407_ (.B(_1761_),
    .A(net1683),
    .X(_2546_));
 sg13g2_a21oi_1 _6408_ (.A1(net771),
    .A2(_2546_),
    .Y(_0500_),
    .B1(net964));
 sg13g2_o21ai_1 _6409_ (.B1(net1706),
    .Y(_2547_),
    .A1(net1683),
    .A2(_1761_));
 sg13g2_nor2b_1 _6410_ (.A(_1762_),
    .B_N(_2547_),
    .Y(_2548_));
 sg13g2_a21oi_1 _6411_ (.A1(net768),
    .A2(_2548_),
    .Y(_0501_),
    .B1(net964));
 sg13g2_xnor2_1 _6412_ (.Y(_2549_),
    .A(net1624),
    .B(_1762_));
 sg13g2_a21oi_1 _6413_ (.A1(net770),
    .A2(net1625),
    .Y(_0502_),
    .B1(net963));
 sg13g2_xor2_1 _6414_ (.B(_1763_),
    .A(net1681),
    .X(_2550_));
 sg13g2_a21oi_1 _6415_ (.A1(net768),
    .A2(net1682),
    .Y(_0503_),
    .B1(net963));
 sg13g2_o21ai_1 _6416_ (.B1(net1712),
    .Y(_2551_),
    .A1(\C1.counter2[11] ),
    .A2(_1763_));
 sg13g2_nor2b_1 _6417_ (.A(net1713),
    .B_N(_2551_),
    .Y(_2552_));
 sg13g2_a21oi_1 _6418_ (.A1(net768),
    .A2(net1714),
    .Y(_0504_),
    .B1(net963));
 sg13g2_xnor2_1 _6419_ (.Y(_2553_),
    .A(net1584),
    .B(_1764_));
 sg13g2_a21oi_1 _6420_ (.A1(net769),
    .A2(net1585),
    .Y(_0505_),
    .B1(net963));
 sg13g2_xor2_1 _6421_ (.B(_1765_),
    .A(net1694),
    .X(_2554_));
 sg13g2_a21oi_1 _6422_ (.A1(net769),
    .A2(net1695),
    .Y(_0506_),
    .B1(net965));
 sg13g2_o21ai_1 _6423_ (.B1(net1715),
    .Y(_2555_),
    .A1(\C1.counter2[14] ),
    .A2(_1765_));
 sg13g2_nor2b_1 _6424_ (.A(net1716),
    .B_N(_2555_),
    .Y(_2556_));
 sg13g2_a21oi_1 _6425_ (.A1(net769),
    .A2(net1717),
    .Y(_0507_),
    .B1(net965));
 sg13g2_xnor2_1 _6426_ (.Y(_2557_),
    .A(net1591),
    .B(_1766_));
 sg13g2_a21oi_1 _6427_ (.A1(net769),
    .A2(net1592),
    .Y(_0508_),
    .B1(net965));
 sg13g2_xor2_1 _6428_ (.B(_1767_),
    .A(net1696),
    .X(_2558_));
 sg13g2_a21oi_1 _6429_ (.A1(net771),
    .A2(net1697),
    .Y(_0509_),
    .B1(net965));
 sg13g2_o21ai_1 _6430_ (.B1(net1702),
    .Y(_2559_),
    .A1(net1696),
    .A2(_1767_));
 sg13g2_nor2b_1 _6431_ (.A(net1703),
    .B_N(_2559_),
    .Y(_2560_));
 sg13g2_a21oi_1 _6432_ (.A1(net769),
    .A2(_2560_),
    .Y(_0510_),
    .B1(net965));
 sg13g2_xnor2_1 _6433_ (.Y(_2561_),
    .A(net1576),
    .B(_1768_));
 sg13g2_a21oi_1 _6434_ (.A1(net769),
    .A2(net1577),
    .Y(_0511_),
    .B1(net965));
 sg13g2_xor2_1 _6435_ (.B(_1769_),
    .A(net1672),
    .X(_2562_));
 sg13g2_a21oi_1 _6436_ (.A1(net769),
    .A2(net1673),
    .Y(_0512_),
    .B1(net965));
 sg13g2_o21ai_1 _6437_ (.B1(net1704),
    .Y(_2563_),
    .A1(\C1.counter2[20] ),
    .A2(_1769_));
 sg13g2_nor2b_1 _6438_ (.A(_1770_),
    .B_N(_2563_),
    .Y(_2564_));
 sg13g2_a21oi_1 _6439_ (.A1(net769),
    .A2(net1705),
    .Y(_0513_),
    .B1(net965));
 sg13g2_nor2_1 _6440_ (.A(_2243_),
    .B(_2358_),
    .Y(_2565_));
 sg13g2_nor2_1 _6441_ (.A(net1047),
    .B(net826),
    .Y(_2566_));
 sg13g2_a21oi_1 _6442_ (.A1(net872),
    .A2(_2565_),
    .Y(_0514_),
    .B1(_2566_));
 sg13g2_nor2_1 _6443_ (.A(net1224),
    .B(net825),
    .Y(_2567_));
 sg13g2_a21oi_1 _6444_ (.A1(net869),
    .A2(net825),
    .Y(_0515_),
    .B1(_2567_));
 sg13g2_nor2_1 _6445_ (.A(net1214),
    .B(net825),
    .Y(_2568_));
 sg13g2_a21oi_1 _6446_ (.A1(net866),
    .A2(net825),
    .Y(_0516_),
    .B1(_2568_));
 sg13g2_nor2_1 _6447_ (.A(net1257),
    .B(net825),
    .Y(_2569_));
 sg13g2_a21oi_1 _6448_ (.A1(net863),
    .A2(net825),
    .Y(_0517_),
    .B1(_2569_));
 sg13g2_nor2_1 _6449_ (.A(net1268),
    .B(net825),
    .Y(_2570_));
 sg13g2_a21oi_1 _6450_ (.A1(net856),
    .A2(net825),
    .Y(_0518_),
    .B1(_2570_));
 sg13g2_nor2_1 _6451_ (.A(net1090),
    .B(net826),
    .Y(_2571_));
 sg13g2_a21oi_1 _6452_ (.A1(net862),
    .A2(net826),
    .Y(_0519_),
    .B1(_2571_));
 sg13g2_nor2_1 _6453_ (.A(net1216),
    .B(net826),
    .Y(_2572_));
 sg13g2_a21oi_1 _6454_ (.A1(net853),
    .A2(net826),
    .Y(_0520_),
    .B1(_2572_));
 sg13g2_nor2_1 _6455_ (.A(net1101),
    .B(net826),
    .Y(_2573_));
 sg13g2_a21oi_1 _6456_ (.A1(net850),
    .A2(net826),
    .Y(_0521_),
    .B1(_2573_));
 sg13g2_nand3_1 _6457_ (.B(net1387),
    .C(net1243),
    .A(\FpgaPins_Fpga_GAME_wait_counter_a2[14] ),
    .Y(_2574_));
 sg13g2_a21o_1 _6458_ (.A2(_2424_),
    .A1(_2422_),
    .B1(_2574_),
    .X(_2575_));
 sg13g2_a21oi_1 _6459_ (.A1(_2426_),
    .A2(_2575_),
    .Y(_2576_),
    .B1(_0726_));
 sg13g2_nor3_1 _6460_ (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[21] ),
    .B(\FpgaPins_Fpga_GAME_wait_counter_a2[20] ),
    .C(_2576_),
    .Y(_2577_));
 sg13g2_nor2_1 _6461_ (.A(net1755),
    .B(_2427_),
    .Y(_2578_));
 sg13g2_o21ai_1 _6462_ (.B1(_2578_),
    .Y(_2579_),
    .A1(_2425_),
    .A2(_2577_));
 sg13g2_inv_2 _6463_ (.Y(_2580_),
    .A(_2579_));
 sg13g2_and2_1 _6464_ (.A(net709),
    .B(_2580_),
    .X(_0522_));
 sg13g2_xnor2_1 _6465_ (.Y(_2581_),
    .A(\FpgaPins_Fpga_GAME_wait_counter_a2[0] ),
    .B(net1538));
 sg13g2_nor2_1 _6466_ (.A(net901),
    .B(net1539),
    .Y(_0523_));
 sg13g2_and3_1 _6467_ (.X(_2582_),
    .A(\FpgaPins_Fpga_GAME_wait_counter_a2[0] ),
    .B(\FpgaPins_Fpga_GAME_wait_counter_a2[1] ),
    .C(net1175));
 sg13g2_a21oi_1 _6468_ (.A1(\FpgaPins_Fpga_GAME_wait_counter_a2[0] ),
    .A2(\FpgaPins_Fpga_GAME_wait_counter_a2[1] ),
    .Y(_2583_),
    .B1(net1175));
 sg13g2_nor3_1 _6469_ (.A(net901),
    .B(_2582_),
    .C(net1176),
    .Y(_0524_));
 sg13g2_and2_1 _6470_ (.A(net1480),
    .B(_2582_),
    .X(_2584_));
 sg13g2_nor2_1 _6471_ (.A(net1480),
    .B(_2582_),
    .Y(_2585_));
 sg13g2_nor3_1 _6472_ (.A(net901),
    .B(_2584_),
    .C(net1481),
    .Y(_0525_));
 sg13g2_and2_1 _6473_ (.A(net1501),
    .B(_2584_),
    .X(_2586_));
 sg13g2_nor2_1 _6474_ (.A(net1501),
    .B(_2584_),
    .Y(_2587_));
 sg13g2_nor3_1 _6475_ (.A(net901),
    .B(_2586_),
    .C(_2587_),
    .Y(_0526_));
 sg13g2_and2_1 _6476_ (.A(net1482),
    .B(_2586_),
    .X(_2588_));
 sg13g2_nor2_1 _6477_ (.A(net1482),
    .B(_2586_),
    .Y(_2589_));
 sg13g2_nor3_1 _6478_ (.A(net901),
    .B(_2588_),
    .C(net1483),
    .Y(_0527_));
 sg13g2_and2_1 _6479_ (.A(net1375),
    .B(_2588_),
    .X(_2590_));
 sg13g2_nor2_1 _6480_ (.A(net1375),
    .B(_2588_),
    .Y(_2591_));
 sg13g2_nor3_1 _6481_ (.A(net900),
    .B(_2590_),
    .C(net1376),
    .Y(_0528_));
 sg13g2_and2_1 _6482_ (.A(net1504),
    .B(_2590_),
    .X(_2592_));
 sg13g2_nor2_1 _6483_ (.A(net1504),
    .B(_2590_),
    .Y(_2593_));
 sg13g2_nor3_1 _6484_ (.A(net899),
    .B(_2592_),
    .C(_2593_),
    .Y(_0529_));
 sg13g2_and2_1 _6485_ (.A(net1638),
    .B(_2592_),
    .X(_2594_));
 sg13g2_o21ai_1 _6486_ (.B1(_2580_),
    .Y(_2595_),
    .A1(net1638),
    .A2(_2592_));
 sg13g2_nor2_1 _6487_ (.A(_2594_),
    .B(net1639),
    .Y(_0530_));
 sg13g2_nor2_1 _6488_ (.A(net1524),
    .B(_2594_),
    .Y(_2596_));
 sg13g2_nor2b_1 _6489_ (.A(_2424_),
    .B_N(_2590_),
    .Y(_2597_));
 sg13g2_nor3_1 _6490_ (.A(net899),
    .B(net1525),
    .C(_2597_),
    .Y(_0531_));
 sg13g2_nor2_1 _6491_ (.A(net1602),
    .B(_2597_),
    .Y(_2598_));
 sg13g2_and2_1 _6492_ (.A(net1602),
    .B(_2597_),
    .X(_2599_));
 sg13g2_nor3_1 _6493_ (.A(net899),
    .B(net1603),
    .C(_2599_),
    .Y(_0532_));
 sg13g2_and4_1 _6494_ (.A(net1524),
    .B(net1602),
    .C(net1644),
    .D(_2594_),
    .X(_2600_));
 sg13g2_o21ai_1 _6495_ (.B1(_2580_),
    .Y(_2601_),
    .A1(net1644),
    .A2(_2599_));
 sg13g2_nor2_1 _6496_ (.A(_2600_),
    .B(net1645),
    .Y(_0533_));
 sg13g2_nor2_1 _6497_ (.A(net1529),
    .B(_2600_),
    .Y(_2602_));
 sg13g2_and3_1 _6498_ (.X(_2603_),
    .A(\FpgaPins_Fpga_GAME_wait_counter_a2[11] ),
    .B(net1529),
    .C(_2599_));
 sg13g2_nor3_1 _6499_ (.A(net899),
    .B(net1530),
    .C(_2603_),
    .Y(_0534_));
 sg13g2_or2_1 _6500_ (.X(_2604_),
    .B(_2603_),
    .A(net1722));
 sg13g2_nand3_1 _6501_ (.B(net1529),
    .C(_2600_),
    .A(net1722),
    .Y(_2605_));
 sg13g2_and3_1 _6502_ (.X(_0535_),
    .A(_2580_),
    .B(net1723),
    .C(_2605_));
 sg13g2_a21oi_1 _6503_ (.A1(\FpgaPins_Fpga_GAME_wait_counter_a2[13] ),
    .A2(_2603_),
    .Y(_2606_),
    .B1(net1495));
 sg13g2_nor2_2 _6504_ (.A(_0725_),
    .B(_2605_),
    .Y(_2607_));
 sg13g2_nor3_1 _6505_ (.A(net901),
    .B(net1496),
    .C(_2607_),
    .Y(_0536_));
 sg13g2_o21ai_1 _6506_ (.B1(_2580_),
    .Y(_2608_),
    .A1(net1387),
    .A2(_2607_));
 sg13g2_a21oi_1 _6507_ (.A1(net1387),
    .A2(_2607_),
    .Y(_0537_),
    .B1(_2608_));
 sg13g2_a21oi_1 _6508_ (.A1(\FpgaPins_Fpga_GAME_wait_counter_a2[15] ),
    .A2(_2607_),
    .Y(_2609_),
    .B1(net1243));
 sg13g2_nor2_1 _6509_ (.A(_2574_),
    .B(_2605_),
    .Y(_2610_));
 sg13g2_nor3_1 _6510_ (.A(net899),
    .B(net1244),
    .C(_2610_),
    .Y(_0538_));
 sg13g2_nor2_1 _6511_ (.A(net1448),
    .B(_2610_),
    .Y(_2611_));
 sg13g2_and2_1 _6512_ (.A(net1448),
    .B(_2610_),
    .X(_2612_));
 sg13g2_nor3_1 _6513_ (.A(net899),
    .B(net1449),
    .C(_2612_),
    .Y(_0539_));
 sg13g2_nor2_1 _6514_ (.A(net1451),
    .B(_2612_),
    .Y(_2613_));
 sg13g2_and2_1 _6515_ (.A(net1451),
    .B(_2612_),
    .X(_2614_));
 sg13g2_nor3_1 _6516_ (.A(net900),
    .B(_2613_),
    .C(_2614_),
    .Y(_0540_));
 sg13g2_nor2_1 _6517_ (.A(net1548),
    .B(_2614_),
    .Y(_2615_));
 sg13g2_and2_1 _6518_ (.A(net1548),
    .B(_2614_),
    .X(_2616_));
 sg13g2_nor3_1 _6519_ (.A(net900),
    .B(_2615_),
    .C(_2616_),
    .Y(_0541_));
 sg13g2_nor2_1 _6520_ (.A(net1536),
    .B(_2616_),
    .Y(_2617_));
 sg13g2_and2_1 _6521_ (.A(net1536),
    .B(_2616_),
    .X(_2618_));
 sg13g2_nor3_1 _6522_ (.A(net900),
    .B(net1537),
    .C(_2618_),
    .Y(_0542_));
 sg13g2_nor2_1 _6523_ (.A(net1597),
    .B(_2618_),
    .Y(_2619_));
 sg13g2_and2_1 _6524_ (.A(net1597),
    .B(_2618_),
    .X(_2620_));
 sg13g2_nor3_1 _6525_ (.A(net900),
    .B(_2619_),
    .C(_2620_),
    .Y(_0543_));
 sg13g2_nor2_1 _6526_ (.A(net1567),
    .B(_2620_),
    .Y(_2621_));
 sg13g2_and2_1 _6527_ (.A(net1567),
    .B(_2620_),
    .X(_2622_));
 sg13g2_nor3_1 _6528_ (.A(net899),
    .B(net1568),
    .C(_2622_),
    .Y(_0544_));
 sg13g2_o21ai_1 _6529_ (.B1(_2580_),
    .Y(_2623_),
    .A1(net1412),
    .A2(_2622_));
 sg13g2_a21oi_1 _6530_ (.A1(net1412),
    .A2(_2622_),
    .Y(_0545_),
    .B1(_2623_));
 sg13g2_a21oi_1 _6531_ (.A1(\FpgaPins_Fpga_GAME_wait_counter_a2[23] ),
    .A2(_2622_),
    .Y(_2624_),
    .B1(net1107));
 sg13g2_nor2_1 _6532_ (.A(net899),
    .B(net1108),
    .Y(_0546_));
 sg13g2_nor3_1 _6533_ (.A(_0686_),
    .B(net991),
    .C(_2368_),
    .Y(_2625_));
 sg13g2_nor2_1 _6534_ (.A(net1140),
    .B(net823),
    .Y(_2626_));
 sg13g2_a21oi_1 _6535_ (.A1(net874),
    .A2(net823),
    .Y(_0547_),
    .B1(_2626_));
 sg13g2_nor2_1 _6536_ (.A(net1218),
    .B(net823),
    .Y(_2627_));
 sg13g2_a21oi_1 _6537_ (.A1(net871),
    .A2(net823),
    .Y(_0548_),
    .B1(_2627_));
 sg13g2_nor2_1 _6538_ (.A(net1209),
    .B(net824),
    .Y(_2628_));
 sg13g2_a21oi_1 _6539_ (.A1(net866),
    .A2(net824),
    .Y(_0549_),
    .B1(_2628_));
 sg13g2_nor2_1 _6540_ (.A(net1184),
    .B(net824),
    .Y(_2629_));
 sg13g2_a21oi_1 _6541_ (.A1(net863),
    .A2(net824),
    .Y(_0550_),
    .B1(_2629_));
 sg13g2_nor2_1 _6542_ (.A(net1119),
    .B(net824),
    .Y(_2630_));
 sg13g2_a21oi_1 _6543_ (.A1(net856),
    .A2(_2625_),
    .Y(_0551_),
    .B1(_2630_));
 sg13g2_nor2_1 _6544_ (.A(net1070),
    .B(net824),
    .Y(_2631_));
 sg13g2_a21oi_1 _6545_ (.A1(net860),
    .A2(net823),
    .Y(_0552_),
    .B1(_2631_));
 sg13g2_nor2_1 _6546_ (.A(net1407),
    .B(net824),
    .Y(_2632_));
 sg13g2_a21oi_1 _6547_ (.A1(net853),
    .A2(net823),
    .Y(_0553_),
    .B1(_2632_));
 sg13g2_nor2_1 _6548_ (.A(net1029),
    .B(net823),
    .Y(_2633_));
 sg13g2_a21oi_1 _6549_ (.A1(net852),
    .A2(net823),
    .Y(_0554_),
    .B1(_2633_));
 sg13g2_nand3b_1 _6550_ (.B(net994),
    .C(_1739_),
    .Y(_2634_),
    .A_N(_2125_));
 sg13g2_o21ai_1 _6551_ (.B1(_1735_),
    .Y(_2635_),
    .A1(_0015_),
    .A2(_1739_));
 sg13g2_nor2b_1 _6552_ (.A(_2635_),
    .B_N(_2634_),
    .Y(_2636_));
 sg13g2_inv_1 _6553_ (.Y(_2637_),
    .A(_2636_));
 sg13g2_nor2_1 _6554_ (.A(_0710_),
    .B(_2637_),
    .Y(_2638_));
 sg13g2_nor2_1 _6555_ (.A(_1858_),
    .B(_2225_),
    .Y(_2639_));
 sg13g2_nand3_1 _6556_ (.B(net849),
    .C(_2235_),
    .A(_2161_),
    .Y(_2640_));
 sg13g2_a21oi_1 _6557_ (.A1(_2205_),
    .A2(_2640_),
    .Y(_2641_),
    .B1(_1921_));
 sg13g2_or2_1 _6558_ (.X(_2642_),
    .B(_2641_),
    .A(_2639_));
 sg13g2_a22oi_1 _6559_ (.Y(_2643_),
    .B1(_2638_),
    .B2(_2642_),
    .A2(_2637_),
    .A1(net1411));
 sg13g2_nor2_1 _6560_ (.A(net967),
    .B(_2643_),
    .Y(_0555_));
 sg13g2_nand2_1 _6561_ (.Y(_2644_),
    .A(net1333),
    .B(_2637_));
 sg13g2_o21ai_1 _6562_ (.B1(_2225_),
    .Y(_2645_),
    .A1(_2214_),
    .A2(_2222_));
 sg13g2_nand2b_1 _6563_ (.Y(_2646_),
    .B(_1807_),
    .A_N(_2199_));
 sg13g2_nand2b_1 _6564_ (.Y(_2647_),
    .B(_2192_),
    .A_N(_1879_));
 sg13g2_nand3_1 _6565_ (.B(_2646_),
    .C(_2647_),
    .A(_2184_),
    .Y(_2648_));
 sg13g2_nand4_1 _6566_ (.B(_2205_),
    .C(_2640_),
    .A(_1825_),
    .Y(_2649_),
    .D(_2648_));
 sg13g2_nand3_1 _6567_ (.B(_2645_),
    .C(_2649_),
    .A(_1820_),
    .Y(_2650_));
 sg13g2_a21o_1 _6568_ (.A2(_2650_),
    .A1(_2230_),
    .B1(_1843_),
    .X(_2651_));
 sg13g2_nand3_1 _6569_ (.B(_2638_),
    .C(_2651_),
    .A(_2238_),
    .Y(_2652_));
 sg13g2_a21oi_1 _6570_ (.A1(net1334),
    .A2(_2652_),
    .Y(_0556_),
    .B1(net967));
 sg13g2_nor2_1 _6571_ (.A(_0016_),
    .B(_1755_),
    .Y(_2653_));
 sg13g2_nor2_1 _6572_ (.A(net1414),
    .B(_2653_),
    .Y(_2654_));
 sg13g2_nor2_1 _6573_ (.A(net967),
    .B(net1415),
    .Y(_0557_));
 sg13g2_nor2_1 _6574_ (.A(net1014),
    .B(_1755_),
    .Y(_2655_));
 sg13g2_nor2_1 _6575_ (.A(net1309),
    .B(_2655_),
    .Y(_2656_));
 sg13g2_nor2_1 _6576_ (.A(net966),
    .B(_2656_),
    .Y(_0558_));
 sg13g2_nor2_1 _6577_ (.A(net969),
    .B(net1666),
    .Y(_0559_));
 sg13g2_nor2_1 _6578_ (.A(net969),
    .B(net1749),
    .Y(_0560_));
 sg13g2_and2_1 _6579_ (.A(net974),
    .B(_1895_),
    .X(_0561_));
 sg13g2_nor2_1 _6580_ (.A(net966),
    .B(_1888_),
    .Y(_0562_));
 sg13g2_and2_1 _6581_ (.A(net974),
    .B(net1746),
    .X(_0563_));
 sg13g2_nor2_1 _6582_ (.A(net966),
    .B(_1926_),
    .Y(_0564_));
 sg13g2_and2_1 _6583_ (.A(net970),
    .B(_1857_),
    .X(_0565_));
 sg13g2_a21oi_1 _6584_ (.A1(_1828_),
    .A2(net1727),
    .Y(_0566_),
    .B1(net967));
 sg13g2_and2_1 _6585_ (.A(net970),
    .B(_1869_),
    .X(_0567_));
 sg13g2_and2_1 _6586_ (.A(net970),
    .B(_1842_),
    .X(_0568_));
 sg13g2_nor2_1 _6587_ (.A(net966),
    .B(net1701),
    .Y(_0569_));
 sg13g2_and2_1 _6588_ (.A(net970),
    .B(_1878_),
    .X(_0570_));
 sg13g2_nor2_1 _6589_ (.A(\C1.next_state_var[1] ),
    .B(net993),
    .Y(_2657_));
 sg13g2_a221oi_1 _6590_ (.B2(\C1.next_state_var[2] ),
    .C1(_1226_),
    .B1(_1266_),
    .A1(net993),
    .Y(_2658_),
    .A2(_1218_));
 sg13g2_a21oi_1 _6591_ (.A1(_0087_),
    .A2(_2657_),
    .Y(_2659_),
    .B1(_2658_));
 sg13g2_nor2_1 _6592_ (.A(\C1.next_state_var[4] ),
    .B(\C1.next_state_var[2] ),
    .Y(_2660_));
 sg13g2_a21oi_1 _6593_ (.A1(_2657_),
    .A2(_2660_),
    .Y(_2661_),
    .B1(net1001));
 sg13g2_nand4_1 _6594_ (.B(_0674_),
    .C(_0087_),
    .A(_0673_),
    .Y(_2662_),
    .D(_2657_));
 sg13g2_nand3_1 _6595_ (.B(_2661_),
    .C(_2662_),
    .A(_1189_),
    .Y(_2663_));
 sg13g2_nor2_1 _6596_ (.A(net1379),
    .B(_2661_),
    .Y(_2664_));
 sg13g2_o21ai_1 _6597_ (.B1(net971),
    .Y(_2665_),
    .A1(_2659_),
    .A2(_2663_));
 sg13g2_nor2_1 _6598_ (.A(_2664_),
    .B(_2665_),
    .Y(_0571_));
 sg13g2_o21ai_1 _6599_ (.B1(net997),
    .Y(_2666_),
    .A1(net995),
    .A2(\C1.next_state_var[4] ));
 sg13g2_o21ai_1 _6600_ (.B1(net971),
    .Y(_2667_),
    .A1(_0015_),
    .A2(_2666_));
 sg13g2_a21oi_1 _6601_ (.A1(_0680_),
    .A2(_2666_),
    .Y(_0572_),
    .B1(_2667_));
 sg13g2_o21ai_1 _6602_ (.B1(net997),
    .Y(_2668_),
    .A1(\C1.next_state_var[3] ),
    .A2(net993));
 sg13g2_o21ai_1 _6603_ (.B1(net973),
    .Y(_2669_),
    .A1(_0016_),
    .A2(_2668_));
 sg13g2_a21oi_1 _6604_ (.A1(_0679_),
    .A2(_2668_),
    .Y(_0573_),
    .B1(_2669_));
 sg13g2_o21ai_1 _6605_ (.B1(net997),
    .Y(_2670_),
    .A1(\C1.next_state_var[3] ),
    .A2(\C1.next_state_var[2] ));
 sg13g2_o21ai_1 _6606_ (.B1(net973),
    .Y(_2671_),
    .A1(_0016_),
    .A2(_2670_));
 sg13g2_a21oi_1 _6607_ (.A1(_0678_),
    .A2(_2670_),
    .Y(_0574_),
    .B1(_2671_));
 sg13g2_nand2_2 _6608_ (.Y(_2672_),
    .A(net997),
    .B(_1260_));
 sg13g2_a21oi_2 _6609_ (.B1(_2672_),
    .Y(_2673_),
    .A2(_0724_),
    .A1(_0709_));
 sg13g2_o21ai_1 _6610_ (.B1(net971),
    .Y(_2674_),
    .A1(net1569),
    .A2(_2673_));
 sg13g2_a21oi_1 _6611_ (.A1(_0677_),
    .A2(_2673_),
    .Y(_0575_),
    .B1(_2674_));
 sg13g2_nand2b_2 _6612_ (.Y(_2675_),
    .B(_2673_),
    .A_N(_1268_));
 sg13g2_a21oi_2 _6613_ (.B1(_0677_),
    .Y(_2676_),
    .A2(net4),
    .A1(_0723_));
 sg13g2_o21ai_1 _6614_ (.B1(net971),
    .Y(_2677_),
    .A1(_2675_),
    .A2(_2676_));
 sg13g2_a21oi_1 _6615_ (.A1(_0676_),
    .A2(_2675_),
    .Y(_0576_),
    .B1(_2677_));
 sg13g2_nor2_2 _6616_ (.A(net992),
    .B(net3),
    .Y(_2678_));
 sg13g2_o21ai_1 _6617_ (.B1(net971),
    .Y(_2679_),
    .A1(_2675_),
    .A2(_2678_));
 sg13g2_a21oi_1 _6618_ (.A1(_0675_),
    .A2(_2675_),
    .Y(_0577_),
    .B1(_2679_));
 sg13g2_o21ai_1 _6619_ (.B1(_1194_),
    .Y(_2680_),
    .A1(_0709_),
    .A2(\C1.next_state_var[4] ));
 sg13g2_nand2b_1 _6620_ (.Y(_2681_),
    .B(_2680_),
    .A_N(_2672_));
 sg13g2_o21ai_1 _6621_ (.B1(net972),
    .Y(_2682_),
    .A1(_2676_),
    .A2(_2681_));
 sg13g2_a21oi_1 _6622_ (.A1(_0674_),
    .A2(_2681_),
    .Y(_0578_),
    .B1(_2682_));
 sg13g2_o21ai_1 _6623_ (.B1(net972),
    .Y(_2683_),
    .A1(_2678_),
    .A2(_2681_));
 sg13g2_a21oi_1 _6624_ (.A1(_0673_),
    .A2(_2681_),
    .Y(_0579_),
    .B1(_2683_));
 sg13g2_a21oi_1 _6625_ (.A1(\C1.next_state_var[2] ),
    .A2(_1189_),
    .Y(_2684_),
    .B1(_2672_));
 sg13g2_o21ai_1 _6626_ (.B1(_2684_),
    .Y(_2685_),
    .A1(net992),
    .A2(\C1.next_state_var[2] ));
 sg13g2_o21ai_1 _6627_ (.B1(net972),
    .Y(_2686_),
    .A1(_2676_),
    .A2(_2685_));
 sg13g2_a21oi_1 _6628_ (.A1(_0672_),
    .A2(_2685_),
    .Y(_0580_),
    .B1(_2686_));
 sg13g2_o21ai_1 _6629_ (.B1(net972),
    .Y(_2687_),
    .A1(_2678_),
    .A2(_2685_));
 sg13g2_a21oi_1 _6630_ (.A1(_0671_),
    .A2(_2685_),
    .Y(_0581_),
    .B1(_2687_));
 sg13g2_a21oi_1 _6631_ (.A1(net993),
    .A2(_1189_),
    .Y(_2688_),
    .B1(_2672_));
 sg13g2_o21ai_1 _6632_ (.B1(_2688_),
    .Y(_2689_),
    .A1(net992),
    .A2(net993));
 sg13g2_o21ai_1 _6633_ (.B1(net971),
    .Y(_2690_),
    .A1(_2676_),
    .A2(_2689_));
 sg13g2_a21oi_1 _6634_ (.A1(_0670_),
    .A2(_2689_),
    .Y(_0582_),
    .B1(_2690_));
 sg13g2_o21ai_1 _6635_ (.B1(net971),
    .Y(_2691_),
    .A1(_2678_),
    .A2(_2689_));
 sg13g2_a21oi_1 _6636_ (.A1(_0669_),
    .A2(_2689_),
    .Y(_0583_),
    .B1(_2691_));
 sg13g2_nor4_1 _6637_ (.A(\uart_rx_1.r_Clock_Count[27] ),
    .B(\uart_rx_1.r_Clock_Count[26] ),
    .C(\uart_rx_1.r_Clock_Count[25] ),
    .D(\uart_rx_1.r_Clock_Count[24] ),
    .Y(_2692_));
 sg13g2_nor4_1 _6638_ (.A(\uart_rx_1.r_Clock_Count[31] ),
    .B(\uart_rx_1.r_Clock_Count[30] ),
    .C(\uart_rx_1.r_Clock_Count[29] ),
    .D(\uart_rx_1.r_Clock_Count[28] ),
    .Y(_2693_));
 sg13g2_nand2_1 _6639_ (.Y(_2694_),
    .A(_2692_),
    .B(_2693_));
 sg13g2_nor4_1 _6640_ (.A(\uart_rx_1.r_Clock_Count[19] ),
    .B(\uart_rx_1.r_Clock_Count[18] ),
    .C(\uart_rx_1.r_Clock_Count[17] ),
    .D(\uart_rx_1.r_Clock_Count[16] ),
    .Y(_2695_));
 sg13g2_nor4_1 _6641_ (.A(\uart_rx_1.r_Clock_Count[23] ),
    .B(\uart_rx_1.r_Clock_Count[22] ),
    .C(\uart_rx_1.r_Clock_Count[21] ),
    .D(\uart_rx_1.r_Clock_Count[20] ),
    .Y(_2696_));
 sg13g2_nor4_1 _6642_ (.A(\uart_rx_1.r_Clock_Count[11] ),
    .B(\uart_rx_1.r_Clock_Count[10] ),
    .C(\uart_rx_1.r_Clock_Count[9] ),
    .D(\uart_rx_1.r_Clock_Count[8] ),
    .Y(_2697_));
 sg13g2_nor4_1 _6643_ (.A(\uart_rx_1.r_Clock_Count[15] ),
    .B(\uart_rx_1.r_Clock_Count[14] ),
    .C(\uart_rx_1.r_Clock_Count[13] ),
    .D(\uart_rx_1.r_Clock_Count[12] ),
    .Y(_2698_));
 sg13g2_nand4_1 _6644_ (.B(_2696_),
    .C(_2697_),
    .A(_2695_),
    .Y(_2699_),
    .D(_2698_));
 sg13g2_nor2_1 _6645_ (.A(_2694_),
    .B(_2699_),
    .Y(_2700_));
 sg13g2_nor2b_1 _6646_ (.A(\uart_rx_1.r_Clock_Count[4] ),
    .B_N(\uart_rx_1.r_Clock_Count[5] ),
    .Y(_2701_));
 sg13g2_nor2_1 _6647_ (.A(\uart_rx_1.r_Clock_Count[1] ),
    .B(\uart_rx_1.r_Clock_Count[0] ),
    .Y(_2702_));
 sg13g2_nand2_1 _6648_ (.Y(_2703_),
    .A(_2701_),
    .B(_2702_));
 sg13g2_nand2_1 _6649_ (.Y(_2704_),
    .A(\uart_rx_1.r_Clock_Count[3] ),
    .B(\uart_rx_1.r_Clock_Count[2] ));
 sg13g2_a22oi_1 _6650_ (.Y(_2705_),
    .B1(_2704_),
    .B2(_2701_),
    .A2(_2703_),
    .A1(_0100_));
 sg13g2_o21ai_1 _6651_ (.B1(\uart_rx_1.r_Clock_Count[7] ),
    .Y(_2706_),
    .A1(\uart_rx_1.r_Clock_Count[6] ),
    .A2(_2705_));
 sg13g2_nand2_1 _6652_ (.Y(_2707_),
    .A(_2700_),
    .B(_2706_));
 sg13g2_nand2_1 _6653_ (.Y(_2708_),
    .A(\uart_rx_1.r_SM_Main[1] ),
    .B(_0099_));
 sg13g2_nand4_1 _6654_ (.B(net1637),
    .C(_0099_),
    .A(\uart_rx_1.r_SM_Main[1] ),
    .Y(_2709_),
    .D(_2707_));
 sg13g2_nor2_1 _6655_ (.A(\uart_rx_1.r_SM_Main[1] ),
    .B(net1637),
    .Y(_2710_));
 sg13g2_or2_1 _6656_ (.X(_2711_),
    .B(_0099_),
    .A(net1408));
 sg13g2_a221oi_1 _6657_ (.B2(_2711_),
    .C1(net948),
    .B1(_2710_),
    .A1(_0668_),
    .Y(_0584_),
    .A2(_2709_));
 sg13g2_or2_1 _6658_ (.X(_2712_),
    .B(\uart_rx_1.r_Bit_Index[0] ),
    .A(\uart_rx_1.r_Bit_Index[1] ));
 sg13g2_or2_1 _6659_ (.X(_2713_),
    .B(_2712_),
    .A(\uart_rx_1.r_Bit_Index[2] ));
 sg13g2_nor3_2 _6660_ (.A(\uart_rx_1.r_Bit_Index[4] ),
    .B(\uart_rx_1.r_Bit_Index[3] ),
    .C(_2713_),
    .Y(_2714_));
 sg13g2_o21ai_1 _6661_ (.B1(\uart_rx_1.r_Bit_Index[4] ),
    .Y(_2715_),
    .A1(\uart_rx_1.r_Bit_Index[3] ),
    .A2(_2713_));
 sg13g2_nand2b_1 _6662_ (.Y(_2716_),
    .B(_2715_),
    .A_N(_2714_));
 sg13g2_nand2b_1 _6663_ (.Y(_2717_),
    .B(\uart_rx_1.r_Bit_Index[5] ),
    .A_N(_2714_));
 sg13g2_or4_1 _6664_ (.A(\uart_rx_1.r_Bit_Index[9] ),
    .B(\uart_rx_1.r_Bit_Index[8] ),
    .C(\uart_rx_1.r_Bit_Index[7] ),
    .D(\uart_rx_1.r_Bit_Index[6] ),
    .X(_2718_));
 sg13g2_nor3_1 _6665_ (.A(\uart_rx_1.r_Bit_Index[11] ),
    .B(\uart_rx_1.r_Bit_Index[10] ),
    .C(_2718_),
    .Y(_2719_));
 sg13g2_nor4_1 _6666_ (.A(\uart_rx_1.r_Bit_Index[23] ),
    .B(\uart_rx_1.r_Bit_Index[22] ),
    .C(\uart_rx_1.r_Bit_Index[21] ),
    .D(\uart_rx_1.r_Bit_Index[20] ),
    .Y(_2720_));
 sg13g2_nor2_1 _6667_ (.A(\uart_rx_1.r_Bit_Index[19] ),
    .B(\uart_rx_1.r_Bit_Index[18] ),
    .Y(_2721_));
 sg13g2_or4_1 _6668_ (.A(\uart_rx_1.r_Bit_Index[28] ),
    .B(\uart_rx_1.r_Bit_Index[27] ),
    .C(\uart_rx_1.r_Bit_Index[17] ),
    .D(\uart_rx_1.r_Bit_Index[16] ),
    .X(_2722_));
 sg13g2_nand3_1 _6669_ (.B(_2720_),
    .C(_2721_),
    .A(_2719_),
    .Y(_2723_));
 sg13g2_nor4_2 _6670_ (.A(\uart_rx_1.r_Bit_Index[15] ),
    .B(\uart_rx_1.r_Bit_Index[12] ),
    .C(_2722_),
    .Y(_2724_),
    .D(_2723_));
 sg13g2_nor3_2 _6671_ (.A(\uart_rx_1.r_Bit_Index[26] ),
    .B(\uart_rx_1.r_Bit_Index[25] ),
    .C(\uart_rx_1.r_Bit_Index[24] ),
    .Y(_2725_));
 sg13g2_nand2b_1 _6672_ (.Y(_2726_),
    .B(_2725_),
    .A_N(\uart_rx_1.r_Bit_Index[14] ));
 sg13g2_a21oi_1 _6673_ (.A1(_0663_),
    .A2(_2714_),
    .Y(_2727_),
    .B1(_2726_));
 sg13g2_nor2_1 _6674_ (.A(\uart_rx_1.r_SM_Main[0] ),
    .B(_2708_),
    .Y(_2728_));
 sg13g2_and2_1 _6675_ (.A(_2707_),
    .B(_2728_),
    .X(_2729_));
 sg13g2_or3_1 _6676_ (.A(\uart_rx_1.r_Bit_Index[31] ),
    .B(\uart_rx_1.r_Bit_Index[30] ),
    .C(\uart_rx_1.r_Bit_Index[29] ),
    .X(_2730_));
 sg13g2_nor4_1 _6677_ (.A(\uart_rx_1.r_Bit_Index[30] ),
    .B(\uart_rx_1.r_Bit_Index[29] ),
    .C(\uart_rx_1.r_Bit_Index[14] ),
    .D(\uart_rx_1.r_Bit_Index[13] ),
    .Y(_2731_));
 sg13g2_nand3_1 _6678_ (.B(_2725_),
    .C(_2731_),
    .A(_0661_),
    .Y(_2732_));
 sg13g2_nor4_1 _6679_ (.A(\uart_rx_1.r_Bit_Index[5] ),
    .B(\uart_rx_1.r_Bit_Index[4] ),
    .C(\uart_rx_1.r_Bit_Index[3] ),
    .D(_2732_),
    .Y(_2733_));
 sg13g2_and2_1 _6680_ (.A(_2724_),
    .B(_2733_),
    .X(_2734_));
 sg13g2_and3_1 _6681_ (.X(_2735_),
    .A(_2714_),
    .B(_2729_),
    .C(_2734_));
 sg13g2_nand4_1 _6682_ (.B(_2714_),
    .C(_2729_),
    .A(net982),
    .Y(_2736_),
    .D(_2734_));
 sg13g2_o21ai_1 _6683_ (.B1(_2736_),
    .Y(_2737_),
    .A1(net1674),
    .A2(_2735_));
 sg13g2_nor2_1 _6684_ (.A(net950),
    .B(_2737_),
    .Y(_0585_));
 sg13g2_a21oi_1 _6685_ (.A1(\uart_rx_1.r_Bit_Index[2] ),
    .A2(_2712_),
    .Y(_2738_),
    .B1(\uart_rx_1.r_Bit_Index[3] ));
 sg13g2_nand3_1 _6686_ (.B(_2729_),
    .C(_2738_),
    .A(_2713_),
    .Y(_2739_));
 sg13g2_nand2_1 _6687_ (.Y(_2740_),
    .A(\uart_rx_1.r_Bit_Index[1] ),
    .B(\uart_rx_1.r_Bit_Index[0] ));
 sg13g2_and2_1 _6688_ (.A(_2712_),
    .B(_2740_),
    .X(_2741_));
 sg13g2_nand4_1 _6689_ (.B(\uart_rx_1.r_Bit_Index[30] ),
    .C(\uart_rx_1.r_Bit_Index[29] ),
    .A(\uart_rx_1.r_Bit_Index[31] ),
    .Y(_2742_),
    .D(\uart_rx_1.r_Bit_Index[28] ));
 sg13g2_a221oi_1 _6690_ (.B2(_2742_),
    .C1(_2716_),
    .B1(_2730_),
    .A1(\uart_rx_1.r_Bit_Index[13] ),
    .Y(_2743_),
    .A2(_0662_));
 sg13g2_nand4_1 _6691_ (.B(_2724_),
    .C(_2727_),
    .A(_2717_),
    .Y(_2744_),
    .D(_2743_));
 sg13g2_nor2_1 _6692_ (.A(_0205_),
    .B(_2744_),
    .Y(_2745_));
 sg13g2_nand2_1 _6693_ (.Y(_2746_),
    .A(_2741_),
    .B(_2745_));
 sg13g2_nor2_1 _6694_ (.A(_2739_),
    .B(_2746_),
    .Y(_2747_));
 sg13g2_a21oi_1 _6695_ (.A1(net982),
    .A2(_2747_),
    .Y(_2748_),
    .B1(net950));
 sg13g2_o21ai_1 _6696_ (.B1(_2748_),
    .Y(_2749_),
    .A1(net1698),
    .A2(_2747_));
 sg13g2_inv_1 _6697_ (.Y(_0586_),
    .A(net1699));
 sg13g2_nor3_1 _6698_ (.A(_0664_),
    .B(\uart_rx_1.r_Bit_Index[0] ),
    .C(_2744_),
    .Y(_2750_));
 sg13g2_nor2b_1 _6699_ (.A(_2739_),
    .B_N(_2750_),
    .Y(_2751_));
 sg13g2_o21ai_1 _6700_ (.B1(net955),
    .Y(_2752_),
    .A1(net1667),
    .A2(_2751_));
 sg13g2_a21oi_1 _6701_ (.A1(net982),
    .A2(_2751_),
    .Y(_0587_),
    .B1(_2752_));
 sg13g2_nand2b_1 _6702_ (.Y(_2753_),
    .B(_2745_),
    .A_N(_2741_));
 sg13g2_o21ai_1 _6703_ (.B1(net1628),
    .Y(_2754_),
    .A1(_2739_),
    .A2(_2753_));
 sg13g2_nor2_1 _6704_ (.A(net982),
    .B(_2753_),
    .Y(_2755_));
 sg13g2_nand2b_1 _6705_ (.Y(_2756_),
    .B(_2755_),
    .A_N(_2739_));
 sg13g2_a21oi_1 _6706_ (.A1(net1629),
    .A2(_2756_),
    .Y(_0588_),
    .B1(net950));
 sg13g2_nor3_1 _6707_ (.A(_2712_),
    .B(_2739_),
    .C(_2744_),
    .Y(_2757_));
 sg13g2_o21ai_1 _6708_ (.B1(net955),
    .Y(_2758_),
    .A1(net1595),
    .A2(_2757_));
 sg13g2_a21oi_1 _6709_ (.A1(net982),
    .A2(_2757_),
    .Y(_0589_),
    .B1(_2758_));
 sg13g2_a21oi_1 _6710_ (.A1(\uart_rx_1.r_Bit_Index[3] ),
    .A2(_2713_),
    .Y(_2759_),
    .B1(_2738_));
 sg13g2_nand2_1 _6711_ (.Y(_2760_),
    .A(_2729_),
    .B(_2759_));
 sg13g2_inv_1 _6712_ (.Y(_2761_),
    .A(_2760_));
 sg13g2_nor2_1 _6713_ (.A(_2746_),
    .B(_2760_),
    .Y(_2762_));
 sg13g2_o21ai_1 _6714_ (.B1(net953),
    .Y(_2763_),
    .A1(net1515),
    .A2(_2762_));
 sg13g2_a21oi_1 _6715_ (.A1(net982),
    .A2(_2762_),
    .Y(_0590_),
    .B1(net1516));
 sg13g2_a21oi_1 _6716_ (.A1(_2750_),
    .A2(_2761_),
    .Y(_2764_),
    .B1(net1352));
 sg13g2_and3_1 _6717_ (.X(_2765_),
    .A(net982),
    .B(_2750_),
    .C(_2761_));
 sg13g2_nor3_1 _6718_ (.A(net950),
    .B(net1353),
    .C(_2765_),
    .Y(_0591_));
 sg13g2_o21ai_1 _6719_ (.B1(net1419),
    .Y(_2766_),
    .A1(_2753_),
    .A2(_2760_));
 sg13g2_nand2_1 _6720_ (.Y(_2767_),
    .A(_2755_),
    .B(_2761_));
 sg13g2_a21oi_1 _6721_ (.A1(net1420),
    .A2(_2767_),
    .Y(_0592_),
    .B1(net950));
 sg13g2_nand2_1 _6722_ (.Y(_2768_),
    .A(_0099_),
    .B(_2710_));
 sg13g2_nor2b_1 _6723_ (.A(_2729_),
    .B_N(_2768_),
    .Y(_2769_));
 sg13g2_inv_1 _6724_ (.Y(_2770_),
    .A(net886));
 sg13g2_nand4_1 _6725_ (.B(\uart_rx_1.r_Bit_Index[2] ),
    .C(\uart_rx_1.r_Bit_Index[1] ),
    .A(_0661_),
    .Y(_2771_),
    .D(\uart_rx_1.r_Bit_Index[0] ));
 sg13g2_nand3_1 _6726_ (.B(_2734_),
    .C(_2771_),
    .A(_2728_),
    .Y(_2772_));
 sg13g2_nor2_1 _6727_ (.A(net886),
    .B(_2772_),
    .Y(_2773_));
 sg13g2_o21ai_1 _6728_ (.B1(net953),
    .Y(_2774_),
    .A1(net1598),
    .A2(_2773_));
 sg13g2_a21oi_1 _6729_ (.A1(net1598),
    .A2(_2770_),
    .Y(_0593_),
    .B1(_2774_));
 sg13g2_a22oi_1 _6730_ (.Y(_2775_),
    .B1(_2773_),
    .B2(_2741_),
    .A2(net886),
    .A1(net1608));
 sg13g2_nor2_1 _6731_ (.A(net949),
    .B(_2775_),
    .Y(_0594_));
 sg13g2_xor2_1 _6732_ (.B(_2740_),
    .A(net1435),
    .X(_2776_));
 sg13g2_a22oi_1 _6733_ (.Y(_2777_),
    .B1(_2773_),
    .B2(net1436),
    .A2(net886),
    .A1(\uart_rx_1.r_Bit_Index[2] ));
 sg13g2_nor2_1 _6734_ (.A(net948),
    .B(net1437),
    .Y(_0595_));
 sg13g2_and3_1 _6735_ (.X(_0596_),
    .A(net1535),
    .B(net953),
    .C(net886));
 sg13g2_and3_1 _6736_ (.X(_0597_),
    .A(net1418),
    .B(net954),
    .C(net886));
 sg13g2_nor3_1 _6737_ (.A(_0663_),
    .B(net948),
    .C(_2770_),
    .Y(_0598_));
 sg13g2_and3_1 _6738_ (.X(_0599_),
    .A(net731),
    .B(net958),
    .C(net887));
 sg13g2_and3_1 _6739_ (.X(_0600_),
    .A(net732),
    .B(net958),
    .C(net887));
 sg13g2_and3_1 _6740_ (.X(_0601_),
    .A(net756),
    .B(net958),
    .C(net887));
 sg13g2_and3_1 _6741_ (.X(_0602_),
    .A(net741),
    .B(net958),
    .C(net887));
 sg13g2_and3_1 _6742_ (.X(_0603_),
    .A(net733),
    .B(net959),
    .C(net887));
 sg13g2_and3_1 _6743_ (.X(_0604_),
    .A(net752),
    .B(net959),
    .C(net887));
 sg13g2_nor3_1 _6744_ (.A(_0662_),
    .B(net951),
    .C(_2770_),
    .Y(_0605_));
 sg13g2_and3_1 _6745_ (.X(_0606_),
    .A(net1017),
    .B(net954),
    .C(net890));
 sg13g2_and3_1 _6746_ (.X(_0607_),
    .A(net1054),
    .B(net954),
    .C(net890));
 sg13g2_and3_1 _6747_ (.X(_0608_),
    .A(net1012),
    .B(net956),
    .C(net889));
 sg13g2_and3_1 _6748_ (.X(_0609_),
    .A(net755),
    .B(net958),
    .C(net889));
 sg13g2_and3_1 _6749_ (.X(_0610_),
    .A(net747),
    .B(net956),
    .C(net889));
 sg13g2_and3_1 _6750_ (.X(_0611_),
    .A(net734),
    .B(net959),
    .C(net888));
 sg13g2_and3_1 _6751_ (.X(_0612_),
    .A(net1005),
    .B(net959),
    .C(net888));
 sg13g2_and3_1 _6752_ (.X(_0613_),
    .A(net1003),
    .B(net959),
    .C(net888));
 sg13g2_and3_1 _6753_ (.X(_0614_),
    .A(net1007),
    .B(net959),
    .C(net887));
 sg13g2_and3_1 _6754_ (.X(_0615_),
    .A(net738),
    .B(net958),
    .C(net887));
 sg13g2_and3_1 _6755_ (.X(_0616_),
    .A(net743),
    .B(net958),
    .C(net888));
 sg13g2_and3_1 _6756_ (.X(_0617_),
    .A(net1011),
    .B(net956),
    .C(net889));
 sg13g2_and3_1 _6757_ (.X(_0618_),
    .A(net1028),
    .B(net956),
    .C(net889));
 sg13g2_and3_1 _6758_ (.X(_0619_),
    .A(net1016),
    .B(net956),
    .C(net889));
 sg13g2_and3_1 _6759_ (.X(_0620_),
    .A(net748),
    .B(net958),
    .C(net889));
 sg13g2_and3_1 _6760_ (.X(_0621_),
    .A(net1330),
    .B(net956),
    .C(net889));
 sg13g2_and3_1 _6761_ (.X(_0622_),
    .A(net1277),
    .B(net954),
    .C(net886));
 sg13g2_and3_1 _6762_ (.X(_0623_),
    .A(net1178),
    .B(net954),
    .C(net886));
 sg13g2_nor3_1 _6763_ (.A(_0661_),
    .B(net948),
    .C(_2770_),
    .Y(_0624_));
 sg13g2_nor2b_1 _6764_ (.A(\uart_rx_1.r_SM_Main[1] ),
    .B_N(\uart_rx_1.r_SM_Main[0] ),
    .Y(_2778_));
 sg13g2_nand2b_1 _6765_ (.Y(_2779_),
    .B(\uart_rx_1.r_SM_Main[0] ),
    .A_N(\uart_rx_1.r_SM_Main[1] ));
 sg13g2_nand2_1 _6766_ (.Y(_2780_),
    .A(_0099_),
    .B(_2779_));
 sg13g2_nand2b_1 _6767_ (.Y(_2781_),
    .B(\uart_rx_1.r_Clock_Count[4] ),
    .A_N(\uart_rx_1.r_Clock_Count[5] ));
 sg13g2_nand4_1 _6768_ (.B(\uart_rx_1.r_Clock_Count[6] ),
    .C(\uart_rx_1.r_Clock_Count[2] ),
    .A(_0660_),
    .Y(_2782_),
    .D(\uart_rx_1.r_Clock_Count[1] ));
 sg13g2_nor4_1 _6769_ (.A(\uart_rx_1.r_Clock_Count[3] ),
    .B(\uart_rx_1.r_Clock_Count[0] ),
    .C(_2781_),
    .D(_2782_),
    .Y(_2783_));
 sg13g2_and2_1 _6770_ (.A(_2700_),
    .B(_2783_),
    .X(_2784_));
 sg13g2_inv_1 _6771_ (.Y(_2785_),
    .A(_2784_));
 sg13g2_nor2_2 _6772_ (.A(_0101_),
    .B(_2785_),
    .Y(_2786_));
 sg13g2_a21o_1 _6773_ (.A2(_2786_),
    .A1(_2778_),
    .B1(_0727_),
    .X(_2787_));
 sg13g2_o21ai_1 _6774_ (.B1(_2780_),
    .Y(_2788_),
    .A1(_0727_),
    .A2(_2786_));
 sg13g2_and2_1 _6775_ (.A(net1508),
    .B(net883),
    .X(_2789_));
 sg13g2_nor2_1 _6776_ (.A(_2707_),
    .B(_2708_),
    .Y(_2790_));
 sg13g2_nor2_2 _6777_ (.A(_0727_),
    .B(_2779_),
    .Y(_2791_));
 sg13g2_nand2_2 _6778_ (.Y(_2792_),
    .A(_0099_),
    .B(_2778_));
 sg13g2_a21oi_2 _6779_ (.B1(_2790_),
    .Y(_2793_),
    .A2(net935),
    .A1(_2785_));
 sg13g2_nor2b_1 _6780_ (.A(net1508),
    .B_N(_2793_),
    .Y(_2794_));
 sg13g2_nor3_1 _6781_ (.A(net948),
    .B(_2789_),
    .C(_2794_),
    .Y(_0625_));
 sg13g2_a21o_2 _6782_ (.A2(_2793_),
    .A1(net883),
    .B1(net948),
    .X(_2795_));
 sg13g2_xnor2_1 _6783_ (.Y(_2796_),
    .A(net1661),
    .B(_2789_));
 sg13g2_nor2_1 _6784_ (.A(_2795_),
    .B(_2796_),
    .Y(_0626_));
 sg13g2_a21oi_1 _6785_ (.A1(\uart_rx_1.r_Clock_Count[1] ),
    .A2(_2789_),
    .Y(_2797_),
    .B1(net1356));
 sg13g2_and3_1 _6786_ (.X(_2798_),
    .A(net1356),
    .B(\uart_rx_1.r_Clock_Count[1] ),
    .C(_2789_));
 sg13g2_nor3_1 _6787_ (.A(_2795_),
    .B(net1357),
    .C(_2798_),
    .Y(_0627_));
 sg13g2_o21ai_1 _6788_ (.B1(net954),
    .Y(_2799_),
    .A1(_2780_),
    .A2(_2790_));
 sg13g2_xnor2_1 _6789_ (.Y(_2800_),
    .A(net1582),
    .B(_2798_));
 sg13g2_nor2_1 _6790_ (.A(_2799_),
    .B(net1583),
    .Y(_0628_));
 sg13g2_a21oi_1 _6791_ (.A1(\uart_rx_1.r_Clock_Count[3] ),
    .A2(_2798_),
    .Y(_2801_),
    .B1(net1429));
 sg13g2_nand3_1 _6792_ (.B(\uart_rx_1.r_Clock_Count[1] ),
    .C(\uart_rx_1.r_Clock_Count[0] ),
    .A(\uart_rx_1.r_Clock_Count[4] ),
    .Y(_2802_));
 sg13g2_or2_1 _6793_ (.X(_2803_),
    .B(_2802_),
    .A(_2704_));
 sg13g2_nor2_1 _6794_ (.A(net884),
    .B(_2803_),
    .Y(_2804_));
 sg13g2_nor3_1 _6795_ (.A(_2795_),
    .B(net1430),
    .C(_2804_),
    .Y(_0629_));
 sg13g2_xor2_1 _6796_ (.B(_2803_),
    .A(_0100_),
    .X(_2805_));
 sg13g2_nor2_1 _6797_ (.A(net884),
    .B(_2805_),
    .Y(_2806_));
 sg13g2_nor2_1 _6798_ (.A(net1622),
    .B(net883),
    .Y(_2807_));
 sg13g2_nor3_1 _6799_ (.A(_2795_),
    .B(_2806_),
    .C(_2807_),
    .Y(_0630_));
 sg13g2_a21oi_1 _6800_ (.A1(\uart_rx_1.r_Clock_Count[5] ),
    .A2(_2804_),
    .Y(_2808_),
    .B1(net1505));
 sg13g2_and3_1 _6801_ (.X(_2809_),
    .A(net1505),
    .B(\uart_rx_1.r_Clock_Count[5] ),
    .C(_2804_));
 sg13g2_nor3_1 _6802_ (.A(_2795_),
    .B(net1506),
    .C(_2809_),
    .Y(_0631_));
 sg13g2_xnor2_1 _6803_ (.Y(_2810_),
    .A(net1619),
    .B(_2809_));
 sg13g2_nor2_1 _6804_ (.A(_2799_),
    .B(net1620),
    .Y(_0632_));
 sg13g2_nand4_1 _6805_ (.B(\uart_rx_1.r_Clock_Count[7] ),
    .C(\uart_rx_1.r_Clock_Count[6] ),
    .A(net1173),
    .Y(_2811_),
    .D(\uart_rx_1.r_Clock_Count[5] ));
 sg13g2_nor2_1 _6806_ (.A(_2803_),
    .B(_2811_),
    .Y(_2812_));
 sg13g2_inv_1 _6807_ (.Y(_2813_),
    .A(_2812_));
 sg13g2_a21oi_1 _6808_ (.A1(net935),
    .A2(_2813_),
    .Y(_2814_),
    .B1(net884));
 sg13g2_a21oi_1 _6809_ (.A1(\uart_rx_1.r_Clock_Count[7] ),
    .A2(_2809_),
    .Y(_2815_),
    .B1(net1173));
 sg13g2_nor3_1 _6810_ (.A(net948),
    .B(_2814_),
    .C(net1174),
    .Y(_0633_));
 sg13g2_nand3b_1 _6811_ (.B(net953),
    .C(net1471),
    .Y(_2816_),
    .A_N(_2814_));
 sg13g2_nor2_2 _6812_ (.A(_2786_),
    .B(_2792_),
    .Y(_2817_));
 sg13g2_nand3b_1 _6813_ (.B(_2812_),
    .C(net881),
    .Y(_2818_),
    .A_N(net1471));
 sg13g2_o21ai_1 _6814_ (.B1(_2816_),
    .Y(_0634_),
    .A1(net949),
    .A2(_2818_));
 sg13g2_and2_1 _6815_ (.A(\uart_rx_1.r_Clock_Count[9] ),
    .B(_2812_),
    .X(_2819_));
 sg13g2_a21oi_1 _6816_ (.A1(net883),
    .A2(_2819_),
    .Y(_2820_),
    .B1(net1167));
 sg13g2_and2_1 _6817_ (.A(net1167),
    .B(_2819_),
    .X(_2821_));
 sg13g2_inv_1 _6818_ (.Y(_2822_),
    .A(_2821_));
 sg13g2_a21oi_1 _6819_ (.A1(net935),
    .A2(_2822_),
    .Y(_2823_),
    .B1(net884));
 sg13g2_nor3_1 _6820_ (.A(net949),
    .B(net1168),
    .C(_2823_),
    .Y(_0635_));
 sg13g2_a21oi_1 _6821_ (.A1(net881),
    .A2(_2821_),
    .Y(_2824_),
    .B1(net1655));
 sg13g2_a21oi_1 _6822_ (.A1(net1655),
    .A2(_2823_),
    .Y(_2825_),
    .B1(_2824_));
 sg13g2_and2_1 _6823_ (.A(net953),
    .B(_2825_),
    .X(_0636_));
 sg13g2_and2_1 _6824_ (.A(\uart_rx_1.r_Clock_Count[11] ),
    .B(_2821_),
    .X(_2826_));
 sg13g2_and2_1 _6825_ (.A(\uart_rx_1.r_Clock_Count[12] ),
    .B(_2826_),
    .X(_2827_));
 sg13g2_nor2_1 _6826_ (.A(_2792_),
    .B(_2827_),
    .Y(_2828_));
 sg13g2_nor2_1 _6827_ (.A(net885),
    .B(_2828_),
    .Y(_2829_));
 sg13g2_a21oi_1 _6828_ (.A1(net882),
    .A2(_2826_),
    .Y(_2830_),
    .B1(net1097));
 sg13g2_nor3_1 _6829_ (.A(net951),
    .B(_2829_),
    .C(net1098),
    .Y(_0637_));
 sg13g2_a21oi_1 _6830_ (.A1(net881),
    .A2(_2827_),
    .Y(_2831_),
    .B1(net1080));
 sg13g2_nand2b_1 _6831_ (.Y(_2832_),
    .B(net955),
    .A_N(_2831_));
 sg13g2_a21oi_1 _6832_ (.A1(net1080),
    .A2(_2829_),
    .Y(_0638_),
    .B1(_2832_));
 sg13g2_and2_1 _6833_ (.A(net1080),
    .B(_2827_),
    .X(_2833_));
 sg13g2_and2_1 _6834_ (.A(net1144),
    .B(_2833_),
    .X(_2834_));
 sg13g2_inv_1 _6835_ (.Y(_2835_),
    .A(_2834_));
 sg13g2_a21oi_1 _6836_ (.A1(_2791_),
    .A2(_2835_),
    .Y(_2836_),
    .B1(net885));
 sg13g2_a21oi_1 _6837_ (.A1(net882),
    .A2(_2833_),
    .Y(_2837_),
    .B1(net1144));
 sg13g2_nor3_1 _6838_ (.A(net951),
    .B(_2836_),
    .C(_2837_),
    .Y(_0639_));
 sg13g2_a21oi_1 _6839_ (.A1(_2817_),
    .A2(_2834_),
    .Y(_2838_),
    .B1(net1169));
 sg13g2_nand2b_1 _6840_ (.Y(_2839_),
    .B(net956),
    .A_N(_2838_));
 sg13g2_a21oi_1 _6841_ (.A1(net1169),
    .A2(_2836_),
    .Y(_0640_),
    .B1(_2839_));
 sg13g2_and2_1 _6842_ (.A(\uart_rx_1.r_Clock_Count[15] ),
    .B(_2834_),
    .X(_2840_));
 sg13g2_and2_1 _6843_ (.A(\uart_rx_1.r_Clock_Count[16] ),
    .B(_2840_),
    .X(_2841_));
 sg13g2_inv_1 _6844_ (.Y(_2842_),
    .A(_2841_));
 sg13g2_a21oi_1 _6845_ (.A1(_2791_),
    .A2(_2842_),
    .Y(_2843_),
    .B1(net885));
 sg13g2_a21oi_1 _6846_ (.A1(net882),
    .A2(_2840_),
    .Y(_2844_),
    .B1(net1094));
 sg13g2_nor3_1 _6847_ (.A(net951),
    .B(_2843_),
    .C(net1095),
    .Y(_0641_));
 sg13g2_a21oi_1 _6848_ (.A1(_2817_),
    .A2(_2841_),
    .Y(_2845_),
    .B1(net1302));
 sg13g2_nand2b_1 _6849_ (.Y(_2846_),
    .B(net957),
    .A_N(_2845_));
 sg13g2_a21oi_1 _6850_ (.A1(net1302),
    .A2(_2843_),
    .Y(_0642_),
    .B1(_2846_));
 sg13g2_and3_1 _6851_ (.X(_2847_),
    .A(\uart_rx_1.r_Clock_Count[18] ),
    .B(\uart_rx_1.r_Clock_Count[17] ),
    .C(_2841_));
 sg13g2_nor2_1 _6852_ (.A(_2792_),
    .B(_2847_),
    .Y(_2848_));
 sg13g2_nor2_1 _6853_ (.A(net885),
    .B(_2848_),
    .Y(_2849_));
 sg13g2_nand3_1 _6854_ (.B(net882),
    .C(_2841_),
    .A(net1302),
    .Y(_2850_));
 sg13g2_nor2b_1 _6855_ (.A(net1351),
    .B_N(_2850_),
    .Y(_2851_));
 sg13g2_nor3_1 _6856_ (.A(net951),
    .B(_2849_),
    .C(_2851_),
    .Y(_0643_));
 sg13g2_a21oi_1 _6857_ (.A1(net881),
    .A2(_2847_),
    .Y(_2852_),
    .B1(net1120));
 sg13g2_nand2b_1 _6858_ (.Y(_2853_),
    .B(net957),
    .A_N(_2852_));
 sg13g2_a21oi_1 _6859_ (.A1(net1120),
    .A2(_2849_),
    .Y(_0644_),
    .B1(_2853_));
 sg13g2_and2_1 _6860_ (.A(\uart_rx_1.r_Clock_Count[19] ),
    .B(_2847_),
    .X(_2854_));
 sg13g2_and2_1 _6861_ (.A(\uart_rx_1.r_Clock_Count[20] ),
    .B(_2854_),
    .X(_2855_));
 sg13g2_inv_1 _6862_ (.Y(_2856_),
    .A(_2855_));
 sg13g2_a21oi_1 _6863_ (.A1(net935),
    .A2(_2856_),
    .Y(_2857_),
    .B1(net885));
 sg13g2_a21oi_1 _6864_ (.A1(net883),
    .A2(_2854_),
    .Y(_2858_),
    .B1(net1082));
 sg13g2_nor3_1 _6865_ (.A(net951),
    .B(_2857_),
    .C(net1083),
    .Y(_0645_));
 sg13g2_a21oi_1 _6866_ (.A1(net881),
    .A2(_2855_),
    .Y(_2859_),
    .B1(net1067));
 sg13g2_nand2b_1 _6867_ (.Y(_2860_),
    .B(net957),
    .A_N(_2859_));
 sg13g2_a21oi_1 _6868_ (.A1(net1067),
    .A2(_2857_),
    .Y(_0646_),
    .B1(_2860_));
 sg13g2_and2_1 _6869_ (.A(net1067),
    .B(_2855_),
    .X(_2861_));
 sg13g2_and2_1 _6870_ (.A(\uart_rx_1.r_Clock_Count[22] ),
    .B(_2861_),
    .X(_2862_));
 sg13g2_inv_1 _6871_ (.Y(_2863_),
    .A(_2862_));
 sg13g2_a21oi_1 _6872_ (.A1(net935),
    .A2(_2863_),
    .Y(_2864_),
    .B1(net884));
 sg13g2_a21oi_1 _6873_ (.A1(net882),
    .A2(_2861_),
    .Y(_2865_),
    .B1(net1139));
 sg13g2_nor3_1 _6874_ (.A(net952),
    .B(_2864_),
    .C(_2865_),
    .Y(_0647_));
 sg13g2_a21oi_1 _6875_ (.A1(net881),
    .A2(_2862_),
    .Y(_2866_),
    .B1(net1487));
 sg13g2_nand2b_1 _6876_ (.Y(_2867_),
    .B(net957),
    .A_N(_2866_));
 sg13g2_a21oi_1 _6877_ (.A1(net1487),
    .A2(_2864_),
    .Y(_0648_),
    .B1(_2867_));
 sg13g2_and3_1 _6878_ (.X(_2868_),
    .A(\uart_rx_1.r_Clock_Count[24] ),
    .B(\uart_rx_1.r_Clock_Count[23] ),
    .C(_2862_));
 sg13g2_nor2_1 _6879_ (.A(_2792_),
    .B(_2868_),
    .Y(_2869_));
 sg13g2_nor2_1 _6880_ (.A(net884),
    .B(_2869_),
    .Y(_2870_));
 sg13g2_nand3_1 _6881_ (.B(net882),
    .C(_2862_),
    .A(\uart_rx_1.r_Clock_Count[23] ),
    .Y(_2871_));
 sg13g2_nor2b_1 _6882_ (.A(net1462),
    .B_N(_2871_),
    .Y(_2872_));
 sg13g2_nor3_1 _6883_ (.A(net951),
    .B(_2870_),
    .C(net1463),
    .Y(_0649_));
 sg13g2_a21oi_1 _6884_ (.A1(net881),
    .A2(_2868_),
    .Y(_2873_),
    .B1(net1156));
 sg13g2_nand2b_1 _6885_ (.Y(_2874_),
    .B(net956),
    .A_N(_2873_));
 sg13g2_a21oi_1 _6886_ (.A1(net1156),
    .A2(_2870_),
    .Y(_0650_),
    .B1(_2874_));
 sg13g2_and2_1 _6887_ (.A(net1156),
    .B(_2868_),
    .X(_2875_));
 sg13g2_and2_1 _6888_ (.A(\uart_rx_1.r_Clock_Count[26] ),
    .B(_2875_),
    .X(_2876_));
 sg13g2_inv_1 _6889_ (.Y(_2877_),
    .A(_2876_));
 sg13g2_a21oi_1 _6890_ (.A1(net935),
    .A2(_2877_),
    .Y(_2878_),
    .B1(net885));
 sg13g2_a21oi_1 _6891_ (.A1(net882),
    .A2(_2875_),
    .Y(_2879_),
    .B1(net1170));
 sg13g2_nor3_1 _6892_ (.A(net951),
    .B(_2878_),
    .C(_2879_),
    .Y(_0651_));
 sg13g2_a21oi_1 _6893_ (.A1(_2817_),
    .A2(_2876_),
    .Y(_2880_),
    .B1(net1142));
 sg13g2_nand2b_1 _6894_ (.Y(_2881_),
    .B(net954),
    .A_N(_2880_));
 sg13g2_a21oi_1 _6895_ (.A1(net1142),
    .A2(_2878_),
    .Y(_0652_),
    .B1(_2881_));
 sg13g2_and2_1 _6896_ (.A(net1142),
    .B(_2876_),
    .X(_2882_));
 sg13g2_and2_1 _6897_ (.A(\uart_rx_1.r_Clock_Count[28] ),
    .B(_2882_),
    .X(_2883_));
 sg13g2_inv_1 _6898_ (.Y(_2884_),
    .A(_2883_));
 sg13g2_a21oi_1 _6899_ (.A1(net935),
    .A2(_2884_),
    .Y(_2885_),
    .B1(net884));
 sg13g2_a21oi_1 _6900_ (.A1(net882),
    .A2(_2882_),
    .Y(_2886_),
    .B1(net1204));
 sg13g2_nor3_1 _6901_ (.A(net949),
    .B(_2885_),
    .C(_2886_),
    .Y(_0653_));
 sg13g2_a21oi_1 _6902_ (.A1(net881),
    .A2(_2883_),
    .Y(_2887_),
    .B1(net1397));
 sg13g2_nand2b_1 _6903_ (.Y(_2888_),
    .B(net955),
    .A_N(_2887_));
 sg13g2_a21oi_1 _6904_ (.A1(net1397),
    .A2(_2885_),
    .Y(_0654_),
    .B1(_2888_));
 sg13g2_nand3_1 _6905_ (.B(\uart_rx_1.r_Clock_Count[29] ),
    .C(_2883_),
    .A(\uart_rx_1.r_Clock_Count[30] ),
    .Y(_2889_));
 sg13g2_a21oi_1 _6906_ (.A1(net935),
    .A2(_2889_),
    .Y(_2890_),
    .B1(net884));
 sg13g2_nand3_1 _6907_ (.B(net883),
    .C(_2883_),
    .A(\uart_rx_1.r_Clock_Count[29] ),
    .Y(_2891_));
 sg13g2_nor2b_1 _6908_ (.A(net1338),
    .B_N(_2891_),
    .Y(_2892_));
 sg13g2_nor3_1 _6909_ (.A(net949),
    .B(_2890_),
    .C(net1339),
    .Y(_0655_));
 sg13g2_nor3_1 _6910_ (.A(_2786_),
    .B(_2792_),
    .C(_2889_),
    .Y(_2893_));
 sg13g2_o21ai_1 _6911_ (.B1(net953),
    .Y(_2894_),
    .A1(net1075),
    .A2(_2893_));
 sg13g2_a21oi_1 _6912_ (.A1(net1075),
    .A2(_2890_),
    .Y(_0656_),
    .B1(_2894_));
 sg13g2_o21ai_1 _6913_ (.B1(_2793_),
    .Y(_2895_),
    .A1(net982),
    .A2(_2768_));
 sg13g2_nor2b_2 _6914_ (.A(_2895_),
    .B_N(_2772_),
    .Y(_2896_));
 sg13g2_o21ai_1 _6915_ (.B1(_2896_),
    .Y(_2897_),
    .A1(net1408),
    .A2(net1637));
 sg13g2_o21ai_1 _6916_ (.B1(net953),
    .Y(_2898_),
    .A1(net1637),
    .A2(_2896_));
 sg13g2_nor2b_1 _6917_ (.A(_2898_),
    .B_N(_2897_),
    .Y(_0657_));
 sg13g2_nor2_1 _6918_ (.A(\uart_rx_1.r_Rx_Data ),
    .B(_2792_),
    .Y(_2899_));
 sg13g2_nor3_1 _6919_ (.A(_2728_),
    .B(_2895_),
    .C(_2899_),
    .Y(_2900_));
 sg13g2_o21ai_1 _6920_ (.B1(net953),
    .Y(_2901_),
    .A1(net1662),
    .A2(_2896_));
 sg13g2_nor2_1 _6921_ (.A(_2900_),
    .B(_2901_),
    .Y(_0658_));
 sg13g2_nand2b_1 _6922_ (.Y(_2902_),
    .B(net1408),
    .A_N(_2896_));
 sg13g2_a21oi_1 _6923_ (.A1(_2709_),
    .A2(_2902_),
    .Y(_0659_),
    .B1(net948));
 sg13g2_dfrbp_1 _6924_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net27),
    .D(_0209_),
    .Q_N(_3203_),
    .Q(\C1.spinning ));
 sg13g2_dfrbp_1 _6925_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net28),
    .D(_0000_),
    .Q_N(_3204_),
    .Q(\C1.counter_status[0] ));
 sg13g2_dfrbp_1 _6926_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net101),
    .D(_0001_),
    .Q_N(_3205_),
    .Q(\C1.counter_status[1] ));
 sg13g2_dfrbp_1 _6927_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net26),
    .D(_0002_),
    .Q_N(_3202_),
    .Q(\C1.counter_status[2] ));
 sg13g2_dfrbp_1 _6928_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net421),
    .D(_0210_),
    .Q_N(_0043_),
    .Q(\instrs[10][0] ));
 sg13g2_dfrbp_1 _6929_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net420),
    .D(_0211_),
    .Q_N(_3201_),
    .Q(\instrs[10][1] ));
 sg13g2_dfrbp_1 _6930_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net419),
    .D(_0212_),
    .Q_N(_3200_),
    .Q(\instrs[10][2] ));
 sg13g2_dfrbp_1 _6931_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net418),
    .D(_0213_),
    .Q_N(_3199_),
    .Q(\instrs[10][3] ));
 sg13g2_dfrbp_1 _6932_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net417),
    .D(net1199),
    .Q_N(_3198_),
    .Q(\instrs[10][4] ));
 sg13g2_dfrbp_1 _6933_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net416),
    .D(_0215_),
    .Q_N(_0063_),
    .Q(\instrs[10][5] ));
 sg13g2_dfrbp_1 _6934_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net415),
    .D(_0216_),
    .Q_N(_3197_),
    .Q(\instrs[10][6] ));
 sg13g2_dfrbp_1 _6935_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net414),
    .D(_0217_),
    .Q_N(_0079_),
    .Q(\instrs[10][7] ));
 sg13g2_dfrbp_1 _6936_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net413),
    .D(_0218_),
    .Q_N(_0120_),
    .Q(\datam[14][0] ));
 sg13g2_dfrbp_1 _6937_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net412),
    .D(_0219_),
    .Q_N(_0138_),
    .Q(\datam[14][1] ));
 sg13g2_dfrbp_1 _6938_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net411),
    .D(_0220_),
    .Q_N(_0154_),
    .Q(\datam[14][2] ));
 sg13g2_dfrbp_1 _6939_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net410),
    .D(_0221_),
    .Q_N(_0170_),
    .Q(\datam[14][3] ));
 sg13g2_dfrbp_1 _6940_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net409),
    .D(_0222_),
    .Q_N(_0187_),
    .Q(\datam[14][4] ));
 sg13g2_dfrbp_1 _6941_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net408),
    .D(_0223_),
    .Q_N(_3196_),
    .Q(\datam[14][5] ));
 sg13g2_dfrbp_1 _6942_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net407),
    .D(_0224_),
    .Q_N(_3195_),
    .Q(\datam[14][6] ));
 sg13g2_dfrbp_1 _6943_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net406),
    .D(_0225_),
    .Q_N(_3194_),
    .Q(\datam[14][7] ));
 sg13g2_dfrbp_1 _6944_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net405),
    .D(_0226_),
    .Q_N(_0033_),
    .Q(\instrs[0][0] ));
 sg13g2_dfrbp_1 _6945_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net404),
    .D(_0227_),
    .Q_N(_3193_),
    .Q(\instrs[0][1] ));
 sg13g2_dfrbp_1 _6946_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net403),
    .D(_0228_),
    .Q_N(_3192_),
    .Q(\instrs[0][2] ));
 sg13g2_dfrbp_1 _6947_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net402),
    .D(_0229_),
    .Q_N(_3191_),
    .Q(\instrs[0][3] ));
 sg13g2_dfrbp_1 _6948_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net401),
    .D(net1223),
    .Q_N(_3190_),
    .Q(\instrs[0][4] ));
 sg13g2_dfrbp_1 _6949_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net400),
    .D(_0231_),
    .Q_N(_0053_),
    .Q(\instrs[0][5] ));
 sg13g2_dfrbp_1 _6950_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net399),
    .D(_0232_),
    .Q_N(_3189_),
    .Q(\instrs[0][6] ));
 sg13g2_dfrbp_1 _6951_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net398),
    .D(_0233_),
    .Q_N(_0069_),
    .Q(\instrs[0][7] ));
 sg13g2_dfrbp_1 _6952_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net397),
    .D(_0234_),
    .Q_N(_0041_),
    .Q(\instrs[8][0] ));
 sg13g2_dfrbp_1 _6953_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net396),
    .D(_0235_),
    .Q_N(_3188_),
    .Q(\instrs[8][1] ));
 sg13g2_dfrbp_1 _6954_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net395),
    .D(_0236_),
    .Q_N(_3187_),
    .Q(\instrs[8][2] ));
 sg13g2_dfrbp_1 _6955_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net394),
    .D(_0237_),
    .Q_N(_3186_),
    .Q(\instrs[8][3] ));
 sg13g2_dfrbp_1 _6956_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net393),
    .D(net1183),
    .Q_N(_3185_),
    .Q(\instrs[8][4] ));
 sg13g2_dfrbp_1 _6957_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net392),
    .D(_0239_),
    .Q_N(_0061_),
    .Q(\instrs[8][5] ));
 sg13g2_dfrbp_1 _6958_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net391),
    .D(_0240_),
    .Q_N(_3184_),
    .Q(\instrs[8][6] ));
 sg13g2_dfrbp_1 _6959_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net390),
    .D(_0241_),
    .Q_N(_0077_),
    .Q(\instrs[8][7] ));
 sg13g2_dfrbp_1 _6960_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net389),
    .D(_0242_),
    .Q_N(_0040_),
    .Q(\instrs[7][0] ));
 sg13g2_dfrbp_1 _6961_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net388),
    .D(_0243_),
    .Q_N(_3183_),
    .Q(\instrs[7][1] ));
 sg13g2_dfrbp_1 _6962_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net387),
    .D(_0244_),
    .Q_N(_3182_),
    .Q(\instrs[7][2] ));
 sg13g2_dfrbp_1 _6963_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net386),
    .D(_0245_),
    .Q_N(_3181_),
    .Q(\instrs[7][3] ));
 sg13g2_dfrbp_1 _6964_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net385),
    .D(net1041),
    .Q_N(_3180_),
    .Q(\instrs[7][4] ));
 sg13g2_dfrbp_1 _6965_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net384),
    .D(_0247_),
    .Q_N(_0060_),
    .Q(\instrs[7][5] ));
 sg13g2_dfrbp_1 _6966_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net383),
    .D(_0248_),
    .Q_N(_3179_),
    .Q(\instrs[7][6] ));
 sg13g2_dfrbp_1 _6967_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net382),
    .D(_0249_),
    .Q_N(_0076_),
    .Q(\instrs[7][7] ));
 sg13g2_dfrbp_1 _6968_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net381),
    .D(_0250_),
    .Q_N(_0109_),
    .Q(\datam[3][0] ));
 sg13g2_dfrbp_1 _6969_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net380),
    .D(_0251_),
    .Q_N(_0127_),
    .Q(\datam[3][1] ));
 sg13g2_dfrbp_1 _6970_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net379),
    .D(_0252_),
    .Q_N(_0143_),
    .Q(\datam[3][2] ));
 sg13g2_dfrbp_1 _6971_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net378),
    .D(_0253_),
    .Q_N(_0159_),
    .Q(\datam[3][3] ));
 sg13g2_dfrbp_1 _6972_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net377),
    .D(_0254_),
    .Q_N(_0176_),
    .Q(\datam[3][4] ));
 sg13g2_dfrbp_1 _6973_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net286),
    .D(_0255_),
    .Q_N(_3178_),
    .Q(\datam[3][5] ));
 sg13g2_dfrbp_1 _6974_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net266),
    .D(_0256_),
    .Q_N(_3177_),
    .Q(\datam[3][6] ));
 sg13g2_dfrbp_1 _6975_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net265),
    .D(_0257_),
    .Q_N(_3176_),
    .Q(\datam[3][7] ));
 sg13g2_dfrbp_1 _6976_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net264),
    .D(_0258_),
    .Q_N(_0110_),
    .Q(\datam[4][0] ));
 sg13g2_dfrbp_1 _6977_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net263),
    .D(_0259_),
    .Q_N(_0128_),
    .Q(\datam[4][1] ));
 sg13g2_dfrbp_1 _6978_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net262),
    .D(_0260_),
    .Q_N(_0144_),
    .Q(\datam[4][2] ));
 sg13g2_dfrbp_1 _6979_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net261),
    .D(_0261_),
    .Q_N(_0160_),
    .Q(\datam[4][3] ));
 sg13g2_dfrbp_1 _6980_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net260),
    .D(_0262_),
    .Q_N(_0177_),
    .Q(\datam[4][4] ));
 sg13g2_dfrbp_1 _6981_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net259),
    .D(_0263_),
    .Q_N(_3175_),
    .Q(\datam[4][5] ));
 sg13g2_dfrbp_1 _6982_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net242),
    .D(_0264_),
    .Q_N(_3174_),
    .Q(\datam[4][6] ));
 sg13g2_dfrbp_1 _6983_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net241),
    .D(_0265_),
    .Q_N(_3173_),
    .Q(\datam[4][7] ));
 sg13g2_dfrbp_1 _6984_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net236),
    .D(_0266_),
    .Q_N(_0044_),
    .Q(\instrs[11][0] ));
 sg13g2_dfrbp_1 _6985_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net227),
    .D(_0267_),
    .Q_N(_3172_),
    .Q(\instrs[11][1] ));
 sg13g2_dfrbp_1 _6986_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net170),
    .D(_0268_),
    .Q_N(_3171_),
    .Q(\instrs[11][2] ));
 sg13g2_dfrbp_1 _6987_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net169),
    .D(_0269_),
    .Q_N(_3170_),
    .Q(\instrs[11][3] ));
 sg13g2_dfrbp_1 _6988_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net168),
    .D(net1062),
    .Q_N(_3169_),
    .Q(\instrs[11][4] ));
 sg13g2_dfrbp_1 _6989_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net167),
    .D(_0271_),
    .Q_N(_0064_),
    .Q(\instrs[11][5] ));
 sg13g2_dfrbp_1 _6990_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net166),
    .D(_0272_),
    .Q_N(_3168_),
    .Q(\instrs[11][6] ));
 sg13g2_dfrbp_1 _6991_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net165),
    .D(_0273_),
    .Q_N(_0080_),
    .Q(\instrs[11][7] ));
 sg13g2_dfrbp_1 _6992_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net164),
    .D(_0274_),
    .Q_N(_0108_),
    .Q(\datam[2][0] ));
 sg13g2_dfrbp_1 _6993_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net163),
    .D(_0275_),
    .Q_N(_0126_),
    .Q(\datam[2][1] ));
 sg13g2_dfrbp_1 _6994_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net162),
    .D(_0276_),
    .Q_N(_0142_),
    .Q(\datam[2][2] ));
 sg13g2_dfrbp_1 _6995_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net161),
    .D(_0277_),
    .Q_N(_0158_),
    .Q(\datam[2][3] ));
 sg13g2_dfrbp_1 _6996_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net160),
    .D(_0278_),
    .Q_N(_0175_),
    .Q(\datam[2][4] ));
 sg13g2_dfrbp_1 _6997_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net159),
    .D(_0279_),
    .Q_N(_3167_),
    .Q(\datam[2][5] ));
 sg13g2_dfrbp_1 _6998_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net158),
    .D(_0280_),
    .Q_N(_3166_),
    .Q(\datam[2][6] ));
 sg13g2_dfrbp_1 _6999_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net102),
    .D(_0281_),
    .Q_N(_3206_),
    .Q(\datam[2][7] ));
 sg13g2_dfrbp_1 _7000_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net103),
    .D(net1181),
    .Q_N(_3207_),
    .Q(\C1.next_state_var[0] ));
 sg13g2_dfrbp_1 _7001_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net104),
    .D(net1547),
    .Q_N(_3208_),
    .Q(\C1.next_state_var[1] ));
 sg13g2_dfrbp_1 _7002_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net105),
    .D(net1693),
    .Q_N(_0087_),
    .Q(\C1.next_state_var[2] ));
 sg13g2_dfrbp_1 _7003_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net106),
    .D(net1534),
    .Q_N(_0016_),
    .Q(\C1.next_state_var[3] ));
 sg13g2_dfrbp_1 _7004_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net107),
    .D(net1459),
    .Q_N(_3209_),
    .Q(\C1.next_state_var[4] ));
 sg13g2_dfrbp_1 _7005_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net108),
    .D(_0008_),
    .Q_N(_0015_),
    .Q(\C1.next_state_var[5] ));
 sg13g2_dfrbp_1 _7006_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net156),
    .D(_0009_),
    .Q_N(_3210_),
    .Q(\C1.next_state_var[6] ));
 sg13g2_dfrbp_1 _7007_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net157),
    .D(_0010_),
    .Q_N(_0014_),
    .Q(\C1.next_state_var[7] ));
 sg13g2_dfrbp_1 _7008_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net155),
    .D(_0282_),
    .Q_N(_0103_),
    .Q(\datam[1][0] ));
 sg13g2_dfrbp_1 _7009_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net154),
    .D(_0283_),
    .Q_N(_0125_),
    .Q(\datam[1][1] ));
 sg13g2_dfrbp_1 _7010_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net153),
    .D(_0284_),
    .Q_N(_0141_),
    .Q(\datam[1][2] ));
 sg13g2_dfrbp_1 _7011_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net152),
    .D(_0285_),
    .Q_N(_0157_),
    .Q(\datam[1][3] ));
 sg13g2_dfrbp_1 _7012_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net151),
    .D(_0286_),
    .Q_N(_0174_),
    .Q(\datam[1][4] ));
 sg13g2_dfrbp_1 _7013_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net150),
    .D(_0287_),
    .Q_N(_3165_),
    .Q(\datam[1][5] ));
 sg13g2_dfrbp_1 _7014_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net149),
    .D(_0288_),
    .Q_N(_3164_),
    .Q(\datam[1][6] ));
 sg13g2_dfrbp_1 _7015_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net148),
    .D(_0289_),
    .Q_N(_3163_),
    .Q(\datam[1][7] ));
 sg13g2_dfrbp_1 _7016_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net147),
    .D(_0290_),
    .Q_N(_3162_),
    .Q(\C1.max_count[1] ));
 sg13g2_dfrbp_1 _7017_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net145),
    .D(_0291_),
    .Q_N(_3161_),
    .Q(\C1.max_count[2] ));
 sg13g2_dfrbp_1 _7018_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net143),
    .D(_0292_),
    .Q_N(_3160_),
    .Q(\C1.max_count[3] ));
 sg13g2_dfrbp_1 _7019_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net141),
    .D(_0293_),
    .Q_N(_3159_),
    .Q(\C1.max_count[4] ));
 sg13g2_dfrbp_1 _7020_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net139),
    .D(_0294_),
    .Q_N(_3158_),
    .Q(\C1.max_count[5] ));
 sg13g2_dfrbp_1 _7021_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net137),
    .D(_0295_),
    .Q_N(_3157_),
    .Q(\C1.max_count[6] ));
 sg13g2_dfrbp_1 _7022_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net135),
    .D(_0296_),
    .Q_N(_3156_),
    .Q(\C1.max_count[7] ));
 sg13g2_dfrbp_1 _7023_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net133),
    .D(_0297_),
    .Q_N(_3155_),
    .Q(\C1.max_count[8] ));
 sg13g2_dfrbp_1 _7024_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net131),
    .D(_0298_),
    .Q_N(_3154_),
    .Q(\C1.max_count[9] ));
 sg13g2_dfrbp_1 _7025_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net129),
    .D(_0299_),
    .Q_N(_3153_),
    .Q(\C1.max_count[10] ));
 sg13g2_dfrbp_1 _7026_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net127),
    .D(_0300_),
    .Q_N(_3152_),
    .Q(\C1.max_count[11] ));
 sg13g2_dfrbp_1 _7027_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net125),
    .D(_0301_),
    .Q_N(_0121_),
    .Q(\datam[15][0] ));
 sg13g2_dfrbp_1 _7028_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net124),
    .D(_0302_),
    .Q_N(_0139_),
    .Q(\datam[15][1] ));
 sg13g2_dfrbp_1 _7029_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net123),
    .D(_0303_),
    .Q_N(_0155_),
    .Q(\datam[15][2] ));
 sg13g2_dfrbp_1 _7030_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net122),
    .D(_0304_),
    .Q_N(_0171_),
    .Q(\datam[15][3] ));
 sg13g2_dfrbp_1 _7031_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net121),
    .D(_0305_),
    .Q_N(_0188_),
    .Q(\datam[15][4] ));
 sg13g2_dfrbp_1 _7032_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net120),
    .D(_0306_),
    .Q_N(_3151_),
    .Q(\datam[15][5] ));
 sg13g2_dfrbp_1 _7033_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net119),
    .D(_0307_),
    .Q_N(_3150_),
    .Q(\datam[15][6] ));
 sg13g2_dfrbp_1 _7034_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net118),
    .D(_0308_),
    .Q_N(_3149_),
    .Q(\datam[15][7] ));
 sg13g2_dfrbp_1 _7035_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net117),
    .D(_0309_),
    .Q_N(_0045_),
    .Q(\instrs[12][0] ));
 sg13g2_dfrbp_1 _7036_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net116),
    .D(_0310_),
    .Q_N(_3148_),
    .Q(\instrs[12][1] ));
 sg13g2_dfrbp_1 _7037_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net115),
    .D(_0311_),
    .Q_N(_3147_),
    .Q(\instrs[12][2] ));
 sg13g2_dfrbp_1 _7038_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net114),
    .D(_0312_),
    .Q_N(_3146_),
    .Q(\instrs[12][3] ));
 sg13g2_dfrbp_1 _7039_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net113),
    .D(_0313_),
    .Q_N(_3145_),
    .Q(\instrs[12][4] ));
 sg13g2_dfrbp_1 _7040_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net112),
    .D(_0314_),
    .Q_N(_0065_),
    .Q(\instrs[12][5] ));
 sg13g2_dfrbp_1 _7041_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net111),
    .D(_0315_),
    .Q_N(_3144_),
    .Q(\instrs[12][6] ));
 sg13g2_dfrbp_1 _7042_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net110),
    .D(_0316_),
    .Q_N(_0081_),
    .Q(\instrs[12][7] ));
 sg13g2_dfrbp_1 _7043_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net109),
    .D(_0317_),
    .Q_N(_0046_),
    .Q(\instrs[13][0] ));
 sg13g2_dfrbp_1 _7044_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net100),
    .D(_0318_),
    .Q_N(_3143_),
    .Q(\instrs[13][1] ));
 sg13g2_dfrbp_1 _7045_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net99),
    .D(_0319_),
    .Q_N(_3142_),
    .Q(\instrs[13][2] ));
 sg13g2_dfrbp_1 _7046_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net98),
    .D(_0320_),
    .Q_N(_3141_),
    .Q(\instrs[13][3] ));
 sg13g2_dfrbp_1 _7047_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net97),
    .D(_0321_),
    .Q_N(_3140_),
    .Q(\instrs[13][4] ));
 sg13g2_dfrbp_1 _7048_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net96),
    .D(_0322_),
    .Q_N(_0066_),
    .Q(\instrs[13][5] ));
 sg13g2_dfrbp_1 _7049_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net95),
    .D(_0323_),
    .Q_N(_3139_),
    .Q(\instrs[13][6] ));
 sg13g2_dfrbp_1 _7050_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net94),
    .D(_0324_),
    .Q_N(_0082_),
    .Q(\instrs[13][7] ));
 sg13g2_dfrbp_1 _7051_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net93),
    .D(net1043),
    .Q_N(_0208_),
    .Q(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[0] ));
 sg13g2_dfrbp_1 _7052_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net91),
    .D(_0326_),
    .Q_N(_3138_),
    .Q(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[1] ));
 sg13g2_dfrbp_1 _7053_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net89),
    .D(_0327_),
    .Q_N(_3137_),
    .Q(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[2] ));
 sg13g2_dfrbp_1 _7054_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net171),
    .D(_0328_),
    .Q_N(_3211_),
    .Q(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[3] ));
 sg13g2_dfrbp_1 _7055_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net87),
    .D(net1676),
    .Q_N(_3136_),
    .Q(FpgaPins_Fpga_UART_is_enter_a2));
 sg13g2_dfrbp_1 _7056_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net85),
    .D(net1273),
    .Q_N(_3135_),
    .Q(\C1.counter2[22] ));
 sg13g2_dfrbp_1 _7057_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net84),
    .D(_0330_),
    .Q_N(_3134_),
    .Q(\C1.counter2[23] ));
 sg13g2_dfrbp_1 _7058_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net83),
    .D(_0331_),
    .Q_N(_3133_),
    .Q(\C1.counter2[24] ));
 sg13g2_dfrbp_1 _7059_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net82),
    .D(net1188),
    .Q_N(_3132_),
    .Q(\C1.counter2[25] ));
 sg13g2_dfrbp_1 _7060_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net81),
    .D(_0333_),
    .Q_N(_3131_),
    .Q(\C1.counter2[26] ));
 sg13g2_dfrbp_1 _7061_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net80),
    .D(_0334_),
    .Q_N(_3130_),
    .Q(\C1.counter2[27] ));
 sg13g2_dfrbp_1 _7062_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net79),
    .D(net1288),
    .Q_N(_3129_),
    .Q(\C1.counter2[28] ));
 sg13g2_dfrbp_1 _7063_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net78),
    .D(_0336_),
    .Q_N(_3128_),
    .Q(\C1.counter2[29] ));
 sg13g2_dfrbp_1 _7064_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net77),
    .D(_0337_),
    .Q_N(_3127_),
    .Q(\C1.counter2[30] ));
 sg13g2_dfrbp_1 _7065_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net76),
    .D(net754),
    .Q_N(_3126_),
    .Q(\C1.counter2[31] ));
 sg13g2_dfrbp_1 _7066_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net75),
    .D(net727),
    .Q_N(_0207_),
    .Q(\FpgaPins_Fpga_UART_dptr_a2[0] ));
 sg13g2_dfrbp_1 _7067_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net73),
    .D(_0340_),
    .Q_N(_3125_),
    .Q(\FpgaPins_Fpga_UART_dptr_a2[1] ));
 sg13g2_dfrbp_1 _7068_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net71),
    .D(net746),
    .Q_N(_0203_),
    .Q(\FpgaPins_Fpga_UART_dptr_a2[2] ));
 sg13g2_dfrbp_1 _7069_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net172),
    .D(net730),
    .Q_N(_0204_),
    .Q(\FpgaPins_Fpga_UART_dptr_a2[3] ));
 sg13g2_dfrbp_1 _7070_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net173),
    .D(\FpgaPins_Fpga_FSM_instr_wr_a1[0] ),
    .Q_N(_3212_),
    .Q(\FpgaPins_Fpga_UART_data_a2[0] ));
 sg13g2_dfrbp_1 _7071_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net174),
    .D(\FpgaPins_Fpga_FSM_instr_wr_a1[1] ),
    .Q_N(_3213_),
    .Q(\FpgaPins_Fpga_UART_data_a2[1] ));
 sg13g2_dfrbp_1 _7072_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net175),
    .D(\FpgaPins_Fpga_FSM_instr_wr_a1[2] ),
    .Q_N(_3214_),
    .Q(\FpgaPins_Fpga_UART_data_a2[2] ));
 sg13g2_dfrbp_1 _7073_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net176),
    .D(\FpgaPins_Fpga_FSM_instr_wr_a1[3] ),
    .Q_N(_3215_),
    .Q(\FpgaPins_Fpga_UART_data_a2[3] ));
 sg13g2_dfrbp_1 _7074_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net177),
    .D(\FpgaPins_Fpga_FSM_instr_wr_a1[4] ),
    .Q_N(_3216_),
    .Q(\FpgaPins_Fpga_UART_data_a2[4] ));
 sg13g2_dfrbp_1 _7075_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net178),
    .D(\FpgaPins_Fpga_FSM_instr_wr_a1[5] ),
    .Q_N(_3217_),
    .Q(\FpgaPins_Fpga_UART_data_a2[5] ));
 sg13g2_dfrbp_1 _7076_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net179),
    .D(\FpgaPins_Fpga_FSM_instr_wr_a1[6] ),
    .Q_N(_3218_),
    .Q(\FpgaPins_Fpga_UART_data_a2[6] ));
 sg13g2_dfrbp_1 _7077_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net180),
    .D(\FpgaPins_Fpga_FSM_instr_wr_a1[7] ),
    .Q_N(_3219_),
    .Q(\FpgaPins_Fpga_UART_data_a2[7] ));
 sg13g2_dfrbp_1 _7078_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net181),
    .D(FpgaPins_Fpga_UART_comment_a1),
    .Q_N(_3220_),
    .Q(FpgaPins_Fpga_UART_comment_a2));
 sg13g2_dfrbp_1 _7079_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net182),
    .D(FpgaPins_Fpga_LIPSI_z_a1),
    .Q_N(_3221_),
    .Q(FpgaPins_Fpga_LIPSI_z_a2));
 sg13g2_dfrbp_1 _7080_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net183),
    .D(net944),
    .Q_N(_3222_),
    .Q(FpgaPins_Fpga_LIPSI_reset_a2));
 sg13g2_dfrbp_1 _7081_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net184),
    .D(net911),
    .Q_N(_0020_),
    .Q(\FpgaPins_Fpga_LIPSI_pc_a2[0] ));
 sg13g2_dfrbp_1 _7082_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net185),
    .D(net918),
    .Q_N(_0023_),
    .Q(\FpgaPins_Fpga_LIPSI_pc_a2[1] ));
 sg13g2_dfrbp_1 _7083_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net186),
    .D(\FpgaPins_Fpga_FSM_imem_rd_addr_a1[2] ),
    .Q_N(_0026_),
    .Q(\FpgaPins_Fpga_LIPSI_pc_a2[2] ));
 sg13g2_dfrbp_1 _7084_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net187),
    .D(net891),
    .Q_N(_0029_),
    .Q(\FpgaPins_Fpga_LIPSI_pc_a2[3] ));
 sg13g2_dfrbp_1 _7085_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net188),
    .D(net1104),
    .Q_N(_0194_),
    .Q(\FpgaPins_Fpga_LIPSI_pc_a2[4] ));
 sg13g2_dfrbp_1 _7086_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net189),
    .D(net740),
    .Q_N(_0196_),
    .Q(\FpgaPins_Fpga_LIPSI_pc_a2[5] ));
 sg13g2_dfrbp_1 _7087_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net190),
    .D(net718),
    .Q_N(_0198_),
    .Q(\FpgaPins_Fpga_LIPSI_pc_a2[6] ));
 sg13g2_dfrbp_1 _7088_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net191),
    .D(net736),
    .Q_N(_0200_),
    .Q(\FpgaPins_Fpga_LIPSI_pc_a2[7] ));
 sg13g2_dfrbp_1 _7089_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net192),
    .D(FpgaPins_Fpga_LIPSI_is_st_ind_a1),
    .Q_N(_3223_),
    .Q(FpgaPins_Fpga_LIPSI_is_st_ind_a2));
 sg13g2_dfrbp_1 _7090_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net193),
    .D(FpgaPins_Fpga_LIPSI_is_ret_a1),
    .Q_N(_3224_),
    .Q(FpgaPins_Fpga_LIPSI_is_ret_a2));
 sg13g2_dfrbp_1 _7091_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net194),
    .D(FpgaPins_Fpga_LIPSI_is_ld_ind_a1),
    .Q_N(_3225_),
    .Q(FpgaPins_Fpga_LIPSI_is_ld_ind_a2));
 sg13g2_dfrbp_1 _7092_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net195),
    .D(net692),
    .Q_N(_3226_),
    .Q(FpgaPins_Fpga_LIPSI_is_brz_a3));
 sg13g2_dfrbp_1 _7093_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net196),
    .D(FpgaPins_Fpga_LIPSI_is_brz_a1),
    .Q_N(_3227_),
    .Q(FpgaPins_Fpga_LIPSI_is_brz_a2));
 sg13g2_dfrbp_1 _7094_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net197),
    .D(net701),
    .Q_N(_3228_),
    .Q(FpgaPins_Fpga_LIPSI_is_brnz_a3));
 sg13g2_dfrbp_1 _7095_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net198),
    .D(FpgaPins_Fpga_LIPSI_is_brnz_a1),
    .Q_N(_3229_),
    .Q(FpgaPins_Fpga_LIPSI_is_brnz_a2));
 sg13g2_dfrbp_1 _7096_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net199),
    .D(FpgaPins_Fpga_LIPSI_is_brl_a1),
    .Q_N(_3230_),
    .Q(FpgaPins_Fpga_LIPSI_is_brl_a2));
 sg13g2_dfrbp_1 _7097_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net200),
    .D(net695),
    .Q_N(_3231_),
    .Q(FpgaPins_Fpga_LIPSI_is_br_a3));
 sg13g2_dfrbp_1 _7098_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net201),
    .D(FpgaPins_Fpga_LIPSI_is_br_a1),
    .Q_N(_3232_),
    .Q(FpgaPins_Fpga_LIPSI_is_br_a2));
 sg13g2_dfrbp_1 _7099_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net202),
    .D(FpgaPins_Fpga_LIPSI_is_ALU_imm_a1),
    .Q_N(_3233_),
    .Q(FpgaPins_Fpga_LIPSI_is_ALU_imm_a2));
 sg13g2_dfrbp_1 _7100_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net203),
    .D(FpgaPins_Fpga_LIPSI_is_2cyc_a1),
    .Q_N(_3234_),
    .Q(FpgaPins_Fpga_LIPSI_is_2cyc_a2));
 sg13g2_dfrbp_1 _7101_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net204),
    .D(net859),
    .Q_N(_0021_),
    .Q(\FpgaPins_Fpga_LIPSI_instr_a2[0] ));
 sg13g2_dfrbp_1 _7102_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net205),
    .D(\FpgaPins_Fpga_FSM_instr_a1[1] ),
    .Q_N(_0024_),
    .Q(\FpgaPins_Fpga_LIPSI_instr_a2[1] ));
 sg13g2_dfrbp_1 _7103_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net206),
    .D(\FpgaPins_Fpga_FSM_instr_a1[2] ),
    .Q_N(_0027_),
    .Q(\FpgaPins_Fpga_LIPSI_instr_a2[2] ));
 sg13g2_dfrbp_1 _7104_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net207),
    .D(\FpgaPins_Fpga_FSM_instr_a1[3] ),
    .Q_N(_0030_),
    .Q(\FpgaPins_Fpga_LIPSI_instr_a2[3] ));
 sg13g2_dfrbp_1 _7105_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net208),
    .D(\FpgaPins_Fpga_FSM_instr_a1[4] ),
    .Q_N(_0195_),
    .Q(\FpgaPins_Fpga_LIPSI_instr_a2[4] ));
 sg13g2_dfrbp_1 _7106_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net209),
    .D(net875),
    .Q_N(_0197_),
    .Q(\FpgaPins_Fpga_LIPSI_instr_a2[5] ));
 sg13g2_dfrbp_1 _7107_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net210),
    .D(\FpgaPins_Fpga_FSM_instr_a1[6] ),
    .Q_N(_0199_),
    .Q(\FpgaPins_Fpga_LIPSI_instr_a2[6] ));
 sg13g2_dfrbp_1 _7108_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net211),
    .D(\FpgaPins_Fpga_FSM_instr_a1[7] ),
    .Q_N(_0201_),
    .Q(\FpgaPins_Fpga_LIPSI_instr_a2[7] ));
 sg13g2_dfrbp_1 _7109_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net212),
    .D(FpgaPins_Fpga_LIPSI_exit_a1),
    .Q_N(_3235_),
    .Q(FpgaPins_Fpga_LIPSI_exit_a2));
 sg13g2_dfrbp_1 _7110_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net213),
    .D(\FpgaPins_Fpga_LIPSI_data_wr_a1[0] ),
    .Q_N(_3236_),
    .Q(\FpgaPins_Fpga_LIPSI_data_wr_a2[0] ));
 sg13g2_dfrbp_1 _7111_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net214),
    .D(\FpgaPins_Fpga_LIPSI_data_wr_a1[1] ),
    .Q_N(_3237_),
    .Q(\FpgaPins_Fpga_LIPSI_data_wr_a2[1] ));
 sg13g2_dfrbp_1 _7112_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net215),
    .D(\FpgaPins_Fpga_LIPSI_data_wr_a1[2] ),
    .Q_N(_3238_),
    .Q(\FpgaPins_Fpga_LIPSI_data_wr_a2[2] ));
 sg13g2_dfrbp_1 _7113_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net216),
    .D(\FpgaPins_Fpga_LIPSI_data_wr_a1[3] ),
    .Q_N(_3239_),
    .Q(\FpgaPins_Fpga_LIPSI_data_wr_a2[3] ));
 sg13g2_dfrbp_1 _7114_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net217),
    .D(\FpgaPins_Fpga_LIPSI_data_wr_a1[4] ),
    .Q_N(_3240_),
    .Q(\FpgaPins_Fpga_LIPSI_data_wr_a2[4] ));
 sg13g2_dfrbp_1 _7115_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net218),
    .D(\FpgaPins_Fpga_LIPSI_data_wr_a1[5] ),
    .Q_N(_3241_),
    .Q(\FpgaPins_Fpga_LIPSI_data_wr_a2[5] ));
 sg13g2_dfrbp_1 _7116_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net219),
    .D(\FpgaPins_Fpga_LIPSI_data_wr_a1[6] ),
    .Q_N(_3242_),
    .Q(\FpgaPins_Fpga_LIPSI_data_wr_a2[6] ));
 sg13g2_dfrbp_1 _7117_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net220),
    .D(\FpgaPins_Fpga_LIPSI_data_wr_a1[7] ),
    .Q_N(_3243_),
    .Q(\FpgaPins_Fpga_LIPSI_data_wr_a2[7] ));
 sg13g2_dfrbp_1 _7118_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net221),
    .D(net1643),
    .Q_N(_0104_),
    .Q(\FpgaPins_Fpga_LIPSI_data_a2[0] ));
 sg13g2_dfrbp_1 _7119_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net222),
    .D(\FpgaPins_Fpga_FSM_data_a1[1] ),
    .Q_N(_0106_),
    .Q(\FpgaPins_Fpga_LIPSI_data_a2[1] ));
 sg13g2_dfrbp_1 _7120_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net223),
    .D(\FpgaPins_Fpga_FSM_data_a1[2] ),
    .Q_N(_3244_),
    .Q(\FpgaPins_Fpga_LIPSI_data_a2[2] ));
 sg13g2_dfrbp_1 _7121_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net224),
    .D(\FpgaPins_Fpga_FSM_data_a1[3] ),
    .Q_N(_0032_),
    .Q(\FpgaPins_Fpga_LIPSI_data_a2[3] ));
 sg13g2_dfrbp_1 _7122_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net225),
    .D(\FpgaPins_Fpga_FSM_data_a1[4] ),
    .Q_N(_3245_),
    .Q(\FpgaPins_Fpga_LIPSI_data_a2[4] ));
 sg13g2_dfrbp_1 _7123_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net226),
    .D(\FpgaPins_Fpga_FSM_data_a1[5] ),
    .Q_N(_3246_),
    .Q(\FpgaPins_Fpga_LIPSI_data_a2[5] ));
 sg13g2_dfrbp_1 _7124_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net228),
    .D(\FpgaPins_Fpga_FSM_data_a1[6] ),
    .Q_N(_3247_),
    .Q(\FpgaPins_Fpga_LIPSI_data_a2[6] ));
 sg13g2_dfrbp_1 _7125_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net69),
    .D(\FpgaPins_Fpga_FSM_data_a1[7] ),
    .Q_N(_3124_),
    .Q(\FpgaPins_Fpga_LIPSI_data_a2[7] ));
 sg13g2_dfrbp_1 _7126_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net229),
    .D(_0343_),
    .Q_N(_0122_),
    .Q(FpgaPins_Fpga_LIPSI_c_a2));
 sg13g2_dfrbp_1 _7127_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net230),
    .D(\FpgaPins_Fpga_LIPSI_acc_a1[0] ),
    .Q_N(_0022_),
    .Q(\FpgaPins_Fpga_LIPSI_acc_a2[0] ));
 sg13g2_dfrbp_1 _7128_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net231),
    .D(\FpgaPins_Fpga_LIPSI_acc_a1[1] ),
    .Q_N(_0025_),
    .Q(\FpgaPins_Fpga_LIPSI_acc_a2[1] ));
 sg13g2_dfrbp_1 _7129_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net232),
    .D(\FpgaPins_Fpga_LIPSI_acc_a1[2] ),
    .Q_N(_0028_),
    .Q(\FpgaPins_Fpga_LIPSI_acc_a2[2] ));
 sg13g2_dfrbp_1 _7130_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net233),
    .D(\FpgaPins_Fpga_LIPSI_acc_a1[3] ),
    .Q_N(_0031_),
    .Q(\FpgaPins_Fpga_LIPSI_acc_a2[3] ));
 sg13g2_dfrbp_1 _7131_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net234),
    .D(\FpgaPins_Fpga_LIPSI_acc_a1[4] ),
    .Q_N(_0172_),
    .Q(\FpgaPins_Fpga_LIPSI_acc_a2[4] ));
 sg13g2_dfrbp_1 _7132_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net235),
    .D(\FpgaPins_Fpga_LIPSI_acc_a1[5] ),
    .Q_N(_0189_),
    .Q(\FpgaPins_Fpga_LIPSI_acc_a2[5] ));
 sg13g2_dfrbp_1 _7133_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net237),
    .D(\FpgaPins_Fpga_LIPSI_acc_a1[6] ),
    .Q_N(_0190_),
    .Q(\FpgaPins_Fpga_LIPSI_acc_a2[6] ));
 sg13g2_dfrbp_1 _7134_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net67),
    .D(\FpgaPins_Fpga_LIPSI_acc_a1[7] ),
    .Q_N(_0123_),
    .Q(\FpgaPins_Fpga_LIPSI_acc_a2[7] ));
 sg13g2_dfrbp_1 _7135_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net238),
    .D(_0344_),
    .Q_N(_0191_),
    .Q(FpgaPins_Fpga_UART_first_byte_a2));
 sg13g2_dfrbp_1 _7136_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net239),
    .D(net708),
    .Q_N(_3248_),
    .Q(\FpgaPins_Fpga_GAME_state_a4[0] ));
 sg13g2_dfrbp_1 _7137_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net240),
    .D(net707),
    .Q_N(_3249_),
    .Q(\FpgaPins_Fpga_GAME_state_a4[1] ));
 sg13g2_dfrbp_1 _7138_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net243),
    .D(net706),
    .Q_N(_3250_),
    .Q(\FpgaPins_Fpga_GAME_state_a3[0] ));
 sg13g2_dfrbp_1 _7139_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net65),
    .D(net704),
    .Q_N(_3123_),
    .Q(\FpgaPins_Fpga_GAME_state_a3[1] ));
 sg13g2_dfrbp_1 _7140_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net64),
    .D(_0345_),
    .Q_N(_3122_),
    .Q(\FpgaPins_Fpga_GAME_state_a2[0] ));
 sg13g2_dfrbp_1 _7141_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net244),
    .D(_0346_),
    .Q_N(_3251_),
    .Q(\FpgaPins_Fpga_GAME_state_a2[1] ));
 sg13g2_dfrbp_1 _7142_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net245),
    .D(net697),
    .Q_N(_3252_),
    .Q(\FpgaPins_Fpga_GAME_score_a4[0] ));
 sg13g2_dfrbp_1 _7143_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net246),
    .D(net693),
    .Q_N(_3253_),
    .Q(\FpgaPins_Fpga_GAME_score_a4[1] ));
 sg13g2_dfrbp_1 _7144_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net247),
    .D(net698),
    .Q_N(_3254_),
    .Q(\FpgaPins_Fpga_GAME_score_a4[2] ));
 sg13g2_dfrbp_1 _7145_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net248),
    .D(net703),
    .Q_N(_3255_),
    .Q(\FpgaPins_Fpga_GAME_score_a4[3] ));
 sg13g2_dfrbp_1 _7146_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net249),
    .D(net702),
    .Q_N(_3256_),
    .Q(\FpgaPins_Fpga_GAME_score_a4[4] ));
 sg13g2_dfrbp_1 _7147_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net250),
    .D(net700),
    .Q_N(_3257_),
    .Q(\FpgaPins_Fpga_GAME_score_a4[5] ));
 sg13g2_dfrbp_1 _7148_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net251),
    .D(net696),
    .Q_N(_3258_),
    .Q(\FpgaPins_Fpga_GAME_score_a4[6] ));
 sg13g2_dfrbp_1 _7149_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net252),
    .D(net699),
    .Q_N(_3259_),
    .Q(\FpgaPins_Fpga_GAME_score_a4[7] ));
 sg13g2_dfrbp_1 _7150_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net253),
    .D(net720),
    .Q_N(_3260_),
    .Q(\FpgaPins_Fpga_GAME_score_a3[0] ));
 sg13g2_dfrbp_1 _7151_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net254),
    .D(net712),
    .Q_N(_3261_),
    .Q(\FpgaPins_Fpga_GAME_score_a3[1] ));
 sg13g2_dfrbp_1 _7152_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net255),
    .D(net713),
    .Q_N(_3262_),
    .Q(\FpgaPins_Fpga_GAME_score_a3[2] ));
 sg13g2_dfrbp_1 _7153_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net256),
    .D(net715),
    .Q_N(_3263_),
    .Q(\FpgaPins_Fpga_GAME_score_a3[3] ));
 sg13g2_dfrbp_1 _7154_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net257),
    .D(net716),
    .Q_N(_3264_),
    .Q(\FpgaPins_Fpga_GAME_score_a3[4] ));
 sg13g2_dfrbp_1 _7155_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net258),
    .D(net710),
    .Q_N(_3265_),
    .Q(\FpgaPins_Fpga_GAME_score_a3[5] ));
 sg13g2_dfrbp_1 _7156_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net267),
    .D(net721),
    .Q_N(_3266_),
    .Q(\FpgaPins_Fpga_GAME_score_a3[6] ));
 sg13g2_dfrbp_1 _7157_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net62),
    .D(net714),
    .Q_N(_3121_),
    .Q(\FpgaPins_Fpga_GAME_score_a3[7] ));
 sg13g2_dfrbp_1 _7158_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net60),
    .D(_0347_),
    .Q_N(_3120_),
    .Q(\FpgaPins_Fpga_GAME_score_a2[0] ));
 sg13g2_dfrbp_1 _7159_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net58),
    .D(_0348_),
    .Q_N(_3119_),
    .Q(\FpgaPins_Fpga_GAME_score_a2[1] ));
 sg13g2_dfrbp_1 _7160_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net56),
    .D(_0349_),
    .Q_N(_3118_),
    .Q(\FpgaPins_Fpga_GAME_score_a2[2] ));
 sg13g2_dfrbp_1 _7161_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net54),
    .D(_0350_),
    .Q_N(_3117_),
    .Q(\FpgaPins_Fpga_GAME_score_a2[3] ));
 sg13g2_dfrbp_1 _7162_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net52),
    .D(_0351_),
    .Q_N(_3116_),
    .Q(\FpgaPins_Fpga_GAME_score_a2[4] ));
 sg13g2_dfrbp_1 _7163_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net50),
    .D(_0352_),
    .Q_N(_3115_),
    .Q(\FpgaPins_Fpga_GAME_score_a2[5] ));
 sg13g2_dfrbp_1 _7164_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net48),
    .D(_0353_),
    .Q_N(_3114_),
    .Q(\FpgaPins_Fpga_GAME_score_a2[6] ));
 sg13g2_dfrbp_1 _7165_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net268),
    .D(net1493),
    .Q_N(_3267_),
    .Q(\FpgaPins_Fpga_GAME_score_a2[7] ));
 sg13g2_dfrbp_1 _7166_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net269),
    .D(net1000),
    .Q_N(_3268_),
    .Q(FpgaPins_Fpga_GAME_right_btn_a2));
 sg13g2_dfrbp_1 _7167_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net270),
    .D(FpgaPins_Fpga_GAME_reset_a1),
    .Q_N(_0017_),
    .Q(FpgaPins_Fpga_GAME_reset_a2));
 sg13g2_dfrbp_1 _7168_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net271),
    .D(net4),
    .Q_N(_3269_),
    .Q(FpgaPins_Fpga_GAME_left_btn_a2));
 sg13g2_dfrbp_1 _7169_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net272),
    .D(net719),
    .Q_N(_3270_),
    .Q(\FpgaPins_Fpga_GAME_led_output_a3[0] ));
 sg13g2_dfrbp_1 _7170_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net273),
    .D(net723),
    .Q_N(_3271_),
    .Q(\FpgaPins_Fpga_GAME_led_output_a3[1] ));
 sg13g2_dfrbp_1 _7171_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net274),
    .D(net711),
    .Q_N(_3272_),
    .Q(\FpgaPins_Fpga_GAME_led_output_a3[2] ));
 sg13g2_dfrbp_1 _7172_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net275),
    .D(net722),
    .Q_N(_3273_),
    .Q(\FpgaPins_Fpga_GAME_led_output_a3[3] ));
 sg13g2_dfrbp_1 _7173_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net276),
    .D(net1006),
    .Q_N(_3274_),
    .Q(\FpgaPins_Fpga_GAME_led_output_a3[4] ));
 sg13g2_dfrbp_1 _7174_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net277),
    .D(net1013),
    .Q_N(_3275_),
    .Q(\FpgaPins_Fpga_GAME_led_output_a3[5] ));
 sg13g2_dfrbp_1 _7175_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net278),
    .D(net742),
    .Q_N(_3276_),
    .Q(\FpgaPins_Fpga_GAME_led_output_a3[6] ));
 sg13g2_dfrbp_1 _7176_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net279),
    .D(net724),
    .Q_N(_3277_),
    .Q(\FpgaPins_Fpga_GAME_led_output_a3[7] ));
 sg13g2_dfrbp_1 _7177_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net280),
    .D(\FpgaPins_Fpga_GAME_led_output_a1[0] ),
    .Q_N(_3278_),
    .Q(\FpgaPins_Fpga_GAME_led_output_a2[0] ));
 sg13g2_dfrbp_1 _7178_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net281),
    .D(\FpgaPins_Fpga_GAME_led_output_a1[1] ),
    .Q_N(_3279_),
    .Q(\FpgaPins_Fpga_GAME_led_output_a2[1] ));
 sg13g2_dfrbp_1 _7179_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net282),
    .D(net1670),
    .Q_N(_3280_),
    .Q(\FpgaPins_Fpga_GAME_led_output_a2[2] ));
 sg13g2_dfrbp_1 _7180_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net283),
    .D(\FpgaPins_Fpga_GAME_led_output_a1[3] ),
    .Q_N(_3281_),
    .Q(\FpgaPins_Fpga_GAME_led_output_a2[3] ));
 sg13g2_dfrbp_1 _7181_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net284),
    .D(net1688),
    .Q_N(_3282_),
    .Q(\FpgaPins_Fpga_GAME_led_output_a2[4] ));
 sg13g2_dfrbp_1 _7182_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net285),
    .D(\FpgaPins_Fpga_GAME_led_output_a1[5] ),
    .Q_N(_3283_),
    .Q(\FpgaPins_Fpga_GAME_led_output_a2[5] ));
 sg13g2_dfrbp_1 _7183_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net287),
    .D(\FpgaPins_Fpga_GAME_led_output_a1[6] ),
    .Q_N(_3284_),
    .Q(\FpgaPins_Fpga_GAME_led_output_a2[6] ));
 sg13g2_dfrbp_1 _7184_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net46),
    .D(\FpgaPins_Fpga_GAME_led_output_a1[7] ),
    .Q_N(_3113_),
    .Q(\FpgaPins_Fpga_GAME_led_output_a2[7] ));
 sg13g2_dfrbp_1 _7185_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net288),
    .D(net1730),
    .Q_N(_3285_),
    .Q(FpgaPins_Fpga_GAME_forward_a2));
 sg13g2_dfrbp_1 _7186_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net289),
    .D(\FpgaPins_Fpga_GAME_count_speed4_a1[0] ),
    .Q_N(_3286_),
    .Q(\FpgaPins_Fpga_GAME_count_speed4_a2[0] ));
 sg13g2_dfrbp_1 _7187_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net290),
    .D(\FpgaPins_Fpga_GAME_count_speed4_a1[1] ),
    .Q_N(_3287_),
    .Q(\FpgaPins_Fpga_GAME_count_speed4_a2[1] ));
 sg13g2_dfrbp_1 _7188_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net291),
    .D(net1166),
    .Q_N(_3288_),
    .Q(\FpgaPins_Fpga_GAME_count_speed4_a2[2] ));
 sg13g2_dfrbp_1 _7189_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net292),
    .D(\FpgaPins_Fpga_GAME_count_speed4_a1[3] ),
    .Q_N(_3289_),
    .Q(\FpgaPins_Fpga_GAME_count_speed4_a2[3] ));
 sg13g2_dfrbp_1 _7190_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net293),
    .D(\FpgaPins_Fpga_GAME_count_speed4_a1[4] ),
    .Q_N(_3290_),
    .Q(\FpgaPins_Fpga_GAME_count_speed4_a2[4] ));
 sg13g2_dfrbp_1 _7191_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net294),
    .D(\FpgaPins_Fpga_GAME_count_speed4_a1[5] ),
    .Q_N(_3291_),
    .Q(\FpgaPins_Fpga_GAME_count_speed4_a2[5] ));
 sg13g2_dfrbp_1 _7192_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net295),
    .D(\FpgaPins_Fpga_GAME_count_speed4_a1[6] ),
    .Q_N(_3292_),
    .Q(\FpgaPins_Fpga_GAME_count_speed4_a2[6] ));
 sg13g2_dfrbp_1 _7193_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net296),
    .D(\FpgaPins_Fpga_GAME_count_speed4_a1[7] ),
    .Q_N(_3293_),
    .Q(\FpgaPins_Fpga_GAME_count_speed4_a2[7] ));
 sg13g2_dfrbp_1 _7194_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net297),
    .D(\FpgaPins_Fpga_GAME_count_speed4_a1[8] ),
    .Q_N(_3294_),
    .Q(\FpgaPins_Fpga_GAME_count_speed4_a2[8] ));
 sg13g2_dfrbp_1 _7195_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net298),
    .D(\FpgaPins_Fpga_GAME_count_speed4_a1[9] ),
    .Q_N(_3295_),
    .Q(\FpgaPins_Fpga_GAME_count_speed4_a2[9] ));
 sg13g2_dfrbp_1 _7196_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net299),
    .D(\FpgaPins_Fpga_GAME_count_speed4_a1[10] ),
    .Q_N(_3296_),
    .Q(\FpgaPins_Fpga_GAME_count_speed4_a2[10] ));
 sg13g2_dfrbp_1 _7197_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net300),
    .D(\FpgaPins_Fpga_GAME_count_speed4_a1[11] ),
    .Q_N(_3297_),
    .Q(\FpgaPins_Fpga_GAME_count_speed4_a2[11] ));
 sg13g2_dfrbp_1 _7198_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net301),
    .D(\FpgaPins_Fpga_GAME_count_speed4_a1[12] ),
    .Q_N(_3298_),
    .Q(\FpgaPins_Fpga_GAME_count_speed4_a2[12] ));
 sg13g2_dfrbp_1 _7199_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net302),
    .D(\FpgaPins_Fpga_GAME_count_speed4_a1[13] ),
    .Q_N(_3299_),
    .Q(\FpgaPins_Fpga_GAME_count_speed4_a2[13] ));
 sg13g2_dfrbp_1 _7200_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net303),
    .D(\FpgaPins_Fpga_GAME_count_speed4_a1[14] ),
    .Q_N(_0049_),
    .Q(\FpgaPins_Fpga_GAME_count_speed4_a2[14] ));
 sg13g2_dfrbp_1 _7201_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net304),
    .D(net1499),
    .Q_N(_3300_),
    .Q(\FpgaPins_Fpga_GAME_count_speed4_a2[15] ));
 sg13g2_dfrbp_1 _7202_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net305),
    .D(\FpgaPins_Fpga_GAME_count_speed4_a1[16] ),
    .Q_N(_3301_),
    .Q(\FpgaPins_Fpga_GAME_count_speed4_a2[16] ));
 sg13g2_dfrbp_1 _7203_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net306),
    .D(\FpgaPins_Fpga_GAME_count_speed4_a1[17] ),
    .Q_N(_3302_),
    .Q(\FpgaPins_Fpga_GAME_count_speed4_a2[17] ));
 sg13g2_dfrbp_1 _7204_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net307),
    .D(net1031),
    .Q_N(_3303_),
    .Q(\FpgaPins_Fpga_GAME_count_speed4_a2[18] ));
 sg13g2_dfrbp_1 _7205_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net308),
    .D(\FpgaPins_Fpga_GAME_count_speed3_a1[0] ),
    .Q_N(_3304_),
    .Q(\FpgaPins_Fpga_GAME_count_speed3_a2[0] ));
 sg13g2_dfrbp_1 _7206_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net309),
    .D(net1092),
    .Q_N(_3305_),
    .Q(\FpgaPins_Fpga_GAME_count_speed3_a2[1] ));
 sg13g2_dfrbp_1 _7207_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net310),
    .D(\FpgaPins_Fpga_GAME_count_speed3_a1[2] ),
    .Q_N(_3306_),
    .Q(\FpgaPins_Fpga_GAME_count_speed3_a2[2] ));
 sg13g2_dfrbp_1 _7208_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net311),
    .D(\FpgaPins_Fpga_GAME_count_speed3_a1[3] ),
    .Q_N(_3307_),
    .Q(\FpgaPins_Fpga_GAME_count_speed3_a2[3] ));
 sg13g2_dfrbp_1 _7209_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net312),
    .D(\FpgaPins_Fpga_GAME_count_speed3_a1[4] ),
    .Q_N(_3308_),
    .Q(\FpgaPins_Fpga_GAME_count_speed3_a2[4] ));
 sg13g2_dfrbp_1 _7210_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net313),
    .D(\FpgaPins_Fpga_GAME_count_speed3_a1[5] ),
    .Q_N(_3309_),
    .Q(\FpgaPins_Fpga_GAME_count_speed3_a2[5] ));
 sg13g2_dfrbp_1 _7211_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net314),
    .D(\FpgaPins_Fpga_GAME_count_speed3_a1[6] ),
    .Q_N(_3310_),
    .Q(\FpgaPins_Fpga_GAME_count_speed3_a2[6] ));
 sg13g2_dfrbp_1 _7212_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net315),
    .D(\FpgaPins_Fpga_GAME_count_speed3_a1[7] ),
    .Q_N(_3311_),
    .Q(\FpgaPins_Fpga_GAME_count_speed3_a2[7] ));
 sg13g2_dfrbp_1 _7213_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net316),
    .D(\FpgaPins_Fpga_GAME_count_speed3_a1[8] ),
    .Q_N(_3312_),
    .Q(\FpgaPins_Fpga_GAME_count_speed3_a2[8] ));
 sg13g2_dfrbp_1 _7214_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net317),
    .D(net1559),
    .Q_N(_3313_),
    .Q(\FpgaPins_Fpga_GAME_count_speed3_a2[9] ));
 sg13g2_dfrbp_1 _7215_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net318),
    .D(\FpgaPins_Fpga_GAME_count_speed3_a1[10] ),
    .Q_N(_3314_),
    .Q(\FpgaPins_Fpga_GAME_count_speed3_a2[10] ));
 sg13g2_dfrbp_1 _7216_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net319),
    .D(\FpgaPins_Fpga_GAME_count_speed3_a1[11] ),
    .Q_N(_3315_),
    .Q(\FpgaPins_Fpga_GAME_count_speed3_a2[11] ));
 sg13g2_dfrbp_1 _7217_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net320),
    .D(net1396),
    .Q_N(_3316_),
    .Q(\FpgaPins_Fpga_GAME_count_speed3_a2[12] ));
 sg13g2_dfrbp_1 _7218_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net321),
    .D(\FpgaPins_Fpga_GAME_count_speed3_a1[13] ),
    .Q_N(_3317_),
    .Q(\FpgaPins_Fpga_GAME_count_speed3_a2[13] ));
 sg13g2_dfrbp_1 _7219_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net322),
    .D(\FpgaPins_Fpga_GAME_count_speed3_a1[14] ),
    .Q_N(_0050_),
    .Q(\FpgaPins_Fpga_GAME_count_speed3_a2[14] ));
 sg13g2_dfrbp_1 _7220_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net323),
    .D(\FpgaPins_Fpga_GAME_count_speed3_a1[15] ),
    .Q_N(_3318_),
    .Q(\FpgaPins_Fpga_GAME_count_speed3_a2[15] ));
 sg13g2_dfrbp_1 _7221_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net324),
    .D(\FpgaPins_Fpga_GAME_count_speed3_a1[16] ),
    .Q_N(_3319_),
    .Q(\FpgaPins_Fpga_GAME_count_speed3_a2[16] ));
 sg13g2_dfrbp_1 _7222_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net325),
    .D(\FpgaPins_Fpga_GAME_count_speed3_a1[17] ),
    .Q_N(_3320_),
    .Q(\FpgaPins_Fpga_GAME_count_speed3_a2[17] ));
 sg13g2_dfrbp_1 _7223_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net326),
    .D(\FpgaPins_Fpga_GAME_count_speed3_a1[18] ),
    .Q_N(_3321_),
    .Q(\FpgaPins_Fpga_GAME_count_speed3_a2[18] ));
 sg13g2_dfrbp_1 _7224_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net327),
    .D(net1267),
    .Q_N(_3322_),
    .Q(\FpgaPins_Fpga_GAME_count_speed3_a2[19] ));
 sg13g2_dfrbp_1 _7225_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net328),
    .D(\FpgaPins_Fpga_GAME_count_speed2_a1[0] ),
    .Q_N(_3323_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[0] ));
 sg13g2_dfrbp_1 _7226_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net329),
    .D(\FpgaPins_Fpga_GAME_count_speed2_a1[1] ),
    .Q_N(_3324_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[1] ));
 sg13g2_dfrbp_1 _7227_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net330),
    .D(net1129),
    .Q_N(_3325_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[2] ));
 sg13g2_dfrbp_1 _7228_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net331),
    .D(\FpgaPins_Fpga_GAME_count_speed2_a1[3] ),
    .Q_N(_3326_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[3] ));
 sg13g2_dfrbp_1 _7229_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net332),
    .D(\FpgaPins_Fpga_GAME_count_speed2_a1[4] ),
    .Q_N(_3327_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[4] ));
 sg13g2_dfrbp_1 _7230_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net333),
    .D(\FpgaPins_Fpga_GAME_count_speed2_a1[5] ),
    .Q_N(_3328_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[5] ));
 sg13g2_dfrbp_1 _7231_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net334),
    .D(\FpgaPins_Fpga_GAME_count_speed2_a1[6] ),
    .Q_N(_3329_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[6] ));
 sg13g2_dfrbp_1 _7232_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net335),
    .D(\FpgaPins_Fpga_GAME_count_speed2_a1[7] ),
    .Q_N(_3330_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[7] ));
 sg13g2_dfrbp_1 _7233_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net336),
    .D(\FpgaPins_Fpga_GAME_count_speed2_a1[8] ),
    .Q_N(_3331_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[8] ));
 sg13g2_dfrbp_1 _7234_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net337),
    .D(\FpgaPins_Fpga_GAME_count_speed2_a1[9] ),
    .Q_N(_3332_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[9] ));
 sg13g2_dfrbp_1 _7235_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net338),
    .D(\FpgaPins_Fpga_GAME_count_speed2_a1[10] ),
    .Q_N(_3333_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[10] ));
 sg13g2_dfrbp_1 _7236_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net339),
    .D(\FpgaPins_Fpga_GAME_count_speed2_a1[11] ),
    .Q_N(_3334_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[11] ));
 sg13g2_dfrbp_1 _7237_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net340),
    .D(\FpgaPins_Fpga_GAME_count_speed2_a1[12] ),
    .Q_N(_3335_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[12] ));
 sg13g2_dfrbp_1 _7238_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net341),
    .D(\FpgaPins_Fpga_GAME_count_speed2_a1[13] ),
    .Q_N(_3336_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[13] ));
 sg13g2_dfrbp_1 _7239_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net342),
    .D(net1348),
    .Q_N(_0051_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[14] ));
 sg13g2_dfrbp_1 _7240_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net343),
    .D(\FpgaPins_Fpga_GAME_count_speed2_a1[15] ),
    .Q_N(_3337_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[15] ));
 sg13g2_dfrbp_1 _7241_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net344),
    .D(\FpgaPins_Fpga_GAME_count_speed2_a1[16] ),
    .Q_N(_3338_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[16] ));
 sg13g2_dfrbp_1 _7242_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net345),
    .D(net1445),
    .Q_N(_3339_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[17] ));
 sg13g2_dfrbp_1 _7243_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net346),
    .D(\FpgaPins_Fpga_GAME_count_speed2_a1[18] ),
    .Q_N(_3340_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[18] ));
 sg13g2_dfrbp_1 _7244_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net347),
    .D(net1195),
    .Q_N(_3341_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[19] ));
 sg13g2_dfrbp_1 _7245_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net348),
    .D(\FpgaPins_Fpga_GAME_count_speed2_a1[20] ),
    .Q_N(_0052_),
    .Q(\FpgaPins_Fpga_GAME_count_speed2_a2[20] ));
 sg13g2_dfrbp_1 _7246_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net349),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a1[0] ),
    .Q_N(_3342_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[0] ));
 sg13g2_dfrbp_1 _7247_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net350),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a1[1] ),
    .Q_N(_3343_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[1] ));
 sg13g2_dfrbp_1 _7248_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net351),
    .D(net1434),
    .Q_N(_3344_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[2] ));
 sg13g2_dfrbp_1 _7249_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net352),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a1[3] ),
    .Q_N(_3345_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[3] ));
 sg13g2_dfrbp_1 _7250_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net353),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a1[4] ),
    .Q_N(_3346_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[4] ));
 sg13g2_dfrbp_1 _7251_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net354),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a1[5] ),
    .Q_N(_3347_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[5] ));
 sg13g2_dfrbp_1 _7252_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net355),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a1[6] ),
    .Q_N(_3348_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[6] ));
 sg13g2_dfrbp_1 _7253_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net356),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a1[7] ),
    .Q_N(_3349_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[7] ));
 sg13g2_dfrbp_1 _7254_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net357),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a1[8] ),
    .Q_N(_3350_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[8] ));
 sg13g2_dfrbp_1 _7255_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net358),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a1[9] ),
    .Q_N(_3351_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[9] ));
 sg13g2_dfrbp_1 _7256_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net359),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a1[10] ),
    .Q_N(_3352_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[10] ));
 sg13g2_dfrbp_1 _7257_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net360),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a1[11] ),
    .Q_N(_3353_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[11] ));
 sg13g2_dfrbp_1 _7258_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net361),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a1[12] ),
    .Q_N(_3354_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[12] ));
 sg13g2_dfrbp_1 _7259_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net362),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a1[13] ),
    .Q_N(_3355_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[13] ));
 sg13g2_dfrbp_1 _7260_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net363),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a1[14] ),
    .Q_N(_3356_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[14] ));
 sg13g2_dfrbp_1 _7261_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net364),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a1[15] ),
    .Q_N(_3357_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[15] ));
 sg13g2_dfrbp_1 _7262_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net365),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a1[16] ),
    .Q_N(_3358_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[16] ));
 sg13g2_dfrbp_1 _7263_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net366),
    .D(net1466),
    .Q_N(_3359_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[17] ));
 sg13g2_dfrbp_1 _7264_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net367),
    .D(net1305),
    .Q_N(_3360_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[18] ));
 sg13g2_dfrbp_1 _7265_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net368),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a1[19] ),
    .Q_N(_3361_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[19] ));
 sg13g2_dfrbp_1 _7266_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net369),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a1[20] ),
    .Q_N(_3362_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[20] ));
 sg13g2_dfrbp_1 _7267_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net370),
    .D(net1362),
    .Q_N(_3363_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[21] ));
 sg13g2_dfrbp_1 _7268_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net371),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a1[22] ),
    .Q_N(_3364_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[22] ));
 sg13g2_dfrbp_1 _7269_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net372),
    .D(\FpgaPins_Fpga_GAME_count_speed1_a1[23] ),
    .Q_N(_3365_),
    .Q(\FpgaPins_Fpga_GAME_count_speed1_a2[23] ));
 sg13g2_dfrbp_1 _7270_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net373),
    .D(net1314),
    .Q_N(_3366_),
    .Q(FpgaPins_Fpga_GAME_clk_pulse4_a2));
 sg13g2_dfrbp_1 _7271_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net374),
    .D(net1160),
    .Q_N(_3367_),
    .Q(FpgaPins_Fpga_GAME_clk_pulse3_a2));
 sg13g2_dfrbp_1 _7272_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net375),
    .D(net1479),
    .Q_N(_3368_),
    .Q(FpgaPins_Fpga_GAME_clk_pulse2_a2));
 sg13g2_dfrbp_1 _7273_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net376),
    .D(net1528),
    .Q_N(_0019_),
    .Q(FpgaPins_Fpga_GAME_clk_pulse1_a2));
 sg13g2_dfrbp_1 _7274_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net543),
    .D(net705),
    .Q_N(_3369_),
    .Q(FpgaPins_Fpga_GAME_clk_pulse_a3));
 sg13g2_dfrbp_1 _7275_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net44),
    .D(FpgaPins_Fpga_GAME_clk_pulse_a1),
    .Q_N(_3112_),
    .Q(FpgaPins_Fpga_GAME_clk_pulse_a2));
 sg13g2_dfrbp_1 _7276_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net42),
    .D(_0356_),
    .Q_N(_0119_),
    .Q(\datam[13][0] ));
 sg13g2_dfrbp_1 _7277_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net41),
    .D(_0357_),
    .Q_N(_0137_),
    .Q(\datam[13][1] ));
 sg13g2_dfrbp_1 _7278_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net40),
    .D(_0358_),
    .Q_N(_0153_),
    .Q(\datam[13][2] ));
 sg13g2_dfrbp_1 _7279_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net39),
    .D(_0359_),
    .Q_N(_0169_),
    .Q(\datam[13][3] ));
 sg13g2_dfrbp_1 _7280_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net38),
    .D(_0360_),
    .Q_N(_0186_),
    .Q(\datam[13][4] ));
 sg13g2_dfrbp_1 _7281_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net37),
    .D(_0361_),
    .Q_N(_3111_),
    .Q(\datam[13][5] ));
 sg13g2_dfrbp_1 _7282_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net36),
    .D(_0362_),
    .Q_N(_3110_),
    .Q(\datam[13][6] ));
 sg13g2_dfrbp_1 _7283_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net35),
    .D(_0363_),
    .Q_N(_3109_),
    .Q(\datam[13][7] ));
 sg13g2_dfrbp_1 _7284_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net34),
    .D(_0364_),
    .Q_N(_0039_),
    .Q(\instrs[6][0] ));
 sg13g2_dfrbp_1 _7285_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net33),
    .D(_0365_),
    .Q_N(_3108_),
    .Q(\instrs[6][1] ));
 sg13g2_dfrbp_1 _7286_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net32),
    .D(_0366_),
    .Q_N(_3107_),
    .Q(\instrs[6][2] ));
 sg13g2_dfrbp_1 _7287_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net31),
    .D(_0367_),
    .Q_N(_3106_),
    .Q(\instrs[6][3] ));
 sg13g2_dfrbp_1 _7288_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net30),
    .D(net1332),
    .Q_N(_3105_),
    .Q(\instrs[6][4] ));
 sg13g2_dfrbp_1 _7289_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net29),
    .D(_0369_),
    .Q_N(_0059_),
    .Q(\instrs[6][5] ));
 sg13g2_dfrbp_1 _7290_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net25),
    .D(_0370_),
    .Q_N(_3104_),
    .Q(\instrs[6][6] ));
 sg13g2_dfrbp_1 _7291_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net691),
    .D(_0371_),
    .Q_N(_0075_),
    .Q(\instrs[6][7] ));
 sg13g2_dfrbp_1 _7292_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net690),
    .D(_0372_),
    .Q_N(_0118_),
    .Q(\datam[12][0] ));
 sg13g2_dfrbp_1 _7293_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net689),
    .D(_0373_),
    .Q_N(_0136_),
    .Q(\datam[12][1] ));
 sg13g2_dfrbp_1 _7294_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net688),
    .D(_0374_),
    .Q_N(_0152_),
    .Q(\datam[12][2] ));
 sg13g2_dfrbp_1 _7295_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net687),
    .D(_0375_),
    .Q_N(_0168_),
    .Q(\datam[12][3] ));
 sg13g2_dfrbp_1 _7296_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net686),
    .D(_0376_),
    .Q_N(_0185_),
    .Q(\datam[12][4] ));
 sg13g2_dfrbp_1 _7297_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net685),
    .D(_0377_),
    .Q_N(_3103_),
    .Q(\datam[12][5] ));
 sg13g2_dfrbp_1 _7298_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net684),
    .D(_0378_),
    .Q_N(_3102_),
    .Q(\datam[12][6] ));
 sg13g2_dfrbp_1 _7299_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net683),
    .D(_0379_),
    .Q_N(_3101_),
    .Q(\datam[12][7] ));
 sg13g2_dfrbp_1 _7300_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net682),
    .D(_0380_),
    .Q_N(_0038_),
    .Q(\instrs[5][0] ));
 sg13g2_dfrbp_1 _7301_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net681),
    .D(_0381_),
    .Q_N(_3100_),
    .Q(\instrs[5][1] ));
 sg13g2_dfrbp_1 _7302_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net680),
    .D(_0382_),
    .Q_N(_3099_),
    .Q(\instrs[5][2] ));
 sg13g2_dfrbp_1 _7303_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net679),
    .D(_0383_),
    .Q_N(_3098_),
    .Q(\instrs[5][3] ));
 sg13g2_dfrbp_1 _7304_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net678),
    .D(_0384_),
    .Q_N(_3097_),
    .Q(\instrs[5][4] ));
 sg13g2_dfrbp_1 _7305_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net677),
    .D(_0385_),
    .Q_N(_0058_),
    .Q(\instrs[5][5] ));
 sg13g2_dfrbp_1 _7306_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net676),
    .D(_0386_),
    .Q_N(_3096_),
    .Q(\instrs[5][6] ));
 sg13g2_dfrbp_1 _7307_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net675),
    .D(_0387_),
    .Q_N(_0074_),
    .Q(\instrs[5][7] ));
 sg13g2_dfrbp_1 _7308_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net674),
    .D(_0388_),
    .Q_N(_0117_),
    .Q(\datam[11][0] ));
 sg13g2_dfrbp_1 _7309_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net673),
    .D(_0389_),
    .Q_N(_0135_),
    .Q(\datam[11][1] ));
 sg13g2_dfrbp_1 _7310_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net672),
    .D(_0390_),
    .Q_N(_0151_),
    .Q(\datam[11][2] ));
 sg13g2_dfrbp_1 _7311_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net671),
    .D(_0391_),
    .Q_N(_0167_),
    .Q(\datam[11][3] ));
 sg13g2_dfrbp_1 _7312_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net670),
    .D(_0392_),
    .Q_N(_0184_),
    .Q(\datam[11][4] ));
 sg13g2_dfrbp_1 _7313_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net669),
    .D(_0393_),
    .Q_N(_3095_),
    .Q(\datam[11][5] ));
 sg13g2_dfrbp_1 _7314_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net668),
    .D(_0394_),
    .Q_N(_3094_),
    .Q(\datam[11][6] ));
 sg13g2_dfrbp_1 _7315_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net667),
    .D(_0395_),
    .Q_N(_3093_),
    .Q(\datam[11][7] ));
 sg13g2_dfrbp_1 _7316_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net666),
    .D(_0396_),
    .Q_N(_0037_),
    .Q(\instrs[4][0] ));
 sg13g2_dfrbp_1 _7317_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net665),
    .D(_0397_),
    .Q_N(_3092_),
    .Q(\instrs[4][1] ));
 sg13g2_dfrbp_1 _7318_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net664),
    .D(_0398_),
    .Q_N(_3091_),
    .Q(\instrs[4][2] ));
 sg13g2_dfrbp_1 _7319_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net663),
    .D(_0399_),
    .Q_N(_3090_),
    .Q(\instrs[4][3] ));
 sg13g2_dfrbp_1 _7320_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net662),
    .D(_0400_),
    .Q_N(_3089_),
    .Q(\instrs[4][4] ));
 sg13g2_dfrbp_1 _7321_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net661),
    .D(_0401_),
    .Q_N(_0057_),
    .Q(\instrs[4][5] ));
 sg13g2_dfrbp_1 _7322_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net660),
    .D(_0402_),
    .Q_N(_3088_),
    .Q(\instrs[4][6] ));
 sg13g2_dfrbp_1 _7323_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net659),
    .D(_0403_),
    .Q_N(_0073_),
    .Q(\instrs[4][7] ));
 sg13g2_dfrbp_1 _7324_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net658),
    .D(_0404_),
    .Q_N(_0116_),
    .Q(\datam[10][0] ));
 sg13g2_dfrbp_1 _7325_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net657),
    .D(_0405_),
    .Q_N(_0134_),
    .Q(\datam[10][1] ));
 sg13g2_dfrbp_1 _7326_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net656),
    .D(_0406_),
    .Q_N(_0150_),
    .Q(\datam[10][2] ));
 sg13g2_dfrbp_1 _7327_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net655),
    .D(_0407_),
    .Q_N(_0166_),
    .Q(\datam[10][3] ));
 sg13g2_dfrbp_1 _7328_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net654),
    .D(_0408_),
    .Q_N(_0183_),
    .Q(\datam[10][4] ));
 sg13g2_dfrbp_1 _7329_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net653),
    .D(_0409_),
    .Q_N(_3087_),
    .Q(\datam[10][5] ));
 sg13g2_dfrbp_1 _7330_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net652),
    .D(_0410_),
    .Q_N(_3086_),
    .Q(\datam[10][6] ));
 sg13g2_dfrbp_1 _7331_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net651),
    .D(_0411_),
    .Q_N(_3085_),
    .Q(\datam[10][7] ));
 sg13g2_dfrbp_1 _7332_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net650),
    .D(_0412_),
    .Q_N(_0036_),
    .Q(\instrs[3][0] ));
 sg13g2_dfrbp_1 _7333_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net649),
    .D(_0413_),
    .Q_N(_3084_),
    .Q(\instrs[3][1] ));
 sg13g2_dfrbp_1 _7334_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net648),
    .D(_0414_),
    .Q_N(_3083_),
    .Q(\instrs[3][2] ));
 sg13g2_dfrbp_1 _7335_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net647),
    .D(_0415_),
    .Q_N(_3082_),
    .Q(\instrs[3][3] ));
 sg13g2_dfrbp_1 _7336_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net646),
    .D(_0416_),
    .Q_N(_3081_),
    .Q(\instrs[3][4] ));
 sg13g2_dfrbp_1 _7337_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net645),
    .D(_0417_),
    .Q_N(_0056_),
    .Q(\instrs[3][5] ));
 sg13g2_dfrbp_1 _7338_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net644),
    .D(_0418_),
    .Q_N(_3080_),
    .Q(\instrs[3][6] ));
 sg13g2_dfrbp_1 _7339_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net643),
    .D(_0419_),
    .Q_N(_0072_),
    .Q(\instrs[3][7] ));
 sg13g2_dfrbp_1 _7340_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net642),
    .D(_0420_),
    .Q_N(_0102_),
    .Q(\datam[0][0] ));
 sg13g2_dfrbp_1 _7341_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net641),
    .D(_0421_),
    .Q_N(_0124_),
    .Q(\datam[0][1] ));
 sg13g2_dfrbp_1 _7342_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net640),
    .D(_0422_),
    .Q_N(_0140_),
    .Q(\datam[0][2] ));
 sg13g2_dfrbp_1 _7343_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net639),
    .D(_0423_),
    .Q_N(_0156_),
    .Q(\datam[0][3] ));
 sg13g2_dfrbp_1 _7344_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net638),
    .D(_0424_),
    .Q_N(_0173_),
    .Q(\datam[0][4] ));
 sg13g2_dfrbp_1 _7345_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net637),
    .D(_0425_),
    .Q_N(_3079_),
    .Q(\datam[0][5] ));
 sg13g2_dfrbp_1 _7346_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net636),
    .D(_0426_),
    .Q_N(_3078_),
    .Q(\datam[0][6] ));
 sg13g2_dfrbp_1 _7347_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net635),
    .D(_0427_),
    .Q_N(_3077_),
    .Q(\datam[0][7] ));
 sg13g2_dfrbp_1 _7348_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net634),
    .D(_0428_),
    .Q_N(_0114_),
    .Q(\datam[8][0] ));
 sg13g2_dfrbp_1 _7349_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net633),
    .D(_0429_),
    .Q_N(_0132_),
    .Q(\datam[8][1] ));
 sg13g2_dfrbp_1 _7350_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net632),
    .D(_0430_),
    .Q_N(_0148_),
    .Q(\datam[8][2] ));
 sg13g2_dfrbp_1 _7351_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net631),
    .D(_0431_),
    .Q_N(_0164_),
    .Q(\datam[8][3] ));
 sg13g2_dfrbp_1 _7352_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net630),
    .D(_0432_),
    .Q_N(_0181_),
    .Q(\datam[8][4] ));
 sg13g2_dfrbp_1 _7353_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net629),
    .D(_0433_),
    .Q_N(_3076_),
    .Q(\datam[8][5] ));
 sg13g2_dfrbp_1 _7354_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net628),
    .D(_0434_),
    .Q_N(_3075_),
    .Q(\datam[8][6] ));
 sg13g2_dfrbp_1 _7355_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net627),
    .D(_0435_),
    .Q_N(_3074_),
    .Q(\datam[8][7] ));
 sg13g2_dfrbp_1 _7356_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net626),
    .D(_0436_),
    .Q_N(_0113_),
    .Q(\datam[7][0] ));
 sg13g2_dfrbp_1 _7357_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net625),
    .D(_0437_),
    .Q_N(_0131_),
    .Q(\datam[7][1] ));
 sg13g2_dfrbp_1 _7358_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net624),
    .D(_0438_),
    .Q_N(_0147_),
    .Q(\datam[7][2] ));
 sg13g2_dfrbp_1 _7359_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net623),
    .D(_0439_),
    .Q_N(_0163_),
    .Q(\datam[7][3] ));
 sg13g2_dfrbp_1 _7360_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net622),
    .D(_0440_),
    .Q_N(_0180_),
    .Q(\datam[7][4] ));
 sg13g2_dfrbp_1 _7361_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net621),
    .D(_0441_),
    .Q_N(_3073_),
    .Q(\datam[7][5] ));
 sg13g2_dfrbp_1 _7362_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net620),
    .D(_0442_),
    .Q_N(_3072_),
    .Q(\datam[7][6] ));
 sg13g2_dfrbp_1 _7363_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net619),
    .D(_0443_),
    .Q_N(_3071_),
    .Q(\datam[7][7] ));
 sg13g2_dfrbp_1 _7364_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net618),
    .D(_0444_),
    .Q_N(_0112_),
    .Q(\datam[6][0] ));
 sg13g2_dfrbp_1 _7365_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net617),
    .D(_0445_),
    .Q_N(_0130_),
    .Q(\datam[6][1] ));
 sg13g2_dfrbp_1 _7366_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net616),
    .D(_0446_),
    .Q_N(_0146_),
    .Q(\datam[6][2] ));
 sg13g2_dfrbp_1 _7367_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net613),
    .D(_0447_),
    .Q_N(_0162_),
    .Q(\datam[6][3] ));
 sg13g2_dfrbp_1 _7368_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net612),
    .D(_0448_),
    .Q_N(_0179_),
    .Q(\datam[6][4] ));
 sg13g2_dfrbp_1 _7369_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net611),
    .D(_0449_),
    .Q_N(_3070_),
    .Q(\datam[6][5] ));
 sg13g2_dfrbp_1 _7370_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net610),
    .D(_0450_),
    .Q_N(_3069_),
    .Q(\datam[6][6] ));
 sg13g2_dfrbp_1 _7371_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net609),
    .D(_0451_),
    .Q_N(_3068_),
    .Q(\datam[6][7] ));
 sg13g2_dfrbp_1 _7372_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net608),
    .D(_0452_),
    .Q_N(_0035_),
    .Q(\instrs[2][0] ));
 sg13g2_dfrbp_1 _7373_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net607),
    .D(_0453_),
    .Q_N(_3067_),
    .Q(\instrs[2][1] ));
 sg13g2_dfrbp_1 _7374_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net606),
    .D(_0454_),
    .Q_N(_3066_),
    .Q(\instrs[2][2] ));
 sg13g2_dfrbp_1 _7375_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net605),
    .D(_0455_),
    .Q_N(_3065_),
    .Q(\instrs[2][3] ));
 sg13g2_dfrbp_1 _7376_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net604),
    .D(_0456_),
    .Q_N(_3064_),
    .Q(\instrs[2][4] ));
 sg13g2_dfrbp_1 _7377_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net603),
    .D(_0457_),
    .Q_N(_0055_),
    .Q(\instrs[2][5] ));
 sg13g2_dfrbp_1 _7378_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net602),
    .D(_0458_),
    .Q_N(_3063_),
    .Q(\instrs[2][6] ));
 sg13g2_dfrbp_1 _7379_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net601),
    .D(_0459_),
    .Q_N(_0071_),
    .Q(\instrs[2][7] ));
 sg13g2_dfrbp_1 _7380_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net600),
    .D(_0460_),
    .Q_N(_0034_),
    .Q(\instrs[1][0] ));
 sg13g2_dfrbp_1 _7381_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net599),
    .D(_0461_),
    .Q_N(_3062_),
    .Q(\instrs[1][1] ));
 sg13g2_dfrbp_1 _7382_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net598),
    .D(_0462_),
    .Q_N(_3061_),
    .Q(\instrs[1][2] ));
 sg13g2_dfrbp_1 _7383_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net597),
    .D(_0463_),
    .Q_N(_3060_),
    .Q(\instrs[1][3] ));
 sg13g2_dfrbp_1 _7384_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net596),
    .D(_0464_),
    .Q_N(_3059_),
    .Q(\instrs[1][4] ));
 sg13g2_dfrbp_1 _7385_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net595),
    .D(_0465_),
    .Q_N(_0054_),
    .Q(\instrs[1][5] ));
 sg13g2_dfrbp_1 _7386_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net594),
    .D(_0466_),
    .Q_N(_3058_),
    .Q(\instrs[1][6] ));
 sg13g2_dfrbp_1 _7387_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net593),
    .D(_0467_),
    .Q_N(_0070_),
    .Q(\instrs[1][7] ));
 sg13g2_dfrbp_1 _7388_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net592),
    .D(_0468_),
    .Q_N(_0048_),
    .Q(\instrs[15][0] ));
 sg13g2_dfrbp_1 _7389_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net591),
    .D(_0469_),
    .Q_N(_3057_),
    .Q(\instrs[15][1] ));
 sg13g2_dfrbp_1 _7390_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net590),
    .D(_0470_),
    .Q_N(_3056_),
    .Q(\instrs[15][2] ));
 sg13g2_dfrbp_1 _7391_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net589),
    .D(_0471_),
    .Q_N(_3055_),
    .Q(\instrs[15][3] ));
 sg13g2_dfrbp_1 _7392_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net588),
    .D(net1371),
    .Q_N(_3054_),
    .Q(\instrs[15][4] ));
 sg13g2_dfrbp_1 _7393_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net587),
    .D(_0473_),
    .Q_N(_0068_),
    .Q(\instrs[15][5] ));
 sg13g2_dfrbp_1 _7394_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net586),
    .D(_0474_),
    .Q_N(_3053_),
    .Q(\instrs[15][6] ));
 sg13g2_dfrbp_1 _7395_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net585),
    .D(_0475_),
    .Q_N(_0084_),
    .Q(\instrs[15][7] ));
 sg13g2_dfrbp_1 _7396_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net584),
    .D(_0476_),
    .Q_N(_0111_),
    .Q(\datam[5][0] ));
 sg13g2_dfrbp_1 _7397_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net583),
    .D(_0477_),
    .Q_N(_0129_),
    .Q(\datam[5][1] ));
 sg13g2_dfrbp_1 _7398_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net582),
    .D(_0478_),
    .Q_N(_0145_),
    .Q(\datam[5][2] ));
 sg13g2_dfrbp_1 _7399_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net581),
    .D(_0479_),
    .Q_N(_0161_),
    .Q(\datam[5][3] ));
 sg13g2_dfrbp_1 _7400_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net580),
    .D(_0480_),
    .Q_N(_0178_),
    .Q(\datam[5][4] ));
 sg13g2_dfrbp_1 _7401_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net579),
    .D(_0481_),
    .Q_N(_3052_),
    .Q(\datam[5][5] ));
 sg13g2_dfrbp_1 _7402_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net578),
    .D(_0482_),
    .Q_N(_3051_),
    .Q(\datam[5][6] ));
 sg13g2_dfrbp_1 _7403_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net577),
    .D(_0483_),
    .Q_N(_3050_),
    .Q(\datam[5][7] ));
 sg13g2_dfrbp_1 _7404_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net576),
    .D(_0484_),
    .Q_N(_0115_),
    .Q(\datam[9][0] ));
 sg13g2_dfrbp_1 _7405_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net575),
    .D(_0485_),
    .Q_N(_0133_),
    .Q(\datam[9][1] ));
 sg13g2_dfrbp_1 _7406_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net574),
    .D(_0486_),
    .Q_N(_0149_),
    .Q(\datam[9][2] ));
 sg13g2_dfrbp_1 _7407_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net573),
    .D(_0487_),
    .Q_N(_0165_),
    .Q(\datam[9][3] ));
 sg13g2_dfrbp_1 _7408_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net572),
    .D(_0488_),
    .Q_N(_0182_),
    .Q(\datam[9][4] ));
 sg13g2_dfrbp_1 _7409_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net571),
    .D(_0489_),
    .Q_N(_3049_),
    .Q(\datam[9][5] ));
 sg13g2_dfrbp_1 _7410_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net570),
    .D(_0490_),
    .Q_N(_3048_),
    .Q(\datam[9][6] ));
 sg13g2_dfrbp_1 _7411_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net569),
    .D(_0491_),
    .Q_N(_3047_),
    .Q(\datam[9][7] ));
 sg13g2_dfrbp_1 _7412_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net568),
    .D(_0492_),
    .Q_N(_3046_),
    .Q(\C1.counter2[0] ));
 sg13g2_dfrbp_1 _7413_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net567),
    .D(_0493_),
    .Q_N(_3045_),
    .Q(\C1.counter2[1] ));
 sg13g2_dfrbp_1 _7414_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net566),
    .D(_0494_),
    .Q_N(_3044_),
    .Q(\C1.counter2[2] ));
 sg13g2_dfrbp_1 _7415_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net565),
    .D(_0495_),
    .Q_N(_3043_),
    .Q(\C1.counter2[3] ));
 sg13g2_dfrbp_1 _7416_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net564),
    .D(_0496_),
    .Q_N(_3042_),
    .Q(\C1.counter2[4] ));
 sg13g2_dfrbp_1 _7417_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net563),
    .D(_0497_),
    .Q_N(_3041_),
    .Q(\C1.counter2[5] ));
 sg13g2_dfrbp_1 _7418_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net562),
    .D(_0498_),
    .Q_N(_3040_),
    .Q(\C1.counter2[6] ));
 sg13g2_dfrbp_1 _7419_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net561),
    .D(_0499_),
    .Q_N(_3039_),
    .Q(\C1.counter2[7] ));
 sg13g2_dfrbp_1 _7420_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net560),
    .D(_0500_),
    .Q_N(_3038_),
    .Q(\C1.counter2[8] ));
 sg13g2_dfrbp_1 _7421_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net559),
    .D(_0501_),
    .Q_N(_3037_),
    .Q(\C1.counter2[9] ));
 sg13g2_dfrbp_1 _7422_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net558),
    .D(_0502_),
    .Q_N(_3036_),
    .Q(\C1.counter2[10] ));
 sg13g2_dfrbp_1 _7423_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net557),
    .D(_0503_),
    .Q_N(_3035_),
    .Q(\C1.counter2[11] ));
 sg13g2_dfrbp_1 _7424_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net556),
    .D(_0504_),
    .Q_N(_3034_),
    .Q(\C1.counter2[12] ));
 sg13g2_dfrbp_1 _7425_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net555),
    .D(_0505_),
    .Q_N(_3033_),
    .Q(\C1.counter2[13] ));
 sg13g2_dfrbp_1 _7426_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net554),
    .D(_0506_),
    .Q_N(_3032_),
    .Q(\C1.counter2[14] ));
 sg13g2_dfrbp_1 _7427_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net553),
    .D(_0507_),
    .Q_N(_3031_),
    .Q(\C1.counter2[15] ));
 sg13g2_dfrbp_1 _7428_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net552),
    .D(_0508_),
    .Q_N(_3030_),
    .Q(\C1.counter2[16] ));
 sg13g2_dfrbp_1 _7429_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net542),
    .D(_0509_),
    .Q_N(_3029_),
    .Q(\C1.counter2[17] ));
 sg13g2_dfrbp_1 _7430_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net541),
    .D(_0510_),
    .Q_N(_3028_),
    .Q(\C1.counter2[18] ));
 sg13g2_dfrbp_1 _7431_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net540),
    .D(_0511_),
    .Q_N(_3027_),
    .Q(\C1.counter2[19] ));
 sg13g2_dfrbp_1 _7432_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net539),
    .D(_0512_),
    .Q_N(_3026_),
    .Q(\C1.counter2[20] ));
 sg13g2_dfrbp_1 _7433_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net538),
    .D(_0513_),
    .Q_N(_3025_),
    .Q(\C1.counter2[21] ));
 sg13g2_dfrbp_1 _7434_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net537),
    .D(net1048),
    .Q_N(_0047_),
    .Q(\instrs[14][0] ));
 sg13g2_dfrbp_1 _7435_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net536),
    .D(_0515_),
    .Q_N(_3024_),
    .Q(\instrs[14][1] ));
 sg13g2_dfrbp_1 _7436_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net535),
    .D(_0516_),
    .Q_N(_3023_),
    .Q(\instrs[14][2] ));
 sg13g2_dfrbp_1 _7437_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net534),
    .D(_0517_),
    .Q_N(_3022_),
    .Q(\instrs[14][3] ));
 sg13g2_dfrbp_1 _7438_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net533),
    .D(_0518_),
    .Q_N(_3021_),
    .Q(\instrs[14][4] ));
 sg13g2_dfrbp_1 _7439_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net532),
    .D(_0519_),
    .Q_N(_0067_),
    .Q(\instrs[14][5] ));
 sg13g2_dfrbp_1 _7440_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net531),
    .D(_0520_),
    .Q_N(_3020_),
    .Q(\instrs[14][6] ));
 sg13g2_dfrbp_1 _7441_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net544),
    .D(_0521_),
    .Q_N(_0083_),
    .Q(\instrs[14][7] ));
 sg13g2_dfrbp_1 _7442_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net545),
    .D(net798),
    .Q_N(_0105_),
    .Q(\FpgaPins_Fpga_LIPSI_dptr_a2[0] ));
 sg13g2_dfrbp_1 _7443_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net546),
    .D(net818),
    .Q_N(_0107_),
    .Q(\FpgaPins_Fpga_LIPSI_dptr_a2[1] ));
 sg13g2_dfrbp_1 _7444_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net547),
    .D(net797),
    .Q_N(_3370_),
    .Q(\FpgaPins_Fpga_LIPSI_dptr_a2[2] ));
 sg13g2_dfrbp_1 _7445_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net548),
    .D(net794),
    .Q_N(_3371_),
    .Q(\FpgaPins_Fpga_LIPSI_dptr_a2[3] ));
 sg13g2_dfrbp_1 _7446_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net549),
    .D(\FpgaPins_Fpga_GAME_win_a1[1] ),
    .Q_N(_0086_),
    .Q(\FpgaPins_Fpga_GAME_win_a2[1] ));
 sg13g2_dfrbp_1 _7447_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net550),
    .D(\FpgaPins_Fpga_GAME_win_a1[0] ),
    .Q_N(_0018_),
    .Q(\FpgaPins_Fpga_GAME_win_a2[2] ));
 sg13g2_dfrbp_1 _7448_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net551),
    .D(_0011_),
    .Q_N(_3372_),
    .Q(\FpgaPins_Fpga_GAME_speed_level_a2[1] ));
 sg13g2_dfrbp_1 _7449_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net614),
    .D(_0012_),
    .Q_N(_3373_),
    .Q(\FpgaPins_Fpga_GAME_speed_level_a2[2] ));
 sg13g2_dfrbp_1 _7450_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net530),
    .D(_0013_),
    .Q_N(_3019_),
    .Q(\FpgaPins_Fpga_GAME_speed_level_a2[3] ));
 sg13g2_dfrbp_1 _7451_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net529),
    .D(_0522_),
    .Q_N(_0206_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[0] ));
 sg13g2_dfrbp_1 _7452_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net528),
    .D(_0523_),
    .Q_N(_3018_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[1] ));
 sg13g2_dfrbp_1 _7453_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net527),
    .D(net1177),
    .Q_N(_3017_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[2] ));
 sg13g2_dfrbp_1 _7454_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net526),
    .D(_0525_),
    .Q_N(_3016_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[3] ));
 sg13g2_dfrbp_1 _7455_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net525),
    .D(_0526_),
    .Q_N(_3015_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[4] ));
 sg13g2_dfrbp_1 _7456_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net524),
    .D(_0527_),
    .Q_N(_3014_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[5] ));
 sg13g2_dfrbp_1 _7457_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net523),
    .D(_0528_),
    .Q_N(_3013_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[6] ));
 sg13g2_dfrbp_1 _7458_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net522),
    .D(_0529_),
    .Q_N(_3012_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[7] ));
 sg13g2_dfrbp_1 _7459_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net521),
    .D(_0530_),
    .Q_N(_3011_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[8] ));
 sg13g2_dfrbp_1 _7460_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net520),
    .D(net1526),
    .Q_N(_3010_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[9] ));
 sg13g2_dfrbp_1 _7461_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net519),
    .D(_0532_),
    .Q_N(_3009_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[10] ));
 sg13g2_dfrbp_1 _7462_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net518),
    .D(_0533_),
    .Q_N(_3008_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[11] ));
 sg13g2_dfrbp_1 _7463_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net517),
    .D(net1531),
    .Q_N(_3007_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[12] ));
 sg13g2_dfrbp_1 _7464_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net516),
    .D(net1724),
    .Q_N(_3006_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[13] ));
 sg13g2_dfrbp_1 _7465_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net515),
    .D(net1497),
    .Q_N(_3005_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[14] ));
 sg13g2_dfrbp_1 _7466_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net514),
    .D(net1388),
    .Q_N(_3004_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[15] ));
 sg13g2_dfrbp_1 _7467_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net513),
    .D(net1245),
    .Q_N(_3003_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[16] ));
 sg13g2_dfrbp_1 _7468_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net512),
    .D(_0539_),
    .Q_N(_3002_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[17] ));
 sg13g2_dfrbp_1 _7469_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net511),
    .D(_0540_),
    .Q_N(_3001_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[18] ));
 sg13g2_dfrbp_1 _7470_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net510),
    .D(_0541_),
    .Q_N(_3000_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[19] ));
 sg13g2_dfrbp_1 _7471_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net509),
    .D(_0542_),
    .Q_N(_2999_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[20] ));
 sg13g2_dfrbp_1 _7472_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net508),
    .D(_0543_),
    .Q_N(_2998_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[21] ));
 sg13g2_dfrbp_1 _7473_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net507),
    .D(_0544_),
    .Q_N(_2997_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[22] ));
 sg13g2_dfrbp_1 _7474_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net506),
    .D(net1413),
    .Q_N(_2996_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[23] ));
 sg13g2_dfrbp_1 _7475_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net505),
    .D(_0546_),
    .Q_N(_2995_),
    .Q(\FpgaPins_Fpga_GAME_wait_counter_a2[24] ));
 sg13g2_dfrbp_1 _7476_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net504),
    .D(_0547_),
    .Q_N(_0042_),
    .Q(\instrs[9][0] ));
 sg13g2_dfrbp_1 _7477_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net503),
    .D(_0548_),
    .Q_N(_2994_),
    .Q(\instrs[9][1] ));
 sg13g2_dfrbp_1 _7478_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net502),
    .D(_0549_),
    .Q_N(_2993_),
    .Q(\instrs[9][2] ));
 sg13g2_dfrbp_1 _7479_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net501),
    .D(_0550_),
    .Q_N(_2992_),
    .Q(\instrs[9][3] ));
 sg13g2_dfrbp_1 _7480_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net500),
    .D(_0551_),
    .Q_N(_2991_),
    .Q(\instrs[9][4] ));
 sg13g2_dfrbp_1 _7481_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net499),
    .D(_0552_),
    .Q_N(_0062_),
    .Q(\instrs[9][5] ));
 sg13g2_dfrbp_1 _7482_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net498),
    .D(_0553_),
    .Q_N(_2990_),
    .Q(\instrs[9][6] ));
 sg13g2_dfrbp_1 _7483_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net497),
    .D(_0554_),
    .Q_N(_0078_),
    .Q(\instrs[9][7] ));
 sg13g2_dfrbp_1 _7484_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net496),
    .D(_0555_),
    .Q_N(_2989_),
    .Q(\C1.heating ));
 sg13g2_dfrbp_1 _7485_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net494),
    .D(_0556_),
    .Q_N(_2988_),
    .Q(\C1.pouring ));
 sg13g2_dfrbp_1 _7486_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net492),
    .D(_0557_),
    .Q_N(_2987_),
    .Q(\C1.rinse_status ));
 sg13g2_dfrbp_1 _7487_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net490),
    .D(_0558_),
    .Q_N(_2986_),
    .Q(\C1.dry_status ));
 sg13g2_dfrbp_1 _7488_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net488),
    .D(_0559_),
    .Q_N(_0085_),
    .Q(\C1.counter1[0] ));
 sg13g2_dfrbp_1 _7489_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net487),
    .D(_0560_),
    .Q_N(_0088_),
    .Q(\C1.counter1[1] ));
 sg13g2_dfrbp_1 _7490_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net486),
    .D(_0561_),
    .Q_N(_0089_),
    .Q(\C1.counter1[2] ));
 sg13g2_dfrbp_1 _7491_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net485),
    .D(_0562_),
    .Q_N(_0090_),
    .Q(\C1.counter1[3] ));
 sg13g2_dfrbp_1 _7492_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net484),
    .D(_0563_),
    .Q_N(_0091_),
    .Q(\C1.counter1[4] ));
 sg13g2_dfrbp_1 _7493_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net483),
    .D(_0564_),
    .Q_N(_0092_),
    .Q(\C1.counter1[5] ));
 sg13g2_dfrbp_1 _7494_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net482),
    .D(_0565_),
    .Q_N(_0093_),
    .Q(\C1.counter1[6] ));
 sg13g2_dfrbp_1 _7495_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net481),
    .D(_0566_),
    .Q_N(_0094_),
    .Q(\C1.counter1[7] ));
 sg13g2_dfrbp_1 _7496_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net480),
    .D(_0567_),
    .Q_N(_0095_),
    .Q(\C1.counter1[8] ));
 sg13g2_dfrbp_1 _7497_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net479),
    .D(_0568_),
    .Q_N(_0096_),
    .Q(\C1.counter1[9] ));
 sg13g2_dfrbp_1 _7498_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net478),
    .D(_0569_),
    .Q_N(_0097_),
    .Q(\C1.counter1[10] ));
 sg13g2_dfrbp_1 _7499_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net477),
    .D(_0570_),
    .Q_N(_0098_),
    .Q(\C1.counter1[11] ));
 sg13g2_dfrbp_1 _7500_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net476),
    .D(net1380),
    .Q_N(_2985_),
    .Q(\C1.waiting ));
 sg13g2_dfrbp_1 _7501_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net474),
    .D(net1236),
    .Q_N(_2984_),
    .Q(\C1.prog_op ));
 sg13g2_dfrbp_1 _7502_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net472),
    .D(net1110),
    .Q_N(_2983_),
    .Q(\C1.level_op ));
 sg13g2_dfrbp_1 _7503_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net470),
    .D(net1124),
    .Q_N(_2982_),
    .Q(\C1.temp_op ));
 sg13g2_dfrbp_1 _7504_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net468),
    .D(_0575_),
    .Q_N(_2981_),
    .Q(\C1.dura_op ));
 sg13g2_dfrbp_1 _7505_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net466),
    .D(_0576_),
    .Q_N(_2980_),
    .Q(\C1.timer[0] ));
 sg13g2_dfrbp_1 _7506_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net464),
    .D(_0577_),
    .Q_N(_2979_),
    .Q(\C1.timer[1] ));
 sg13g2_dfrbp_1 _7507_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net462),
    .D(_0578_),
    .Q_N(_2978_),
    .Q(\C1.Program[0] ));
 sg13g2_dfrbp_1 _7508_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net460),
    .D(_0579_),
    .Q_N(_2977_),
    .Q(\C1.Program[1] ));
 sg13g2_dfrbp_1 _7509_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net458),
    .D(_0580_),
    .Q_N(_2976_),
    .Q(\C1.temp[0] ));
 sg13g2_dfrbp_1 _7510_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net456),
    .D(_0581_),
    .Q_N(_2975_),
    .Q(\C1.temp[1] ));
 sg13g2_dfrbp_1 _7511_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net454),
    .D(_0582_),
    .Q_N(_2974_),
    .Q(\C1.level[0] ));
 sg13g2_dfrbp_1 _7512_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net615),
    .D(_0583_),
    .Q_N(_3374_),
    .Q(\C1.level[1] ));
 sg13g2_dfrbp_1 _7513_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net425),
    .D(net694),
    .Q_N(_0101_),
    .Q(\uart_rx_1.r_Rx_Data ));
 sg13g2_dfrbp_1 _7514_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net452),
    .D(net7),
    .Q_N(_2973_),
    .Q(\uart_rx_1.r_Rx_Data_R ));
 sg13g2_dfrbp_1 _7515_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net450),
    .D(net1660),
    .Q_N(_2972_),
    .Q(\uart_rx_1.r_Rx_DV ));
 sg13g2_dfrbp_1 _7516_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net448),
    .D(_0585_),
    .Q_N(_0192_),
    .Q(\uart_rx_1.r_Rx_Byte[0] ));
 sg13g2_dfrbp_1 _7517_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net446),
    .D(_0586_),
    .Q_N(_2971_),
    .Q(\uart_rx_1.r_Rx_Byte[1] ));
 sg13g2_dfrbp_1 _7518_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net444),
    .D(net1668),
    .Q_N(_0193_),
    .Q(\uart_rx_1.r_Rx_Byte[2] ));
 sg13g2_dfrbp_1 _7519_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net442),
    .D(net1630),
    .Q_N(_2970_),
    .Q(\uart_rx_1.r_Rx_Byte[3] ));
 sg13g2_dfrbp_1 _7520_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net440),
    .D(net1596),
    .Q_N(_2969_),
    .Q(\uart_rx_1.r_Rx_Byte[4] ));
 sg13g2_dfrbp_1 _7521_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net438),
    .D(net1517),
    .Q_N(_2968_),
    .Q(\uart_rx_1.r_Rx_Byte[5] ));
 sg13g2_dfrbp_1 _7522_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net436),
    .D(net1354),
    .Q_N(_2967_),
    .Q(\uart_rx_1.r_Rx_Byte[6] ));
 sg13g2_dfrbp_1 _7523_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net434),
    .D(net1421),
    .Q_N(_2966_),
    .Q(\uart_rx_1.r_Rx_Byte[7] ));
 sg13g2_dfrbp_1 _7524_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net432),
    .D(_0593_),
    .Q_N(_0205_),
    .Q(\uart_rx_1.r_Bit_Index[0] ));
 sg13g2_dfrbp_1 _7525_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net430),
    .D(_0594_),
    .Q_N(_2965_),
    .Q(\uart_rx_1.r_Bit_Index[1] ));
 sg13g2_dfrbp_1 _7526_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net428),
    .D(_0595_),
    .Q_N(_0202_),
    .Q(\uart_rx_1.r_Bit_Index[2] ));
 sg13g2_dfrbp_1 _7527_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net426),
    .D(_0596_),
    .Q_N(_2964_),
    .Q(\uart_rx_1.r_Bit_Index[3] ));
 sg13g2_dfrbp_1 _7528_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net424),
    .D(_0597_),
    .Q_N(_2963_),
    .Q(\uart_rx_1.r_Bit_Index[4] ));
 sg13g2_dfrbp_1 _7529_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net422),
    .D(_0598_),
    .Q_N(_2962_),
    .Q(\uart_rx_1.r_Bit_Index[5] ));
 sg13g2_dfrbp_1 _7530_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net144),
    .D(_0599_),
    .Q_N(_2961_),
    .Q(\uart_rx_1.r_Bit_Index[6] ));
 sg13g2_dfrbp_1 _7531_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net140),
    .D(_0600_),
    .Q_N(_2960_),
    .Q(\uart_rx_1.r_Bit_Index[7] ));
 sg13g2_dfrbp_1 _7532_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net136),
    .D(_0601_),
    .Q_N(_2959_),
    .Q(\uart_rx_1.r_Bit_Index[8] ));
 sg13g2_dfrbp_1 _7533_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net132),
    .D(_0602_),
    .Q_N(_2958_),
    .Q(\uart_rx_1.r_Bit_Index[9] ));
 sg13g2_dfrbp_1 _7534_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net128),
    .D(_0603_),
    .Q_N(_2957_),
    .Q(\uart_rx_1.r_Bit_Index[10] ));
 sg13g2_dfrbp_1 _7535_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net92),
    .D(_0604_),
    .Q_N(_2956_),
    .Q(\uart_rx_1.r_Bit_Index[11] ));
 sg13g2_dfrbp_1 _7536_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net88),
    .D(_0605_),
    .Q_N(_2955_),
    .Q(\uart_rx_1.r_Bit_Index[12] ));
 sg13g2_dfrbp_1 _7537_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net74),
    .D(_0606_),
    .Q_N(_2954_),
    .Q(\uart_rx_1.r_Bit_Index[13] ));
 sg13g2_dfrbp_1 _7538_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net70),
    .D(_0607_),
    .Q_N(_2953_),
    .Q(\uart_rx_1.r_Bit_Index[14] ));
 sg13g2_dfrbp_1 _7539_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net66),
    .D(_0608_),
    .Q_N(_2952_),
    .Q(\uart_rx_1.r_Bit_Index[15] ));
 sg13g2_dfrbp_1 _7540_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net61),
    .D(_0609_),
    .Q_N(_2951_),
    .Q(\uart_rx_1.r_Bit_Index[16] ));
 sg13g2_dfrbp_1 _7541_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net57),
    .D(_0610_),
    .Q_N(_2950_),
    .Q(\uart_rx_1.r_Bit_Index[17] ));
 sg13g2_dfrbp_1 _7542_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net53),
    .D(_0611_),
    .Q_N(_2949_),
    .Q(\uart_rx_1.r_Bit_Index[18] ));
 sg13g2_dfrbp_1 _7543_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net49),
    .D(_0612_),
    .Q_N(_2948_),
    .Q(\uart_rx_1.r_Bit_Index[19] ));
 sg13g2_dfrbp_1 _7544_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net45),
    .D(_0613_),
    .Q_N(_2947_),
    .Q(\uart_rx_1.r_Bit_Index[20] ));
 sg13g2_dfrbp_1 _7545_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net495),
    .D(_0614_),
    .Q_N(_2946_),
    .Q(\uart_rx_1.r_Bit_Index[21] ));
 sg13g2_dfrbp_1 _7546_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net491),
    .D(_0615_),
    .Q_N(_2945_),
    .Q(\uart_rx_1.r_Bit_Index[22] ));
 sg13g2_dfrbp_1 _7547_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net475),
    .D(_0616_),
    .Q_N(_2944_),
    .Q(\uart_rx_1.r_Bit_Index[23] ));
 sg13g2_dfrbp_1 _7548_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net471),
    .D(_0617_),
    .Q_N(_2943_),
    .Q(\uart_rx_1.r_Bit_Index[24] ));
 sg13g2_dfrbp_1 _7549_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net467),
    .D(_0618_),
    .Q_N(_2942_),
    .Q(\uart_rx_1.r_Bit_Index[25] ));
 sg13g2_dfrbp_1 _7550_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net463),
    .D(_0619_),
    .Q_N(_2941_),
    .Q(\uart_rx_1.r_Bit_Index[26] ));
 sg13g2_dfrbp_1 _7551_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net459),
    .D(_0620_),
    .Q_N(_2940_),
    .Q(\uart_rx_1.r_Bit_Index[27] ));
 sg13g2_dfrbp_1 _7552_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net455),
    .D(_0621_),
    .Q_N(_2939_),
    .Q(\uart_rx_1.r_Bit_Index[28] ));
 sg13g2_dfrbp_1 _7553_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net451),
    .D(_0622_),
    .Q_N(_2938_),
    .Q(\uart_rx_1.r_Bit_Index[29] ));
 sg13g2_dfrbp_1 _7554_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net447),
    .D(_0623_),
    .Q_N(_2937_),
    .Q(\uart_rx_1.r_Bit_Index[30] ));
 sg13g2_dfrbp_1 _7555_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net443),
    .D(_0624_),
    .Q_N(_2936_),
    .Q(\uart_rx_1.r_Bit_Index[31] ));
 sg13g2_dfrbp_1 _7556_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net439),
    .D(_0625_),
    .Q_N(_2935_),
    .Q(\uart_rx_1.r_Clock_Count[0] ));
 sg13g2_dfrbp_1 _7557_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net435),
    .D(_0626_),
    .Q_N(_2934_),
    .Q(\uart_rx_1.r_Clock_Count[1] ));
 sg13g2_dfrbp_1 _7558_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net431),
    .D(net1358),
    .Q_N(_2933_),
    .Q(\uart_rx_1.r_Clock_Count[2] ));
 sg13g2_dfrbp_1 _7559_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net427),
    .D(_0628_),
    .Q_N(_2932_),
    .Q(\uart_rx_1.r_Clock_Count[3] ));
 sg13g2_dfrbp_1 _7560_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net423),
    .D(_0629_),
    .Q_N(_2931_),
    .Q(\uart_rx_1.r_Clock_Count[4] ));
 sg13g2_dfrbp_1 _7561_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net142),
    .D(net1623),
    .Q_N(_0100_),
    .Q(\uart_rx_1.r_Clock_Count[5] ));
 sg13g2_dfrbp_1 _7562_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net134),
    .D(net1507),
    .Q_N(_2930_),
    .Q(\uart_rx_1.r_Clock_Count[6] ));
 sg13g2_dfrbp_1 _7563_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net126),
    .D(_0632_),
    .Q_N(_2929_),
    .Q(\uart_rx_1.r_Clock_Count[7] ));
 sg13g2_dfrbp_1 _7564_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net86),
    .D(_0633_),
    .Q_N(_2928_),
    .Q(\uart_rx_1.r_Clock_Count[8] ));
 sg13g2_dfrbp_1 _7565_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net68),
    .D(net1472),
    .Q_N(_2927_),
    .Q(\uart_rx_1.r_Clock_Count[9] ));
 sg13g2_dfrbp_1 _7566_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net59),
    .D(_0635_),
    .Q_N(_2926_),
    .Q(\uart_rx_1.r_Clock_Count[10] ));
 sg13g2_dfrbp_1 _7567_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net51),
    .D(_0636_),
    .Q_N(_2925_),
    .Q(\uart_rx_1.r_Clock_Count[11] ));
 sg13g2_dfrbp_1 _7568_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net43),
    .D(_0637_),
    .Q_N(_2924_),
    .Q(\uart_rx_1.r_Clock_Count[12] ));
 sg13g2_dfrbp_1 _7569_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net489),
    .D(net1081),
    .Q_N(_2923_),
    .Q(\uart_rx_1.r_Clock_Count[13] ));
 sg13g2_dfrbp_1 _7570_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net469),
    .D(_0639_),
    .Q_N(_2922_),
    .Q(\uart_rx_1.r_Clock_Count[14] ));
 sg13g2_dfrbp_1 _7571_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net461),
    .D(_0640_),
    .Q_N(_2921_),
    .Q(\uart_rx_1.r_Clock_Count[15] ));
 sg13g2_dfrbp_1 _7572_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net453),
    .D(_0641_),
    .Q_N(_2920_),
    .Q(\uart_rx_1.r_Clock_Count[16] ));
 sg13g2_dfrbp_1 _7573_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net445),
    .D(_0642_),
    .Q_N(_2919_),
    .Q(\uart_rx_1.r_Clock_Count[17] ));
 sg13g2_dfrbp_1 _7574_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net437),
    .D(_0643_),
    .Q_N(_2918_),
    .Q(\uart_rx_1.r_Clock_Count[18] ));
 sg13g2_dfrbp_1 _7575_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net429),
    .D(net1121),
    .Q_N(_2917_),
    .Q(\uart_rx_1.r_Clock_Count[19] ));
 sg13g2_dfrbp_1 _7576_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net146),
    .D(_0645_),
    .Q_N(_2916_),
    .Q(\uart_rx_1.r_Clock_Count[20] ));
 sg13g2_dfrbp_1 _7577_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net130),
    .D(net1068),
    .Q_N(_2915_),
    .Q(\uart_rx_1.r_Clock_Count[21] ));
 sg13g2_dfrbp_1 _7578_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net72),
    .D(_0647_),
    .Q_N(_2914_),
    .Q(\uart_rx_1.r_Clock_Count[22] ));
 sg13g2_dfrbp_1 _7579_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net55),
    .D(_0648_),
    .Q_N(_2913_),
    .Q(\uart_rx_1.r_Clock_Count[23] ));
 sg13g2_dfrbp_1 _7580_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net493),
    .D(_0649_),
    .Q_N(_2912_),
    .Q(\uart_rx_1.r_Clock_Count[24] ));
 sg13g2_dfrbp_1 _7581_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net465),
    .D(net1157),
    .Q_N(_2911_),
    .Q(\uart_rx_1.r_Clock_Count[25] ));
 sg13g2_dfrbp_1 _7582_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net449),
    .D(_0651_),
    .Q_N(_2910_),
    .Q(\uart_rx_1.r_Clock_Count[26] ));
 sg13g2_dfrbp_1 _7583_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net433),
    .D(net1143),
    .Q_N(_2909_),
    .Q(\uart_rx_1.r_Clock_Count[27] ));
 sg13g2_dfrbp_1 _7584_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net138),
    .D(_0653_),
    .Q_N(_2908_),
    .Q(\uart_rx_1.r_Clock_Count[28] ));
 sg13g2_dfrbp_1 _7585_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net63),
    .D(net1398),
    .Q_N(_2907_),
    .Q(\uart_rx_1.r_Clock_Count[29] ));
 sg13g2_dfrbp_1 _7586_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net473),
    .D(net1340),
    .Q_N(_2906_),
    .Q(\uart_rx_1.r_Clock_Count[30] ));
 sg13g2_dfrbp_1 _7587_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net441),
    .D(net1076),
    .Q_N(_2905_),
    .Q(\uart_rx_1.r_Clock_Count[31] ));
 sg13g2_dfrbp_1 _7588_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net90),
    .D(_0657_),
    .Q_N(_2904_),
    .Q(\uart_rx_1.r_SM_Main[0] ));
 sg13g2_dfrbp_1 _7589_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net457),
    .D(net1663),
    .Q_N(_2903_),
    .Q(\uart_rx_1.r_SM_Main[1] ));
 sg13g2_dfrbp_1 _7590_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net47),
    .D(net1409),
    .Q_N(_0099_),
    .Q(\uart_rx_1.r_SM_Main[2] ));
 sg13g2_tiehi _6927__26 (.L_HI(net26));
 sg13g2_tiehi _6924__27 (.L_HI(net27));
 sg13g2_tiehi _6925__28 (.L_HI(net28));
 sg13g2_tiehi _7289__29 (.L_HI(net29));
 sg13g2_tiehi _7288__30 (.L_HI(net30));
 sg13g2_tiehi _7287__31 (.L_HI(net31));
 sg13g2_tiehi _7286__32 (.L_HI(net32));
 sg13g2_tiehi _7285__33 (.L_HI(net33));
 sg13g2_tiehi _7284__34 (.L_HI(net34));
 sg13g2_tiehi _7283__35 (.L_HI(net35));
 sg13g2_tiehi _7282__36 (.L_HI(net36));
 sg13g2_tiehi _7281__37 (.L_HI(net37));
 sg13g2_tiehi _7280__38 (.L_HI(net38));
 sg13g2_tiehi _7279__39 (.L_HI(net39));
 sg13g2_tiehi _7278__40 (.L_HI(net40));
 sg13g2_tiehi _7277__41 (.L_HI(net41));
 sg13g2_tiehi _7276__42 (.L_HI(net42));
 sg13g2_tiehi _7568__43 (.L_HI(net43));
 sg13g2_tiehi _7275__44 (.L_HI(net44));
 sg13g2_tiehi _7544__45 (.L_HI(net45));
 sg13g2_tiehi _7184__46 (.L_HI(net46));
 sg13g2_tiehi _7590__47 (.L_HI(net47));
 sg13g2_tiehi _7164__48 (.L_HI(net48));
 sg13g2_tiehi _7543__49 (.L_HI(net49));
 sg13g2_tiehi _7163__50 (.L_HI(net50));
 sg13g2_tiehi _7567__51 (.L_HI(net51));
 sg13g2_tiehi _7162__52 (.L_HI(net52));
 sg13g2_tiehi _7542__53 (.L_HI(net53));
 sg13g2_tiehi _7161__54 (.L_HI(net54));
 sg13g2_tiehi _7579__55 (.L_HI(net55));
 sg13g2_tiehi _7160__56 (.L_HI(net56));
 sg13g2_tiehi _7541__57 (.L_HI(net57));
 sg13g2_tiehi _7159__58 (.L_HI(net58));
 sg13g2_tiehi _7566__59 (.L_HI(net59));
 sg13g2_tiehi _7158__60 (.L_HI(net60));
 sg13g2_tiehi _7540__61 (.L_HI(net61));
 sg13g2_tiehi _7157__62 (.L_HI(net62));
 sg13g2_tiehi _7585__63 (.L_HI(net63));
 sg13g2_tiehi _7140__64 (.L_HI(net64));
 sg13g2_tiehi _7139__65 (.L_HI(net65));
 sg13g2_tiehi _7539__66 (.L_HI(net66));
 sg13g2_tiehi _7134__67 (.L_HI(net67));
 sg13g2_tiehi _7565__68 (.L_HI(net68));
 sg13g2_tiehi _7125__69 (.L_HI(net69));
 sg13g2_tiehi _7538__70 (.L_HI(net70));
 sg13g2_tiehi _7068__71 (.L_HI(net71));
 sg13g2_tiehi _7578__72 (.L_HI(net72));
 sg13g2_tiehi _7067__73 (.L_HI(net73));
 sg13g2_tiehi _7537__74 (.L_HI(net74));
 sg13g2_tiehi _7066__75 (.L_HI(net75));
 sg13g2_tiehi _7065__76 (.L_HI(net76));
 sg13g2_tiehi _7064__77 (.L_HI(net77));
 sg13g2_tiehi _7063__78 (.L_HI(net78));
 sg13g2_tiehi _7062__79 (.L_HI(net79));
 sg13g2_tiehi _7061__80 (.L_HI(net80));
 sg13g2_tiehi _7060__81 (.L_HI(net81));
 sg13g2_tiehi _7059__82 (.L_HI(net82));
 sg13g2_tiehi _7058__83 (.L_HI(net83));
 sg13g2_tiehi _7057__84 (.L_HI(net84));
 sg13g2_tiehi _7056__85 (.L_HI(net85));
 sg13g2_tiehi _7564__86 (.L_HI(net86));
 sg13g2_tiehi _7055__87 (.L_HI(net87));
 sg13g2_tiehi _7536__88 (.L_HI(net88));
 sg13g2_tiehi _7053__89 (.L_HI(net89));
 sg13g2_tiehi _7588__90 (.L_HI(net90));
 sg13g2_tiehi _7052__91 (.L_HI(net91));
 sg13g2_tiehi _7535__92 (.L_HI(net92));
 sg13g2_tiehi _7051__93 (.L_HI(net93));
 sg13g2_tiehi _7050__94 (.L_HI(net94));
 sg13g2_tiehi _7049__95 (.L_HI(net95));
 sg13g2_tiehi _7048__96 (.L_HI(net96));
 sg13g2_tiehi _7047__97 (.L_HI(net97));
 sg13g2_tiehi _7046__98 (.L_HI(net98));
 sg13g2_tiehi _7045__99 (.L_HI(net99));
 sg13g2_tiehi _7044__100 (.L_HI(net100));
 sg13g2_tiehi _6926__101 (.L_HI(net101));
 sg13g2_tiehi _6999__102 (.L_HI(net102));
 sg13g2_tiehi _7000__103 (.L_HI(net103));
 sg13g2_tiehi _7001__104 (.L_HI(net104));
 sg13g2_tiehi _7002__105 (.L_HI(net105));
 sg13g2_tiehi _7003__106 (.L_HI(net106));
 sg13g2_tiehi _7004__107 (.L_HI(net107));
 sg13g2_tiehi _7005__108 (.L_HI(net108));
 sg13g2_tiehi _7043__109 (.L_HI(net109));
 sg13g2_tiehi _7042__110 (.L_HI(net110));
 sg13g2_tiehi _7041__111 (.L_HI(net111));
 sg13g2_tiehi _7040__112 (.L_HI(net112));
 sg13g2_tiehi _7039__113 (.L_HI(net113));
 sg13g2_tiehi _7038__114 (.L_HI(net114));
 sg13g2_tiehi _7037__115 (.L_HI(net115));
 sg13g2_tiehi _7036__116 (.L_HI(net116));
 sg13g2_tiehi _7035__117 (.L_HI(net117));
 sg13g2_tiehi _7034__118 (.L_HI(net118));
 sg13g2_tiehi _7033__119 (.L_HI(net119));
 sg13g2_tiehi _7032__120 (.L_HI(net120));
 sg13g2_tiehi _7031__121 (.L_HI(net121));
 sg13g2_tiehi _7030__122 (.L_HI(net122));
 sg13g2_tiehi _7029__123 (.L_HI(net123));
 sg13g2_tiehi _7028__124 (.L_HI(net124));
 sg13g2_tiehi _7027__125 (.L_HI(net125));
 sg13g2_tiehi _7563__126 (.L_HI(net126));
 sg13g2_tiehi _7026__127 (.L_HI(net127));
 sg13g2_tiehi _7534__128 (.L_HI(net128));
 sg13g2_tiehi _7025__129 (.L_HI(net129));
 sg13g2_tiehi _7577__130 (.L_HI(net130));
 sg13g2_tiehi _7024__131 (.L_HI(net131));
 sg13g2_tiehi _7533__132 (.L_HI(net132));
 sg13g2_tiehi _7023__133 (.L_HI(net133));
 sg13g2_tiehi _7562__134 (.L_HI(net134));
 sg13g2_tiehi _7022__135 (.L_HI(net135));
 sg13g2_tiehi _7532__136 (.L_HI(net136));
 sg13g2_tiehi _7021__137 (.L_HI(net137));
 sg13g2_tiehi _7584__138 (.L_HI(net138));
 sg13g2_tiehi _7020__139 (.L_HI(net139));
 sg13g2_tiehi _7531__140 (.L_HI(net140));
 sg13g2_tiehi _7019__141 (.L_HI(net141));
 sg13g2_tiehi _7561__142 (.L_HI(net142));
 sg13g2_tiehi _7018__143 (.L_HI(net143));
 sg13g2_tiehi _7530__144 (.L_HI(net144));
 sg13g2_tiehi _7017__145 (.L_HI(net145));
 sg13g2_tiehi _7576__146 (.L_HI(net146));
 sg13g2_tiehi _7016__147 (.L_HI(net147));
 sg13g2_tiehi _7015__148 (.L_HI(net148));
 sg13g2_tiehi _7014__149 (.L_HI(net149));
 sg13g2_tiehi _7013__150 (.L_HI(net150));
 sg13g2_tiehi _7012__151 (.L_HI(net151));
 sg13g2_tiehi _7011__152 (.L_HI(net152));
 sg13g2_tiehi _7010__153 (.L_HI(net153));
 sg13g2_tiehi _7009__154 (.L_HI(net154));
 sg13g2_tiehi _7008__155 (.L_HI(net155));
 sg13g2_tiehi _7006__156 (.L_HI(net156));
 sg13g2_tiehi _7007__157 (.L_HI(net157));
 sg13g2_tiehi _6998__158 (.L_HI(net158));
 sg13g2_tiehi _6997__159 (.L_HI(net159));
 sg13g2_tiehi _6996__160 (.L_HI(net160));
 sg13g2_tiehi _6995__161 (.L_HI(net161));
 sg13g2_tiehi _6994__162 (.L_HI(net162));
 sg13g2_tiehi _6993__163 (.L_HI(net163));
 sg13g2_tiehi _6992__164 (.L_HI(net164));
 sg13g2_tiehi _6991__165 (.L_HI(net165));
 sg13g2_tiehi _6990__166 (.L_HI(net166));
 sg13g2_tiehi _6989__167 (.L_HI(net167));
 sg13g2_tiehi _6988__168 (.L_HI(net168));
 sg13g2_tiehi _6987__169 (.L_HI(net169));
 sg13g2_tiehi _6986__170 (.L_HI(net170));
 sg13g2_tiehi _7054__171 (.L_HI(net171));
 sg13g2_tiehi _7069__172 (.L_HI(net172));
 sg13g2_tiehi _7070__173 (.L_HI(net173));
 sg13g2_tiehi _7071__174 (.L_HI(net174));
 sg13g2_tiehi _7072__175 (.L_HI(net175));
 sg13g2_tiehi _7073__176 (.L_HI(net176));
 sg13g2_tiehi _7074__177 (.L_HI(net177));
 sg13g2_tiehi _7075__178 (.L_HI(net178));
 sg13g2_tiehi _7076__179 (.L_HI(net179));
 sg13g2_tiehi _7077__180 (.L_HI(net180));
 sg13g2_tiehi _7078__181 (.L_HI(net181));
 sg13g2_tiehi _7079__182 (.L_HI(net182));
 sg13g2_tiehi _7080__183 (.L_HI(net183));
 sg13g2_tiehi _7081__184 (.L_HI(net184));
 sg13g2_tiehi _7082__185 (.L_HI(net185));
 sg13g2_tiehi _7083__186 (.L_HI(net186));
 sg13g2_tiehi _7084__187 (.L_HI(net187));
 sg13g2_tiehi _7085__188 (.L_HI(net188));
 sg13g2_tiehi _7086__189 (.L_HI(net189));
 sg13g2_tiehi _7087__190 (.L_HI(net190));
 sg13g2_tiehi _7088__191 (.L_HI(net191));
 sg13g2_tiehi _7089__192 (.L_HI(net192));
 sg13g2_tiehi _7090__193 (.L_HI(net193));
 sg13g2_tiehi _7091__194 (.L_HI(net194));
 sg13g2_tiehi _7092__195 (.L_HI(net195));
 sg13g2_tiehi _7093__196 (.L_HI(net196));
 sg13g2_tiehi _7094__197 (.L_HI(net197));
 sg13g2_tiehi _7095__198 (.L_HI(net198));
 sg13g2_tiehi _7096__199 (.L_HI(net199));
 sg13g2_tiehi _7097__200 (.L_HI(net200));
 sg13g2_tiehi _7098__201 (.L_HI(net201));
 sg13g2_tiehi _7099__202 (.L_HI(net202));
 sg13g2_tiehi _7100__203 (.L_HI(net203));
 sg13g2_tiehi _7101__204 (.L_HI(net204));
 sg13g2_tiehi _7102__205 (.L_HI(net205));
 sg13g2_tiehi _7103__206 (.L_HI(net206));
 sg13g2_tiehi _7104__207 (.L_HI(net207));
 sg13g2_tiehi _7105__208 (.L_HI(net208));
 sg13g2_tiehi _7106__209 (.L_HI(net209));
 sg13g2_tiehi _7107__210 (.L_HI(net210));
 sg13g2_tiehi _7108__211 (.L_HI(net211));
 sg13g2_tiehi _7109__212 (.L_HI(net212));
 sg13g2_tiehi _7110__213 (.L_HI(net213));
 sg13g2_tiehi _7111__214 (.L_HI(net214));
 sg13g2_tiehi _7112__215 (.L_HI(net215));
 sg13g2_tiehi _7113__216 (.L_HI(net216));
 sg13g2_tiehi _7114__217 (.L_HI(net217));
 sg13g2_tiehi _7115__218 (.L_HI(net218));
 sg13g2_tiehi _7116__219 (.L_HI(net219));
 sg13g2_tiehi _7117__220 (.L_HI(net220));
 sg13g2_tiehi _7118__221 (.L_HI(net221));
 sg13g2_tiehi _7119__222 (.L_HI(net222));
 sg13g2_tiehi _7120__223 (.L_HI(net223));
 sg13g2_tiehi _7121__224 (.L_HI(net224));
 sg13g2_tiehi _7122__225 (.L_HI(net225));
 sg13g2_tiehi _7123__226 (.L_HI(net226));
 sg13g2_tiehi _6985__227 (.L_HI(net227));
 sg13g2_tiehi _7124__228 (.L_HI(net228));
 sg13g2_tiehi _7126__229 (.L_HI(net229));
 sg13g2_tiehi _7127__230 (.L_HI(net230));
 sg13g2_tiehi _7128__231 (.L_HI(net231));
 sg13g2_tiehi _7129__232 (.L_HI(net232));
 sg13g2_tiehi _7130__233 (.L_HI(net233));
 sg13g2_tiehi _7131__234 (.L_HI(net234));
 sg13g2_tiehi _7132__235 (.L_HI(net235));
 sg13g2_tiehi _6984__236 (.L_HI(net236));
 sg13g2_tiehi _7133__237 (.L_HI(net237));
 sg13g2_tiehi _7135__238 (.L_HI(net238));
 sg13g2_tiehi _7136__239 (.L_HI(net239));
 sg13g2_tiehi _7137__240 (.L_HI(net240));
 sg13g2_tiehi _6983__241 (.L_HI(net241));
 sg13g2_tiehi _6982__242 (.L_HI(net242));
 sg13g2_tiehi _7138__243 (.L_HI(net243));
 sg13g2_tiehi _7141__244 (.L_HI(net244));
 sg13g2_tiehi _7142__245 (.L_HI(net245));
 sg13g2_tiehi _7143__246 (.L_HI(net246));
 sg13g2_tiehi _7144__247 (.L_HI(net247));
 sg13g2_tiehi _7145__248 (.L_HI(net248));
 sg13g2_tiehi _7146__249 (.L_HI(net249));
 sg13g2_tiehi _7147__250 (.L_HI(net250));
 sg13g2_tiehi _7148__251 (.L_HI(net251));
 sg13g2_tiehi _7149__252 (.L_HI(net252));
 sg13g2_tiehi _7150__253 (.L_HI(net253));
 sg13g2_tiehi _7151__254 (.L_HI(net254));
 sg13g2_tiehi _7152__255 (.L_HI(net255));
 sg13g2_tiehi _7153__256 (.L_HI(net256));
 sg13g2_tiehi _7154__257 (.L_HI(net257));
 sg13g2_tiehi _7155__258 (.L_HI(net258));
 sg13g2_tiehi _6981__259 (.L_HI(net259));
 sg13g2_tiehi _6980__260 (.L_HI(net260));
 sg13g2_tiehi _6979__261 (.L_HI(net261));
 sg13g2_tiehi _6978__262 (.L_HI(net262));
 sg13g2_tiehi _6977__263 (.L_HI(net263));
 sg13g2_tiehi _6976__264 (.L_HI(net264));
 sg13g2_tiehi _6975__265 (.L_HI(net265));
 sg13g2_tiehi _6974__266 (.L_HI(net266));
 sg13g2_tiehi _7156__267 (.L_HI(net267));
 sg13g2_tiehi _7165__268 (.L_HI(net268));
 sg13g2_tiehi _7166__269 (.L_HI(net269));
 sg13g2_tiehi _7167__270 (.L_HI(net270));
 sg13g2_tiehi _7168__271 (.L_HI(net271));
 sg13g2_tiehi _7169__272 (.L_HI(net272));
 sg13g2_tiehi _7170__273 (.L_HI(net273));
 sg13g2_tiehi _7171__274 (.L_HI(net274));
 sg13g2_tiehi _7172__275 (.L_HI(net275));
 sg13g2_tiehi _7173__276 (.L_HI(net276));
 sg13g2_tiehi _7174__277 (.L_HI(net277));
 sg13g2_tiehi _7175__278 (.L_HI(net278));
 sg13g2_tiehi _7176__279 (.L_HI(net279));
 sg13g2_tiehi _7177__280 (.L_HI(net280));
 sg13g2_tiehi _7178__281 (.L_HI(net281));
 sg13g2_tiehi _7179__282 (.L_HI(net282));
 sg13g2_tiehi _7180__283 (.L_HI(net283));
 sg13g2_tiehi _7181__284 (.L_HI(net284));
 sg13g2_tiehi _7182__285 (.L_HI(net285));
 sg13g2_tiehi _6973__286 (.L_HI(net286));
 sg13g2_tiehi _7183__287 (.L_HI(net287));
 sg13g2_tiehi _7185__288 (.L_HI(net288));
 sg13g2_tiehi _7186__289 (.L_HI(net289));
 sg13g2_tiehi _7187__290 (.L_HI(net290));
 sg13g2_tiehi _7188__291 (.L_HI(net291));
 sg13g2_tiehi _7189__292 (.L_HI(net292));
 sg13g2_tiehi _7190__293 (.L_HI(net293));
 sg13g2_tiehi _7191__294 (.L_HI(net294));
 sg13g2_tiehi _7192__295 (.L_HI(net295));
 sg13g2_tiehi _7193__296 (.L_HI(net296));
 sg13g2_tiehi _7194__297 (.L_HI(net297));
 sg13g2_tiehi _7195__298 (.L_HI(net298));
 sg13g2_tiehi _7196__299 (.L_HI(net299));
 sg13g2_tiehi _7197__300 (.L_HI(net300));
 sg13g2_tiehi _7198__301 (.L_HI(net301));
 sg13g2_tiehi _7199__302 (.L_HI(net302));
 sg13g2_tiehi _7200__303 (.L_HI(net303));
 sg13g2_tiehi _7201__304 (.L_HI(net304));
 sg13g2_tiehi _7202__305 (.L_HI(net305));
 sg13g2_tiehi _7203__306 (.L_HI(net306));
 sg13g2_tiehi _7204__307 (.L_HI(net307));
 sg13g2_tiehi _7205__308 (.L_HI(net308));
 sg13g2_tiehi _7206__309 (.L_HI(net309));
 sg13g2_tiehi _7207__310 (.L_HI(net310));
 sg13g2_tiehi _7208__311 (.L_HI(net311));
 sg13g2_tiehi _7209__312 (.L_HI(net312));
 sg13g2_tiehi _7210__313 (.L_HI(net313));
 sg13g2_tiehi _7211__314 (.L_HI(net314));
 sg13g2_tiehi _7212__315 (.L_HI(net315));
 sg13g2_tiehi _7213__316 (.L_HI(net316));
 sg13g2_tiehi _7214__317 (.L_HI(net317));
 sg13g2_tiehi _7215__318 (.L_HI(net318));
 sg13g2_tiehi _7216__319 (.L_HI(net319));
 sg13g2_tiehi _7217__320 (.L_HI(net320));
 sg13g2_tiehi _7218__321 (.L_HI(net321));
 sg13g2_tiehi _7219__322 (.L_HI(net322));
 sg13g2_tiehi _7220__323 (.L_HI(net323));
 sg13g2_tiehi _7221__324 (.L_HI(net324));
 sg13g2_tiehi _7222__325 (.L_HI(net325));
 sg13g2_tiehi _7223__326 (.L_HI(net326));
 sg13g2_tiehi _7224__327 (.L_HI(net327));
 sg13g2_tiehi _7225__328 (.L_HI(net328));
 sg13g2_tiehi _7226__329 (.L_HI(net329));
 sg13g2_tiehi _7227__330 (.L_HI(net330));
 sg13g2_tiehi _7228__331 (.L_HI(net331));
 sg13g2_tiehi _7229__332 (.L_HI(net332));
 sg13g2_tiehi _7230__333 (.L_HI(net333));
 sg13g2_tiehi _7231__334 (.L_HI(net334));
 sg13g2_tiehi _7232__335 (.L_HI(net335));
 sg13g2_tiehi _7233__336 (.L_HI(net336));
 sg13g2_tiehi _7234__337 (.L_HI(net337));
 sg13g2_tiehi _7235__338 (.L_HI(net338));
 sg13g2_tiehi _7236__339 (.L_HI(net339));
 sg13g2_tiehi _7237__340 (.L_HI(net340));
 sg13g2_tiehi _7238__341 (.L_HI(net341));
 sg13g2_tiehi _7239__342 (.L_HI(net342));
 sg13g2_tiehi _7240__343 (.L_HI(net343));
 sg13g2_tiehi _7241__344 (.L_HI(net344));
 sg13g2_tiehi _7242__345 (.L_HI(net345));
 sg13g2_tiehi _7243__346 (.L_HI(net346));
 sg13g2_tiehi _7244__347 (.L_HI(net347));
 sg13g2_tiehi _7245__348 (.L_HI(net348));
 sg13g2_tiehi _7246__349 (.L_HI(net349));
 sg13g2_tiehi _7247__350 (.L_HI(net350));
 sg13g2_tiehi _7248__351 (.L_HI(net351));
 sg13g2_tiehi _7249__352 (.L_HI(net352));
 sg13g2_tiehi _7250__353 (.L_HI(net353));
 sg13g2_tiehi _7251__354 (.L_HI(net354));
 sg13g2_tiehi _7252__355 (.L_HI(net355));
 sg13g2_tiehi _7253__356 (.L_HI(net356));
 sg13g2_tiehi _7254__357 (.L_HI(net357));
 sg13g2_tiehi _7255__358 (.L_HI(net358));
 sg13g2_tiehi _7256__359 (.L_HI(net359));
 sg13g2_tiehi _7257__360 (.L_HI(net360));
 sg13g2_tiehi _7258__361 (.L_HI(net361));
 sg13g2_tiehi _7259__362 (.L_HI(net362));
 sg13g2_tiehi _7260__363 (.L_HI(net363));
 sg13g2_tiehi _7261__364 (.L_HI(net364));
 sg13g2_tiehi _7262__365 (.L_HI(net365));
 sg13g2_tiehi _7263__366 (.L_HI(net366));
 sg13g2_tiehi _7264__367 (.L_HI(net367));
 sg13g2_tiehi _7265__368 (.L_HI(net368));
 sg13g2_tiehi _7266__369 (.L_HI(net369));
 sg13g2_tiehi _7267__370 (.L_HI(net370));
 sg13g2_tiehi _7268__371 (.L_HI(net371));
 sg13g2_tiehi _7269__372 (.L_HI(net372));
 sg13g2_tiehi _7270__373 (.L_HI(net373));
 sg13g2_tiehi _7271__374 (.L_HI(net374));
 sg13g2_tiehi _7272__375 (.L_HI(net375));
 sg13g2_tiehi _7273__376 (.L_HI(net376));
 sg13g2_tiehi _6972__377 (.L_HI(net377));
 sg13g2_tiehi _6971__378 (.L_HI(net378));
 sg13g2_tiehi _6970__379 (.L_HI(net379));
 sg13g2_tiehi _6969__380 (.L_HI(net380));
 sg13g2_tiehi _6968__381 (.L_HI(net381));
 sg13g2_tiehi _6967__382 (.L_HI(net382));
 sg13g2_tiehi _6966__383 (.L_HI(net383));
 sg13g2_tiehi _6965__384 (.L_HI(net384));
 sg13g2_tiehi _6964__385 (.L_HI(net385));
 sg13g2_tiehi _6963__386 (.L_HI(net386));
 sg13g2_tiehi _6962__387 (.L_HI(net387));
 sg13g2_tiehi _6961__388 (.L_HI(net388));
 sg13g2_tiehi _6960__389 (.L_HI(net389));
 sg13g2_tiehi _6959__390 (.L_HI(net390));
 sg13g2_tiehi _6958__391 (.L_HI(net391));
 sg13g2_tiehi _6957__392 (.L_HI(net392));
 sg13g2_tiehi _6956__393 (.L_HI(net393));
 sg13g2_tiehi _6955__394 (.L_HI(net394));
 sg13g2_tiehi _6954__395 (.L_HI(net395));
 sg13g2_tiehi _6953__396 (.L_HI(net396));
 sg13g2_tiehi _6952__397 (.L_HI(net397));
 sg13g2_tiehi _6951__398 (.L_HI(net398));
 sg13g2_tiehi _6950__399 (.L_HI(net399));
 sg13g2_tiehi _6949__400 (.L_HI(net400));
 sg13g2_tiehi _6948__401 (.L_HI(net401));
 sg13g2_tiehi _6947__402 (.L_HI(net402));
 sg13g2_tiehi _6946__403 (.L_HI(net403));
 sg13g2_tiehi _6945__404 (.L_HI(net404));
 sg13g2_tiehi _6944__405 (.L_HI(net405));
 sg13g2_tiehi _6943__406 (.L_HI(net406));
 sg13g2_tiehi _6942__407 (.L_HI(net407));
 sg13g2_tiehi _6941__408 (.L_HI(net408));
 sg13g2_tiehi _6940__409 (.L_HI(net409));
 sg13g2_tiehi _6939__410 (.L_HI(net410));
 sg13g2_tiehi _6938__411 (.L_HI(net411));
 sg13g2_tiehi _6937__412 (.L_HI(net412));
 sg13g2_tiehi _6936__413 (.L_HI(net413));
 sg13g2_tiehi _6935__414 (.L_HI(net414));
 sg13g2_tiehi _6934__415 (.L_HI(net415));
 sg13g2_tiehi _6933__416 (.L_HI(net416));
 sg13g2_tiehi _6932__417 (.L_HI(net417));
 sg13g2_tiehi _6931__418 (.L_HI(net418));
 sg13g2_tiehi _6930__419 (.L_HI(net419));
 sg13g2_tiehi _6929__420 (.L_HI(net420));
 sg13g2_tiehi _6928__421 (.L_HI(net421));
 sg13g2_tiehi _7529__422 (.L_HI(net422));
 sg13g2_tiehi _7560__423 (.L_HI(net423));
 sg13g2_tiehi _7528__424 (.L_HI(net424));
 sg13g2_tiehi _7513__425 (.L_HI(net425));
 sg13g2_tiehi _7527__426 (.L_HI(net426));
 sg13g2_tiehi _7559__427 (.L_HI(net427));
 sg13g2_tiehi _7526__428 (.L_HI(net428));
 sg13g2_tiehi _7575__429 (.L_HI(net429));
 sg13g2_tiehi _7525__430 (.L_HI(net430));
 sg13g2_tiehi _7558__431 (.L_HI(net431));
 sg13g2_tiehi _7524__432 (.L_HI(net432));
 sg13g2_tiehi _7583__433 (.L_HI(net433));
 sg13g2_tiehi _7523__434 (.L_HI(net434));
 sg13g2_tiehi _7557__435 (.L_HI(net435));
 sg13g2_tiehi _7522__436 (.L_HI(net436));
 sg13g2_tiehi _7574__437 (.L_HI(net437));
 sg13g2_tiehi _7521__438 (.L_HI(net438));
 sg13g2_tiehi _7556__439 (.L_HI(net439));
 sg13g2_tiehi _7520__440 (.L_HI(net440));
 sg13g2_tiehi _7587__441 (.L_HI(net441));
 sg13g2_tiehi _7519__442 (.L_HI(net442));
 sg13g2_tiehi _7555__443 (.L_HI(net443));
 sg13g2_tiehi _7518__444 (.L_HI(net444));
 sg13g2_tiehi _7573__445 (.L_HI(net445));
 sg13g2_tiehi _7517__446 (.L_HI(net446));
 sg13g2_tiehi _7554__447 (.L_HI(net447));
 sg13g2_tiehi _7516__448 (.L_HI(net448));
 sg13g2_tiehi _7582__449 (.L_HI(net449));
 sg13g2_tiehi _7515__450 (.L_HI(net450));
 sg13g2_tiehi _7553__451 (.L_HI(net451));
 sg13g2_tiehi _7514__452 (.L_HI(net452));
 sg13g2_tiehi _7572__453 (.L_HI(net453));
 sg13g2_tiehi _7511__454 (.L_HI(net454));
 sg13g2_tiehi _7552__455 (.L_HI(net455));
 sg13g2_tiehi _7510__456 (.L_HI(net456));
 sg13g2_tiehi _7589__457 (.L_HI(net457));
 sg13g2_tiehi _7509__458 (.L_HI(net458));
 sg13g2_tiehi _7551__459 (.L_HI(net459));
 sg13g2_tiehi _7508__460 (.L_HI(net460));
 sg13g2_tiehi _7571__461 (.L_HI(net461));
 sg13g2_tiehi _7507__462 (.L_HI(net462));
 sg13g2_tiehi _7550__463 (.L_HI(net463));
 sg13g2_tiehi _7506__464 (.L_HI(net464));
 sg13g2_tiehi _7581__465 (.L_HI(net465));
 sg13g2_tiehi _7505__466 (.L_HI(net466));
 sg13g2_tiehi _7549__467 (.L_HI(net467));
 sg13g2_tiehi _7504__468 (.L_HI(net468));
 sg13g2_tiehi _7570__469 (.L_HI(net469));
 sg13g2_tiehi _7503__470 (.L_HI(net470));
 sg13g2_tiehi _7548__471 (.L_HI(net471));
 sg13g2_tiehi _7502__472 (.L_HI(net472));
 sg13g2_tiehi _7586__473 (.L_HI(net473));
 sg13g2_tiehi _7501__474 (.L_HI(net474));
 sg13g2_tiehi _7547__475 (.L_HI(net475));
 sg13g2_tiehi _7500__476 (.L_HI(net476));
 sg13g2_tiehi _7499__477 (.L_HI(net477));
 sg13g2_tiehi _7498__478 (.L_HI(net478));
 sg13g2_tiehi _7497__479 (.L_HI(net479));
 sg13g2_tiehi _7496__480 (.L_HI(net480));
 sg13g2_tiehi _7495__481 (.L_HI(net481));
 sg13g2_tiehi _7494__482 (.L_HI(net482));
 sg13g2_tiehi _7493__483 (.L_HI(net483));
 sg13g2_tiehi _7492__484 (.L_HI(net484));
 sg13g2_tiehi _7491__485 (.L_HI(net485));
 sg13g2_tiehi _7490__486 (.L_HI(net486));
 sg13g2_tiehi _7489__487 (.L_HI(net487));
 sg13g2_tiehi _7488__488 (.L_HI(net488));
 sg13g2_tiehi _7569__489 (.L_HI(net489));
 sg13g2_tiehi _7487__490 (.L_HI(net490));
 sg13g2_tiehi _7546__491 (.L_HI(net491));
 sg13g2_tiehi _7486__492 (.L_HI(net492));
 sg13g2_tiehi _7580__493 (.L_HI(net493));
 sg13g2_tiehi _7485__494 (.L_HI(net494));
 sg13g2_tiehi _7545__495 (.L_HI(net495));
 sg13g2_tiehi _7484__496 (.L_HI(net496));
 sg13g2_tiehi _7483__497 (.L_HI(net497));
 sg13g2_tiehi _7482__498 (.L_HI(net498));
 sg13g2_tiehi _7481__499 (.L_HI(net499));
 sg13g2_tiehi _7480__500 (.L_HI(net500));
 sg13g2_tiehi _7479__501 (.L_HI(net501));
 sg13g2_tiehi _7478__502 (.L_HI(net502));
 sg13g2_tiehi _7477__503 (.L_HI(net503));
 sg13g2_tiehi _7476__504 (.L_HI(net504));
 sg13g2_tiehi _7475__505 (.L_HI(net505));
 sg13g2_tiehi _7474__506 (.L_HI(net506));
 sg13g2_tiehi _7473__507 (.L_HI(net507));
 sg13g2_tiehi _7472__508 (.L_HI(net508));
 sg13g2_tiehi _7471__509 (.L_HI(net509));
 sg13g2_tiehi _7470__510 (.L_HI(net510));
 sg13g2_tiehi _7469__511 (.L_HI(net511));
 sg13g2_tiehi _7468__512 (.L_HI(net512));
 sg13g2_tiehi _7467__513 (.L_HI(net513));
 sg13g2_tiehi _7466__514 (.L_HI(net514));
 sg13g2_tiehi _7465__515 (.L_HI(net515));
 sg13g2_tiehi _7464__516 (.L_HI(net516));
 sg13g2_tiehi _7463__517 (.L_HI(net517));
 sg13g2_tiehi _7462__518 (.L_HI(net518));
 sg13g2_tiehi _7461__519 (.L_HI(net519));
 sg13g2_tiehi _7460__520 (.L_HI(net520));
 sg13g2_tiehi _7459__521 (.L_HI(net521));
 sg13g2_tiehi _7458__522 (.L_HI(net522));
 sg13g2_tiehi _7457__523 (.L_HI(net523));
 sg13g2_tiehi _7456__524 (.L_HI(net524));
 sg13g2_tiehi _7455__525 (.L_HI(net525));
 sg13g2_tiehi _7454__526 (.L_HI(net526));
 sg13g2_tiehi _7453__527 (.L_HI(net527));
 sg13g2_tiehi _7452__528 (.L_HI(net528));
 sg13g2_tiehi _7451__529 (.L_HI(net529));
 sg13g2_tiehi _7450__530 (.L_HI(net530));
 sg13g2_tiehi _7440__531 (.L_HI(net531));
 sg13g2_tiehi _7439__532 (.L_HI(net532));
 sg13g2_tiehi _7438__533 (.L_HI(net533));
 sg13g2_tiehi _7437__534 (.L_HI(net534));
 sg13g2_tiehi _7436__535 (.L_HI(net535));
 sg13g2_tiehi _7435__536 (.L_HI(net536));
 sg13g2_tiehi _7434__537 (.L_HI(net537));
 sg13g2_tiehi _7433__538 (.L_HI(net538));
 sg13g2_tiehi _7432__539 (.L_HI(net539));
 sg13g2_tiehi _7431__540 (.L_HI(net540));
 sg13g2_tiehi _7430__541 (.L_HI(net541));
 sg13g2_tiehi _7429__542 (.L_HI(net542));
 sg13g2_tiehi _7274__543 (.L_HI(net543));
 sg13g2_tiehi _7441__544 (.L_HI(net544));
 sg13g2_tiehi _7442__545 (.L_HI(net545));
 sg13g2_tiehi _7443__546 (.L_HI(net546));
 sg13g2_tiehi _7444__547 (.L_HI(net547));
 sg13g2_tiehi _7445__548 (.L_HI(net548));
 sg13g2_tiehi _7446__549 (.L_HI(net549));
 sg13g2_tiehi _7447__550 (.L_HI(net550));
 sg13g2_tiehi _7448__551 (.L_HI(net551));
 sg13g2_tiehi _7428__552 (.L_HI(net552));
 sg13g2_tiehi _7427__553 (.L_HI(net553));
 sg13g2_tiehi _7426__554 (.L_HI(net554));
 sg13g2_tiehi _7425__555 (.L_HI(net555));
 sg13g2_tiehi _7424__556 (.L_HI(net556));
 sg13g2_tiehi _7423__557 (.L_HI(net557));
 sg13g2_tiehi _7422__558 (.L_HI(net558));
 sg13g2_tiehi _7421__559 (.L_HI(net559));
 sg13g2_tiehi _7420__560 (.L_HI(net560));
 sg13g2_tiehi _7419__561 (.L_HI(net561));
 sg13g2_tiehi _7418__562 (.L_HI(net562));
 sg13g2_tiehi _7417__563 (.L_HI(net563));
 sg13g2_tiehi _7416__564 (.L_HI(net564));
 sg13g2_tiehi _7415__565 (.L_HI(net565));
 sg13g2_tiehi _7414__566 (.L_HI(net566));
 sg13g2_tiehi _7413__567 (.L_HI(net567));
 sg13g2_tiehi _7412__568 (.L_HI(net568));
 sg13g2_tiehi _7411__569 (.L_HI(net569));
 sg13g2_tiehi _7410__570 (.L_HI(net570));
 sg13g2_tiehi _7409__571 (.L_HI(net571));
 sg13g2_tiehi _7408__572 (.L_HI(net572));
 sg13g2_tiehi _7407__573 (.L_HI(net573));
 sg13g2_tiehi _7406__574 (.L_HI(net574));
 sg13g2_tiehi _7405__575 (.L_HI(net575));
 sg13g2_tiehi _7404__576 (.L_HI(net576));
 sg13g2_tiehi _7403__577 (.L_HI(net577));
 sg13g2_tiehi _7402__578 (.L_HI(net578));
 sg13g2_tiehi _7401__579 (.L_HI(net579));
 sg13g2_tiehi _7400__580 (.L_HI(net580));
 sg13g2_tiehi _7399__581 (.L_HI(net581));
 sg13g2_tiehi _7398__582 (.L_HI(net582));
 sg13g2_tiehi _7397__583 (.L_HI(net583));
 sg13g2_tiehi _7396__584 (.L_HI(net584));
 sg13g2_tiehi _7395__585 (.L_HI(net585));
 sg13g2_tiehi _7394__586 (.L_HI(net586));
 sg13g2_tiehi _7393__587 (.L_HI(net587));
 sg13g2_tiehi _7392__588 (.L_HI(net588));
 sg13g2_tiehi _7391__589 (.L_HI(net589));
 sg13g2_tiehi _7390__590 (.L_HI(net590));
 sg13g2_tiehi _7389__591 (.L_HI(net591));
 sg13g2_tiehi _7388__592 (.L_HI(net592));
 sg13g2_tiehi _7387__593 (.L_HI(net593));
 sg13g2_tiehi _7386__594 (.L_HI(net594));
 sg13g2_tiehi _7385__595 (.L_HI(net595));
 sg13g2_tiehi _7384__596 (.L_HI(net596));
 sg13g2_tiehi _7383__597 (.L_HI(net597));
 sg13g2_tiehi _7382__598 (.L_HI(net598));
 sg13g2_tiehi _7381__599 (.L_HI(net599));
 sg13g2_tiehi _7380__600 (.L_HI(net600));
 sg13g2_tiehi _7379__601 (.L_HI(net601));
 sg13g2_tiehi _7378__602 (.L_HI(net602));
 sg13g2_tiehi _7377__603 (.L_HI(net603));
 sg13g2_tiehi _7376__604 (.L_HI(net604));
 sg13g2_tiehi _7375__605 (.L_HI(net605));
 sg13g2_tiehi _7374__606 (.L_HI(net606));
 sg13g2_tiehi _7373__607 (.L_HI(net607));
 sg13g2_tiehi _7372__608 (.L_HI(net608));
 sg13g2_tiehi _7371__609 (.L_HI(net609));
 sg13g2_tiehi _7370__610 (.L_HI(net610));
 sg13g2_tiehi _7369__611 (.L_HI(net611));
 sg13g2_tiehi _7368__612 (.L_HI(net612));
 sg13g2_tiehi _7367__613 (.L_HI(net613));
 sg13g2_tiehi _7449__614 (.L_HI(net614));
 sg13g2_tiehi _7512__615 (.L_HI(net615));
 sg13g2_tiehi _7366__616 (.L_HI(net616));
 sg13g2_tiehi _7365__617 (.L_HI(net617));
 sg13g2_tiehi _7364__618 (.L_HI(net618));
 sg13g2_tiehi _7363__619 (.L_HI(net619));
 sg13g2_tiehi _7362__620 (.L_HI(net620));
 sg13g2_tiehi _7361__621 (.L_HI(net621));
 sg13g2_tiehi _7360__622 (.L_HI(net622));
 sg13g2_tiehi _7359__623 (.L_HI(net623));
 sg13g2_tiehi _7358__624 (.L_HI(net624));
 sg13g2_tiehi _7357__625 (.L_HI(net625));
 sg13g2_tiehi _7356__626 (.L_HI(net626));
 sg13g2_tiehi _7355__627 (.L_HI(net627));
 sg13g2_tiehi _7354__628 (.L_HI(net628));
 sg13g2_tiehi _7353__629 (.L_HI(net629));
 sg13g2_tiehi _7352__630 (.L_HI(net630));
 sg13g2_tiehi _7351__631 (.L_HI(net631));
 sg13g2_tiehi _7350__632 (.L_HI(net632));
 sg13g2_tiehi _7349__633 (.L_HI(net633));
 sg13g2_tiehi _7348__634 (.L_HI(net634));
 sg13g2_tiehi _7347__635 (.L_HI(net635));
 sg13g2_tiehi _7346__636 (.L_HI(net636));
 sg13g2_tiehi _7345__637 (.L_HI(net637));
 sg13g2_tiehi _7344__638 (.L_HI(net638));
 sg13g2_tiehi _7343__639 (.L_HI(net639));
 sg13g2_tiehi _7342__640 (.L_HI(net640));
 sg13g2_tiehi _7341__641 (.L_HI(net641));
 sg13g2_tiehi _7340__642 (.L_HI(net642));
 sg13g2_tiehi _7339__643 (.L_HI(net643));
 sg13g2_tiehi _7338__644 (.L_HI(net644));
 sg13g2_tiehi _7337__645 (.L_HI(net645));
 sg13g2_tiehi _7336__646 (.L_HI(net646));
 sg13g2_tiehi _7335__647 (.L_HI(net647));
 sg13g2_tiehi _7334__648 (.L_HI(net648));
 sg13g2_tiehi _7333__649 (.L_HI(net649));
 sg13g2_tiehi _7332__650 (.L_HI(net650));
 sg13g2_tiehi _7331__651 (.L_HI(net651));
 sg13g2_tiehi _7330__652 (.L_HI(net652));
 sg13g2_tiehi _7329__653 (.L_HI(net653));
 sg13g2_tiehi _7328__654 (.L_HI(net654));
 sg13g2_tiehi _7327__655 (.L_HI(net655));
 sg13g2_tiehi _7326__656 (.L_HI(net656));
 sg13g2_tiehi _7325__657 (.L_HI(net657));
 sg13g2_tiehi _7324__658 (.L_HI(net658));
 sg13g2_tiehi _7323__659 (.L_HI(net659));
 sg13g2_tiehi _7322__660 (.L_HI(net660));
 sg13g2_tiehi _7321__661 (.L_HI(net661));
 sg13g2_tiehi _7320__662 (.L_HI(net662));
 sg13g2_tiehi _7319__663 (.L_HI(net663));
 sg13g2_tiehi _7318__664 (.L_HI(net664));
 sg13g2_tiehi _7317__665 (.L_HI(net665));
 sg13g2_tiehi _7316__666 (.L_HI(net666));
 sg13g2_tiehi _7315__667 (.L_HI(net667));
 sg13g2_tiehi _7314__668 (.L_HI(net668));
 sg13g2_tiehi _7313__669 (.L_HI(net669));
 sg13g2_tiehi _7312__670 (.L_HI(net670));
 sg13g2_tiehi _7311__671 (.L_HI(net671));
 sg13g2_tiehi _7310__672 (.L_HI(net672));
 sg13g2_tiehi _7309__673 (.L_HI(net673));
 sg13g2_tiehi _7308__674 (.L_HI(net674));
 sg13g2_tiehi _7307__675 (.L_HI(net675));
 sg13g2_tiehi _7306__676 (.L_HI(net676));
 sg13g2_tiehi _7305__677 (.L_HI(net677));
 sg13g2_tiehi _7304__678 (.L_HI(net678));
 sg13g2_tiehi _7303__679 (.L_HI(net679));
 sg13g2_tiehi _7302__680 (.L_HI(net680));
 sg13g2_tiehi _7301__681 (.L_HI(net681));
 sg13g2_tiehi _7300__682 (.L_HI(net682));
 sg13g2_tiehi _7299__683 (.L_HI(net683));
 sg13g2_tiehi _7298__684 (.L_HI(net684));
 sg13g2_tiehi _7297__685 (.L_HI(net685));
 sg13g2_tiehi _7296__686 (.L_HI(net686));
 sg13g2_tiehi _7295__687 (.L_HI(net687));
 sg13g2_tiehi _7294__688 (.L_HI(net688));
 sg13g2_tiehi _7293__689 (.L_HI(net689));
 sg13g2_tiehi _7292__690 (.L_HI(net690));
 sg13g2_tiehi _7291__691 (.L_HI(net691));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_iitbbs_10 (.L_LO(net10));
 sg13g2_tielo tt_um_iitbbs_11 (.L_LO(net11));
 sg13g2_tielo tt_um_iitbbs_12 (.L_LO(net12));
 sg13g2_tielo tt_um_iitbbs_13 (.L_LO(net13));
 sg13g2_tielo tt_um_iitbbs_14 (.L_LO(net14));
 sg13g2_tielo tt_um_iitbbs_15 (.L_LO(net15));
 sg13g2_tielo tt_um_iitbbs_16 (.L_LO(net16));
 sg13g2_tielo tt_um_iitbbs_17 (.L_LO(net17));
 sg13g2_tielo tt_um_iitbbs_18 (.L_LO(net18));
 sg13g2_tielo tt_um_iitbbs_19 (.L_LO(net19));
 sg13g2_tielo tt_um_iitbbs_20 (.L_LO(net20));
 sg13g2_tielo tt_um_iitbbs_21 (.L_LO(net21));
 sg13g2_tielo tt_um_iitbbs_22 (.L_LO(net22));
 sg13g2_tielo tt_um_iitbbs_23 (.L_LO(net23));
 sg13g2_tielo tt_um_iitbbs_24 (.L_LO(net24));
 sg13g2_tiehi _7290__25 (.L_HI(net25));
 sg13g2_buf_2 _8274_ (.A(\L1_Digit[0].L2_Leds[7].L2_viz_lit_a0 ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout757 (.A(_2282_),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(_2282_),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(_2280_),
    .X(net759));
 sg13g2_buf_4 fanout760 (.X(net760),
    .A(_2280_));
 sg13g2_buf_4 fanout761 (.X(net761),
    .A(_2274_));
 sg13g2_buf_4 fanout762 (.X(net762),
    .A(_2274_));
 sg13g2_buf_2 fanout763 (.A(_2384_),
    .X(net763));
 sg13g2_buf_4 fanout764 (.X(net764),
    .A(_2278_));
 sg13g2_buf_4 fanout765 (.X(net765),
    .A(_2278_));
 sg13g2_buf_2 fanout766 (.A(_2276_),
    .X(net766));
 sg13g2_buf_4 fanout767 (.X(net767),
    .A(_2276_));
 sg13g2_buf_2 fanout768 (.A(net770),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(net771),
    .X(net769));
 sg13g2_buf_1 fanout770 (.A(net771),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(_2383_),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(_2272_),
    .X(net772));
 sg13g2_buf_2 fanout773 (.A(_2272_),
    .X(net773));
 sg13g2_buf_2 fanout774 (.A(_2270_),
    .X(net774));
 sg13g2_buf_4 fanout775 (.X(net775),
    .A(_2270_));
 sg13g2_buf_4 fanout776 (.X(net776),
    .A(_2268_));
 sg13g2_buf_4 fanout777 (.X(net777),
    .A(_2268_));
 sg13g2_buf_4 fanout778 (.X(net778),
    .A(_2463_));
 sg13g2_buf_4 fanout779 (.X(net779),
    .A(_2320_));
 sg13g2_buf_2 fanout780 (.A(_1382_),
    .X(net780));
 sg13g2_buf_2 fanout781 (.A(_1357_),
    .X(net781));
 sg13g2_buf_1 fanout782 (.A(_1357_),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(_1952_),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(_1385_),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(_1376_),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(_1373_),
    .X(net786));
 sg13g2_buf_2 fanout787 (.A(_1373_),
    .X(net787));
 sg13g2_buf_2 fanout788 (.A(net789),
    .X(net788));
 sg13g2_buf_2 fanout789 (.A(_1366_),
    .X(net789));
 sg13g2_buf_2 fanout790 (.A(_1359_),
    .X(net790));
 sg13g2_buf_2 fanout791 (.A(_1351_),
    .X(net791));
 sg13g2_buf_2 fanout792 (.A(_1344_),
    .X(net792));
 sg13g2_buf_2 fanout793 (.A(_1339_),
    .X(net793));
 sg13g2_buf_4 fanout794 (.X(net794),
    .A(\FpgaPins_Fpga_FSM_idata_rd_addr_a1[3] ));
 sg13g2_buf_2 fanout795 (.A(net796),
    .X(net795));
 sg13g2_buf_1 fanout796 (.A(net797),
    .X(net796));
 sg13g2_buf_2 fanout797 (.A(\FpgaPins_Fpga_FSM_idata_rd_addr_a1[2] ),
    .X(net797));
 sg13g2_buf_2 fanout798 (.A(\FpgaPins_Fpga_FSM_idata_rd_addr_a1[0] ),
    .X(net798));
 sg13g2_buf_4 fanout799 (.X(net799),
    .A(\FpgaPins_Fpga_FSM_idata_rd_addr_a1[0] ));
 sg13g2_buf_2 fanout800 (.A(_1298_),
    .X(net800));
 sg13g2_buf_2 fanout801 (.A(_1372_),
    .X(net801));
 sg13g2_buf_2 fanout802 (.A(_1316_),
    .X(net802));
 sg13g2_buf_4 fanout803 (.X(net803),
    .A(_1316_));
 sg13g2_buf_8 fanout804 (.A(net806),
    .X(net804));
 sg13g2_buf_4 fanout805 (.X(net805),
    .A(net806));
 sg13g2_buf_4 fanout806 (.X(net806),
    .A(_1310_));
 sg13g2_buf_4 fanout807 (.X(net807),
    .A(net808));
 sg13g2_buf_4 fanout808 (.X(net808),
    .A(_1310_));
 sg13g2_buf_4 fanout809 (.X(net809),
    .A(net811));
 sg13g2_buf_4 fanout810 (.X(net810),
    .A(net811));
 sg13g2_buf_2 fanout811 (.A(_1310_),
    .X(net811));
 sg13g2_buf_4 fanout812 (.X(net812),
    .A(net814));
 sg13g2_buf_4 fanout813 (.X(net813),
    .A(net814));
 sg13g2_buf_2 fanout814 (.A(\FpgaPins_Fpga_FSM_idata_rd_addr_a1[1] ),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(net817),
    .X(net815));
 sg13g2_buf_1 fanout816 (.A(net817),
    .X(net816));
 sg13g2_buf_2 fanout817 (.A(\FpgaPins_Fpga_FSM_idata_rd_addr_a1[1] ),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(net819),
    .X(net818));
 sg13g2_buf_2 fanout819 (.A(\FpgaPins_Fpga_FSM_idata_rd_addr_a1[1] ),
    .X(net819));
 sg13g2_buf_2 fanout820 (.A(_2381_),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(_2381_),
    .X(net821));
 sg13g2_buf_2 fanout822 (.A(_1285_),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(net824),
    .X(net823));
 sg13g2_buf_2 fanout824 (.A(_2625_),
    .X(net824));
 sg13g2_buf_2 fanout825 (.A(net826),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(_2565_),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(net828),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(_2519_),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(_2497_),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(_2497_),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(net832),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(_2487_),
    .X(net832));
 sg13g2_buf_4 fanout833 (.X(net833),
    .A(_2476_));
 sg13g2_buf_2 fanout834 (.A(_2476_),
    .X(net834));
 sg13g2_buf_2 fanout835 (.A(net836),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(_2466_),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(net838),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(_2369_),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(net840),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(_2359_),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(net842),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(_2322_),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(net844),
    .X(net843));
 sg13g2_buf_4 fanout844 (.X(net844),
    .A(_2305_));
 sg13g2_buf_2 fanout845 (.A(net846),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(_2293_),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(net848),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(_2248_),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(_2163_),
    .X(net849));
 sg13g2_buf_4 fanout850 (.X(net850),
    .A(_2040_));
 sg13g2_buf_2 fanout851 (.A(net852),
    .X(net851));
 sg13g2_buf_4 fanout852 (.X(net852),
    .A(_2040_));
 sg13g2_buf_4 fanout853 (.X(net853),
    .A(net854));
 sg13g2_buf_4 fanout854 (.X(net854),
    .A(_2029_));
 sg13g2_buf_1 fanout855 (.A(_2029_),
    .X(net855));
 sg13g2_buf_4 fanout856 (.X(net856),
    .A(net858));
 sg13g2_buf_4 fanout857 (.X(net857),
    .A(net858));
 sg13g2_buf_4 fanout858 (.X(net858),
    .A(_2006_));
 sg13g2_buf_2 fanout859 (.A(\FpgaPins_Fpga_FSM_instr_a1[0] ),
    .X(net859));
 sg13g2_buf_4 fanout860 (.X(net860),
    .A(net862));
 sg13g2_buf_4 fanout861 (.X(net861),
    .A(net862));
 sg13g2_buf_4 fanout862 (.X(net862),
    .A(_2018_));
 sg13g2_buf_4 fanout863 (.X(net863),
    .A(net865));
 sg13g2_buf_2 fanout864 (.A(net865),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(_1992_),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(net868),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(net868),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(_1985_),
    .X(net868));
 sg13g2_buf_2 fanout869 (.A(_1975_),
    .X(net869));
 sg13g2_buf_1 fanout870 (.A(net871),
    .X(net870));
 sg13g2_buf_4 fanout871 (.X(net871),
    .A(_1975_));
 sg13g2_buf_2 fanout872 (.A(net874),
    .X(net872));
 sg13g2_buf_1 fanout873 (.A(net874),
    .X(net873));
 sg13g2_buf_4 fanout874 (.X(net874),
    .A(_1967_));
 sg13g2_buf_4 fanout875 (.X(net875),
    .A(\FpgaPins_Fpga_FSM_instr_a1[5] ));
 sg13g2_buf_2 fanout876 (.A(net877),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(_2510_),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(_2284_),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(_2284_),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(_2166_),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(_2817_),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(net883),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(_2788_),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(_2787_),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(_2787_),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(net890),
    .X(net886));
 sg13g2_buf_2 fanout887 (.A(net888),
    .X(net887));
 sg13g2_buf_1 fanout888 (.A(net890),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(net890),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(_2769_),
    .X(net890));
 sg13g2_buf_4 fanout891 (.X(net891),
    .A(\FpgaPins_Fpga_FSM_imem_rd_addr_a1[3] ));
 sg13g2_buf_2 fanout892 (.A(_0780_),
    .X(net892));
 sg13g2_buf_1 fanout893 (.A(_0780_),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(_0922_),
    .X(net894));
 sg13g2_buf_1 fanout895 (.A(_0922_),
    .X(net895));
 sg13g2_buf_4 fanout896 (.X(net896),
    .A(_0840_));
 sg13g2_buf_2 fanout897 (.A(_0779_),
    .X(net897));
 sg13g2_buf_1 fanout898 (.A(_0779_),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(net901),
    .X(net899));
 sg13g2_buf_1 fanout900 (.A(net901),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(_2579_),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(_1956_),
    .X(net902));
 sg13g2_buf_2 fanout903 (.A(net905),
    .X(net903));
 sg13g2_buf_2 fanout904 (.A(net905),
    .X(net904));
 sg13g2_buf_2 fanout905 (.A(_0963_),
    .X(net905));
 sg13g2_buf_2 fanout906 (.A(net907),
    .X(net906));
 sg13g2_buf_2 fanout907 (.A(_0823_),
    .X(net907));
 sg13g2_buf_2 fanout908 (.A(net910),
    .X(net908));
 sg13g2_buf_1 fanout909 (.A(net910),
    .X(net909));
 sg13g2_buf_2 fanout910 (.A(_0823_),
    .X(net910));
 sg13g2_buf_4 fanout911 (.X(net911),
    .A(\FpgaPins_Fpga_FSM_imem_rd_addr_a1[0] ));
 sg13g2_buf_2 fanout912 (.A(\FpgaPins_Fpga_FSM_imem_rd_addr_a1[0] ),
    .X(net912));
 sg13g2_buf_2 fanout913 (.A(net915),
    .X(net913));
 sg13g2_buf_4 fanout914 (.X(net914),
    .A(net915));
 sg13g2_buf_2 fanout915 (.A(\FpgaPins_Fpga_FSM_imem_rd_addr_a1[0] ),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(_0889_),
    .X(net916));
 sg13g2_buf_1 fanout917 (.A(_0889_),
    .X(net917));
 sg13g2_buf_4 fanout918 (.X(net918),
    .A(net920));
 sg13g2_buf_1 fanout919 (.A(net920),
    .X(net919));
 sg13g2_buf_4 fanout920 (.X(net920),
    .A(net924));
 sg13g2_buf_2 fanout921 (.A(net922),
    .X(net921));
 sg13g2_buf_4 fanout922 (.X(net922),
    .A(net923));
 sg13g2_buf_4 fanout923 (.X(net923),
    .A(net924));
 sg13g2_buf_4 fanout924 (.X(net924),
    .A(\FpgaPins_Fpga_FSM_imem_rd_addr_a1[1] ));
 sg13g2_buf_2 fanout925 (.A(net927),
    .X(net925));
 sg13g2_buf_8 fanout926 (.A(net927),
    .X(net926));
 sg13g2_buf_2 fanout927 (.A(net932),
    .X(net927));
 sg13g2_buf_2 fanout928 (.A(net929),
    .X(net928));
 sg13g2_buf_2 fanout929 (.A(net931),
    .X(net929));
 sg13g2_buf_4 fanout930 (.X(net930),
    .A(net931));
 sg13g2_buf_8 fanout931 (.A(net932),
    .X(net931));
 sg13g2_buf_4 fanout932 (.X(net932),
    .A(_0808_));
 sg13g2_buf_2 fanout933 (.A(_1737_),
    .X(net933));
 sg13g2_buf_2 fanout934 (.A(_1737_),
    .X(net934));
 sg13g2_buf_4 fanout935 (.X(net935),
    .A(_2791_));
 sg13g2_buf_4 fanout936 (.X(net936),
    .A(_1837_));
 sg13g2_buf_2 fanout937 (.A(_1837_),
    .X(net937));
 sg13g2_buf_2 fanout938 (.A(net939),
    .X(net938));
 sg13g2_buf_2 fanout939 (.A(_1741_),
    .X(net939));
 sg13g2_buf_2 fanout940 (.A(net941),
    .X(net940));
 sg13g2_buf_2 fanout941 (.A(_0802_),
    .X(net941));
 sg13g2_buf_2 fanout942 (.A(_0799_),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(_0799_),
    .X(net943));
 sg13g2_buf_2 fanout944 (.A(net946),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(net946),
    .X(net945));
 sg13g2_buf_2 fanout946 (.A(net947),
    .X(net946));
 sg13g2_buf_4 fanout947 (.X(net947),
    .A(FpgaPins_Fpga_LIPSI_reset_a1));
 sg13g2_buf_4 fanout948 (.X(net948),
    .A(net952));
 sg13g2_buf_2 fanout949 (.A(net950),
    .X(net949));
 sg13g2_buf_2 fanout950 (.A(net952),
    .X(net950));
 sg13g2_buf_4 fanout951 (.X(net951),
    .A(net952));
 sg13g2_buf_4 fanout952 (.X(net952),
    .A(_1940_));
 sg13g2_buf_2 fanout953 (.A(net954),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(net955),
    .X(net954));
 sg13g2_buf_4 fanout955 (.X(net955),
    .A(net962));
 sg13g2_buf_2 fanout956 (.A(net960),
    .X(net956));
 sg13g2_buf_1 fanout957 (.A(net960),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(net960),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(net960),
    .X(net959));
 sg13g2_buf_1 fanout960 (.A(net961),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(net962),
    .X(net961));
 sg13g2_buf_4 fanout962 (.X(net962),
    .A(_1939_));
 sg13g2_buf_2 fanout963 (.A(net964),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(net966),
    .X(net964));
 sg13g2_buf_2 fanout965 (.A(net966),
    .X(net965));
 sg13g2_buf_4 fanout966 (.X(net966),
    .A(net969));
 sg13g2_buf_2 fanout967 (.A(net968),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(net969),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(_1188_),
    .X(net969));
 sg13g2_buf_2 fanout970 (.A(net974),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(net973),
    .X(net971));
 sg13g2_buf_1 fanout972 (.A(net973),
    .X(net972));
 sg13g2_buf_1 fanout973 (.A(net974),
    .X(net973));
 sg13g2_buf_4 fanout974 (.X(net974),
    .A(_1187_));
 sg13g2_buf_2 fanout975 (.A(net976),
    .X(net975));
 sg13g2_buf_4 fanout976 (.X(net976),
    .A(net977));
 sg13g2_buf_4 fanout977 (.X(net977),
    .A(_0796_));
 sg13g2_buf_2 fanout978 (.A(_0785_),
    .X(net978));
 sg13g2_buf_1 fanout979 (.A(_0785_),
    .X(net979));
 sg13g2_buf_2 fanout980 (.A(_0784_),
    .X(net980));
 sg13g2_buf_4 fanout981 (.X(net981),
    .A(_0728_));
 sg13g2_buf_2 fanout982 (.A(_0101_),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(net984),
    .X(net983));
 sg13g2_buf_2 fanout984 (.A(FpgaPins_Fpga_GAME_forward_a2),
    .X(net984));
 sg13g2_buf_4 fanout985 (.X(net985),
    .A(_0017_));
 sg13g2_buf_2 fanout986 (.A(net987),
    .X(net986));
 sg13g2_buf_2 fanout987 (.A(FpgaPins_Fpga_LIPSI_is_brl_a2),
    .X(net987));
 sg13g2_buf_2 fanout988 (.A(net989),
    .X(net988));
 sg13g2_buf_2 fanout989 (.A(FpgaPins_Fpga_LIPSI_is_ld_ind_a2),
    .X(net989));
 sg13g2_buf_4 fanout990 (.X(net990),
    .A(FpgaPins_Fpga_LIPSI_is_ret_a2));
 sg13g2_buf_2 fanout991 (.A(net1753),
    .X(net991));
 sg13g2_buf_4 fanout992 (.X(net992),
    .A(net1179));
 sg13g2_buf_2 fanout993 (.A(net1732),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(net995),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(net1733),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(_1186_),
    .X(net996));
 sg13g2_buf_4 fanout997 (.X(net997),
    .A(_0722_));
 sg13g2_buf_2 fanout998 (.A(net8),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(net1000),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(net1001),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(net1002),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(ui_in[1]),
    .X(net1002));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_4 input2 (.X(net2),
    .A(ui_in[0]));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[3]));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_iitbbs_9 (.L_LO(net9));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_leaf_62_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_2 clkbuf_leaf_63_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_2 clkbuf_leaf_64_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_2 clkbuf_leaf_65_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_2 clkbuf_leaf_66_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_2 clkbuf_leaf_67_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_2 clkbuf_leaf_68_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_2 clkbuf_leaf_69_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_2 clkbuf_leaf_70_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_2 clkbuf_leaf_71_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_2 clkbuf_leaf_72_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_2 clkbuf_leaf_73_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_2 clkbuf_leaf_74_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_2 clkbuf_leaf_75_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_2 clkbuf_leaf_76_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_2 clkbuf_leaf_77_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_2 clkbuf_leaf_78_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_2 clkbuf_leaf_79_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_2 clkbuf_leaf_80_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_2 clkbuf_leaf_81_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_2 clkbuf_leaf_82_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_2 clkbuf_leaf_83_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_2 clkbuf_leaf_84_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_2 clkbuf_leaf_85_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_2 clkbuf_leaf_86_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_2 clkbuf_leaf_87_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_2 clkbuf_leaf_88_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_2 clkbuf_leaf_89_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_2 clkbuf_leaf_90_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_4_7_0_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_4_11_0_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_4_13_0_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_leaf_4_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_5_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_6_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_10_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_16_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_17_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_27_clk));
 sg13g2_inv_4 clkload12 (.A(clknet_leaf_11_clk));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_12_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_leaf_15_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_33_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_28_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_29_clk));
 sg13g2_inv_4 clkload18 (.A(clknet_leaf_32_clk));
 sg13g2_inv_1 clkload19 (.A(clknet_leaf_70_clk));
 sg13g2_inv_2 clkload20 (.A(clknet_leaf_61_clk));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_62_clk));
 sg13g2_inv_2 clkload22 (.A(clknet_leaf_78_clk));
 sg13g2_inv_1 clkload23 (.A(clknet_leaf_57_clk));
 sg13g2_inv_4 clkload24 (.A(clknet_leaf_68_clk));
 sg13g2_inv_8 clkload25 (.A(clknet_leaf_67_clk));
 sg13g2_inv_1 clkload26 (.A(clknet_leaf_41_clk));
 sg13g2_inv_4 clkload27 (.A(clknet_leaf_42_clk));
 sg13g2_inv_1 clkload28 (.A(clknet_leaf_43_clk));
 sg13g2_inv_1 clkload29 (.A(clknet_leaf_44_clk));
 sg13g2_inv_4 clkload30 (.A(clknet_leaf_51_clk));
 sg13g2_inv_4 clkload31 (.A(clknet_leaf_58_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(FpgaPins_Fpga_LIPSI_is_brz_a2),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold2 (.A(\FpgaPins_Fpga_GAME_score_a3[1] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold3 (.A(\uart_rx_1.r_Rx_Data_R ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold4 (.A(FpgaPins_Fpga_LIPSI_is_br_a2),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold5 (.A(\FpgaPins_Fpga_GAME_score_a3[6] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold6 (.A(\FpgaPins_Fpga_GAME_score_a3[0] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold7 (.A(\FpgaPins_Fpga_GAME_score_a3[2] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold8 (.A(\FpgaPins_Fpga_GAME_score_a3[7] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold9 (.A(\FpgaPins_Fpga_GAME_score_a3[5] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold10 (.A(FpgaPins_Fpga_LIPSI_is_brnz_a2),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold11 (.A(\FpgaPins_Fpga_GAME_score_a3[4] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold12 (.A(\FpgaPins_Fpga_GAME_score_a3[3] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold13 (.A(\FpgaPins_Fpga_GAME_state_a2[1] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold14 (.A(FpgaPins_Fpga_GAME_clk_pulse_a2),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold15 (.A(\FpgaPins_Fpga_GAME_state_a2[0] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold16 (.A(\FpgaPins_Fpga_GAME_state_a3[1] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold17 (.A(\FpgaPins_Fpga_GAME_state_a3[0] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0206_),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold19 (.A(\FpgaPins_Fpga_GAME_score_a2[5] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold20 (.A(\FpgaPins_Fpga_GAME_led_output_a2[2] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold21 (.A(\FpgaPins_Fpga_GAME_score_a2[1] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold22 (.A(\FpgaPins_Fpga_GAME_score_a2[2] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold23 (.A(\FpgaPins_Fpga_GAME_score_a2[7] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold24 (.A(\FpgaPins_Fpga_GAME_score_a2[3] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold25 (.A(\FpgaPins_Fpga_GAME_score_a2[4] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0198_),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold27 (.A(\FpgaPins_Fpga_LIPSI_pc_a1[6] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold28 (.A(\FpgaPins_Fpga_GAME_led_output_a2[0] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold29 (.A(\FpgaPins_Fpga_GAME_score_a2[0] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold30 (.A(\FpgaPins_Fpga_GAME_score_a2[6] ),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold31 (.A(\FpgaPins_Fpga_GAME_led_output_a2[3] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold32 (.A(\FpgaPins_Fpga_GAME_led_output_a2[1] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold33 (.A(\FpgaPins_Fpga_GAME_led_output_a2[7] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold34 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[0] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0207_),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0339_),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold37 (.A(\instrs[11][5] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold38 (.A(\FpgaPins_Fpga_UART_dptr_a2[3] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0342_),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold40 (.A(\uart_rx_1.r_Bit_Index[6] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold41 (.A(\uart_rx_1.r_Bit_Index[7] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold42 (.A(\uart_rx_1.r_Bit_Index[10] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold43 (.A(\uart_rx_1.r_Bit_Index[18] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0200_),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold45 (.A(\FpgaPins_Fpga_LIPSI_pc_a1[7] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold46 (.A(\instrs[7][0] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold47 (.A(\uart_rx_1.r_Bit_Index[22] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0196_),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold49 (.A(\FpgaPins_Fpga_LIPSI_pc_a1[5] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold50 (.A(\uart_rx_1.r_Bit_Index[9] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold51 (.A(\FpgaPins_Fpga_GAME_led_output_a2[6] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold52 (.A(\uart_rx_1.r_Bit_Index[23] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold53 (.A(\instrs[3][0] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold54 (.A(\FpgaPins_Fpga_UART_dptr_a2[2] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0341_),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold56 (.A(\uart_rx_1.r_Bit_Index[17] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold57 (.A(\uart_rx_1.r_Bit_Index[27] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold58 (.A(\instrs[3][7] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold59 (.A(\instrs[7][7] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold60 (.A(\C1.counter_status[2] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold61 (.A(\uart_rx_1.r_Bit_Index[11] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold62 (.A(\C1.counter2[31] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0338_),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold64 (.A(\uart_rx_1.r_Bit_Index[16] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold65 (.A(\uart_rx_1.r_Bit_Index[8] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold66 (.A(\uart_rx_1.r_Bit_Index[20] ),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold67 (.A(\instrs[3][5] ),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold68 (.A(\uart_rx_1.r_Bit_Index[19] ),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold69 (.A(\FpgaPins_Fpga_GAME_led_output_a2[4] ),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold70 (.A(\uart_rx_1.r_Bit_Index[21] ),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold71 (.A(\instrs[11][7] ),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold72 (.A(\instrs[11][0] ),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold73 (.A(\instrs[7][5] ),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold74 (.A(\uart_rx_1.r_Bit_Index[24] ),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold75 (.A(\uart_rx_1.r_Bit_Index[15] ),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold76 (.A(\FpgaPins_Fpga_GAME_led_output_a2[5] ),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0014_),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold78 (.A(\instrs[7][3] ),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold79 (.A(\uart_rx_1.r_Bit_Index[26] ),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold80 (.A(\uart_rx_1.r_Bit_Index[13] ),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold81 (.A(\instrs[11][2] ),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold82 (.A(\instrs[11][3] ),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold83 (.A(\instrs[10][0] ),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold84 (.A(\instrs[3][2] ),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold85 (.A(\instrs[3][6] ),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold86 (.A(\instrs[3][3] ),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold87 (.A(\instrs[1][7] ),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold88 (.A(\instrs[13][5] ),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold89 (.A(\instrs[7][6] ),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold90 (.A(\instrs[11][1] ),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold91 (.A(\uart_rx_1.r_Bit_Index[25] ),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold92 (.A(\instrs[9][7] ),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold93 (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[18] ),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold94 (.A(\FpgaPins_Fpga_GAME_count_speed4_a1[18] ),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold95 (.A(\instrs[15][5] ),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold96 (.A(\instrs[3][4] ),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold97 (.A(\instrs[4][5] ),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold98 (.A(\instrs[4][0] ),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold99 (.A(\instrs[5][7] ),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold100 (.A(\instrs[7][2] ),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold101 (.A(\datam[8][3] ),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold102 (.A(\instrs[0][0] ),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold103 (.A(\instrs[7][4] ),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0246_),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0208_),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0325_),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold107 (.A(\instrs[0][7] ),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold108 (.A(\datam[12][4] ),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold109 (.A(\instrs[15][0] ),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold110 (.A(\instrs[14][0] ),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0514_),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold112 (.A(\instrs[6][0] ),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold113 (.A(\datam[12][3] ),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold114 (.A(\instrs[6][5] ),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold115 (.A(\datam[0][1] ),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold116 (.A(\datam[4][0] ),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold117 (.A(\uart_rx_1.r_Bit_Index[14] ),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold118 (.A(\datam[8][1] ),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold119 (.A(\datam[4][4] ),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold120 (.A(\datam[0][4] ),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold121 (.A(\datam[8][0] ),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold122 (.A(\datam[4][2] ),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold123 (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[0] ),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold124 (.A(\instrs[11][4] ),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0270_),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold126 (.A(\datam[8][4] ),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold127 (.A(\datam[8][2] ),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold128 (.A(\datam[4][1] ),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold129 (.A(\instrs[1][5] ),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold130 (.A(\uart_rx_1.r_Clock_Count[21] ),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0646_),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold132 (.A(\instrs[13][7] ),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold133 (.A(\instrs[9][5] ),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold134 (.A(\instrs[6][7] ),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold135 (.A(\datam[12][1] ),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold136 (.A(\datam[0][3] ),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold137 (.A(\datam[12][0] ),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold138 (.A(\uart_rx_1.r_Clock_Count[31] ),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0656_),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold140 (.A(\instrs[10][7] ),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold141 (.A(\datam[0][0] ),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold142 (.A(\instrs[7][1] ),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold143 (.A(\uart_rx_1.r_Clock_Count[13] ),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0638_),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold145 (.A(\uart_rx_1.r_Clock_Count[20] ),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold146 (.A(_2858_),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold147 (.A(\instrs[4][7] ),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold148 (.A(\datam[0][2] ),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold149 (.A(\instrs[1][0] ),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold150 (.A(\datam[4][3] ),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold151 (.A(\datam[12][2] ),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold152 (.A(\instrs[10][5] ),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold153 (.A(\instrs[14][5] ),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold154 (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[1] ),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold155 (.A(\FpgaPins_Fpga_GAME_count_speed3_a1[1] ),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold156 (.A(\instrs[8][5] ),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold157 (.A(\uart_rx_1.r_Clock_Count[16] ),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold158 (.A(_2844_),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold159 (.A(\instrs[12][5] ),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold160 (.A(\uart_rx_1.r_Clock_Count[12] ),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold161 (.A(_2830_),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold162 (.A(\datam[13][5] ),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold163 (.A(\instrs[8][0] ),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold164 (.A(\instrs[14][7] ),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0194_),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold166 (.A(_2000_),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold167 (.A(\FpgaPins_Fpga_LIPSI_pc_a1[4] ),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold168 (.A(\FpgaPins_Fpga_LIPSI_data_wr_a2[0] ),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold169 (.A(\instrs[5][5] ),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold170 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[24] ),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold171 (.A(_2624_),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold172 (.A(\C1.level_op ),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0573_),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold174 (.A(\instrs[12][7] ),
    .X(net1111));
 sg13g2_dlygate4sd3_1 hold175 (.A(\instrs[5][6] ),
    .X(net1112));
 sg13g2_dlygate4sd3_1 hold176 (.A(\instrs[0][1] ),
    .X(net1113));
 sg13g2_dlygate4sd3_1 hold177 (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[16] ),
    .X(net1114));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0899_),
    .X(net1115));
 sg13g2_dlygate4sd3_1 hold179 (.A(\FpgaPins_Fpga_LIPSI_data_wr_a2[1] ),
    .X(net1116));
 sg13g2_dlygate4sd3_1 hold180 (.A(\FpgaPins_Fpga_LIPSI_data_wr_a2[2] ),
    .X(net1117));
 sg13g2_dlygate4sd3_1 hold181 (.A(\instrs[13][0] ),
    .X(net1118));
 sg13g2_dlygate4sd3_1 hold182 (.A(\instrs[9][4] ),
    .X(net1119));
 sg13g2_dlygate4sd3_1 hold183 (.A(\uart_rx_1.r_Clock_Count[19] ),
    .X(net1120));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0644_),
    .X(net1121));
 sg13g2_dlygate4sd3_1 hold185 (.A(\instrs[0][5] ),
    .X(net1122));
 sg13g2_dlygate4sd3_1 hold186 (.A(\C1.temp_op ),
    .X(net1123));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0574_),
    .X(net1124));
 sg13g2_dlygate4sd3_1 hold188 (.A(\instrs[1][3] ),
    .X(net1125));
 sg13g2_dlygate4sd3_1 hold189 (.A(\instrs[12][2] ),
    .X(net1126));
 sg13g2_dlygate4sd3_1 hold190 (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[2] ),
    .X(net1127));
 sg13g2_dlygate4sd3_1 hold191 (.A(_1115_),
    .X(net1128));
 sg13g2_dlygate4sd3_1 hold192 (.A(\FpgaPins_Fpga_GAME_count_speed2_a1[2] ),
    .X(net1129));
 sg13g2_dlygate4sd3_1 hold193 (.A(\FpgaPins_Fpga_LIPSI_data_wr_a2[3] ),
    .X(net1130));
 sg13g2_dlygate4sd3_1 hold194 (.A(\instrs[8][7] ),
    .X(net1131));
 sg13g2_dlygate4sd3_1 hold195 (.A(\instrs[6][6] ),
    .X(net1132));
 sg13g2_dlygate4sd3_1 hold196 (.A(\instrs[4][6] ),
    .X(net1133));
 sg13g2_dlygate4sd3_1 hold197 (.A(\instrs[2][5] ),
    .X(net1134));
 sg13g2_dlygate4sd3_1 hold198 (.A(\FpgaPins_Fpga_LIPSI_data_wr_a2[5] ),
    .X(net1135));
 sg13g2_dlygate4sd3_1 hold199 (.A(\instrs[2][0] ),
    .X(net1136));
 sg13g2_dlygate4sd3_1 hold200 (.A(\instrs[1][4] ),
    .X(net1137));
 sg13g2_dlygate4sd3_1 hold201 (.A(\instrs[15][7] ),
    .X(net1138));
 sg13g2_dlygate4sd3_1 hold202 (.A(\uart_rx_1.r_Clock_Count[22] ),
    .X(net1139));
 sg13g2_dlygate4sd3_1 hold203 (.A(\instrs[9][0] ),
    .X(net1140));
 sg13g2_dlygate4sd3_1 hold204 (.A(\instrs[6][3] ),
    .X(net1141));
 sg13g2_dlygate4sd3_1 hold205 (.A(\uart_rx_1.r_Clock_Count[27] ),
    .X(net1142));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0652_),
    .X(net1143));
 sg13g2_dlygate4sd3_1 hold207 (.A(\uart_rx_1.r_Clock_Count[14] ),
    .X(net1144));
 sg13g2_dlygate4sd3_1 hold208 (.A(\instrs[1][1] ),
    .X(net1145));
 sg13g2_dlygate4sd3_1 hold209 (.A(\instrs[8][6] ),
    .X(net1146));
 sg13g2_dlygate4sd3_1 hold210 (.A(\instrs[5][0] ),
    .X(net1147));
 sg13g2_dlygate4sd3_1 hold211 (.A(\instrs[12][1] ),
    .X(net1148));
 sg13g2_dlygate4sd3_1 hold212 (.A(\instrs[12][3] ),
    .X(net1149));
 sg13g2_dlygate4sd3_1 hold213 (.A(\instrs[13][3] ),
    .X(net1150));
 sg13g2_dlygate4sd3_1 hold214 (.A(\instrs[12][4] ),
    .X(net1151));
 sg13g2_dlygate4sd3_1 hold215 (.A(\instrs[0][3] ),
    .X(net1152));
 sg13g2_dlygate4sd3_1 hold216 (.A(\instrs[12][0] ),
    .X(net1153));
 sg13g2_dlygate4sd3_1 hold217 (.A(_2360_),
    .X(net1154));
 sg13g2_dlygate4sd3_1 hold218 (.A(\instrs[12][6] ),
    .X(net1155));
 sg13g2_dlygate4sd3_1 hold219 (.A(\uart_rx_1.r_Clock_Count[25] ),
    .X(net1156));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0650_),
    .X(net1157));
 sg13g2_dlygate4sd3_1 hold221 (.A(\instrs[5][1] ),
    .X(net1158));
 sg13g2_dlygate4sd3_1 hold222 (.A(FpgaPins_Fpga_GAME_clk_pulse3_a2),
    .X(net1159));
 sg13g2_dlygate4sd3_1 hold223 (.A(FpgaPins_Fpga_GAME_clk_pulse3_a1),
    .X(net1160));
 sg13g2_dlygate4sd3_1 hold224 (.A(\instrs[10][2] ),
    .X(net1161));
 sg13g2_dlygate4sd3_1 hold225 (.A(\instrs[3][1] ),
    .X(net1162));
 sg13g2_dlygate4sd3_1 hold226 (.A(\instrs[2][7] ),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold227 (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[2] ),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold228 (.A(_1094_),
    .X(net1165));
 sg13g2_dlygate4sd3_1 hold229 (.A(\FpgaPins_Fpga_GAME_count_speed4_a1[2] ),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold230 (.A(\uart_rx_1.r_Clock_Count[10] ),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold231 (.A(_2820_),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold232 (.A(\uart_rx_1.r_Clock_Count[15] ),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold233 (.A(\uart_rx_1.r_Clock_Count[26] ),
    .X(net1170));
 sg13g2_dlygate4sd3_1 hold234 (.A(\instrs[8][1] ),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold235 (.A(\instrs[10][1] ),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold236 (.A(\uart_rx_1.r_Clock_Count[8] ),
    .X(net1173));
 sg13g2_dlygate4sd3_1 hold237 (.A(_2815_),
    .X(net1174));
 sg13g2_dlygate4sd3_1 hold238 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[2] ),
    .X(net1175));
 sg13g2_dlygate4sd3_1 hold239 (.A(_2583_),
    .X(net1176));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0524_),
    .X(net1177));
 sg13g2_dlygate4sd3_1 hold241 (.A(\uart_rx_1.r_Bit_Index[30] ),
    .X(net1178));
 sg13g2_dlygate4sd3_1 hold242 (.A(\C1.next_state_var[7] ),
    .X(net1179));
 sg13g2_dlygate4sd3_1 hold243 (.A(_1228_),
    .X(net1180));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0003_),
    .X(net1181));
 sg13g2_dlygate4sd3_1 hold245 (.A(\instrs[8][4] ),
    .X(net1182));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0238_),
    .X(net1183));
 sg13g2_dlygate4sd3_1 hold247 (.A(\instrs[9][3] ),
    .X(net1184));
 sg13g2_dlygate4sd3_1 hold248 (.A(\FpgaPins_Fpga_LIPSI_data_wr_a2[4] ),
    .X(net1185));
 sg13g2_dlygate4sd3_1 hold249 (.A(\C1.counter2[25] ),
    .X(net1186));
 sg13g2_dlygate4sd3_1 hold250 (.A(_2389_),
    .X(net1187));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0332_),
    .X(net1188));
 sg13g2_dlygate4sd3_1 hold252 (.A(\instrs[15][3] ),
    .X(net1189));
 sg13g2_dlygate4sd3_1 hold253 (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[0] ),
    .X(net1190));
 sg13g2_dlygate4sd3_1 hold254 (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[2] ),
    .X(net1191));
 sg13g2_dlygate4sd3_1 hold255 (.A(\instrs[0][6] ),
    .X(net1192));
 sg13g2_dlygate4sd3_1 hold256 (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[19] ),
    .X(net1193));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0975_),
    .X(net1194));
 sg13g2_dlygate4sd3_1 hold258 (.A(\FpgaPins_Fpga_GAME_count_speed2_a1[19] ),
    .X(net1195));
 sg13g2_dlygate4sd3_1 hold259 (.A(\instrs[0][2] ),
    .X(net1196));
 sg13g2_dlygate4sd3_1 hold260 (.A(\datam[0][7] ),
    .X(net1197));
 sg13g2_dlygate4sd3_1 hold261 (.A(\instrs[10][4] ),
    .X(net1198));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0214_),
    .X(net1199));
 sg13g2_dlygate4sd3_1 hold263 (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[13] ),
    .X(net1200));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0926_),
    .X(net1201));
 sg13g2_dlygate4sd3_1 hold265 (.A(\instrs[15][2] ),
    .X(net1202));
 sg13g2_dlygate4sd3_1 hold266 (.A(\instrs[15][6] ),
    .X(net1203));
 sg13g2_dlygate4sd3_1 hold267 (.A(\uart_rx_1.r_Clock_Count[28] ),
    .X(net1204));
 sg13g2_dlygate4sd3_1 hold268 (.A(\datam[0][5] ),
    .X(net1205));
 sg13g2_dlygate4sd3_1 hold269 (.A(\instrs[11][6] ),
    .X(net1206));
 sg13g2_dlygate4sd3_1 hold270 (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[0] ),
    .X(net1207));
 sg13g2_dlygate4sd3_1 hold271 (.A(\datam[4][6] ),
    .X(net1208));
 sg13g2_dlygate4sd3_1 hold272 (.A(\instrs[9][2] ),
    .X(net1209));
 sg13g2_dlygate4sd3_1 hold273 (.A(\instrs[2][2] ),
    .X(net1210));
 sg13g2_dlygate4sd3_1 hold274 (.A(_2513_),
    .X(net1211));
 sg13g2_dlygate4sd3_1 hold275 (.A(\instrs[2][1] ),
    .X(net1212));
 sg13g2_dlygate4sd3_1 hold276 (.A(\instrs[8][2] ),
    .X(net1213));
 sg13g2_dlygate4sd3_1 hold277 (.A(\instrs[14][2] ),
    .X(net1214));
 sg13g2_dlygate4sd3_1 hold278 (.A(\datam[1][3] ),
    .X(net1215));
 sg13g2_dlygate4sd3_1 hold279 (.A(\instrs[14][6] ),
    .X(net1216));
 sg13g2_dlygate4sd3_1 hold280 (.A(\datam[4][7] ),
    .X(net1217));
 sg13g2_dlygate4sd3_1 hold281 (.A(\instrs[9][1] ),
    .X(net1218));
 sg13g2_dlygate4sd3_1 hold282 (.A(\datam[8][5] ),
    .X(net1219));
 sg13g2_dlygate4sd3_1 hold283 (.A(\datam[12][5] ),
    .X(net1220));
 sg13g2_dlygate4sd3_1 hold284 (.A(\instrs[13][2] ),
    .X(net1221));
 sg13g2_dlygate4sd3_1 hold285 (.A(\instrs[0][4] ),
    .X(net1222));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0230_),
    .X(net1223));
 sg13g2_dlygate4sd3_1 hold287 (.A(\instrs[14][1] ),
    .X(net1224));
 sg13g2_dlygate4sd3_1 hold288 (.A(\datam[3][2] ),
    .X(net1225));
 sg13g2_dlygate4sd3_1 hold289 (.A(\datam[1][2] ),
    .X(net1226));
 sg13g2_dlygate4sd3_1 hold290 (.A(\datam[14][4] ),
    .X(net1227));
 sg13g2_dlygate4sd3_1 hold291 (.A(\datam[9][2] ),
    .X(net1228));
 sg13g2_dlygate4sd3_1 hold292 (.A(\instrs[5][2] ),
    .X(net1229));
 sg13g2_dlygate4sd3_1 hold293 (.A(\instrs[13][4] ),
    .X(net1230));
 sg13g2_dlygate4sd3_1 hold294 (.A(\datam[2][2] ),
    .X(net1231));
 sg13g2_dlygate4sd3_1 hold295 (.A(\datam[11][0] ),
    .X(net1232));
 sg13g2_dlygate4sd3_1 hold296 (.A(\datam[10][2] ),
    .X(net1233));
 sg13g2_dlygate4sd3_1 hold297 (.A(\datam[3][4] ),
    .X(net1234));
 sg13g2_dlygate4sd3_1 hold298 (.A(\C1.prog_op ),
    .X(net1235));
 sg13g2_dlygate4sd3_1 hold299 (.A(_0572_),
    .X(net1236));
 sg13g2_dlygate4sd3_1 hold300 (.A(\datam[12][7] ),
    .X(net1237));
 sg13g2_dlygate4sd3_1 hold301 (.A(\datam[15][0] ),
    .X(net1238));
 sg13g2_dlygate4sd3_1 hold302 (.A(\datam[15][4] ),
    .X(net1239));
 sg13g2_dlygate4sd3_1 hold303 (.A(\datam[10][3] ),
    .X(net1240));
 sg13g2_dlygate4sd3_1 hold304 (.A(\datam[11][1] ),
    .X(net1241));
 sg13g2_dlygate4sd3_1 hold305 (.A(\datam[9][3] ),
    .X(net1242));
 sg13g2_dlygate4sd3_1 hold306 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[16] ),
    .X(net1243));
 sg13g2_dlygate4sd3_1 hold307 (.A(_2609_),
    .X(net1244));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0538_),
    .X(net1245));
 sg13g2_dlygate4sd3_1 hold309 (.A(\datam[13][3] ),
    .X(net1246));
 sg13g2_dlygate4sd3_1 hold310 (.A(\datam[13][4] ),
    .X(net1247));
 sg13g2_dlygate4sd3_1 hold311 (.A(\instrs[13][6] ),
    .X(net1248));
 sg13g2_dlygate4sd3_1 hold312 (.A(\datam[0][6] ),
    .X(net1249));
 sg13g2_dlygate4sd3_1 hold313 (.A(\datam[14][0] ),
    .X(net1250));
 sg13g2_dlygate4sd3_1 hold314 (.A(\instrs[10][3] ),
    .X(net1251));
 sg13g2_dlygate4sd3_1 hold315 (.A(\datam[3][1] ),
    .X(net1252));
 sg13g2_dlygate4sd3_1 hold316 (.A(\datam[2][0] ),
    .X(net1253));
 sg13g2_dlygate4sd3_1 hold317 (.A(\instrs[4][1] ),
    .X(net1254));
 sg13g2_dlygate4sd3_1 hold318 (.A(\instrs[2][6] ),
    .X(net1255));
 sg13g2_dlygate4sd3_1 hold319 (.A(\instrs[6][2] ),
    .X(net1256));
 sg13g2_dlygate4sd3_1 hold320 (.A(\instrs[14][3] ),
    .X(net1257));
 sg13g2_dlygate4sd3_1 hold321 (.A(\datam[1][1] ),
    .X(net1258));
 sg13g2_dlygate4sd3_1 hold322 (.A(\datam[1][0] ),
    .X(net1259));
 sg13g2_dlygate4sd3_1 hold323 (.A(\datam[10][4] ),
    .X(net1260));
 sg13g2_dlygate4sd3_1 hold324 (.A(\datam[11][3] ),
    .X(net1261));
 sg13g2_dlygate4sd3_1 hold325 (.A(\uart_rx_1.r_Bit_Index[5] ),
    .X(net1262));
 sg13g2_dlygate4sd3_1 hold326 (.A(\datam[15][1] ),
    .X(net1263));
 sg13g2_dlygate4sd3_1 hold327 (.A(\instrs[4][3] ),
    .X(net1264));
 sg13g2_dlygate4sd3_1 hold328 (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[19] ),
    .X(net1265));
 sg13g2_dlygate4sd3_1 hold329 (.A(_0936_),
    .X(net1266));
 sg13g2_dlygate4sd3_1 hold330 (.A(\FpgaPins_Fpga_GAME_count_speed3_a1[19] ),
    .X(net1267));
 sg13g2_dlygate4sd3_1 hold331 (.A(\instrs[14][4] ),
    .X(net1268));
 sg13g2_dlygate4sd3_1 hold332 (.A(\datam[5][1] ),
    .X(net1269));
 sg13g2_dlygate4sd3_1 hold333 (.A(\datam[6][2] ),
    .X(net1270));
 sg13g2_dlygate4sd3_1 hold334 (.A(\C1.counter2[22] ),
    .X(net1271));
 sg13g2_dlygate4sd3_1 hold335 (.A(_2385_),
    .X(net1272));
 sg13g2_dlygate4sd3_1 hold336 (.A(_0329_),
    .X(net1273));
 sg13g2_dlygate4sd3_1 hold337 (.A(\datam[10][0] ),
    .X(net1274));
 sg13g2_dlygate4sd3_1 hold338 (.A(\datam[8][6] ),
    .X(net1275));
 sg13g2_dlygate4sd3_1 hold339 (.A(\datam[10][1] ),
    .X(net1276));
 sg13g2_dlygate4sd3_1 hold340 (.A(\uart_rx_1.r_Bit_Index[29] ),
    .X(net1277));
 sg13g2_dlygate4sd3_1 hold341 (.A(\datam[3][3] ),
    .X(net1278));
 sg13g2_dlygate4sd3_1 hold342 (.A(\datam[11][4] ),
    .X(net1279));
 sg13g2_dlygate4sd3_1 hold343 (.A(\instrs[2][3] ),
    .X(net1280));
 sg13g2_dlygate4sd3_1 hold344 (.A(\datam[9][0] ),
    .X(net1281));
 sg13g2_dlygate4sd3_1 hold345 (.A(\FpgaPins_Fpga_LIPSI_data_wr_a2[7] ),
    .X(net1282));
 sg13g2_dlygate4sd3_1 hold346 (.A(\datam[4][5] ),
    .X(net1283));
 sg13g2_dlygate4sd3_1 hold347 (.A(\datam[14][1] ),
    .X(net1284));
 sg13g2_dlygate4sd3_1 hold348 (.A(\datam[9][1] ),
    .X(net1285));
 sg13g2_dlygate4sd3_1 hold349 (.A(\C1.counter2[28] ),
    .X(net1286));
 sg13g2_dlygate4sd3_1 hold350 (.A(_2393_),
    .X(net1287));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0335_),
    .X(net1288));
 sg13g2_dlygate4sd3_1 hold352 (.A(\datam[6][3] ),
    .X(net1289));
 sg13g2_dlygate4sd3_1 hold353 (.A(\datam[11][2] ),
    .X(net1290));
 sg13g2_dlygate4sd3_1 hold354 (.A(\datam[5][4] ),
    .X(net1291));
 sg13g2_dlygate4sd3_1 hold355 (.A(\datam[9][4] ),
    .X(net1292));
 sg13g2_dlygate4sd3_1 hold356 (.A(\datam[15][3] ),
    .X(net1293));
 sg13g2_dlygate4sd3_1 hold357 (.A(\instrs[5][3] ),
    .X(net1294));
 sg13g2_dlygate4sd3_1 hold358 (.A(\datam[3][0] ),
    .X(net1295));
 sg13g2_dlygate4sd3_1 hold359 (.A(\datam[7][2] ),
    .X(net1296));
 sg13g2_dlygate4sd3_1 hold360 (.A(\datam[13][2] ),
    .X(net1297));
 sg13g2_dlygate4sd3_1 hold361 (.A(\instrs[1][6] ),
    .X(net1298));
 sg13g2_dlygate4sd3_1 hold362 (.A(\datam[2][4] ),
    .X(net1299));
 sg13g2_dlygate4sd3_1 hold363 (.A(\FpgaPins_Fpga_LIPSI_data_wr_a2[6] ),
    .X(net1300));
 sg13g2_dlygate4sd3_1 hold364 (.A(\instrs[15][1] ),
    .X(net1301));
 sg13g2_dlygate4sd3_1 hold365 (.A(\uart_rx_1.r_Clock_Count[17] ),
    .X(net1302));
 sg13g2_dlygate4sd3_1 hold366 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[18] ),
    .X(net1303));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0992_),
    .X(net1304));
 sg13g2_dlygate4sd3_1 hold368 (.A(\FpgaPins_Fpga_GAME_count_speed1_a1[18] ),
    .X(net1305));
 sg13g2_dlygate4sd3_1 hold369 (.A(\datam[14][3] ),
    .X(net1306));
 sg13g2_dlygate4sd3_1 hold370 (.A(\datam[7][1] ),
    .X(net1307));
 sg13g2_dlygate4sd3_1 hold371 (.A(\datam[6][1] ),
    .X(net1308));
 sg13g2_dlygate4sd3_1 hold372 (.A(\C1.dry_status ),
    .X(net1309));
 sg13g2_dlygate4sd3_1 hold373 (.A(\datam[2][3] ),
    .X(net1310));
 sg13g2_dlygate4sd3_1 hold374 (.A(\datam[14][2] ),
    .X(net1311));
 sg13g2_dlygate4sd3_1 hold375 (.A(\datam[13][0] ),
    .X(net1312));
 sg13g2_dlygate4sd3_1 hold376 (.A(FpgaPins_Fpga_GAME_clk_pulse4_a2),
    .X(net1313));
 sg13g2_dlygate4sd3_1 hold377 (.A(FpgaPins_Fpga_GAME_clk_pulse4_a1),
    .X(net1314));
 sg13g2_dlygate4sd3_1 hold378 (.A(\datam[5][3] ),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold379 (.A(\datam[13][1] ),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold380 (.A(\datam[2][1] ),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold381 (.A(\datam[6][0] ),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold382 (.A(\datam[6][4] ),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold383 (.A(\datam[1][4] ),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold384 (.A(\datam[5][0] ),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold385 (.A(\datam[12][6] ),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold386 (.A(\datam[15][2] ),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold387 (.A(\datam[7][4] ),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold388 (.A(\datam[5][2] ),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold389 (.A(\datam[7][0] ),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold390 (.A(\datam[7][5] ),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold391 (.A(\instrs[4][2] ),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold392 (.A(\instrs[10][6] ),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold393 (.A(\uart_rx_1.r_Bit_Index[28] ),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold394 (.A(\instrs[6][4] ),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold395 (.A(_0368_),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold396 (.A(\C1.pouring ),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold397 (.A(_2644_),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold398 (.A(\instrs[5][4] ),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold399 (.A(\instrs[2][4] ),
    .X(net1336));
 sg13g2_dlygate4sd3_1 hold400 (.A(\datam[15][5] ),
    .X(net1337));
 sg13g2_dlygate4sd3_1 hold401 (.A(\uart_rx_1.r_Clock_Count[30] ),
    .X(net1338));
 sg13g2_dlygate4sd3_1 hold402 (.A(_2892_),
    .X(net1339));
 sg13g2_dlygate4sd3_1 hold403 (.A(_0655_),
    .X(net1340));
 sg13g2_dlygate4sd3_1 hold404 (.A(\instrs[13][1] ),
    .X(net1341));
 sg13g2_dlygate4sd3_1 hold405 (.A(\datam[8][7] ),
    .X(net1342));
 sg13g2_dlygate4sd3_1 hold406 (.A(\datam[7][7] ),
    .X(net1343));
 sg13g2_dlygate4sd3_1 hold407 (.A(\instrs[6][1] ),
    .X(net1344));
 sg13g2_dlygate4sd3_1 hold408 (.A(\datam[7][3] ),
    .X(net1345));
 sg13g2_dlygate4sd3_1 hold409 (.A(_0051_),
    .X(net1346));
 sg13g2_dlygate4sd3_1 hold410 (.A(_0967_),
    .X(net1347));
 sg13g2_dlygate4sd3_1 hold411 (.A(\FpgaPins_Fpga_GAME_count_speed2_a1[14] ),
    .X(net1348));
 sg13g2_dlygate4sd3_1 hold412 (.A(\instrs[1][2] ),
    .X(net1349));
 sg13g2_dlygate4sd3_1 hold413 (.A(_2522_),
    .X(net1350));
 sg13g2_dlygate4sd3_1 hold414 (.A(\uart_rx_1.r_Clock_Count[18] ),
    .X(net1351));
 sg13g2_dlygate4sd3_1 hold415 (.A(\uart_rx_1.r_Rx_Byte[6] ),
    .X(net1352));
 sg13g2_dlygate4sd3_1 hold416 (.A(_2764_),
    .X(net1353));
 sg13g2_dlygate4sd3_1 hold417 (.A(_0591_),
    .X(net1354));
 sg13g2_dlygate4sd3_1 hold418 (.A(\datam[11][6] ),
    .X(net1355));
 sg13g2_dlygate4sd3_1 hold419 (.A(\uart_rx_1.r_Clock_Count[2] ),
    .X(net1356));
 sg13g2_dlygate4sd3_1 hold420 (.A(_2797_),
    .X(net1357));
 sg13g2_dlygate4sd3_1 hold421 (.A(_0627_),
    .X(net1358));
 sg13g2_dlygate4sd3_1 hold422 (.A(\C1.Program[1] ),
    .X(net1359));
 sg13g2_dlygate4sd3_1 hold423 (.A(\instrs[4][4] ),
    .X(net1360));
 sg13g2_dlygate4sd3_1 hold424 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[21] ),
    .X(net1361));
 sg13g2_dlygate4sd3_1 hold425 (.A(\FpgaPins_Fpga_GAME_count_speed1_a1[21] ),
    .X(net1362));
 sg13g2_dlygate4sd3_1 hold426 (.A(\datam[7][6] ),
    .X(net1363));
 sg13g2_dlygate4sd3_1 hold427 (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[6] ),
    .X(net1364));
 sg13g2_dlygate4sd3_1 hold428 (.A(_1109_),
    .X(net1365));
 sg13g2_dlygate4sd3_1 hold429 (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[4] ),
    .X(net1366));
 sg13g2_dlygate4sd3_1 hold430 (.A(_1096_),
    .X(net1367));
 sg13g2_dlygate4sd3_1 hold431 (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[4] ),
    .X(net1368));
 sg13g2_dlygate4sd3_1 hold432 (.A(_1117_),
    .X(net1369));
 sg13g2_dlygate4sd3_1 hold433 (.A(\instrs[15][4] ),
    .X(net1370));
 sg13g2_dlygate4sd3_1 hold434 (.A(_0472_),
    .X(net1371));
 sg13g2_dlygate4sd3_1 hold435 (.A(\datam[15][7] ),
    .X(net1372));
 sg13g2_dlygate4sd3_1 hold436 (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[16] ),
    .X(net1373));
 sg13g2_dlygate4sd3_1 hold437 (.A(_0939_),
    .X(net1374));
 sg13g2_dlygate4sd3_1 hold438 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[6] ),
    .X(net1375));
 sg13g2_dlygate4sd3_1 hold439 (.A(_2591_),
    .X(net1376));
 sg13g2_dlygate4sd3_1 hold440 (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[9] ),
    .X(net1377));
 sg13g2_dlygate4sd3_1 hold441 (.A(_1120_),
    .X(net1378));
 sg13g2_dlygate4sd3_1 hold442 (.A(\C1.waiting ),
    .X(net1379));
 sg13g2_dlygate4sd3_1 hold443 (.A(_0571_),
    .X(net1380));
 sg13g2_dlygate4sd3_1 hold444 (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[4] ),
    .X(net1381));
 sg13g2_dlygate4sd3_1 hold445 (.A(_1108_),
    .X(net1382));
 sg13g2_dlygate4sd3_1 hold446 (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[8] ),
    .X(net1383));
 sg13g2_dlygate4sd3_1 hold447 (.A(_0930_),
    .X(net1384));
 sg13g2_dlygate4sd3_1 hold448 (.A(_0050_),
    .X(net1385));
 sg13g2_dlygate4sd3_1 hold449 (.A(_1112_),
    .X(net1386));
 sg13g2_dlygate4sd3_1 hold450 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[15] ),
    .X(net1387));
 sg13g2_dlygate4sd3_1 hold451 (.A(_0537_),
    .X(net1388));
 sg13g2_dlygate4sd3_1 hold452 (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[6] ),
    .X(net1389));
 sg13g2_dlygate4sd3_1 hold453 (.A(_1097_),
    .X(net1390));
 sg13g2_dlygate4sd3_1 hold454 (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[5] ),
    .X(net1391));
 sg13g2_dlygate4sd3_1 hold455 (.A(\instrs[8][3] ),
    .X(net1392));
 sg13g2_dlygate4sd3_1 hold456 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[6] ),
    .X(net1393));
 sg13g2_dlygate4sd3_1 hold457 (.A(_1129_),
    .X(net1394));
 sg13g2_dlygate4sd3_1 hold458 (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[12] ),
    .X(net1395));
 sg13g2_dlygate4sd3_1 hold459 (.A(\FpgaPins_Fpga_GAME_count_speed3_a1[12] ),
    .X(net1396));
 sg13g2_dlygate4sd3_1 hold460 (.A(\uart_rx_1.r_Clock_Count[29] ),
    .X(net1397));
 sg13g2_dlygate4sd3_1 hold461 (.A(_0654_),
    .X(net1398));
 sg13g2_dlygate4sd3_1 hold462 (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[3] ),
    .X(net1399));
 sg13g2_dlygate4sd3_1 hold463 (.A(\uart_rx_1.r_Bit_Index[12] ),
    .X(net1400));
 sg13g2_dlygate4sd3_1 hold464 (.A(\datam[5][5] ),
    .X(net1401));
 sg13g2_dlygate4sd3_1 hold465 (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[11] ),
    .X(net1402));
 sg13g2_dlygate4sd3_1 hold466 (.A(_1122_),
    .X(net1403));
 sg13g2_dlygate4sd3_1 hold467 (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[5] ),
    .X(net1404));
 sg13g2_dlygate4sd3_1 hold468 (.A(_0049_),
    .X(net1405));
 sg13g2_dlygate4sd3_1 hold469 (.A(_1103_),
    .X(net1406));
 sg13g2_dlygate4sd3_1 hold470 (.A(\instrs[9][6] ),
    .X(net1407));
 sg13g2_dlygate4sd3_1 hold471 (.A(\uart_rx_1.r_SM_Main[2] ),
    .X(net1408));
 sg13g2_dlygate4sd3_1 hold472 (.A(_0659_),
    .X(net1409));
 sg13g2_dlygate4sd3_1 hold473 (.A(\datam[5][6] ),
    .X(net1410));
 sg13g2_dlygate4sd3_1 hold474 (.A(\C1.heating ),
    .X(net1411));
 sg13g2_dlygate4sd3_1 hold475 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[23] ),
    .X(net1412));
 sg13g2_dlygate4sd3_1 hold476 (.A(_0545_),
    .X(net1413));
 sg13g2_dlygate4sd3_1 hold477 (.A(\C1.rinse_status ),
    .X(net1414));
 sg13g2_dlygate4sd3_1 hold478 (.A(_2654_),
    .X(net1415));
 sg13g2_dlygate4sd3_1 hold479 (.A(\datam[3][5] ),
    .X(net1416));
 sg13g2_dlygate4sd3_1 hold480 (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[7] ),
    .X(net1417));
 sg13g2_dlygate4sd3_1 hold481 (.A(\uart_rx_1.r_Bit_Index[4] ),
    .X(net1418));
 sg13g2_dlygate4sd3_1 hold482 (.A(\uart_rx_1.r_Rx_Byte[7] ),
    .X(net1419));
 sg13g2_dlygate4sd3_1 hold483 (.A(_2766_),
    .X(net1420));
 sg13g2_dlygate4sd3_1 hold484 (.A(_0592_),
    .X(net1421));
 sg13g2_dlygate4sd3_1 hold485 (.A(_0052_),
    .X(net1422));
 sg13g2_dlygate4sd3_1 hold486 (.A(_0980_),
    .X(net1423));
 sg13g2_dlygate4sd3_1 hold487 (.A(\C1.Program[0] ),
    .X(net1424));
 sg13g2_dlygate4sd3_1 hold488 (.A(\datam[11][5] ),
    .X(net1425));
 sg13g2_dlygate4sd3_1 hold489 (.A(\datam[14][6] ),
    .X(net1426));
 sg13g2_dlygate4sd3_1 hold490 (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[17] ),
    .X(net1427));
 sg13g2_dlygate4sd3_1 hold491 (.A(_1113_),
    .X(net1428));
 sg13g2_dlygate4sd3_1 hold492 (.A(\uart_rx_1.r_Clock_Count[4] ),
    .X(net1429));
 sg13g2_dlygate4sd3_1 hold493 (.A(_2801_),
    .X(net1430));
 sg13g2_dlygate4sd3_1 hold494 (.A(\datam[15][6] ),
    .X(net1431));
 sg13g2_dlygate4sd3_1 hold495 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[2] ),
    .X(net1432));
 sg13g2_dlygate4sd3_1 hold496 (.A(_1125_),
    .X(net1433));
 sg13g2_dlygate4sd3_1 hold497 (.A(\FpgaPins_Fpga_GAME_count_speed1_a1[2] ),
    .X(net1434));
 sg13g2_dlygate4sd3_1 hold498 (.A(_0202_),
    .X(net1435));
 sg13g2_dlygate4sd3_1 hold499 (.A(_2776_),
    .X(net1436));
 sg13g2_dlygate4sd3_1 hold500 (.A(_2777_),
    .X(net1437));
 sg13g2_dlygate4sd3_1 hold501 (.A(\datam[14][5] ),
    .X(net1438));
 sg13g2_dlygate4sd3_1 hold502 (.A(\datam[11][7] ),
    .X(net1439));
 sg13g2_dlygate4sd3_1 hold503 (.A(\C1.max_count[6] ),
    .X(net1440));
 sg13g2_dlygate4sd3_1 hold504 (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[10] ),
    .X(net1441));
 sg13g2_dlygate4sd3_1 hold505 (.A(\datam[1][6] ),
    .X(net1442));
 sg13g2_dlygate4sd3_1 hold506 (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[17] ),
    .X(net1443));
 sg13g2_dlygate4sd3_1 hold507 (.A(_1123_),
    .X(net1444));
 sg13g2_dlygate4sd3_1 hold508 (.A(\FpgaPins_Fpga_GAME_count_speed2_a1[17] ),
    .X(net1445));
 sg13g2_dlygate4sd3_1 hold509 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[3] ),
    .X(net1446));
 sg13g2_dlygate4sd3_1 hold510 (.A(\datam[13][6] ),
    .X(net1447));
 sg13g2_dlygate4sd3_1 hold511 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[17] ),
    .X(net1448));
 sg13g2_dlygate4sd3_1 hold512 (.A(_2611_),
    .X(net1449));
 sg13g2_dlygate4sd3_1 hold513 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[4] ),
    .X(net1450));
 sg13g2_dlygate4sd3_1 hold514 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[18] ),
    .X(net1451));
 sg13g2_dlygate4sd3_1 hold515 (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[3] ),
    .X(net1452));
 sg13g2_dlygate4sd3_1 hold516 (.A(_1116_),
    .X(net1453));
 sg13g2_dlygate4sd3_1 hold517 (.A(\datam[10][7] ),
    .X(net1454));
 sg13g2_dlygate4sd3_1 hold518 (.A(\datam[10][6] ),
    .X(net1455));
 sg13g2_dlygate4sd3_1 hold519 (.A(\datam[9][6] ),
    .X(net1456));
 sg13g2_dlygate4sd3_1 hold520 (.A(_0087_),
    .X(net1457));
 sg13g2_dlygate4sd3_1 hold521 (.A(_1193_),
    .X(net1458));
 sg13g2_dlygate4sd3_1 hold522 (.A(_0007_),
    .X(net1459));
 sg13g2_dlygate4sd3_1 hold523 (.A(\datam[10][5] ),
    .X(net1460));
 sg13g2_dlygate4sd3_1 hold524 (.A(\datam[3][7] ),
    .X(net1461));
 sg13g2_dlygate4sd3_1 hold525 (.A(\uart_rx_1.r_Clock_Count[24] ),
    .X(net1462));
 sg13g2_dlygate4sd3_1 hold526 (.A(_2872_),
    .X(net1463));
 sg13g2_dlygate4sd3_1 hold527 (.A(\datam[6][6] ),
    .X(net1464));
 sg13g2_dlygate4sd3_1 hold528 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[17] ),
    .X(net1465));
 sg13g2_dlygate4sd3_1 hold529 (.A(\FpgaPins_Fpga_GAME_count_speed1_a1[17] ),
    .X(net1466));
 sg13g2_dlygate4sd3_1 hold530 (.A(\datam[5][7] ),
    .X(net1467));
 sg13g2_dlygate4sd3_1 hold531 (.A(\datam[9][7] ),
    .X(net1468));
 sg13g2_dlygate4sd3_1 hold532 (.A(\datam[9][5] ),
    .X(net1469));
 sg13g2_dlygate4sd3_1 hold533 (.A(\datam[1][7] ),
    .X(net1470));
 sg13g2_dlygate4sd3_1 hold534 (.A(\uart_rx_1.r_Clock_Count[9] ),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold535 (.A(_0634_),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold536 (.A(\C1.max_count[9] ),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold537 (.A(\datam[2][6] ),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold538 (.A(\datam[1][5] ),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold539 (.A(\datam[2][5] ),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold540 (.A(\datam[2][7] ),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold541 (.A(FpgaPins_Fpga_GAME_clk_pulse2_a2),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold542 (.A(FpgaPins_Fpga_GAME_clk_pulse2_a1),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold543 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[3] ),
    .X(net1480));
 sg13g2_dlygate4sd3_1 hold544 (.A(_2585_),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold545 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[5] ),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold546 (.A(_2589_),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold547 (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[7] ),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold548 (.A(_0970_),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold549 (.A(\datam[3][6] ),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold550 (.A(\uart_rx_1.r_Clock_Count[23] ),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold551 (.A(\datam[6][5] ),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold552 (.A(\C1.max_count[2] ),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold553 (.A(\datam[14][7] ),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold554 (.A(\datam[13][7] ),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold555 (.A(FpgaPins_Fpga_GAME_reset_a2),
    .X(net1492));
 sg13g2_dlygate4sd3_1 hold556 (.A(_0354_),
    .X(net1493));
 sg13g2_dlygate4sd3_1 hold557 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[5] ),
    .X(net1494));
 sg13g2_dlygate4sd3_1 hold558 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[14] ),
    .X(net1495));
 sg13g2_dlygate4sd3_1 hold559 (.A(_2606_),
    .X(net1496));
 sg13g2_dlygate4sd3_1 hold560 (.A(_0536_),
    .X(net1497));
 sg13g2_dlygate4sd3_1 hold561 (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[15] ),
    .X(net1498));
 sg13g2_dlygate4sd3_1 hold562 (.A(\FpgaPins_Fpga_GAME_count_speed4_a1[15] ),
    .X(net1499));
 sg13g2_dlygate4sd3_1 hold563 (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[8] ),
    .X(net1500));
 sg13g2_dlygate4sd3_1 hold564 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[4] ),
    .X(net1501));
 sg13g2_dlygate4sd3_1 hold565 (.A(\datam[6][7] ),
    .X(net1502));
 sg13g2_dlygate4sd3_1 hold566 (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[17] ),
    .X(net1503));
 sg13g2_dlygate4sd3_1 hold567 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[7] ),
    .X(net1504));
 sg13g2_dlygate4sd3_1 hold568 (.A(\uart_rx_1.r_Clock_Count[6] ),
    .X(net1505));
 sg13g2_dlygate4sd3_1 hold569 (.A(_2808_),
    .X(net1506));
 sg13g2_dlygate4sd3_1 hold570 (.A(_0631_),
    .X(net1507));
 sg13g2_dlygate4sd3_1 hold571 (.A(\uart_rx_1.r_Clock_Count[0] ),
    .X(net1508));
 sg13g2_dlygate4sd3_1 hold572 (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[16] ),
    .X(net1509));
 sg13g2_dlygate4sd3_1 hold573 (.A(_0978_),
    .X(net1510));
 sg13g2_dlygate4sd3_1 hold574 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[19] ),
    .X(net1511));
 sg13g2_dlygate4sd3_1 hold575 (.A(\C1.max_count[1] ),
    .X(net1512));
 sg13g2_dlygate4sd3_1 hold576 (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[3] ),
    .X(net1513));
 sg13g2_dlygate4sd3_1 hold577 (.A(_1095_),
    .X(net1514));
 sg13g2_dlygate4sd3_1 hold578 (.A(\uart_rx_1.r_Rx_Byte[5] ),
    .X(net1515));
 sg13g2_dlygate4sd3_1 hold579 (.A(_2763_),
    .X(net1516));
 sg13g2_dlygate4sd3_1 hold580 (.A(_0590_),
    .X(net1517));
 sg13g2_dlygate4sd3_1 hold581 (.A(\C1.max_count[4] ),
    .X(net1518));
 sg13g2_dlygate4sd3_1 hold582 (.A(\uart_rx_1.r_Bit_Index[31] ),
    .X(net1519));
 sg13g2_dlygate4sd3_1 hold583 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[20] ),
    .X(net1520));
 sg13g2_dlygate4sd3_1 hold584 (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[6] ),
    .X(net1521));
 sg13g2_dlygate4sd3_1 hold585 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[23] ),
    .X(net1522));
 sg13g2_dlygate4sd3_1 hold586 (.A(_1140_),
    .X(net1523));
 sg13g2_dlygate4sd3_1 hold587 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[9] ),
    .X(net1524));
 sg13g2_dlygate4sd3_1 hold588 (.A(_2596_),
    .X(net1525));
 sg13g2_dlygate4sd3_1 hold589 (.A(_0531_),
    .X(net1526));
 sg13g2_dlygate4sd3_1 hold590 (.A(_0019_),
    .X(net1527));
 sg13g2_dlygate4sd3_1 hold591 (.A(FpgaPins_Fpga_GAME_clk_pulse1_a1),
    .X(net1528));
 sg13g2_dlygate4sd3_1 hold592 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[12] ),
    .X(net1529));
 sg13g2_dlygate4sd3_1 hold593 (.A(_2602_),
    .X(net1530));
 sg13g2_dlygate4sd3_1 hold594 (.A(_0534_),
    .X(net1531));
 sg13g2_dlygate4sd3_1 hold595 (.A(\C1.counter_status[1] ),
    .X(net1532));
 sg13g2_dlygate4sd3_1 hold596 (.A(_1270_),
    .X(net1533));
 sg13g2_dlygate4sd3_1 hold597 (.A(_0006_),
    .X(net1534));
 sg13g2_dlygate4sd3_1 hold598 (.A(\uart_rx_1.r_Bit_Index[3] ),
    .X(net1535));
 sg13g2_dlygate4sd3_1 hold599 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[20] ),
    .X(net1536));
 sg13g2_dlygate4sd3_1 hold600 (.A(_2617_),
    .X(net1537));
 sg13g2_dlygate4sd3_1 hold601 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[1] ),
    .X(net1538));
 sg13g2_dlygate4sd3_1 hold602 (.A(_2581_),
    .X(net1539));
 sg13g2_dlygate4sd3_1 hold603 (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[15] ),
    .X(net1540));
 sg13g2_dlygate4sd3_1 hold604 (.A(_0966_),
    .X(net1541));
 sg13g2_dlygate4sd3_1 hold605 (.A(\C1.max_count[7] ),
    .X(net1542));
 sg13g2_dlygate4sd3_1 hold606 (.A(FpgaPins_Fpga_UART_is_enter_a2),
    .X(net1543));
 sg13g2_dlygate4sd3_1 hold607 (.A(_1941_),
    .X(net1544));
 sg13g2_dlygate4sd3_1 hold608 (.A(\C1.counter2[0] ),
    .X(net1545));
 sg13g2_dlygate4sd3_1 hold609 (.A(\C1.next_state_var[1] ),
    .X(net1546));
 sg13g2_dlygate4sd3_1 hold610 (.A(_0004_),
    .X(net1547));
 sg13g2_dlygate4sd3_1 hold611 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[19] ),
    .X(net1548));
 sg13g2_dlygate4sd3_1 hold612 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[16] ),
    .X(net1549));
 sg13g2_dlygate4sd3_1 hold613 (.A(_1136_),
    .X(net1550));
 sg13g2_dlygate4sd3_1 hold614 (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[5] ),
    .X(net1551));
 sg13g2_dlygate4sd3_1 hold615 (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[10] ),
    .X(net1552));
 sg13g2_dlygate4sd3_1 hold616 (.A(_1111_),
    .X(net1553));
 sg13g2_dlygate4sd3_1 hold617 (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[11] ),
    .X(net1554));
 sg13g2_dlygate4sd3_1 hold618 (.A(_1101_),
    .X(net1555));
 sg13g2_dlygate4sd3_1 hold619 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[9] ),
    .X(net1556));
 sg13g2_dlygate4sd3_1 hold620 (.A(_1131_),
    .X(net1557));
 sg13g2_dlygate4sd3_1 hold621 (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[9] ),
    .X(net1558));
 sg13g2_dlygate4sd3_1 hold622 (.A(\FpgaPins_Fpga_GAME_count_speed3_a1[9] ),
    .X(net1559));
 sg13g2_dlygate4sd3_1 hold623 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[14] ),
    .X(net1560));
 sg13g2_dlygate4sd3_1 hold624 (.A(_1135_),
    .X(net1561));
 sg13g2_dlygate4sd3_1 hold625 (.A(\FpgaPins_Fpga_GAME_led_output_a3[0] ),
    .X(net1562));
 sg13g2_dlygate4sd3_1 hold626 (.A(\C1.max_count[11] ),
    .X(net1563));
 sg13g2_dlygate4sd3_1 hold627 (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[12] ),
    .X(net1564));
 sg13g2_dlygate4sd3_1 hold628 (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[12] ),
    .X(net1565));
 sg13g2_dlygate4sd3_1 hold629 (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[13] ),
    .X(net1566));
 sg13g2_dlygate4sd3_1 hold630 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[22] ),
    .X(net1567));
 sg13g2_dlygate4sd3_1 hold631 (.A(_2621_),
    .X(net1568));
 sg13g2_dlygate4sd3_1 hold632 (.A(\C1.dura_op ),
    .X(net1569));
 sg13g2_dlygate4sd3_1 hold633 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[15] ),
    .X(net1570));
 sg13g2_dlygate4sd3_1 hold634 (.A(\FpgaPins_Fpga_GAME_led_output_a3[7] ),
    .X(net1571));
 sg13g2_dlygate4sd3_1 hold635 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[11] ),
    .X(net1572));
 sg13g2_dlygate4sd3_1 hold636 (.A(_1132_),
    .X(net1573));
 sg13g2_dlygate4sd3_1 hold637 (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[9] ),
    .X(net1574));
 sg13g2_dlygate4sd3_1 hold638 (.A(_1099_),
    .X(net1575));
 sg13g2_dlygate4sd3_1 hold639 (.A(\C1.counter2[19] ),
    .X(net1576));
 sg13g2_dlygate4sd3_1 hold640 (.A(_2561_),
    .X(net1577));
 sg13g2_dlygate4sd3_1 hold641 (.A(\FpgaPins_Fpga_GAME_speed_level_a2[2] ),
    .X(net1578));
 sg13g2_dlygate4sd3_1 hold642 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[8] ),
    .X(net1579));
 sg13g2_dlygate4sd3_1 hold643 (.A(_1130_),
    .X(net1580));
 sg13g2_dlygate4sd3_1 hold644 (.A(\FpgaPins_Fpga_GAME_score_a2[1] ),
    .X(net1581));
 sg13g2_dlygate4sd3_1 hold645 (.A(\uart_rx_1.r_Clock_Count[3] ),
    .X(net1582));
 sg13g2_dlygate4sd3_1 hold646 (.A(_2800_),
    .X(net1583));
 sg13g2_dlygate4sd3_1 hold647 (.A(\C1.counter2[13] ),
    .X(net1584));
 sg13g2_dlygate4sd3_1 hold648 (.A(_2553_),
    .X(net1585));
 sg13g2_dlygate4sd3_1 hold649 (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[18] ),
    .X(net1586));
 sg13g2_dlygate4sd3_1 hold650 (.A(\FpgaPins_Fpga_UART_dptr_a2[1] ),
    .X(net1587));
 sg13g2_dlygate4sd3_1 hold651 (.A(_2400_),
    .X(net1588));
 sg13g2_dlygate4sd3_1 hold652 (.A(\FpgaPins_Fpga_GAME_win_a2[2] ),
    .X(net1589));
 sg13g2_dlygate4sd3_1 hold653 (.A(_1214_),
    .X(net1590));
 sg13g2_dlygate4sd3_1 hold654 (.A(\C1.counter2[16] ),
    .X(net1591));
 sg13g2_dlygate4sd3_1 hold655 (.A(_2557_),
    .X(net1592));
 sg13g2_dlygate4sd3_1 hold656 (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[1] ),
    .X(net1593));
 sg13g2_dlygate4sd3_1 hold657 (.A(\C1.next_state_var[3] ),
    .X(net1594));
 sg13g2_dlygate4sd3_1 hold658 (.A(\uart_rx_1.r_Rx_Byte[4] ),
    .X(net1595));
 sg13g2_dlygate4sd3_1 hold659 (.A(_0589_),
    .X(net1596));
 sg13g2_dlygate4sd3_1 hold660 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[21] ),
    .X(net1597));
 sg13g2_dlygate4sd3_1 hold661 (.A(\uart_rx_1.r_Bit_Index[0] ),
    .X(net1598));
 sg13g2_dlygate4sd3_1 hold662 (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[13] ),
    .X(net1599));
 sg13g2_dlygate4sd3_1 hold663 (.A(\C1.counter2[6] ),
    .X(net1600));
 sg13g2_dlygate4sd3_1 hold664 (.A(_2544_),
    .X(net1601));
 sg13g2_dlygate4sd3_1 hold665 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[10] ),
    .X(net1602));
 sg13g2_dlygate4sd3_1 hold666 (.A(_2598_),
    .X(net1603));
 sg13g2_dlygate4sd3_1 hold667 (.A(\C1.counter2[4] ),
    .X(net1604));
 sg13g2_dlygate4sd3_1 hold668 (.A(_2542_),
    .X(net1605));
 sg13g2_dlygate4sd3_1 hold669 (.A(\C1.max_count[3] ),
    .X(net1606));
 sg13g2_dlygate4sd3_1 hold670 (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[8] ),
    .X(net1607));
 sg13g2_dlygate4sd3_1 hold671 (.A(\uart_rx_1.r_Bit_Index[1] ),
    .X(net1608));
 sg13g2_dlygate4sd3_1 hold672 (.A(\FpgaPins_Fpga_GAME_count_speed2_a2[18] ),
    .X(net1609));
 sg13g2_dlygate4sd3_1 hold673 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[13] ),
    .X(net1610));
 sg13g2_dlygate4sd3_1 hold674 (.A(_1134_),
    .X(net1611));
 sg13g2_dlygate4sd3_1 hold675 (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[1] ),
    .X(net1612));
 sg13g2_dlygate4sd3_1 hold676 (.A(\C1.counter2[29] ),
    .X(net1613));
 sg13g2_dlygate4sd3_1 hold677 (.A(_2394_),
    .X(net1614));
 sg13g2_dlygate4sd3_1 hold678 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[10] ),
    .X(net1615));
 sg13g2_dlygate4sd3_1 hold679 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[1] ),
    .X(net1616));
 sg13g2_dlygate4sd3_1 hold680 (.A(\C1.counter2[23] ),
    .X(net1617));
 sg13g2_dlygate4sd3_1 hold681 (.A(_2386_),
    .X(net1618));
 sg13g2_dlygate4sd3_1 hold682 (.A(\uart_rx_1.r_Clock_Count[7] ),
    .X(net1619));
 sg13g2_dlygate4sd3_1 hold683 (.A(_2810_),
    .X(net1620));
 sg13g2_dlygate4sd3_1 hold684 (.A(\FpgaPins_Fpga_GAME_count_speed4_a2[10] ),
    .X(net1621));
 sg13g2_dlygate4sd3_1 hold685 (.A(\uart_rx_1.r_Clock_Count[5] ),
    .X(net1622));
 sg13g2_dlygate4sd3_1 hold686 (.A(_0630_),
    .X(net1623));
 sg13g2_dlygate4sd3_1 hold687 (.A(\C1.counter2[10] ),
    .X(net1624));
 sg13g2_dlygate4sd3_1 hold688 (.A(_2549_),
    .X(net1625));
 sg13g2_dlygate4sd3_1 hold689 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[12] ),
    .X(net1626));
 sg13g2_dlygate4sd3_1 hold690 (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[11] ),
    .X(net1627));
 sg13g2_dlygate4sd3_1 hold691 (.A(\uart_rx_1.r_Rx_Byte[3] ),
    .X(net1628));
 sg13g2_dlygate4sd3_1 hold692 (.A(_2754_),
    .X(net1629));
 sg13g2_dlygate4sd3_1 hold693 (.A(_0588_),
    .X(net1630));
 sg13g2_dlygate4sd3_1 hold694 (.A(\C1.max_count[8] ),
    .X(net1631));
 sg13g2_dlygate4sd3_1 hold695 (.A(\C1.counter2[26] ),
    .X(net1632));
 sg13g2_dlygate4sd3_1 hold696 (.A(_2390_),
    .X(net1633));
 sg13g2_dlygate4sd3_1 hold697 (.A(\C1.counter2[5] ),
    .X(net1634));
 sg13g2_dlygate4sd3_1 hold698 (.A(\C1.max_count[10] ),
    .X(net1635));
 sg13g2_dlygate4sd3_1 hold699 (.A(\FpgaPins_Fpga_GAME_win_a2[1] ),
    .X(net1636));
 sg13g2_dlygate4sd3_1 hold700 (.A(\uart_rx_1.r_SM_Main[0] ),
    .X(net1637));
 sg13g2_dlygate4sd3_1 hold701 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[8] ),
    .X(net1638));
 sg13g2_dlygate4sd3_1 hold702 (.A(_2595_),
    .X(net1639));
 sg13g2_dlygate4sd3_1 hold703 (.A(_0118_),
    .X(net1640));
 sg13g2_dlygate4sd3_1 hold704 (.A(_1318_),
    .X(net1641));
 sg13g2_dlygate4sd3_1 hold705 (.A(_1327_),
    .X(net1642));
 sg13g2_dlygate4sd3_1 hold706 (.A(\FpgaPins_Fpga_FSM_data_a1[0] ),
    .X(net1643));
 sg13g2_dlygate4sd3_1 hold707 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[11] ),
    .X(net1644));
 sg13g2_dlygate4sd3_1 hold708 (.A(_2601_),
    .X(net1645));
 sg13g2_dlygate4sd3_1 hold709 (.A(\C1.max_count[5] ),
    .X(net1646));
 sg13g2_dlygate4sd3_1 hold710 (.A(\C1.counter2[3] ),
    .X(net1647));
 sg13g2_dlygate4sd3_1 hold711 (.A(_2541_),
    .X(net1648));
 sg13g2_dlygate4sd3_1 hold712 (.A(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[1] ),
    .X(net1649));
 sg13g2_dlygate4sd3_1 hold713 (.A(_2379_),
    .X(net1650));
 sg13g2_dlygate4sd3_1 hold714 (.A(\C1.counter2[24] ),
    .X(net1651));
 sg13g2_dlygate4sd3_1 hold715 (.A(_1772_),
    .X(net1652));
 sg13g2_dlygate4sd3_1 hold716 (.A(FpgaPins_Fpga_LIPSI_c_a2),
    .X(net1653));
 sg13g2_dlygate4sd3_1 hold717 (.A(\C1.timer[1] ),
    .X(net1654));
 sg13g2_dlygate4sd3_1 hold718 (.A(\uart_rx_1.r_Clock_Count[11] ),
    .X(net1655));
 sg13g2_dlygate4sd3_1 hold719 (.A(\C1.counter2[30] ),
    .X(net1656));
 sg13g2_dlygate4sd3_1 hold720 (.A(_1776_),
    .X(net1657));
 sg13g2_dlygate4sd3_1 hold721 (.A(\C1.counter2[27] ),
    .X(net1658));
 sg13g2_dlygate4sd3_1 hold722 (.A(\uart_rx_1.r_Rx_DV ),
    .X(net1659));
 sg13g2_dlygate4sd3_1 hold723 (.A(_0584_),
    .X(net1660));
 sg13g2_dlygate4sd3_1 hold724 (.A(\uart_rx_1.r_Clock_Count[1] ),
    .X(net1661));
 sg13g2_dlygate4sd3_1 hold725 (.A(\uart_rx_1.r_SM_Main[1] ),
    .X(net1662));
 sg13g2_dlygate4sd3_1 hold726 (.A(_0658_),
    .X(net1663));
 sg13g2_dlygate4sd3_1 hold727 (.A(FpgaPins_Fpga_UART_first_byte_a2),
    .X(net1664));
 sg13g2_dlygate4sd3_1 hold728 (.A(_0085_),
    .X(net1665));
 sg13g2_dlygate4sd3_1 hold729 (.A(_1906_),
    .X(net1666));
 sg13g2_dlygate4sd3_1 hold730 (.A(\uart_rx_1.r_Rx_Byte[2] ),
    .X(net1667));
 sg13g2_dlygate4sd3_1 hold731 (.A(_0587_),
    .X(net1668));
 sg13g2_dlygate4sd3_1 hold732 (.A(FpgaPins_Fpga_GAME_clk_pulse1_a2),
    .X(net1669));
 sg13g2_dlygate4sd3_1 hold733 (.A(\FpgaPins_Fpga_GAME_led_output_a1[2] ),
    .X(net1670));
 sg13g2_dlygate4sd3_1 hold734 (.A(_0086_),
    .X(net1671));
 sg13g2_dlygate4sd3_1 hold735 (.A(\C1.counter2[20] ),
    .X(net1672));
 sg13g2_dlygate4sd3_1 hold736 (.A(_2562_),
    .X(net1673));
 sg13g2_dlygate4sd3_1 hold737 (.A(\uart_rx_1.r_Rx_Byte[0] ),
    .X(net1674));
 sg13g2_dlygate4sd3_1 hold738 (.A(_1932_),
    .X(net1675));
 sg13g2_dlygate4sd3_1 hold739 (.A(FpgaPins_Fpga_UART_is_enter_a1),
    .X(net1676));
 sg13g2_dlygate4sd3_1 hold740 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[22] ),
    .X(net1677));
 sg13g2_dlygate4sd3_1 hold741 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[15] ),
    .X(net1678));
 sg13g2_dlygate4sd3_1 hold742 (.A(_2436_),
    .X(net1679));
 sg13g2_dlygate4sd3_1 hold743 (.A(_2438_),
    .X(net1680));
 sg13g2_dlygate4sd3_1 hold744 (.A(\C1.counter2[11] ),
    .X(net1681));
 sg13g2_dlygate4sd3_1 hold745 (.A(_2550_),
    .X(net1682));
 sg13g2_dlygate4sd3_1 hold746 (.A(\C1.counter2[8] ),
    .X(net1683));
 sg13g2_dlygate4sd3_1 hold747 (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[15] ),
    .X(net1684));
 sg13g2_dlygate4sd3_1 hold748 (.A(\C1.counter2[7] ),
    .X(net1685));
 sg13g2_dlygate4sd3_1 hold749 (.A(\FpgaPins_Fpga_GAME_speed_level_a2[3] ),
    .X(net1686));
 sg13g2_dlygate4sd3_1 hold750 (.A(_0018_),
    .X(net1687));
 sg13g2_dlygate4sd3_1 hold751 (.A(\FpgaPins_Fpga_GAME_led_output_a1[4] ),
    .X(net1688));
 sg13g2_dlygate4sd3_1 hold752 (.A(\C1.counter2[1] ),
    .X(net1689));
 sg13g2_dlygate4sd3_1 hold753 (.A(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[3] ),
    .X(net1690));
 sg13g2_dlygate4sd3_1 hold754 (.A(\FpgaPins_Fpga_GAME_score_a4[5] ),
    .X(net1691));
 sg13g2_dlygate4sd3_1 hold755 (.A(\C1.next_state_var[2] ),
    .X(net1692));
 sg13g2_dlygate4sd3_1 hold756 (.A(_0005_),
    .X(net1693));
 sg13g2_dlygate4sd3_1 hold757 (.A(\C1.counter2[14] ),
    .X(net1694));
 sg13g2_dlygate4sd3_1 hold758 (.A(_2554_),
    .X(net1695));
 sg13g2_dlygate4sd3_1 hold759 (.A(\C1.counter2[17] ),
    .X(net1696));
 sg13g2_dlygate4sd3_1 hold760 (.A(_2558_),
    .X(net1697));
 sg13g2_dlygate4sd3_1 hold761 (.A(\uart_rx_1.r_Rx_Byte[1] ),
    .X(net1698));
 sg13g2_dlygate4sd3_1 hold762 (.A(_2749_),
    .X(net1699));
 sg13g2_dlygate4sd3_1 hold763 (.A(\C1.counter1[10] ),
    .X(net1700));
 sg13g2_dlygate4sd3_1 hold764 (.A(_1801_),
    .X(net1701));
 sg13g2_dlygate4sd3_1 hold765 (.A(\C1.counter2[18] ),
    .X(net1702));
 sg13g2_dlygate4sd3_1 hold766 (.A(_1768_),
    .X(net1703));
 sg13g2_dlygate4sd3_1 hold767 (.A(\C1.counter2[21] ),
    .X(net1704));
 sg13g2_dlygate4sd3_1 hold768 (.A(_2564_),
    .X(net1705));
 sg13g2_dlygate4sd3_1 hold769 (.A(\C1.counter2[9] ),
    .X(net1706));
 sg13g2_dlygate4sd3_1 hold770 (.A(\C1.next_state_var[0] ),
    .X(net1707));
 sg13g2_dlygate4sd3_1 hold771 (.A(_2123_),
    .X(net1708));
 sg13g2_dlygate4sd3_1 hold772 (.A(_2242_),
    .X(net1709));
 sg13g2_dlygate4sd3_1 hold773 (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[7] ),
    .X(net1710));
 sg13g2_dlygate4sd3_1 hold774 (.A(_0931_),
    .X(net1711));
 sg13g2_dlygate4sd3_1 hold775 (.A(\C1.counter2[12] ),
    .X(net1712));
 sg13g2_dlygate4sd3_1 hold776 (.A(_1764_),
    .X(net1713));
 sg13g2_dlygate4sd3_1 hold777 (.A(_2552_),
    .X(net1714));
 sg13g2_dlygate4sd3_1 hold778 (.A(\C1.counter2[15] ),
    .X(net1715));
 sg13g2_dlygate4sd3_1 hold779 (.A(_1766_),
    .X(net1716));
 sg13g2_dlygate4sd3_1 hold780 (.A(_2556_),
    .X(net1717));
 sg13g2_dlygate4sd3_1 hold781 (.A(_0168_),
    .X(net1718));
 sg13g2_dlygate4sd3_1 hold782 (.A(_1491_),
    .X(net1719));
 sg13g2_dlygate4sd3_1 hold783 (.A(\FpgaPins_Fpga_GAME_speed_level_a2[1] ),
    .X(net1720));
 sg13g2_dlygate4sd3_1 hold784 (.A(\FpgaPins_Fpga_GAME_count_speed1_a2[7] ),
    .X(net1721));
 sg13g2_dlygate4sd3_1 hold785 (.A(\FpgaPins_Fpga_GAME_wait_counter_a2[13] ),
    .X(net1722));
 sg13g2_dlygate4sd3_1 hold786 (.A(_2604_),
    .X(net1723));
 sg13g2_dlygate4sd3_1 hold787 (.A(_0535_),
    .X(net1724));
 sg13g2_dlygate4sd3_1 hold788 (.A(\FpgaPins_Fpga_GAME_score_a4[0] ),
    .X(net1725));
 sg13g2_dlygate4sd3_1 hold789 (.A(_0094_),
    .X(net1726));
 sg13g2_dlygate4sd3_1 hold790 (.A(_1829_),
    .X(net1727));
 sg13g2_dlygate4sd3_1 hold791 (.A(FpgaPins_Fpga_GAME_right_btn_a2),
    .X(net1728));
 sg13g2_dlygate4sd3_1 hold792 (.A(_2461_),
    .X(net1729));
 sg13g2_dlygate4sd3_1 hold793 (.A(_0355_),
    .X(net1730));
 sg13g2_dlygate4sd3_1 hold794 (.A(FpgaPins_Fpga_LIPSI_is_2cyc_a2),
    .X(net1731));
 sg13g2_dlygate4sd3_1 hold795 (.A(\C1.next_state_var[6] ),
    .X(net1732));
 sg13g2_dlygate4sd3_1 hold796 (.A(\C1.next_state_var[5] ),
    .X(net1733));
 sg13g2_dlygate4sd3_1 hold797 (.A(\C1.counter2[2] ),
    .X(net1734));
 sg13g2_dlygate4sd3_1 hold798 (.A(_2540_),
    .X(net1735));
 sg13g2_dlygate4sd3_1 hold799 (.A(\C1.timer[0] ),
    .X(net1736));
 sg13g2_dlygate4sd3_1 hold800 (.A(_0136_),
    .X(net1737));
 sg13g2_dlygate4sd3_1 hold801 (.A(_0153_),
    .X(net1738));
 sg13g2_dlygate4sd3_1 hold802 (.A(_1447_),
    .X(net1739));
 sg13g2_dlygate4sd3_1 hold803 (.A(\C1.counter1[3] ),
    .X(net1740));
 sg13g2_dlygate4sd3_1 hold804 (.A(\C1.temp[0] ),
    .X(net1741));
 sg13g2_dlygate4sd3_1 hold805 (.A(\C1.temp[1] ),
    .X(net1742));
 sg13g2_dlygate4sd3_1 hold806 (.A(_0092_),
    .X(net1743));
 sg13g2_dlygate4sd3_1 hold807 (.A(\C1.level[1] ),
    .X(net1744));
 sg13g2_dlygate4sd3_1 hold808 (.A(\C1.counter1[4] ),
    .X(net1745));
 sg13g2_dlygate4sd3_1 hold809 (.A(_1917_),
    .X(net1746));
 sg13g2_dlygate4sd3_1 hold810 (.A(\C1.next_state_var[3] ),
    .X(net1747));
 sg13g2_dlygate4sd3_1 hold811 (.A(\C1.counter1[1] ),
    .X(net1748));
 sg13g2_dlygate4sd3_1 hold812 (.A(_1903_),
    .X(net1749));
 sg13g2_dlygate4sd3_1 hold813 (.A(\C1.level[0] ),
    .X(net1750));
 sg13g2_dlygate4sd3_1 hold814 (.A(\C1.counter1[9] ),
    .X(net1751));
 sg13g2_dlygate4sd3_1 hold815 (.A(_0029_),
    .X(net1752));
 sg13g2_dlygate4sd3_1 hold816 (.A(\FpgaPins_Fpga_FSM_imem_wr_addr_a1[2] ),
    .X(net1753));
 sg13g2_dlygate4sd3_1 hold817 (.A(\C1.counter2[7] ),
    .X(net1754));
 sg13g2_dlygate4sd3_1 hold818 (.A(FpgaPins_Fpga_GAME_reset_a2),
    .X(net1755));
 sg13g2_dlygate4sd3_1 hold819 (.A(\FpgaPins_Fpga_GAME_count_speed3_a2[12] ),
    .X(net1756));
 sg13g2_dlygate4sd3_1 hold820 (.A(FpgaPins_Fpga_LIPSI_is_2cyc_a2),
    .X(net1757));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_88 ();
 sg13g2_decap_8 FILLER_10_95 ();
 sg13g2_fill_2 FILLER_10_102 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_fill_1 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_135 ();
 sg13g2_decap_8 FILLER_10_142 ();
 sg13g2_decap_8 FILLER_10_149 ();
 sg13g2_decap_8 FILLER_10_156 ();
 sg13g2_decap_8 FILLER_10_163 ();
 sg13g2_decap_8 FILLER_10_170 ();
 sg13g2_decap_8 FILLER_10_177 ();
 sg13g2_decap_8 FILLER_10_184 ();
 sg13g2_decap_8 FILLER_10_191 ();
 sg13g2_decap_8 FILLER_10_198 ();
 sg13g2_decap_8 FILLER_10_205 ();
 sg13g2_decap_8 FILLER_10_212 ();
 sg13g2_decap_8 FILLER_10_219 ();
 sg13g2_decap_8 FILLER_10_226 ();
 sg13g2_decap_8 FILLER_10_233 ();
 sg13g2_decap_8 FILLER_10_240 ();
 sg13g2_decap_8 FILLER_10_247 ();
 sg13g2_decap_8 FILLER_10_254 ();
 sg13g2_decap_8 FILLER_10_261 ();
 sg13g2_decap_8 FILLER_10_268 ();
 sg13g2_decap_8 FILLER_10_275 ();
 sg13g2_decap_8 FILLER_10_282 ();
 sg13g2_decap_8 FILLER_10_289 ();
 sg13g2_decap_8 FILLER_10_296 ();
 sg13g2_decap_8 FILLER_10_303 ();
 sg13g2_decap_8 FILLER_10_310 ();
 sg13g2_decap_8 FILLER_10_317 ();
 sg13g2_decap_8 FILLER_10_324 ();
 sg13g2_decap_8 FILLER_10_331 ();
 sg13g2_decap_8 FILLER_10_338 ();
 sg13g2_decap_8 FILLER_10_345 ();
 sg13g2_decap_8 FILLER_10_352 ();
 sg13g2_decap_8 FILLER_10_359 ();
 sg13g2_decap_8 FILLER_10_366 ();
 sg13g2_decap_8 FILLER_10_373 ();
 sg13g2_decap_8 FILLER_10_380 ();
 sg13g2_decap_8 FILLER_10_387 ();
 sg13g2_decap_8 FILLER_10_394 ();
 sg13g2_decap_8 FILLER_10_401 ();
 sg13g2_decap_8 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_10_415 ();
 sg13g2_decap_8 FILLER_10_422 ();
 sg13g2_decap_8 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_10_436 ();
 sg13g2_decap_8 FILLER_10_443 ();
 sg13g2_decap_8 FILLER_10_450 ();
 sg13g2_decap_8 FILLER_10_457 ();
 sg13g2_decap_8 FILLER_10_464 ();
 sg13g2_decap_8 FILLER_10_471 ();
 sg13g2_decap_8 FILLER_10_478 ();
 sg13g2_decap_8 FILLER_10_485 ();
 sg13g2_decap_8 FILLER_10_492 ();
 sg13g2_decap_8 FILLER_10_499 ();
 sg13g2_decap_8 FILLER_10_506 ();
 sg13g2_decap_8 FILLER_10_513 ();
 sg13g2_decap_8 FILLER_10_520 ();
 sg13g2_decap_8 FILLER_10_527 ();
 sg13g2_decap_8 FILLER_10_534 ();
 sg13g2_decap_8 FILLER_10_541 ();
 sg13g2_decap_8 FILLER_10_548 ();
 sg13g2_decap_8 FILLER_10_555 ();
 sg13g2_decap_8 FILLER_10_562 ();
 sg13g2_decap_8 FILLER_10_569 ();
 sg13g2_decap_8 FILLER_10_576 ();
 sg13g2_decap_8 FILLER_10_583 ();
 sg13g2_decap_8 FILLER_10_590 ();
 sg13g2_decap_8 FILLER_10_597 ();
 sg13g2_decap_8 FILLER_10_604 ();
 sg13g2_decap_8 FILLER_10_611 ();
 sg13g2_decap_8 FILLER_10_618 ();
 sg13g2_decap_8 FILLER_10_625 ();
 sg13g2_decap_8 FILLER_10_632 ();
 sg13g2_decap_8 FILLER_10_639 ();
 sg13g2_decap_8 FILLER_10_646 ();
 sg13g2_decap_8 FILLER_10_653 ();
 sg13g2_decap_8 FILLER_10_660 ();
 sg13g2_decap_8 FILLER_10_667 ();
 sg13g2_decap_8 FILLER_10_674 ();
 sg13g2_decap_8 FILLER_10_681 ();
 sg13g2_decap_8 FILLER_10_688 ();
 sg13g2_decap_8 FILLER_10_695 ();
 sg13g2_decap_8 FILLER_10_702 ();
 sg13g2_decap_8 FILLER_10_709 ();
 sg13g2_decap_8 FILLER_10_716 ();
 sg13g2_decap_8 FILLER_10_723 ();
 sg13g2_decap_8 FILLER_10_730 ();
 sg13g2_decap_8 FILLER_10_737 ();
 sg13g2_decap_8 FILLER_10_744 ();
 sg13g2_decap_8 FILLER_10_751 ();
 sg13g2_decap_8 FILLER_10_758 ();
 sg13g2_decap_8 FILLER_10_765 ();
 sg13g2_decap_8 FILLER_10_772 ();
 sg13g2_decap_8 FILLER_10_779 ();
 sg13g2_decap_8 FILLER_10_786 ();
 sg13g2_decap_8 FILLER_10_793 ();
 sg13g2_decap_8 FILLER_10_800 ();
 sg13g2_decap_8 FILLER_10_807 ();
 sg13g2_decap_8 FILLER_10_814 ();
 sg13g2_decap_8 FILLER_10_821 ();
 sg13g2_decap_8 FILLER_10_828 ();
 sg13g2_decap_8 FILLER_10_835 ();
 sg13g2_decap_8 FILLER_10_842 ();
 sg13g2_decap_8 FILLER_10_849 ();
 sg13g2_decap_4 FILLER_10_856 ();
 sg13g2_fill_2 FILLER_10_860 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_fill_1 FILLER_11_49 ();
 sg13g2_decap_4 FILLER_11_54 ();
 sg13g2_fill_2 FILLER_11_58 ();
 sg13g2_fill_2 FILLER_11_64 ();
 sg13g2_fill_1 FILLER_11_74 ();
 sg13g2_fill_2 FILLER_11_84 ();
 sg13g2_fill_1 FILLER_11_98 ();
 sg13g2_fill_1 FILLER_11_109 ();
 sg13g2_fill_1 FILLER_11_124 ();
 sg13g2_decap_8 FILLER_11_142 ();
 sg13g2_decap_8 FILLER_11_149 ();
 sg13g2_decap_8 FILLER_11_156 ();
 sg13g2_decap_8 FILLER_11_163 ();
 sg13g2_decap_8 FILLER_11_170 ();
 sg13g2_decap_8 FILLER_11_177 ();
 sg13g2_decap_8 FILLER_11_184 ();
 sg13g2_decap_8 FILLER_11_191 ();
 sg13g2_decap_8 FILLER_11_198 ();
 sg13g2_decap_8 FILLER_11_205 ();
 sg13g2_decap_8 FILLER_11_212 ();
 sg13g2_decap_8 FILLER_11_219 ();
 sg13g2_decap_8 FILLER_11_226 ();
 sg13g2_decap_8 FILLER_11_233 ();
 sg13g2_decap_8 FILLER_11_240 ();
 sg13g2_decap_8 FILLER_11_247 ();
 sg13g2_decap_8 FILLER_11_254 ();
 sg13g2_decap_8 FILLER_11_261 ();
 sg13g2_decap_8 FILLER_11_268 ();
 sg13g2_decap_8 FILLER_11_275 ();
 sg13g2_decap_8 FILLER_11_282 ();
 sg13g2_decap_8 FILLER_11_289 ();
 sg13g2_decap_8 FILLER_11_296 ();
 sg13g2_decap_4 FILLER_11_303 ();
 sg13g2_fill_1 FILLER_11_307 ();
 sg13g2_decap_8 FILLER_11_321 ();
 sg13g2_decap_8 FILLER_11_328 ();
 sg13g2_decap_8 FILLER_11_335 ();
 sg13g2_decap_8 FILLER_11_342 ();
 sg13g2_decap_8 FILLER_11_349 ();
 sg13g2_decap_8 FILLER_11_356 ();
 sg13g2_decap_8 FILLER_11_363 ();
 sg13g2_decap_8 FILLER_11_370 ();
 sg13g2_decap_4 FILLER_11_377 ();
 sg13g2_fill_1 FILLER_11_381 ();
 sg13g2_fill_2 FILLER_11_392 ();
 sg13g2_fill_1 FILLER_11_407 ();
 sg13g2_fill_1 FILLER_11_418 ();
 sg13g2_fill_2 FILLER_11_423 ();
 sg13g2_decap_8 FILLER_11_435 ();
 sg13g2_fill_2 FILLER_11_442 ();
 sg13g2_fill_1 FILLER_11_444 ();
 sg13g2_decap_8 FILLER_11_454 ();
 sg13g2_decap_4 FILLER_11_461 ();
 sg13g2_fill_2 FILLER_11_465 ();
 sg13g2_fill_1 FILLER_11_502 ();
 sg13g2_fill_1 FILLER_11_507 ();
 sg13g2_fill_2 FILLER_11_518 ();
 sg13g2_fill_1 FILLER_11_520 ();
 sg13g2_decap_4 FILLER_11_531 ();
 sg13g2_decap_8 FILLER_11_544 ();
 sg13g2_fill_2 FILLER_11_551 ();
 sg13g2_decap_8 FILLER_11_563 ();
 sg13g2_decap_8 FILLER_11_570 ();
 sg13g2_decap_8 FILLER_11_577 ();
 sg13g2_decap_8 FILLER_11_584 ();
 sg13g2_decap_8 FILLER_11_591 ();
 sg13g2_decap_8 FILLER_11_598 ();
 sg13g2_decap_8 FILLER_11_605 ();
 sg13g2_decap_8 FILLER_11_612 ();
 sg13g2_decap_8 FILLER_11_619 ();
 sg13g2_decap_8 FILLER_11_626 ();
 sg13g2_decap_8 FILLER_11_633 ();
 sg13g2_decap_8 FILLER_11_640 ();
 sg13g2_decap_8 FILLER_11_647 ();
 sg13g2_decap_8 FILLER_11_654 ();
 sg13g2_decap_8 FILLER_11_661 ();
 sg13g2_decap_8 FILLER_11_668 ();
 sg13g2_decap_8 FILLER_11_675 ();
 sg13g2_decap_8 FILLER_11_682 ();
 sg13g2_decap_8 FILLER_11_689 ();
 sg13g2_decap_8 FILLER_11_696 ();
 sg13g2_decap_8 FILLER_11_703 ();
 sg13g2_decap_8 FILLER_11_710 ();
 sg13g2_decap_8 FILLER_11_717 ();
 sg13g2_decap_8 FILLER_11_724 ();
 sg13g2_decap_8 FILLER_11_731 ();
 sg13g2_decap_8 FILLER_11_738 ();
 sg13g2_decap_8 FILLER_11_745 ();
 sg13g2_decap_8 FILLER_11_752 ();
 sg13g2_decap_8 FILLER_11_759 ();
 sg13g2_decap_8 FILLER_11_766 ();
 sg13g2_decap_8 FILLER_11_773 ();
 sg13g2_decap_8 FILLER_11_780 ();
 sg13g2_decap_8 FILLER_11_787 ();
 sg13g2_decap_8 FILLER_11_794 ();
 sg13g2_decap_8 FILLER_11_801 ();
 sg13g2_decap_8 FILLER_11_808 ();
 sg13g2_decap_8 FILLER_11_815 ();
 sg13g2_decap_8 FILLER_11_822 ();
 sg13g2_decap_8 FILLER_11_829 ();
 sg13g2_decap_8 FILLER_11_836 ();
 sg13g2_decap_8 FILLER_11_843 ();
 sg13g2_decap_8 FILLER_11_850 ();
 sg13g2_decap_4 FILLER_11_857 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_4 FILLER_12_35 ();
 sg13g2_fill_2 FILLER_12_122 ();
 sg13g2_fill_1 FILLER_12_124 ();
 sg13g2_fill_2 FILLER_12_151 ();
 sg13g2_decap_8 FILLER_12_157 ();
 sg13g2_decap_8 FILLER_12_164 ();
 sg13g2_decap_8 FILLER_12_171 ();
 sg13g2_decap_8 FILLER_12_178 ();
 sg13g2_decap_8 FILLER_12_185 ();
 sg13g2_decap_8 FILLER_12_192 ();
 sg13g2_decap_8 FILLER_12_199 ();
 sg13g2_decap_8 FILLER_12_206 ();
 sg13g2_decap_8 FILLER_12_213 ();
 sg13g2_decap_8 FILLER_12_220 ();
 sg13g2_decap_8 FILLER_12_227 ();
 sg13g2_decap_8 FILLER_12_234 ();
 sg13g2_decap_8 FILLER_12_241 ();
 sg13g2_decap_8 FILLER_12_248 ();
 sg13g2_decap_8 FILLER_12_255 ();
 sg13g2_decap_8 FILLER_12_262 ();
 sg13g2_decap_8 FILLER_12_269 ();
 sg13g2_decap_8 FILLER_12_276 ();
 sg13g2_decap_8 FILLER_12_283 ();
 sg13g2_decap_4 FILLER_12_294 ();
 sg13g2_fill_2 FILLER_12_298 ();
 sg13g2_fill_2 FILLER_12_326 ();
 sg13g2_fill_1 FILLER_12_338 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_fill_1 FILLER_12_382 ();
 sg13g2_fill_2 FILLER_12_461 ();
 sg13g2_fill_1 FILLER_12_463 ();
 sg13g2_fill_2 FILLER_12_478 ();
 sg13g2_fill_2 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_596 ();
 sg13g2_fill_2 FILLER_12_603 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_fill_2 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_628 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_fill_2 FILLER_13_35 ();
 sg13g2_fill_2 FILLER_13_59 ();
 sg13g2_fill_1 FILLER_13_61 ();
 sg13g2_fill_1 FILLER_13_96 ();
 sg13g2_fill_2 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_4 FILLER_13_273 ();
 sg13g2_fill_2 FILLER_13_277 ();
 sg13g2_fill_2 FILLER_13_315 ();
 sg13g2_fill_1 FILLER_13_317 ();
 sg13g2_fill_2 FILLER_13_328 ();
 sg13g2_fill_2 FILLER_13_392 ();
 sg13g2_fill_1 FILLER_13_394 ();
 sg13g2_decap_8 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_13_415 ();
 sg13g2_fill_1 FILLER_13_441 ();
 sg13g2_fill_2 FILLER_13_468 ();
 sg13g2_fill_2 FILLER_13_513 ();
 sg13g2_decap_4 FILLER_13_524 ();
 sg13g2_fill_1 FILLER_13_528 ();
 sg13g2_decap_4 FILLER_13_533 ();
 sg13g2_fill_1 FILLER_13_537 ();
 sg13g2_fill_2 FILLER_13_564 ();
 sg13g2_fill_1 FILLER_13_593 ();
 sg13g2_fill_2 FILLER_13_620 ();
 sg13g2_decap_8 FILLER_13_661 ();
 sg13g2_decap_8 FILLER_13_668 ();
 sg13g2_decap_8 FILLER_13_675 ();
 sg13g2_decap_8 FILLER_13_682 ();
 sg13g2_decap_8 FILLER_13_689 ();
 sg13g2_decap_8 FILLER_13_696 ();
 sg13g2_decap_8 FILLER_13_703 ();
 sg13g2_decap_8 FILLER_13_710 ();
 sg13g2_decap_8 FILLER_13_717 ();
 sg13g2_decap_8 FILLER_13_724 ();
 sg13g2_decap_8 FILLER_13_731 ();
 sg13g2_decap_8 FILLER_13_738 ();
 sg13g2_decap_8 FILLER_13_745 ();
 sg13g2_decap_8 FILLER_13_752 ();
 sg13g2_decap_8 FILLER_13_759 ();
 sg13g2_decap_8 FILLER_13_766 ();
 sg13g2_decap_8 FILLER_13_773 ();
 sg13g2_decap_8 FILLER_13_780 ();
 sg13g2_decap_8 FILLER_13_787 ();
 sg13g2_decap_8 FILLER_13_794 ();
 sg13g2_decap_8 FILLER_13_801 ();
 sg13g2_decap_8 FILLER_13_808 ();
 sg13g2_decap_8 FILLER_13_815 ();
 sg13g2_decap_8 FILLER_13_822 ();
 sg13g2_decap_8 FILLER_13_829 ();
 sg13g2_decap_8 FILLER_13_836 ();
 sg13g2_decap_8 FILLER_13_843 ();
 sg13g2_decap_8 FILLER_13_850 ();
 sg13g2_decap_4 FILLER_13_857 ();
 sg13g2_fill_1 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_fill_2 FILLER_14_28 ();
 sg13g2_fill_2 FILLER_14_56 ();
 sg13g2_fill_1 FILLER_14_58 ();
 sg13g2_fill_2 FILLER_14_78 ();
 sg13g2_fill_2 FILLER_14_120 ();
 sg13g2_fill_1 FILLER_14_122 ();
 sg13g2_fill_1 FILLER_14_128 ();
 sg13g2_decap_8 FILLER_14_170 ();
 sg13g2_decap_8 FILLER_14_177 ();
 sg13g2_decap_8 FILLER_14_184 ();
 sg13g2_decap_8 FILLER_14_191 ();
 sg13g2_decap_8 FILLER_14_198 ();
 sg13g2_decap_8 FILLER_14_205 ();
 sg13g2_decap_8 FILLER_14_212 ();
 sg13g2_decap_8 FILLER_14_219 ();
 sg13g2_decap_8 FILLER_14_226 ();
 sg13g2_decap_8 FILLER_14_233 ();
 sg13g2_decap_8 FILLER_14_240 ();
 sg13g2_decap_8 FILLER_14_247 ();
 sg13g2_decap_8 FILLER_14_254 ();
 sg13g2_fill_2 FILLER_14_261 ();
 sg13g2_decap_4 FILLER_14_342 ();
 sg13g2_fill_2 FILLER_14_367 ();
 sg13g2_fill_1 FILLER_14_369 ();
 sg13g2_fill_1 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_433 ();
 sg13g2_fill_1 FILLER_14_440 ();
 sg13g2_fill_1 FILLER_14_445 ();
 sg13g2_fill_1 FILLER_14_450 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_4 FILLER_14_476 ();
 sg13g2_fill_1 FILLER_14_480 ();
 sg13g2_decap_4 FILLER_14_485 ();
 sg13g2_fill_1 FILLER_14_489 ();
 sg13g2_fill_1 FILLER_14_505 ();
 sg13g2_decap_8 FILLER_14_516 ();
 sg13g2_fill_1 FILLER_14_523 ();
 sg13g2_fill_2 FILLER_14_534 ();
 sg13g2_fill_2 FILLER_14_558 ();
 sg13g2_fill_1 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_621 ();
 sg13g2_decap_8 FILLER_14_668 ();
 sg13g2_decap_8 FILLER_14_675 ();
 sg13g2_decap_8 FILLER_14_682 ();
 sg13g2_decap_8 FILLER_14_689 ();
 sg13g2_decap_8 FILLER_14_696 ();
 sg13g2_decap_8 FILLER_14_703 ();
 sg13g2_decap_8 FILLER_14_710 ();
 sg13g2_decap_8 FILLER_14_717 ();
 sg13g2_decap_8 FILLER_14_724 ();
 sg13g2_decap_8 FILLER_14_731 ();
 sg13g2_decap_8 FILLER_14_738 ();
 sg13g2_decap_8 FILLER_14_745 ();
 sg13g2_decap_8 FILLER_14_752 ();
 sg13g2_decap_8 FILLER_14_759 ();
 sg13g2_decap_8 FILLER_14_766 ();
 sg13g2_decap_8 FILLER_14_773 ();
 sg13g2_decap_8 FILLER_14_780 ();
 sg13g2_decap_8 FILLER_14_787 ();
 sg13g2_decap_8 FILLER_14_794 ();
 sg13g2_decap_8 FILLER_14_801 ();
 sg13g2_decap_8 FILLER_14_808 ();
 sg13g2_decap_8 FILLER_14_815 ();
 sg13g2_decap_8 FILLER_14_822 ();
 sg13g2_decap_8 FILLER_14_829 ();
 sg13g2_decap_8 FILLER_14_836 ();
 sg13g2_decap_8 FILLER_14_843 ();
 sg13g2_decap_8 FILLER_14_850 ();
 sg13g2_decap_4 FILLER_14_857 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_fill_2 FILLER_15_35 ();
 sg13g2_fill_1 FILLER_15_37 ();
 sg13g2_fill_2 FILLER_15_64 ();
 sg13g2_fill_1 FILLER_15_99 ();
 sg13g2_decap_8 FILLER_15_172 ();
 sg13g2_decap_4 FILLER_15_179 ();
 sg13g2_fill_2 FILLER_15_187 ();
 sg13g2_fill_2 FILLER_15_192 ();
 sg13g2_fill_1 FILLER_15_194 ();
 sg13g2_decap_8 FILLER_15_207 ();
 sg13g2_decap_8 FILLER_15_214 ();
 sg13g2_decap_8 FILLER_15_221 ();
 sg13g2_decap_8 FILLER_15_228 ();
 sg13g2_decap_8 FILLER_15_235 ();
 sg13g2_decap_8 FILLER_15_242 ();
 sg13g2_decap_8 FILLER_15_249 ();
 sg13g2_decap_4 FILLER_15_256 ();
 sg13g2_fill_2 FILLER_15_260 ();
 sg13g2_fill_2 FILLER_15_272 ();
 sg13g2_fill_1 FILLER_15_274 ();
 sg13g2_decap_8 FILLER_15_311 ();
 sg13g2_fill_2 FILLER_15_318 ();
 sg13g2_fill_1 FILLER_15_320 ();
 sg13g2_decap_4 FILLER_15_383 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_481 ();
 sg13g2_decap_4 FILLER_15_514 ();
 sg13g2_decap_4 FILLER_15_544 ();
 sg13g2_fill_1 FILLER_15_563 ();
 sg13g2_fill_2 FILLER_15_583 ();
 sg13g2_decap_4 FILLER_15_621 ();
 sg13g2_fill_1 FILLER_15_625 ();
 sg13g2_decap_4 FILLER_15_669 ();
 sg13g2_decap_8 FILLER_15_682 ();
 sg13g2_decap_8 FILLER_15_689 ();
 sg13g2_decap_8 FILLER_15_696 ();
 sg13g2_decap_8 FILLER_15_703 ();
 sg13g2_decap_8 FILLER_15_710 ();
 sg13g2_decap_8 FILLER_15_717 ();
 sg13g2_decap_8 FILLER_15_724 ();
 sg13g2_decap_8 FILLER_15_731 ();
 sg13g2_decap_8 FILLER_15_738 ();
 sg13g2_decap_8 FILLER_15_745 ();
 sg13g2_decap_8 FILLER_15_752 ();
 sg13g2_decap_8 FILLER_15_759 ();
 sg13g2_decap_8 FILLER_15_766 ();
 sg13g2_decap_8 FILLER_15_773 ();
 sg13g2_decap_8 FILLER_15_780 ();
 sg13g2_decap_8 FILLER_15_787 ();
 sg13g2_decap_8 FILLER_15_794 ();
 sg13g2_decap_8 FILLER_15_801 ();
 sg13g2_decap_8 FILLER_15_808 ();
 sg13g2_decap_8 FILLER_15_815 ();
 sg13g2_decap_8 FILLER_15_822 ();
 sg13g2_decap_8 FILLER_15_829 ();
 sg13g2_decap_8 FILLER_15_836 ();
 sg13g2_decap_8 FILLER_15_843 ();
 sg13g2_decap_8 FILLER_15_850 ();
 sg13g2_decap_4 FILLER_15_857 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_fill_1 FILLER_16_35 ();
 sg13g2_fill_2 FILLER_16_160 ();
 sg13g2_fill_1 FILLER_16_162 ();
 sg13g2_fill_2 FILLER_16_168 ();
 sg13g2_fill_2 FILLER_16_178 ();
 sg13g2_fill_1 FILLER_16_180 ();
 sg13g2_fill_2 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_230 ();
 sg13g2_decap_8 FILLER_16_237 ();
 sg13g2_decap_8 FILLER_16_244 ();
 sg13g2_decap_8 FILLER_16_251 ();
 sg13g2_fill_2 FILLER_16_272 ();
 sg13g2_fill_1 FILLER_16_274 ();
 sg13g2_decap_4 FILLER_16_324 ();
 sg13g2_fill_2 FILLER_16_328 ();
 sg13g2_fill_2 FILLER_16_354 ();
 sg13g2_fill_1 FILLER_16_405 ();
 sg13g2_decap_4 FILLER_16_419 ();
 sg13g2_fill_2 FILLER_16_423 ();
 sg13g2_fill_2 FILLER_16_461 ();
 sg13g2_fill_1 FILLER_16_463 ();
 sg13g2_fill_2 FILLER_16_472 ();
 sg13g2_decap_4 FILLER_16_535 ();
 sg13g2_fill_1 FILLER_16_539 ();
 sg13g2_decap_4 FILLER_16_545 ();
 sg13g2_decap_8 FILLER_16_688 ();
 sg13g2_decap_8 FILLER_16_695 ();
 sg13g2_decap_8 FILLER_16_702 ();
 sg13g2_decap_8 FILLER_16_709 ();
 sg13g2_decap_8 FILLER_16_716 ();
 sg13g2_decap_8 FILLER_16_723 ();
 sg13g2_decap_8 FILLER_16_730 ();
 sg13g2_decap_8 FILLER_16_737 ();
 sg13g2_decap_8 FILLER_16_744 ();
 sg13g2_decap_8 FILLER_16_751 ();
 sg13g2_decap_8 FILLER_16_758 ();
 sg13g2_decap_8 FILLER_16_765 ();
 sg13g2_decap_8 FILLER_16_772 ();
 sg13g2_decap_8 FILLER_16_779 ();
 sg13g2_decap_8 FILLER_16_786 ();
 sg13g2_decap_8 FILLER_16_793 ();
 sg13g2_decap_8 FILLER_16_800 ();
 sg13g2_decap_8 FILLER_16_807 ();
 sg13g2_decap_8 FILLER_16_814 ();
 sg13g2_decap_8 FILLER_16_821 ();
 sg13g2_decap_8 FILLER_16_828 ();
 sg13g2_decap_8 FILLER_16_835 ();
 sg13g2_decap_8 FILLER_16_842 ();
 sg13g2_decap_8 FILLER_16_849 ();
 sg13g2_decap_4 FILLER_16_856 ();
 sg13g2_fill_2 FILLER_16_860 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_7 ();
 sg13g2_fill_2 FILLER_17_11 ();
 sg13g2_decap_4 FILLER_17_17 ();
 sg13g2_decap_8 FILLER_17_29 ();
 sg13g2_fill_1 FILLER_17_36 ();
 sg13g2_fill_2 FILLER_17_82 ();
 sg13g2_fill_1 FILLER_17_84 ();
 sg13g2_fill_2 FILLER_17_108 ();
 sg13g2_fill_2 FILLER_17_130 ();
 sg13g2_fill_2 FILLER_17_213 ();
 sg13g2_fill_2 FILLER_17_241 ();
 sg13g2_fill_1 FILLER_17_243 ();
 sg13g2_decap_8 FILLER_17_309 ();
 sg13g2_decap_4 FILLER_17_342 ();
 sg13g2_fill_2 FILLER_17_372 ();
 sg13g2_fill_1 FILLER_17_374 ();
 sg13g2_fill_2 FILLER_17_394 ();
 sg13g2_decap_4 FILLER_17_422 ();
 sg13g2_decap_4 FILLER_17_431 ();
 sg13g2_fill_1 FILLER_17_435 ();
 sg13g2_decap_4 FILLER_17_458 ();
 sg13g2_fill_1 FILLER_17_466 ();
 sg13g2_decap_8 FILLER_17_481 ();
 sg13g2_fill_1 FILLER_17_488 ();
 sg13g2_fill_2 FILLER_17_493 ();
 sg13g2_decap_8 FILLER_17_505 ();
 sg13g2_fill_2 FILLER_17_512 ();
 sg13g2_fill_1 FILLER_17_514 ();
 sg13g2_fill_1 FILLER_17_541 ();
 sg13g2_decap_4 FILLER_17_555 ();
 sg13g2_fill_1 FILLER_17_559 ();
 sg13g2_fill_2 FILLER_17_564 ();
 sg13g2_fill_1 FILLER_17_566 ();
 sg13g2_fill_2 FILLER_17_571 ();
 sg13g2_fill_2 FILLER_17_583 ();
 sg13g2_fill_1 FILLER_17_598 ();
 sg13g2_decap_4 FILLER_17_634 ();
 sg13g2_fill_2 FILLER_17_667 ();
 sg13g2_fill_1 FILLER_17_669 ();
 sg13g2_decap_8 FILLER_17_674 ();
 sg13g2_decap_8 FILLER_17_681 ();
 sg13g2_decap_8 FILLER_17_688 ();
 sg13g2_decap_8 FILLER_17_695 ();
 sg13g2_decap_8 FILLER_17_702 ();
 sg13g2_decap_8 FILLER_17_709 ();
 sg13g2_decap_8 FILLER_17_716 ();
 sg13g2_decap_8 FILLER_17_723 ();
 sg13g2_decap_8 FILLER_17_730 ();
 sg13g2_decap_8 FILLER_17_737 ();
 sg13g2_decap_8 FILLER_17_744 ();
 sg13g2_decap_8 FILLER_17_751 ();
 sg13g2_decap_8 FILLER_17_758 ();
 sg13g2_decap_8 FILLER_17_765 ();
 sg13g2_decap_8 FILLER_17_772 ();
 sg13g2_decap_8 FILLER_17_779 ();
 sg13g2_decap_8 FILLER_17_786 ();
 sg13g2_decap_8 FILLER_17_793 ();
 sg13g2_decap_8 FILLER_17_800 ();
 sg13g2_decap_8 FILLER_17_807 ();
 sg13g2_decap_8 FILLER_17_814 ();
 sg13g2_decap_8 FILLER_17_821 ();
 sg13g2_decap_8 FILLER_17_828 ();
 sg13g2_decap_8 FILLER_17_835 ();
 sg13g2_decap_8 FILLER_17_842 ();
 sg13g2_decap_8 FILLER_17_849 ();
 sg13g2_decap_4 FILLER_17_856 ();
 sg13g2_fill_2 FILLER_17_860 ();
 sg13g2_decap_4 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_30 ();
 sg13g2_fill_1 FILLER_18_78 ();
 sg13g2_fill_2 FILLER_18_134 ();
 sg13g2_fill_1 FILLER_18_136 ();
 sg13g2_fill_1 FILLER_18_163 ();
 sg13g2_fill_2 FILLER_18_183 ();
 sg13g2_fill_2 FILLER_18_200 ();
 sg13g2_decap_8 FILLER_18_246 ();
 sg13g2_decap_4 FILLER_18_253 ();
 sg13g2_fill_2 FILLER_18_257 ();
 sg13g2_fill_1 FILLER_18_263 ();
 sg13g2_fill_2 FILLER_18_277 ();
 sg13g2_fill_2 FILLER_18_284 ();
 sg13g2_fill_1 FILLER_18_286 ();
 sg13g2_fill_2 FILLER_18_349 ();
 sg13g2_fill_2 FILLER_18_426 ();
 sg13g2_fill_2 FILLER_18_438 ();
 sg13g2_fill_1 FILLER_18_440 ();
 sg13g2_decap_4 FILLER_18_445 ();
 sg13g2_fill_2 FILLER_18_449 ();
 sg13g2_fill_2 FILLER_18_477 ();
 sg13g2_fill_2 FILLER_18_510 ();
 sg13g2_decap_8 FILLER_18_538 ();
 sg13g2_fill_1 FILLER_18_545 ();
 sg13g2_decap_4 FILLER_18_555 ();
 sg13g2_fill_1 FILLER_18_559 ();
 sg13g2_decap_4 FILLER_18_570 ();
 sg13g2_fill_1 FILLER_18_574 ();
 sg13g2_decap_8 FILLER_18_649 ();
 sg13g2_fill_1 FILLER_18_656 ();
 sg13g2_decap_8 FILLER_18_683 ();
 sg13g2_decap_8 FILLER_18_690 ();
 sg13g2_decap_8 FILLER_18_697 ();
 sg13g2_decap_8 FILLER_18_704 ();
 sg13g2_decap_8 FILLER_18_711 ();
 sg13g2_decap_8 FILLER_18_718 ();
 sg13g2_decap_8 FILLER_18_725 ();
 sg13g2_decap_8 FILLER_18_732 ();
 sg13g2_decap_8 FILLER_18_739 ();
 sg13g2_decap_8 FILLER_18_746 ();
 sg13g2_decap_8 FILLER_18_753 ();
 sg13g2_decap_8 FILLER_18_760 ();
 sg13g2_decap_8 FILLER_18_767 ();
 sg13g2_decap_8 FILLER_18_774 ();
 sg13g2_decap_8 FILLER_18_781 ();
 sg13g2_decap_8 FILLER_18_788 ();
 sg13g2_decap_8 FILLER_18_795 ();
 sg13g2_decap_8 FILLER_18_802 ();
 sg13g2_decap_8 FILLER_18_809 ();
 sg13g2_decap_8 FILLER_18_816 ();
 sg13g2_decap_8 FILLER_18_823 ();
 sg13g2_decap_8 FILLER_18_830 ();
 sg13g2_decap_8 FILLER_18_837 ();
 sg13g2_decap_8 FILLER_18_844 ();
 sg13g2_decap_8 FILLER_18_851 ();
 sg13g2_decap_4 FILLER_18_858 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_24 ();
 sg13g2_fill_1 FILLER_19_61 ();
 sg13g2_fill_2 FILLER_19_148 ();
 sg13g2_fill_2 FILLER_19_185 ();
 sg13g2_fill_1 FILLER_19_187 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_fill_1 FILLER_19_266 ();
 sg13g2_fill_2 FILLER_19_271 ();
 sg13g2_fill_1 FILLER_19_283 ();
 sg13g2_decap_4 FILLER_19_294 ();
 sg13g2_fill_2 FILLER_19_307 ();
 sg13g2_fill_2 FILLER_19_319 ();
 sg13g2_fill_1 FILLER_19_321 ();
 sg13g2_decap_4 FILLER_19_356 ();
 sg13g2_fill_1 FILLER_19_360 ();
 sg13g2_fill_1 FILLER_19_371 ();
 sg13g2_fill_2 FILLER_19_386 ();
 sg13g2_fill_1 FILLER_19_388 ();
 sg13g2_fill_2 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_405 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_fill_2 FILLER_19_465 ();
 sg13g2_fill_2 FILLER_19_472 ();
 sg13g2_fill_2 FILLER_19_491 ();
 sg13g2_fill_2 FILLER_19_520 ();
 sg13g2_fill_1 FILLER_19_522 ();
 sg13g2_fill_2 FILLER_19_536 ();
 sg13g2_decap_4 FILLER_19_543 ();
 sg13g2_fill_2 FILLER_19_595 ();
 sg13g2_decap_4 FILLER_19_605 ();
 sg13g2_fill_2 FILLER_19_609 ();
 sg13g2_decap_4 FILLER_19_621 ();
 sg13g2_fill_1 FILLER_19_633 ();
 sg13g2_fill_2 FILLER_19_638 ();
 sg13g2_decap_8 FILLER_19_650 ();
 sg13g2_decap_8 FILLER_19_689 ();
 sg13g2_decap_8 FILLER_19_696 ();
 sg13g2_decap_8 FILLER_19_703 ();
 sg13g2_decap_8 FILLER_19_710 ();
 sg13g2_decap_8 FILLER_19_717 ();
 sg13g2_decap_8 FILLER_19_724 ();
 sg13g2_decap_8 FILLER_19_731 ();
 sg13g2_decap_8 FILLER_19_738 ();
 sg13g2_decap_8 FILLER_19_745 ();
 sg13g2_decap_8 FILLER_19_752 ();
 sg13g2_decap_8 FILLER_19_759 ();
 sg13g2_decap_8 FILLER_19_766 ();
 sg13g2_decap_8 FILLER_19_773 ();
 sg13g2_decap_8 FILLER_19_780 ();
 sg13g2_decap_8 FILLER_19_787 ();
 sg13g2_decap_8 FILLER_19_794 ();
 sg13g2_decap_8 FILLER_19_801 ();
 sg13g2_decap_8 FILLER_19_808 ();
 sg13g2_decap_8 FILLER_19_815 ();
 sg13g2_decap_8 FILLER_19_822 ();
 sg13g2_decap_8 FILLER_19_829 ();
 sg13g2_decap_8 FILLER_19_836 ();
 sg13g2_decap_8 FILLER_19_843 ();
 sg13g2_decap_8 FILLER_19_850 ();
 sg13g2_decap_4 FILLER_19_857 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_30 ();
 sg13g2_fill_1 FILLER_20_50 ();
 sg13g2_fill_1 FILLER_20_67 ();
 sg13g2_fill_1 FILLER_20_94 ();
 sg13g2_fill_1 FILLER_20_152 ();
 sg13g2_fill_2 FILLER_20_172 ();
 sg13g2_fill_1 FILLER_20_174 ();
 sg13g2_fill_2 FILLER_20_184 ();
 sg13g2_fill_2 FILLER_20_217 ();
 sg13g2_fill_1 FILLER_20_219 ();
 sg13g2_decap_8 FILLER_20_246 ();
 sg13g2_fill_2 FILLER_20_253 ();
 sg13g2_fill_1 FILLER_20_255 ();
 sg13g2_fill_2 FILLER_20_360 ();
 sg13g2_decap_8 FILLER_20_388 ();
 sg13g2_decap_4 FILLER_20_439 ();
 sg13g2_fill_1 FILLER_20_443 ();
 sg13g2_fill_1 FILLER_20_465 ();
 sg13g2_fill_1 FILLER_20_475 ();
 sg13g2_fill_1 FILLER_20_490 ();
 sg13g2_decap_4 FILLER_20_495 ();
 sg13g2_fill_2 FILLER_20_504 ();
 sg13g2_fill_1 FILLER_20_506 ();
 sg13g2_fill_2 FILLER_20_556 ();
 sg13g2_fill_2 FILLER_20_576 ();
 sg13g2_decap_4 FILLER_20_643 ();
 sg13g2_fill_2 FILLER_20_647 ();
 sg13g2_fill_2 FILLER_20_680 ();
 sg13g2_decap_8 FILLER_20_695 ();
 sg13g2_decap_8 FILLER_20_702 ();
 sg13g2_decap_8 FILLER_20_709 ();
 sg13g2_decap_8 FILLER_20_716 ();
 sg13g2_decap_8 FILLER_20_723 ();
 sg13g2_decap_8 FILLER_20_730 ();
 sg13g2_decap_8 FILLER_20_737 ();
 sg13g2_decap_8 FILLER_20_744 ();
 sg13g2_decap_8 FILLER_20_751 ();
 sg13g2_decap_8 FILLER_20_758 ();
 sg13g2_decap_8 FILLER_20_765 ();
 sg13g2_decap_8 FILLER_20_772 ();
 sg13g2_decap_8 FILLER_20_779 ();
 sg13g2_decap_8 FILLER_20_786 ();
 sg13g2_decap_8 FILLER_20_793 ();
 sg13g2_decap_8 FILLER_20_800 ();
 sg13g2_decap_8 FILLER_20_807 ();
 sg13g2_decap_8 FILLER_20_814 ();
 sg13g2_decap_8 FILLER_20_821 ();
 sg13g2_decap_8 FILLER_20_828 ();
 sg13g2_decap_8 FILLER_20_835 ();
 sg13g2_decap_8 FILLER_20_842 ();
 sg13g2_decap_8 FILLER_20_849 ();
 sg13g2_decap_4 FILLER_20_856 ();
 sg13g2_fill_2 FILLER_20_860 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_2 ();
 sg13g2_fill_2 FILLER_21_29 ();
 sg13g2_fill_1 FILLER_21_31 ();
 sg13g2_fill_2 FILLER_21_84 ();
 sg13g2_fill_2 FILLER_21_96 ();
 sg13g2_fill_2 FILLER_21_133 ();
 sg13g2_fill_1 FILLER_21_176 ();
 sg13g2_fill_1 FILLER_21_230 ();
 sg13g2_fill_2 FILLER_21_330 ();
 sg13g2_fill_1 FILLER_21_332 ();
 sg13g2_decap_8 FILLER_21_361 ();
 sg13g2_fill_2 FILLER_21_368 ();
 sg13g2_fill_1 FILLER_21_370 ();
 sg13g2_fill_2 FILLER_21_385 ();
 sg13g2_fill_1 FILLER_21_400 ();
 sg13g2_decap_4 FILLER_21_458 ();
 sg13g2_fill_2 FILLER_21_462 ();
 sg13g2_decap_4 FILLER_21_470 ();
 sg13g2_fill_2 FILLER_21_524 ();
 sg13g2_decap_4 FILLER_21_543 ();
 sg13g2_fill_1 FILLER_21_547 ();
 sg13g2_decap_4 FILLER_21_584 ();
 sg13g2_fill_2 FILLER_21_588 ();
 sg13g2_decap_4 FILLER_21_612 ();
 sg13g2_fill_1 FILLER_21_616 ();
 sg13g2_fill_1 FILLER_21_626 ();
 sg13g2_decap_8 FILLER_21_631 ();
 sg13g2_fill_1 FILLER_21_638 ();
 sg13g2_decap_8 FILLER_21_649 ();
 sg13g2_fill_2 FILLER_21_656 ();
 sg13g2_decap_8 FILLER_21_698 ();
 sg13g2_decap_8 FILLER_21_705 ();
 sg13g2_decap_8 FILLER_21_712 ();
 sg13g2_decap_8 FILLER_21_719 ();
 sg13g2_decap_8 FILLER_21_726 ();
 sg13g2_decap_8 FILLER_21_733 ();
 sg13g2_decap_8 FILLER_21_740 ();
 sg13g2_decap_8 FILLER_21_747 ();
 sg13g2_decap_8 FILLER_21_754 ();
 sg13g2_decap_8 FILLER_21_761 ();
 sg13g2_decap_8 FILLER_21_768 ();
 sg13g2_decap_8 FILLER_21_775 ();
 sg13g2_decap_8 FILLER_21_782 ();
 sg13g2_decap_8 FILLER_21_789 ();
 sg13g2_decap_8 FILLER_21_796 ();
 sg13g2_decap_8 FILLER_21_803 ();
 sg13g2_decap_8 FILLER_21_810 ();
 sg13g2_decap_8 FILLER_21_817 ();
 sg13g2_decap_8 FILLER_21_824 ();
 sg13g2_decap_8 FILLER_21_831 ();
 sg13g2_decap_8 FILLER_21_838 ();
 sg13g2_decap_8 FILLER_21_845 ();
 sg13g2_decap_8 FILLER_21_852 ();
 sg13g2_fill_2 FILLER_21_859 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_7 ();
 sg13g2_fill_2 FILLER_22_26 ();
 sg13g2_fill_1 FILLER_22_28 ();
 sg13g2_fill_2 FILLER_22_59 ();
 sg13g2_fill_1 FILLER_22_61 ();
 sg13g2_fill_2 FILLER_22_115 ();
 sg13g2_fill_1 FILLER_22_206 ();
 sg13g2_fill_1 FILLER_22_243 ();
 sg13g2_fill_1 FILLER_22_253 ();
 sg13g2_fill_2 FILLER_22_268 ();
 sg13g2_decap_4 FILLER_22_300 ();
 sg13g2_fill_2 FILLER_22_304 ();
 sg13g2_decap_4 FILLER_22_332 ();
 sg13g2_decap_4 FILLER_22_371 ();
 sg13g2_fill_1 FILLER_22_375 ();
 sg13g2_decap_4 FILLER_22_423 ();
 sg13g2_fill_1 FILLER_22_427 ();
 sg13g2_decap_4 FILLER_22_436 ();
 sg13g2_fill_2 FILLER_22_440 ();
 sg13g2_decap_4 FILLER_22_455 ();
 sg13g2_fill_2 FILLER_22_459 ();
 sg13g2_fill_2 FILLER_22_466 ();
 sg13g2_decap_8 FILLER_22_486 ();
 sg13g2_decap_4 FILLER_22_493 ();
 sg13g2_decap_8 FILLER_22_542 ();
 sg13g2_decap_8 FILLER_22_549 ();
 sg13g2_decap_4 FILLER_22_556 ();
 sg13g2_fill_1 FILLER_22_560 ();
 sg13g2_fill_2 FILLER_22_569 ();
 sg13g2_fill_1 FILLER_22_571 ();
 sg13g2_fill_1 FILLER_22_576 ();
 sg13g2_fill_2 FILLER_22_582 ();
 sg13g2_fill_2 FILLER_22_589 ();
 sg13g2_fill_2 FILLER_22_594 ();
 sg13g2_fill_1 FILLER_22_596 ();
 sg13g2_fill_2 FILLER_22_606 ();
 sg13g2_fill_1 FILLER_22_608 ();
 sg13g2_decap_8 FILLER_22_619 ();
 sg13g2_fill_2 FILLER_22_626 ();
 sg13g2_decap_4 FILLER_22_642 ();
 sg13g2_fill_1 FILLER_22_646 ();
 sg13g2_fill_2 FILLER_22_680 ();
 sg13g2_fill_1 FILLER_22_682 ();
 sg13g2_decap_8 FILLER_22_709 ();
 sg13g2_decap_8 FILLER_22_716 ();
 sg13g2_decap_8 FILLER_22_723 ();
 sg13g2_decap_8 FILLER_22_730 ();
 sg13g2_decap_8 FILLER_22_737 ();
 sg13g2_decap_8 FILLER_22_744 ();
 sg13g2_decap_8 FILLER_22_751 ();
 sg13g2_decap_8 FILLER_22_758 ();
 sg13g2_decap_8 FILLER_22_765 ();
 sg13g2_decap_8 FILLER_22_772 ();
 sg13g2_decap_8 FILLER_22_779 ();
 sg13g2_decap_8 FILLER_22_786 ();
 sg13g2_decap_8 FILLER_22_793 ();
 sg13g2_decap_8 FILLER_22_800 ();
 sg13g2_decap_8 FILLER_22_807 ();
 sg13g2_decap_8 FILLER_22_814 ();
 sg13g2_decap_8 FILLER_22_821 ();
 sg13g2_decap_8 FILLER_22_828 ();
 sg13g2_decap_8 FILLER_22_835 ();
 sg13g2_decap_8 FILLER_22_842 ();
 sg13g2_decap_8 FILLER_22_849 ();
 sg13g2_decap_4 FILLER_22_856 ();
 sg13g2_fill_2 FILLER_22_860 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_fill_2 FILLER_23_14 ();
 sg13g2_fill_2 FILLER_23_126 ();
 sg13g2_fill_2 FILLER_23_153 ();
 sg13g2_fill_1 FILLER_23_294 ();
 sg13g2_decap_4 FILLER_23_320 ();
 sg13g2_fill_1 FILLER_23_324 ();
 sg13g2_fill_2 FILLER_23_365 ();
 sg13g2_fill_1 FILLER_23_367 ();
 sg13g2_fill_2 FILLER_23_394 ();
 sg13g2_fill_1 FILLER_23_410 ();
 sg13g2_decap_4 FILLER_23_417 ();
 sg13g2_decap_4 FILLER_23_457 ();
 sg13g2_fill_2 FILLER_23_467 ();
 sg13g2_fill_2 FILLER_23_494 ();
 sg13g2_fill_1 FILLER_23_525 ();
 sg13g2_decap_8 FILLER_23_705 ();
 sg13g2_decap_8 FILLER_23_712 ();
 sg13g2_decap_8 FILLER_23_719 ();
 sg13g2_decap_8 FILLER_23_726 ();
 sg13g2_decap_8 FILLER_23_733 ();
 sg13g2_decap_8 FILLER_23_740 ();
 sg13g2_decap_8 FILLER_23_747 ();
 sg13g2_decap_8 FILLER_23_754 ();
 sg13g2_decap_8 FILLER_23_761 ();
 sg13g2_decap_8 FILLER_23_768 ();
 sg13g2_decap_8 FILLER_23_775 ();
 sg13g2_decap_8 FILLER_23_782 ();
 sg13g2_decap_8 FILLER_23_789 ();
 sg13g2_decap_8 FILLER_23_796 ();
 sg13g2_decap_8 FILLER_23_803 ();
 sg13g2_decap_8 FILLER_23_810 ();
 sg13g2_decap_8 FILLER_23_817 ();
 sg13g2_decap_8 FILLER_23_824 ();
 sg13g2_decap_8 FILLER_23_831 ();
 sg13g2_decap_8 FILLER_23_838 ();
 sg13g2_decap_8 FILLER_23_845 ();
 sg13g2_decap_8 FILLER_23_852 ();
 sg13g2_fill_2 FILLER_23_859 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_58 ();
 sg13g2_fill_1 FILLER_24_60 ();
 sg13g2_fill_1 FILLER_24_161 ();
 sg13g2_fill_2 FILLER_24_185 ();
 sg13g2_fill_2 FILLER_24_205 ();
 sg13g2_fill_1 FILLER_24_207 ();
 sg13g2_fill_2 FILLER_24_222 ();
 sg13g2_decap_4 FILLER_24_237 ();
 sg13g2_fill_1 FILLER_24_245 ();
 sg13g2_fill_2 FILLER_24_283 ();
 sg13g2_fill_2 FILLER_24_341 ();
 sg13g2_fill_1 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_365 ();
 sg13g2_decap_4 FILLER_24_372 ();
 sg13g2_fill_2 FILLER_24_429 ();
 sg13g2_fill_2 FILLER_24_439 ();
 sg13g2_fill_2 FILLER_24_460 ();
 sg13g2_decap_8 FILLER_24_468 ();
 sg13g2_fill_2 FILLER_24_475 ();
 sg13g2_fill_1 FILLER_24_477 ();
 sg13g2_fill_2 FILLER_24_488 ();
 sg13g2_fill_1 FILLER_24_506 ();
 sg13g2_fill_1 FILLER_24_551 ();
 sg13g2_fill_2 FILLER_24_584 ();
 sg13g2_fill_2 FILLER_24_613 ();
 sg13g2_fill_1 FILLER_24_615 ();
 sg13g2_fill_2 FILLER_24_643 ();
 sg13g2_fill_1 FILLER_24_645 ();
 sg13g2_decap_4 FILLER_24_655 ();
 sg13g2_fill_2 FILLER_24_659 ();
 sg13g2_fill_1 FILLER_24_693 ();
 sg13g2_decap_8 FILLER_24_698 ();
 sg13g2_decap_8 FILLER_24_705 ();
 sg13g2_decap_8 FILLER_24_712 ();
 sg13g2_decap_8 FILLER_24_719 ();
 sg13g2_decap_8 FILLER_24_726 ();
 sg13g2_decap_8 FILLER_24_733 ();
 sg13g2_decap_8 FILLER_24_740 ();
 sg13g2_decap_8 FILLER_24_747 ();
 sg13g2_decap_8 FILLER_24_754 ();
 sg13g2_decap_8 FILLER_24_761 ();
 sg13g2_decap_8 FILLER_24_768 ();
 sg13g2_decap_8 FILLER_24_775 ();
 sg13g2_decap_8 FILLER_24_782 ();
 sg13g2_decap_8 FILLER_24_789 ();
 sg13g2_decap_8 FILLER_24_796 ();
 sg13g2_decap_8 FILLER_24_803 ();
 sg13g2_decap_8 FILLER_24_810 ();
 sg13g2_decap_8 FILLER_24_817 ();
 sg13g2_decap_8 FILLER_24_824 ();
 sg13g2_decap_8 FILLER_24_831 ();
 sg13g2_decap_8 FILLER_24_838 ();
 sg13g2_decap_8 FILLER_24_845 ();
 sg13g2_decap_8 FILLER_24_852 ();
 sg13g2_fill_2 FILLER_24_859 ();
 sg13g2_fill_1 FILLER_24_861 ();
 sg13g2_fill_2 FILLER_25_35 ();
 sg13g2_fill_1 FILLER_25_37 ();
 sg13g2_fill_2 FILLER_25_47 ();
 sg13g2_fill_1 FILLER_25_49 ();
 sg13g2_fill_2 FILLER_25_73 ();
 sg13g2_fill_1 FILLER_25_94 ();
 sg13g2_fill_1 FILLER_25_101 ();
 sg13g2_fill_1 FILLER_25_137 ();
 sg13g2_fill_2 FILLER_25_164 ();
 sg13g2_fill_2 FILLER_25_183 ();
 sg13g2_fill_1 FILLER_25_191 ();
 sg13g2_decap_8 FILLER_25_232 ();
 sg13g2_fill_1 FILLER_25_239 ();
 sg13g2_decap_4 FILLER_25_266 ();
 sg13g2_fill_1 FILLER_25_300 ();
 sg13g2_decap_4 FILLER_25_327 ();
 sg13g2_fill_1 FILLER_25_357 ();
 sg13g2_decap_4 FILLER_25_363 ();
 sg13g2_fill_1 FILLER_25_367 ();
 sg13g2_fill_2 FILLER_25_395 ();
 sg13g2_fill_2 FILLER_25_421 ();
 sg13g2_fill_1 FILLER_25_428 ();
 sg13g2_fill_2 FILLER_25_433 ();
 sg13g2_decap_4 FILLER_25_444 ();
 sg13g2_fill_2 FILLER_25_466 ();
 sg13g2_fill_1 FILLER_25_468 ();
 sg13g2_fill_1 FILLER_25_473 ();
 sg13g2_decap_8 FILLER_25_489 ();
 sg13g2_fill_2 FILLER_25_496 ();
 sg13g2_fill_2 FILLER_25_528 ();
 sg13g2_fill_1 FILLER_25_548 ();
 sg13g2_fill_2 FILLER_25_598 ();
 sg13g2_fill_1 FILLER_25_634 ();
 sg13g2_fill_2 FILLER_25_681 ();
 sg13g2_fill_1 FILLER_25_683 ();
 sg13g2_fill_2 FILLER_25_688 ();
 sg13g2_decap_8 FILLER_25_716 ();
 sg13g2_decap_8 FILLER_25_723 ();
 sg13g2_decap_8 FILLER_25_730 ();
 sg13g2_decap_8 FILLER_25_737 ();
 sg13g2_decap_8 FILLER_25_744 ();
 sg13g2_decap_8 FILLER_25_751 ();
 sg13g2_decap_8 FILLER_25_758 ();
 sg13g2_decap_8 FILLER_25_765 ();
 sg13g2_decap_8 FILLER_25_772 ();
 sg13g2_decap_8 FILLER_25_779 ();
 sg13g2_decap_8 FILLER_25_786 ();
 sg13g2_decap_8 FILLER_25_793 ();
 sg13g2_decap_8 FILLER_25_800 ();
 sg13g2_decap_8 FILLER_25_807 ();
 sg13g2_decap_8 FILLER_25_814 ();
 sg13g2_decap_8 FILLER_25_821 ();
 sg13g2_decap_8 FILLER_25_828 ();
 sg13g2_decap_8 FILLER_25_835 ();
 sg13g2_decap_8 FILLER_25_842 ();
 sg13g2_decap_8 FILLER_25_849 ();
 sg13g2_decap_4 FILLER_25_856 ();
 sg13g2_fill_2 FILLER_25_860 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_110 ();
 sg13g2_fill_1 FILLER_26_121 ();
 sg13g2_fill_1 FILLER_26_141 ();
 sg13g2_fill_2 FILLER_26_218 ();
 sg13g2_decap_8 FILLER_26_228 ();
 sg13g2_decap_8 FILLER_26_235 ();
 sg13g2_decap_4 FILLER_26_242 ();
 sg13g2_fill_2 FILLER_26_246 ();
 sg13g2_fill_1 FILLER_26_256 ();
 sg13g2_fill_2 FILLER_26_276 ();
 sg13g2_decap_8 FILLER_26_309 ();
 sg13g2_decap_4 FILLER_26_316 ();
 sg13g2_fill_1 FILLER_26_320 ();
 sg13g2_fill_1 FILLER_26_343 ();
 sg13g2_decap_4 FILLER_26_357 ();
 sg13g2_fill_1 FILLER_26_361 ();
 sg13g2_fill_1 FILLER_26_388 ();
 sg13g2_fill_2 FILLER_26_456 ();
 sg13g2_fill_2 FILLER_26_499 ();
 sg13g2_decap_4 FILLER_26_621 ();
 sg13g2_fill_2 FILLER_26_625 ();
 sg13g2_decap_4 FILLER_26_641 ();
 sg13g2_fill_1 FILLER_26_645 ();
 sg13g2_decap_8 FILLER_26_650 ();
 sg13g2_decap_4 FILLER_26_657 ();
 sg13g2_fill_2 FILLER_26_661 ();
 sg13g2_fill_1 FILLER_26_673 ();
 sg13g2_decap_8 FILLER_26_713 ();
 sg13g2_decap_8 FILLER_26_720 ();
 sg13g2_decap_8 FILLER_26_727 ();
 sg13g2_decap_8 FILLER_26_734 ();
 sg13g2_decap_8 FILLER_26_741 ();
 sg13g2_decap_8 FILLER_26_748 ();
 sg13g2_decap_8 FILLER_26_755 ();
 sg13g2_decap_8 FILLER_26_762 ();
 sg13g2_decap_8 FILLER_26_769 ();
 sg13g2_decap_8 FILLER_26_776 ();
 sg13g2_decap_8 FILLER_26_783 ();
 sg13g2_decap_8 FILLER_26_790 ();
 sg13g2_decap_8 FILLER_26_797 ();
 sg13g2_decap_8 FILLER_26_804 ();
 sg13g2_decap_8 FILLER_26_811 ();
 sg13g2_decap_8 FILLER_26_818 ();
 sg13g2_decap_8 FILLER_26_825 ();
 sg13g2_decap_8 FILLER_26_832 ();
 sg13g2_decap_8 FILLER_26_839 ();
 sg13g2_decap_8 FILLER_26_846 ();
 sg13g2_decap_8 FILLER_26_853 ();
 sg13g2_fill_2 FILLER_26_860 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_17 ();
 sg13g2_fill_1 FILLER_27_36 ();
 sg13g2_fill_1 FILLER_27_134 ();
 sg13g2_fill_2 FILLER_27_235 ();
 sg13g2_decap_4 FILLER_27_263 ();
 sg13g2_fill_2 FILLER_27_302 ();
 sg13g2_fill_1 FILLER_27_304 ();
 sg13g2_fill_2 FILLER_27_331 ();
 sg13g2_decap_8 FILLER_27_361 ();
 sg13g2_decap_4 FILLER_27_368 ();
 sg13g2_fill_1 FILLER_27_372 ();
 sg13g2_fill_2 FILLER_27_387 ();
 sg13g2_fill_1 FILLER_27_389 ();
 sg13g2_fill_1 FILLER_27_395 ();
 sg13g2_fill_1 FILLER_27_410 ();
 sg13g2_decap_4 FILLER_27_425 ();
 sg13g2_decap_8 FILLER_27_444 ();
 sg13g2_decap_8 FILLER_27_461 ();
 sg13g2_decap_4 FILLER_27_468 ();
 sg13g2_fill_1 FILLER_27_472 ();
 sg13g2_fill_1 FILLER_27_554 ();
 sg13g2_fill_2 FILLER_27_588 ();
 sg13g2_fill_1 FILLER_27_590 ();
 sg13g2_fill_2 FILLER_27_613 ();
 sg13g2_fill_1 FILLER_27_615 ();
 sg13g2_fill_1 FILLER_27_652 ();
 sg13g2_decap_4 FILLER_27_657 ();
 sg13g2_fill_2 FILLER_27_680 ();
 sg13g2_decap_8 FILLER_27_708 ();
 sg13g2_decap_8 FILLER_27_715 ();
 sg13g2_decap_8 FILLER_27_722 ();
 sg13g2_decap_8 FILLER_27_729 ();
 sg13g2_decap_8 FILLER_27_736 ();
 sg13g2_decap_8 FILLER_27_743 ();
 sg13g2_decap_8 FILLER_27_750 ();
 sg13g2_decap_8 FILLER_27_757 ();
 sg13g2_decap_8 FILLER_27_764 ();
 sg13g2_decap_8 FILLER_27_771 ();
 sg13g2_decap_8 FILLER_27_778 ();
 sg13g2_decap_8 FILLER_27_785 ();
 sg13g2_decap_8 FILLER_27_792 ();
 sg13g2_decap_8 FILLER_27_799 ();
 sg13g2_decap_8 FILLER_27_806 ();
 sg13g2_decap_8 FILLER_27_813 ();
 sg13g2_decap_8 FILLER_27_820 ();
 sg13g2_decap_8 FILLER_27_827 ();
 sg13g2_decap_8 FILLER_27_834 ();
 sg13g2_decap_8 FILLER_27_841 ();
 sg13g2_decap_8 FILLER_27_848 ();
 sg13g2_decap_8 FILLER_27_855 ();
 sg13g2_fill_2 FILLER_28_38 ();
 sg13g2_fill_1 FILLER_28_40 ();
 sg13g2_fill_2 FILLER_28_79 ();
 sg13g2_fill_1 FILLER_28_81 ();
 sg13g2_fill_2 FILLER_28_101 ();
 sg13g2_fill_2 FILLER_28_108 ();
 sg13g2_fill_2 FILLER_28_141 ();
 sg13g2_fill_1 FILLER_28_195 ();
 sg13g2_decap_4 FILLER_28_230 ();
 sg13g2_fill_2 FILLER_28_234 ();
 sg13g2_fill_2 FILLER_28_309 ();
 sg13g2_decap_4 FILLER_28_330 ();
 sg13g2_fill_1 FILLER_28_334 ();
 sg13g2_decap_8 FILLER_28_387 ();
 sg13g2_decap_8 FILLER_28_394 ();
 sg13g2_fill_1 FILLER_28_401 ();
 sg13g2_decap_8 FILLER_28_428 ();
 sg13g2_decap_4 FILLER_28_435 ();
 sg13g2_fill_2 FILLER_28_439 ();
 sg13g2_fill_2 FILLER_28_451 ();
 sg13g2_fill_1 FILLER_28_453 ();
 sg13g2_fill_1 FILLER_28_570 ();
 sg13g2_decap_4 FILLER_28_612 ();
 sg13g2_fill_1 FILLER_28_616 ();
 sg13g2_decap_8 FILLER_28_709 ();
 sg13g2_decap_8 FILLER_28_716 ();
 sg13g2_decap_8 FILLER_28_723 ();
 sg13g2_decap_8 FILLER_28_730 ();
 sg13g2_decap_8 FILLER_28_737 ();
 sg13g2_decap_8 FILLER_28_744 ();
 sg13g2_decap_8 FILLER_28_751 ();
 sg13g2_decap_8 FILLER_28_758 ();
 sg13g2_decap_8 FILLER_28_765 ();
 sg13g2_decap_8 FILLER_28_772 ();
 sg13g2_decap_8 FILLER_28_779 ();
 sg13g2_decap_8 FILLER_28_786 ();
 sg13g2_decap_8 FILLER_28_793 ();
 sg13g2_decap_8 FILLER_28_800 ();
 sg13g2_decap_8 FILLER_28_807 ();
 sg13g2_decap_8 FILLER_28_814 ();
 sg13g2_decap_8 FILLER_28_821 ();
 sg13g2_decap_8 FILLER_28_828 ();
 sg13g2_decap_8 FILLER_28_835 ();
 sg13g2_decap_8 FILLER_28_842 ();
 sg13g2_decap_8 FILLER_28_849 ();
 sg13g2_decap_4 FILLER_28_856 ();
 sg13g2_fill_2 FILLER_28_860 ();
 sg13g2_fill_2 FILLER_29_31 ();
 sg13g2_fill_1 FILLER_29_33 ();
 sg13g2_fill_1 FILLER_29_128 ();
 sg13g2_fill_2 FILLER_29_155 ();
 sg13g2_decap_8 FILLER_29_227 ();
 sg13g2_decap_8 FILLER_29_234 ();
 sg13g2_decap_4 FILLER_29_241 ();
 sg13g2_fill_2 FILLER_29_245 ();
 sg13g2_fill_1 FILLER_29_259 ();
 sg13g2_fill_1 FILLER_29_305 ();
 sg13g2_fill_2 FILLER_29_341 ();
 sg13g2_fill_1 FILLER_29_343 ();
 sg13g2_decap_4 FILLER_29_367 ();
 sg13g2_fill_1 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_fill_2 FILLER_29_405 ();
 sg13g2_fill_2 FILLER_29_412 ();
 sg13g2_decap_8 FILLER_29_450 ();
 sg13g2_fill_2 FILLER_29_471 ();
 sg13g2_fill_1 FILLER_29_473 ();
 sg13g2_decap_8 FILLER_29_488 ();
 sg13g2_fill_1 FILLER_29_495 ();
 sg13g2_fill_1 FILLER_29_500 ();
 sg13g2_fill_1 FILLER_29_515 ();
 sg13g2_fill_1 FILLER_29_542 ();
 sg13g2_fill_2 FILLER_29_588 ();
 sg13g2_fill_1 FILLER_29_600 ();
 sg13g2_fill_2 FILLER_29_627 ();
 sg13g2_decap_4 FILLER_29_652 ();
 sg13g2_fill_2 FILLER_29_656 ();
 sg13g2_decap_8 FILLER_29_691 ();
 sg13g2_decap_8 FILLER_29_702 ();
 sg13g2_decap_8 FILLER_29_709 ();
 sg13g2_decap_8 FILLER_29_716 ();
 sg13g2_decap_8 FILLER_29_723 ();
 sg13g2_decap_8 FILLER_29_730 ();
 sg13g2_decap_8 FILLER_29_737 ();
 sg13g2_decap_8 FILLER_29_744 ();
 sg13g2_decap_8 FILLER_29_751 ();
 sg13g2_decap_8 FILLER_29_758 ();
 sg13g2_decap_8 FILLER_29_765 ();
 sg13g2_decap_8 FILLER_29_772 ();
 sg13g2_decap_8 FILLER_29_779 ();
 sg13g2_decap_8 FILLER_29_786 ();
 sg13g2_decap_8 FILLER_29_793 ();
 sg13g2_decap_8 FILLER_29_800 ();
 sg13g2_decap_8 FILLER_29_807 ();
 sg13g2_decap_8 FILLER_29_814 ();
 sg13g2_decap_8 FILLER_29_821 ();
 sg13g2_decap_8 FILLER_29_828 ();
 sg13g2_decap_8 FILLER_29_835 ();
 sg13g2_decap_8 FILLER_29_842 ();
 sg13g2_decap_8 FILLER_29_849 ();
 sg13g2_decap_4 FILLER_29_856 ();
 sg13g2_fill_2 FILLER_29_860 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_33 ();
 sg13g2_fill_1 FILLER_30_35 ();
 sg13g2_fill_2 FILLER_30_62 ();
 sg13g2_fill_1 FILLER_30_64 ();
 sg13g2_fill_2 FILLER_30_86 ();
 sg13g2_fill_1 FILLER_30_160 ();
 sg13g2_fill_1 FILLER_30_196 ();
 sg13g2_fill_1 FILLER_30_202 ();
 sg13g2_fill_2 FILLER_30_211 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_4 FILLER_30_224 ();
 sg13g2_fill_2 FILLER_30_228 ();
 sg13g2_fill_1 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_fill_2 FILLER_30_334 ();
 sg13g2_fill_2 FILLER_30_362 ();
 sg13g2_fill_1 FILLER_30_385 ();
 sg13g2_fill_2 FILLER_30_412 ();
 sg13g2_decap_4 FILLER_30_426 ();
 sg13g2_fill_2 FILLER_30_443 ();
 sg13g2_decap_8 FILLER_30_497 ();
 sg13g2_fill_2 FILLER_30_504 ();
 sg13g2_fill_1 FILLER_30_506 ();
 sg13g2_fill_2 FILLER_30_533 ();
 sg13g2_decap_4 FILLER_30_630 ();
 sg13g2_fill_2 FILLER_30_644 ();
 sg13g2_fill_1 FILLER_30_646 ();
 sg13g2_decap_8 FILLER_30_683 ();
 sg13g2_decap_8 FILLER_30_690 ();
 sg13g2_decap_8 FILLER_30_697 ();
 sg13g2_decap_8 FILLER_30_704 ();
 sg13g2_decap_8 FILLER_30_711 ();
 sg13g2_decap_8 FILLER_30_718 ();
 sg13g2_decap_8 FILLER_30_725 ();
 sg13g2_decap_8 FILLER_30_732 ();
 sg13g2_decap_8 FILLER_30_739 ();
 sg13g2_decap_8 FILLER_30_746 ();
 sg13g2_decap_8 FILLER_30_753 ();
 sg13g2_decap_8 FILLER_30_760 ();
 sg13g2_decap_8 FILLER_30_767 ();
 sg13g2_decap_8 FILLER_30_774 ();
 sg13g2_decap_8 FILLER_30_781 ();
 sg13g2_decap_8 FILLER_30_788 ();
 sg13g2_decap_8 FILLER_30_795 ();
 sg13g2_decap_8 FILLER_30_802 ();
 sg13g2_decap_8 FILLER_30_809 ();
 sg13g2_decap_8 FILLER_30_816 ();
 sg13g2_decap_8 FILLER_30_823 ();
 sg13g2_decap_8 FILLER_30_830 ();
 sg13g2_decap_8 FILLER_30_837 ();
 sg13g2_decap_8 FILLER_30_844 ();
 sg13g2_decap_8 FILLER_30_851 ();
 sg13g2_decap_4 FILLER_30_858 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_14 ();
 sg13g2_fill_2 FILLER_31_29 ();
 sg13g2_fill_1 FILLER_31_31 ();
 sg13g2_fill_2 FILLER_31_41 ();
 sg13g2_fill_2 FILLER_31_48 ();
 sg13g2_fill_1 FILLER_31_50 ();
 sg13g2_fill_2 FILLER_31_82 ();
 sg13g2_fill_1 FILLER_31_84 ();
 sg13g2_fill_1 FILLER_31_107 ();
 sg13g2_fill_2 FILLER_31_115 ();
 sg13g2_fill_1 FILLER_31_171 ();
 sg13g2_fill_2 FILLER_31_243 ();
 sg13g2_fill_1 FILLER_31_245 ();
 sg13g2_fill_1 FILLER_31_251 ();
 sg13g2_fill_1 FILLER_31_262 ();
 sg13g2_fill_2 FILLER_31_319 ();
 sg13g2_fill_1 FILLER_31_321 ();
 sg13g2_decap_4 FILLER_31_335 ();
 sg13g2_fill_2 FILLER_31_339 ();
 sg13g2_decap_4 FILLER_31_377 ();
 sg13g2_fill_2 FILLER_31_381 ();
 sg13g2_fill_1 FILLER_31_404 ();
 sg13g2_fill_2 FILLER_31_422 ();
 sg13g2_fill_1 FILLER_31_424 ();
 sg13g2_decap_8 FILLER_31_447 ();
 sg13g2_decap_8 FILLER_31_467 ();
 sg13g2_fill_2 FILLER_31_474 ();
 sg13g2_fill_1 FILLER_31_476 ();
 sg13g2_decap_8 FILLER_31_502 ();
 sg13g2_fill_2 FILLER_31_517 ();
 sg13g2_decap_8 FILLER_31_586 ();
 sg13g2_decap_8 FILLER_31_593 ();
 sg13g2_decap_4 FILLER_31_626 ();
 sg13g2_fill_2 FILLER_31_630 ();
 sg13g2_fill_2 FILLER_31_658 ();
 sg13g2_fill_1 FILLER_31_660 ();
 sg13g2_decap_8 FILLER_31_674 ();
 sg13g2_decap_8 FILLER_31_681 ();
 sg13g2_decap_8 FILLER_31_688 ();
 sg13g2_decap_8 FILLER_31_695 ();
 sg13g2_decap_8 FILLER_31_702 ();
 sg13g2_decap_8 FILLER_31_709 ();
 sg13g2_decap_8 FILLER_31_716 ();
 sg13g2_decap_8 FILLER_31_723 ();
 sg13g2_decap_8 FILLER_31_730 ();
 sg13g2_decap_8 FILLER_31_737 ();
 sg13g2_decap_8 FILLER_31_744 ();
 sg13g2_decap_8 FILLER_31_751 ();
 sg13g2_decap_8 FILLER_31_758 ();
 sg13g2_decap_8 FILLER_31_765 ();
 sg13g2_decap_8 FILLER_31_772 ();
 sg13g2_decap_8 FILLER_31_779 ();
 sg13g2_decap_8 FILLER_31_786 ();
 sg13g2_decap_8 FILLER_31_793 ();
 sg13g2_decap_8 FILLER_31_800 ();
 sg13g2_decap_8 FILLER_31_807 ();
 sg13g2_decap_8 FILLER_31_814 ();
 sg13g2_decap_8 FILLER_31_821 ();
 sg13g2_decap_8 FILLER_31_828 ();
 sg13g2_decap_8 FILLER_31_835 ();
 sg13g2_decap_8 FILLER_31_842 ();
 sg13g2_decap_8 FILLER_31_849 ();
 sg13g2_decap_4 FILLER_31_856 ();
 sg13g2_fill_2 FILLER_31_860 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_4 FILLER_32_14 ();
 sg13g2_fill_2 FILLER_32_63 ();
 sg13g2_fill_1 FILLER_32_65 ();
 sg13g2_fill_1 FILLER_32_176 ();
 sg13g2_fill_2 FILLER_32_182 ();
 sg13g2_fill_2 FILLER_32_210 ();
 sg13g2_fill_1 FILLER_32_230 ();
 sg13g2_fill_2 FILLER_32_275 ();
 sg13g2_fill_1 FILLER_32_277 ();
 sg13g2_fill_1 FILLER_32_356 ();
 sg13g2_fill_1 FILLER_32_370 ();
 sg13g2_fill_2 FILLER_32_384 ();
 sg13g2_fill_2 FILLER_32_412 ();
 sg13g2_fill_1 FILLER_32_414 ();
 sg13g2_fill_2 FILLER_32_469 ();
 sg13g2_fill_1 FILLER_32_471 ();
 sg13g2_decap_8 FILLER_32_519 ();
 sg13g2_fill_2 FILLER_32_526 ();
 sg13g2_decap_8 FILLER_32_575 ();
 sg13g2_decap_8 FILLER_32_582 ();
 sg13g2_decap_8 FILLER_32_615 ();
 sg13g2_decap_8 FILLER_32_626 ();
 sg13g2_fill_1 FILLER_32_633 ();
 sg13g2_fill_1 FILLER_32_642 ();
 sg13g2_fill_1 FILLER_32_647 ();
 sg13g2_decap_8 FILLER_32_657 ();
 sg13g2_decap_8 FILLER_32_664 ();
 sg13g2_decap_8 FILLER_32_671 ();
 sg13g2_decap_8 FILLER_32_678 ();
 sg13g2_decap_8 FILLER_32_685 ();
 sg13g2_decap_8 FILLER_32_692 ();
 sg13g2_decap_8 FILLER_32_699 ();
 sg13g2_decap_8 FILLER_32_706 ();
 sg13g2_decap_8 FILLER_32_713 ();
 sg13g2_decap_8 FILLER_32_720 ();
 sg13g2_decap_8 FILLER_32_727 ();
 sg13g2_decap_8 FILLER_32_734 ();
 sg13g2_decap_8 FILLER_32_741 ();
 sg13g2_decap_8 FILLER_32_748 ();
 sg13g2_decap_8 FILLER_32_755 ();
 sg13g2_decap_8 FILLER_32_762 ();
 sg13g2_decap_8 FILLER_32_769 ();
 sg13g2_decap_8 FILLER_32_776 ();
 sg13g2_decap_8 FILLER_32_783 ();
 sg13g2_decap_8 FILLER_32_790 ();
 sg13g2_decap_8 FILLER_32_797 ();
 sg13g2_decap_8 FILLER_32_804 ();
 sg13g2_decap_8 FILLER_32_811 ();
 sg13g2_decap_8 FILLER_32_818 ();
 sg13g2_decap_8 FILLER_32_825 ();
 sg13g2_decap_8 FILLER_32_832 ();
 sg13g2_decap_8 FILLER_32_839 ();
 sg13g2_decap_8 FILLER_32_846 ();
 sg13g2_decap_8 FILLER_32_853 ();
 sg13g2_fill_2 FILLER_32_860 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_fill_1 FILLER_33_76 ();
 sg13g2_fill_2 FILLER_33_86 ();
 sg13g2_fill_1 FILLER_33_88 ();
 sg13g2_fill_2 FILLER_33_120 ();
 sg13g2_fill_2 FILLER_33_164 ();
 sg13g2_fill_1 FILLER_33_166 ();
 sg13g2_fill_1 FILLER_33_205 ();
 sg13g2_fill_2 FILLER_33_248 ();
 sg13g2_fill_2 FILLER_33_303 ();
 sg13g2_fill_2 FILLER_33_314 ();
 sg13g2_fill_1 FILLER_33_316 ();
 sg13g2_decap_8 FILLER_33_321 ();
 sg13g2_decap_4 FILLER_33_328 ();
 sg13g2_fill_2 FILLER_33_332 ();
 sg13g2_decap_8 FILLER_33_342 ();
 sg13g2_fill_2 FILLER_33_349 ();
 sg13g2_decap_8 FILLER_33_377 ();
 sg13g2_decap_8 FILLER_33_384 ();
 sg13g2_decap_4 FILLER_33_391 ();
 sg13g2_fill_1 FILLER_33_395 ();
 sg13g2_fill_2 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_fill_1 FILLER_33_409 ();
 sg13g2_fill_2 FILLER_33_429 ();
 sg13g2_fill_1 FILLER_33_431 ();
 sg13g2_fill_1 FILLER_33_441 ();
 sg13g2_fill_2 FILLER_33_478 ();
 sg13g2_fill_1 FILLER_33_480 ();
 sg13g2_fill_1 FILLER_33_516 ();
 sg13g2_decap_4 FILLER_33_552 ();
 sg13g2_fill_1 FILLER_33_556 ();
 sg13g2_decap_8 FILLER_33_561 ();
 sg13g2_decap_4 FILLER_33_568 ();
 sg13g2_fill_2 FILLER_33_597 ();
 sg13g2_fill_1 FILLER_33_599 ();
 sg13g2_fill_2 FILLER_33_604 ();
 sg13g2_decap_8 FILLER_33_637 ();
 sg13g2_decap_8 FILLER_33_644 ();
 sg13g2_decap_8 FILLER_33_651 ();
 sg13g2_decap_8 FILLER_33_658 ();
 sg13g2_decap_8 FILLER_33_665 ();
 sg13g2_decap_8 FILLER_33_672 ();
 sg13g2_decap_8 FILLER_33_679 ();
 sg13g2_decap_8 FILLER_33_686 ();
 sg13g2_decap_8 FILLER_33_693 ();
 sg13g2_decap_8 FILLER_33_700 ();
 sg13g2_decap_8 FILLER_33_707 ();
 sg13g2_decap_8 FILLER_33_714 ();
 sg13g2_decap_8 FILLER_33_721 ();
 sg13g2_decap_8 FILLER_33_728 ();
 sg13g2_decap_8 FILLER_33_735 ();
 sg13g2_decap_8 FILLER_33_742 ();
 sg13g2_decap_8 FILLER_33_749 ();
 sg13g2_decap_8 FILLER_33_756 ();
 sg13g2_decap_8 FILLER_33_763 ();
 sg13g2_decap_8 FILLER_33_770 ();
 sg13g2_decap_8 FILLER_33_777 ();
 sg13g2_decap_8 FILLER_33_784 ();
 sg13g2_decap_8 FILLER_33_791 ();
 sg13g2_decap_8 FILLER_33_798 ();
 sg13g2_decap_8 FILLER_33_805 ();
 sg13g2_decap_8 FILLER_33_812 ();
 sg13g2_decap_8 FILLER_33_819 ();
 sg13g2_decap_8 FILLER_33_826 ();
 sg13g2_decap_8 FILLER_33_833 ();
 sg13g2_decap_8 FILLER_33_840 ();
 sg13g2_decap_8 FILLER_33_847 ();
 sg13g2_decap_8 FILLER_33_854 ();
 sg13g2_fill_1 FILLER_33_861 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_7 ();
 sg13g2_fill_2 FILLER_34_11 ();
 sg13g2_fill_1 FILLER_34_121 ();
 sg13g2_fill_1 FILLER_34_148 ();
 sg13g2_fill_1 FILLER_34_202 ();
 sg13g2_fill_2 FILLER_34_298 ();
 sg13g2_fill_1 FILLER_34_300 ();
 sg13g2_decap_8 FILLER_34_306 ();
 sg13g2_decap_8 FILLER_34_313 ();
 sg13g2_decap_4 FILLER_34_320 ();
 sg13g2_fill_1 FILLER_34_324 ();
 sg13g2_fill_1 FILLER_34_355 ();
 sg13g2_fill_1 FILLER_34_361 ();
 sg13g2_decap_4 FILLER_34_366 ();
 sg13g2_fill_2 FILLER_34_400 ();
 sg13g2_fill_1 FILLER_34_407 ();
 sg13g2_decap_4 FILLER_34_443 ();
 sg13g2_fill_2 FILLER_34_456 ();
 sg13g2_decap_8 FILLER_34_471 ();
 sg13g2_fill_1 FILLER_34_478 ();
 sg13g2_decap_8 FILLER_34_494 ();
 sg13g2_fill_2 FILLER_34_505 ();
 sg13g2_fill_1 FILLER_34_517 ();
 sg13g2_fill_2 FILLER_34_528 ();
 sg13g2_fill_2 FILLER_34_543 ();
 sg13g2_fill_1 FILLER_34_545 ();
 sg13g2_fill_2 FILLER_34_572 ();
 sg13g2_decap_8 FILLER_34_602 ();
 sg13g2_fill_1 FILLER_34_609 ();
 sg13g2_decap_8 FILLER_34_615 ();
 sg13g2_fill_2 FILLER_34_622 ();
 sg13g2_fill_1 FILLER_34_624 ();
 sg13g2_decap_8 FILLER_34_635 ();
 sg13g2_decap_8 FILLER_34_642 ();
 sg13g2_decap_8 FILLER_34_649 ();
 sg13g2_decap_8 FILLER_34_656 ();
 sg13g2_decap_8 FILLER_34_663 ();
 sg13g2_decap_8 FILLER_34_670 ();
 sg13g2_decap_8 FILLER_34_677 ();
 sg13g2_decap_8 FILLER_34_684 ();
 sg13g2_decap_8 FILLER_34_691 ();
 sg13g2_decap_8 FILLER_34_698 ();
 sg13g2_decap_8 FILLER_34_705 ();
 sg13g2_decap_8 FILLER_34_712 ();
 sg13g2_decap_8 FILLER_34_719 ();
 sg13g2_decap_8 FILLER_34_726 ();
 sg13g2_decap_8 FILLER_34_733 ();
 sg13g2_decap_8 FILLER_34_740 ();
 sg13g2_decap_8 FILLER_34_747 ();
 sg13g2_decap_8 FILLER_34_754 ();
 sg13g2_decap_8 FILLER_34_761 ();
 sg13g2_decap_8 FILLER_34_768 ();
 sg13g2_decap_8 FILLER_34_775 ();
 sg13g2_decap_8 FILLER_34_782 ();
 sg13g2_decap_8 FILLER_34_789 ();
 sg13g2_decap_8 FILLER_34_796 ();
 sg13g2_decap_8 FILLER_34_803 ();
 sg13g2_decap_8 FILLER_34_810 ();
 sg13g2_decap_8 FILLER_34_817 ();
 sg13g2_decap_8 FILLER_34_824 ();
 sg13g2_decap_8 FILLER_34_831 ();
 sg13g2_decap_8 FILLER_34_838 ();
 sg13g2_decap_8 FILLER_34_845 ();
 sg13g2_decap_8 FILLER_34_852 ();
 sg13g2_fill_2 FILLER_34_859 ();
 sg13g2_fill_1 FILLER_34_861 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_31 ();
 sg13g2_fill_2 FILLER_35_59 ();
 sg13g2_fill_1 FILLER_35_61 ();
 sg13g2_decap_8 FILLER_35_114 ();
 sg13g2_decap_4 FILLER_35_121 ();
 sg13g2_fill_1 FILLER_35_125 ();
 sg13g2_fill_2 FILLER_35_181 ();
 sg13g2_fill_2 FILLER_35_193 ();
 sg13g2_fill_2 FILLER_35_229 ();
 sg13g2_fill_2 FILLER_35_247 ();
 sg13g2_fill_2 FILLER_35_284 ();
 sg13g2_fill_1 FILLER_35_286 ();
 sg13g2_decap_4 FILLER_35_300 ();
 sg13g2_fill_2 FILLER_35_319 ();
 sg13g2_fill_2 FILLER_35_334 ();
 sg13g2_fill_1 FILLER_35_346 ();
 sg13g2_fill_1 FILLER_35_414 ();
 sg13g2_fill_2 FILLER_35_419 ();
 sg13g2_decap_4 FILLER_35_442 ();
 sg13g2_decap_4 FILLER_35_465 ();
 sg13g2_fill_1 FILLER_35_469 ();
 sg13g2_fill_2 FILLER_35_480 ();
 sg13g2_decap_8 FILLER_35_519 ();
 sg13g2_fill_2 FILLER_35_526 ();
 sg13g2_decap_4 FILLER_35_558 ();
 sg13g2_fill_2 FILLER_35_580 ();
 sg13g2_fill_2 FILLER_35_592 ();
 sg13g2_decap_4 FILLER_35_650 ();
 sg13g2_fill_1 FILLER_35_663 ();
 sg13g2_decap_8 FILLER_35_668 ();
 sg13g2_decap_8 FILLER_35_675 ();
 sg13g2_decap_8 FILLER_35_682 ();
 sg13g2_decap_8 FILLER_35_689 ();
 sg13g2_decap_8 FILLER_35_696 ();
 sg13g2_decap_8 FILLER_35_703 ();
 sg13g2_decap_8 FILLER_35_710 ();
 sg13g2_decap_8 FILLER_35_717 ();
 sg13g2_decap_8 FILLER_35_724 ();
 sg13g2_decap_8 FILLER_35_731 ();
 sg13g2_decap_8 FILLER_35_738 ();
 sg13g2_decap_8 FILLER_35_745 ();
 sg13g2_decap_8 FILLER_35_752 ();
 sg13g2_decap_8 FILLER_35_759 ();
 sg13g2_decap_8 FILLER_35_766 ();
 sg13g2_decap_8 FILLER_35_773 ();
 sg13g2_decap_8 FILLER_35_780 ();
 sg13g2_decap_8 FILLER_35_787 ();
 sg13g2_decap_8 FILLER_35_794 ();
 sg13g2_decap_8 FILLER_35_801 ();
 sg13g2_decap_8 FILLER_35_808 ();
 sg13g2_decap_8 FILLER_35_815 ();
 sg13g2_decap_8 FILLER_35_822 ();
 sg13g2_decap_8 FILLER_35_829 ();
 sg13g2_decap_8 FILLER_35_836 ();
 sg13g2_decap_8 FILLER_35_843 ();
 sg13g2_decap_8 FILLER_35_850 ();
 sg13g2_decap_4 FILLER_35_857 ();
 sg13g2_fill_1 FILLER_35_861 ();
 sg13g2_fill_1 FILLER_36_44 ();
 sg13g2_fill_2 FILLER_36_50 ();
 sg13g2_fill_2 FILLER_36_117 ();
 sg13g2_fill_1 FILLER_36_119 ();
 sg13g2_fill_1 FILLER_36_146 ();
 sg13g2_fill_1 FILLER_36_178 ();
 sg13g2_fill_2 FILLER_36_224 ();
 sg13g2_fill_1 FILLER_36_226 ();
 sg13g2_decap_4 FILLER_36_275 ();
 sg13g2_fill_1 FILLER_36_300 ();
 sg13g2_fill_1 FILLER_36_335 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_fill_1 FILLER_36_357 ();
 sg13g2_fill_1 FILLER_36_389 ();
 sg13g2_fill_2 FILLER_36_467 ();
 sg13g2_fill_1 FILLER_36_469 ();
 sg13g2_fill_2 FILLER_36_475 ();
 sg13g2_decap_8 FILLER_36_515 ();
 sg13g2_decap_8 FILLER_36_522 ();
 sg13g2_decap_8 FILLER_36_529 ();
 sg13g2_fill_1 FILLER_36_536 ();
 sg13g2_decap_4 FILLER_36_552 ();
 sg13g2_fill_1 FILLER_36_556 ();
 sg13g2_fill_2 FILLER_36_571 ();
 sg13g2_decap_8 FILLER_36_595 ();
 sg13g2_fill_2 FILLER_36_602 ();
 sg13g2_fill_2 FILLER_36_612 ();
 sg13g2_fill_1 FILLER_36_614 ();
 sg13g2_fill_2 FILLER_36_620 ();
 sg13g2_fill_2 FILLER_36_626 ();
 sg13g2_decap_8 FILLER_36_680 ();
 sg13g2_decap_8 FILLER_36_687 ();
 sg13g2_decap_8 FILLER_36_694 ();
 sg13g2_decap_8 FILLER_36_701 ();
 sg13g2_decap_8 FILLER_36_708 ();
 sg13g2_decap_8 FILLER_36_715 ();
 sg13g2_decap_8 FILLER_36_722 ();
 sg13g2_decap_8 FILLER_36_729 ();
 sg13g2_decap_8 FILLER_36_736 ();
 sg13g2_decap_8 FILLER_36_743 ();
 sg13g2_decap_8 FILLER_36_750 ();
 sg13g2_decap_8 FILLER_36_757 ();
 sg13g2_decap_8 FILLER_36_764 ();
 sg13g2_decap_8 FILLER_36_771 ();
 sg13g2_decap_8 FILLER_36_778 ();
 sg13g2_decap_8 FILLER_36_785 ();
 sg13g2_decap_8 FILLER_36_792 ();
 sg13g2_decap_8 FILLER_36_799 ();
 sg13g2_decap_8 FILLER_36_806 ();
 sg13g2_decap_8 FILLER_36_813 ();
 sg13g2_decap_8 FILLER_36_820 ();
 sg13g2_decap_8 FILLER_36_827 ();
 sg13g2_decap_8 FILLER_36_834 ();
 sg13g2_decap_8 FILLER_36_841 ();
 sg13g2_decap_8 FILLER_36_848 ();
 sg13g2_decap_8 FILLER_36_855 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_120 ();
 sg13g2_fill_1 FILLER_37_122 ();
 sg13g2_fill_2 FILLER_37_149 ();
 sg13g2_fill_1 FILLER_37_151 ();
 sg13g2_fill_2 FILLER_37_167 ();
 sg13g2_fill_1 FILLER_37_169 ();
 sg13g2_fill_2 FILLER_37_185 ();
 sg13g2_fill_2 FILLER_37_192 ();
 sg13g2_fill_1 FILLER_37_194 ();
 sg13g2_fill_1 FILLER_37_223 ();
 sg13g2_fill_1 FILLER_37_230 ();
 sg13g2_decap_8 FILLER_37_270 ();
 sg13g2_decap_4 FILLER_37_277 ();
 sg13g2_fill_1 FILLER_37_281 ();
 sg13g2_fill_2 FILLER_37_299 ();
 sg13g2_decap_4 FILLER_37_319 ();
 sg13g2_fill_1 FILLER_37_323 ();
 sg13g2_decap_4 FILLER_37_335 ();
 sg13g2_decap_8 FILLER_37_352 ();
 sg13g2_decap_8 FILLER_37_359 ();
 sg13g2_decap_4 FILLER_37_366 ();
 sg13g2_decap_4 FILLER_37_385 ();
 sg13g2_fill_1 FILLER_37_389 ();
 sg13g2_decap_4 FILLER_37_397 ();
 sg13g2_fill_2 FILLER_37_401 ();
 sg13g2_decap_8 FILLER_37_416 ();
 sg13g2_fill_2 FILLER_37_427 ();
 sg13g2_fill_2 FILLER_37_433 ();
 sg13g2_decap_8 FILLER_37_441 ();
 sg13g2_decap_4 FILLER_37_448 ();
 sg13g2_fill_1 FILLER_37_452 ();
 sg13g2_decap_4 FILLER_37_457 ();
 sg13g2_decap_4 FILLER_37_465 ();
 sg13g2_fill_2 FILLER_37_497 ();
 sg13g2_fill_1 FILLER_37_499 ();
 sg13g2_fill_2 FILLER_37_507 ();
 sg13g2_fill_1 FILLER_37_509 ();
 sg13g2_decap_8 FILLER_37_594 ();
 sg13g2_fill_2 FILLER_37_601 ();
 sg13g2_fill_1 FILLER_37_603 ();
 sg13g2_fill_1 FILLER_37_621 ();
 sg13g2_decap_8 FILLER_37_648 ();
 sg13g2_decap_4 FILLER_37_664 ();
 sg13g2_fill_2 FILLER_37_668 ();
 sg13g2_decap_8 FILLER_37_679 ();
 sg13g2_decap_8 FILLER_37_686 ();
 sg13g2_decap_8 FILLER_37_693 ();
 sg13g2_decap_8 FILLER_37_700 ();
 sg13g2_decap_8 FILLER_37_707 ();
 sg13g2_decap_8 FILLER_37_714 ();
 sg13g2_decap_8 FILLER_37_721 ();
 sg13g2_decap_8 FILLER_37_728 ();
 sg13g2_decap_8 FILLER_37_735 ();
 sg13g2_decap_8 FILLER_37_742 ();
 sg13g2_decap_8 FILLER_37_749 ();
 sg13g2_decap_8 FILLER_37_756 ();
 sg13g2_decap_8 FILLER_37_763 ();
 sg13g2_decap_8 FILLER_37_770 ();
 sg13g2_decap_8 FILLER_37_777 ();
 sg13g2_decap_8 FILLER_37_784 ();
 sg13g2_decap_8 FILLER_37_791 ();
 sg13g2_decap_8 FILLER_37_798 ();
 sg13g2_decap_8 FILLER_37_805 ();
 sg13g2_decap_8 FILLER_37_812 ();
 sg13g2_decap_8 FILLER_37_819 ();
 sg13g2_decap_8 FILLER_37_826 ();
 sg13g2_decap_8 FILLER_37_833 ();
 sg13g2_decap_8 FILLER_37_840 ();
 sg13g2_decap_8 FILLER_37_847 ();
 sg13g2_decap_8 FILLER_37_854 ();
 sg13g2_fill_1 FILLER_37_861 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_28 ();
 sg13g2_fill_1 FILLER_38_38 ();
 sg13g2_fill_2 FILLER_38_84 ();
 sg13g2_fill_2 FILLER_38_121 ();
 sg13g2_fill_1 FILLER_38_123 ();
 sg13g2_fill_2 FILLER_38_132 ();
 sg13g2_fill_1 FILLER_38_138 ();
 sg13g2_fill_1 FILLER_38_148 ();
 sg13g2_fill_1 FILLER_38_167 ();
 sg13g2_fill_2 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_296 ();
 sg13g2_decap_8 FILLER_38_303 ();
 sg13g2_decap_8 FILLER_38_310 ();
 sg13g2_fill_2 FILLER_38_317 ();
 sg13g2_decap_8 FILLER_38_359 ();
 sg13g2_fill_2 FILLER_38_366 ();
 sg13g2_fill_1 FILLER_38_368 ();
 sg13g2_fill_2 FILLER_38_402 ();
 sg13g2_decap_4 FILLER_38_410 ();
 sg13g2_fill_2 FILLER_38_440 ();
 sg13g2_fill_2 FILLER_38_481 ();
 sg13g2_fill_1 FILLER_38_493 ();
 sg13g2_decap_8 FILLER_38_513 ();
 sg13g2_decap_4 FILLER_38_520 ();
 sg13g2_fill_2 FILLER_38_529 ();
 sg13g2_decap_4 FILLER_38_539 ();
 sg13g2_fill_1 FILLER_38_543 ();
 sg13g2_decap_4 FILLER_38_552 ();
 sg13g2_fill_1 FILLER_38_556 ();
 sg13g2_decap_8 FILLER_38_561 ();
 sg13g2_fill_1 FILLER_38_568 ();
 sg13g2_decap_4 FILLER_38_627 ();
 sg13g2_fill_2 FILLER_38_631 ();
 sg13g2_decap_8 FILLER_38_637 ();
 sg13g2_decap_8 FILLER_38_696 ();
 sg13g2_decap_8 FILLER_38_703 ();
 sg13g2_decap_8 FILLER_38_710 ();
 sg13g2_decap_8 FILLER_38_717 ();
 sg13g2_decap_8 FILLER_38_724 ();
 sg13g2_decap_8 FILLER_38_731 ();
 sg13g2_decap_8 FILLER_38_738 ();
 sg13g2_decap_8 FILLER_38_745 ();
 sg13g2_decap_8 FILLER_38_752 ();
 sg13g2_decap_8 FILLER_38_759 ();
 sg13g2_decap_8 FILLER_38_766 ();
 sg13g2_decap_8 FILLER_38_773 ();
 sg13g2_decap_8 FILLER_38_780 ();
 sg13g2_decap_8 FILLER_38_787 ();
 sg13g2_decap_8 FILLER_38_794 ();
 sg13g2_decap_8 FILLER_38_801 ();
 sg13g2_decap_8 FILLER_38_808 ();
 sg13g2_decap_8 FILLER_38_815 ();
 sg13g2_decap_8 FILLER_38_822 ();
 sg13g2_decap_8 FILLER_38_829 ();
 sg13g2_decap_8 FILLER_38_836 ();
 sg13g2_decap_8 FILLER_38_843 ();
 sg13g2_decap_8 FILLER_38_850 ();
 sg13g2_decap_4 FILLER_38_857 ();
 sg13g2_fill_1 FILLER_38_861 ();
 sg13g2_fill_1 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_27 ();
 sg13g2_fill_1 FILLER_39_29 ();
 sg13g2_fill_1 FILLER_39_58 ();
 sg13g2_fill_2 FILLER_39_73 ();
 sg13g2_fill_1 FILLER_39_75 ();
 sg13g2_fill_2 FILLER_39_102 ();
 sg13g2_fill_1 FILLER_39_104 ();
 sg13g2_decap_8 FILLER_39_139 ();
 sg13g2_fill_2 FILLER_39_172 ();
 sg13g2_fill_2 FILLER_39_225 ();
 sg13g2_fill_2 FILLER_39_236 ();
 sg13g2_fill_1 FILLER_39_280 ();
 sg13g2_decap_8 FILLER_39_313 ();
 sg13g2_fill_2 FILLER_39_320 ();
 sg13g2_fill_2 FILLER_39_335 ();
 sg13g2_fill_2 FILLER_39_352 ();
 sg13g2_fill_1 FILLER_39_354 ();
 sg13g2_decap_4 FILLER_39_360 ();
 sg13g2_decap_8 FILLER_39_367 ();
 sg13g2_decap_4 FILLER_39_374 ();
 sg13g2_fill_1 FILLER_39_378 ();
 sg13g2_fill_2 FILLER_39_395 ();
 sg13g2_fill_1 FILLER_39_397 ();
 sg13g2_decap_8 FILLER_39_404 ();
 sg13g2_fill_1 FILLER_39_411 ();
 sg13g2_decap_4 FILLER_39_420 ();
 sg13g2_fill_1 FILLER_39_424 ();
 sg13g2_decap_8 FILLER_39_429 ();
 sg13g2_fill_2 FILLER_39_436 ();
 sg13g2_decap_4 FILLER_39_441 ();
 sg13g2_fill_2 FILLER_39_453 ();
 sg13g2_decap_8 FILLER_39_461 ();
 sg13g2_fill_1 FILLER_39_468 ();
 sg13g2_fill_2 FILLER_39_476 ();
 sg13g2_decap_4 FILLER_39_522 ();
 sg13g2_decap_4 FILLER_39_543 ();
 sg13g2_fill_2 FILLER_39_573 ();
 sg13g2_fill_1 FILLER_39_575 ();
 sg13g2_decap_4 FILLER_39_580 ();
 sg13g2_fill_1 FILLER_39_589 ();
 sg13g2_decap_8 FILLER_39_593 ();
 sg13g2_decap_8 FILLER_39_600 ();
 sg13g2_fill_2 FILLER_39_607 ();
 sg13g2_fill_1 FILLER_39_609 ();
 sg13g2_decap_4 FILLER_39_628 ();
 sg13g2_fill_1 FILLER_39_632 ();
 sg13g2_fill_1 FILLER_39_659 ();
 sg13g2_decap_8 FILLER_39_688 ();
 sg13g2_decap_8 FILLER_39_695 ();
 sg13g2_decap_8 FILLER_39_702 ();
 sg13g2_decap_8 FILLER_39_709 ();
 sg13g2_decap_8 FILLER_39_716 ();
 sg13g2_decap_8 FILLER_39_723 ();
 sg13g2_decap_8 FILLER_39_730 ();
 sg13g2_decap_8 FILLER_39_737 ();
 sg13g2_decap_8 FILLER_39_744 ();
 sg13g2_decap_8 FILLER_39_751 ();
 sg13g2_decap_8 FILLER_39_758 ();
 sg13g2_decap_8 FILLER_39_765 ();
 sg13g2_decap_8 FILLER_39_772 ();
 sg13g2_decap_8 FILLER_39_779 ();
 sg13g2_decap_8 FILLER_39_786 ();
 sg13g2_decap_8 FILLER_39_793 ();
 sg13g2_decap_8 FILLER_39_800 ();
 sg13g2_decap_8 FILLER_39_807 ();
 sg13g2_decap_8 FILLER_39_814 ();
 sg13g2_decap_8 FILLER_39_821 ();
 sg13g2_decap_8 FILLER_39_828 ();
 sg13g2_decap_8 FILLER_39_835 ();
 sg13g2_decap_8 FILLER_39_842 ();
 sg13g2_decap_8 FILLER_39_849 ();
 sg13g2_decap_4 FILLER_39_856 ();
 sg13g2_fill_2 FILLER_39_860 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_67 ();
 sg13g2_fill_2 FILLER_40_84 ();
 sg13g2_fill_1 FILLER_40_86 ();
 sg13g2_fill_1 FILLER_40_156 ();
 sg13g2_fill_2 FILLER_40_161 ();
 sg13g2_fill_1 FILLER_40_163 ();
 sg13g2_fill_1 FILLER_40_186 ();
 sg13g2_fill_1 FILLER_40_230 ();
 sg13g2_fill_1 FILLER_40_257 ();
 sg13g2_fill_2 FILLER_40_261 ();
 sg13g2_fill_1 FILLER_40_263 ();
 sg13g2_fill_2 FILLER_40_297 ();
 sg13g2_fill_1 FILLER_40_299 ();
 sg13g2_decap_4 FILLER_40_317 ();
 sg13g2_fill_1 FILLER_40_321 ();
 sg13g2_fill_2 FILLER_40_327 ();
 sg13g2_decap_4 FILLER_40_334 ();
 sg13g2_decap_8 FILLER_40_346 ();
 sg13g2_decap_8 FILLER_40_381 ();
 sg13g2_decap_4 FILLER_40_388 ();
 sg13g2_fill_2 FILLER_40_392 ();
 sg13g2_fill_2 FILLER_40_404 ();
 sg13g2_fill_1 FILLER_40_406 ();
 sg13g2_fill_2 FILLER_40_418 ();
 sg13g2_fill_1 FILLER_40_420 ();
 sg13g2_fill_2 FILLER_40_433 ();
 sg13g2_fill_1 FILLER_40_435 ();
 sg13g2_decap_4 FILLER_40_462 ();
 sg13g2_fill_1 FILLER_40_466 ();
 sg13g2_decap_4 FILLER_40_487 ();
 sg13g2_fill_1 FILLER_40_491 ();
 sg13g2_decap_4 FILLER_40_500 ();
 sg13g2_fill_2 FILLER_40_504 ();
 sg13g2_decap_4 FILLER_40_515 ();
 sg13g2_fill_2 FILLER_40_528 ();
 sg13g2_decap_4 FILLER_40_533 ();
 sg13g2_decap_8 FILLER_40_543 ();
 sg13g2_decap_8 FILLER_40_648 ();
 sg13g2_fill_1 FILLER_40_655 ();
 sg13g2_decap_8 FILLER_40_691 ();
 sg13g2_decap_8 FILLER_40_698 ();
 sg13g2_decap_8 FILLER_40_705 ();
 sg13g2_decap_8 FILLER_40_712 ();
 sg13g2_decap_8 FILLER_40_719 ();
 sg13g2_decap_8 FILLER_40_726 ();
 sg13g2_decap_8 FILLER_40_733 ();
 sg13g2_decap_8 FILLER_40_740 ();
 sg13g2_decap_8 FILLER_40_747 ();
 sg13g2_decap_8 FILLER_40_754 ();
 sg13g2_decap_8 FILLER_40_761 ();
 sg13g2_decap_8 FILLER_40_768 ();
 sg13g2_decap_8 FILLER_40_775 ();
 sg13g2_decap_8 FILLER_40_782 ();
 sg13g2_decap_8 FILLER_40_789 ();
 sg13g2_decap_8 FILLER_40_796 ();
 sg13g2_decap_8 FILLER_40_803 ();
 sg13g2_decap_8 FILLER_40_810 ();
 sg13g2_decap_8 FILLER_40_817 ();
 sg13g2_decap_8 FILLER_40_824 ();
 sg13g2_decap_8 FILLER_40_831 ();
 sg13g2_decap_8 FILLER_40_838 ();
 sg13g2_decap_8 FILLER_40_845 ();
 sg13g2_decap_8 FILLER_40_852 ();
 sg13g2_fill_2 FILLER_40_859 ();
 sg13g2_fill_1 FILLER_40_861 ();
 sg13g2_fill_1 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_27 ();
 sg13g2_fill_2 FILLER_41_38 ();
 sg13g2_fill_1 FILLER_41_58 ();
 sg13g2_fill_1 FILLER_41_68 ();
 sg13g2_fill_2 FILLER_41_107 ();
 sg13g2_fill_1 FILLER_41_109 ();
 sg13g2_fill_2 FILLER_41_146 ();
 sg13g2_fill_1 FILLER_41_162 ();
 sg13g2_fill_2 FILLER_41_198 ();
 sg13g2_fill_1 FILLER_41_200 ();
 sg13g2_fill_1 FILLER_41_211 ();
 sg13g2_decap_8 FILLER_41_251 ();
 sg13g2_decap_8 FILLER_41_258 ();
 sg13g2_fill_2 FILLER_41_265 ();
 sg13g2_fill_1 FILLER_41_267 ();
 sg13g2_fill_2 FILLER_41_283 ();
 sg13g2_fill_1 FILLER_41_285 ();
 sg13g2_decap_4 FILLER_41_295 ();
 sg13g2_fill_2 FILLER_41_299 ();
 sg13g2_fill_1 FILLER_41_321 ();
 sg13g2_fill_1 FILLER_41_327 ();
 sg13g2_decap_4 FILLER_41_349 ();
 sg13g2_fill_1 FILLER_41_353 ();
 sg13g2_fill_2 FILLER_41_380 ();
 sg13g2_decap_8 FILLER_41_413 ();
 sg13g2_decap_4 FILLER_41_425 ();
 sg13g2_fill_2 FILLER_41_429 ();
 sg13g2_fill_2 FILLER_41_435 ();
 sg13g2_fill_2 FILLER_41_447 ();
 sg13g2_fill_1 FILLER_41_449 ();
 sg13g2_fill_1 FILLER_41_455 ();
 sg13g2_fill_2 FILLER_41_461 ();
 sg13g2_fill_1 FILLER_41_463 ();
 sg13g2_decap_8 FILLER_41_469 ();
 sg13g2_fill_1 FILLER_41_476 ();
 sg13g2_fill_1 FILLER_41_497 ();
 sg13g2_fill_2 FILLER_41_501 ();
 sg13g2_fill_1 FILLER_41_503 ();
 sg13g2_decap_8 FILLER_41_508 ();
 sg13g2_decap_4 FILLER_41_519 ();
 sg13g2_fill_2 FILLER_41_523 ();
 sg13g2_decap_4 FILLER_41_569 ();
 sg13g2_fill_1 FILLER_41_573 ();
 sg13g2_decap_8 FILLER_41_578 ();
 sg13g2_decap_4 FILLER_41_585 ();
 sg13g2_fill_1 FILLER_41_595 ();
 sg13g2_fill_2 FILLER_41_606 ();
 sg13g2_decap_4 FILLER_41_623 ();
 sg13g2_fill_2 FILLER_41_627 ();
 sg13g2_decap_4 FILLER_41_633 ();
 sg13g2_fill_1 FILLER_41_648 ();
 sg13g2_decap_8 FILLER_41_675 ();
 sg13g2_decap_8 FILLER_41_682 ();
 sg13g2_decap_8 FILLER_41_689 ();
 sg13g2_decap_8 FILLER_41_696 ();
 sg13g2_decap_8 FILLER_41_703 ();
 sg13g2_decap_8 FILLER_41_710 ();
 sg13g2_fill_1 FILLER_41_717 ();
 sg13g2_decap_8 FILLER_41_744 ();
 sg13g2_decap_8 FILLER_41_751 ();
 sg13g2_decap_8 FILLER_41_758 ();
 sg13g2_decap_8 FILLER_41_765 ();
 sg13g2_decap_8 FILLER_41_772 ();
 sg13g2_decap_8 FILLER_41_779 ();
 sg13g2_decap_8 FILLER_41_786 ();
 sg13g2_decap_8 FILLER_41_793 ();
 sg13g2_decap_8 FILLER_41_800 ();
 sg13g2_decap_8 FILLER_41_807 ();
 sg13g2_decap_8 FILLER_41_814 ();
 sg13g2_decap_8 FILLER_41_821 ();
 sg13g2_decap_8 FILLER_41_828 ();
 sg13g2_decap_8 FILLER_41_835 ();
 sg13g2_decap_8 FILLER_41_842 ();
 sg13g2_decap_8 FILLER_41_849 ();
 sg13g2_decap_4 FILLER_41_856 ();
 sg13g2_fill_2 FILLER_41_860 ();
 sg13g2_decap_4 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_4 ();
 sg13g2_fill_2 FILLER_42_35 ();
 sg13g2_fill_1 FILLER_42_56 ();
 sg13g2_fill_1 FILLER_42_62 ();
 sg13g2_fill_1 FILLER_42_177 ();
 sg13g2_decap_8 FILLER_42_183 ();
 sg13g2_decap_4 FILLER_42_213 ();
 sg13g2_fill_1 FILLER_42_217 ();
 sg13g2_decap_8 FILLER_42_261 ();
 sg13g2_fill_1 FILLER_42_268 ();
 sg13g2_fill_2 FILLER_42_296 ();
 sg13g2_decap_8 FILLER_42_313 ();
 sg13g2_fill_1 FILLER_42_320 ();
 sg13g2_fill_1 FILLER_42_325 ();
 sg13g2_fill_1 FILLER_42_344 ();
 sg13g2_fill_1 FILLER_42_371 ();
 sg13g2_decap_8 FILLER_42_377 ();
 sg13g2_fill_2 FILLER_42_384 ();
 sg13g2_fill_1 FILLER_42_396 ();
 sg13g2_fill_2 FILLER_42_412 ();
 sg13g2_fill_1 FILLER_42_414 ();
 sg13g2_decap_4 FILLER_42_426 ();
 sg13g2_decap_8 FILLER_42_461 ();
 sg13g2_fill_2 FILLER_42_468 ();
 sg13g2_fill_1 FILLER_42_470 ();
 sg13g2_decap_8 FILLER_42_478 ();
 sg13g2_fill_1 FILLER_42_485 ();
 sg13g2_decap_8 FILLER_42_542 ();
 sg13g2_decap_4 FILLER_42_549 ();
 sg13g2_fill_2 FILLER_42_553 ();
 sg13g2_decap_8 FILLER_42_580 ();
 sg13g2_decap_4 FILLER_42_587 ();
 sg13g2_fill_1 FILLER_42_591 ();
 sg13g2_decap_4 FILLER_42_610 ();
 sg13g2_fill_2 FILLER_42_614 ();
 sg13g2_fill_2 FILLER_42_637 ();
 sg13g2_decap_8 FILLER_42_647 ();
 sg13g2_decap_4 FILLER_42_654 ();
 sg13g2_fill_2 FILLER_42_658 ();
 sg13g2_fill_2 FILLER_42_674 ();
 sg13g2_decap_4 FILLER_42_681 ();
 sg13g2_decap_4 FILLER_42_689 ();
 sg13g2_fill_2 FILLER_42_719 ();
 sg13g2_fill_2 FILLER_42_726 ();
 sg13g2_fill_1 FILLER_42_728 ();
 sg13g2_fill_2 FILLER_42_737 ();
 sg13g2_decap_8 FILLER_42_748 ();
 sg13g2_decap_4 FILLER_42_755 ();
 sg13g2_decap_8 FILLER_42_764 ();
 sg13g2_decap_4 FILLER_42_771 ();
 sg13g2_fill_1 FILLER_42_797 ();
 sg13g2_decap_4 FILLER_42_803 ();
 sg13g2_decap_8 FILLER_42_811 ();
 sg13g2_decap_8 FILLER_42_818 ();
 sg13g2_decap_8 FILLER_42_825 ();
 sg13g2_decap_8 FILLER_42_832 ();
 sg13g2_decap_8 FILLER_42_839 ();
 sg13g2_decap_8 FILLER_42_846 ();
 sg13g2_decap_8 FILLER_42_853 ();
 sg13g2_fill_2 FILLER_42_860 ();
 sg13g2_fill_1 FILLER_43_35 ();
 sg13g2_fill_2 FILLER_43_110 ();
 sg13g2_fill_1 FILLER_43_112 ();
 sg13g2_decap_4 FILLER_43_139 ();
 sg13g2_fill_2 FILLER_43_143 ();
 sg13g2_fill_2 FILLER_43_157 ();
 sg13g2_decap_4 FILLER_43_194 ();
 sg13g2_fill_2 FILLER_43_202 ();
 sg13g2_fill_1 FILLER_43_204 ();
 sg13g2_fill_1 FILLER_43_209 ();
 sg13g2_decap_4 FILLER_43_240 ();
 sg13g2_fill_2 FILLER_43_244 ();
 sg13g2_decap_8 FILLER_43_250 ();
 sg13g2_decap_8 FILLER_43_257 ();
 sg13g2_fill_1 FILLER_43_264 ();
 sg13g2_decap_4 FILLER_43_278 ();
 sg13g2_fill_2 FILLER_43_289 ();
 sg13g2_fill_2 FILLER_43_296 ();
 sg13g2_fill_1 FILLER_43_313 ();
 sg13g2_decap_8 FILLER_43_347 ();
 sg13g2_decap_8 FILLER_43_354 ();
 sg13g2_decap_8 FILLER_43_361 ();
 sg13g2_fill_1 FILLER_43_416 ();
 sg13g2_fill_2 FILLER_43_426 ();
 sg13g2_fill_1 FILLER_43_428 ();
 sg13g2_fill_2 FILLER_43_441 ();
 sg13g2_fill_1 FILLER_43_477 ();
 sg13g2_decap_4 FILLER_43_488 ();
 sg13g2_fill_1 FILLER_43_506 ();
 sg13g2_fill_2 FILLER_43_520 ();
 sg13g2_fill_1 FILLER_43_537 ();
 sg13g2_fill_2 FILLER_43_558 ();
 sg13g2_fill_1 FILLER_43_560 ();
 sg13g2_fill_1 FILLER_43_589 ();
 sg13g2_fill_2 FILLER_43_612 ();
 sg13g2_fill_1 FILLER_43_614 ();
 sg13g2_fill_2 FILLER_43_623 ();
 sg13g2_fill_1 FILLER_43_625 ();
 sg13g2_decap_4 FILLER_43_643 ();
 sg13g2_fill_1 FILLER_43_673 ();
 sg13g2_fill_1 FILLER_43_700 ();
 sg13g2_fill_2 FILLER_43_728 ();
 sg13g2_fill_1 FILLER_43_730 ();
 sg13g2_decap_8 FILLER_43_735 ();
 sg13g2_fill_2 FILLER_43_794 ();
 sg13g2_decap_8 FILLER_43_822 ();
 sg13g2_decap_8 FILLER_43_829 ();
 sg13g2_decap_8 FILLER_43_836 ();
 sg13g2_decap_8 FILLER_43_843 ();
 sg13g2_decap_8 FILLER_43_850 ();
 sg13g2_decap_4 FILLER_43_857 ();
 sg13g2_fill_1 FILLER_43_861 ();
 sg13g2_fill_1 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_23 ();
 sg13g2_fill_1 FILLER_44_25 ();
 sg13g2_fill_2 FILLER_44_45 ();
 sg13g2_fill_2 FILLER_44_65 ();
 sg13g2_fill_1 FILLER_44_67 ();
 sg13g2_fill_1 FILLER_44_73 ();
 sg13g2_fill_2 FILLER_44_87 ();
 sg13g2_fill_1 FILLER_44_89 ();
 sg13g2_fill_2 FILLER_44_191 ();
 sg13g2_fill_1 FILLER_44_193 ();
 sg13g2_fill_2 FILLER_44_220 ();
 sg13g2_decap_4 FILLER_44_231 ();
 sg13g2_fill_2 FILLER_44_235 ();
 sg13g2_decap_4 FILLER_44_263 ();
 sg13g2_fill_1 FILLER_44_267 ();
 sg13g2_fill_2 FILLER_44_304 ();
 sg13g2_decap_8 FILLER_44_311 ();
 sg13g2_fill_2 FILLER_44_318 ();
 sg13g2_fill_1 FILLER_44_320 ();
 sg13g2_fill_1 FILLER_44_337 ();
 sg13g2_fill_2 FILLER_44_355 ();
 sg13g2_decap_8 FILLER_44_375 ();
 sg13g2_decap_4 FILLER_44_382 ();
 sg13g2_fill_1 FILLER_44_386 ();
 sg13g2_decap_8 FILLER_44_424 ();
 sg13g2_decap_8 FILLER_44_431 ();
 sg13g2_decap_8 FILLER_44_438 ();
 sg13g2_decap_8 FILLER_44_445 ();
 sg13g2_decap_8 FILLER_44_452 ();
 sg13g2_fill_2 FILLER_44_459 ();
 sg13g2_fill_1 FILLER_44_461 ();
 sg13g2_decap_4 FILLER_44_466 ();
 sg13g2_fill_2 FILLER_44_470 ();
 sg13g2_fill_2 FILLER_44_506 ();
 sg13g2_decap_4 FILLER_44_526 ();
 sg13g2_fill_1 FILLER_44_543 ();
 sg13g2_decap_8 FILLER_44_559 ();
 sg13g2_decap_4 FILLER_44_566 ();
 sg13g2_fill_2 FILLER_44_570 ();
 sg13g2_decap_8 FILLER_44_582 ();
 sg13g2_decap_8 FILLER_44_589 ();
 sg13g2_fill_1 FILLER_44_596 ();
 sg13g2_fill_2 FILLER_44_626 ();
 sg13g2_fill_1 FILLER_44_628 ();
 sg13g2_decap_4 FILLER_44_642 ();
 sg13g2_decap_4 FILLER_44_650 ();
 sg13g2_fill_2 FILLER_44_664 ();
 sg13g2_fill_1 FILLER_44_666 ();
 sg13g2_fill_1 FILLER_44_689 ();
 sg13g2_fill_2 FILLER_44_716 ();
 sg13g2_fill_1 FILLER_44_718 ();
 sg13g2_fill_1 FILLER_44_766 ();
 sg13g2_fill_2 FILLER_44_780 ();
 sg13g2_fill_1 FILLER_44_782 ();
 sg13g2_fill_1 FILLER_44_796 ();
 sg13g2_fill_2 FILLER_44_805 ();
 sg13g2_fill_1 FILLER_44_807 ();
 sg13g2_decap_8 FILLER_44_834 ();
 sg13g2_decap_8 FILLER_44_841 ();
 sg13g2_decap_8 FILLER_44_848 ();
 sg13g2_decap_8 FILLER_44_855 ();
 sg13g2_fill_1 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_83 ();
 sg13g2_fill_1 FILLER_45_108 ();
 sg13g2_fill_2 FILLER_45_134 ();
 sg13g2_fill_1 FILLER_45_162 ();
 sg13g2_fill_2 FILLER_45_172 ();
 sg13g2_fill_2 FILLER_45_197 ();
 sg13g2_fill_1 FILLER_45_199 ();
 sg13g2_decap_4 FILLER_45_204 ();
 sg13g2_fill_2 FILLER_45_208 ();
 sg13g2_decap_8 FILLER_45_256 ();
 sg13g2_decap_4 FILLER_45_263 ();
 sg13g2_decap_8 FILLER_45_271 ();
 sg13g2_fill_2 FILLER_45_278 ();
 sg13g2_fill_1 FILLER_45_280 ();
 sg13g2_fill_1 FILLER_45_292 ();
 sg13g2_fill_1 FILLER_45_312 ();
 sg13g2_fill_2 FILLER_45_318 ();
 sg13g2_fill_1 FILLER_45_347 ();
 sg13g2_decap_4 FILLER_45_363 ();
 sg13g2_fill_2 FILLER_45_367 ();
 sg13g2_decap_8 FILLER_45_398 ();
 sg13g2_decap_4 FILLER_45_405 ();
 sg13g2_fill_1 FILLER_45_461 ();
 sg13g2_fill_1 FILLER_45_466 ();
 sg13g2_fill_1 FILLER_45_476 ();
 sg13g2_fill_1 FILLER_45_492 ();
 sg13g2_decap_4 FILLER_45_524 ();
 sg13g2_fill_2 FILLER_45_591 ();
 sg13g2_fill_1 FILLER_45_593 ();
 sg13g2_fill_1 FILLER_45_620 ();
 sg13g2_fill_2 FILLER_45_652 ();
 sg13g2_decap_4 FILLER_45_660 ();
 sg13g2_fill_1 FILLER_45_664 ();
 sg13g2_fill_2 FILLER_45_699 ();
 sg13g2_fill_1 FILLER_45_701 ();
 sg13g2_decap_4 FILLER_45_753 ();
 sg13g2_fill_1 FILLER_45_770 ();
 sg13g2_decap_8 FILLER_45_850 ();
 sg13g2_decap_4 FILLER_45_857 ();
 sg13g2_fill_1 FILLER_45_861 ();
 sg13g2_decap_4 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_4 ();
 sg13g2_fill_2 FILLER_46_31 ();
 sg13g2_fill_1 FILLER_46_33 ();
 sg13g2_fill_2 FILLER_46_66 ();
 sg13g2_fill_1 FILLER_46_68 ();
 sg13g2_fill_1 FILLER_46_78 ();
 sg13g2_fill_1 FILLER_46_114 ();
 sg13g2_fill_2 FILLER_46_167 ();
 sg13g2_fill_1 FILLER_46_169 ();
 sg13g2_fill_2 FILLER_46_187 ();
 sg13g2_fill_1 FILLER_46_221 ();
 sg13g2_fill_2 FILLER_46_231 ();
 sg13g2_fill_1 FILLER_46_233 ();
 sg13g2_decap_4 FILLER_46_251 ();
 sg13g2_fill_1 FILLER_46_255 ();
 sg13g2_decap_8 FILLER_46_282 ();
 sg13g2_decap_8 FILLER_46_289 ();
 sg13g2_fill_2 FILLER_46_296 ();
 sg13g2_decap_8 FILLER_46_312 ();
 sg13g2_decap_8 FILLER_46_319 ();
 sg13g2_decap_4 FILLER_46_326 ();
 sg13g2_decap_8 FILLER_46_358 ();
 sg13g2_decap_8 FILLER_46_365 ();
 sg13g2_decap_8 FILLER_46_372 ();
 sg13g2_fill_1 FILLER_46_379 ();
 sg13g2_fill_1 FILLER_46_393 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_fill_2 FILLER_46_413 ();
 sg13g2_fill_1 FILLER_46_415 ();
 sg13g2_decap_8 FILLER_46_428 ();
 sg13g2_fill_2 FILLER_46_435 ();
 sg13g2_decap_8 FILLER_46_490 ();
 sg13g2_fill_1 FILLER_46_497 ();
 sg13g2_decap_4 FILLER_46_524 ();
 sg13g2_fill_2 FILLER_46_528 ();
 sg13g2_decap_4 FILLER_46_570 ();
 sg13g2_decap_8 FILLER_46_587 ();
 sg13g2_decap_8 FILLER_46_594 ();
 sg13g2_fill_1 FILLER_46_601 ();
 sg13g2_decap_8 FILLER_46_614 ();
 sg13g2_decap_4 FILLER_46_621 ();
 sg13g2_fill_2 FILLER_46_625 ();
 sg13g2_decap_8 FILLER_46_670 ();
 sg13g2_fill_2 FILLER_46_677 ();
 sg13g2_fill_2 FILLER_46_683 ();
 sg13g2_fill_1 FILLER_46_685 ();
 sg13g2_fill_1 FILLER_46_712 ();
 sg13g2_decap_4 FILLER_46_717 ();
 sg13g2_fill_2 FILLER_46_721 ();
 sg13g2_fill_2 FILLER_46_732 ();
 sg13g2_fill_2 FILLER_46_744 ();
 sg13g2_fill_1 FILLER_46_746 ();
 sg13g2_fill_2 FILLER_46_755 ();
 sg13g2_fill_1 FILLER_46_757 ();
 sg13g2_fill_1 FILLER_46_781 ();
 sg13g2_fill_2 FILLER_46_803 ();
 sg13g2_fill_1 FILLER_46_805 ();
 sg13g2_fill_1 FILLER_46_811 ();
 sg13g2_fill_2 FILLER_46_826 ();
 sg13g2_fill_1 FILLER_46_828 ();
 sg13g2_fill_2 FILLER_46_859 ();
 sg13g2_fill_1 FILLER_46_861 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_4 FILLER_47_7 ();
 sg13g2_fill_1 FILLER_47_11 ();
 sg13g2_fill_2 FILLER_47_16 ();
 sg13g2_fill_1 FILLER_47_18 ();
 sg13g2_fill_2 FILLER_47_91 ();
 sg13g2_fill_2 FILLER_47_133 ();
 sg13g2_fill_1 FILLER_47_135 ();
 sg13g2_decap_8 FILLER_47_144 ();
 sg13g2_fill_1 FILLER_47_151 ();
 sg13g2_decap_4 FILLER_47_156 ();
 sg13g2_fill_1 FILLER_47_160 ();
 sg13g2_fill_1 FILLER_47_166 ();
 sg13g2_decap_8 FILLER_47_181 ();
 sg13g2_fill_2 FILLER_47_188 ();
 sg13g2_decap_8 FILLER_47_197 ();
 sg13g2_decap_8 FILLER_47_204 ();
 sg13g2_fill_2 FILLER_47_211 ();
 sg13g2_fill_1 FILLER_47_213 ();
 sg13g2_fill_2 FILLER_47_218 ();
 sg13g2_fill_2 FILLER_47_246 ();
 sg13g2_fill_1 FILLER_47_278 ();
 sg13g2_fill_1 FILLER_47_285 ();
 sg13g2_decap_8 FILLER_47_312 ();
 sg13g2_decap_8 FILLER_47_319 ();
 sg13g2_fill_2 FILLER_47_326 ();
 sg13g2_decap_8 FILLER_47_347 ();
 sg13g2_decap_8 FILLER_47_354 ();
 sg13g2_fill_1 FILLER_47_404 ();
 sg13g2_decap_4 FILLER_47_417 ();
 sg13g2_decap_8 FILLER_47_457 ();
 sg13g2_fill_2 FILLER_47_464 ();
 sg13g2_fill_1 FILLER_47_466 ();
 sg13g2_decap_4 FILLER_47_471 ();
 sg13g2_fill_1 FILLER_47_475 ();
 sg13g2_fill_2 FILLER_47_488 ();
 sg13g2_fill_1 FILLER_47_525 ();
 sg13g2_fill_1 FILLER_47_559 ();
 sg13g2_decap_8 FILLER_47_595 ();
 sg13g2_fill_1 FILLER_47_602 ();
 sg13g2_decap_4 FILLER_47_613 ();
 sg13g2_fill_1 FILLER_47_617 ();
 sg13g2_decap_8 FILLER_47_622 ();
 sg13g2_decap_8 FILLER_47_629 ();
 sg13g2_decap_4 FILLER_47_636 ();
 sg13g2_decap_8 FILLER_47_670 ();
 sg13g2_fill_1 FILLER_47_682 ();
 sg13g2_fill_1 FILLER_47_691 ();
 sg13g2_decap_4 FILLER_47_719 ();
 sg13g2_fill_1 FILLER_47_723 ();
 sg13g2_fill_2 FILLER_47_754 ();
 sg13g2_decap_4 FILLER_47_761 ();
 sg13g2_fill_2 FILLER_47_795 ();
 sg13g2_fill_1 FILLER_47_832 ();
 sg13g2_fill_2 FILLER_47_859 ();
 sg13g2_fill_1 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_fill_2 FILLER_48_14 ();
 sg13g2_decap_4 FILLER_48_20 ();
 sg13g2_fill_2 FILLER_48_37 ();
 sg13g2_fill_1 FILLER_48_39 ();
 sg13g2_fill_1 FILLER_48_68 ();
 sg13g2_fill_2 FILLER_48_100 ();
 sg13g2_fill_2 FILLER_48_136 ();
 sg13g2_fill_2 FILLER_48_176 ();
 sg13g2_fill_2 FILLER_48_198 ();
 sg13g2_fill_2 FILLER_48_229 ();
 sg13g2_fill_1 FILLER_48_231 ();
 sg13g2_fill_1 FILLER_48_258 ();
 sg13g2_decap_8 FILLER_48_285 ();
 sg13g2_decap_4 FILLER_48_292 ();
 sg13g2_fill_1 FILLER_48_296 ();
 sg13g2_decap_8 FILLER_48_301 ();
 sg13g2_decap_8 FILLER_48_308 ();
 sg13g2_decap_4 FILLER_48_315 ();
 sg13g2_fill_2 FILLER_48_319 ();
 sg13g2_fill_2 FILLER_48_353 ();
 sg13g2_fill_1 FILLER_48_355 ();
 sg13g2_fill_2 FILLER_48_382 ();
 sg13g2_fill_2 FILLER_48_393 ();
 sg13g2_fill_2 FILLER_48_400 ();
 sg13g2_fill_1 FILLER_48_407 ();
 sg13g2_fill_1 FILLER_48_431 ();
 sg13g2_decap_8 FILLER_48_440 ();
 sg13g2_fill_2 FILLER_48_447 ();
 sg13g2_fill_2 FILLER_48_454 ();
 sg13g2_decap_8 FILLER_48_515 ();
 sg13g2_decap_4 FILLER_48_547 ();
 sg13g2_fill_2 FILLER_48_551 ();
 sg13g2_fill_1 FILLER_48_561 ();
 sg13g2_decap_4 FILLER_48_570 ();
 sg13g2_fill_1 FILLER_48_574 ();
 sg13g2_fill_1 FILLER_48_606 ();
 sg13g2_decap_8 FILLER_48_641 ();
 sg13g2_fill_2 FILLER_48_648 ();
 sg13g2_fill_2 FILLER_48_671 ();
 sg13g2_fill_1 FILLER_48_673 ();
 sg13g2_fill_1 FILLER_48_726 ();
 sg13g2_fill_2 FILLER_48_736 ();
 sg13g2_fill_1 FILLER_48_738 ();
 sg13g2_fill_2 FILLER_48_747 ();
 sg13g2_fill_1 FILLER_48_749 ();
 sg13g2_fill_2 FILLER_48_759 ();
 sg13g2_fill_1 FILLER_48_761 ();
 sg13g2_fill_1 FILLER_48_774 ();
 sg13g2_fill_1 FILLER_48_798 ();
 sg13g2_fill_2 FILLER_48_812 ();
 sg13g2_fill_1 FILLER_48_829 ();
 sg13g2_fill_2 FILLER_48_835 ();
 sg13g2_fill_2 FILLER_48_846 ();
 sg13g2_fill_1 FILLER_48_861 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_fill_2 FILLER_49_36 ();
 sg13g2_fill_1 FILLER_49_38 ();
 sg13g2_fill_2 FILLER_49_99 ();
 sg13g2_fill_1 FILLER_49_105 ();
 sg13g2_fill_1 FILLER_49_141 ();
 sg13g2_fill_2 FILLER_49_156 ();
 sg13g2_fill_1 FILLER_49_173 ();
 sg13g2_fill_2 FILLER_49_184 ();
 sg13g2_decap_8 FILLER_49_195 ();
 sg13g2_fill_2 FILLER_49_202 ();
 sg13g2_decap_4 FILLER_49_224 ();
 sg13g2_fill_2 FILLER_49_228 ();
 sg13g2_fill_2 FILLER_49_256 ();
 sg13g2_fill_1 FILLER_49_258 ();
 sg13g2_fill_1 FILLER_49_298 ();
 sg13g2_decap_8 FILLER_49_317 ();
 sg13g2_decap_8 FILLER_49_324 ();
 sg13g2_decap_8 FILLER_49_347 ();
 sg13g2_decap_4 FILLER_49_354 ();
 sg13g2_fill_2 FILLER_49_374 ();
 sg13g2_fill_2 FILLER_49_389 ();
 sg13g2_fill_2 FILLER_49_456 ();
 sg13g2_fill_1 FILLER_49_466 ();
 sg13g2_fill_2 FILLER_49_472 ();
 sg13g2_fill_1 FILLER_49_474 ();
 sg13g2_decap_4 FILLER_49_479 ();
 sg13g2_fill_2 FILLER_49_483 ();
 sg13g2_fill_1 FILLER_49_490 ();
 sg13g2_decap_4 FILLER_49_495 ();
 sg13g2_fill_1 FILLER_49_499 ();
 sg13g2_fill_2 FILLER_49_534 ();
 sg13g2_fill_1 FILLER_49_536 ();
 sg13g2_decap_4 FILLER_49_551 ();
 sg13g2_fill_2 FILLER_49_555 ();
 sg13g2_fill_2 FILLER_49_562 ();
 sg13g2_decap_4 FILLER_49_575 ();
 sg13g2_fill_2 FILLER_49_584 ();
 sg13g2_decap_4 FILLER_49_599 ();
 sg13g2_fill_1 FILLER_49_603 ();
 sg13g2_fill_2 FILLER_49_609 ();
 sg13g2_decap_4 FILLER_49_615 ();
 sg13g2_fill_1 FILLER_49_619 ();
 sg13g2_fill_1 FILLER_49_629 ();
 sg13g2_fill_2 FILLER_49_646 ();
 sg13g2_fill_1 FILLER_49_663 ();
 sg13g2_decap_4 FILLER_49_673 ();
 sg13g2_fill_1 FILLER_49_682 ();
 sg13g2_decap_4 FILLER_49_688 ();
 sg13g2_fill_2 FILLER_49_692 ();
 sg13g2_fill_1 FILLER_49_702 ();
 sg13g2_fill_2 FILLER_49_725 ();
 sg13g2_fill_1 FILLER_49_727 ();
 sg13g2_fill_2 FILLER_49_736 ();
 sg13g2_fill_1 FILLER_49_738 ();
 sg13g2_decap_8 FILLER_49_803 ();
 sg13g2_fill_1 FILLER_49_810 ();
 sg13g2_fill_1 FILLER_49_830 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_fill_2 FILLER_50_14 ();
 sg13g2_fill_1 FILLER_50_16 ();
 sg13g2_fill_1 FILLER_50_84 ();
 sg13g2_fill_1 FILLER_50_89 ();
 sg13g2_fill_2 FILLER_50_133 ();
 sg13g2_fill_2 FILLER_50_262 ();
 sg13g2_fill_1 FILLER_50_264 ();
 sg13g2_decap_4 FILLER_50_287 ();
 sg13g2_fill_2 FILLER_50_291 ();
 sg13g2_fill_1 FILLER_50_323 ();
 sg13g2_fill_1 FILLER_50_401 ();
 sg13g2_decap_8 FILLER_50_410 ();
 sg13g2_fill_2 FILLER_50_417 ();
 sg13g2_fill_2 FILLER_50_423 ();
 sg13g2_fill_1 FILLER_50_425 ();
 sg13g2_fill_2 FILLER_50_430 ();
 sg13g2_decap_8 FILLER_50_436 ();
 sg13g2_fill_2 FILLER_50_448 ();
 sg13g2_fill_1 FILLER_50_458 ();
 sg13g2_decap_4 FILLER_50_494 ();
 sg13g2_decap_4 FILLER_50_506 ();
 sg13g2_fill_1 FILLER_50_510 ();
 sg13g2_fill_2 FILLER_50_519 ();
 sg13g2_fill_1 FILLER_50_548 ();
 sg13g2_fill_2 FILLER_50_590 ();
 sg13g2_fill_1 FILLER_50_592 ();
 sg13g2_decap_4 FILLER_50_628 ();
 sg13g2_fill_1 FILLER_50_632 ();
 sg13g2_fill_2 FILLER_50_667 ();
 sg13g2_fill_1 FILLER_50_695 ();
 sg13g2_decap_4 FILLER_50_727 ();
 sg13g2_fill_2 FILLER_50_731 ();
 sg13g2_fill_2 FILLER_50_742 ();
 sg13g2_fill_1 FILLER_50_744 ();
 sg13g2_fill_2 FILLER_50_759 ();
 sg13g2_fill_1 FILLER_50_761 ();
 sg13g2_fill_2 FILLER_50_783 ();
 sg13g2_fill_2 FILLER_50_808 ();
 sg13g2_fill_1 FILLER_50_810 ();
 sg13g2_fill_1 FILLER_50_820 ();
 sg13g2_fill_2 FILLER_50_860 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_fill_1 FILLER_51_28 ();
 sg13g2_fill_1 FILLER_51_64 ();
 sg13g2_fill_2 FILLER_51_90 ();
 sg13g2_fill_1 FILLER_51_100 ();
 sg13g2_fill_1 FILLER_51_149 ();
 sg13g2_fill_1 FILLER_51_160 ();
 sg13g2_fill_1 FILLER_51_181 ();
 sg13g2_fill_2 FILLER_51_199 ();
 sg13g2_fill_1 FILLER_51_201 ();
 sg13g2_fill_2 FILLER_51_211 ();
 sg13g2_fill_1 FILLER_51_213 ();
 sg13g2_fill_2 FILLER_51_229 ();
 sg13g2_decap_4 FILLER_51_235 ();
 sg13g2_decap_8 FILLER_51_278 ();
 sg13g2_fill_2 FILLER_51_285 ();
 sg13g2_fill_1 FILLER_51_287 ();
 sg13g2_fill_1 FILLER_51_315 ();
 sg13g2_decap_4 FILLER_51_343 ();
 sg13g2_decap_8 FILLER_51_351 ();
 sg13g2_fill_1 FILLER_51_358 ();
 sg13g2_fill_1 FILLER_51_369 ();
 sg13g2_decap_8 FILLER_51_375 ();
 sg13g2_decap_8 FILLER_51_382 ();
 sg13g2_fill_1 FILLER_51_389 ();
 sg13g2_decap_8 FILLER_51_401 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_fill_2 FILLER_51_433 ();
 sg13g2_fill_2 FILLER_51_504 ();
 sg13g2_fill_2 FILLER_51_557 ();
 sg13g2_fill_1 FILLER_51_559 ();
 sg13g2_decap_4 FILLER_51_569 ();
 sg13g2_fill_2 FILLER_51_573 ();
 sg13g2_fill_2 FILLER_51_584 ();
 sg13g2_fill_1 FILLER_51_586 ();
 sg13g2_decap_4 FILLER_51_592 ();
 sg13g2_fill_1 FILLER_51_606 ();
 sg13g2_fill_1 FILLER_51_612 ();
 sg13g2_decap_4 FILLER_51_621 ();
 sg13g2_fill_1 FILLER_51_625 ();
 sg13g2_fill_1 FILLER_51_639 ();
 sg13g2_fill_1 FILLER_51_657 ();
 sg13g2_fill_2 FILLER_51_681 ();
 sg13g2_fill_1 FILLER_51_683 ();
 sg13g2_fill_2 FILLER_51_689 ();
 sg13g2_fill_2 FILLER_51_723 ();
 sg13g2_fill_1 FILLER_51_782 ();
 sg13g2_fill_2 FILLER_51_832 ();
 sg13g2_fill_2 FILLER_51_860 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_7 ();
 sg13g2_fill_1 FILLER_52_9 ();
 sg13g2_fill_2 FILLER_52_19 ();
 sg13g2_fill_1 FILLER_52_21 ();
 sg13g2_fill_1 FILLER_52_55 ();
 sg13g2_fill_1 FILLER_52_66 ();
 sg13g2_fill_1 FILLER_52_92 ();
 sg13g2_fill_1 FILLER_52_151 ();
 sg13g2_fill_1 FILLER_52_188 ();
 sg13g2_fill_1 FILLER_52_201 ();
 sg13g2_fill_1 FILLER_52_235 ();
 sg13g2_decap_8 FILLER_52_262 ();
 sg13g2_decap_4 FILLER_52_269 ();
 sg13g2_fill_2 FILLER_52_273 ();
 sg13g2_fill_1 FILLER_52_280 ();
 sg13g2_fill_1 FILLER_52_326 ();
 sg13g2_fill_2 FILLER_52_337 ();
 sg13g2_fill_1 FILLER_52_339 ();
 sg13g2_fill_2 FILLER_52_345 ();
 sg13g2_decap_8 FILLER_52_352 ();
 sg13g2_fill_1 FILLER_52_359 ();
 sg13g2_decap_8 FILLER_52_365 ();
 sg13g2_decap_8 FILLER_52_372 ();
 sg13g2_fill_1 FILLER_52_379 ();
 sg13g2_decap_4 FILLER_52_428 ();
 sg13g2_fill_2 FILLER_52_432 ();
 sg13g2_fill_2 FILLER_52_439 ();
 sg13g2_decap_8 FILLER_52_461 ();
 sg13g2_decap_8 FILLER_52_468 ();
 sg13g2_decap_8 FILLER_52_475 ();
 sg13g2_fill_1 FILLER_52_482 ();
 sg13g2_decap_8 FILLER_52_492 ();
 sg13g2_fill_1 FILLER_52_499 ();
 sg13g2_fill_2 FILLER_52_509 ();
 sg13g2_fill_2 FILLER_52_515 ();
 sg13g2_decap_4 FILLER_52_521 ();
 sg13g2_fill_1 FILLER_52_525 ();
 sg13g2_fill_2 FILLER_52_530 ();
 sg13g2_fill_1 FILLER_52_532 ();
 sg13g2_decap_4 FILLER_52_573 ();
 sg13g2_decap_4 FILLER_52_643 ();
 sg13g2_fill_2 FILLER_52_657 ();
 sg13g2_fill_1 FILLER_52_659 ();
 sg13g2_fill_1 FILLER_52_674 ();
 sg13g2_fill_1 FILLER_52_683 ();
 sg13g2_fill_2 FILLER_52_723 ();
 sg13g2_fill_1 FILLER_52_725 ();
 sg13g2_fill_2 FILLER_52_731 ();
 sg13g2_decap_4 FILLER_52_742 ();
 sg13g2_fill_2 FILLER_52_746 ();
 sg13g2_fill_2 FILLER_52_761 ();
 sg13g2_fill_1 FILLER_52_763 ();
 sg13g2_fill_1 FILLER_52_785 ();
 sg13g2_decap_8 FILLER_52_812 ();
 sg13g2_fill_1 FILLER_52_819 ();
 sg13g2_fill_2 FILLER_52_829 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_fill_2 FILLER_53_47 ();
 sg13g2_fill_2 FILLER_53_66 ();
 sg13g2_fill_2 FILLER_53_91 ();
 sg13g2_fill_1 FILLER_53_149 ();
 sg13g2_fill_1 FILLER_53_165 ();
 sg13g2_fill_2 FILLER_53_179 ();
 sg13g2_decap_4 FILLER_53_206 ();
 sg13g2_fill_1 FILLER_53_210 ();
 sg13g2_fill_1 FILLER_53_220 ();
 sg13g2_fill_2 FILLER_53_232 ();
 sg13g2_fill_1 FILLER_53_234 ();
 sg13g2_decap_4 FILLER_53_261 ();
 sg13g2_fill_1 FILLER_53_265 ();
 sg13g2_fill_1 FILLER_53_284 ();
 sg13g2_fill_2 FILLER_53_297 ();
 sg13g2_fill_2 FILLER_53_318 ();
 sg13g2_fill_1 FILLER_53_320 ();
 sg13g2_fill_1 FILLER_53_339 ();
 sg13g2_fill_2 FILLER_53_376 ();
 sg13g2_fill_1 FILLER_53_378 ();
 sg13g2_fill_1 FILLER_53_389 ();
 sg13g2_fill_1 FILLER_53_394 ();
 sg13g2_fill_2 FILLER_53_411 ();
 sg13g2_fill_2 FILLER_53_498 ();
 sg13g2_fill_1 FILLER_53_500 ();
 sg13g2_fill_2 FILLER_53_541 ();
 sg13g2_fill_1 FILLER_53_543 ();
 sg13g2_fill_2 FILLER_53_553 ();
 sg13g2_fill_1 FILLER_53_555 ();
 sg13g2_decap_4 FILLER_53_577 ();
 sg13g2_fill_2 FILLER_53_581 ();
 sg13g2_fill_2 FILLER_53_601 ();
 sg13g2_decap_8 FILLER_53_631 ();
 sg13g2_decap_8 FILLER_53_638 ();
 sg13g2_fill_1 FILLER_53_711 ();
 sg13g2_fill_2 FILLER_53_730 ();
 sg13g2_decap_4 FILLER_53_741 ();
 sg13g2_fill_1 FILLER_53_745 ();
 sg13g2_fill_1 FILLER_53_807 ();
 sg13g2_fill_2 FILLER_53_813 ();
 sg13g2_fill_1 FILLER_53_815 ();
 sg13g2_fill_2 FILLER_53_825 ();
 sg13g2_fill_1 FILLER_53_827 ();
 sg13g2_fill_2 FILLER_53_833 ();
 sg13g2_fill_1 FILLER_53_835 ();
 sg13g2_fill_2 FILLER_53_841 ();
 sg13g2_fill_1 FILLER_53_861 ();
 sg13g2_fill_1 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_27 ();
 sg13g2_fill_2 FILLER_54_34 ();
 sg13g2_fill_1 FILLER_54_75 ();
 sg13g2_fill_2 FILLER_54_89 ();
 sg13g2_fill_2 FILLER_54_135 ();
 sg13g2_fill_1 FILLER_54_137 ();
 sg13g2_decap_8 FILLER_54_213 ();
 sg13g2_decap_8 FILLER_54_224 ();
 sg13g2_fill_2 FILLER_54_248 ();
 sg13g2_fill_1 FILLER_54_250 ();
 sg13g2_decap_8 FILLER_54_266 ();
 sg13g2_fill_2 FILLER_54_278 ();
 sg13g2_decap_8 FILLER_54_285 ();
 sg13g2_decap_4 FILLER_54_309 ();
 sg13g2_fill_1 FILLER_54_313 ();
 sg13g2_decap_4 FILLER_54_334 ();
 sg13g2_decap_8 FILLER_54_345 ();
 sg13g2_fill_1 FILLER_54_352 ();
 sg13g2_fill_2 FILLER_54_362 ();
 sg13g2_fill_2 FILLER_54_372 ();
 sg13g2_fill_1 FILLER_54_374 ();
 sg13g2_fill_1 FILLER_54_389 ();
 sg13g2_fill_2 FILLER_54_398 ();
 sg13g2_fill_1 FILLER_54_400 ();
 sg13g2_fill_1 FILLER_54_427 ();
 sg13g2_decap_8 FILLER_54_432 ();
 sg13g2_fill_2 FILLER_54_439 ();
 sg13g2_fill_1 FILLER_54_445 ();
 sg13g2_decap_8 FILLER_54_459 ();
 sg13g2_decap_8 FILLER_54_466 ();
 sg13g2_decap_4 FILLER_54_473 ();
 sg13g2_decap_4 FILLER_54_481 ();
 sg13g2_fill_1 FILLER_54_485 ();
 sg13g2_decap_4 FILLER_54_516 ();
 sg13g2_fill_1 FILLER_54_520 ();
 sg13g2_fill_2 FILLER_54_546 ();
 sg13g2_fill_1 FILLER_54_548 ();
 sg13g2_fill_2 FILLER_54_597 ();
 sg13g2_decap_8 FILLER_54_618 ();
 sg13g2_fill_2 FILLER_54_625 ();
 sg13g2_fill_1 FILLER_54_656 ();
 sg13g2_fill_1 FILLER_54_661 ();
 sg13g2_fill_1 FILLER_54_675 ();
 sg13g2_fill_2 FILLER_54_694 ();
 sg13g2_fill_2 FILLER_54_769 ();
 sg13g2_fill_1 FILLER_54_784 ();
 sg13g2_fill_1 FILLER_54_861 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_4 FILLER_55_14 ();
 sg13g2_fill_1 FILLER_55_18 ();
 sg13g2_fill_1 FILLER_55_55 ();
 sg13g2_fill_2 FILLER_55_168 ();
 sg13g2_fill_1 FILLER_55_179 ();
 sg13g2_fill_1 FILLER_55_232 ();
 sg13g2_decap_8 FILLER_55_298 ();
 sg13g2_fill_1 FILLER_55_305 ();
 sg13g2_decap_8 FILLER_55_310 ();
 sg13g2_decap_4 FILLER_55_317 ();
 sg13g2_fill_1 FILLER_55_321 ();
 sg13g2_fill_2 FILLER_55_327 ();
 sg13g2_decap_8 FILLER_55_367 ();
 sg13g2_decap_4 FILLER_55_374 ();
 sg13g2_fill_1 FILLER_55_378 ();
 sg13g2_decap_4 FILLER_55_395 ();
 sg13g2_fill_1 FILLER_55_399 ();
 sg13g2_decap_8 FILLER_55_404 ();
 sg13g2_fill_1 FILLER_55_411 ();
 sg13g2_decap_8 FILLER_55_416 ();
 sg13g2_decap_8 FILLER_55_423 ();
 sg13g2_fill_2 FILLER_55_430 ();
 sg13g2_fill_1 FILLER_55_432 ();
 sg13g2_fill_1 FILLER_55_448 ();
 sg13g2_fill_1 FILLER_55_454 ();
 sg13g2_fill_1 FILLER_55_481 ();
 sg13g2_fill_2 FILLER_55_487 ();
 sg13g2_fill_1 FILLER_55_503 ();
 sg13g2_fill_2 FILLER_55_565 ();
 sg13g2_fill_2 FILLER_55_581 ();
 sg13g2_fill_1 FILLER_55_583 ();
 sg13g2_fill_1 FILLER_55_627 ();
 sg13g2_fill_2 FILLER_55_658 ();
 sg13g2_fill_1 FILLER_55_660 ();
 sg13g2_fill_2 FILLER_55_666 ();
 sg13g2_fill_1 FILLER_55_668 ();
 sg13g2_fill_1 FILLER_55_682 ();
 sg13g2_fill_1 FILLER_55_722 ();
 sg13g2_fill_1 FILLER_55_727 ();
 sg13g2_decap_4 FILLER_55_732 ();
 sg13g2_fill_2 FILLER_55_749 ();
 sg13g2_fill_1 FILLER_55_768 ();
 sg13g2_fill_2 FILLER_55_783 ();
 sg13g2_fill_1 FILLER_55_785 ();
 sg13g2_decap_4 FILLER_55_811 ();
 sg13g2_fill_1 FILLER_55_819 ();
 sg13g2_fill_2 FILLER_55_824 ();
 sg13g2_fill_1 FILLER_55_826 ();
 sg13g2_fill_1 FILLER_55_861 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_4 FILLER_56_7 ();
 sg13g2_fill_1 FILLER_56_11 ();
 sg13g2_decap_8 FILLER_56_16 ();
 sg13g2_decap_8 FILLER_56_23 ();
 sg13g2_decap_8 FILLER_56_34 ();
 sg13g2_fill_1 FILLER_56_41 ();
 sg13g2_fill_2 FILLER_56_62 ();
 sg13g2_fill_2 FILLER_56_74 ();
 sg13g2_fill_1 FILLER_56_86 ();
 sg13g2_fill_2 FILLER_56_113 ();
 sg13g2_fill_2 FILLER_56_124 ();
 sg13g2_fill_1 FILLER_56_126 ();
 sg13g2_fill_2 FILLER_56_153 ();
 sg13g2_fill_1 FILLER_56_155 ();
 sg13g2_fill_2 FILLER_56_182 ();
 sg13g2_fill_1 FILLER_56_184 ();
 sg13g2_decap_8 FILLER_56_188 ();
 sg13g2_decap_8 FILLER_56_195 ();
 sg13g2_decap_4 FILLER_56_202 ();
 sg13g2_fill_2 FILLER_56_206 ();
 sg13g2_decap_4 FILLER_56_213 ();
 sg13g2_decap_8 FILLER_56_221 ();
 sg13g2_fill_2 FILLER_56_228 ();
 sg13g2_fill_2 FILLER_56_245 ();
 sg13g2_fill_2 FILLER_56_255 ();
 sg13g2_fill_2 FILLER_56_270 ();
 sg13g2_fill_2 FILLER_56_333 ();
 sg13g2_fill_1 FILLER_56_335 ();
 sg13g2_decap_8 FILLER_56_345 ();
 sg13g2_decap_4 FILLER_56_356 ();
 sg13g2_fill_1 FILLER_56_415 ();
 sg13g2_decap_4 FILLER_56_425 ();
 sg13g2_decap_8 FILLER_56_433 ();
 sg13g2_decap_8 FILLER_56_440 ();
 sg13g2_fill_2 FILLER_56_447 ();
 sg13g2_decap_4 FILLER_56_462 ();
 sg13g2_fill_1 FILLER_56_470 ();
 sg13g2_fill_1 FILLER_56_474 ();
 sg13g2_fill_1 FILLER_56_505 ();
 sg13g2_decap_8 FILLER_56_535 ();
 sg13g2_decap_4 FILLER_56_555 ();
 sg13g2_fill_2 FILLER_56_559 ();
 sg13g2_fill_2 FILLER_56_626 ();
 sg13g2_fill_1 FILLER_56_628 ();
 sg13g2_fill_1 FILLER_56_643 ();
 sg13g2_fill_2 FILLER_56_653 ();
 sg13g2_fill_1 FILLER_56_655 ();
 sg13g2_fill_1 FILLER_56_665 ();
 sg13g2_fill_1 FILLER_56_702 ();
 sg13g2_fill_2 FILLER_56_707 ();
 sg13g2_decap_4 FILLER_56_718 ();
 sg13g2_fill_2 FILLER_56_722 ();
 sg13g2_decap_8 FILLER_56_762 ();
 sg13g2_fill_2 FILLER_56_808 ();
 sg13g2_fill_1 FILLER_56_810 ();
 sg13g2_fill_2 FILLER_56_821 ();
 sg13g2_fill_2 FILLER_56_828 ();
 sg13g2_fill_1 FILLER_56_835 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_fill_2 FILLER_57_42 ();
 sg13g2_fill_2 FILLER_57_70 ();
 sg13g2_decap_4 FILLER_57_89 ();
 sg13g2_fill_2 FILLER_57_145 ();
 sg13g2_fill_1 FILLER_57_147 ();
 sg13g2_fill_2 FILLER_57_157 ();
 sg13g2_decap_4 FILLER_57_175 ();
 sg13g2_fill_1 FILLER_57_179 ();
 sg13g2_fill_1 FILLER_57_293 ();
 sg13g2_fill_2 FILLER_57_303 ();
 sg13g2_decap_4 FILLER_57_370 ();
 sg13g2_fill_1 FILLER_57_374 ();
 sg13g2_decap_8 FILLER_57_379 ();
 sg13g2_decap_8 FILLER_57_386 ();
 sg13g2_fill_1 FILLER_57_393 ();
 sg13g2_decap_4 FILLER_57_444 ();
 sg13g2_fill_1 FILLER_57_448 ();
 sg13g2_decap_8 FILLER_57_472 ();
 sg13g2_decap_8 FILLER_57_479 ();
 sg13g2_fill_1 FILLER_57_490 ();
 sg13g2_fill_2 FILLER_57_531 ();
 sg13g2_decap_4 FILLER_57_568 ();
 sg13g2_fill_2 FILLER_57_576 ();
 sg13g2_fill_1 FILLER_57_578 ();
 sg13g2_decap_4 FILLER_57_587 ();
 sg13g2_fill_1 FILLER_57_591 ();
 sg13g2_fill_1 FILLER_57_623 ();
 sg13g2_fill_1 FILLER_57_650 ();
 sg13g2_decap_4 FILLER_57_683 ();
 sg13g2_fill_2 FILLER_57_687 ();
 sg13g2_fill_2 FILLER_57_720 ();
 sg13g2_fill_2 FILLER_57_732 ();
 sg13g2_fill_1 FILLER_57_734 ();
 sg13g2_decap_4 FILLER_57_739 ();
 sg13g2_decap_8 FILLER_57_791 ();
 sg13g2_fill_1 FILLER_57_798 ();
 sg13g2_fill_2 FILLER_57_859 ();
 sg13g2_fill_1 FILLER_57_861 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_4 FILLER_58_35 ();
 sg13g2_fill_1 FILLER_58_39 ();
 sg13g2_decap_4 FILLER_58_50 ();
 sg13g2_fill_1 FILLER_58_54 ();
 sg13g2_fill_1 FILLER_58_59 ();
 sg13g2_fill_2 FILLER_58_64 ();
 sg13g2_fill_1 FILLER_58_92 ();
 sg13g2_fill_2 FILLER_58_102 ();
 sg13g2_fill_1 FILLER_58_104 ();
 sg13g2_fill_1 FILLER_58_118 ();
 sg13g2_fill_1 FILLER_58_132 ();
 sg13g2_fill_2 FILLER_58_194 ();
 sg13g2_decap_4 FILLER_58_207 ();
 sg13g2_fill_2 FILLER_58_211 ();
 sg13g2_fill_1 FILLER_58_225 ();
 sg13g2_fill_1 FILLER_58_235 ();
 sg13g2_fill_2 FILLER_58_242 ();
 sg13g2_fill_2 FILLER_58_253 ();
 sg13g2_fill_2 FILLER_58_275 ();
 sg13g2_fill_1 FILLER_58_277 ();
 sg13g2_fill_1 FILLER_58_292 ();
 sg13g2_decap_4 FILLER_58_392 ();
 sg13g2_decap_4 FILLER_58_431 ();
 sg13g2_fill_2 FILLER_58_435 ();
 sg13g2_fill_1 FILLER_58_442 ();
 sg13g2_decap_4 FILLER_58_446 ();
 sg13g2_fill_1 FILLER_58_492 ();
 sg13g2_fill_2 FILLER_58_510 ();
 sg13g2_fill_1 FILLER_58_512 ();
 sg13g2_fill_2 FILLER_58_522 ();
 sg13g2_fill_1 FILLER_58_524 ();
 sg13g2_fill_2 FILLER_58_539 ();
 sg13g2_fill_1 FILLER_58_541 ();
 sg13g2_fill_2 FILLER_58_572 ();
 sg13g2_decap_8 FILLER_58_578 ();
 sg13g2_decap_4 FILLER_58_593 ();
 sg13g2_fill_1 FILLER_58_597 ();
 sg13g2_decap_8 FILLER_58_602 ();
 sg13g2_decap_8 FILLER_58_609 ();
 sg13g2_fill_1 FILLER_58_616 ();
 sg13g2_fill_2 FILLER_58_627 ();
 sg13g2_fill_2 FILLER_58_634 ();
 sg13g2_fill_1 FILLER_58_679 ();
 sg13g2_decap_4 FILLER_58_692 ();
 sg13g2_fill_2 FILLER_58_709 ();
 sg13g2_decap_4 FILLER_58_742 ();
 sg13g2_fill_2 FILLER_58_746 ();
 sg13g2_fill_2 FILLER_58_757 ();
 sg13g2_fill_2 FILLER_58_763 ();
 sg13g2_fill_1 FILLER_58_810 ();
 sg13g2_fill_1 FILLER_58_824 ();
 sg13g2_fill_2 FILLER_58_860 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_4 FILLER_59_21 ();
 sg13g2_fill_2 FILLER_59_25 ();
 sg13g2_fill_1 FILLER_59_61 ();
 sg13g2_fill_1 FILLER_59_70 ();
 sg13g2_fill_1 FILLER_59_92 ();
 sg13g2_decap_8 FILLER_59_149 ();
 sg13g2_decap_8 FILLER_59_156 ();
 sg13g2_decap_8 FILLER_59_163 ();
 sg13g2_fill_1 FILLER_59_220 ();
 sg13g2_fill_2 FILLER_59_251 ();
 sg13g2_fill_1 FILLER_59_253 ();
 sg13g2_fill_2 FILLER_59_264 ();
 sg13g2_fill_1 FILLER_59_266 ();
 sg13g2_fill_2 FILLER_59_280 ();
 sg13g2_fill_1 FILLER_59_282 ();
 sg13g2_fill_1 FILLER_59_289 ();
 sg13g2_fill_1 FILLER_59_295 ();
 sg13g2_fill_1 FILLER_59_357 ();
 sg13g2_decap_4 FILLER_59_371 ();
 sg13g2_fill_2 FILLER_59_375 ();
 sg13g2_fill_2 FILLER_59_381 ();
 sg13g2_fill_2 FILLER_59_438 ();
 sg13g2_fill_1 FILLER_59_440 ();
 sg13g2_decap_8 FILLER_59_461 ();
 sg13g2_decap_8 FILLER_59_468 ();
 sg13g2_decap_4 FILLER_59_475 ();
 sg13g2_fill_2 FILLER_59_479 ();
 sg13g2_fill_1 FILLER_59_507 ();
 sg13g2_fill_2 FILLER_59_560 ();
 sg13g2_fill_1 FILLER_59_562 ();
 sg13g2_fill_2 FILLER_59_645 ();
 sg13g2_fill_1 FILLER_59_647 ();
 sg13g2_fill_2 FILLER_59_700 ();
 sg13g2_fill_2 FILLER_59_711 ();
 sg13g2_fill_1 FILLER_59_722 ();
 sg13g2_fill_1 FILLER_59_767 ();
 sg13g2_fill_2 FILLER_59_819 ();
 sg13g2_fill_1 FILLER_59_821 ();
 sg13g2_fill_2 FILLER_59_835 ();
 sg13g2_fill_1 FILLER_59_837 ();
 sg13g2_fill_1 FILLER_59_861 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_7 ();
 sg13g2_fill_1 FILLER_60_35 ();
 sg13g2_fill_2 FILLER_60_68 ();
 sg13g2_decap_8 FILLER_60_148 ();
 sg13g2_fill_2 FILLER_60_159 ();
 sg13g2_fill_2 FILLER_60_187 ();
 sg13g2_fill_1 FILLER_60_207 ();
 sg13g2_fill_2 FILLER_60_237 ();
 sg13g2_fill_1 FILLER_60_239 ();
 sg13g2_fill_2 FILLER_60_250 ();
 sg13g2_fill_1 FILLER_60_252 ();
 sg13g2_fill_1 FILLER_60_297 ();
 sg13g2_fill_1 FILLER_60_308 ();
 sg13g2_fill_2 FILLER_60_339 ();
 sg13g2_decap_8 FILLER_60_376 ();
 sg13g2_decap_4 FILLER_60_388 ();
 sg13g2_fill_2 FILLER_60_392 ();
 sg13g2_decap_8 FILLER_60_398 ();
 sg13g2_fill_2 FILLER_60_405 ();
 sg13g2_fill_2 FILLER_60_429 ();
 sg13g2_decap_4 FILLER_60_434 ();
 sg13g2_fill_2 FILLER_60_448 ();
 sg13g2_decap_8 FILLER_60_460 ();
 sg13g2_fill_2 FILLER_60_467 ();
 sg13g2_decap_8 FILLER_60_482 ();
 sg13g2_fill_2 FILLER_60_489 ();
 sg13g2_fill_2 FILLER_60_500 ();
 sg13g2_fill_2 FILLER_60_528 ();
 sg13g2_fill_1 FILLER_60_530 ();
 sg13g2_fill_2 FILLER_60_545 ();
 sg13g2_fill_1 FILLER_60_547 ();
 sg13g2_decap_4 FILLER_60_592 ();
 sg13g2_fill_2 FILLER_60_649 ();
 sg13g2_fill_1 FILLER_60_651 ();
 sg13g2_fill_1 FILLER_60_666 ();
 sg13g2_decap_4 FILLER_60_742 ();
 sg13g2_fill_1 FILLER_60_746 ();
 sg13g2_fill_2 FILLER_60_761 ();
 sg13g2_decap_4 FILLER_60_776 ();
 sg13g2_fill_1 FILLER_60_785 ();
 sg13g2_fill_1 FILLER_60_795 ();
 sg13g2_fill_2 FILLER_60_810 ();
 sg13g2_fill_1 FILLER_60_812 ();
 sg13g2_fill_2 FILLER_60_834 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_58 ();
 sg13g2_fill_1 FILLER_61_60 ();
 sg13g2_fill_1 FILLER_61_89 ();
 sg13g2_fill_2 FILLER_61_112 ();
 sg13g2_fill_2 FILLER_61_123 ();
 sg13g2_fill_1 FILLER_61_125 ();
 sg13g2_fill_1 FILLER_61_232 ();
 sg13g2_fill_2 FILLER_61_255 ();
 sg13g2_fill_2 FILLER_61_276 ();
 sg13g2_fill_1 FILLER_61_278 ();
 sg13g2_fill_2 FILLER_61_287 ();
 sg13g2_fill_1 FILLER_61_297 ();
 sg13g2_fill_1 FILLER_61_321 ();
 sg13g2_fill_2 FILLER_61_362 ();
 sg13g2_decap_8 FILLER_61_368 ();
 sg13g2_fill_2 FILLER_61_432 ();
 sg13g2_fill_2 FILLER_61_437 ();
 sg13g2_decap_8 FILLER_61_459 ();
 sg13g2_fill_2 FILLER_61_466 ();
 sg13g2_decap_4 FILLER_61_484 ();
 sg13g2_fill_1 FILLER_61_488 ();
 sg13g2_fill_1 FILLER_61_515 ();
 sg13g2_fill_2 FILLER_61_565 ();
 sg13g2_decap_4 FILLER_61_601 ();
 sg13g2_fill_2 FILLER_61_605 ();
 sg13g2_fill_1 FILLER_61_615 ();
 sg13g2_fill_2 FILLER_61_647 ();
 sg13g2_decap_4 FILLER_61_697 ();
 sg13g2_fill_2 FILLER_61_723 ();
 sg13g2_fill_1 FILLER_61_725 ();
 sg13g2_fill_1 FILLER_61_773 ();
 sg13g2_fill_2 FILLER_61_778 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_80 ();
 sg13g2_fill_1 FILLER_62_139 ();
 sg13g2_fill_2 FILLER_62_149 ();
 sg13g2_fill_1 FILLER_62_151 ();
 sg13g2_fill_2 FILLER_62_204 ();
 sg13g2_fill_1 FILLER_62_232 ();
 sg13g2_fill_2 FILLER_62_263 ();
 sg13g2_fill_1 FILLER_62_265 ();
 sg13g2_fill_2 FILLER_62_271 ();
 sg13g2_fill_1 FILLER_62_273 ();
 sg13g2_fill_1 FILLER_62_304 ();
 sg13g2_fill_2 FILLER_62_319 ();
 sg13g2_fill_1 FILLER_62_379 ();
 sg13g2_fill_2 FILLER_62_406 ();
 sg13g2_fill_1 FILLER_62_436 ();
 sg13g2_decap_8 FILLER_62_476 ();
 sg13g2_fill_2 FILLER_62_483 ();
 sg13g2_fill_1 FILLER_62_485 ();
 sg13g2_decap_4 FILLER_62_490 ();
 sg13g2_fill_1 FILLER_62_499 ();
 sg13g2_decap_8 FILLER_62_504 ();
 sg13g2_fill_2 FILLER_62_511 ();
 sg13g2_fill_1 FILLER_62_513 ();
 sg13g2_fill_2 FILLER_62_535 ();
 sg13g2_fill_1 FILLER_62_537 ();
 sg13g2_fill_1 FILLER_62_622 ();
 sg13g2_fill_1 FILLER_62_628 ();
 sg13g2_fill_1 FILLER_62_659 ();
 sg13g2_fill_2 FILLER_62_669 ();
 sg13g2_fill_1 FILLER_62_671 ();
 sg13g2_fill_2 FILLER_62_684 ();
 sg13g2_fill_1 FILLER_62_686 ();
 sg13g2_fill_2 FILLER_62_709 ();
 sg13g2_decap_4 FILLER_62_721 ();
 sg13g2_fill_1 FILLER_62_725 ();
 sg13g2_fill_1 FILLER_62_744 ();
 sg13g2_fill_2 FILLER_62_754 ();
 sg13g2_fill_1 FILLER_62_756 ();
 sg13g2_decap_4 FILLER_62_801 ();
 sg13g2_fill_1 FILLER_62_805 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_fill_1 FILLER_63_70 ();
 sg13g2_fill_1 FILLER_63_89 ();
 sg13g2_fill_1 FILLER_63_117 ();
 sg13g2_fill_1 FILLER_63_179 ();
 sg13g2_fill_2 FILLER_63_186 ();
 sg13g2_fill_1 FILLER_63_188 ();
 sg13g2_fill_2 FILLER_63_195 ();
 sg13g2_fill_1 FILLER_63_207 ();
 sg13g2_fill_1 FILLER_63_275 ();
 sg13g2_decap_4 FILLER_63_311 ();
 sg13g2_decap_4 FILLER_63_320 ();
 sg13g2_fill_1 FILLER_63_324 ();
 sg13g2_decap_8 FILLER_63_333 ();
 sg13g2_fill_1 FILLER_63_340 ();
 sg13g2_decap_8 FILLER_63_354 ();
 sg13g2_decap_8 FILLER_63_361 ();
 sg13g2_decap_4 FILLER_63_368 ();
 sg13g2_fill_1 FILLER_63_372 ();
 sg13g2_fill_2 FILLER_63_404 ();
 sg13g2_fill_2 FILLER_63_454 ();
 sg13g2_fill_1 FILLER_63_460 ();
 sg13g2_decap_8 FILLER_63_465 ();
 sg13g2_fill_2 FILLER_63_472 ();
 sg13g2_fill_1 FILLER_63_474 ();
 sg13g2_fill_2 FILLER_63_531 ();
 sg13g2_fill_1 FILLER_63_533 ();
 sg13g2_fill_1 FILLER_63_555 ();
 sg13g2_fill_2 FILLER_63_561 ();
 sg13g2_fill_1 FILLER_63_563 ();
 sg13g2_fill_2 FILLER_63_604 ();
 sg13g2_fill_1 FILLER_63_606 ();
 sg13g2_fill_2 FILLER_63_633 ();
 sg13g2_fill_1 FILLER_63_684 ();
 sg13g2_decap_8 FILLER_63_715 ();
 sg13g2_decap_4 FILLER_63_722 ();
 sg13g2_fill_2 FILLER_63_726 ();
 sg13g2_fill_2 FILLER_63_763 ();
 sg13g2_fill_2 FILLER_63_774 ();
 sg13g2_fill_1 FILLER_63_776 ();
 sg13g2_fill_2 FILLER_63_782 ();
 sg13g2_fill_1 FILLER_63_784 ();
 sg13g2_fill_1 FILLER_63_824 ();
 sg13g2_fill_1 FILLER_63_848 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_39 ();
 sg13g2_fill_2 FILLER_64_111 ();
 sg13g2_fill_1 FILLER_64_113 ();
 sg13g2_fill_1 FILLER_64_128 ();
 sg13g2_fill_1 FILLER_64_133 ();
 sg13g2_fill_2 FILLER_64_160 ();
 sg13g2_fill_2 FILLER_64_191 ();
 sg13g2_fill_1 FILLER_64_219 ();
 sg13g2_fill_1 FILLER_64_227 ();
 sg13g2_fill_2 FILLER_64_255 ();
 sg13g2_fill_2 FILLER_64_315 ();
 sg13g2_fill_1 FILLER_64_317 ();
 sg13g2_fill_2 FILLER_64_333 ();
 sg13g2_fill_1 FILLER_64_335 ();
 sg13g2_fill_2 FILLER_64_366 ();
 sg13g2_fill_1 FILLER_64_415 ();
 sg13g2_decap_8 FILLER_64_480 ();
 sg13g2_decap_4 FILLER_64_487 ();
 sg13g2_fill_1 FILLER_64_500 ();
 sg13g2_fill_1 FILLER_64_515 ();
 sg13g2_fill_2 FILLER_64_525 ();
 sg13g2_fill_2 FILLER_64_540 ();
 sg13g2_fill_1 FILLER_64_542 ();
 sg13g2_fill_2 FILLER_64_577 ();
 sg13g2_fill_1 FILLER_64_579 ();
 sg13g2_fill_1 FILLER_64_610 ();
 sg13g2_fill_2 FILLER_64_682 ();
 sg13g2_fill_1 FILLER_64_706 ();
 sg13g2_fill_1 FILLER_64_733 ();
 sg13g2_fill_2 FILLER_64_774 ();
 sg13g2_fill_2 FILLER_64_811 ();
 sg13g2_fill_1 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_49 ();
 sg13g2_fill_2 FILLER_65_80 ();
 sg13g2_fill_1 FILLER_65_82 ();
 sg13g2_fill_2 FILLER_65_88 ();
 sg13g2_fill_2 FILLER_65_137 ();
 sg13g2_decap_8 FILLER_65_169 ();
 sg13g2_fill_2 FILLER_65_176 ();
 sg13g2_fill_1 FILLER_65_178 ();
 sg13g2_fill_1 FILLER_65_184 ();
 sg13g2_fill_2 FILLER_65_194 ();
 sg13g2_fill_2 FILLER_65_210 ();
 sg13g2_fill_1 FILLER_65_212 ();
 sg13g2_fill_1 FILLER_65_221 ();
 sg13g2_fill_2 FILLER_65_240 ();
 sg13g2_fill_2 FILLER_65_248 ();
 sg13g2_fill_1 FILLER_65_281 ();
 sg13g2_decap_8 FILLER_65_308 ();
 sg13g2_fill_2 FILLER_65_336 ();
 sg13g2_decap_4 FILLER_65_373 ();
 sg13g2_fill_1 FILLER_65_377 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_fill_2 FILLER_65_423 ();
 sg13g2_fill_2 FILLER_65_439 ();
 sg13g2_fill_2 FILLER_65_450 ();
 sg13g2_fill_1 FILLER_65_452 ();
 sg13g2_fill_2 FILLER_65_545 ();
 sg13g2_fill_1 FILLER_65_547 ();
 sg13g2_fill_2 FILLER_65_579 ();
 sg13g2_fill_1 FILLER_65_595 ();
 sg13g2_decap_4 FILLER_65_631 ();
 sg13g2_fill_2 FILLER_65_635 ();
 sg13g2_fill_1 FILLER_65_651 ();
 sg13g2_fill_2 FILLER_65_678 ();
 sg13g2_fill_2 FILLER_65_745 ();
 sg13g2_fill_1 FILLER_65_747 ();
 sg13g2_fill_2 FILLER_65_791 ();
 sg13g2_fill_1 FILLER_65_817 ();
 sg13g2_fill_1 FILLER_65_844 ();
 sg13g2_decap_4 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_4 ();
 sg13g2_fill_1 FILLER_66_48 ();
 sg13g2_fill_1 FILLER_66_94 ();
 sg13g2_fill_1 FILLER_66_99 ();
 sg13g2_fill_1 FILLER_66_128 ();
 sg13g2_fill_1 FILLER_66_141 ();
 sg13g2_fill_2 FILLER_66_148 ();
 sg13g2_fill_2 FILLER_66_163 ();
 sg13g2_fill_2 FILLER_66_214 ();
 sg13g2_fill_2 FILLER_66_234 ();
 sg13g2_fill_1 FILLER_66_236 ();
 sg13g2_fill_2 FILLER_66_259 ();
 sg13g2_fill_1 FILLER_66_261 ();
 sg13g2_decap_4 FILLER_66_272 ();
 sg13g2_fill_1 FILLER_66_276 ();
 sg13g2_decap_4 FILLER_66_300 ();
 sg13g2_fill_2 FILLER_66_304 ();
 sg13g2_fill_2 FILLER_66_338 ();
 sg13g2_fill_1 FILLER_66_340 ();
 sg13g2_decap_4 FILLER_66_366 ();
 sg13g2_fill_1 FILLER_66_370 ();
 sg13g2_fill_1 FILLER_66_481 ();
 sg13g2_decap_4 FILLER_66_486 ();
 sg13g2_fill_1 FILLER_66_490 ();
 sg13g2_fill_1 FILLER_66_500 ();
 sg13g2_fill_1 FILLER_66_514 ();
 sg13g2_fill_2 FILLER_66_554 ();
 sg13g2_fill_1 FILLER_66_556 ();
 sg13g2_fill_2 FILLER_66_592 ();
 sg13g2_fill_2 FILLER_66_619 ();
 sg13g2_decap_4 FILLER_66_630 ();
 sg13g2_fill_2 FILLER_66_647 ();
 sg13g2_fill_1 FILLER_66_649 ();
 sg13g2_decap_8 FILLER_66_668 ();
 sg13g2_decap_8 FILLER_66_675 ();
 sg13g2_decap_4 FILLER_66_682 ();
 sg13g2_fill_2 FILLER_66_686 ();
 sg13g2_fill_2 FILLER_66_817 ();
 sg13g2_fill_1 FILLER_66_831 ();
 sg13g2_fill_2 FILLER_66_837 ();
 sg13g2_fill_1 FILLER_66_839 ();
 sg13g2_decap_4 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_4 ();
 sg13g2_fill_1 FILLER_67_36 ();
 sg13g2_fill_1 FILLER_67_154 ();
 sg13g2_fill_1 FILLER_67_159 ();
 sg13g2_decap_8 FILLER_67_165 ();
 sg13g2_fill_2 FILLER_67_192 ();
 sg13g2_decap_4 FILLER_67_198 ();
 sg13g2_fill_1 FILLER_67_202 ();
 sg13g2_fill_1 FILLER_67_231 ();
 sg13g2_fill_2 FILLER_67_254 ();
 sg13g2_fill_1 FILLER_67_256 ();
 sg13g2_fill_2 FILLER_67_280 ();
 sg13g2_decap_8 FILLER_67_287 ();
 sg13g2_decap_4 FILLER_67_294 ();
 sg13g2_fill_1 FILLER_67_298 ();
 sg13g2_fill_1 FILLER_67_342 ();
 sg13g2_decap_4 FILLER_67_369 ();
 sg13g2_fill_1 FILLER_67_399 ();
 sg13g2_fill_2 FILLER_67_446 ();
 sg13g2_decap_4 FILLER_67_529 ();
 sg13g2_fill_2 FILLER_67_538 ();
 sg13g2_fill_1 FILLER_67_540 ();
 sg13g2_fill_1 FILLER_67_550 ();
 sg13g2_fill_2 FILLER_67_563 ();
 sg13g2_fill_1 FILLER_67_578 ();
 sg13g2_decap_4 FILLER_67_627 ();
 sg13g2_fill_2 FILLER_67_631 ();
 sg13g2_fill_1 FILLER_67_763 ();
 sg13g2_fill_1 FILLER_67_794 ();
 sg13g2_fill_2 FILLER_67_800 ();
 sg13g2_fill_2 FILLER_67_810 ();
 sg13g2_fill_1 FILLER_67_812 ();
 sg13g2_fill_2 FILLER_67_834 ();
 sg13g2_decap_4 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_35 ();
 sg13g2_fill_1 FILLER_68_45 ();
 sg13g2_fill_1 FILLER_68_77 ();
 sg13g2_decap_4 FILLER_68_121 ();
 sg13g2_fill_2 FILLER_68_142 ();
 sg13g2_decap_4 FILLER_68_170 ();
 sg13g2_fill_2 FILLER_68_200 ();
 sg13g2_fill_1 FILLER_68_202 ();
 sg13g2_decap_8 FILLER_68_209 ();
 sg13g2_decap_4 FILLER_68_216 ();
 sg13g2_fill_1 FILLER_68_220 ();
 sg13g2_decap_4 FILLER_68_226 ();
 sg13g2_fill_2 FILLER_68_230 ();
 sg13g2_fill_1 FILLER_68_242 ();
 sg13g2_fill_2 FILLER_68_252 ();
 sg13g2_fill_1 FILLER_68_254 ();
 sg13g2_fill_1 FILLER_68_293 ();
 sg13g2_fill_1 FILLER_68_339 ();
 sg13g2_fill_1 FILLER_68_344 ();
 sg13g2_fill_2 FILLER_68_351 ();
 sg13g2_fill_1 FILLER_68_353 ();
 sg13g2_decap_4 FILLER_68_363 ();
 sg13g2_fill_2 FILLER_68_367 ();
 sg13g2_fill_1 FILLER_68_457 ();
 sg13g2_decap_8 FILLER_68_485 ();
 sg13g2_decap_4 FILLER_68_501 ();
 sg13g2_fill_2 FILLER_68_505 ();
 sg13g2_decap_4 FILLER_68_521 ();
 sg13g2_fill_1 FILLER_68_567 ();
 sg13g2_decap_8 FILLER_68_594 ();
 sg13g2_decap_4 FILLER_68_601 ();
 sg13g2_decap_8 FILLER_68_640 ();
 sg13g2_fill_2 FILLER_68_669 ();
 sg13g2_decap_4 FILLER_68_684 ();
 sg13g2_fill_2 FILLER_68_723 ();
 sg13g2_fill_1 FILLER_68_748 ();
 sg13g2_fill_2 FILLER_68_770 ();
 sg13g2_fill_1 FILLER_68_791 ();
 sg13g2_fill_1 FILLER_68_832 ();
 sg13g2_fill_2 FILLER_68_859 ();
 sg13g2_fill_1 FILLER_68_861 ();
 sg13g2_fill_2 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_28 ();
 sg13g2_decap_4 FILLER_69_92 ();
 sg13g2_decap_4 FILLER_69_100 ();
 sg13g2_fill_2 FILLER_69_104 ();
 sg13g2_decap_8 FILLER_69_110 ();
 sg13g2_fill_1 FILLER_69_117 ();
 sg13g2_fill_2 FILLER_69_131 ();
 sg13g2_fill_1 FILLER_69_133 ();
 sg13g2_fill_2 FILLER_69_157 ();
 sg13g2_fill_1 FILLER_69_159 ();
 sg13g2_fill_1 FILLER_69_181 ();
 sg13g2_fill_2 FILLER_69_192 ();
 sg13g2_fill_1 FILLER_69_194 ();
 sg13g2_fill_2 FILLER_69_244 ();
 sg13g2_fill_2 FILLER_69_251 ();
 sg13g2_decap_4 FILLER_69_265 ();
 sg13g2_fill_1 FILLER_69_269 ();
 sg13g2_fill_1 FILLER_69_287 ();
 sg13g2_decap_8 FILLER_69_293 ();
 sg13g2_fill_2 FILLER_69_300 ();
 sg13g2_fill_2 FILLER_69_307 ();
 sg13g2_fill_2 FILLER_69_324 ();
 sg13g2_fill_1 FILLER_69_347 ();
 sg13g2_fill_1 FILLER_69_374 ();
 sg13g2_fill_2 FILLER_69_410 ();
 sg13g2_fill_2 FILLER_69_446 ();
 sg13g2_fill_1 FILLER_69_448 ();
 sg13g2_fill_1 FILLER_69_479 ();
 sg13g2_fill_1 FILLER_69_511 ();
 sg13g2_decap_4 FILLER_69_533 ();
 sg13g2_decap_8 FILLER_69_581 ();
 sg13g2_decap_4 FILLER_69_588 ();
 sg13g2_decap_4 FILLER_69_622 ();
 sg13g2_decap_4 FILLER_69_709 ();
 sg13g2_fill_2 FILLER_69_769 ();
 sg13g2_fill_1 FILLER_69_771 ();
 sg13g2_decap_4 FILLER_69_798 ();
 sg13g2_fill_1 FILLER_69_806 ();
 sg13g2_fill_2 FILLER_69_842 ();
 sg13g2_decap_4 FILLER_69_856 ();
 sg13g2_fill_2 FILLER_69_860 ();
 sg13g2_decap_4 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_4 ();
 sg13g2_fill_2 FILLER_70_41 ();
 sg13g2_fill_2 FILLER_70_52 ();
 sg13g2_decap_8 FILLER_70_86 ();
 sg13g2_fill_2 FILLER_70_93 ();
 sg13g2_decap_4 FILLER_70_121 ();
 sg13g2_fill_2 FILLER_70_142 ();
 sg13g2_fill_1 FILLER_70_144 ();
 sg13g2_fill_2 FILLER_70_154 ();
 sg13g2_fill_2 FILLER_70_161 ();
 sg13g2_fill_2 FILLER_70_182 ();
 sg13g2_fill_1 FILLER_70_202 ();
 sg13g2_fill_2 FILLER_70_212 ();
 sg13g2_fill_1 FILLER_70_214 ();
 sg13g2_decap_4 FILLER_70_219 ();
 sg13g2_fill_2 FILLER_70_223 ();
 sg13g2_fill_2 FILLER_70_234 ();
 sg13g2_fill_1 FILLER_70_236 ();
 sg13g2_decap_4 FILLER_70_242 ();
 sg13g2_fill_2 FILLER_70_251 ();
 sg13g2_fill_1 FILLER_70_253 ();
 sg13g2_decap_4 FILLER_70_267 ();
 sg13g2_fill_1 FILLER_70_283 ();
 sg13g2_fill_1 FILLER_70_289 ();
 sg13g2_decap_8 FILLER_70_295 ();
 sg13g2_decap_4 FILLER_70_302 ();
 sg13g2_fill_2 FILLER_70_320 ();
 sg13g2_fill_1 FILLER_70_322 ();
 sg13g2_decap_4 FILLER_70_343 ();
 sg13g2_fill_2 FILLER_70_347 ();
 sg13g2_decap_8 FILLER_70_362 ();
 sg13g2_fill_2 FILLER_70_369 ();
 sg13g2_fill_1 FILLER_70_371 ();
 sg13g2_fill_2 FILLER_70_430 ();
 sg13g2_fill_1 FILLER_70_489 ();
 sg13g2_decap_4 FILLER_70_503 ();
 sg13g2_fill_1 FILLER_70_515 ();
 sg13g2_decap_4 FILLER_70_521 ();
 sg13g2_decap_4 FILLER_70_551 ();
 sg13g2_fill_2 FILLER_70_590 ();
 sg13g2_decap_4 FILLER_70_597 ();
 sg13g2_fill_2 FILLER_70_601 ();
 sg13g2_fill_2 FILLER_70_607 ();
 sg13g2_fill_1 FILLER_70_609 ();
 sg13g2_fill_2 FILLER_70_644 ();
 sg13g2_fill_2 FILLER_70_661 ();
 sg13g2_fill_1 FILLER_70_679 ();
 sg13g2_fill_2 FILLER_70_684 ();
 sg13g2_fill_1 FILLER_70_686 ();
 sg13g2_fill_2 FILLER_70_696 ();
 sg13g2_fill_1 FILLER_70_702 ();
 sg13g2_fill_2 FILLER_70_742 ();
 sg13g2_fill_1 FILLER_70_744 ();
 sg13g2_fill_1 FILLER_70_757 ();
 sg13g2_fill_1 FILLER_70_776 ();
 sg13g2_decap_4 FILLER_70_807 ();
 sg13g2_fill_2 FILLER_70_811 ();
 sg13g2_fill_1 FILLER_70_822 ();
 sg13g2_fill_1 FILLER_70_827 ();
 sg13g2_decap_8 FILLER_70_833 ();
 sg13g2_decap_8 FILLER_70_840 ();
 sg13g2_decap_8 FILLER_70_847 ();
 sg13g2_decap_8 FILLER_70_854 ();
 sg13g2_fill_1 FILLER_70_861 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_2 ();
 sg13g2_decap_4 FILLER_71_110 ();
 sg13g2_fill_1 FILLER_71_114 ();
 sg13g2_fill_2 FILLER_71_132 ();
 sg13g2_fill_2 FILLER_71_161 ();
 sg13g2_fill_2 FILLER_71_172 ();
 sg13g2_decap_4 FILLER_71_193 ();
 sg13g2_fill_2 FILLER_71_203 ();
 sg13g2_fill_1 FILLER_71_205 ();
 sg13g2_fill_2 FILLER_71_216 ();
 sg13g2_fill_1 FILLER_71_218 ();
 sg13g2_fill_2 FILLER_71_239 ();
 sg13g2_fill_1 FILLER_71_241 ();
 sg13g2_fill_1 FILLER_71_252 ();
 sg13g2_fill_2 FILLER_71_272 ();
 sg13g2_fill_2 FILLER_71_289 ();
 sg13g2_fill_2 FILLER_71_296 ();
 sg13g2_fill_1 FILLER_71_298 ();
 sg13g2_decap_8 FILLER_71_320 ();
 sg13g2_fill_2 FILLER_71_333 ();
 sg13g2_fill_1 FILLER_71_340 ();
 sg13g2_decap_8 FILLER_71_353 ();
 sg13g2_decap_8 FILLER_71_360 ();
 sg13g2_fill_1 FILLER_71_367 ();
 sg13g2_fill_2 FILLER_71_437 ();
 sg13g2_fill_1 FILLER_71_439 ();
 sg13g2_fill_2 FILLER_71_449 ();
 sg13g2_fill_1 FILLER_71_451 ();
 sg13g2_fill_2 FILLER_71_572 ();
 sg13g2_fill_1 FILLER_71_574 ();
 sg13g2_fill_1 FILLER_71_604 ();
 sg13g2_fill_1 FILLER_71_656 ();
 sg13g2_fill_2 FILLER_71_673 ();
 sg13g2_decap_4 FILLER_71_683 ();
 sg13g2_decap_4 FILLER_71_722 ();
 sg13g2_fill_2 FILLER_71_726 ();
 sg13g2_fill_2 FILLER_71_772 ();
 sg13g2_fill_1 FILLER_71_774 ();
 sg13g2_decap_8 FILLER_71_806 ();
 sg13g2_decap_8 FILLER_71_813 ();
 sg13g2_decap_8 FILLER_71_820 ();
 sg13g2_decap_8 FILLER_71_827 ();
 sg13g2_decap_8 FILLER_71_834 ();
 sg13g2_decap_8 FILLER_71_841 ();
 sg13g2_decap_8 FILLER_71_848 ();
 sg13g2_decap_8 FILLER_71_855 ();
 sg13g2_decap_4 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_63 ();
 sg13g2_fill_1 FILLER_72_65 ();
 sg13g2_fill_1 FILLER_72_71 ();
 sg13g2_decap_4 FILLER_72_98 ();
 sg13g2_fill_1 FILLER_72_102 ();
 sg13g2_fill_2 FILLER_72_129 ();
 sg13g2_fill_1 FILLER_72_131 ();
 sg13g2_fill_2 FILLER_72_155 ();
 sg13g2_fill_1 FILLER_72_157 ();
 sg13g2_fill_1 FILLER_72_184 ();
 sg13g2_fill_1 FILLER_72_212 ();
 sg13g2_fill_1 FILLER_72_233 ();
 sg13g2_fill_1 FILLER_72_244 ();
 sg13g2_fill_2 FILLER_72_258 ();
 sg13g2_fill_1 FILLER_72_260 ();
 sg13g2_fill_2 FILLER_72_303 ();
 sg13g2_fill_2 FILLER_72_326 ();
 sg13g2_fill_1 FILLER_72_334 ();
 sg13g2_decap_8 FILLER_72_356 ();
 sg13g2_fill_2 FILLER_72_363 ();
 sg13g2_fill_1 FILLER_72_365 ();
 sg13g2_fill_2 FILLER_72_392 ();
 sg13g2_fill_1 FILLER_72_394 ();
 sg13g2_fill_1 FILLER_72_419 ();
 sg13g2_fill_2 FILLER_72_493 ();
 sg13g2_fill_1 FILLER_72_495 ();
 sg13g2_fill_1 FILLER_72_518 ();
 sg13g2_fill_2 FILLER_72_554 ();
 sg13g2_fill_1 FILLER_72_556 ();
 sg13g2_decap_8 FILLER_72_561 ();
 sg13g2_fill_2 FILLER_72_586 ();
 sg13g2_fill_1 FILLER_72_588 ();
 sg13g2_fill_1 FILLER_72_620 ();
 sg13g2_fill_2 FILLER_72_669 ();
 sg13g2_fill_2 FILLER_72_702 ();
 sg13g2_fill_1 FILLER_72_704 ();
 sg13g2_fill_2 FILLER_72_788 ();
 sg13g2_fill_1 FILLER_72_790 ();
 sg13g2_decap_8 FILLER_72_795 ();
 sg13g2_decap_8 FILLER_72_802 ();
 sg13g2_decap_8 FILLER_72_809 ();
 sg13g2_decap_8 FILLER_72_816 ();
 sg13g2_decap_8 FILLER_72_823 ();
 sg13g2_decap_8 FILLER_72_830 ();
 sg13g2_decap_8 FILLER_72_837 ();
 sg13g2_decap_8 FILLER_72_844 ();
 sg13g2_decap_8 FILLER_72_851 ();
 sg13g2_decap_4 FILLER_72_858 ();
 sg13g2_fill_1 FILLER_73_74 ();
 sg13g2_fill_1 FILLER_73_106 ();
 sg13g2_fill_2 FILLER_73_133 ();
 sg13g2_fill_1 FILLER_73_152 ();
 sg13g2_fill_1 FILLER_73_190 ();
 sg13g2_fill_1 FILLER_73_196 ();
 sg13g2_fill_1 FILLER_73_230 ();
 sg13g2_decap_8 FILLER_73_242 ();
 sg13g2_decap_8 FILLER_73_249 ();
 sg13g2_fill_2 FILLER_73_256 ();
 sg13g2_decap_4 FILLER_73_278 ();
 sg13g2_fill_2 FILLER_73_292 ();
 sg13g2_fill_1 FILLER_73_294 ();
 sg13g2_fill_2 FILLER_73_300 ();
 sg13g2_fill_1 FILLER_73_302 ();
 sg13g2_fill_1 FILLER_73_308 ();
 sg13g2_decap_8 FILLER_73_323 ();
 sg13g2_fill_1 FILLER_73_330 ();
 sg13g2_fill_2 FILLER_73_336 ();
 sg13g2_fill_1 FILLER_73_338 ();
 sg13g2_decap_8 FILLER_73_351 ();
 sg13g2_fill_2 FILLER_73_419 ();
 sg13g2_fill_1 FILLER_73_435 ();
 sg13g2_fill_2 FILLER_73_450 ();
 sg13g2_decap_4 FILLER_73_458 ();
 sg13g2_fill_1 FILLER_73_462 ();
 sg13g2_fill_1 FILLER_73_468 ();
 sg13g2_fill_1 FILLER_73_532 ();
 sg13g2_fill_2 FILLER_73_625 ();
 sg13g2_fill_1 FILLER_73_635 ();
 sg13g2_decap_8 FILLER_73_640 ();
 sg13g2_decap_8 FILLER_73_647 ();
 sg13g2_fill_1 FILLER_73_719 ();
 sg13g2_fill_2 FILLER_73_729 ();
 sg13g2_fill_2 FILLER_73_738 ();
 sg13g2_fill_1 FILLER_73_740 ();
 sg13g2_fill_2 FILLER_73_774 ();
 sg13g2_fill_1 FILLER_73_776 ();
 sg13g2_decap_8 FILLER_73_794 ();
 sg13g2_decap_8 FILLER_73_801 ();
 sg13g2_decap_8 FILLER_73_808 ();
 sg13g2_decap_8 FILLER_73_815 ();
 sg13g2_decap_8 FILLER_73_822 ();
 sg13g2_decap_8 FILLER_73_829 ();
 sg13g2_decap_8 FILLER_73_836 ();
 sg13g2_decap_8 FILLER_73_843 ();
 sg13g2_decap_8 FILLER_73_850 ();
 sg13g2_decap_4 FILLER_73_857 ();
 sg13g2_fill_1 FILLER_73_861 ();
 sg13g2_fill_2 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_2 ();
 sg13g2_fill_2 FILLER_74_86 ();
 sg13g2_fill_1 FILLER_74_88 ();
 sg13g2_fill_2 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_122 ();
 sg13g2_fill_1 FILLER_74_129 ();
 sg13g2_fill_2 FILLER_74_174 ();
 sg13g2_fill_2 FILLER_74_193 ();
 sg13g2_decap_4 FILLER_74_213 ();
 sg13g2_fill_1 FILLER_74_217 ();
 sg13g2_decap_8 FILLER_74_269 ();
 sg13g2_fill_2 FILLER_74_276 ();
 sg13g2_fill_1 FILLER_74_278 ();
 sg13g2_fill_2 FILLER_74_317 ();
 sg13g2_fill_1 FILLER_74_319 ();
 sg13g2_decap_8 FILLER_74_353 ();
 sg13g2_decap_8 FILLER_74_360 ();
 sg13g2_fill_2 FILLER_74_367 ();
 sg13g2_decap_4 FILLER_74_373 ();
 sg13g2_fill_2 FILLER_74_466 ();
 sg13g2_fill_2 FILLER_74_482 ();
 sg13g2_fill_1 FILLER_74_484 ();
 sg13g2_fill_2 FILLER_74_494 ();
 sg13g2_fill_1 FILLER_74_496 ();
 sg13g2_fill_2 FILLER_74_530 ();
 sg13g2_fill_2 FILLER_74_538 ();
 sg13g2_fill_1 FILLER_74_540 ();
 sg13g2_fill_2 FILLER_74_568 ();
 sg13g2_fill_1 FILLER_74_570 ();
 sg13g2_decap_4 FILLER_74_577 ();
 sg13g2_fill_1 FILLER_74_591 ();
 sg13g2_fill_2 FILLER_74_613 ();
 sg13g2_fill_1 FILLER_74_624 ();
 sg13g2_fill_1 FILLER_74_733 ();
 sg13g2_fill_2 FILLER_74_760 ();
 sg13g2_decap_8 FILLER_74_788 ();
 sg13g2_decap_8 FILLER_74_795 ();
 sg13g2_decap_8 FILLER_74_802 ();
 sg13g2_decap_8 FILLER_74_809 ();
 sg13g2_decap_8 FILLER_74_816 ();
 sg13g2_decap_8 FILLER_74_823 ();
 sg13g2_decap_8 FILLER_74_830 ();
 sg13g2_decap_8 FILLER_74_837 ();
 sg13g2_decap_8 FILLER_74_844 ();
 sg13g2_decap_8 FILLER_74_851 ();
 sg13g2_decap_4 FILLER_74_858 ();
 sg13g2_fill_2 FILLER_75_52 ();
 sg13g2_fill_1 FILLER_75_54 ();
 sg13g2_fill_2 FILLER_75_77 ();
 sg13g2_fill_2 FILLER_75_96 ();
 sg13g2_decap_8 FILLER_75_220 ();
 sg13g2_decap_4 FILLER_75_227 ();
 sg13g2_decap_4 FILLER_75_282 ();
 sg13g2_fill_1 FILLER_75_286 ();
 sg13g2_fill_2 FILLER_75_292 ();
 sg13g2_fill_1 FILLER_75_294 ();
 sg13g2_fill_2 FILLER_75_304 ();
 sg13g2_decap_8 FILLER_75_309 ();
 sg13g2_fill_1 FILLER_75_316 ();
 sg13g2_decap_8 FILLER_75_344 ();
 sg13g2_decap_8 FILLER_75_457 ();
 sg13g2_fill_1 FILLER_75_464 ();
 sg13g2_fill_1 FILLER_75_473 ();
 sg13g2_fill_1 FILLER_75_590 ();
 sg13g2_fill_1 FILLER_75_603 ();
 sg13g2_fill_2 FILLER_75_651 ();
 sg13g2_fill_2 FILLER_75_675 ();
 sg13g2_fill_2 FILLER_75_682 ();
 sg13g2_fill_1 FILLER_75_691 ();
 sg13g2_fill_1 FILLER_75_696 ();
 sg13g2_fill_2 FILLER_75_706 ();
 sg13g2_fill_1 FILLER_75_720 ();
 sg13g2_decap_4 FILLER_75_763 ();
 sg13g2_fill_2 FILLER_75_775 ();
 sg13g2_decap_8 FILLER_75_803 ();
 sg13g2_decap_8 FILLER_75_810 ();
 sg13g2_decap_8 FILLER_75_817 ();
 sg13g2_decap_8 FILLER_75_824 ();
 sg13g2_decap_8 FILLER_75_831 ();
 sg13g2_decap_8 FILLER_75_838 ();
 sg13g2_decap_8 FILLER_75_845 ();
 sg13g2_decap_8 FILLER_75_852 ();
 sg13g2_fill_2 FILLER_75_859 ();
 sg13g2_fill_1 FILLER_75_861 ();
 sg13g2_fill_2 FILLER_76_36 ();
 sg13g2_fill_1 FILLER_76_38 ();
 sg13g2_fill_1 FILLER_76_48 ();
 sg13g2_fill_1 FILLER_76_63 ();
 sg13g2_fill_1 FILLER_76_90 ();
 sg13g2_decap_8 FILLER_76_157 ();
 sg13g2_decap_8 FILLER_76_164 ();
 sg13g2_fill_1 FILLER_76_171 ();
 sg13g2_decap_4 FILLER_76_176 ();
 sg13g2_fill_2 FILLER_76_212 ();
 sg13g2_decap_4 FILLER_76_227 ();
 sg13g2_fill_1 FILLER_76_231 ();
 sg13g2_fill_2 FILLER_76_240 ();
 sg13g2_fill_1 FILLER_76_251 ();
 sg13g2_fill_2 FILLER_76_257 ();
 sg13g2_fill_1 FILLER_76_259 ();
 sg13g2_fill_1 FILLER_76_286 ();
 sg13g2_fill_2 FILLER_76_327 ();
 sg13g2_fill_1 FILLER_76_346 ();
 sg13g2_fill_1 FILLER_76_372 ();
 sg13g2_fill_2 FILLER_76_477 ();
 sg13g2_fill_1 FILLER_76_479 ();
 sg13g2_fill_1 FILLER_76_500 ();
 sg13g2_fill_2 FILLER_76_551 ();
 sg13g2_fill_2 FILLER_76_573 ();
 sg13g2_fill_2 FILLER_76_593 ();
 sg13g2_fill_2 FILLER_76_634 ();
 sg13g2_decap_4 FILLER_76_695 ();
 sg13g2_decap_4 FILLER_76_734 ();
 sg13g2_fill_2 FILLER_76_751 ();
 sg13g2_fill_1 FILLER_76_753 ();
 sg13g2_fill_1 FILLER_76_766 ();
 sg13g2_fill_2 FILLER_76_783 ();
 sg13g2_fill_1 FILLER_76_785 ();
 sg13g2_decap_8 FILLER_76_799 ();
 sg13g2_decap_8 FILLER_76_806 ();
 sg13g2_decap_8 FILLER_76_813 ();
 sg13g2_decap_8 FILLER_76_820 ();
 sg13g2_decap_8 FILLER_76_827 ();
 sg13g2_decap_8 FILLER_76_834 ();
 sg13g2_decap_8 FILLER_76_841 ();
 sg13g2_decap_8 FILLER_76_848 ();
 sg13g2_decap_8 FILLER_76_855 ();
 sg13g2_fill_2 FILLER_77_26 ();
 sg13g2_fill_1 FILLER_77_28 ();
 sg13g2_fill_1 FILLER_77_81 ();
 sg13g2_fill_2 FILLER_77_102 ();
 sg13g2_decap_8 FILLER_77_113 ();
 sg13g2_decap_4 FILLER_77_120 ();
 sg13g2_fill_1 FILLER_77_124 ();
 sg13g2_decap_8 FILLER_77_159 ();
 sg13g2_fill_2 FILLER_77_166 ();
 sg13g2_fill_1 FILLER_77_168 ();
 sg13g2_fill_2 FILLER_77_182 ();
 sg13g2_fill_1 FILLER_77_219 ();
 sg13g2_fill_2 FILLER_77_238 ();
 sg13g2_fill_1 FILLER_77_240 ();
 sg13g2_fill_2 FILLER_77_254 ();
 sg13g2_decap_4 FILLER_77_264 ();
 sg13g2_fill_2 FILLER_77_268 ();
 sg13g2_decap_8 FILLER_77_275 ();
 sg13g2_fill_2 FILLER_77_287 ();
 sg13g2_fill_1 FILLER_77_289 ();
 sg13g2_fill_1 FILLER_77_307 ();
 sg13g2_fill_2 FILLER_77_325 ();
 sg13g2_fill_1 FILLER_77_342 ();
 sg13g2_fill_1 FILLER_77_558 ();
 sg13g2_fill_1 FILLER_77_603 ();
 sg13g2_fill_2 FILLER_77_627 ();
 sg13g2_fill_2 FILLER_77_712 ();
 sg13g2_fill_1 FILLER_77_714 ();
 sg13g2_decap_8 FILLER_77_741 ();
 sg13g2_fill_2 FILLER_77_748 ();
 sg13g2_decap_8 FILLER_77_802 ();
 sg13g2_decap_8 FILLER_77_809 ();
 sg13g2_decap_8 FILLER_77_816 ();
 sg13g2_decap_8 FILLER_77_823 ();
 sg13g2_decap_8 FILLER_77_830 ();
 sg13g2_decap_8 FILLER_77_837 ();
 sg13g2_decap_8 FILLER_77_844 ();
 sg13g2_decap_8 FILLER_77_851 ();
 sg13g2_decap_4 FILLER_77_858 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_7 ();
 sg13g2_fill_1 FILLER_78_34 ();
 sg13g2_fill_2 FILLER_78_44 ();
 sg13g2_fill_1 FILLER_78_46 ();
 sg13g2_fill_2 FILLER_78_59 ();
 sg13g2_decap_8 FILLER_78_92 ();
 sg13g2_fill_2 FILLER_78_99 ();
 sg13g2_fill_1 FILLER_78_101 ();
 sg13g2_decap_8 FILLER_78_106 ();
 sg13g2_decap_8 FILLER_78_113 ();
 sg13g2_decap_8 FILLER_78_151 ();
 sg13g2_decap_4 FILLER_78_158 ();
 sg13g2_decap_4 FILLER_78_188 ();
 sg13g2_fill_1 FILLER_78_201 ();
 sg13g2_fill_1 FILLER_78_214 ();
 sg13g2_fill_2 FILLER_78_224 ();
 sg13g2_fill_1 FILLER_78_235 ();
 sg13g2_decap_4 FILLER_78_244 ();
 sg13g2_fill_1 FILLER_78_248 ();
 sg13g2_decap_8 FILLER_78_258 ();
 sg13g2_fill_1 FILLER_78_305 ();
 sg13g2_fill_2 FILLER_78_353 ();
 sg13g2_fill_1 FILLER_78_394 ();
 sg13g2_fill_2 FILLER_78_421 ();
 sg13g2_fill_1 FILLER_78_479 ();
 sg13g2_fill_1 FILLER_78_506 ();
 sg13g2_fill_1 FILLER_78_533 ();
 sg13g2_fill_1 FILLER_78_612 ();
 sg13g2_fill_2 FILLER_78_625 ();
 sg13g2_fill_1 FILLER_78_646 ();
 sg13g2_decap_8 FILLER_78_673 ();
 sg13g2_fill_2 FILLER_78_680 ();
 sg13g2_fill_1 FILLER_78_682 ();
 sg13g2_fill_2 FILLER_78_709 ();
 sg13g2_fill_1 FILLER_78_711 ();
 sg13g2_decap_8 FILLER_78_738 ();
 sg13g2_decap_8 FILLER_78_745 ();
 sg13g2_decap_8 FILLER_78_752 ();
 sg13g2_fill_2 FILLER_78_759 ();
 sg13g2_fill_2 FILLER_78_765 ();
 sg13g2_fill_1 FILLER_78_767 ();
 sg13g2_decap_8 FILLER_78_775 ();
 sg13g2_decap_4 FILLER_78_782 ();
 sg13g2_decap_8 FILLER_78_799 ();
 sg13g2_decap_8 FILLER_78_806 ();
 sg13g2_decap_8 FILLER_78_813 ();
 sg13g2_decap_8 FILLER_78_820 ();
 sg13g2_decap_8 FILLER_78_827 ();
 sg13g2_decap_8 FILLER_78_834 ();
 sg13g2_decap_8 FILLER_78_841 ();
 sg13g2_decap_8 FILLER_78_848 ();
 sg13g2_decap_8 FILLER_78_855 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_fill_1 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_83 ();
 sg13g2_decap_8 FILLER_79_90 ();
 sg13g2_decap_8 FILLER_79_97 ();
 sg13g2_decap_8 FILLER_79_104 ();
 sg13g2_decap_8 FILLER_79_111 ();
 sg13g2_decap_8 FILLER_79_118 ();
 sg13g2_decap_8 FILLER_79_125 ();
 sg13g2_decap_8 FILLER_79_132 ();
 sg13g2_decap_8 FILLER_79_139 ();
 sg13g2_decap_8 FILLER_79_146 ();
 sg13g2_fill_1 FILLER_79_179 ();
 sg13g2_fill_2 FILLER_79_215 ();
 sg13g2_fill_1 FILLER_79_217 ();
 sg13g2_fill_2 FILLER_79_222 ();
 sg13g2_fill_1 FILLER_79_224 ();
 sg13g2_fill_1 FILLER_79_251 ();
 sg13g2_fill_1 FILLER_79_307 ();
 sg13g2_fill_1 FILLER_79_317 ();
 sg13g2_fill_1 FILLER_79_327 ();
 sg13g2_fill_2 FILLER_79_377 ();
 sg13g2_fill_2 FILLER_79_388 ();
 sg13g2_fill_1 FILLER_79_390 ();
 sg13g2_fill_2 FILLER_79_408 ();
 sg13g2_fill_2 FILLER_79_431 ();
 sg13g2_fill_1 FILLER_79_433 ();
 sg13g2_fill_1 FILLER_79_538 ();
 sg13g2_fill_1 FILLER_79_585 ();
 sg13g2_fill_2 FILLER_79_595 ();
 sg13g2_decap_8 FILLER_79_680 ();
 sg13g2_decap_8 FILLER_79_700 ();
 sg13g2_decap_4 FILLER_79_707 ();
 sg13g2_fill_2 FILLER_79_711 ();
 sg13g2_decap_8 FILLER_79_726 ();
 sg13g2_decap_8 FILLER_79_733 ();
 sg13g2_decap_8 FILLER_79_740 ();
 sg13g2_decap_8 FILLER_79_747 ();
 sg13g2_decap_8 FILLER_79_754 ();
 sg13g2_decap_8 FILLER_79_761 ();
 sg13g2_decap_8 FILLER_79_768 ();
 sg13g2_decap_8 FILLER_79_775 ();
 sg13g2_decap_8 FILLER_79_782 ();
 sg13g2_decap_8 FILLER_79_789 ();
 sg13g2_decap_8 FILLER_79_796 ();
 sg13g2_decap_8 FILLER_79_803 ();
 sg13g2_decap_8 FILLER_79_810 ();
 sg13g2_decap_8 FILLER_79_817 ();
 sg13g2_decap_8 FILLER_79_824 ();
 sg13g2_decap_8 FILLER_79_831 ();
 sg13g2_decap_8 FILLER_79_838 ();
 sg13g2_decap_8 FILLER_79_845 ();
 sg13g2_decap_8 FILLER_79_852 ();
 sg13g2_fill_2 FILLER_79_859 ();
 sg13g2_fill_1 FILLER_79_861 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_fill_1 FILLER_80_21 ();
 sg13g2_fill_1 FILLER_80_36 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_4 FILLER_80_194 ();
 sg13g2_fill_2 FILLER_80_198 ();
 sg13g2_fill_2 FILLER_80_204 ();
 sg13g2_fill_1 FILLER_80_206 ();
 sg13g2_decap_8 FILLER_80_233 ();
 sg13g2_fill_1 FILLER_80_279 ();
 sg13g2_fill_1 FILLER_80_297 ();
 sg13g2_fill_1 FILLER_80_359 ();
 sg13g2_fill_2 FILLER_80_399 ();
 sg13g2_fill_1 FILLER_80_454 ();
 sg13g2_fill_1 FILLER_80_519 ();
 sg13g2_fill_2 FILLER_80_546 ();
 sg13g2_fill_1 FILLER_80_548 ();
 sg13g2_fill_1 FILLER_80_605 ();
 sg13g2_decap_8 FILLER_80_672 ();
 sg13g2_decap_8 FILLER_80_679 ();
 sg13g2_decap_8 FILLER_80_686 ();
 sg13g2_decap_8 FILLER_80_693 ();
 sg13g2_decap_8 FILLER_80_700 ();
 sg13g2_decap_8 FILLER_80_707 ();
 sg13g2_decap_8 FILLER_80_714 ();
 sg13g2_decap_8 FILLER_80_721 ();
 sg13g2_decap_8 FILLER_80_728 ();
 sg13g2_decap_8 FILLER_80_735 ();
 sg13g2_decap_8 FILLER_80_742 ();
 sg13g2_decap_8 FILLER_80_749 ();
 sg13g2_decap_8 FILLER_80_756 ();
 sg13g2_decap_8 FILLER_80_763 ();
 sg13g2_decap_8 FILLER_80_770 ();
 sg13g2_decap_8 FILLER_80_777 ();
 sg13g2_decap_8 FILLER_80_784 ();
 sg13g2_decap_8 FILLER_80_791 ();
 sg13g2_decap_8 FILLER_80_798 ();
 sg13g2_decap_8 FILLER_80_805 ();
 sg13g2_decap_8 FILLER_80_812 ();
 sg13g2_decap_8 FILLER_80_819 ();
 sg13g2_decap_8 FILLER_80_826 ();
 sg13g2_decap_8 FILLER_80_833 ();
 sg13g2_decap_8 FILLER_80_840 ();
 sg13g2_decap_8 FILLER_80_847 ();
 sg13g2_decap_8 FILLER_80_854 ();
 sg13g2_fill_1 FILLER_80_861 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule

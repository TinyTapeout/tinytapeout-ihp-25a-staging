module tt_um_log_afpm (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \A[0] ;
 wire \A[10] ;
 wire \A[11] ;
 wire \A[12] ;
 wire \A[13] ;
 wire \A[14] ;
 wire \A[15] ;
 wire \A[1] ;
 wire \A[2] ;
 wire \A[3] ;
 wire \A[4] ;
 wire \A[5] ;
 wire \A[6] ;
 wire \A[7] ;
 wire \A[8] ;
 wire \A[9] ;
 wire \B[0] ;
 wire \B[10] ;
 wire \B[11] ;
 wire \B[12] ;
 wire \B[13] ;
 wire \B[14] ;
 wire \B[15] ;
 wire \B[1] ;
 wire \B[2] ;
 wire \B[3] ;
 wire \B[4] ;
 wire \B[5] ;
 wire \B[6] ;
 wire \B[7] ;
 wire \B[8] ;
 wire \B[9] ;
 wire Ce;
 wire \Ea[0] ;
 wire \Ea[1] ;
 wire \Ea[2] ;
 wire \Ea[3] ;
 wire \Ea[4] ;
 wire \Eb[0] ;
 wire \Eb[1] ;
 wire \Eb[2] ;
 wire \Eb[3] ;
 wire \Eb[4] ;
 wire \Eout[0] ;
 wire \Eout[1] ;
 wire \Eout[2] ;
 wire \Eout[3] ;
 wire \Eout[4] ;
 wire \M1addout[0] ;
 wire \M1addout[10] ;
 wire \M1addout[1] ;
 wire \M1addout[2] ;
 wire \M1addout[3] ;
 wire \M1addout[4] ;
 wire \M1addout[5] ;
 wire \M1addout[6] ;
 wire \M1addout[7] ;
 wire \M1addout[8] ;
 wire \M1addout[9] ;
 wire \M1aout[0] ;
 wire \M1aout[1] ;
 wire \M1aout[2] ;
 wire \M1aout[3] ;
 wire \M1aout[4] ;
 wire \M1aout[5] ;
 wire \M1aout[6] ;
 wire \M1aout[7] ;
 wire \M1aout[8] ;
 wire \M1aout[9] ;
 wire \M1bout[0] ;
 wire \M1bout[1] ;
 wire \M1bout[2] ;
 wire \M1bout[3] ;
 wire \M1bout[4] ;
 wire \M1bout[5] ;
 wire \M1bout[6] ;
 wire \M1bout[7] ;
 wire \M1bout[8] ;
 wire \M1bout[9] ;
 wire \Ma[0] ;
 wire \Ma[1] ;
 wire \Ma[2] ;
 wire \Ma[3] ;
 wire \Ma[4] ;
 wire \Ma[5] ;
 wire \Ma[6] ;
 wire \Ma[7] ;
 wire \Ma[8] ;
 wire \Ma[9] ;
 wire \Mb[0] ;
 wire \Mb[1] ;
 wire \Mb[2] ;
 wire \Mb[3] ;
 wire \Mb[4] ;
 wire \Mb[5] ;
 wire \Mb[6] ;
 wire \Mb[7] ;
 wire \Mb[8] ;
 wire \Mb[9] ;
 wire \Mout[0] ;
 wire \Mout[1] ;
 wire \Mout[2] ;
 wire \Mout[3] ;
 wire \Mout[4] ;
 wire \Mout[5] ;
 wire \Mout[6] ;
 wire \Mout[7] ;
 wire \Mout[8] ;
 wire \Mout[9] ;
 wire Sa;
 wire Sb;
 wire Sout;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire clknet_0_clk;
 wire \byte_count[0] ;
 wire \byte_count[1] ;
 wire \result[0] ;
 wire \result[10] ;
 wire \result[11] ;
 wire \result[12] ;
 wire \result[13] ;
 wire \result[14] ;
 wire \result[15] ;
 wire \result[1] ;
 wire \result[2] ;
 wire \result[3] ;
 wire \result[4] ;
 wire \result[5] ;
 wire \result[6] ;
 wire \result[7] ;
 wire \result[8] ;
 wire \result[9] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire \state[4] ;
 wire \state[5] ;
 wire \state[6] ;
 wire \state[7] ;
 wire \state[8] ;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;

 sg13g2_inv_1 _1128_ (.Y(_0268_),
    .A(\result[15] ));
 sg13g2_inv_1 _1129_ (.Y(_0269_),
    .A(net212));
 sg13g2_inv_1 _1130_ (.Y(_0270_),
    .A(\result[14] ));
 sg13g2_inv_1 _1131_ (.Y(_0271_),
    .A(net190));
 sg13g2_inv_1 _1132_ (.Y(_0272_),
    .A(net261));
 sg13g2_inv_1 _1133_ (.Y(_0273_),
    .A(net185));
 sg13g2_inv_1 _1134_ (.Y(_0274_),
    .A(\result[12] ));
 sg13g2_inv_1 _1135_ (.Y(_0275_),
    .A(net214));
 sg13g2_inv_1 _1136_ (.Y(_0276_),
    .A(\result[11] ));
 sg13g2_inv_1 _1137_ (.Y(_0277_),
    .A(net183));
 sg13g2_inv_1 _1138_ (.Y(_0278_),
    .A(\result[10] ));
 sg13g2_inv_1 _1139_ (.Y(_0279_),
    .A(net188));
 sg13g2_inv_1 _1140_ (.Y(_0280_),
    .A(\result[9] ));
 sg13g2_inv_1 _1141_ (.Y(_0281_),
    .A(net236));
 sg13g2_inv_1 _1142_ (.Y(_0282_),
    .A(\result[8] ));
 sg13g2_inv_1 _1143_ (.Y(_0283_),
    .A(net201));
 sg13g2_inv_1 _1144_ (.Y(_0284_),
    .A(net239));
 sg13g2_inv_1 _1145_ (.Y(_0285_),
    .A(net247));
 sg13g2_inv_1 _1146_ (.Y(_0286_),
    .A(net257));
 sg13g2_inv_1 _1147_ (.Y(_0287_),
    .A(net410));
 sg13g2_inv_1 _1148_ (.Y(_0288_),
    .A(net238));
 sg13g2_inv_1 _1149_ (.Y(_0289_),
    .A(net366));
 sg13g2_inv_1 _1150_ (.Y(_0290_),
    .A(net352));
 sg13g2_inv_1 _1151_ (.Y(_0291_),
    .A(net220));
 sg13g2_inv_1 _1152_ (.Y(_0292_),
    .A(net209));
 sg13g2_inv_1 _1153_ (.Y(_0293_),
    .A(net348));
 sg13g2_inv_1 _1154_ (.Y(_0294_),
    .A(net3));
 sg13g2_inv_1 _1155_ (.Y(_0295_),
    .A(net2));
 sg13g2_inv_1 _1156_ (.Y(_0296_),
    .A(net5));
 sg13g2_inv_1 _1157_ (.Y(_0297_),
    .A(net4));
 sg13g2_inv_1 _1158_ (.Y(_0298_),
    .A(net7));
 sg13g2_inv_1 _1159_ (.Y(_0299_),
    .A(net6));
 sg13g2_inv_1 _1160_ (.Y(_0300_),
    .A(net9));
 sg13g2_inv_1 _1161_ (.Y(_0301_),
    .A(net8));
 sg13g2_inv_1 _1162_ (.Y(_0302_),
    .A(net229));
 sg13g2_inv_1 _1163_ (.Y(_0303_),
    .A(net308));
 sg13g2_inv_2 _1164_ (.Y(_0304_),
    .A(net312));
 sg13g2_inv_1 _1165_ (.Y(_0305_),
    .A(\Ma[7] ));
 sg13g2_inv_1 _1166_ (.Y(_0306_),
    .A(_0014_));
 sg13g2_inv_1 _1167_ (.Y(_0307_),
    .A(_0010_));
 sg13g2_inv_1 _1168_ (.Y(_0308_),
    .A(net299));
 sg13g2_inv_2 _1169_ (.Y(_0309_),
    .A(net302));
 sg13g2_inv_1 _1170_ (.Y(_0310_),
    .A(net411));
 sg13g2_inv_1 _1171_ (.Y(_0311_),
    .A(_0016_));
 sg13g2_inv_1 _1172_ (.Y(_0312_),
    .A(net318));
 sg13g2_inv_1 _1173_ (.Y(_0313_),
    .A(net325));
 sg13g2_inv_1 _1174_ (.Y(_0314_),
    .A(net322));
 sg13g2_inv_1 _1175_ (.Y(_0315_),
    .A(net414));
 sg13g2_inv_1 _1176_ (.Y(_0316_),
    .A(net379));
 sg13g2_inv_1 _1177_ (.Y(_0317_),
    .A(net427));
 sg13g2_inv_1 _1178_ (.Y(_0318_),
    .A(net429));
 sg13g2_inv_1 _1179_ (.Y(_0319_),
    .A(net392));
 sg13g2_inv_1 _1180_ (.Y(_0320_),
    .A(net422));
 sg13g2_inv_1 _1181_ (.Y(_0321_),
    .A(net365));
 sg13g2_inv_1 _1182_ (.Y(_0322_),
    .A(net407));
 sg13g2_inv_1 _1183_ (.Y(_0323_),
    .A(net428));
 sg13g2_inv_1 _1184_ (.Y(_0324_),
    .A(net425));
 sg13g2_inv_1 _1185_ (.Y(_0325_),
    .A(net408));
 sg13g2_inv_1 _1186_ (.Y(_0326_),
    .A(net420));
 sg13g2_inv_1 _1187_ (.Y(_0327_),
    .A(net418));
 sg13g2_inv_1 _1188_ (.Y(_0328_),
    .A(net423));
 sg13g2_inv_1 _1189_ (.Y(_0329_),
    .A(net416));
 sg13g2_inv_1 _1190_ (.Y(_0330_),
    .A(net437));
 sg13g2_inv_1 _1191_ (.Y(_0331_),
    .A(net376));
 sg13g2_inv_1 _1192_ (.Y(_0332_),
    .A(net388));
 sg13g2_inv_1 _1193_ (.Y(_0333_),
    .A(net435));
 sg13g2_inv_1 _1194_ (.Y(_0334_),
    .A(\M1aout[9] ));
 sg13g2_inv_1 _1195_ (.Y(_0335_),
    .A(net10));
 sg13g2_inv_1 _1196_ (.Y(_0336_),
    .A(net11));
 sg13g2_inv_1 _1197_ (.Y(_0337_),
    .A(net12));
 sg13g2_inv_1 _1198_ (.Y(_0338_),
    .A(net13));
 sg13g2_inv_1 _1199_ (.Y(_0339_),
    .A(net14));
 sg13g2_inv_1 _1200_ (.Y(_0340_),
    .A(net15));
 sg13g2_inv_1 _1201_ (.Y(_0341_),
    .A(net16));
 sg13g2_inv_1 _1202_ (.Y(_0342_),
    .A(net17));
 sg13g2_nor2b_1 _1203_ (.A(net368),
    .B_N(net332),
    .Y(_0343_));
 sg13g2_nand2b_1 _1204_ (.Y(_0344_),
    .B(net332),
    .A_N(net373));
 sg13g2_a21oi_1 _1205_ (.A1(net333),
    .A2(_0344_),
    .Y(_0345_),
    .B1(net340));
 sg13g2_nor2_1 _1206_ (.A(net342),
    .B(_0345_),
    .Y(_0007_));
 sg13g2_nor4_1 _1207_ (.A(net7),
    .B(net6),
    .C(net9),
    .D(net8),
    .Y(_0346_));
 sg13g2_nor3_1 _1208_ (.A(net3),
    .B(net2),
    .C(net5),
    .Y(_0347_));
 sg13g2_nand3_1 _1209_ (.B(_0346_),
    .C(_0347_),
    .A(_0297_),
    .Y(_0348_));
 sg13g2_a22oi_1 _1210_ (.Y(_0349_),
    .B1(_0348_),
    .B2(net229),
    .A2(_0344_),
    .A1(net209));
 sg13g2_nor2_1 _1211_ (.A(net341),
    .B(net230),
    .Y(_0008_));
 sg13g2_a21oi_1 _1212_ (.A1(net334),
    .A2(_0343_),
    .Y(_0350_),
    .B1(net341));
 sg13g2_o21ai_1 _1213_ (.B1(_0350_),
    .Y(_0006_),
    .A1(_0302_),
    .A2(_0348_));
 sg13g2_nand2_1 _1214_ (.Y(_0351_),
    .A(net351),
    .B(\state[7] ));
 sg13g2_inv_1 _1215_ (.Y(_0001_),
    .A(net288));
 sg13g2_nand2_1 _1216_ (.Y(_0352_),
    .A(net348),
    .B(\state[3] ));
 sg13g2_inv_1 _1217_ (.Y(_0002_),
    .A(net286));
 sg13g2_nand2_1 _1218_ (.Y(_0353_),
    .A(net348),
    .B(net205));
 sg13g2_inv_1 _1219_ (.Y(_0000_),
    .A(net279));
 sg13g2_nand2_1 _1220_ (.Y(_0354_),
    .A(net351),
    .B(\state[4] ));
 sg13g2_inv_2 _1221_ (.Y(_0005_),
    .A(net277));
 sg13g2_nand2_1 _1222_ (.Y(_0355_),
    .A(net209),
    .B(_0343_));
 sg13g2_nor2_1 _1223_ (.A(net341),
    .B(net274),
    .Y(_0004_));
 sg13g2_and2_1 _1224_ (.A(net348),
    .B(net186),
    .X(_0003_));
 sg13g2_and2_1 _1225_ (.A(net329),
    .B(\M1addout[0] ),
    .X(_0356_));
 sg13g2_xor2_1 _1226_ (.B(\M1addout[0] ),
    .A(net329),
    .X(_0357_));
 sg13g2_xnor2_1 _1227_ (.Y(_0358_),
    .A(net327),
    .B(_0357_));
 sg13g2_or2_1 _1228_ (.X(_0359_),
    .B(_0358_),
    .A(_0313_));
 sg13g2_a21oi_1 _1229_ (.A1(_0313_),
    .A2(_0358_),
    .Y(_0360_),
    .B1(net295));
 sg13g2_nand2_2 _1230_ (.Y(_0361_),
    .A(\M1addout[2] ),
    .B(\M1addout[1] ));
 sg13g2_or2_1 _1231_ (.X(_0362_),
    .B(\M1addout[1] ),
    .A(\M1addout[2] ));
 sg13g2_nand3_1 _1232_ (.B(_0361_),
    .C(_0362_),
    .A(net328),
    .Y(_0363_));
 sg13g2_a21oi_1 _1233_ (.A1(_0361_),
    .A2(_0362_),
    .Y(_0364_),
    .B1(net328));
 sg13g2_nor2_1 _1234_ (.A(net318),
    .B(_0364_),
    .Y(_0365_));
 sg13g2_a221oi_1 _1235_ (.B2(_0365_),
    .C1(net281),
    .B1(_0363_),
    .A1(_0359_),
    .Y(_0366_),
    .A2(_0360_));
 sg13g2_a21oi_1 _1236_ (.A1(_0291_),
    .A2(net281),
    .Y(_0023_),
    .B1(_0366_));
 sg13g2_a21oi_1 _1237_ (.A1(net326),
    .A2(_0357_),
    .Y(_0367_),
    .B1(_0356_));
 sg13g2_and2_1 _1238_ (.A(\M1addout[1] ),
    .B(\M1addout[4] ),
    .X(_0368_));
 sg13g2_xor2_1 _1239_ (.B(net328),
    .A(\M1addout[1] ),
    .X(_0369_));
 sg13g2_xnor2_1 _1240_ (.Y(_0370_),
    .A(net324),
    .B(_0369_));
 sg13g2_nor2_1 _1241_ (.A(_0367_),
    .B(_0370_),
    .Y(_0371_));
 sg13g2_xor2_1 _1242_ (.B(_0370_),
    .A(_0367_),
    .X(_0372_));
 sg13g2_xnor2_1 _1243_ (.Y(_0373_),
    .A(net322),
    .B(_0372_));
 sg13g2_or2_1 _1244_ (.X(_0374_),
    .B(_0373_),
    .A(_0359_));
 sg13g2_a21oi_1 _1245_ (.A1(_0359_),
    .A2(_0373_),
    .Y(_0375_),
    .B1(net296));
 sg13g2_and2_1 _1246_ (.A(\M1addout[2] ),
    .B(\M1addout[3] ),
    .X(_0376_));
 sg13g2_xor2_1 _1247_ (.B(net329),
    .A(\M1addout[2] ),
    .X(_0377_));
 sg13g2_xnor2_1 _1248_ (.Y(_0378_),
    .A(net327),
    .B(_0377_));
 sg13g2_a21oi_2 _1249_ (.B1(_0378_),
    .Y(_0379_),
    .A2(_0363_),
    .A1(_0361_));
 sg13g2_nand3_1 _1250_ (.B(_0363_),
    .C(_0378_),
    .A(_0361_),
    .Y(_0380_));
 sg13g2_nand2_1 _1251_ (.Y(_0381_),
    .A(net296),
    .B(_0380_));
 sg13g2_o21ai_1 _1252_ (.B1(net275),
    .Y(_0382_),
    .A1(_0379_),
    .A2(_0381_));
 sg13g2_a21oi_1 _1253_ (.A1(_0374_),
    .A2(_0375_),
    .Y(_0383_),
    .B1(_0382_));
 sg13g2_a21oi_1 _1254_ (.A1(_0290_),
    .A2(net281),
    .Y(_0024_),
    .B1(_0383_));
 sg13g2_a21oi_1 _1255_ (.A1(net324),
    .A2(_0369_),
    .Y(_0384_),
    .B1(_0368_));
 sg13g2_and2_1 _1256_ (.A(\M1addout[2] ),
    .B(net327),
    .X(_0385_));
 sg13g2_xor2_1 _1257_ (.B(net327),
    .A(\M1addout[2] ),
    .X(_0386_));
 sg13g2_xnor2_1 _1258_ (.Y(_0387_),
    .A(net323),
    .B(_0386_));
 sg13g2_nor2_1 _1259_ (.A(_0384_),
    .B(_0387_),
    .Y(_0388_));
 sg13g2_xor2_1 _1260_ (.B(_0387_),
    .A(_0384_),
    .X(_0389_));
 sg13g2_and2_1 _1261_ (.A(net320),
    .B(_0389_),
    .X(_0390_));
 sg13g2_xnor2_1 _1262_ (.Y(_0391_),
    .A(net320),
    .B(_0389_));
 sg13g2_a21oi_1 _1263_ (.A1(net322),
    .A2(_0372_),
    .Y(_0392_),
    .B1(_0371_));
 sg13g2_nor2_1 _1264_ (.A(_0391_),
    .B(_0392_),
    .Y(_0393_));
 sg13g2_xnor2_1 _1265_ (.Y(_0394_),
    .A(_0391_),
    .B(_0392_));
 sg13g2_nor2_1 _1266_ (.A(_0374_),
    .B(_0394_),
    .Y(_0395_));
 sg13g2_a21oi_1 _1267_ (.A1(_0374_),
    .A2(_0394_),
    .Y(_0396_),
    .B1(net296));
 sg13g2_nand2b_1 _1268_ (.Y(_0397_),
    .B(_0396_),
    .A_N(_0395_));
 sg13g2_and2_1 _1269_ (.A(\M1addout[4] ),
    .B(net329),
    .X(_0398_));
 sg13g2_xor2_1 _1270_ (.B(net329),
    .A(\M1addout[4] ),
    .X(_0399_));
 sg13g2_xnor2_1 _1271_ (.Y(_0400_),
    .A(net324),
    .B(_0399_));
 sg13g2_a21oi_1 _1272_ (.A1(net326),
    .A2(_0377_),
    .Y(_0401_),
    .B1(_0376_));
 sg13g2_nor2_1 _1273_ (.A(_0400_),
    .B(_0401_),
    .Y(_0402_));
 sg13g2_nand2_1 _1274_ (.Y(_0403_),
    .A(_0400_),
    .B(_0401_));
 sg13g2_nand2b_1 _1275_ (.Y(_0404_),
    .B(_0403_),
    .A_N(_0402_));
 sg13g2_xnor2_1 _1276_ (.Y(_0405_),
    .A(_0379_),
    .B(_0404_));
 sg13g2_a21oi_1 _1277_ (.A1(net296),
    .A2(_0405_),
    .Y(_0406_),
    .B1(net281));
 sg13g2_a22oi_1 _1278_ (.Y(_0025_),
    .B1(_0397_),
    .B2(_0406_),
    .A2(net281),
    .A1(_0289_));
 sg13g2_a21oi_1 _1279_ (.A1(net320),
    .A2(_0389_),
    .Y(_0407_),
    .B1(_0388_));
 sg13g2_and2_1 _1280_ (.A(net329),
    .B(net324),
    .X(_0408_));
 sg13g2_xor2_1 _1281_ (.B(net324),
    .A(net329),
    .X(_0409_));
 sg13g2_xnor2_1 _1282_ (.Y(_0410_),
    .A(net320),
    .B(_0409_));
 sg13g2_a21oi_2 _1283_ (.B1(_0385_),
    .Y(_0411_),
    .A2(_0386_),
    .A1(net322));
 sg13g2_nor2_1 _1284_ (.A(_0410_),
    .B(_0411_),
    .Y(_0412_));
 sg13g2_xor2_1 _1285_ (.B(_0411_),
    .A(_0410_),
    .X(_0413_));
 sg13g2_xnor2_1 _1286_ (.Y(_0414_),
    .A(_0022_),
    .B(_0413_));
 sg13g2_nor2b_1 _1287_ (.A(_0407_),
    .B_N(_0414_),
    .Y(_0415_));
 sg13g2_or3_1 _1288_ (.A(_0388_),
    .B(_0390_),
    .C(_0414_),
    .X(_0416_));
 sg13g2_xor2_1 _1289_ (.B(_0414_),
    .A(_0407_),
    .X(_0417_));
 sg13g2_nor2_1 _1290_ (.A(_0393_),
    .B(_0395_),
    .Y(_0418_));
 sg13g2_xor2_1 _1291_ (.B(_0418_),
    .A(_0417_),
    .X(_0419_));
 sg13g2_a21oi_2 _1292_ (.B1(_0402_),
    .Y(_0420_),
    .A2(_0403_),
    .A1(_0379_));
 sg13g2_and2_1 _1293_ (.A(net328),
    .B(net326),
    .X(_0421_));
 sg13g2_xor2_1 _1294_ (.B(net326),
    .A(net328),
    .X(_0422_));
 sg13g2_xnor2_1 _1295_ (.Y(_0423_),
    .A(net322),
    .B(_0422_));
 sg13g2_a21oi_2 _1296_ (.B1(_0398_),
    .Y(_0424_),
    .A2(_0399_),
    .A1(net325));
 sg13g2_or2_1 _1297_ (.X(_0425_),
    .B(_0424_),
    .A(_0423_));
 sg13g2_xnor2_1 _1298_ (.Y(_0426_),
    .A(_0423_),
    .B(_0424_));
 sg13g2_nand2_1 _1299_ (.Y(_0427_),
    .A(_0420_),
    .B(_0426_));
 sg13g2_o21ai_1 _1300_ (.B1(net295),
    .Y(_0428_),
    .A1(_0420_),
    .A2(_0426_));
 sg13g2_inv_1 _1301_ (.Y(_0429_),
    .A(_0428_));
 sg13g2_a221oi_1 _1302_ (.B2(_0429_),
    .C1(net280),
    .B1(_0427_),
    .A1(net318),
    .Y(_0430_),
    .A2(_0419_));
 sg13g2_a21oi_1 _1303_ (.A1(_0288_),
    .A2(net281),
    .Y(_0026_),
    .B1(_0430_));
 sg13g2_and2_1 _1304_ (.A(net328),
    .B(net322),
    .X(_0431_));
 sg13g2_xor2_1 _1305_ (.B(net322),
    .A(net328),
    .X(_0432_));
 sg13g2_xnor2_1 _1306_ (.Y(_0433_),
    .A(net319),
    .B(_0432_));
 sg13g2_a21oi_1 _1307_ (.A1(net320),
    .A2(_0409_),
    .Y(_0434_),
    .B1(_0408_));
 sg13g2_nor2_1 _1308_ (.A(_0433_),
    .B(_0434_),
    .Y(_0435_));
 sg13g2_xnor2_1 _1309_ (.Y(_0436_),
    .A(_0433_),
    .B(_0434_));
 sg13g2_a21oi_1 _1310_ (.A1(_0410_),
    .A2(_0411_),
    .Y(_0437_),
    .B1(net295));
 sg13g2_nor2_1 _1311_ (.A(_0412_),
    .B(_0437_),
    .Y(_0438_));
 sg13g2_nor2_1 _1312_ (.A(_0436_),
    .B(_0438_),
    .Y(_0439_));
 sg13g2_xnor2_1 _1313_ (.Y(_0440_),
    .A(_0436_),
    .B(_0438_));
 sg13g2_or3_1 _1314_ (.A(_0374_),
    .B(_0394_),
    .C(_0417_),
    .X(_0441_));
 sg13g2_a21oi_1 _1315_ (.A1(_0393_),
    .A2(_0416_),
    .Y(_0442_),
    .B1(_0415_));
 sg13g2_nand3_1 _1316_ (.B(_0441_),
    .C(_0442_),
    .A(_0440_),
    .Y(_0443_));
 sg13g2_a21oi_1 _1317_ (.A1(_0441_),
    .A2(_0442_),
    .Y(_0444_),
    .B1(_0440_));
 sg13g2_nand3b_1 _1318_ (.B(net317),
    .C(_0443_),
    .Y(_0445_),
    .A_N(_0444_));
 sg13g2_o21ai_1 _1319_ (.B1(_0425_),
    .Y(_0446_),
    .A1(_0420_),
    .A2(_0426_));
 sg13g2_and2_1 _1320_ (.A(net326),
    .B(net325),
    .X(_0447_));
 sg13g2_xor2_1 _1321_ (.B(net325),
    .A(net326),
    .X(_0448_));
 sg13g2_xnor2_1 _1322_ (.Y(_0449_),
    .A(net321),
    .B(_0448_));
 sg13g2_a21oi_1 _1323_ (.A1(net322),
    .A2(_0422_),
    .Y(_0450_),
    .B1(_0421_));
 sg13g2_or2_1 _1324_ (.X(_0451_),
    .B(_0450_),
    .A(_0449_));
 sg13g2_inv_1 _1325_ (.Y(_0452_),
    .A(_0451_));
 sg13g2_nand2_1 _1326_ (.Y(_0453_),
    .A(_0449_),
    .B(_0450_));
 sg13g2_nand2_1 _1327_ (.Y(_0454_),
    .A(_0451_),
    .B(_0453_));
 sg13g2_xnor2_1 _1328_ (.Y(_0455_),
    .A(_0446_),
    .B(_0454_));
 sg13g2_a21oi_1 _1329_ (.A1(net295),
    .A2(_0455_),
    .Y(_0456_),
    .B1(net280));
 sg13g2_a22oi_1 _1330_ (.Y(_0027_),
    .B1(_0445_),
    .B2(_0456_),
    .A2(net280),
    .A1(_0287_));
 sg13g2_nor2_1 _1331_ (.A(_0439_),
    .B(_0444_),
    .Y(_0457_));
 sg13g2_nand2_1 _1332_ (.Y(_0458_),
    .A(net326),
    .B(net321));
 sg13g2_xor2_1 _1333_ (.B(net320),
    .A(net326),
    .X(_0459_));
 sg13g2_a21oi_1 _1334_ (.A1(net319),
    .A2(_0432_),
    .Y(_0460_),
    .B1(_0431_));
 sg13g2_nand2b_1 _1335_ (.Y(_0461_),
    .B(_0459_),
    .A_N(_0460_));
 sg13g2_xnor2_1 _1336_ (.Y(_0462_),
    .A(_0459_),
    .B(_0460_));
 sg13g2_or2_1 _1337_ (.X(_0463_),
    .B(_0462_),
    .A(_0435_));
 sg13g2_nand2_1 _1338_ (.Y(_0464_),
    .A(_0435_),
    .B(_0462_));
 sg13g2_nand2_1 _1339_ (.Y(_0465_),
    .A(_0463_),
    .B(_0464_));
 sg13g2_xor2_1 _1340_ (.B(_0465_),
    .A(_0457_),
    .X(_0466_));
 sg13g2_a21oi_1 _1341_ (.A1(_0446_),
    .A2(_0453_),
    .Y(_0467_),
    .B1(_0452_));
 sg13g2_xor2_1 _1342_ (.B(net323),
    .A(net324),
    .X(_0468_));
 sg13g2_xnor2_1 _1343_ (.Y(_0469_),
    .A(net317),
    .B(_0468_));
 sg13g2_a21oi_1 _1344_ (.A1(net321),
    .A2(_0448_),
    .Y(_0470_),
    .B1(_0447_));
 sg13g2_or2_1 _1345_ (.X(_0471_),
    .B(_0470_),
    .A(_0469_));
 sg13g2_xnor2_1 _1346_ (.Y(_0472_),
    .A(_0469_),
    .B(_0470_));
 sg13g2_nand2_1 _1347_ (.Y(_0473_),
    .A(_0467_),
    .B(_0472_));
 sg13g2_nor2_1 _1348_ (.A(_0467_),
    .B(_0472_),
    .Y(_0474_));
 sg13g2_nor2_1 _1349_ (.A(net317),
    .B(_0474_),
    .Y(_0475_));
 sg13g2_a221oi_1 _1350_ (.B2(_0475_),
    .C1(net279),
    .B1(_0473_),
    .A1(net317),
    .Y(_0476_),
    .A2(_0466_));
 sg13g2_a21oi_1 _1351_ (.A1(_0286_),
    .A2(net280),
    .Y(_0028_),
    .B1(_0476_));
 sg13g2_o21ai_1 _1352_ (.B1(_0464_),
    .Y(_0477_),
    .A1(_0436_),
    .A2(_0438_));
 sg13g2_o21ai_1 _1353_ (.B1(_0463_),
    .Y(_0478_),
    .A1(_0444_),
    .A2(_0477_));
 sg13g2_nand2_1 _1354_ (.Y(_0479_),
    .A(net295),
    .B(_0313_));
 sg13g2_xnor2_1 _1355_ (.Y(_0480_),
    .A(net319),
    .B(net324));
 sg13g2_nand3b_1 _1356_ (.B(_0461_),
    .C(_0458_),
    .Y(_0481_),
    .A_N(_0480_));
 sg13g2_nor2b_1 _1357_ (.A(_0458_),
    .B_N(_0480_),
    .Y(_0482_));
 sg13g2_inv_1 _1358_ (.Y(_0483_),
    .A(_0482_));
 sg13g2_nand2b_1 _1359_ (.Y(_0484_),
    .B(_0480_),
    .A_N(_0461_));
 sg13g2_nand3_1 _1360_ (.B(_0483_),
    .C(_0484_),
    .A(_0481_),
    .Y(_0485_));
 sg13g2_xor2_1 _1361_ (.B(_0485_),
    .A(_0478_),
    .X(_0486_));
 sg13g2_o21ai_1 _1362_ (.B1(_0471_),
    .Y(_0487_),
    .A1(_0467_),
    .A2(_0472_));
 sg13g2_xnor2_1 _1363_ (.Y(_0488_),
    .A(net323),
    .B(net321));
 sg13g2_nand2_1 _1364_ (.Y(_0489_),
    .A(net317),
    .B(net323));
 sg13g2_nand2_1 _1365_ (.Y(_0490_),
    .A(net323),
    .B(_0479_));
 sg13g2_a22oi_1 _1366_ (.Y(_0491_),
    .B1(_0479_),
    .B2(net323),
    .A2(_0468_),
    .A1(net318));
 sg13g2_nor2_1 _1367_ (.A(_0488_),
    .B(_0491_),
    .Y(_0492_));
 sg13g2_xor2_1 _1368_ (.B(_0491_),
    .A(_0488_),
    .X(_0493_));
 sg13g2_o21ai_1 _1369_ (.B1(net295),
    .Y(_0494_),
    .A1(_0487_),
    .A2(_0493_));
 sg13g2_a21o_1 _1370_ (.A2(_0493_),
    .A1(_0487_),
    .B1(_0494_),
    .X(_0495_));
 sg13g2_a21oi_1 _1371_ (.A1(net317),
    .A2(_0486_),
    .Y(_0496_),
    .B1(net279));
 sg13g2_a22oi_1 _1372_ (.Y(_0029_),
    .B1(_0495_),
    .B2(_0496_),
    .A2(net279),
    .A1(_0285_));
 sg13g2_o21ai_1 _1373_ (.B1(_0489_),
    .Y(_0497_),
    .A1(net317),
    .A2(_0468_));
 sg13g2_inv_1 _1374_ (.Y(_0498_),
    .A(_0497_));
 sg13g2_xor2_1 _1375_ (.B(_0497_),
    .A(_0482_),
    .X(_0499_));
 sg13g2_o21ai_1 _1376_ (.B1(_0484_),
    .Y(_0500_),
    .A1(_0478_),
    .A2(_0485_));
 sg13g2_xnor2_1 _1377_ (.Y(_0501_),
    .A(_0499_),
    .B(_0500_));
 sg13g2_nand2_1 _1378_ (.Y(_0502_),
    .A(net317),
    .B(_0501_));
 sg13g2_a21oi_1 _1379_ (.A1(_0487_),
    .A2(_0493_),
    .Y(_0503_),
    .B1(_0492_));
 sg13g2_o21ai_1 _1380_ (.B1(_0314_),
    .Y(_0504_),
    .A1(net319),
    .A2(net320));
 sg13g2_o21ai_1 _1381_ (.B1(net295),
    .Y(_0505_),
    .A1(_0503_),
    .A2(_0504_));
 sg13g2_a21oi_1 _1382_ (.A1(_0503_),
    .A2(_0504_),
    .Y(_0506_),
    .B1(_0505_));
 sg13g2_nor2_1 _1383_ (.A(net279),
    .B(_0506_),
    .Y(_0507_));
 sg13g2_a22oi_1 _1384_ (.Y(_0030_),
    .B1(_0502_),
    .B2(_0507_),
    .A2(net279),
    .A1(_0284_));
 sg13g2_nor2_1 _1385_ (.A(_0283_),
    .B(net275),
    .Y(_0508_));
 sg13g2_a21o_1 _1386_ (.A2(net321),
    .A1(net323),
    .B1(_0505_),
    .X(_0509_));
 sg13g2_or2_1 _1387_ (.X(_0510_),
    .B(_0499_),
    .A(_0485_));
 sg13g2_o21ai_1 _1388_ (.B1(_0484_),
    .Y(_0511_),
    .A1(_0483_),
    .A2(_0497_));
 sg13g2_o21ai_1 _1389_ (.B1(_0511_),
    .Y(_0512_),
    .A1(_0482_),
    .A2(_0498_));
 sg13g2_o21ai_1 _1390_ (.B1(_0512_),
    .Y(_0513_),
    .A1(_0478_),
    .A2(_0510_));
 sg13g2_xnor2_1 _1391_ (.Y(_0514_),
    .A(net321),
    .B(_0490_));
 sg13g2_or2_1 _1392_ (.X(_0515_),
    .B(_0514_),
    .A(_0513_));
 sg13g2_a21oi_1 _1393_ (.A1(_0513_),
    .A2(_0514_),
    .Y(_0516_),
    .B1(net295));
 sg13g2_a21oi_1 _1394_ (.A1(_0515_),
    .A2(_0516_),
    .Y(_0517_),
    .B1(net279));
 sg13g2_a21o_1 _1395_ (.A2(_0517_),
    .A1(_0509_),
    .B1(_0508_),
    .X(_0031_));
 sg13g2_nand2_1 _1396_ (.Y(_0518_),
    .A(net318),
    .B(net321));
 sg13g2_a22oi_1 _1397_ (.Y(_0032_),
    .B1(_0517_),
    .B2(_0518_),
    .A2(net279),
    .A1(_0281_));
 sg13g2_nor3_2 _1398_ (.A(\byte_count[1] ),
    .B(net332),
    .C(_0292_),
    .Y(_0519_));
 sg13g2_o21ai_1 _1399_ (.B1(net350),
    .Y(_0520_),
    .A1(net264),
    .A2(net271));
 sg13g2_a21oi_1 _1400_ (.A1(_0295_),
    .A2(net270),
    .Y(_0033_),
    .B1(_0520_));
 sg13g2_o21ai_1 _1401_ (.B1(net350),
    .Y(_0521_),
    .A1(net354),
    .A2(net271));
 sg13g2_a21oi_1 _1402_ (.A1(_0294_),
    .A2(net270),
    .Y(_0034_),
    .B1(_0521_));
 sg13g2_o21ai_1 _1403_ (.B1(net350),
    .Y(_0522_),
    .A1(net241),
    .A2(net271));
 sg13g2_a21oi_1 _1404_ (.A1(_0297_),
    .A2(net271),
    .Y(_0035_),
    .B1(_0522_));
 sg13g2_o21ai_1 _1405_ (.B1(net1),
    .Y(_0523_),
    .A1(net249),
    .A2(net271));
 sg13g2_a21oi_1 _1406_ (.A1(_0296_),
    .A2(net271),
    .Y(_0036_),
    .B1(_0523_));
 sg13g2_o21ai_1 _1407_ (.B1(net350),
    .Y(_0524_),
    .A1(net251),
    .A2(net271));
 sg13g2_a21oi_1 _1408_ (.A1(_0299_),
    .A2(net270),
    .Y(_0037_),
    .B1(_0524_));
 sg13g2_o21ai_1 _1409_ (.B1(net350),
    .Y(_0525_),
    .A1(net234),
    .A2(net270));
 sg13g2_a21oi_1 _1410_ (.A1(_0298_),
    .A2(net270),
    .Y(_0038_),
    .B1(_0525_));
 sg13g2_o21ai_1 _1411_ (.B1(net350),
    .Y(_0526_),
    .A1(net374),
    .A2(net270));
 sg13g2_a21oi_1 _1412_ (.A1(_0301_),
    .A2(net270),
    .Y(_0039_),
    .B1(_0526_));
 sg13g2_o21ai_1 _1413_ (.B1(net350),
    .Y(_0527_),
    .A1(net381),
    .A2(net270));
 sg13g2_a21oi_1 _1414_ (.A1(_0300_),
    .A2(net272),
    .Y(_0040_),
    .B1(_0527_));
 sg13g2_xnor2_1 _1415_ (.Y(_0528_),
    .A(net368),
    .B(net332));
 sg13g2_nor3_1 _1416_ (.A(_0292_),
    .B(net181),
    .C(_0528_),
    .Y(_0529_));
 sg13g2_a22oi_1 _1417_ (.Y(_0530_),
    .B1(net266),
    .B2(net2),
    .A2(net273),
    .A1(net396));
 sg13g2_nor2_1 _1418_ (.A(net343),
    .B(_0530_),
    .Y(_0041_));
 sg13g2_a22oi_1 _1419_ (.Y(_0531_),
    .B1(net266),
    .B2(net3),
    .A2(net273),
    .A1(net406));
 sg13g2_nor2_1 _1420_ (.A(net343),
    .B(_0531_),
    .Y(_0042_));
 sg13g2_a22oi_1 _1421_ (.Y(_0532_),
    .B1(net266),
    .B2(net4),
    .A2(net273),
    .A1(net246));
 sg13g2_nor2_1 _1422_ (.A(net343),
    .B(_0532_),
    .Y(_0043_));
 sg13g2_a22oi_1 _1423_ (.Y(_0533_),
    .B1(net266),
    .B2(net5),
    .A2(net273),
    .A1(net194));
 sg13g2_nor2_1 _1424_ (.A(net344),
    .B(_0533_),
    .Y(_0044_));
 sg13g2_a22oi_1 _1425_ (.Y(_0534_),
    .B1(net266),
    .B2(net6),
    .A2(net273),
    .A1(net208));
 sg13g2_nor2_1 _1426_ (.A(net343),
    .B(_0534_),
    .Y(_0045_));
 sg13g2_a22oi_1 _1427_ (.Y(_0535_),
    .B1(net266),
    .B2(net7),
    .A2(net273),
    .A1(net195));
 sg13g2_nor2_1 _1428_ (.A(net343),
    .B(_0535_),
    .Y(_0046_));
 sg13g2_a22oi_1 _1429_ (.Y(_0536_),
    .B1(net266),
    .B2(net8),
    .A2(net273),
    .A1(net222));
 sg13g2_nor2_1 _1430_ (.A(net343),
    .B(_0536_),
    .Y(_0047_));
 sg13g2_a22oi_1 _1431_ (.Y(_0537_),
    .B1(net266),
    .B2(net9),
    .A2(net273),
    .A1(net197));
 sg13g2_nor2_1 _1432_ (.A(net343),
    .B(_0537_),
    .Y(_0048_));
 sg13g2_o21ai_1 _1433_ (.B1(net350),
    .Y(_0538_),
    .A1(net243),
    .A2(net272));
 sg13g2_a21oi_1 _1434_ (.A1(_0335_),
    .A2(net272),
    .Y(_0049_),
    .B1(_0538_));
 sg13g2_o21ai_1 _1435_ (.B1(net351),
    .Y(_0539_),
    .A1(net259),
    .A2(net269));
 sg13g2_a21oi_1 _1436_ (.A1(_0336_),
    .A2(net269),
    .Y(_0050_),
    .B1(_0539_));
 sg13g2_o21ai_1 _1437_ (.B1(net351),
    .Y(_0540_),
    .A1(net192),
    .A2(net268));
 sg13g2_a21oi_1 _1438_ (.A1(_0337_),
    .A2(net268),
    .Y(_0051_),
    .B1(_0540_));
 sg13g2_o21ai_1 _1439_ (.B1(net351),
    .Y(_0541_),
    .A1(net210),
    .A2(net269));
 sg13g2_a21oi_1 _1440_ (.A1(_0338_),
    .A2(net269),
    .Y(_0052_),
    .B1(_0541_));
 sg13g2_o21ai_1 _1441_ (.B1(net351),
    .Y(_0542_),
    .A1(net363),
    .A2(net268));
 sg13g2_a21oi_1 _1442_ (.A1(_0339_),
    .A2(net269),
    .Y(_0053_),
    .B1(_0542_));
 sg13g2_o21ai_1 _1443_ (.B1(net351),
    .Y(_0543_),
    .A1(net386),
    .A2(net268));
 sg13g2_a21oi_1 _1444_ (.A1(_0340_),
    .A2(net269),
    .Y(_0054_),
    .B1(_0543_));
 sg13g2_o21ai_1 _1445_ (.B1(net348),
    .Y(_0544_),
    .A1(net218),
    .A2(net268));
 sg13g2_a21oi_1 _1446_ (.A1(_0341_),
    .A2(net268),
    .Y(_0055_),
    .B1(_0544_));
 sg13g2_o21ai_1 _1447_ (.B1(net348),
    .Y(_0545_),
    .A1(net399),
    .A2(net268));
 sg13g2_a21oi_1 _1448_ (.A1(_0342_),
    .A2(net268),
    .Y(_0056_),
    .B1(_0545_));
 sg13g2_a22oi_1 _1449_ (.Y(_0546_),
    .B1(net267),
    .B2(net10),
    .A2(net274),
    .A1(net263));
 sg13g2_nor2_1 _1450_ (.A(net344),
    .B(_0546_),
    .Y(_0057_));
 sg13g2_a22oi_1 _1451_ (.Y(_0547_),
    .B1(net267),
    .B2(net11),
    .A2(net274),
    .A1(net378));
 sg13g2_nor2_1 _1452_ (.A(net341),
    .B(_0547_),
    .Y(_0058_));
 sg13g2_a22oi_1 _1453_ (.Y(_0548_),
    .B1(net267),
    .B2(net12),
    .A2(net274),
    .A1(net203));
 sg13g2_nor2_1 _1454_ (.A(net341),
    .B(_0548_),
    .Y(_0059_));
 sg13g2_a22oi_1 _1455_ (.Y(_0549_),
    .B1(net267),
    .B2(net13),
    .A2(net274),
    .A1(net199));
 sg13g2_nor2_1 _1456_ (.A(net344),
    .B(_0549_),
    .Y(_0060_));
 sg13g2_a22oi_1 _1457_ (.Y(_0550_),
    .B1(net267),
    .B2(net14),
    .A2(net274),
    .A1(net217));
 sg13g2_nor2_1 _1458_ (.A(net344),
    .B(_0550_),
    .Y(_0061_));
 sg13g2_a22oi_1 _1459_ (.Y(_0551_),
    .B1(net267),
    .B2(net15),
    .A2(net274),
    .A1(net226));
 sg13g2_nor2_1 _1460_ (.A(net344),
    .B(_0551_),
    .Y(_0062_));
 sg13g2_a22oi_1 _1461_ (.Y(_0552_),
    .B1(_0529_),
    .B2(net16),
    .A2(_0355_),
    .A1(net360));
 sg13g2_nor2_1 _1462_ (.A(net343),
    .B(_0552_),
    .Y(_0063_));
 sg13g2_a22oi_1 _1463_ (.Y(_0553_),
    .B1(net267),
    .B2(net17),
    .A2(net274),
    .A1(net187));
 sg13g2_nor2_1 _1464_ (.A(net341),
    .B(_0553_),
    .Y(_0064_));
 sg13g2_nand2b_1 _1465_ (.Y(_0554_),
    .B(net404),
    .A_N(net334));
 sg13g2_nand2b_2 _1466_ (.Y(_0555_),
    .B(net333),
    .A_N(\byte_count[1] ));
 sg13g2_a21oi_1 _1467_ (.A1(net330),
    .A2(_0282_),
    .Y(_0556_),
    .B1(_0555_));
 sg13g2_o21ai_1 _1468_ (.B1(_0556_),
    .Y(_0557_),
    .A1(net330),
    .A2(net224));
 sg13g2_a21oi_1 _1469_ (.A1(_0554_),
    .A2(_0557_),
    .Y(_0065_),
    .B1(net345));
 sg13g2_nand2b_1 _1470_ (.Y(_0558_),
    .B(net412),
    .A_N(net334));
 sg13g2_a21oi_1 _1471_ (.A1(net330),
    .A2(_0280_),
    .Y(_0559_),
    .B1(_0555_));
 sg13g2_o21ai_1 _1472_ (.B1(_0559_),
    .Y(_0560_),
    .A1(net331),
    .A2(\result[1] ));
 sg13g2_a21oi_1 _1473_ (.A1(_0558_),
    .A2(_0560_),
    .Y(_0066_),
    .B1(net341));
 sg13g2_nand2b_1 _1474_ (.Y(_0561_),
    .B(net357),
    .A_N(net333));
 sg13g2_a21oi_1 _1475_ (.A1(net332),
    .A2(_0278_),
    .Y(_0562_),
    .B1(_0555_));
 sg13g2_o21ai_1 _1476_ (.B1(_0562_),
    .Y(_0563_),
    .A1(net332),
    .A2(\result[2] ));
 sg13g2_a21oi_1 _1477_ (.A1(net358),
    .A2(_0563_),
    .Y(_0067_),
    .B1(net342));
 sg13g2_nand2b_1 _1478_ (.Y(_0564_),
    .B(net394),
    .A_N(net334));
 sg13g2_a21oi_1 _1479_ (.A1(net330),
    .A2(_0276_),
    .Y(_0565_),
    .B1(_0555_));
 sg13g2_o21ai_1 _1480_ (.B1(_0565_),
    .Y(_0566_),
    .A1(net331),
    .A2(net256));
 sg13g2_a21oi_1 _1481_ (.A1(_0564_),
    .A2(_0566_),
    .Y(_0068_),
    .B1(net342));
 sg13g2_nand2b_1 _1482_ (.Y(_0567_),
    .B(net400),
    .A_N(net333));
 sg13g2_a21oi_1 _1483_ (.A1(net330),
    .A2(_0274_),
    .Y(_0568_),
    .B1(_0555_));
 sg13g2_o21ai_1 _1484_ (.B1(_0568_),
    .Y(_0569_),
    .A1(net330),
    .A2(net383));
 sg13g2_a21oi_1 _1485_ (.A1(_0567_),
    .A2(_0569_),
    .Y(_0069_),
    .B1(net342));
 sg13g2_nand2b_1 _1486_ (.Y(_0570_),
    .B(net402),
    .A_N(net333));
 sg13g2_a21oi_1 _1487_ (.A1(net331),
    .A2(_0272_),
    .Y(_0571_),
    .B1(_0555_));
 sg13g2_o21ai_1 _1488_ (.B1(_0571_),
    .Y(_0572_),
    .A1(net331),
    .A2(\result[5] ));
 sg13g2_a21oi_1 _1489_ (.A1(_0570_),
    .A2(_0572_),
    .Y(_0070_),
    .B1(net342));
 sg13g2_nand2b_1 _1490_ (.Y(_0573_),
    .B(net390),
    .A_N(net333));
 sg13g2_a21oi_1 _1491_ (.A1(net330),
    .A2(_0270_),
    .Y(_0574_),
    .B1(_0555_));
 sg13g2_o21ai_1 _1492_ (.B1(_0574_),
    .Y(_0575_),
    .A1(net330),
    .A2(\result[6] ));
 sg13g2_a21oi_1 _1493_ (.A1(_0573_),
    .A2(_0575_),
    .Y(_0071_),
    .B1(net342));
 sg13g2_nand2b_1 _1494_ (.Y(_0576_),
    .B(net369),
    .A_N(net333));
 sg13g2_a21oi_1 _1495_ (.A1(\byte_count[0] ),
    .A2(_0268_),
    .Y(_0577_),
    .B1(_0555_));
 sg13g2_o21ai_1 _1496_ (.B1(_0577_),
    .Y(_0578_),
    .A1(net331),
    .A2(\result[7] ));
 sg13g2_a21oi_1 _1497_ (.A1(net370),
    .A2(_0578_),
    .Y(_0072_),
    .B1(net342));
 sg13g2_o21ai_1 _1498_ (.B1(net347),
    .Y(_0579_),
    .A1(net335),
    .A2(net224));
 sg13g2_a21oi_1 _1499_ (.A1(net338),
    .A2(_0291_),
    .Y(_0073_),
    .B1(_0579_));
 sg13g2_o21ai_1 _1500_ (.B1(net347),
    .Y(_0580_),
    .A1(net335),
    .A2(\result[1] ));
 sg13g2_a21oi_1 _1501_ (.A1(net338),
    .A2(_0290_),
    .Y(_0074_),
    .B1(_0580_));
 sg13g2_o21ai_1 _1502_ (.B1(net348),
    .Y(_0581_),
    .A1(net339),
    .A2(\result[2] ));
 sg13g2_a21oi_1 _1503_ (.A1(net339),
    .A2(_0289_),
    .Y(_0075_),
    .B1(_0581_));
 sg13g2_o21ai_1 _1504_ (.B1(net347),
    .Y(_0582_),
    .A1(net339),
    .A2(net256));
 sg13g2_a21oi_1 _1505_ (.A1(net339),
    .A2(_0288_),
    .Y(_0076_),
    .B1(_0582_));
 sg13g2_o21ai_1 _1506_ (.B1(net346),
    .Y(_0583_),
    .A1(net337),
    .A2(net383));
 sg13g2_a21oi_1 _1507_ (.A1(net337),
    .A2(_0287_),
    .Y(_0077_),
    .B1(_0583_));
 sg13g2_o21ai_1 _1508_ (.B1(net346),
    .Y(_0584_),
    .A1(net336),
    .A2(\result[5] ));
 sg13g2_a21oi_1 _1509_ (.A1(net336),
    .A2(_0286_),
    .Y(_0078_),
    .B1(_0584_));
 sg13g2_o21ai_1 _1510_ (.B1(net346),
    .Y(_0585_),
    .A1(net336),
    .A2(\result[6] ));
 sg13g2_a21oi_1 _1511_ (.A1(net336),
    .A2(_0285_),
    .Y(_0079_),
    .B1(_0585_));
 sg13g2_o21ai_1 _1512_ (.B1(net346),
    .Y(_0586_),
    .A1(net335),
    .A2(\result[7] ));
 sg13g2_a21oi_1 _1513_ (.A1(net335),
    .A2(_0284_),
    .Y(_0080_),
    .B1(_0586_));
 sg13g2_o21ai_1 _1514_ (.B1(net346),
    .Y(_0587_),
    .A1(net335),
    .A2(\result[8] ));
 sg13g2_a21oi_1 _1515_ (.A1(net335),
    .A2(_0283_),
    .Y(_0081_),
    .B1(_0587_));
 sg13g2_o21ai_1 _1516_ (.B1(net346),
    .Y(_0588_),
    .A1(net335),
    .A2(\result[9] ));
 sg13g2_a21oi_1 _1517_ (.A1(net335),
    .A2(_0281_),
    .Y(_0082_),
    .B1(_0588_));
 sg13g2_o21ai_1 _1518_ (.B1(net349),
    .Y(_0589_),
    .A1(net340),
    .A2(\result[10] ));
 sg13g2_a21oi_1 _1519_ (.A1(net340),
    .A2(_0279_),
    .Y(_0083_),
    .B1(_0589_));
 sg13g2_o21ai_1 _1520_ (.B1(net347),
    .Y(_0590_),
    .A1(net337),
    .A2(\result[11] ));
 sg13g2_a21oi_1 _1521_ (.A1(net337),
    .A2(_0277_),
    .Y(_0084_),
    .B1(_0590_));
 sg13g2_o21ai_1 _1522_ (.B1(net346),
    .Y(_0591_),
    .A1(net336),
    .A2(\result[12] ));
 sg13g2_a21oi_1 _1523_ (.A1(net336),
    .A2(_0275_),
    .Y(_0085_),
    .B1(_0591_));
 sg13g2_o21ai_1 _1524_ (.B1(net347),
    .Y(_0592_),
    .A1(net339),
    .A2(net261));
 sg13g2_a21oi_1 _1525_ (.A1(net339),
    .A2(_0273_),
    .Y(_0086_),
    .B1(_0592_));
 sg13g2_o21ai_1 _1526_ (.B1(net346),
    .Y(_0593_),
    .A1(net336),
    .A2(\result[14] ));
 sg13g2_a21oi_1 _1527_ (.A1(net336),
    .A2(_0271_),
    .Y(_0087_),
    .B1(_0593_));
 sg13g2_o21ai_1 _1528_ (.B1(net348),
    .Y(_0594_),
    .A1(\result[15] ),
    .A2(net339));
 sg13g2_a21oi_1 _1529_ (.A1(_0269_),
    .A2(net339),
    .Y(_0088_),
    .B1(_0594_));
 sg13g2_or2_1 _1530_ (.X(_0595_),
    .B(net439),
    .A(net333));
 sg13g2_nor3_1 _1531_ (.A(net229),
    .B(net206),
    .C(_0595_),
    .Y(_0596_));
 sg13g2_a22oi_1 _1532_ (.Y(_0597_),
    .B1(_0596_),
    .B2(net332),
    .A2(_0595_),
    .A1(net181));
 sg13g2_nor2_1 _1533_ (.A(net341),
    .B(net182),
    .Y(_0089_));
 sg13g2_nor2b_1 _1534_ (.A(_0528_),
    .B_N(_0595_),
    .Y(_0598_));
 sg13g2_a21oi_1 _1535_ (.A1(net368),
    .A2(_0596_),
    .Y(_0599_),
    .B1(_0598_));
 sg13g2_nor2_1 _1536_ (.A(net342),
    .B(_0599_),
    .Y(_0090_));
 sg13g2_nand2_1 _1537_ (.Y(_0600_),
    .A(\Ma[0] ),
    .B(\Ma[2] ));
 sg13g2_xor2_1 _1538_ (.B(\Ma[2] ),
    .A(\Ma[0] ),
    .X(_0601_));
 sg13g2_nor2_1 _1539_ (.A(_0011_),
    .B(net312),
    .Y(_0602_));
 sg13g2_xor2_1 _1540_ (.B(_0602_),
    .A(_0601_),
    .X(_0603_));
 sg13g2_mux2_1 _1541_ (.A0(net316),
    .A1(\Ma[5] ),
    .S(net312),
    .X(_0604_));
 sg13g2_nand2_1 _1542_ (.Y(_0605_),
    .A(\Ma[0] ),
    .B(_0604_));
 sg13g2_o21ai_1 _1543_ (.B1(\Ma[9] ),
    .Y(_0606_),
    .A1(\Ma[0] ),
    .A2(_0604_));
 sg13g2_inv_1 _1544_ (.Y(_0607_),
    .A(_0606_));
 sg13g2_a221oi_1 _1545_ (.B2(_0607_),
    .C1(net286),
    .B1(_0605_),
    .A1(_0303_),
    .Y(_0608_),
    .A2(_0603_));
 sg13g2_a21oi_1 _1546_ (.A1(_0318_),
    .A2(net287),
    .Y(_0091_),
    .B1(_0608_));
 sg13g2_and2_1 _1547_ (.A(\Ma[4] ),
    .B(_0601_),
    .X(_0609_));
 sg13g2_nand2_1 _1548_ (.Y(_0610_),
    .A(net316),
    .B(\Ma[1] ));
 sg13g2_nor2_1 _1549_ (.A(net316),
    .B(\Ma[1] ),
    .Y(_0611_));
 sg13g2_xor2_1 _1550_ (.B(\Ma[1] ),
    .A(net316),
    .X(_0612_));
 sg13g2_xnor2_1 _1551_ (.Y(_0613_),
    .A(_0600_),
    .B(_0612_));
 sg13g2_xnor2_1 _1552_ (.Y(_0614_),
    .A(_0012_),
    .B(_0613_));
 sg13g2_nor2_1 _1553_ (.A(net309),
    .B(net312),
    .Y(_0615_));
 sg13g2_xor2_1 _1554_ (.B(_0614_),
    .A(_0609_),
    .X(_0616_));
 sg13g2_nand2_1 _1555_ (.Y(_0617_),
    .A(net311),
    .B(net313));
 sg13g2_mux2_1 _1556_ (.A0(net315),
    .A1(\Ma[6] ),
    .S(net312),
    .X(_0618_));
 sg13g2_nand2_1 _1557_ (.Y(_0619_),
    .A(\Ma[1] ),
    .B(_0618_));
 sg13g2_xnor2_1 _1558_ (.Y(_0620_),
    .A(\Ma[1] ),
    .B(_0618_));
 sg13g2_and2_1 _1559_ (.A(_0605_),
    .B(_0620_),
    .X(_0621_));
 sg13g2_o21ai_1 _1560_ (.B1(net309),
    .Y(_0622_),
    .A1(_0605_),
    .A2(_0620_));
 sg13g2_nor2_2 _1561_ (.A(\Ma[9] ),
    .B(_0304_),
    .Y(_0623_));
 sg13g2_o21ai_1 _1562_ (.B1(_0002_),
    .Y(_0624_),
    .A1(_0621_),
    .A2(_0622_));
 sg13g2_a221oi_1 _1563_ (.B2(_0613_),
    .C1(_0624_),
    .B1(_0623_),
    .A1(_0615_),
    .Y(_0625_),
    .A2(_0616_));
 sg13g2_a21oi_1 _1564_ (.A1(_0316_),
    .A2(net287),
    .Y(_0092_),
    .B1(_0625_));
 sg13g2_a22oi_1 _1565_ (.Y(_0626_),
    .B1(_0614_),
    .B2(_0609_),
    .A2(_0613_),
    .A1(net314));
 sg13g2_o21ai_1 _1566_ (.B1(_0610_),
    .Y(_0627_),
    .A1(_0600_),
    .A2(_0611_));
 sg13g2_and2_1 _1567_ (.A(\Ma[2] ),
    .B(net315),
    .X(_0628_));
 sg13g2_xor2_1 _1568_ (.B(net315),
    .A(\Ma[2] ),
    .X(_0629_));
 sg13g2_xnor2_1 _1569_ (.Y(_0630_),
    .A(_0627_),
    .B(_0629_));
 sg13g2_xor2_1 _1570_ (.B(_0630_),
    .A(\Ma[6] ),
    .X(_0631_));
 sg13g2_o21ai_1 _1571_ (.B1(_0615_),
    .Y(_0632_),
    .A1(_0626_),
    .A2(_0631_));
 sg13g2_a21o_1 _1572_ (.A2(_0631_),
    .A1(_0626_),
    .B1(_0632_),
    .X(_0633_));
 sg13g2_mux2_1 _1573_ (.A0(net314),
    .A1(\Ma[7] ),
    .S(net312),
    .X(_0634_));
 sg13g2_and2_1 _1574_ (.A(\Ma[2] ),
    .B(_0634_),
    .X(_0635_));
 sg13g2_xnor2_1 _1575_ (.Y(_0636_),
    .A(\Ma[2] ),
    .B(_0634_));
 sg13g2_inv_1 _1576_ (.Y(_0637_),
    .A(_0636_));
 sg13g2_o21ai_1 _1577_ (.B1(_0619_),
    .Y(_0638_),
    .A1(_0605_),
    .A2(_0620_));
 sg13g2_o21ai_1 _1578_ (.B1(net309),
    .Y(_0639_),
    .A1(_0637_),
    .A2(_0638_));
 sg13g2_a21oi_1 _1579_ (.A1(_0637_),
    .A2(_0638_),
    .Y(_0640_),
    .B1(_0639_));
 sg13g2_nor3_1 _1580_ (.A(net309),
    .B(_0304_),
    .C(_0630_),
    .Y(_0641_));
 sg13g2_nor3_1 _1581_ (.A(net286),
    .B(_0640_),
    .C(_0641_),
    .Y(_0642_));
 sg13g2_a22oi_1 _1582_ (.Y(_0093_),
    .B1(_0633_),
    .B2(_0642_),
    .A2(net286),
    .A1(_0320_));
 sg13g2_or2_1 _1583_ (.X(_0643_),
    .B(_0630_),
    .A(_0013_));
 sg13g2_o21ai_1 _1584_ (.B1(_0643_),
    .Y(_0644_),
    .A1(_0626_),
    .A2(_0631_));
 sg13g2_nor2_1 _1585_ (.A(net316),
    .B(net314),
    .Y(_0645_));
 sg13g2_nand2_1 _1586_ (.Y(_0646_),
    .A(net316),
    .B(net314));
 sg13g2_nor2b_1 _1587_ (.A(_0645_),
    .B_N(_0646_),
    .Y(_0647_));
 sg13g2_a21oi_1 _1588_ (.A1(_0627_),
    .A2(_0629_),
    .Y(_0648_),
    .B1(_0628_));
 sg13g2_xnor2_1 _1589_ (.Y(_0649_),
    .A(_0647_),
    .B(_0648_));
 sg13g2_xnor2_1 _1590_ (.Y(_0650_),
    .A(_0305_),
    .B(_0649_));
 sg13g2_xnor2_1 _1591_ (.Y(_0651_),
    .A(_0644_),
    .B(_0650_));
 sg13g2_a21o_1 _1592_ (.A2(_0638_),
    .A1(_0637_),
    .B1(_0635_),
    .X(_0652_));
 sg13g2_nor2_1 _1593_ (.A(net311),
    .B(net313),
    .Y(_0653_));
 sg13g2_o21ai_1 _1594_ (.B1(net316),
    .Y(_0654_),
    .A1(net311),
    .A2(net313));
 sg13g2_inv_1 _1595_ (.Y(_0655_),
    .A(_0654_));
 sg13g2_xnor2_1 _1596_ (.Y(_0656_),
    .A(net316),
    .B(_0653_));
 sg13g2_o21ai_1 _1597_ (.B1(net309),
    .Y(_0657_),
    .A1(_0652_),
    .A2(_0656_));
 sg13g2_a21oi_1 _1598_ (.A1(_0652_),
    .A2(_0656_),
    .Y(_0658_),
    .B1(_0657_));
 sg13g2_nor2_1 _1599_ (.A(net285),
    .B(_0658_),
    .Y(_0659_));
 sg13g2_nor2_1 _1600_ (.A(_0304_),
    .B(_0649_),
    .Y(_0660_));
 sg13g2_a21oi_1 _1601_ (.A1(_0304_),
    .A2(_0651_),
    .Y(_0661_),
    .B1(_0660_));
 sg13g2_nand2_1 _1602_ (.Y(_0662_),
    .A(net298),
    .B(_0661_));
 sg13g2_a22oi_1 _1603_ (.Y(_0094_),
    .B1(_0659_),
    .B2(_0662_),
    .A2(net285),
    .A1(_0322_));
 sg13g2_and2_1 _1604_ (.A(net315),
    .B(net313),
    .X(_0663_));
 sg13g2_or2_1 _1605_ (.X(_0664_),
    .B(net313),
    .A(net315));
 sg13g2_nand2b_1 _1606_ (.Y(_0665_),
    .B(_0664_),
    .A_N(_0663_));
 sg13g2_o21ai_1 _1607_ (.B1(_0646_),
    .Y(_0666_),
    .A1(_0645_),
    .A2(_0648_));
 sg13g2_xnor2_1 _1608_ (.Y(_0667_),
    .A(_0665_),
    .B(_0666_));
 sg13g2_a22oi_1 _1609_ (.Y(_0668_),
    .B1(_0650_),
    .B2(_0644_),
    .A2(_0649_),
    .A1(_0306_));
 sg13g2_nor2_1 _1610_ (.A(net310),
    .B(_0668_),
    .Y(_0669_));
 sg13g2_and2_1 _1611_ (.A(_0667_),
    .B(_0669_),
    .X(_0670_));
 sg13g2_nor2_1 _1612_ (.A(net309),
    .B(_0670_),
    .Y(_0671_));
 sg13g2_o21ai_1 _1613_ (.B1(_0671_),
    .Y(_0672_),
    .A1(_0667_),
    .A2(_0669_));
 sg13g2_a21oi_1 _1614_ (.A1(_0652_),
    .A2(_0656_),
    .Y(_0673_),
    .B1(_0655_));
 sg13g2_a21oi_2 _1615_ (.B1(_0623_),
    .Y(_0674_),
    .A2(_0305_),
    .A1(_0304_));
 sg13g2_xor2_1 _1616_ (.B(_0674_),
    .A(_0011_),
    .X(_0675_));
 sg13g2_or2_1 _1617_ (.X(_0676_),
    .B(_0675_),
    .A(_0673_));
 sg13g2_a21oi_1 _1618_ (.A1(_0673_),
    .A2(_0675_),
    .Y(_0677_),
    .B1(net298));
 sg13g2_a21oi_1 _1619_ (.A1(_0676_),
    .A2(_0677_),
    .Y(_0678_),
    .B1(net286));
 sg13g2_a22oi_1 _1620_ (.Y(_0095_),
    .B1(_0672_),
    .B2(_0678_),
    .A2(net287),
    .A1(_0324_));
 sg13g2_a21o_1 _1621_ (.A2(_0666_),
    .A1(_0664_),
    .B1(_0663_),
    .X(_0679_));
 sg13g2_and2_1 _1622_ (.A(net314),
    .B(\Ma[7] ),
    .X(_0680_));
 sg13g2_or2_1 _1623_ (.X(_0681_),
    .B(\Ma[7] ),
    .A(net314));
 sg13g2_nand2b_1 _1624_ (.Y(_0682_),
    .B(_0681_),
    .A_N(_0680_));
 sg13g2_xor2_1 _1625_ (.B(_0682_),
    .A(_0679_),
    .X(_0683_));
 sg13g2_xnor2_1 _1626_ (.Y(_0684_),
    .A(_0679_),
    .B(_0682_));
 sg13g2_nand2_1 _1627_ (.Y(_0685_),
    .A(net315),
    .B(_0674_));
 sg13g2_nand3_1 _1628_ (.B(_0676_),
    .C(_0685_),
    .A(_0012_),
    .Y(_0686_));
 sg13g2_a21o_1 _1629_ (.A2(_0685_),
    .A1(_0676_),
    .B1(_0012_),
    .X(_0687_));
 sg13g2_nand3_1 _1630_ (.B(_0686_),
    .C(_0687_),
    .A(net309),
    .Y(_0688_));
 sg13g2_nor2_1 _1631_ (.A(net308),
    .B(_0684_),
    .Y(_0689_));
 sg13g2_a221oi_1 _1632_ (.B2(_0670_),
    .C1(net286),
    .B1(_0689_),
    .A1(_0671_),
    .Y(_0690_),
    .A2(_0684_));
 sg13g2_a22oi_1 _1633_ (.Y(_0096_),
    .B1(_0688_),
    .B2(_0690_),
    .A2(net286),
    .A1(_0326_));
 sg13g2_xnor2_1 _1634_ (.Y(_0691_),
    .A(net310),
    .B(net313));
 sg13g2_a21oi_1 _1635_ (.A1(_0679_),
    .A2(_0681_),
    .Y(_0692_),
    .B1(_0680_));
 sg13g2_xnor2_1 _1636_ (.Y(_0693_),
    .A(_0691_),
    .B(_0692_));
 sg13g2_nor2_1 _1637_ (.A(net310),
    .B(_0667_),
    .Y(_0694_));
 sg13g2_a21oi_1 _1638_ (.A1(net308),
    .A2(_0684_),
    .Y(_0695_),
    .B1(_0694_));
 sg13g2_nand2_1 _1639_ (.Y(_0696_),
    .A(net310),
    .B(_0667_));
 sg13g2_a22oi_1 _1640_ (.Y(_0697_),
    .B1(_0696_),
    .B2(_0668_),
    .A2(_0683_),
    .A1(net298));
 sg13g2_a22oi_1 _1641_ (.Y(_0698_),
    .B1(_0695_),
    .B2(_0697_),
    .A2(_0684_),
    .A1(_0307_));
 sg13g2_or3_1 _1642_ (.A(net310),
    .B(_0693_),
    .C(_0698_),
    .X(_0699_));
 sg13g2_o21ai_1 _1643_ (.B1(_0693_),
    .Y(_0700_),
    .A1(net310),
    .A2(_0698_));
 sg13g2_nand3_1 _1644_ (.B(_0699_),
    .C(_0700_),
    .A(net298),
    .Y(_0701_));
 sg13g2_nand3_1 _1645_ (.B(net314),
    .C(_0674_),
    .A(net315),
    .Y(_0702_));
 sg13g2_inv_1 _1646_ (.Y(_0703_),
    .A(_0702_));
 sg13g2_nor3_1 _1647_ (.A(_0012_),
    .B(_0673_),
    .C(_0675_),
    .Y(_0704_));
 sg13g2_nor2_1 _1648_ (.A(net298),
    .B(net311),
    .Y(_0705_));
 sg13g2_xnor2_1 _1649_ (.Y(_0706_),
    .A(_0013_),
    .B(_0705_));
 sg13g2_o21ai_1 _1650_ (.B1(_0706_),
    .Y(_0707_),
    .A1(_0703_),
    .A2(_0704_));
 sg13g2_nor3_1 _1651_ (.A(_0703_),
    .B(_0704_),
    .C(_0706_),
    .Y(_0708_));
 sg13g2_nor2_1 _1652_ (.A(net298),
    .B(_0708_),
    .Y(_0709_));
 sg13g2_a21oi_1 _1653_ (.A1(_0707_),
    .A2(_0709_),
    .Y(_0710_),
    .B1(net285));
 sg13g2_a22oi_1 _1654_ (.Y(_0097_),
    .B1(_0701_),
    .B2(_0710_),
    .A2(net287),
    .A1(_0328_));
 sg13g2_o21ai_1 _1655_ (.B1(_0617_),
    .Y(_0711_),
    .A1(_0653_),
    .A2(_0692_));
 sg13g2_xor2_1 _1656_ (.B(\Ma[7] ),
    .A(net308),
    .X(_0712_));
 sg13g2_and2_1 _1657_ (.A(_0711_),
    .B(_0712_),
    .X(_0713_));
 sg13g2_xnor2_1 _1658_ (.Y(_0714_),
    .A(_0711_),
    .B(_0712_));
 sg13g2_a21oi_1 _1659_ (.A1(_0699_),
    .A2(_0714_),
    .Y(_0715_),
    .B1(net308));
 sg13g2_o21ai_1 _1660_ (.B1(_0715_),
    .Y(_0716_),
    .A1(_0699_),
    .A2(_0714_));
 sg13g2_nand2_1 _1661_ (.Y(_0717_),
    .A(net313),
    .B(_0705_));
 sg13g2_nand3_1 _1662_ (.B(_0707_),
    .C(_0717_),
    .A(_0014_),
    .Y(_0718_));
 sg13g2_a21oi_1 _1663_ (.A1(_0707_),
    .A2(_0717_),
    .Y(_0719_),
    .B1(_0014_));
 sg13g2_nor2_1 _1664_ (.A(net298),
    .B(_0719_),
    .Y(_0720_));
 sg13g2_a21oi_1 _1665_ (.A1(_0718_),
    .A2(_0720_),
    .Y(_0721_),
    .B1(net285));
 sg13g2_a22oi_1 _1666_ (.Y(_0098_),
    .B1(_0716_),
    .B2(_0721_),
    .A2(net285),
    .A1(_0330_));
 sg13g2_nor3_1 _1667_ (.A(_0693_),
    .B(_0698_),
    .C(_0714_),
    .Y(_0722_));
 sg13g2_or3_1 _1668_ (.A(net310),
    .B(_0713_),
    .C(_0722_),
    .X(_0723_));
 sg13g2_a21oi_1 _1669_ (.A1(net310),
    .A2(_0713_),
    .Y(_0724_),
    .B1(net308));
 sg13g2_nand2b_1 _1670_ (.Y(_0725_),
    .B(_0015_),
    .A_N(_0719_));
 sg13g2_a21o_1 _1671_ (.A2(_0015_),
    .A1(net308),
    .B1(_0720_),
    .X(_0726_));
 sg13g2_a21oi_1 _1672_ (.A1(net308),
    .A2(net431),
    .Y(_0727_),
    .B1(_0720_));
 sg13g2_a221oi_1 _1673_ (.B2(_0726_),
    .C1(net285),
    .B1(_0725_),
    .A1(_0723_),
    .Y(_0728_),
    .A2(_0724_));
 sg13g2_a21oi_1 _1674_ (.A1(_0332_),
    .A2(net282),
    .Y(_0099_),
    .B1(_0728_));
 sg13g2_a21oi_1 _1675_ (.A1(_0623_),
    .A2(_0713_),
    .Y(_0729_),
    .B1(net285));
 sg13g2_a22oi_1 _1676_ (.Y(_0100_),
    .B1(net432),
    .B2(_0729_),
    .A2(net285),
    .A1(_0334_));
 sg13g2_nand2_1 _1677_ (.Y(_0730_),
    .A(\Mb[0] ),
    .B(\Mb[2] ));
 sg13g2_xor2_1 _1678_ (.B(\Mb[2] ),
    .A(\Mb[0] ),
    .X(_0731_));
 sg13g2_nor2_1 _1679_ (.A(_0017_),
    .B(net302),
    .Y(_0732_));
 sg13g2_xor2_1 _1680_ (.B(_0732_),
    .A(_0731_),
    .X(_0733_));
 sg13g2_mux2_1 _1681_ (.A0(net307),
    .A1(\Mb[5] ),
    .S(net302),
    .X(_0734_));
 sg13g2_nand2_1 _1682_ (.Y(_0735_),
    .A(\Mb[0] ),
    .B(_0734_));
 sg13g2_o21ai_1 _1683_ (.B1(net300),
    .Y(_0736_),
    .A1(\Mb[0] ),
    .A2(_0734_));
 sg13g2_inv_1 _1684_ (.Y(_0737_),
    .A(_0736_));
 sg13g2_a221oi_1 _1685_ (.B2(_0737_),
    .C1(net284),
    .B1(_0735_),
    .A1(_0308_),
    .Y(_0738_),
    .A2(_0733_));
 sg13g2_a21oi_1 _1686_ (.A1(_0317_),
    .A2(net283),
    .Y(_0101_),
    .B1(_0738_));
 sg13g2_and2_1 _1687_ (.A(net306),
    .B(_0731_),
    .X(_0739_));
 sg13g2_nand2_1 _1688_ (.Y(_0740_),
    .A(\Mb[3] ),
    .B(\Mb[1] ));
 sg13g2_nor2_1 _1689_ (.A(net307),
    .B(\Mb[1] ),
    .Y(_0741_));
 sg13g2_xor2_1 _1690_ (.B(\Mb[1] ),
    .A(net307),
    .X(_0742_));
 sg13g2_xnor2_1 _1691_ (.Y(_0743_),
    .A(_0730_),
    .B(_0742_));
 sg13g2_xnor2_1 _1692_ (.Y(_0744_),
    .A(_0018_),
    .B(_0743_));
 sg13g2_nor2_1 _1693_ (.A(net300),
    .B(net302),
    .Y(_0745_));
 sg13g2_xnor2_1 _1694_ (.Y(_0746_),
    .A(_0739_),
    .B(_0744_));
 sg13g2_nor3_1 _1695_ (.A(net300),
    .B(net303),
    .C(_0746_),
    .Y(_0747_));
 sg13g2_nand2_1 _1696_ (.Y(_0748_),
    .A(net301),
    .B(net304));
 sg13g2_mux2_1 _1697_ (.A0(\Mb[4] ),
    .A1(\Mb[6] ),
    .S(net302),
    .X(_0749_));
 sg13g2_nand2_1 _1698_ (.Y(_0750_),
    .A(\Mb[1] ),
    .B(_0749_));
 sg13g2_xnor2_1 _1699_ (.Y(_0751_),
    .A(\Mb[1] ),
    .B(_0749_));
 sg13g2_o21ai_1 _1700_ (.B1(net300),
    .Y(_0752_),
    .A1(_0735_),
    .A2(_0751_));
 sg13g2_a21oi_1 _1701_ (.A1(_0735_),
    .A2(_0751_),
    .Y(_0753_),
    .B1(_0752_));
 sg13g2_nor2_2 _1702_ (.A(net300),
    .B(_0309_),
    .Y(_0754_));
 sg13g2_nand2_1 _1703_ (.Y(_0755_),
    .A(_0743_),
    .B(_0754_));
 sg13g2_nor3_1 _1704_ (.A(net283),
    .B(_0747_),
    .C(_0753_),
    .Y(_0756_));
 sg13g2_a22oi_1 _1705_ (.Y(_0102_),
    .B1(_0755_),
    .B2(_0756_),
    .A2(net287),
    .A1(_0315_));
 sg13g2_a22oi_1 _1706_ (.Y(_0757_),
    .B1(_0744_),
    .B2(_0739_),
    .A2(_0743_),
    .A1(net305));
 sg13g2_o21ai_1 _1707_ (.B1(_0740_),
    .Y(_0758_),
    .A1(_0730_),
    .A2(_0741_));
 sg13g2_and2_1 _1708_ (.A(\Mb[2] ),
    .B(net306),
    .X(_0759_));
 sg13g2_xor2_1 _1709_ (.B(net306),
    .A(\Mb[2] ),
    .X(_0760_));
 sg13g2_xnor2_1 _1710_ (.Y(_0761_),
    .A(_0758_),
    .B(_0760_));
 sg13g2_xor2_1 _1711_ (.B(_0761_),
    .A(\Mb[6] ),
    .X(_0762_));
 sg13g2_o21ai_1 _1712_ (.B1(_0745_),
    .Y(_0763_),
    .A1(_0757_),
    .A2(_0762_));
 sg13g2_a21o_1 _1713_ (.A2(_0762_),
    .A1(_0757_),
    .B1(_0763_),
    .X(_0764_));
 sg13g2_mux2_1 _1714_ (.A0(net305),
    .A1(\Mb[7] ),
    .S(net303),
    .X(_0765_));
 sg13g2_and2_1 _1715_ (.A(\Mb[2] ),
    .B(_0765_),
    .X(_0766_));
 sg13g2_xnor2_1 _1716_ (.Y(_0767_),
    .A(\Mb[2] ),
    .B(_0765_));
 sg13g2_inv_1 _1717_ (.Y(_0768_),
    .A(_0767_));
 sg13g2_o21ai_1 _1718_ (.B1(_0750_),
    .Y(_0769_),
    .A1(_0735_),
    .A2(_0751_));
 sg13g2_o21ai_1 _1719_ (.B1(net300),
    .Y(_0770_),
    .A1(_0768_),
    .A2(_0769_));
 sg13g2_a21oi_1 _1720_ (.A1(_0768_),
    .A2(_0769_),
    .Y(_0771_),
    .B1(_0770_));
 sg13g2_nor3_1 _1721_ (.A(net300),
    .B(_0309_),
    .C(_0761_),
    .Y(_0772_));
 sg13g2_nor3_1 _1722_ (.A(net284),
    .B(_0771_),
    .C(_0772_),
    .Y(_0773_));
 sg13g2_a22oi_1 _1723_ (.Y(_0103_),
    .B1(_0764_),
    .B2(_0773_),
    .A2(net287),
    .A1(_0319_));
 sg13g2_or2_1 _1724_ (.X(_0774_),
    .B(_0761_),
    .A(_0019_));
 sg13g2_o21ai_1 _1725_ (.B1(_0774_),
    .Y(_0775_),
    .A1(_0757_),
    .A2(_0762_));
 sg13g2_nor2_1 _1726_ (.A(net307),
    .B(net305),
    .Y(_0776_));
 sg13g2_nand2_1 _1727_ (.Y(_0777_),
    .A(net307),
    .B(net305));
 sg13g2_nor2b_1 _1728_ (.A(_0776_),
    .B_N(_0777_),
    .Y(_0778_));
 sg13g2_a21oi_2 _1729_ (.B1(_0759_),
    .Y(_0779_),
    .A2(_0760_),
    .A1(_0758_));
 sg13g2_xnor2_1 _1730_ (.Y(_0780_),
    .A(_0778_),
    .B(_0779_));
 sg13g2_xnor2_1 _1731_ (.Y(_0781_),
    .A(_0310_),
    .B(_0780_));
 sg13g2_nand2_1 _1732_ (.Y(_0782_),
    .A(_0775_),
    .B(_0781_));
 sg13g2_nor2_1 _1733_ (.A(_0775_),
    .B(_0781_),
    .Y(_0783_));
 sg13g2_nor2b_1 _1734_ (.A(_0783_),
    .B_N(_0745_),
    .Y(_0784_));
 sg13g2_a21o_1 _1735_ (.A2(_0769_),
    .A1(_0768_),
    .B1(_0766_),
    .X(_0785_));
 sg13g2_nor2_1 _1736_ (.A(net303),
    .B(net304),
    .Y(_0786_));
 sg13g2_o21ai_1 _1737_ (.B1(net307),
    .Y(_0787_),
    .A1(net302),
    .A2(net304));
 sg13g2_inv_1 _1738_ (.Y(_0788_),
    .A(_0787_));
 sg13g2_xnor2_1 _1739_ (.Y(_0789_),
    .A(net307),
    .B(_0786_));
 sg13g2_nor2_1 _1740_ (.A(_0785_),
    .B(_0789_),
    .Y(_0790_));
 sg13g2_a21o_1 _1741_ (.A2(_0789_),
    .A1(_0785_),
    .B1(net297),
    .X(_0791_));
 sg13g2_o21ai_1 _1742_ (.B1(_0002_),
    .Y(_0792_),
    .A1(_0790_),
    .A2(_0791_));
 sg13g2_a221oi_1 _1743_ (.B2(_0784_),
    .C1(_0792_),
    .B1(_0782_),
    .A1(_0754_),
    .Y(_0793_),
    .A2(_0780_));
 sg13g2_a21oi_1 _1744_ (.A1(_0321_),
    .A2(net283),
    .Y(_0104_),
    .B1(_0793_));
 sg13g2_and2_1 _1745_ (.A(net306),
    .B(net304),
    .X(_0794_));
 sg13g2_or2_1 _1746_ (.X(_0795_),
    .B(net304),
    .A(net306));
 sg13g2_nand2b_1 _1747_ (.Y(_0796_),
    .B(_0795_),
    .A_N(_0794_));
 sg13g2_o21ai_1 _1748_ (.B1(_0777_),
    .Y(_0797_),
    .A1(_0776_),
    .A2(_0779_));
 sg13g2_xnor2_1 _1749_ (.Y(_0798_),
    .A(_0796_),
    .B(_0797_));
 sg13g2_xor2_1 _1750_ (.B(_0797_),
    .A(_0796_),
    .X(_0799_));
 sg13g2_nor2b_1 _1751_ (.A(_0020_),
    .B_N(_0780_),
    .Y(_0800_));
 sg13g2_a21oi_1 _1752_ (.A1(_0775_),
    .A2(_0781_),
    .Y(_0801_),
    .B1(_0800_));
 sg13g2_o21ai_1 _1753_ (.B1(_0799_),
    .Y(_0802_),
    .A1(net302),
    .A2(_0801_));
 sg13g2_nor3_1 _1754_ (.A(net301),
    .B(_0799_),
    .C(_0801_),
    .Y(_0803_));
 sg13g2_nor2_1 _1755_ (.A(net299),
    .B(_0803_),
    .Y(_0804_));
 sg13g2_a21oi_1 _1756_ (.A1(_0785_),
    .A2(_0789_),
    .Y(_0805_),
    .B1(_0788_));
 sg13g2_a21oi_2 _1757_ (.B1(_0754_),
    .Y(_0806_),
    .A2(_0310_),
    .A1(_0309_));
 sg13g2_xor2_1 _1758_ (.B(_0806_),
    .A(_0017_),
    .X(_0807_));
 sg13g2_or2_1 _1759_ (.X(_0808_),
    .B(_0807_),
    .A(_0805_));
 sg13g2_a21oi_1 _1760_ (.A1(_0805_),
    .A2(_0807_),
    .Y(_0809_),
    .B1(net297));
 sg13g2_nand2_1 _1761_ (.Y(_0810_),
    .A(_0808_),
    .B(_0809_));
 sg13g2_a21oi_1 _1762_ (.A1(_0802_),
    .A2(_0804_),
    .Y(_0811_),
    .B1(net283));
 sg13g2_a22oi_1 _1763_ (.Y(_0105_),
    .B1(_0810_),
    .B2(_0811_),
    .A2(net283),
    .A1(_0323_));
 sg13g2_a21o_1 _1764_ (.A2(_0797_),
    .A1(_0795_),
    .B1(_0794_),
    .X(_0812_));
 sg13g2_and2_1 _1765_ (.A(net305),
    .B(\Mb[7] ),
    .X(_0813_));
 sg13g2_or2_1 _1766_ (.X(_0814_),
    .B(\Mb[7] ),
    .A(net305));
 sg13g2_nand2b_1 _1767_ (.Y(_0815_),
    .B(_0814_),
    .A_N(_0813_));
 sg13g2_xnor2_1 _1768_ (.Y(_0816_),
    .A(_0812_),
    .B(_0815_));
 sg13g2_nor2_1 _1769_ (.A(net299),
    .B(_0816_),
    .Y(_0817_));
 sg13g2_nand2_1 _1770_ (.Y(_0818_),
    .A(net306),
    .B(_0806_));
 sg13g2_a21oi_1 _1771_ (.A1(_0808_),
    .A2(_0818_),
    .Y(_0819_),
    .B1(_0018_));
 sg13g2_nand3_1 _1772_ (.B(_0808_),
    .C(_0818_),
    .A(_0018_),
    .Y(_0820_));
 sg13g2_nor2_1 _1773_ (.A(_0308_),
    .B(_0819_),
    .Y(_0821_));
 sg13g2_a21oi_1 _1774_ (.A1(_0820_),
    .A2(_0821_),
    .Y(_0822_),
    .B1(net283));
 sg13g2_a22oi_1 _1775_ (.Y(_0823_),
    .B1(_0817_),
    .B2(_0803_),
    .A2(_0816_),
    .A1(_0804_));
 sg13g2_a22oi_1 _1776_ (.Y(_0106_),
    .B1(_0822_),
    .B2(_0823_),
    .A2(net284),
    .A1(_0325_));
 sg13g2_xnor2_1 _1777_ (.Y(_0824_),
    .A(net301),
    .B(net304));
 sg13g2_a21oi_1 _1778_ (.A1(_0812_),
    .A2(_0814_),
    .Y(_0825_),
    .B1(_0813_));
 sg13g2_xnor2_1 _1779_ (.Y(_0826_),
    .A(_0824_),
    .B(_0825_));
 sg13g2_a221oi_1 _1780_ (.B2(net302),
    .C1(_0800_),
    .B1(_0798_),
    .A1(_0775_),
    .Y(_0827_),
    .A2(_0781_));
 sg13g2_a21oi_1 _1781_ (.A1(_0309_),
    .A2(_0799_),
    .Y(_0828_),
    .B1(_0827_));
 sg13g2_xnor2_1 _1782_ (.Y(_0829_),
    .A(net297),
    .B(_0816_));
 sg13g2_a22oi_1 _1783_ (.Y(_0830_),
    .B1(_0828_),
    .B2(_0829_),
    .A2(_0816_),
    .A1(_0311_));
 sg13g2_or3_1 _1784_ (.A(net301),
    .B(_0826_),
    .C(_0830_),
    .X(_0831_));
 sg13g2_o21ai_1 _1785_ (.B1(_0826_),
    .Y(_0832_),
    .A1(net301),
    .A2(_0830_));
 sg13g2_nand3_1 _1786_ (.B(_0831_),
    .C(_0832_),
    .A(net297),
    .Y(_0833_));
 sg13g2_nand3_1 _1787_ (.B(net305),
    .C(_0806_),
    .A(net306),
    .Y(_0834_));
 sg13g2_inv_1 _1788_ (.Y(_0835_),
    .A(_0834_));
 sg13g2_nor3_1 _1789_ (.A(_0018_),
    .B(_0805_),
    .C(_0807_),
    .Y(_0836_));
 sg13g2_nor2_1 _1790_ (.A(net297),
    .B(net301),
    .Y(_0837_));
 sg13g2_xnor2_1 _1791_ (.Y(_0838_),
    .A(_0019_),
    .B(_0837_));
 sg13g2_o21ai_1 _1792_ (.B1(_0838_),
    .Y(_0839_),
    .A1(_0835_),
    .A2(_0836_));
 sg13g2_nor3_1 _1793_ (.A(_0835_),
    .B(_0836_),
    .C(_0838_),
    .Y(_0840_));
 sg13g2_nor2_1 _1794_ (.A(net297),
    .B(_0840_),
    .Y(_0841_));
 sg13g2_a21oi_1 _1795_ (.A1(_0839_),
    .A2(_0841_),
    .Y(_0842_),
    .B1(net282));
 sg13g2_a22oi_1 _1796_ (.Y(_0107_),
    .B1(_0833_),
    .B2(_0842_),
    .A2(net282),
    .A1(_0327_));
 sg13g2_o21ai_1 _1797_ (.B1(_0748_),
    .Y(_0843_),
    .A1(_0786_),
    .A2(_0825_));
 sg13g2_xor2_1 _1798_ (.B(\Mb[7] ),
    .A(net299),
    .X(_0844_));
 sg13g2_and2_1 _1799_ (.A(_0843_),
    .B(_0844_),
    .X(_0845_));
 sg13g2_xnor2_1 _1800_ (.Y(_0846_),
    .A(_0843_),
    .B(_0844_));
 sg13g2_a21oi_1 _1801_ (.A1(_0831_),
    .A2(_0846_),
    .Y(_0847_),
    .B1(net299));
 sg13g2_o21ai_1 _1802_ (.B1(_0847_),
    .Y(_0161_),
    .A1(_0831_),
    .A2(_0846_));
 sg13g2_nand2_1 _1803_ (.Y(_0162_),
    .A(net304),
    .B(_0837_));
 sg13g2_nand3_1 _1804_ (.B(_0839_),
    .C(_0162_),
    .A(_0020_),
    .Y(_0163_));
 sg13g2_a21oi_1 _1805_ (.A1(_0839_),
    .A2(_0162_),
    .Y(_0164_),
    .B1(_0020_));
 sg13g2_nor2_1 _1806_ (.A(net297),
    .B(_0164_),
    .Y(_0165_));
 sg13g2_a21oi_1 _1807_ (.A1(_0163_),
    .A2(_0165_),
    .Y(_0166_),
    .B1(net282));
 sg13g2_a22oi_1 _1808_ (.Y(_0108_),
    .B1(_0161_),
    .B2(_0166_),
    .A2(net282),
    .A1(_0329_));
 sg13g2_nor3_1 _1809_ (.A(_0826_),
    .B(_0830_),
    .C(_0846_),
    .Y(_0167_));
 sg13g2_or3_1 _1810_ (.A(net301),
    .B(_0845_),
    .C(_0167_),
    .X(_0168_));
 sg13g2_a21oi_1 _1811_ (.A1(net301),
    .A2(_0845_),
    .Y(_0169_),
    .B1(net299));
 sg13g2_nand2b_1 _1812_ (.Y(_0170_),
    .B(_0021_),
    .A_N(_0164_));
 sg13g2_a21o_1 _1813_ (.A2(_0021_),
    .A1(net299),
    .B1(_0165_),
    .X(_0171_));
 sg13g2_a21oi_1 _1814_ (.A1(net299),
    .A2(_0021_),
    .Y(_0172_),
    .B1(_0165_));
 sg13g2_a221oi_1 _1815_ (.B2(_0171_),
    .C1(net282),
    .B1(_0170_),
    .A1(_0168_),
    .Y(_0173_),
    .A2(_0169_));
 sg13g2_a21oi_1 _1816_ (.A1(_0331_),
    .A2(net282),
    .Y(_0109_),
    .B1(_0173_));
 sg13g2_a21oi_1 _1817_ (.A1(_0754_),
    .A2(_0845_),
    .Y(_0174_),
    .B1(net283));
 sg13g2_a22oi_1 _1818_ (.Y(_0110_),
    .B1(_0172_),
    .B2(_0174_),
    .A2(net282),
    .A1(_0333_));
 sg13g2_nand2_1 _1819_ (.Y(_0175_),
    .A(\M1bout[0] ),
    .B(\M1aout[0] ));
 sg13g2_xnor2_1 _1820_ (.Y(_0176_),
    .A(\M1bout[0] ),
    .B(\M1aout[0] ));
 sg13g2_nand2_1 _1821_ (.Y(_0177_),
    .A(net231),
    .B(net277));
 sg13g2_o21ai_1 _1822_ (.B1(_0177_),
    .Y(_0111_),
    .A1(net277),
    .A2(_0176_));
 sg13g2_nand2_1 _1823_ (.Y(_0178_),
    .A(net414),
    .B(net379));
 sg13g2_nor2_1 _1824_ (.A(\M1bout[1] ),
    .B(\M1aout[1] ),
    .Y(_0179_));
 sg13g2_nand2_1 _1825_ (.Y(_0180_),
    .A(_0315_),
    .B(_0316_));
 sg13g2_a22oi_1 _1826_ (.Y(_0181_),
    .B1(_0178_),
    .B2(_0180_),
    .A2(net429),
    .A1(net427));
 sg13g2_nand4_1 _1827_ (.B(net429),
    .C(_0178_),
    .A(net427),
    .Y(_0182_),
    .D(_0180_));
 sg13g2_nor2_1 _1828_ (.A(net278),
    .B(_0181_),
    .Y(_0183_));
 sg13g2_a22oi_1 _1829_ (.Y(_0184_),
    .B1(_0182_),
    .B2(_0183_),
    .A2(net278),
    .A1(net441));
 sg13g2_inv_1 _1830_ (.Y(_0112_),
    .A(net442));
 sg13g2_nor2_1 _1831_ (.A(_0319_),
    .B(_0320_),
    .Y(_0185_));
 sg13g2_nand2_1 _1832_ (.Y(_0186_),
    .A(_0319_),
    .B(_0320_));
 sg13g2_nand2b_1 _1833_ (.Y(_0187_),
    .B(_0186_),
    .A_N(_0185_));
 sg13g2_o21ai_1 _1834_ (.B1(_0178_),
    .Y(_0188_),
    .A1(_0175_),
    .A2(_0179_));
 sg13g2_nor2_1 _1835_ (.A(net356),
    .B(_0005_),
    .Y(_0189_));
 sg13g2_xor2_1 _1836_ (.B(_0188_),
    .A(_0187_),
    .X(_0190_));
 sg13g2_a21oi_1 _1837_ (.A1(_0005_),
    .A2(_0190_),
    .Y(_0113_),
    .B1(_0189_));
 sg13g2_nand2_1 _1838_ (.Y(_0191_),
    .A(net329),
    .B(net277));
 sg13g2_nand2_1 _1839_ (.Y(_0192_),
    .A(\M1bout[3] ),
    .B(\M1aout[3] ));
 sg13g2_xnor2_1 _1840_ (.Y(_0193_),
    .A(\M1bout[3] ),
    .B(\M1aout[3] ));
 sg13g2_a21oi_2 _1841_ (.B1(_0185_),
    .Y(_0194_),
    .A2(_0188_),
    .A1(_0186_));
 sg13g2_xnor2_1 _1842_ (.Y(_0195_),
    .A(_0193_),
    .B(_0194_));
 sg13g2_o21ai_1 _1843_ (.B1(_0191_),
    .Y(_0114_),
    .A1(net277),
    .A2(_0195_));
 sg13g2_nor2_1 _1844_ (.A(_0323_),
    .B(_0324_),
    .Y(_0196_));
 sg13g2_xor2_1 _1845_ (.B(\M1aout[4] ),
    .A(\M1bout[4] ),
    .X(_0197_));
 sg13g2_o21ai_1 _1846_ (.B1(_0192_),
    .Y(_0198_),
    .A1(_0193_),
    .A2(_0194_));
 sg13g2_xnor2_1 _1847_ (.Y(_0199_),
    .A(_0197_),
    .B(_0198_));
 sg13g2_nand2_1 _1848_ (.Y(_0200_),
    .A(net328),
    .B(net276));
 sg13g2_o21ai_1 _1849_ (.B1(_0200_),
    .Y(_0115_),
    .A1(net276),
    .A2(_0199_));
 sg13g2_a21oi_1 _1850_ (.A1(_0197_),
    .A2(_0198_),
    .Y(_0201_),
    .B1(_0196_));
 sg13g2_nor2_1 _1851_ (.A(\M1bout[5] ),
    .B(\M1aout[5] ),
    .Y(_0202_));
 sg13g2_nand2_1 _1852_ (.Y(_0203_),
    .A(\M1bout[5] ),
    .B(\M1aout[5] ));
 sg13g2_nor2b_1 _1853_ (.A(_0202_),
    .B_N(_0203_),
    .Y(_0204_));
 sg13g2_xnor2_1 _1854_ (.Y(_0205_),
    .A(_0201_),
    .B(_0204_));
 sg13g2_mux2_1 _1855_ (.A0(net327),
    .A1(_0205_),
    .S(_0005_),
    .X(_0116_));
 sg13g2_nor2_1 _1856_ (.A(_0327_),
    .B(_0328_),
    .Y(_0206_));
 sg13g2_xor2_1 _1857_ (.B(\M1aout[6] ),
    .A(\M1bout[6] ),
    .X(_0207_));
 sg13g2_o21ai_1 _1858_ (.B1(_0203_),
    .Y(_0208_),
    .A1(_0201_),
    .A2(_0202_));
 sg13g2_xnor2_1 _1859_ (.Y(_0209_),
    .A(_0207_),
    .B(_0208_));
 sg13g2_nand2_1 _1860_ (.Y(_0210_),
    .A(net324),
    .B(net276));
 sg13g2_o21ai_1 _1861_ (.B1(_0210_),
    .Y(_0117_),
    .A1(net276),
    .A2(_0209_));
 sg13g2_nor2_1 _1862_ (.A(_0329_),
    .B(_0330_),
    .Y(_0211_));
 sg13g2_nand2_1 _1863_ (.Y(_0212_),
    .A(_0329_),
    .B(_0330_));
 sg13g2_nand2b_1 _1864_ (.Y(_0213_),
    .B(_0212_),
    .A_N(_0211_));
 sg13g2_a21o_1 _1865_ (.A2(_0208_),
    .A1(_0207_),
    .B1(_0206_),
    .X(_0214_));
 sg13g2_xnor2_1 _1866_ (.Y(_0215_),
    .A(_0213_),
    .B(_0214_));
 sg13g2_nor2_1 _1867_ (.A(net276),
    .B(_0215_),
    .Y(_0216_));
 sg13g2_a21oi_1 _1868_ (.A1(_0314_),
    .A2(net276),
    .Y(_0118_),
    .B1(_0216_));
 sg13g2_xor2_1 _1869_ (.B(net388),
    .A(net376),
    .X(_0217_));
 sg13g2_a21o_1 _1870_ (.A2(_0214_),
    .A1(_0212_),
    .B1(_0211_),
    .X(_0218_));
 sg13g2_nand2_1 _1871_ (.Y(_0219_),
    .A(_0217_),
    .B(_0218_));
 sg13g2_xnor2_1 _1872_ (.Y(_0220_),
    .A(_0217_),
    .B(_0218_));
 sg13g2_nand2_1 _1873_ (.Y(_0221_),
    .A(net320),
    .B(net276));
 sg13g2_o21ai_1 _1874_ (.B1(_0221_),
    .Y(_0119_),
    .A1(net276),
    .A2(_0220_));
 sg13g2_xnor2_1 _1875_ (.Y(_0222_),
    .A(\M1bout[9] ),
    .B(\M1aout[9] ));
 sg13g2_o21ai_1 _1876_ (.B1(_0219_),
    .Y(_0223_),
    .A1(_0331_),
    .A2(_0332_));
 sg13g2_xnor2_1 _1877_ (.Y(_0224_),
    .A(_0222_),
    .B(_0223_));
 sg13g2_mux2_1 _1878_ (.A0(net319),
    .A1(_0224_),
    .S(_0005_),
    .X(_0120_));
 sg13g2_nand2_1 _1879_ (.Y(_0225_),
    .A(net253),
    .B(net278));
 sg13g2_a21oi_1 _1880_ (.A1(\M1bout[9] ),
    .A2(\M1aout[9] ),
    .Y(_0226_),
    .B1(_0223_));
 sg13g2_o21ai_1 _1881_ (.B1(_0005_),
    .Y(_0227_),
    .A1(\M1bout[9] ),
    .A2(\M1aout[9] ));
 sg13g2_o21ai_1 _1882_ (.B1(net254),
    .Y(_0121_),
    .A1(_0226_),
    .A2(_0227_));
 sg13g2_nor2_2 _1883_ (.A(Ce),
    .B(\Ea[0] ),
    .Y(_0228_));
 sg13g2_and2_1 _1884_ (.A(Ce),
    .B(\Ea[0] ),
    .X(_0229_));
 sg13g2_nor3_1 _1885_ (.A(net204),
    .B(_0228_),
    .C(_0229_),
    .Y(_0230_));
 sg13g2_o21ai_1 _1886_ (.B1(net204),
    .Y(_0231_),
    .A1(_0228_),
    .A2(_0229_));
 sg13g2_nor2_1 _1887_ (.A(_0353_),
    .B(_0230_),
    .Y(_0232_));
 sg13g2_a22oi_1 _1888_ (.Y(_0233_),
    .B1(_0231_),
    .B2(_0232_),
    .A2(net281),
    .A1(net188));
 sg13g2_inv_1 _1889_ (.Y(_0122_),
    .A(_0233_));
 sg13g2_nor2_1 _1890_ (.A(net183),
    .B(net275),
    .Y(_0234_));
 sg13g2_nand2_1 _1891_ (.Y(_0235_),
    .A(\Eb[1] ),
    .B(\Ea[1] ));
 sg13g2_xor2_1 _1892_ (.B(\Ea[1] ),
    .A(\Eb[1] ),
    .X(_0236_));
 sg13g2_nand2b_1 _1893_ (.Y(_0237_),
    .B(_0236_),
    .A_N(_0228_));
 sg13g2_xnor2_1 _1894_ (.Y(_0238_),
    .A(_0228_),
    .B(_0236_));
 sg13g2_nand2b_1 _1895_ (.Y(_0239_),
    .B(_0238_),
    .A_N(_0231_));
 sg13g2_xor2_1 _1896_ (.B(_0238_),
    .A(_0231_),
    .X(_0240_));
 sg13g2_a21oi_1 _1897_ (.A1(_0000_),
    .A2(_0240_),
    .Y(_0123_),
    .B1(_0234_));
 sg13g2_nor2_1 _1898_ (.A(net214),
    .B(net275),
    .Y(_0241_));
 sg13g2_and2_1 _1899_ (.A(\Eb[2] ),
    .B(\Ea[2] ),
    .X(_0242_));
 sg13g2_xor2_1 _1900_ (.B(\Ea[2] ),
    .A(\Eb[2] ),
    .X(_0243_));
 sg13g2_nand2b_1 _1901_ (.Y(_0244_),
    .B(_0243_),
    .A_N(_0235_));
 sg13g2_xnor2_1 _1902_ (.Y(_0245_),
    .A(_0235_),
    .B(_0243_));
 sg13g2_nand2_1 _1903_ (.Y(_0246_),
    .A(_0237_),
    .B(_0239_));
 sg13g2_nand2_1 _1904_ (.Y(_0247_),
    .A(_0245_),
    .B(_0246_));
 sg13g2_xnor2_1 _1905_ (.Y(_0248_),
    .A(_0245_),
    .B(_0246_));
 sg13g2_a21oi_1 _1906_ (.A1(net275),
    .A2(_0248_),
    .Y(_0124_),
    .B1(_0241_));
 sg13g2_nand2_1 _1907_ (.Y(_0249_),
    .A(\Eb[3] ),
    .B(\Ea[3] ));
 sg13g2_xor2_1 _1908_ (.B(\Ea[3] ),
    .A(\Eb[3] ),
    .X(_0250_));
 sg13g2_xnor2_1 _1909_ (.Y(_0251_),
    .A(_0242_),
    .B(_0250_));
 sg13g2_a21oi_2 _1910_ (.B1(_0251_),
    .Y(_0252_),
    .A2(_0247_),
    .A1(_0244_));
 sg13g2_nand3_1 _1911_ (.B(_0247_),
    .C(_0251_),
    .A(_0244_),
    .Y(_0253_));
 sg13g2_nand2_1 _1912_ (.Y(_0254_),
    .A(net275),
    .B(_0253_));
 sg13g2_nand2_1 _1913_ (.Y(_0255_),
    .A(net185),
    .B(net281));
 sg13g2_o21ai_1 _1914_ (.B1(_0255_),
    .Y(_0125_),
    .A1(_0252_),
    .A2(_0254_));
 sg13g2_nor2_1 _1915_ (.A(net190),
    .B(net275),
    .Y(_0256_));
 sg13g2_a21oi_1 _1916_ (.A1(_0242_),
    .A2(_0250_),
    .Y(_0257_),
    .B1(_0252_));
 sg13g2_xor2_1 _1917_ (.B(\Ea[4] ),
    .A(\Eb[4] ),
    .X(_0258_));
 sg13g2_xnor2_1 _1918_ (.Y(_0259_),
    .A(_0249_),
    .B(_0258_));
 sg13g2_xnor2_1 _1919_ (.Y(_0260_),
    .A(_0257_),
    .B(_0259_));
 sg13g2_a21oi_1 _1920_ (.A1(net275),
    .A2(_0260_),
    .Y(_0126_),
    .B1(_0256_));
 sg13g2_mux2_1 _1921_ (.A0(net246),
    .A1(net372),
    .S(net290),
    .X(_0127_));
 sg13g2_mux2_1 _1922_ (.A0(net194),
    .A1(net216),
    .S(net293),
    .X(_0128_));
 sg13g2_mux2_1 _1923_ (.A0(net208),
    .A1(net262),
    .S(net293),
    .X(_0129_));
 sg13g2_mux2_1 _1924_ (.A0(net195),
    .A1(\Ea[3] ),
    .S(net293),
    .X(_0130_));
 sg13g2_mux2_1 _1925_ (.A0(net222),
    .A1(net233),
    .S(net293),
    .X(_0131_));
 sg13g2_mux2_1 _1926_ (.A0(net203),
    .A1(net204),
    .S(net290),
    .X(_0132_));
 sg13g2_mux2_1 _1927_ (.A0(net199),
    .A1(net221),
    .S(net293),
    .X(_0133_));
 sg13g2_mux2_1 _1928_ (.A0(net217),
    .A1(net245),
    .S(net293),
    .X(_0134_));
 sg13g2_mux2_1 _1929_ (.A0(net226),
    .A1(net200),
    .S(net293),
    .X(_0135_));
 sg13g2_mux2_1 _1930_ (.A0(net360),
    .A1(\Eb[4] ),
    .S(net294),
    .X(_0136_));
 sg13g2_xor2_1 _1931_ (.B(net227),
    .A(net223),
    .X(_0261_));
 sg13g2_nor2_1 _1932_ (.A(net284),
    .B(_0261_),
    .Y(_0262_));
 sg13g2_a21oi_1 _1933_ (.A1(_0269_),
    .A2(net284),
    .Y(_0137_),
    .B1(_0262_));
 sg13g2_mux2_1 _1934_ (.A0(net197),
    .A1(Sa),
    .S(net293),
    .X(_0138_));
 sg13g2_mux2_1 _1935_ (.A0(net187),
    .A1(net223),
    .S(net290),
    .X(_0139_));
 sg13g2_mux2_1 _1936_ (.A0(net434),
    .A1(net253),
    .S(_0003_),
    .X(_0140_));
 sg13g2_mux2_1 _1937_ (.A0(net264),
    .A1(\Ma[0] ),
    .S(net292),
    .X(_0141_));
 sg13g2_mux2_1 _1938_ (.A0(net354),
    .A1(\Ma[1] ),
    .S(net291),
    .X(_0142_));
 sg13g2_mux2_1 _1939_ (.A0(net241),
    .A1(\Ma[2] ),
    .S(net294),
    .X(_0143_));
 sg13g2_mux2_1 _1940_ (.A0(net249),
    .A1(\Ma[3] ),
    .S(net294),
    .X(_0144_));
 sg13g2_mux2_1 _1941_ (.A0(net251),
    .A1(net315),
    .S(net291),
    .X(_0145_));
 sg13g2_mux2_1 _1942_ (.A0(net234),
    .A1(net314),
    .S(net291),
    .X(_0146_));
 sg13g2_mux2_1 _1943_ (.A0(net374),
    .A1(net313),
    .S(net292),
    .X(_0147_));
 sg13g2_mux2_1 _1944_ (.A0(net381),
    .A1(\Ma[7] ),
    .S(net291),
    .X(_0148_));
 sg13g2_nor2_1 _1945_ (.A(net396),
    .B(net291),
    .Y(_0263_));
 sg13g2_a21oi_1 _1946_ (.A1(_0304_),
    .A2(net291),
    .Y(_0149_),
    .B1(_0263_));
 sg13g2_nor2_1 _1947_ (.A(net406),
    .B(net291),
    .Y(_0264_));
 sg13g2_a21oi_1 _1948_ (.A1(net298),
    .A2(net291),
    .Y(_0150_),
    .B1(_0264_));
 sg13g2_mux2_1 _1949_ (.A0(net243),
    .A1(\Mb[0] ),
    .S(net292),
    .X(_0151_));
 sg13g2_mux2_1 _1950_ (.A0(net259),
    .A1(\Mb[1] ),
    .S(net292),
    .X(_0152_));
 sg13g2_mux2_1 _1951_ (.A0(net192),
    .A1(\Mb[2] ),
    .S(net289),
    .X(_0153_));
 sg13g2_mux2_1 _1952_ (.A0(net210),
    .A1(net307),
    .S(net289),
    .X(_0154_));
 sg13g2_mux2_1 _1953_ (.A0(net363),
    .A1(net306),
    .S(net288),
    .X(_0155_));
 sg13g2_mux2_1 _1954_ (.A0(net386),
    .A1(net305),
    .S(net288),
    .X(_0156_));
 sg13g2_mux2_1 _1955_ (.A0(net218),
    .A1(net304),
    .S(net288),
    .X(_0157_));
 sg13g2_nor2_1 _1956_ (.A(net399),
    .B(net288),
    .Y(_0265_));
 sg13g2_a21oi_1 _1957_ (.A1(_0310_),
    .A2(net288),
    .Y(_0158_),
    .B1(_0265_));
 sg13g2_nor2_1 _1958_ (.A(net263),
    .B(net289),
    .Y(_0266_));
 sg13g2_a21oi_1 _1959_ (.A1(_0309_),
    .A2(net289),
    .Y(_0159_),
    .B1(_0266_));
 sg13g2_nor2_1 _1960_ (.A(net378),
    .B(net288),
    .Y(_0267_));
 sg13g2_a21oi_1 _1961_ (.A1(net297),
    .A2(net288),
    .Y(_0160_),
    .B1(_0267_));
 sg13g2_dfrbp_1 _1962_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net36),
    .D(_0006_),
    .Q_N(_0973_),
    .Q(\state[0] ));
 sg13g2_dfrbp_1 _1963_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net37),
    .D(_0000_),
    .Q_N(_0974_),
    .Q(\state[1] ));
 sg13g2_dfrbp_1 _1964_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net38),
    .D(_0007_),
    .Q_N(_0975_),
    .Q(\state[2] ));
 sg13g2_dfrbp_1 _1965_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net39),
    .D(_0001_),
    .Q_N(_0976_),
    .Q(\state[3] ));
 sg13g2_dfrbp_1 _1966_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net40),
    .D(_0002_),
    .Q_N(_0977_),
    .Q(\state[4] ));
 sg13g2_dfrbp_1 _1967_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net41),
    .D(_0008_),
    .Q_N(_0978_),
    .Q(\state[5] ));
 sg13g2_dfrbp_1 _1968_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net42),
    .D(_0003_),
    .Q_N(_0979_),
    .Q(\state[6] ));
 sg13g2_dfrbp_1 _1969_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net151),
    .D(_0004_),
    .Q_N(_0980_),
    .Q(\state[7] ));
 sg13g2_dfrbp_1 _1970_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net35),
    .D(_0005_),
    .Q_N(_0972_),
    .Q(\state[8] ));
 sg13g2_dfrbp_1 _1971_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net137),
    .D(_0023_),
    .Q_N(_0971_),
    .Q(\Mout[0] ));
 sg13g2_dfrbp_1 _1972_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net136),
    .D(_0024_),
    .Q_N(_0970_),
    .Q(\Mout[1] ));
 sg13g2_dfrbp_1 _1973_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net135),
    .D(_0025_),
    .Q_N(_0969_),
    .Q(\Mout[2] ));
 sg13g2_dfrbp_1 _1974_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net134),
    .D(_0026_),
    .Q_N(_0968_),
    .Q(\Mout[3] ));
 sg13g2_dfrbp_1 _1975_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net133),
    .D(_0027_),
    .Q_N(_0967_),
    .Q(\Mout[4] ));
 sg13g2_dfrbp_1 _1976_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net132),
    .D(_0028_),
    .Q_N(_0966_),
    .Q(\Mout[5] ));
 sg13g2_dfrbp_1 _1977_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net131),
    .D(_0029_),
    .Q_N(_0965_),
    .Q(\Mout[6] ));
 sg13g2_dfrbp_1 _1978_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net130),
    .D(_0030_),
    .Q_N(_0964_),
    .Q(\Mout[7] ));
 sg13g2_dfrbp_1 _1979_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net129),
    .D(_0031_),
    .Q_N(_0963_),
    .Q(\Mout[8] ));
 sg13g2_dfrbp_1 _1980_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net128),
    .D(_0032_),
    .Q_N(_0962_),
    .Q(\Mout[9] ));
 sg13g2_dfrbp_1 _1981_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net127),
    .D(_0033_),
    .Q_N(_0961_),
    .Q(\A[0] ));
 sg13g2_dfrbp_1 _1982_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net125),
    .D(_0034_),
    .Q_N(_0960_),
    .Q(\A[1] ));
 sg13g2_dfrbp_1 _1983_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net123),
    .D(_0035_),
    .Q_N(_0959_),
    .Q(\A[2] ));
 sg13g2_dfrbp_1 _1984_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net121),
    .D(_0036_),
    .Q_N(_0958_),
    .Q(\A[3] ));
 sg13g2_dfrbp_1 _1985_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net119),
    .D(_0037_),
    .Q_N(_0957_),
    .Q(\A[4] ));
 sg13g2_dfrbp_1 _1986_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net117),
    .D(_0038_),
    .Q_N(_0956_),
    .Q(\A[5] ));
 sg13g2_dfrbp_1 _1987_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net115),
    .D(_0039_),
    .Q_N(_0955_),
    .Q(\A[6] ));
 sg13g2_dfrbp_1 _1988_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net113),
    .D(_0040_),
    .Q_N(_0954_),
    .Q(\A[7] ));
 sg13g2_dfrbp_1 _1989_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net111),
    .D(_0041_),
    .Q_N(_0953_),
    .Q(\A[8] ));
 sg13g2_dfrbp_1 _1990_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net109),
    .D(_0042_),
    .Q_N(_0952_),
    .Q(\A[9] ));
 sg13g2_dfrbp_1 _1991_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net107),
    .D(_0043_),
    .Q_N(_0951_),
    .Q(\A[10] ));
 sg13g2_dfrbp_1 _1992_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net105),
    .D(_0044_),
    .Q_N(_0950_),
    .Q(\A[11] ));
 sg13g2_dfrbp_1 _1993_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net103),
    .D(_0045_),
    .Q_N(_0949_),
    .Q(\A[12] ));
 sg13g2_dfrbp_1 _1994_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net101),
    .D(_0046_),
    .Q_N(_0948_),
    .Q(\A[13] ));
 sg13g2_dfrbp_1 _1995_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net99),
    .D(_0047_),
    .Q_N(_0947_),
    .Q(\A[14] ));
 sg13g2_dfrbp_1 _1996_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net97),
    .D(_0048_),
    .Q_N(_0946_),
    .Q(\A[15] ));
 sg13g2_dfrbp_1 _1997_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net95),
    .D(_0049_),
    .Q_N(_0945_),
    .Q(\B[0] ));
 sg13g2_dfrbp_1 _1998_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net93),
    .D(_0050_),
    .Q_N(_0944_),
    .Q(\B[1] ));
 sg13g2_dfrbp_1 _1999_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net91),
    .D(_0051_),
    .Q_N(_0943_),
    .Q(\B[2] ));
 sg13g2_dfrbp_1 _2000_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net89),
    .D(_0052_),
    .Q_N(_0942_),
    .Q(\B[3] ));
 sg13g2_dfrbp_1 _2001_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net87),
    .D(_0053_),
    .Q_N(_0941_),
    .Q(\B[4] ));
 sg13g2_dfrbp_1 _2002_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net85),
    .D(_0054_),
    .Q_N(_0940_),
    .Q(\B[5] ));
 sg13g2_dfrbp_1 _2003_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net83),
    .D(_0055_),
    .Q_N(_0939_),
    .Q(\B[6] ));
 sg13g2_dfrbp_1 _2004_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net81),
    .D(_0056_),
    .Q_N(_0938_),
    .Q(\B[7] ));
 sg13g2_dfrbp_1 _2005_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net79),
    .D(_0057_),
    .Q_N(_0937_),
    .Q(\B[8] ));
 sg13g2_dfrbp_1 _2006_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net77),
    .D(_0058_),
    .Q_N(_0936_),
    .Q(\B[9] ));
 sg13g2_dfrbp_1 _2007_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net75),
    .D(_0059_),
    .Q_N(_0935_),
    .Q(\B[10] ));
 sg13g2_dfrbp_1 _2008_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net73),
    .D(_0060_),
    .Q_N(_0934_),
    .Q(\B[11] ));
 sg13g2_dfrbp_1 _2009_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net71),
    .D(_0061_),
    .Q_N(_0933_),
    .Q(\B[12] ));
 sg13g2_dfrbp_1 _2010_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net69),
    .D(_0062_),
    .Q_N(_0932_),
    .Q(\B[13] ));
 sg13g2_dfrbp_1 _2011_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net67),
    .D(_0063_),
    .Q_N(_0931_),
    .Q(\B[14] ));
 sg13g2_dfrbp_1 _2012_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net65),
    .D(_0064_),
    .Q_N(_0930_),
    .Q(\B[15] ));
 sg13g2_dfrbp_1 _2013_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net63),
    .D(net405),
    .Q_N(_0929_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _2014_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net61),
    .D(net413),
    .Q_N(_0928_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _2015_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net59),
    .D(net359),
    .Q_N(_0927_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _2016_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net57),
    .D(net395),
    .Q_N(_0926_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _2017_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net55),
    .D(net401),
    .Q_N(_0925_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _2018_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net53),
    .D(net403),
    .Q_N(_0924_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _2019_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net51),
    .D(net391),
    .Q_N(_0923_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _2020_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net49),
    .D(net371),
    .Q_N(_0922_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _2021_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net47),
    .D(net225),
    .Q_N(_0921_),
    .Q(\result[0] ));
 sg13g2_dfrbp_1 _2022_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net45),
    .D(net353),
    .Q_N(_0920_),
    .Q(\result[1] ));
 sg13g2_dfrbp_1 _2023_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net43),
    .D(net367),
    .Q_N(_0919_),
    .Q(\result[2] ));
 sg13g2_dfrbp_1 _2024_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net180),
    .D(_0076_),
    .Q_N(_0918_),
    .Q(\result[3] ));
 sg13g2_dfrbp_1 _2025_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net178),
    .D(net384),
    .Q_N(_0917_),
    .Q(\result[4] ));
 sg13g2_dfrbp_1 _2026_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net176),
    .D(net258),
    .Q_N(_0916_),
    .Q(\result[5] ));
 sg13g2_dfrbp_1 _2027_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net174),
    .D(net248),
    .Q_N(_0915_),
    .Q(\result[6] ));
 sg13g2_dfrbp_1 _2028_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net172),
    .D(net240),
    .Q_N(_0914_),
    .Q(\result[7] ));
 sg13g2_dfrbp_1 _2029_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net170),
    .D(net202),
    .Q_N(_0913_),
    .Q(\result[8] ));
 sg13g2_dfrbp_1 _2030_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net168),
    .D(net237),
    .Q_N(_0912_),
    .Q(\result[9] ));
 sg13g2_dfrbp_1 _2031_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net166),
    .D(net189),
    .Q_N(_0911_),
    .Q(\result[10] ));
 sg13g2_dfrbp_1 _2032_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net164),
    .D(net184),
    .Q_N(_0910_),
    .Q(\result[11] ));
 sg13g2_dfrbp_1 _2033_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net162),
    .D(net215),
    .Q_N(_0909_),
    .Q(\result[12] ));
 sg13g2_dfrbp_1 _2034_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net160),
    .D(_0086_),
    .Q_N(_0908_),
    .Q(\result[13] ));
 sg13g2_dfrbp_1 _2035_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net158),
    .D(net191),
    .Q_N(_0907_),
    .Q(\result[14] ));
 sg13g2_dfrbp_1 _2036_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net156),
    .D(net213),
    .Q_N(_0906_),
    .Q(\result[15] ));
 sg13g2_dfrbp_1 _2037_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net154),
    .D(_0089_),
    .Q_N(_0009_),
    .Q(\byte_count[0] ));
 sg13g2_dfrbp_1 _2038_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net152),
    .D(_0090_),
    .Q_N(_0905_),
    .Q(\byte_count[1] ));
 sg13g2_dfrbp_1 _2039_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net150),
    .D(net430),
    .Q_N(_0904_),
    .Q(\M1aout[0] ));
 sg13g2_dfrbp_1 _2040_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net149),
    .D(net380),
    .Q_N(_0903_),
    .Q(\M1aout[1] ));
 sg13g2_dfrbp_1 _2041_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net148),
    .D(_0093_),
    .Q_N(_0902_),
    .Q(\M1aout[2] ));
 sg13g2_dfrbp_1 _2042_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net147),
    .D(_0094_),
    .Q_N(_0901_),
    .Q(\M1aout[3] ));
 sg13g2_dfrbp_1 _2043_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net146),
    .D(net426),
    .Q_N(_0900_),
    .Q(\M1aout[4] ));
 sg13g2_dfrbp_1 _2044_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net145),
    .D(net421),
    .Q_N(_0899_),
    .Q(\M1aout[5] ));
 sg13g2_dfrbp_1 _2045_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net144),
    .D(net424),
    .Q_N(_0898_),
    .Q(\M1aout[6] ));
 sg13g2_dfrbp_1 _2046_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net143),
    .D(net438),
    .Q_N(_0897_),
    .Q(\M1aout[7] ));
 sg13g2_dfrbp_1 _2047_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net142),
    .D(net389),
    .Q_N(_0896_),
    .Q(\M1aout[8] ));
 sg13g2_dfrbp_1 _2048_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net141),
    .D(net433),
    .Q_N(_0895_),
    .Q(\M1aout[9] ));
 sg13g2_dfrbp_1 _2049_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net140),
    .D(_0101_),
    .Q_N(_0894_),
    .Q(\M1bout[0] ));
 sg13g2_dfrbp_1 _2050_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net139),
    .D(net415),
    .Q_N(_0893_),
    .Q(\M1bout[1] ));
 sg13g2_dfrbp_1 _2051_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net138),
    .D(net393),
    .Q_N(_0892_),
    .Q(\M1bout[2] ));
 sg13g2_dfrbp_1 _2052_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net126),
    .D(_0104_),
    .Q_N(_0891_),
    .Q(\M1bout[3] ));
 sg13g2_dfrbp_1 _2053_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net124),
    .D(_0105_),
    .Q_N(_0890_),
    .Q(\M1bout[4] ));
 sg13g2_dfrbp_1 _2054_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net122),
    .D(net409),
    .Q_N(_0889_),
    .Q(\M1bout[5] ));
 sg13g2_dfrbp_1 _2055_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net120),
    .D(net419),
    .Q_N(_0888_),
    .Q(\M1bout[6] ));
 sg13g2_dfrbp_1 _2056_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net118),
    .D(net417),
    .Q_N(_0887_),
    .Q(\M1bout[7] ));
 sg13g2_dfrbp_1 _2057_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net116),
    .D(net377),
    .Q_N(_0886_),
    .Q(\M1bout[8] ));
 sg13g2_dfrbp_1 _2058_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net114),
    .D(net436),
    .Q_N(_0885_),
    .Q(\M1bout[9] ));
 sg13g2_dfrbp_1 _2059_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net112),
    .D(net232),
    .Q_N(_0884_),
    .Q(\M1addout[0] ));
 sg13g2_dfrbp_1 _2060_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net110),
    .D(_0112_),
    .Q_N(_0883_),
    .Q(\M1addout[1] ));
 sg13g2_dfrbp_1 _2061_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net108),
    .D(_0113_),
    .Q_N(_0882_),
    .Q(\M1addout[2] ));
 sg13g2_dfrbp_1 _2062_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net106),
    .D(_0114_),
    .Q_N(_0881_),
    .Q(\M1addout[3] ));
 sg13g2_dfrbp_1 _2063_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net104),
    .D(_0115_),
    .Q_N(_0880_),
    .Q(\M1addout[4] ));
 sg13g2_dfrbp_1 _2064_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net102),
    .D(_0116_),
    .Q_N(_0879_),
    .Q(\M1addout[5] ));
 sg13g2_dfrbp_1 _2065_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net100),
    .D(net444),
    .Q_N(_0878_),
    .Q(\M1addout[6] ));
 sg13g2_dfrbp_1 _2066_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net98),
    .D(_0118_),
    .Q_N(_0877_),
    .Q(\M1addout[7] ));
 sg13g2_dfrbp_1 _2067_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net96),
    .D(_0119_),
    .Q_N(_0876_),
    .Q(\M1addout[8] ));
 sg13g2_dfrbp_1 _2068_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net94),
    .D(_0120_),
    .Q_N(_0022_),
    .Q(\M1addout[9] ));
 sg13g2_dfrbp_1 _2069_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net92),
    .D(net255),
    .Q_N(_0875_),
    .Q(\M1addout[10] ));
 sg13g2_dfrbp_1 _2070_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net90),
    .D(_0122_),
    .Q_N(_0874_),
    .Q(\Eout[0] ));
 sg13g2_dfrbp_1 _2071_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net88),
    .D(_0123_),
    .Q_N(_0873_),
    .Q(\Eout[1] ));
 sg13g2_dfrbp_1 _2072_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net86),
    .D(_0124_),
    .Q_N(_0872_),
    .Q(\Eout[2] ));
 sg13g2_dfrbp_1 _2073_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net84),
    .D(_0125_),
    .Q_N(_0871_),
    .Q(\Eout[3] ));
 sg13g2_dfrbp_1 _2074_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net82),
    .D(_0126_),
    .Q_N(_0870_),
    .Q(\Eout[4] ));
 sg13g2_dfrbp_1 _2075_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net80),
    .D(_0127_),
    .Q_N(_0869_),
    .Q(\Ea[0] ));
 sg13g2_dfrbp_1 _2076_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net78),
    .D(_0128_),
    .Q_N(_0868_),
    .Q(\Ea[1] ));
 sg13g2_dfrbp_1 _2077_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net76),
    .D(_0129_),
    .Q_N(_0867_),
    .Q(\Ea[2] ));
 sg13g2_dfrbp_1 _2078_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net74),
    .D(net196),
    .Q_N(_0866_),
    .Q(\Ea[3] ));
 sg13g2_dfrbp_1 _2079_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net72),
    .D(_0131_),
    .Q_N(_0865_),
    .Q(\Ea[4] ));
 sg13g2_dfrbp_1 _2080_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net70),
    .D(_0132_),
    .Q_N(_0864_),
    .Q(\Eb[0] ));
 sg13g2_dfrbp_1 _2081_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net68),
    .D(_0133_),
    .Q_N(_0863_),
    .Q(\Eb[1] ));
 sg13g2_dfrbp_1 _2082_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net66),
    .D(_0134_),
    .Q_N(_0862_),
    .Q(\Eb[2] ));
 sg13g2_dfrbp_1 _2083_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net64),
    .D(_0135_),
    .Q_N(_0861_),
    .Q(\Eb[3] ));
 sg13g2_dfrbp_1 _2084_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net62),
    .D(net361),
    .Q_N(_0860_),
    .Q(\Eb[4] ));
 sg13g2_dfrbp_1 _2085_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net60),
    .D(net228),
    .Q_N(_0859_),
    .Q(Sout));
 sg13g2_dfrbp_1 _2086_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net58),
    .D(net198),
    .Q_N(_0858_),
    .Q(Sa));
 sg13g2_dfrbp_1 _2087_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net56),
    .D(_0139_),
    .Q_N(_0857_),
    .Q(Sb));
 sg13g2_dfrbp_1 _2088_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net54),
    .D(_0140_),
    .Q_N(_0856_),
    .Q(Ce));
 sg13g2_dfrbp_1 _2089_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net52),
    .D(net265),
    .Q_N(_0855_),
    .Q(\Ma[0] ));
 sg13g2_dfrbp_1 _2090_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net50),
    .D(net355),
    .Q_N(_0854_),
    .Q(\Ma[1] ));
 sg13g2_dfrbp_1 _2091_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net48),
    .D(net242),
    .Q_N(_0853_),
    .Q(\Ma[2] ));
 sg13g2_dfrbp_1 _2092_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net46),
    .D(net250),
    .Q_N(_0852_),
    .Q(\Ma[3] ));
 sg13g2_dfrbp_1 _2093_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net44),
    .D(net252),
    .Q_N(_0011_),
    .Q(\Ma[4] ));
 sg13g2_dfrbp_1 _2094_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net34),
    .D(net235),
    .Q_N(_0012_),
    .Q(\Ma[5] ));
 sg13g2_dfrbp_1 _2095_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net179),
    .D(net375),
    .Q_N(_0013_),
    .Q(\Ma[6] ));
 sg13g2_dfrbp_1 _2096_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net177),
    .D(net382),
    .Q_N(_0014_),
    .Q(\Ma[7] ));
 sg13g2_dfrbp_1 _2097_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net175),
    .D(net397),
    .Q_N(_0015_),
    .Q(\Ma[8] ));
 sg13g2_dfrbp_1 _2098_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net173),
    .D(_0150_),
    .Q_N(_0010_),
    .Q(\Ma[9] ));
 sg13g2_dfrbp_1 _2099_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net171),
    .D(net244),
    .Q_N(_0851_),
    .Q(\Mb[0] ));
 sg13g2_dfrbp_1 _2100_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net169),
    .D(net260),
    .Q_N(_0850_),
    .Q(\Mb[1] ));
 sg13g2_dfrbp_1 _2101_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net167),
    .D(net193),
    .Q_N(_0849_),
    .Q(\Mb[2] ));
 sg13g2_dfrbp_1 _2102_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net165),
    .D(net211),
    .Q_N(_0848_),
    .Q(\Mb[3] ));
 sg13g2_dfrbp_1 _2103_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net163),
    .D(net364),
    .Q_N(_0017_),
    .Q(\Mb[4] ));
 sg13g2_dfrbp_1 _2104_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net161),
    .D(net387),
    .Q_N(_0018_),
    .Q(\Mb[5] ));
 sg13g2_dfrbp_1 _2105_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net159),
    .D(net219),
    .Q_N(_0019_),
    .Q(\Mb[6] ));
 sg13g2_dfrbp_1 _2106_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net157),
    .D(_0158_),
    .Q_N(_0020_),
    .Q(\Mb[7] ));
 sg13g2_dfrbp_1 _2107_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net155),
    .D(_0159_),
    .Q_N(_0021_),
    .Q(\Mb[8] ));
 sg13g2_dfrbp_1 _2108_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net153),
    .D(_0160_),
    .Q_N(_0016_),
    .Q(\Mb[9] ));
 sg13g2_tiehi _1970__35 (.L_HI(net35));
 sg13g2_tiehi _1962__36 (.L_HI(net36));
 sg13g2_tiehi _1963__37 (.L_HI(net37));
 sg13g2_tiehi _1964__38 (.L_HI(net38));
 sg13g2_tiehi _1965__39 (.L_HI(net39));
 sg13g2_tiehi _1966__40 (.L_HI(net40));
 sg13g2_tiehi _1967__41 (.L_HI(net41));
 sg13g2_tiehi _1968__42 (.L_HI(net42));
 sg13g2_tiehi _2023__43 (.L_HI(net43));
 sg13g2_tiehi _2093__44 (.L_HI(net44));
 sg13g2_tiehi _2022__45 (.L_HI(net45));
 sg13g2_tiehi _2092__46 (.L_HI(net46));
 sg13g2_tiehi _2021__47 (.L_HI(net47));
 sg13g2_tiehi _2091__48 (.L_HI(net48));
 sg13g2_tiehi _2020__49 (.L_HI(net49));
 sg13g2_tiehi _2090__50 (.L_HI(net50));
 sg13g2_tiehi _2019__51 (.L_HI(net51));
 sg13g2_tiehi _2089__52 (.L_HI(net52));
 sg13g2_tiehi _2018__53 (.L_HI(net53));
 sg13g2_tiehi _2088__54 (.L_HI(net54));
 sg13g2_tiehi _2017__55 (.L_HI(net55));
 sg13g2_tiehi _2087__56 (.L_HI(net56));
 sg13g2_tiehi _2016__57 (.L_HI(net57));
 sg13g2_tiehi _2086__58 (.L_HI(net58));
 sg13g2_tiehi _2015__59 (.L_HI(net59));
 sg13g2_tiehi _2085__60 (.L_HI(net60));
 sg13g2_tiehi _2014__61 (.L_HI(net61));
 sg13g2_tiehi _2084__62 (.L_HI(net62));
 sg13g2_tiehi _2013__63 (.L_HI(net63));
 sg13g2_tiehi _2083__64 (.L_HI(net64));
 sg13g2_tiehi _2012__65 (.L_HI(net65));
 sg13g2_tiehi _2082__66 (.L_HI(net66));
 sg13g2_tiehi _2011__67 (.L_HI(net67));
 sg13g2_tiehi _2081__68 (.L_HI(net68));
 sg13g2_tiehi _2010__69 (.L_HI(net69));
 sg13g2_tiehi _2080__70 (.L_HI(net70));
 sg13g2_tiehi _2009__71 (.L_HI(net71));
 sg13g2_tiehi _2079__72 (.L_HI(net72));
 sg13g2_tiehi _2008__73 (.L_HI(net73));
 sg13g2_tiehi _2078__74 (.L_HI(net74));
 sg13g2_tiehi _2007__75 (.L_HI(net75));
 sg13g2_tiehi _2077__76 (.L_HI(net76));
 sg13g2_tiehi _2006__77 (.L_HI(net77));
 sg13g2_tiehi _2076__78 (.L_HI(net78));
 sg13g2_tiehi _2005__79 (.L_HI(net79));
 sg13g2_tiehi _2075__80 (.L_HI(net80));
 sg13g2_tiehi _2004__81 (.L_HI(net81));
 sg13g2_tiehi _2074__82 (.L_HI(net82));
 sg13g2_tiehi _2003__83 (.L_HI(net83));
 sg13g2_tiehi _2073__84 (.L_HI(net84));
 sg13g2_tiehi _2002__85 (.L_HI(net85));
 sg13g2_tiehi _2072__86 (.L_HI(net86));
 sg13g2_tiehi _2001__87 (.L_HI(net87));
 sg13g2_tiehi _2071__88 (.L_HI(net88));
 sg13g2_tiehi _2000__89 (.L_HI(net89));
 sg13g2_tiehi _2070__90 (.L_HI(net90));
 sg13g2_tiehi _1999__91 (.L_HI(net91));
 sg13g2_tiehi _2069__92 (.L_HI(net92));
 sg13g2_tiehi _1998__93 (.L_HI(net93));
 sg13g2_tiehi _2068__94 (.L_HI(net94));
 sg13g2_tiehi _1997__95 (.L_HI(net95));
 sg13g2_tiehi _2067__96 (.L_HI(net96));
 sg13g2_tiehi _1996__97 (.L_HI(net97));
 sg13g2_tiehi _2066__98 (.L_HI(net98));
 sg13g2_tiehi _1995__99 (.L_HI(net99));
 sg13g2_tiehi _2065__100 (.L_HI(net100));
 sg13g2_tiehi _1994__101 (.L_HI(net101));
 sg13g2_tiehi _2064__102 (.L_HI(net102));
 sg13g2_tiehi _1993__103 (.L_HI(net103));
 sg13g2_tiehi _2063__104 (.L_HI(net104));
 sg13g2_tiehi _1992__105 (.L_HI(net105));
 sg13g2_tiehi _2062__106 (.L_HI(net106));
 sg13g2_tiehi _1991__107 (.L_HI(net107));
 sg13g2_tiehi _2061__108 (.L_HI(net108));
 sg13g2_tiehi _1990__109 (.L_HI(net109));
 sg13g2_tiehi _2060__110 (.L_HI(net110));
 sg13g2_tiehi _1989__111 (.L_HI(net111));
 sg13g2_tiehi _2059__112 (.L_HI(net112));
 sg13g2_tiehi _1988__113 (.L_HI(net113));
 sg13g2_tiehi _2058__114 (.L_HI(net114));
 sg13g2_tiehi _1987__115 (.L_HI(net115));
 sg13g2_tiehi _2057__116 (.L_HI(net116));
 sg13g2_tiehi _1986__117 (.L_HI(net117));
 sg13g2_tiehi _2056__118 (.L_HI(net118));
 sg13g2_tiehi _1985__119 (.L_HI(net119));
 sg13g2_tiehi _2055__120 (.L_HI(net120));
 sg13g2_tiehi _1984__121 (.L_HI(net121));
 sg13g2_tiehi _2054__122 (.L_HI(net122));
 sg13g2_tiehi _1983__123 (.L_HI(net123));
 sg13g2_tiehi _2053__124 (.L_HI(net124));
 sg13g2_tiehi _1982__125 (.L_HI(net125));
 sg13g2_tiehi _2052__126 (.L_HI(net126));
 sg13g2_tiehi _1981__127 (.L_HI(net127));
 sg13g2_tiehi _1980__128 (.L_HI(net128));
 sg13g2_tiehi _1979__129 (.L_HI(net129));
 sg13g2_tiehi _1978__130 (.L_HI(net130));
 sg13g2_tiehi _1977__131 (.L_HI(net131));
 sg13g2_tiehi _1976__132 (.L_HI(net132));
 sg13g2_tiehi _1975__133 (.L_HI(net133));
 sg13g2_tiehi _1974__134 (.L_HI(net134));
 sg13g2_tiehi _1973__135 (.L_HI(net135));
 sg13g2_tiehi _1972__136 (.L_HI(net136));
 sg13g2_tiehi _1971__137 (.L_HI(net137));
 sg13g2_tiehi _2051__138 (.L_HI(net138));
 sg13g2_tiehi _2050__139 (.L_HI(net139));
 sg13g2_tiehi _2049__140 (.L_HI(net140));
 sg13g2_tiehi _2048__141 (.L_HI(net141));
 sg13g2_tiehi _2047__142 (.L_HI(net142));
 sg13g2_tiehi _2046__143 (.L_HI(net143));
 sg13g2_tiehi _2045__144 (.L_HI(net144));
 sg13g2_tiehi _2044__145 (.L_HI(net145));
 sg13g2_tiehi _2043__146 (.L_HI(net146));
 sg13g2_tiehi _2042__147 (.L_HI(net147));
 sg13g2_tiehi _2041__148 (.L_HI(net148));
 sg13g2_tiehi _2040__149 (.L_HI(net149));
 sg13g2_tiehi _2039__150 (.L_HI(net150));
 sg13g2_tiehi _1969__151 (.L_HI(net151));
 sg13g2_tiehi _2038__152 (.L_HI(net152));
 sg13g2_tiehi _2108__153 (.L_HI(net153));
 sg13g2_tiehi _2037__154 (.L_HI(net154));
 sg13g2_tiehi _2107__155 (.L_HI(net155));
 sg13g2_tiehi _2036__156 (.L_HI(net156));
 sg13g2_tiehi _2106__157 (.L_HI(net157));
 sg13g2_tiehi _2035__158 (.L_HI(net158));
 sg13g2_tiehi _2105__159 (.L_HI(net159));
 sg13g2_tiehi _2034__160 (.L_HI(net160));
 sg13g2_tiehi _2104__161 (.L_HI(net161));
 sg13g2_tiehi _2033__162 (.L_HI(net162));
 sg13g2_tiehi _2103__163 (.L_HI(net163));
 sg13g2_tiehi _2032__164 (.L_HI(net164));
 sg13g2_tiehi _2102__165 (.L_HI(net165));
 sg13g2_tiehi _2031__166 (.L_HI(net166));
 sg13g2_tiehi _2101__167 (.L_HI(net167));
 sg13g2_tiehi _2030__168 (.L_HI(net168));
 sg13g2_tiehi _2100__169 (.L_HI(net169));
 sg13g2_tiehi _2029__170 (.L_HI(net170));
 sg13g2_tiehi _2099__171 (.L_HI(net171));
 sg13g2_tiehi _2028__172 (.L_HI(net172));
 sg13g2_tiehi _2098__173 (.L_HI(net173));
 sg13g2_tiehi _2027__174 (.L_HI(net174));
 sg13g2_tiehi _2097__175 (.L_HI(net175));
 sg13g2_tiehi _2026__176 (.L_HI(net176));
 sg13g2_tiehi _2096__177 (.L_HI(net177));
 sg13g2_tiehi _2025__178 (.L_HI(net178));
 sg13g2_tiehi _2095__179 (.L_HI(net179));
 sg13g2_tiehi _2024__180 (.L_HI(net180));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_log_afpm_19 (.L_LO(net19));
 sg13g2_tielo tt_um_log_afpm_20 (.L_LO(net20));
 sg13g2_tielo tt_um_log_afpm_21 (.L_LO(net21));
 sg13g2_tielo tt_um_log_afpm_22 (.L_LO(net22));
 sg13g2_tielo tt_um_log_afpm_23 (.L_LO(net23));
 sg13g2_tielo tt_um_log_afpm_24 (.L_LO(net24));
 sg13g2_tielo tt_um_log_afpm_25 (.L_LO(net25));
 sg13g2_tielo tt_um_log_afpm_26 (.L_LO(net26));
 sg13g2_tielo tt_um_log_afpm_27 (.L_LO(net27));
 sg13g2_tielo tt_um_log_afpm_28 (.L_LO(net28));
 sg13g2_tielo tt_um_log_afpm_29 (.L_LO(net29));
 sg13g2_tielo tt_um_log_afpm_30 (.L_LO(net30));
 sg13g2_tielo tt_um_log_afpm_31 (.L_LO(net31));
 sg13g2_tielo tt_um_log_afpm_32 (.L_LO(net32));
 sg13g2_tielo tt_um_log_afpm_33 (.L_LO(net33));
 sg13g2_tiehi _2094__34 (.L_HI(net34));
 sg13g2_buf_4 fanout266 (.X(net266),
    .A(net267));
 sg13g2_buf_4 fanout267 (.X(net267),
    .A(_0529_));
 sg13g2_buf_2 fanout268 (.A(net269),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_0519_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(net271),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(net272),
    .X(net271));
 sg13g2_buf_1 fanout272 (.A(_0519_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_0355_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_0355_),
    .X(net274));
 sg13g2_buf_4 fanout275 (.X(net275),
    .A(_0000_));
 sg13g2_buf_2 fanout276 (.A(net278),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(net278),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_0354_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(net280),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_0353_),
    .X(net280));
 sg13g2_buf_4 fanout281 (.X(net281),
    .A(_0353_));
 sg13g2_buf_2 fanout282 (.A(net283),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(net284),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_0352_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(net286),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(net287),
    .X(net286));
 sg13g2_buf_4 fanout287 (.X(net287),
    .A(_0352_));
 sg13g2_buf_2 fanout288 (.A(net290),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(net290),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(net207),
    .X(net290));
 sg13g2_buf_4 fanout291 (.X(net291),
    .A(net292));
 sg13g2_buf_2 fanout292 (.A(net294),
    .X(net292));
 sg13g2_buf_4 fanout293 (.X(net293),
    .A(net294));
 sg13g2_buf_2 fanout294 (.A(_0351_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_0312_),
    .X(net295));
 sg13g2_buf_1 fanout296 (.A(_0312_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_0308_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_0303_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(\Mb[9] ),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(\Mb[9] ),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(net303),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(net303),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(\Mb[8] ),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(\Mb[6] ),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(\Mb[5] ),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(\Mb[4] ),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(\Mb[3] ),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(net309),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(\Ma[9] ),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(net311),
    .X(net310));
 sg13g2_buf_1 fanout311 (.A(net312),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(\Ma[8] ),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(\Ma[6] ),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(\Ma[5] ),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(\Ma[4] ),
    .X(net315));
 sg13g2_buf_4 fanout316 (.X(net316),
    .A(\Ma[3] ));
 sg13g2_buf_2 fanout317 (.A(net318),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(net319),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(net398),
    .X(net319));
 sg13g2_buf_4 fanout320 (.X(net320),
    .A(net362));
 sg13g2_buf_4 fanout321 (.X(net321),
    .A(net362));
 sg13g2_buf_4 fanout322 (.X(net322),
    .A(net323));
 sg13g2_buf_4 fanout323 (.X(net323),
    .A(\M1addout[7] ));
 sg13g2_buf_4 fanout324 (.X(net324),
    .A(net443));
 sg13g2_buf_2 fanout325 (.A(\M1addout[6] ),
    .X(net325));
 sg13g2_buf_4 fanout326 (.X(net326),
    .A(\M1addout[5] ));
 sg13g2_buf_2 fanout327 (.A(net447),
    .X(net327));
 sg13g2_buf_4 fanout328 (.X(net328),
    .A(net446));
 sg13g2_buf_2 fanout329 (.A(net445),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(net331),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(net332),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(\byte_count[0] ),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(net385),
    .X(net333));
 sg13g2_buf_1 fanout334 (.A(net385),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(net338),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(net338),
    .X(net336));
 sg13g2_buf_1 fanout337 (.A(net338),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(net340),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(net340),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(net440),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(net345),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(net345),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(net344),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(net345),
    .X(net344));
 sg13g2_buf_1 fanout345 (.A(_0293_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(net349),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(net349),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(net349),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(net1),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(net351),
    .X(net350));
 sg13g2_buf_4 fanout351 (.X(net351),
    .A(net1));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[0]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[1]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[2]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[3]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[4]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[5]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[6]),
    .X(net16));
 sg13g2_buf_1 input17 (.A(uio_in[7]),
    .X(net17));
 sg13g2_tielo tt_um_log_afpm_18 (.L_LO(net18));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0009_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0597_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold3 (.A(\Eout[1] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0084_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold5 (.A(\Eout[3] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold6 (.A(\state[8] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold7 (.A(\B[15] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold8 (.A(\Eout[0] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0083_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold10 (.A(\Eout[4] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0087_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold12 (.A(\B[2] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0153_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold14 (.A(\A[11] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold15 (.A(\A[13] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0130_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold17 (.A(\A[15] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0138_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold19 (.A(\B[11] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold20 (.A(\Eb[3] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold21 (.A(\Mout[8] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0081_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold23 (.A(\B[10] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold24 (.A(\Eb[0] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold25 (.A(\state[6] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold26 (.A(\state[7] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0351_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold28 (.A(\A[12] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold29 (.A(\state[5] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold30 (.A(\B[3] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0154_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold32 (.A(Sout),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0088_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold34 (.A(\Eout[2] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0085_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold36 (.A(\Ea[1] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold37 (.A(\B[12] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold38 (.A(\B[6] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0157_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold40 (.A(\Mout[0] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold41 (.A(\Eb[1] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold42 (.A(\A[14] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold43 (.A(Sb),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold44 (.A(\result[0] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0073_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold46 (.A(\B[13] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold47 (.A(Sa),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0137_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold49 (.A(\state[0] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0349_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold51 (.A(\M1addout[0] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0111_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold53 (.A(\Ea[4] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold54 (.A(\A[5] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0146_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold56 (.A(\Mout[9] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0082_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold58 (.A(\Mout[3] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold59 (.A(\Mout[7] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0080_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold61 (.A(\A[2] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0143_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold63 (.A(\B[0] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0151_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold65 (.A(\Eb[2] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold66 (.A(\A[10] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold67 (.A(\Mout[6] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0079_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold69 (.A(\A[3] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0144_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold71 (.A(\A[4] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0145_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold73 (.A(\M1addout[10] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0225_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0121_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold76 (.A(\result[3] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold77 (.A(\Mout[5] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0078_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold79 (.A(\B[1] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0152_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold81 (.A(\result[13] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold82 (.A(\Ea[2] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold83 (.A(\B[8] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold84 (.A(\A[0] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0141_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold86 (.A(\Mout[1] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0074_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold88 (.A(\A[1] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0142_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold90 (.A(\M1addout[2] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold91 (.A(uo_out[2]),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0561_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0067_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold94 (.A(\B[14] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0136_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold96 (.A(\M1addout[8] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold97 (.A(\B[4] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0155_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold99 (.A(\M1bout[3] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold100 (.A(\Mout[2] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0075_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold102 (.A(\byte_count[1] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold103 (.A(uo_out[7]),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0576_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0072_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold106 (.A(\Ea[0] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold107 (.A(\byte_count[1] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold108 (.A(\A[6] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0147_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold110 (.A(\M1bout[8] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0109_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold112 (.A(\B[9] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold113 (.A(\M1aout[1] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0092_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold115 (.A(\A[7] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0148_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold117 (.A(\result[4] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0077_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold119 (.A(\state[2] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold120 (.A(\B[5] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0156_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold122 (.A(\M1aout[8] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0099_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold124 (.A(uo_out[6]),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0071_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold126 (.A(\M1bout[2] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0103_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold128 (.A(uo_out[3]),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0068_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold130 (.A(\A[8] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0149_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold132 (.A(\M1addout[9] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold133 (.A(\B[7] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold134 (.A(uo_out[4]),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0069_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold136 (.A(uo_out[5]),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0070_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold138 (.A(uo_out[0]),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0065_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold140 (.A(\A[9] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold141 (.A(\M1aout[3] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold142 (.A(\M1bout[5] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0106_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold144 (.A(\Mout[4] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold145 (.A(\Mb[7] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold146 (.A(uo_out[1]),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0066_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold148 (.A(\M1bout[1] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0102_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold150 (.A(\M1bout[7] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0108_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold152 (.A(\M1bout[6] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0107_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold154 (.A(\M1aout[5] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0096_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold156 (.A(\M1aout[2] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold157 (.A(\M1aout[6] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0097_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold159 (.A(\M1aout[4] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0095_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold161 (.A(\M1bout[0] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold162 (.A(\M1bout[4] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold163 (.A(\M1aout[0] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0091_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0015_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0727_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0100_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold168 (.A(Ce),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold169 (.A(\M1bout[9] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0110_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold171 (.A(\M1aout[7] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0098_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold173 (.A(\state[5] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold174 (.A(\state[1] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold175 (.A(\M1addout[1] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0184_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold177 (.A(\M1addout[6] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0117_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold179 (.A(\M1addout[3] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold180 (.A(\M1addout[4] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold181 (.A(\M1addout[5] ),
    .X(net447));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_4 FILLER_5_140 ();
 sg13g2_fill_2 FILLER_5_144 ();
 sg13g2_decap_8 FILLER_5_151 ();
 sg13g2_decap_8 FILLER_5_158 ();
 sg13g2_decap_8 FILLER_5_165 ();
 sg13g2_decap_8 FILLER_5_172 ();
 sg13g2_decap_8 FILLER_5_179 ();
 sg13g2_decap_8 FILLER_5_186 ();
 sg13g2_decap_8 FILLER_5_193 ();
 sg13g2_decap_8 FILLER_5_200 ();
 sg13g2_decap_8 FILLER_5_207 ();
 sg13g2_decap_8 FILLER_5_214 ();
 sg13g2_decap_8 FILLER_5_221 ();
 sg13g2_decap_8 FILLER_5_228 ();
 sg13g2_decap_8 FILLER_5_235 ();
 sg13g2_decap_8 FILLER_5_242 ();
 sg13g2_decap_8 FILLER_5_249 ();
 sg13g2_decap_8 FILLER_5_256 ();
 sg13g2_decap_8 FILLER_5_263 ();
 sg13g2_decap_8 FILLER_5_270 ();
 sg13g2_decap_8 FILLER_5_277 ();
 sg13g2_decap_8 FILLER_5_284 ();
 sg13g2_decap_8 FILLER_5_291 ();
 sg13g2_decap_8 FILLER_5_298 ();
 sg13g2_decap_8 FILLER_5_305 ();
 sg13g2_decap_8 FILLER_5_312 ();
 sg13g2_decap_8 FILLER_5_319 ();
 sg13g2_decap_8 FILLER_5_326 ();
 sg13g2_decap_8 FILLER_5_333 ();
 sg13g2_decap_8 FILLER_5_340 ();
 sg13g2_decap_8 FILLER_5_347 ();
 sg13g2_decap_8 FILLER_5_354 ();
 sg13g2_decap_8 FILLER_5_361 ();
 sg13g2_decap_8 FILLER_5_368 ();
 sg13g2_decap_8 FILLER_5_375 ();
 sg13g2_decap_8 FILLER_5_382 ();
 sg13g2_decap_8 FILLER_5_389 ();
 sg13g2_decap_8 FILLER_5_396 ();
 sg13g2_decap_4 FILLER_5_403 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_4 FILLER_6_133 ();
 sg13g2_fill_1 FILLER_6_137 ();
 sg13g2_fill_1 FILLER_6_146 ();
 sg13g2_fill_2 FILLER_6_159 ();
 sg13g2_decap_8 FILLER_6_165 ();
 sg13g2_decap_4 FILLER_6_172 ();
 sg13g2_fill_2 FILLER_6_176 ();
 sg13g2_decap_8 FILLER_6_216 ();
 sg13g2_decap_8 FILLER_6_227 ();
 sg13g2_decap_8 FILLER_6_234 ();
 sg13g2_fill_2 FILLER_6_241 ();
 sg13g2_decap_8 FILLER_6_247 ();
 sg13g2_fill_2 FILLER_6_254 ();
 sg13g2_decap_8 FILLER_6_263 ();
 sg13g2_fill_2 FILLER_6_270 ();
 sg13g2_fill_1 FILLER_6_272 ();
 sg13g2_fill_1 FILLER_6_283 ();
 sg13g2_decap_8 FILLER_6_313 ();
 sg13g2_decap_4 FILLER_6_320 ();
 sg13g2_fill_1 FILLER_6_324 ();
 sg13g2_decap_4 FILLER_6_340 ();
 sg13g2_fill_1 FILLER_6_344 ();
 sg13g2_decap_8 FILLER_6_381 ();
 sg13g2_decap_4 FILLER_6_388 ();
 sg13g2_fill_2 FILLER_6_392 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_fill_2 FILLER_7_119 ();
 sg13g2_decap_4 FILLER_7_125 ();
 sg13g2_fill_2 FILLER_7_129 ();
 sg13g2_fill_2 FILLER_7_144 ();
 sg13g2_fill_2 FILLER_7_261 ();
 sg13g2_fill_2 FILLER_7_293 ();
 sg13g2_fill_1 FILLER_7_295 ();
 sg13g2_fill_1 FILLER_7_309 ();
 sg13g2_fill_2 FILLER_7_324 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_4 FILLER_7_350 ();
 sg13g2_fill_2 FILLER_7_354 ();
 sg13g2_fill_1 FILLER_7_360 ();
 sg13g2_fill_1 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_fill_1 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_47 ();
 sg13g2_decap_8 FILLER_8_54 ();
 sg13g2_decap_4 FILLER_8_61 ();
 sg13g2_fill_2 FILLER_8_65 ();
 sg13g2_decap_8 FILLER_8_89 ();
 sg13g2_decap_8 FILLER_8_96 ();
 sg13g2_decap_8 FILLER_8_103 ();
 sg13g2_fill_1 FILLER_8_136 ();
 sg13g2_decap_4 FILLER_8_149 ();
 sg13g2_fill_2 FILLER_8_172 ();
 sg13g2_fill_2 FILLER_8_179 ();
 sg13g2_fill_2 FILLER_8_192 ();
 sg13g2_fill_1 FILLER_8_201 ();
 sg13g2_decap_8 FILLER_8_221 ();
 sg13g2_decap_4 FILLER_8_232 ();
 sg13g2_fill_2 FILLER_8_236 ();
 sg13g2_fill_2 FILLER_8_260 ();
 sg13g2_fill_1 FILLER_8_277 ();
 sg13g2_fill_2 FILLER_8_287 ();
 sg13g2_fill_2 FILLER_8_309 ();
 sg13g2_fill_1 FILLER_8_319 ();
 sg13g2_fill_2 FILLER_8_327 ();
 sg13g2_decap_4 FILLER_8_337 ();
 sg13g2_fill_1 FILLER_8_341 ();
 sg13g2_fill_2 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_4 FILLER_9_28 ();
 sg13g2_fill_2 FILLER_9_67 ();
 sg13g2_fill_1 FILLER_9_69 ();
 sg13g2_decap_4 FILLER_9_162 ();
 sg13g2_fill_1 FILLER_9_185 ();
 sg13g2_fill_1 FILLER_9_205 ();
 sg13g2_fill_2 FILLER_9_215 ();
 sg13g2_decap_4 FILLER_9_243 ();
 sg13g2_fill_1 FILLER_9_247 ();
 sg13g2_fill_2 FILLER_9_300 ();
 sg13g2_fill_1 FILLER_9_329 ();
 sg13g2_decap_4 FILLER_9_343 ();
 sg13g2_fill_1 FILLER_9_347 ();
 sg13g2_fill_2 FILLER_9_371 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_33 ();
 sg13g2_decap_8 FILLER_10_40 ();
 sg13g2_decap_4 FILLER_10_47 ();
 sg13g2_fill_1 FILLER_10_51 ();
 sg13g2_fill_2 FILLER_10_56 ();
 sg13g2_fill_1 FILLER_10_83 ();
 sg13g2_fill_2 FILLER_10_112 ();
 sg13g2_decap_4 FILLER_10_165 ();
 sg13g2_fill_2 FILLER_10_169 ();
 sg13g2_fill_2 FILLER_10_184 ();
 sg13g2_fill_1 FILLER_10_222 ();
 sg13g2_fill_2 FILLER_10_231 ();
 sg13g2_fill_1 FILLER_10_233 ();
 sg13g2_fill_2 FILLER_10_303 ();
 sg13g2_fill_1 FILLER_10_314 ();
 sg13g2_fill_1 FILLER_10_356 ();
 sg13g2_fill_2 FILLER_10_361 ();
 sg13g2_fill_1 FILLER_10_363 ();
 sg13g2_fill_1 FILLER_10_372 ();
 sg13g2_fill_2 FILLER_10_387 ();
 sg13g2_fill_1 FILLER_10_389 ();
 sg13g2_decap_4 FILLER_10_403 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_fill_2 FILLER_11_21 ();
 sg13g2_fill_1 FILLER_11_23 ();
 sg13g2_fill_2 FILLER_11_50 ();
 sg13g2_fill_1 FILLER_11_87 ();
 sg13g2_fill_2 FILLER_11_118 ();
 sg13g2_decap_4 FILLER_11_159 ();
 sg13g2_fill_1 FILLER_11_163 ();
 sg13g2_decap_4 FILLER_11_190 ();
 sg13g2_fill_2 FILLER_11_194 ();
 sg13g2_decap_8 FILLER_11_200 ();
 sg13g2_fill_2 FILLER_11_207 ();
 sg13g2_fill_1 FILLER_11_209 ();
 sg13g2_fill_2 FILLER_11_243 ();
 sg13g2_fill_1 FILLER_11_249 ();
 sg13g2_fill_1 FILLER_11_255 ();
 sg13g2_fill_2 FILLER_11_286 ();
 sg13g2_fill_1 FILLER_11_288 ();
 sg13g2_fill_2 FILLER_11_307 ();
 sg13g2_decap_4 FILLER_11_317 ();
 sg13g2_fill_2 FILLER_11_321 ();
 sg13g2_fill_1 FILLER_11_327 ();
 sg13g2_fill_1 FILLER_11_332 ();
 sg13g2_fill_2 FILLER_11_387 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_fill_1 FILLER_12_39 ();
 sg13g2_fill_1 FILLER_12_44 ();
 sg13g2_fill_2 FILLER_12_58 ();
 sg13g2_fill_1 FILLER_12_60 ();
 sg13g2_fill_2 FILLER_12_71 ();
 sg13g2_fill_1 FILLER_12_95 ();
 sg13g2_fill_1 FILLER_12_105 ();
 sg13g2_fill_2 FILLER_12_127 ();
 sg13g2_fill_2 FILLER_12_191 ();
 sg13g2_decap_4 FILLER_12_208 ();
 sg13g2_fill_2 FILLER_12_232 ();
 sg13g2_fill_1 FILLER_12_234 ();
 sg13g2_fill_2 FILLER_12_339 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_4 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_fill_1 FILLER_13_21 ();
 sg13g2_decap_4 FILLER_13_25 ();
 sg13g2_fill_1 FILLER_13_29 ();
 sg13g2_fill_2 FILLER_13_70 ();
 sg13g2_fill_1 FILLER_13_76 ();
 sg13g2_fill_2 FILLER_13_127 ();
 sg13g2_decap_8 FILLER_13_150 ();
 sg13g2_decap_4 FILLER_13_157 ();
 sg13g2_fill_1 FILLER_13_161 ();
 sg13g2_fill_1 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_202 ();
 sg13g2_fill_2 FILLER_13_209 ();
 sg13g2_fill_1 FILLER_13_216 ();
 sg13g2_fill_2 FILLER_13_237 ();
 sg13g2_decap_8 FILLER_13_244 ();
 sg13g2_decap_4 FILLER_13_255 ();
 sg13g2_fill_1 FILLER_13_259 ();
 sg13g2_fill_1 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_283 ();
 sg13g2_fill_2 FILLER_13_290 ();
 sg13g2_fill_1 FILLER_13_322 ();
 sg13g2_fill_2 FILLER_13_362 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_4 FILLER_14_7 ();
 sg13g2_fill_2 FILLER_14_11 ();
 sg13g2_fill_2 FILLER_14_34 ();
 sg13g2_fill_1 FILLER_14_36 ();
 sg13g2_decap_4 FILLER_14_41 ();
 sg13g2_fill_1 FILLER_14_45 ();
 sg13g2_decap_4 FILLER_14_54 ();
 sg13g2_decap_4 FILLER_14_96 ();
 sg13g2_fill_1 FILLER_14_118 ();
 sg13g2_fill_2 FILLER_14_145 ();
 sg13g2_fill_1 FILLER_14_147 ();
 sg13g2_fill_2 FILLER_14_152 ();
 sg13g2_fill_1 FILLER_14_154 ();
 sg13g2_fill_1 FILLER_14_163 ();
 sg13g2_fill_1 FILLER_14_182 ();
 sg13g2_fill_1 FILLER_14_214 ();
 sg13g2_decap_4 FILLER_14_236 ();
 sg13g2_fill_1 FILLER_14_240 ();
 sg13g2_decap_4 FILLER_14_344 ();
 sg13g2_fill_2 FILLER_14_359 ();
 sg13g2_fill_1 FILLER_14_361 ();
 sg13g2_decap_4 FILLER_14_366 ();
 sg13g2_fill_2 FILLER_14_370 ();
 sg13g2_fill_1 FILLER_14_377 ();
 sg13g2_decap_8 FILLER_14_388 ();
 sg13g2_fill_2 FILLER_14_395 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_7 ();
 sg13g2_fill_1 FILLER_15_9 ();
 sg13g2_decap_4 FILLER_15_15 ();
 sg13g2_fill_1 FILLER_15_19 ();
 sg13g2_fill_1 FILLER_15_38 ();
 sg13g2_fill_2 FILLER_15_47 ();
 sg13g2_decap_8 FILLER_15_94 ();
 sg13g2_fill_1 FILLER_15_114 ();
 sg13g2_fill_1 FILLER_15_177 ();
 sg13g2_fill_1 FILLER_15_186 ();
 sg13g2_decap_4 FILLER_15_205 ();
 sg13g2_decap_8 FILLER_15_221 ();
 sg13g2_decap_4 FILLER_15_233 ();
 sg13g2_fill_2 FILLER_15_237 ();
 sg13g2_fill_2 FILLER_15_263 ();
 sg13g2_fill_1 FILLER_15_265 ();
 sg13g2_fill_2 FILLER_15_341 ();
 sg13g2_decap_4 FILLER_15_347 ();
 sg13g2_fill_1 FILLER_15_351 ();
 sg13g2_decap_8 FILLER_15_362 ();
 sg13g2_fill_1 FILLER_15_369 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_4 ();
 sg13g2_decap_4 FILLER_16_22 ();
 sg13g2_fill_2 FILLER_16_26 ();
 sg13g2_decap_4 FILLER_16_32 ();
 sg13g2_fill_1 FILLER_16_36 ();
 sg13g2_decap_8 FILLER_16_46 ();
 sg13g2_fill_1 FILLER_16_53 ();
 sg13g2_fill_2 FILLER_16_69 ();
 sg13g2_fill_1 FILLER_16_71 ();
 sg13g2_decap_8 FILLER_16_96 ();
 sg13g2_decap_8 FILLER_16_103 ();
 sg13g2_fill_2 FILLER_16_128 ();
 sg13g2_decap_4 FILLER_16_139 ();
 sg13g2_fill_2 FILLER_16_143 ();
 sg13g2_decap_4 FILLER_16_183 ();
 sg13g2_fill_1 FILLER_16_200 ();
 sg13g2_fill_1 FILLER_16_206 ();
 sg13g2_fill_2 FILLER_16_219 ();
 sg13g2_fill_1 FILLER_16_277 ();
 sg13g2_fill_2 FILLER_16_328 ();
 sg13g2_fill_1 FILLER_16_330 ();
 sg13g2_decap_4 FILLER_16_335 ();
 sg13g2_fill_1 FILLER_16_339 ();
 sg13g2_fill_1 FILLER_16_370 ();
 sg13g2_decap_4 FILLER_16_390 ();
 sg13g2_fill_2 FILLER_16_394 ();
 sg13g2_decap_4 FILLER_16_404 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_4 ();
 sg13g2_decap_4 FILLER_17_40 ();
 sg13g2_fill_2 FILLER_17_44 ();
 sg13g2_fill_2 FILLER_17_82 ();
 sg13g2_fill_1 FILLER_17_97 ();
 sg13g2_fill_2 FILLER_17_114 ();
 sg13g2_fill_1 FILLER_17_116 ();
 sg13g2_fill_2 FILLER_17_121 ();
 sg13g2_fill_2 FILLER_17_153 ();
 sg13g2_fill_1 FILLER_17_155 ();
 sg13g2_fill_2 FILLER_17_180 ();
 sg13g2_decap_4 FILLER_17_195 ();
 sg13g2_decap_4 FILLER_17_208 ();
 sg13g2_fill_2 FILLER_17_212 ();
 sg13g2_decap_8 FILLER_17_219 ();
 sg13g2_fill_1 FILLER_17_226 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_4 FILLER_17_238 ();
 sg13g2_fill_2 FILLER_17_242 ();
 sg13g2_decap_4 FILLER_17_257 ();
 sg13g2_fill_1 FILLER_17_261 ();
 sg13g2_fill_2 FILLER_17_270 ();
 sg13g2_fill_1 FILLER_17_272 ();
 sg13g2_fill_1 FILLER_17_310 ();
 sg13g2_fill_1 FILLER_17_324 ();
 sg13g2_fill_1 FILLER_17_328 ();
 sg13g2_fill_2 FILLER_17_362 ();
 sg13g2_fill_1 FILLER_17_364 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_7 ();
 sg13g2_fill_1 FILLER_18_9 ();
 sg13g2_fill_2 FILLER_18_20 ();
 sg13g2_fill_1 FILLER_18_22 ();
 sg13g2_decap_4 FILLER_18_48 ();
 sg13g2_fill_2 FILLER_18_52 ();
 sg13g2_decap_8 FILLER_18_59 ();
 sg13g2_decap_8 FILLER_18_66 ();
 sg13g2_fill_1 FILLER_18_73 ();
 sg13g2_fill_2 FILLER_18_85 ();
 sg13g2_fill_1 FILLER_18_87 ();
 sg13g2_decap_4 FILLER_18_133 ();
 sg13g2_fill_1 FILLER_18_137 ();
 sg13g2_decap_8 FILLER_18_142 ();
 sg13g2_decap_4 FILLER_18_149 ();
 sg13g2_fill_1 FILLER_18_153 ();
 sg13g2_decap_8 FILLER_18_158 ();
 sg13g2_fill_1 FILLER_18_165 ();
 sg13g2_fill_1 FILLER_18_171 ();
 sg13g2_decap_8 FILLER_18_176 ();
 sg13g2_decap_8 FILLER_18_183 ();
 sg13g2_decap_4 FILLER_18_190 ();
 sg13g2_fill_1 FILLER_18_194 ();
 sg13g2_fill_2 FILLER_18_227 ();
 sg13g2_fill_1 FILLER_18_252 ();
 sg13g2_fill_1 FILLER_18_268 ();
 sg13g2_fill_2 FILLER_18_274 ();
 sg13g2_fill_1 FILLER_18_348 ();
 sg13g2_fill_1 FILLER_18_370 ();
 sg13g2_decap_4 FILLER_18_383 ();
 sg13g2_fill_1 FILLER_18_387 ();
 sg13g2_fill_1 FILLER_18_392 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_4 ();
 sg13g2_fill_1 FILLER_19_29 ();
 sg13g2_fill_2 FILLER_19_47 ();
 sg13g2_fill_1 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_67 ();
 sg13g2_fill_1 FILLER_19_74 ();
 sg13g2_fill_1 FILLER_19_83 ();
 sg13g2_fill_2 FILLER_19_94 ();
 sg13g2_fill_2 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_134 ();
 sg13g2_fill_2 FILLER_19_141 ();
 sg13g2_fill_1 FILLER_19_169 ();
 sg13g2_fill_2 FILLER_19_174 ();
 sg13g2_fill_1 FILLER_19_176 ();
 sg13g2_decap_8 FILLER_19_181 ();
 sg13g2_fill_1 FILLER_19_188 ();
 sg13g2_fill_2 FILLER_19_209 ();
 sg13g2_fill_1 FILLER_19_211 ();
 sg13g2_fill_2 FILLER_19_221 ();
 sg13g2_decap_4 FILLER_19_239 ();
 sg13g2_fill_2 FILLER_19_258 ();
 sg13g2_fill_1 FILLER_19_292 ();
 sg13g2_fill_1 FILLER_19_302 ();
 sg13g2_decap_8 FILLER_19_311 ();
 sg13g2_decap_4 FILLER_19_318 ();
 sg13g2_fill_2 FILLER_19_322 ();
 sg13g2_decap_4 FILLER_19_328 ();
 sg13g2_fill_1 FILLER_19_332 ();
 sg13g2_fill_1 FILLER_19_356 ();
 sg13g2_fill_2 FILLER_19_367 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_4 ();
 sg13g2_decap_8 FILLER_20_24 ();
 sg13g2_fill_2 FILLER_20_31 ();
 sg13g2_fill_1 FILLER_20_33 ();
 sg13g2_decap_8 FILLER_20_47 ();
 sg13g2_decap_4 FILLER_20_54 ();
 sg13g2_fill_1 FILLER_20_58 ();
 sg13g2_decap_4 FILLER_20_62 ();
 sg13g2_fill_1 FILLER_20_79 ();
 sg13g2_fill_1 FILLER_20_84 ();
 sg13g2_fill_2 FILLER_20_94 ();
 sg13g2_fill_2 FILLER_20_109 ();
 sg13g2_fill_1 FILLER_20_111 ();
 sg13g2_fill_1 FILLER_20_117 ();
 sg13g2_fill_1 FILLER_20_155 ();
 sg13g2_decap_4 FILLER_20_197 ();
 sg13g2_fill_1 FILLER_20_201 ();
 sg13g2_fill_2 FILLER_20_206 ();
 sg13g2_fill_1 FILLER_20_208 ();
 sg13g2_decap_8 FILLER_20_214 ();
 sg13g2_fill_2 FILLER_20_221 ();
 sg13g2_fill_1 FILLER_20_236 ();
 sg13g2_decap_4 FILLER_20_245 ();
 sg13g2_fill_1 FILLER_20_249 ();
 sg13g2_fill_1 FILLER_20_255 ();
 sg13g2_fill_2 FILLER_20_286 ();
 sg13g2_fill_1 FILLER_20_288 ();
 sg13g2_decap_8 FILLER_20_319 ();
 sg13g2_fill_2 FILLER_20_326 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_20 ();
 sg13g2_fill_1 FILLER_21_34 ();
 sg13g2_fill_1 FILLER_21_40 ();
 sg13g2_decap_4 FILLER_21_67 ();
 sg13g2_fill_1 FILLER_21_71 ();
 sg13g2_fill_2 FILLER_21_77 ();
 sg13g2_fill_2 FILLER_21_90 ();
 sg13g2_fill_1 FILLER_21_92 ();
 sg13g2_decap_4 FILLER_21_98 ();
 sg13g2_fill_2 FILLER_21_102 ();
 sg13g2_decap_4 FILLER_21_109 ();
 sg13g2_fill_2 FILLER_21_113 ();
 sg13g2_fill_2 FILLER_21_135 ();
 sg13g2_fill_2 FILLER_21_175 ();
 sg13g2_fill_1 FILLER_21_177 ();
 sg13g2_fill_1 FILLER_21_238 ();
 sg13g2_fill_2 FILLER_21_247 ();
 sg13g2_fill_1 FILLER_21_249 ();
 sg13g2_fill_2 FILLER_21_262 ();
 sg13g2_decap_8 FILLER_21_272 ();
 sg13g2_fill_1 FILLER_21_296 ();
 sg13g2_fill_2 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_400 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_11 ();
 sg13g2_decap_4 FILLER_22_25 ();
 sg13g2_fill_2 FILLER_22_33 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_fill_2 FILLER_22_56 ();
 sg13g2_fill_2 FILLER_22_66 ();
 sg13g2_fill_1 FILLER_22_68 ();
 sg13g2_fill_1 FILLER_22_99 ();
 sg13g2_fill_1 FILLER_22_152 ();
 sg13g2_fill_2 FILLER_22_215 ();
 sg13g2_fill_1 FILLER_22_217 ();
 sg13g2_decap_4 FILLER_22_227 ();
 sg13g2_fill_2 FILLER_22_231 ();
 sg13g2_decap_4 FILLER_22_251 ();
 sg13g2_fill_1 FILLER_22_255 ();
 sg13g2_decap_8 FILLER_22_260 ();
 sg13g2_fill_2 FILLER_22_267 ();
 sg13g2_fill_2 FILLER_22_338 ();
 sg13g2_fill_1 FILLER_22_340 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_4 ();
 sg13g2_fill_2 FILLER_23_23 ();
 sg13g2_fill_1 FILLER_23_25 ();
 sg13g2_fill_2 FILLER_23_46 ();
 sg13g2_fill_1 FILLER_23_48 ();
 sg13g2_fill_2 FILLER_23_84 ();
 sg13g2_fill_1 FILLER_23_101 ();
 sg13g2_fill_1 FILLER_23_107 ();
 sg13g2_decap_4 FILLER_23_113 ();
 sg13g2_fill_1 FILLER_23_121 ();
 sg13g2_fill_2 FILLER_23_125 ();
 sg13g2_fill_2 FILLER_23_150 ();
 sg13g2_fill_2 FILLER_23_166 ();
 sg13g2_fill_2 FILLER_23_177 ();
 sg13g2_fill_2 FILLER_23_224 ();
 sg13g2_fill_1 FILLER_23_226 ();
 sg13g2_decap_4 FILLER_23_268 ();
 sg13g2_fill_1 FILLER_23_272 ();
 sg13g2_decap_4 FILLER_23_295 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_29 ();
 sg13g2_fill_2 FILLER_24_48 ();
 sg13g2_fill_2 FILLER_24_66 ();
 sg13g2_fill_1 FILLER_24_68 ();
 sg13g2_fill_2 FILLER_24_80 ();
 sg13g2_fill_1 FILLER_24_82 ();
 sg13g2_decap_4 FILLER_24_87 ();
 sg13g2_fill_2 FILLER_24_91 ();
 sg13g2_fill_1 FILLER_24_148 ();
 sg13g2_fill_1 FILLER_24_211 ();
 sg13g2_fill_2 FILLER_24_265 ();
 sg13g2_fill_2 FILLER_24_298 ();
 sg13g2_fill_1 FILLER_24_304 ();
 sg13g2_fill_2 FILLER_24_371 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_9 ();
 sg13g2_fill_2 FILLER_25_25 ();
 sg13g2_decap_4 FILLER_25_68 ();
 sg13g2_fill_1 FILLER_25_98 ();
 sg13g2_fill_2 FILLER_25_131 ();
 sg13g2_fill_2 FILLER_25_201 ();
 sg13g2_fill_2 FILLER_25_207 ();
 sg13g2_fill_1 FILLER_25_223 ();
 sg13g2_fill_1 FILLER_25_233 ();
 sg13g2_fill_1 FILLER_25_270 ();
 sg13g2_decap_4 FILLER_25_285 ();
 sg13g2_fill_2 FILLER_25_381 ();
 sg13g2_decap_4 FILLER_26_59 ();
 sg13g2_decap_4 FILLER_26_92 ();
 sg13g2_fill_1 FILLER_26_122 ();
 sg13g2_fill_1 FILLER_26_132 ();
 sg13g2_decap_4 FILLER_26_156 ();
 sg13g2_fill_2 FILLER_26_184 ();
 sg13g2_fill_1 FILLER_26_191 ();
 sg13g2_decap_8 FILLER_26_234 ();
 sg13g2_decap_4 FILLER_26_241 ();
 sg13g2_decap_4 FILLER_26_249 ();
 sg13g2_fill_1 FILLER_26_253 ();
 sg13g2_decap_8 FILLER_26_295 ();
 sg13g2_fill_1 FILLER_26_302 ();
 sg13g2_fill_2 FILLER_26_308 ();
 sg13g2_fill_1 FILLER_26_310 ();
 sg13g2_fill_2 FILLER_26_329 ();
 sg13g2_fill_2 FILLER_26_339 ();
 sg13g2_fill_1 FILLER_26_365 ();
 sg13g2_fill_2 FILLER_26_371 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_33 ();
 sg13g2_decap_4 FILLER_27_39 ();
 sg13g2_fill_1 FILLER_27_43 ();
 sg13g2_fill_2 FILLER_27_51 ();
 sg13g2_fill_1 FILLER_27_53 ();
 sg13g2_fill_2 FILLER_27_58 ();
 sg13g2_decap_4 FILLER_27_68 ();
 sg13g2_fill_1 FILLER_27_72 ();
 sg13g2_decap_8 FILLER_27_82 ();
 sg13g2_fill_1 FILLER_27_89 ();
 sg13g2_decap_4 FILLER_27_99 ();
 sg13g2_fill_1 FILLER_27_133 ();
 sg13g2_fill_2 FILLER_27_160 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_fill_2 FILLER_27_249 ();
 sg13g2_fill_1 FILLER_27_251 ();
 sg13g2_fill_1 FILLER_27_274 ();
 sg13g2_fill_1 FILLER_27_292 ();
 sg13g2_fill_2 FILLER_27_367 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_9 ();
 sg13g2_fill_2 FILLER_28_21 ();
 sg13g2_fill_1 FILLER_28_23 ();
 sg13g2_fill_2 FILLER_28_50 ();
 sg13g2_fill_2 FILLER_28_86 ();
 sg13g2_fill_1 FILLER_28_106 ();
 sg13g2_fill_2 FILLER_28_111 ();
 sg13g2_fill_2 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_151 ();
 sg13g2_fill_1 FILLER_28_158 ();
 sg13g2_fill_2 FILLER_28_185 ();
 sg13g2_fill_1 FILLER_28_213 ();
 sg13g2_decap_8 FILLER_28_268 ();
 sg13g2_fill_1 FILLER_28_275 ();
 sg13g2_decap_8 FILLER_28_282 ();
 sg13g2_fill_2 FILLER_28_292 ();
 sg13g2_fill_1 FILLER_28_294 ();
 sg13g2_decap_8 FILLER_28_308 ();
 sg13g2_decap_8 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_322 ();
 sg13g2_fill_2 FILLER_28_350 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_44 ();
 sg13g2_fill_1 FILLER_29_109 ();
 sg13g2_fill_2 FILLER_29_114 ();
 sg13g2_fill_1 FILLER_29_116 ();
 sg13g2_fill_1 FILLER_29_156 ();
 sg13g2_fill_1 FILLER_29_163 ();
 sg13g2_fill_1 FILLER_29_205 ();
 sg13g2_fill_2 FILLER_29_226 ();
 sg13g2_fill_2 FILLER_29_232 ();
 sg13g2_decap_4 FILLER_29_244 ();
 sg13g2_fill_2 FILLER_29_261 ();
 sg13g2_fill_1 FILLER_29_263 ();
 sg13g2_decap_4 FILLER_29_303 ();
 sg13g2_fill_1 FILLER_29_397 ();
 sg13g2_fill_2 FILLER_30_56 ();
 sg13g2_fill_2 FILLER_30_235 ();
 sg13g2_fill_1 FILLER_30_237 ();
 sg13g2_decap_4 FILLER_30_274 ();
 sg13g2_fill_2 FILLER_30_278 ();
 sg13g2_fill_1 FILLER_30_284 ();
 sg13g2_fill_1 FILLER_30_311 ();
 sg13g2_fill_2 FILLER_30_347 ();
 sg13g2_fill_2 FILLER_30_355 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_24 ();
 sg13g2_fill_1 FILLER_31_56 ();
 sg13g2_fill_2 FILLER_31_92 ();
 sg13g2_fill_2 FILLER_31_125 ();
 sg13g2_fill_2 FILLER_31_188 ();
 sg13g2_fill_1 FILLER_31_190 ();
 sg13g2_decap_8 FILLER_31_215 ();
 sg13g2_fill_1 FILLER_31_222 ();
 sg13g2_decap_8 FILLER_31_227 ();
 sg13g2_fill_1 FILLER_31_334 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_4 ();
 sg13g2_fill_2 FILLER_32_116 ();
 sg13g2_fill_2 FILLER_32_142 ();
 sg13g2_fill_2 FILLER_32_207 ();
 sg13g2_fill_1 FILLER_32_272 ();
 sg13g2_fill_1 FILLER_32_351 ();
 sg13g2_fill_1 FILLER_32_368 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_14 ();
 sg13g2_fill_2 FILLER_33_96 ();
 sg13g2_fill_2 FILLER_33_108 ();
 sg13g2_fill_2 FILLER_33_130 ();
 sg13g2_fill_2 FILLER_33_225 ();
 sg13g2_decap_4 FILLER_33_235 ();
 sg13g2_fill_2 FILLER_33_305 ();
 sg13g2_fill_1 FILLER_33_319 ();
 sg13g2_fill_2 FILLER_33_356 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_4 ();
 sg13g2_fill_2 FILLER_34_18 ();
 sg13g2_fill_1 FILLER_34_20 ();
 sg13g2_fill_2 FILLER_34_80 ();
 sg13g2_fill_1 FILLER_34_185 ();
 sg13g2_fill_1 FILLER_34_200 ();
 sg13g2_fill_1 FILLER_34_285 ();
 sg13g2_fill_2 FILLER_34_298 ();
 sg13g2_fill_1 FILLER_34_300 ();
 sg13g2_fill_1 FILLER_34_371 ();
 sg13g2_fill_2 FILLER_34_381 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_fill_2 FILLER_35_43 ();
 sg13g2_fill_1 FILLER_35_164 ();
 sg13g2_fill_2 FILLER_35_327 ();
 sg13g2_fill_1 FILLER_36_28 ();
 sg13g2_fill_2 FILLER_36_67 ();
 sg13g2_fill_1 FILLER_36_100 ();
 sg13g2_fill_1 FILLER_36_110 ();
 sg13g2_fill_2 FILLER_36_132 ();
 sg13g2_fill_1 FILLER_36_197 ();
 sg13g2_fill_2 FILLER_36_267 ();
 sg13g2_fill_2 FILLER_36_316 ();
 sg13g2_fill_2 FILLER_36_350 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_57 ();
 sg13g2_fill_2 FILLER_37_83 ();
 sg13g2_fill_2 FILLER_37_151 ();
 sg13g2_fill_1 FILLER_37_167 ();
 sg13g2_fill_2 FILLER_37_177 ();
 sg13g2_fill_1 FILLER_37_261 ();
 sg13g2_fill_2 FILLER_37_333 ();
 sg13g2_fill_1 FILLER_37_335 ();
 sg13g2_fill_2 FILLER_37_388 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_2 ();
 sg13g2_fill_2 FILLER_38_36 ();
 sg13g2_fill_1 FILLER_38_64 ();
 sg13g2_fill_1 FILLER_38_137 ();
 sg13g2_fill_2 FILLER_38_143 ();
 sg13g2_fill_1 FILLER_38_189 ();
 sg13g2_fill_1 FILLER_38_202 ();
 sg13g2_fill_1 FILLER_38_242 ();
 sg13g2_fill_2 FILLER_38_272 ();
 sg13g2_fill_1 FILLER_38_274 ();
 sg13g2_fill_2 FILLER_38_293 ();
 sg13g2_fill_1 FILLER_38_320 ();
 sg13g2_fill_1 FILLER_38_359 ();
 sg13g2_fill_1 FILLER_38_377 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net18;
 assign uio_oe[1] = net19;
 assign uio_oe[2] = net20;
 assign uio_oe[3] = net21;
 assign uio_oe[4] = net22;
 assign uio_oe[5] = net23;
 assign uio_oe[6] = net24;
 assign uio_oe[7] = net25;
 assign uio_out[0] = net26;
 assign uio_out[1] = net27;
 assign uio_out[2] = net28;
 assign uio_out[3] = net29;
 assign uio_out[4] = net30;
 assign uio_out[5] = net31;
 assign uio_out[6] = net32;
 assign uio_out[7] = net33;
endmodule

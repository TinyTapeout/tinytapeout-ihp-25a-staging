module tt_um_monishvr_fifo (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire clknet_0_clk;
 wire dffr1;
 wire dffr2;
 wire dffw1;
 wire dffw2;
 wire empty;
 wire full;
 wire \rd_next[0] ;
 wire \rd_reg[0] ;
 wire \rd_reg[1] ;
 wire \rd_reg[2] ;
 wire \regarray[0][0] ;
 wire \regarray[0][1] ;
 wire \regarray[0][2] ;
 wire \regarray[0][3] ;
 wire \regarray[1][0] ;
 wire \regarray[1][1] ;
 wire \regarray[1][2] ;
 wire \regarray[1][3] ;
 wire \regarray[2][0] ;
 wire \regarray[2][1] ;
 wire \regarray[2][2] ;
 wire \regarray[2][3] ;
 wire \regarray[3][0] ;
 wire \regarray[3][1] ;
 wire \regarray[3][2] ;
 wire \regarray[3][3] ;
 wire \regarray[4][0] ;
 wire \regarray[4][1] ;
 wire \regarray[4][2] ;
 wire \regarray[4][3] ;
 wire \regarray[5][0] ;
 wire \regarray[5][1] ;
 wire \regarray[5][2] ;
 wire \regarray[5][3] ;
 wire \regarray[6][0] ;
 wire \regarray[6][1] ;
 wire \regarray[6][2] ;
 wire \regarray[6][3] ;
 wire \regarray[7][0] ;
 wire \regarray[7][1] ;
 wire \regarray[7][2] ;
 wire \regarray[7][3] ;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire \wr_next[0] ;
 wire \wr_reg[0] ;
 wire \wr_reg[1] ;
 wire \wr_reg[2] ;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;

 sg13g2_nor2_1 _236_ (.A(net44),
    .B(net107),
    .Y(_116_));
 sg13g2_nor3_2 _237_ (.A(net38),
    .B(_115_),
    .C(_116_),
    .Y(_117_));
 sg13g2_nor2b_1 _238_ (.A(net94),
    .B_N(net40),
    .Y(_118_));
 sg13g2_o21ai_1 _239_ (.B1(net36),
    .Y(_119_),
    .A1(net40),
    .A2(\regarray[6][1] ));
 sg13g2_o21ai_1 _240_ (.B1(net35),
    .Y(_120_),
    .A1(_118_),
    .A2(_119_));
 sg13g2_or2_1 _241_ (.X(_121_),
    .B(\regarray[0][1] ),
    .A(net41));
 sg13g2_a21oi_1 _242_ (.A1(net41),
    .A2(_058_),
    .Y(_122_),
    .B1(net38));
 sg13g2_mux2_1 _243_ (.A0(\regarray[2][1] ),
    .A1(\regarray[3][1] ),
    .S(net39),
    .X(_123_));
 sg13g2_a221oi_1 _244_ (.B2(net36),
    .C1(net35),
    .B1(_123_),
    .A1(_121_),
    .Y(_124_),
    .A2(_122_));
 sg13g2_o21ai_1 _245_ (.B1(_065_),
    .Y(_125_),
    .A1(_117_),
    .A2(_120_));
 sg13g2_o21ai_1 _246_ (.B1(_114_),
    .Y(_035_),
    .A1(_124_),
    .A2(_125_));
 sg13g2_nand2_1 _247_ (.Y(_126_),
    .A(net131),
    .B(_066_));
 sg13g2_nor2b_1 _248_ (.A(\regarray[5][2] ),
    .B_N(net42),
    .Y(_127_));
 sg13g2_nor2_1 _249_ (.A(net44),
    .B(\regarray[4][2] ),
    .Y(_128_));
 sg13g2_nor3_2 _250_ (.A(net38),
    .B(_127_),
    .C(_128_),
    .Y(_129_));
 sg13g2_nor2b_1 _251_ (.A(net90),
    .B_N(net40),
    .Y(_130_));
 sg13g2_o21ai_1 _252_ (.B1(net36),
    .Y(_131_),
    .A1(net40),
    .A2(\regarray[6][2] ));
 sg13g2_o21ai_1 _253_ (.B1(net35),
    .Y(_132_),
    .A1(_130_),
    .A2(_131_));
 sg13g2_or2_1 _254_ (.X(_133_),
    .B(\regarray[0][2] ),
    .A(net39));
 sg13g2_a21oi_1 _255_ (.A1(net39),
    .A2(_059_),
    .Y(_134_),
    .B1(net36));
 sg13g2_mux2_1 _256_ (.A0(\regarray[2][2] ),
    .A1(\regarray[3][2] ),
    .S(net39),
    .X(_135_));
 sg13g2_a221oi_1 _257_ (.B2(net36),
    .C1(net35),
    .B1(_135_),
    .A1(_133_),
    .Y(_136_),
    .A2(_134_));
 sg13g2_o21ai_1 _258_ (.B1(_065_),
    .Y(_137_),
    .A1(_129_),
    .A2(_132_));
 sg13g2_o21ai_1 _259_ (.B1(_126_),
    .Y(_036_),
    .A1(_136_),
    .A2(_137_));
 sg13g2_nand2_1 _260_ (.Y(_138_),
    .A(net133),
    .B(_066_));
 sg13g2_or2_1 _261_ (.X(_139_),
    .B(\regarray[0][3] ),
    .A(net39));
 sg13g2_a21oi_1 _262_ (.A1(net39),
    .A2(_060_),
    .Y(_140_),
    .B1(net36));
 sg13g2_mux2_1 _263_ (.A0(\regarray[2][3] ),
    .A1(\regarray[3][3] ),
    .S(net39),
    .X(_141_));
 sg13g2_a221oi_1 _264_ (.B2(net36),
    .C1(net35),
    .B1(_141_),
    .A1(_139_),
    .Y(_142_),
    .A2(_140_));
 sg13g2_nor2b_1 _265_ (.A(\regarray[5][3] ),
    .B_N(net42),
    .Y(_143_));
 sg13g2_nor2_1 _266_ (.A(net42),
    .B(net95),
    .Y(_144_));
 sg13g2_nor3_2 _267_ (.A(net37),
    .B(_143_),
    .C(_144_),
    .Y(_145_));
 sg13g2_nor2b_1 _268_ (.A(net112),
    .B_N(net40),
    .Y(_146_));
 sg13g2_o21ai_1 _269_ (.B1(net36),
    .Y(_147_),
    .A1(net39),
    .A2(\regarray[6][3] ));
 sg13g2_o21ai_1 _270_ (.B1(net35),
    .Y(_148_),
    .A1(_146_),
    .A2(_147_));
 sg13g2_o21ai_1 _271_ (.B1(_065_),
    .Y(_149_),
    .A1(_145_),
    .A2(_148_));
 sg13g2_o21ai_1 _272_ (.B1(_138_),
    .Y(_037_),
    .A1(_142_),
    .A2(_149_));
 sg13g2_nor4_2 _273_ (.A(net45),
    .B(_055_),
    .C(net149),
    .Y(_150_),
    .D(net34));
 sg13g2_mux2_1 _274_ (.A0(net115),
    .A1(net4),
    .S(_150_),
    .X(_038_));
 sg13g2_mux2_1 _275_ (.A0(net108),
    .A1(net5),
    .S(_150_),
    .X(_039_));
 sg13g2_mux2_1 _276_ (.A0(net120),
    .A1(net6),
    .S(_150_),
    .X(_040_));
 sg13g2_mux2_1 _277_ (.A0(net116),
    .A1(net7),
    .S(_150_),
    .X(_041_));
 sg13g2_nor4_2 _278_ (.A(net45),
    .B(_055_),
    .C(\wr_reg[0] ),
    .Y(_151_),
    .D(net34));
 sg13g2_mux2_1 _279_ (.A0(net85),
    .A1(net4),
    .S(_151_),
    .X(_042_));
 sg13g2_mux2_1 _280_ (.A0(net86),
    .A1(net5),
    .S(_151_),
    .X(_043_));
 sg13g2_mux2_1 _281_ (.A0(net87),
    .A1(net6),
    .S(_151_),
    .X(_044_));
 sg13g2_mux2_1 _282_ (.A0(net88),
    .A1(net7),
    .S(_151_),
    .X(_045_));
 sg13g2_inv_1 _283_ (.Y(_003_),
    .A(net1));
 sg13g2_inv_1 _284_ (.Y(_004_),
    .A(net1));
 sg13g2_inv_1 _285_ (.Y(_005_),
    .A(net1));
 sg13g2_inv_1 _286_ (.Y(_006_),
    .A(net1));
 sg13g2_inv_1 _287_ (.Y(_007_),
    .A(net1));
 sg13g2_inv_1 _288_ (.Y(_008_),
    .A(net1));
 sg13g2_inv_1 _289_ (.Y(_009_),
    .A(net1));
 sg13g2_inv_1 _290_ (.Y(_054_),
    .A(net45));
 sg13g2_inv_1 _291_ (.Y(_055_),
    .A(\wr_reg[1] ));
 sg13g2_inv_1 _292_ (.Y(_056_),
    .A(\wr_reg[0] ));
 sg13g2_inv_1 _293_ (.Y(_057_),
    .A(net110));
 sg13g2_inv_1 _294_ (.Y(_058_),
    .A(net101));
 sg13g2_inv_1 _295_ (.Y(_059_),
    .A(net129));
 sg13g2_inv_1 _296_ (.Y(_060_),
    .A(net127));
 sg13g2_inv_1 _297_ (.Y(_002_),
    .A(net1));
 sg13g2_nor2b_1 _298_ (.A(net79),
    .B_N(dffw2),
    .Y(_061_));
 sg13g2_nand2b_2 _299_ (.Y(_062_),
    .B(dffw2),
    .A_N(net79));
 sg13g2_nor2b_2 _300_ (.A(net78),
    .B_N(dffr2),
    .Y(_063_));
 sg13g2_nand2b_2 _301_ (.Y(_064_),
    .B(net146),
    .A_N(net78));
 sg13g2_nor2_2 _302_ (.A(empty),
    .B(_064_),
    .Y(_065_));
 sg13g2_nand2b_2 _303_ (.Y(_066_),
    .B(_063_),
    .A_N(empty));
 sg13g2_nand2_1 _304_ (.Y(_067_),
    .A(_062_),
    .B(_063_));
 sg13g2_nand2_1 _305_ (.Y(_068_),
    .A(_062_),
    .B(_065_));
 sg13g2_xnor2_1 _306_ (.Y(_069_),
    .A(net37),
    .B(\wr_reg[1] ));
 sg13g2_nand2b_1 _307_ (.Y(_070_),
    .B(net43),
    .A_N(\wr_reg[0] ));
 sg13g2_nand2b_1 _308_ (.Y(_071_),
    .B(\wr_reg[0] ),
    .A_N(net43));
 sg13g2_mux2_1 _309_ (.A0(_070_),
    .A1(_071_),
    .S(_069_),
    .X(_072_));
 sg13g2_a21o_1 _310_ (.A2(net42),
    .A1(net37),
    .B1(net35),
    .X(_073_));
 sg13g2_nand3_1 _311_ (.B(net37),
    .C(net43),
    .A(net35),
    .Y(_074_));
 sg13g2_nand3_1 _312_ (.B(_073_),
    .C(_074_),
    .A(net45),
    .Y(_075_));
 sg13g2_a21o_1 _313_ (.A2(_074_),
    .A1(_073_),
    .B1(\wr_reg[2] ),
    .X(_076_));
 sg13g2_a21oi_1 _314_ (.A1(_075_),
    .A2(_076_),
    .Y(_077_),
    .B1(_072_));
 sg13g2_nand3b_1 _315_ (.B(dffw2),
    .C(_000_),
    .Y(_078_),
    .A_N(dffw1));
 sg13g2_nor2_1 _316_ (.A(_063_),
    .B(net34),
    .Y(_079_));
 sg13g2_o21ai_1 _317_ (.B1(_067_),
    .Y(_080_),
    .A1(net135),
    .A2(_079_));
 sg13g2_o21ai_1 _318_ (.B1(net136),
    .Y(_053_),
    .A1(_068_),
    .A2(_077_));
 sg13g2_nand2_1 _319_ (.Y(_081_),
    .A(net45),
    .B(\wr_reg[1] ));
 sg13g2_nand2b_1 _320_ (.Y(_082_),
    .B(_056_),
    .A_N(_081_));
 sg13g2_a21oi_1 _321_ (.A1(_061_),
    .A2(_064_),
    .Y(_083_),
    .B1(net82));
 sg13g2_a221oi_1 _322_ (.B2(_082_),
    .C1(net83),
    .B1(_079_),
    .A1(_062_),
    .Y(_052_),
    .A2(_065_));
 sg13g2_a21oi_2 _323_ (.B1(_064_),
    .Y(_084_),
    .A2(_062_),
    .A1(empty));
 sg13g2_a221oi_1 _324_ (.B2(_074_),
    .C1(_064_),
    .B1(_073_),
    .A1(empty),
    .Y(_085_),
    .A2(_062_));
 sg13g2_nor2_1 _325_ (.A(net138),
    .B(_084_),
    .Y(_086_));
 sg13g2_nor2_1 _326_ (.A(_085_),
    .B(net139),
    .Y(_051_));
 sg13g2_nand2_1 _327_ (.Y(_087_),
    .A(net42),
    .B(net147));
 sg13g2_xnor2_1 _328_ (.Y(_050_),
    .A(net37),
    .B(_087_));
 sg13g2_mux2_1 _329_ (.A0(net42),
    .A1(net80),
    .S(_084_),
    .X(_049_));
 sg13g2_o21ai_1 _330_ (.B1(_061_),
    .Y(_088_),
    .A1(_000_),
    .A2(_063_));
 sg13g2_nand3b_1 _331_ (.B(\wr_reg[0] ),
    .C(\wr_reg[1] ),
    .Y(_089_),
    .A_N(_088_));
 sg13g2_xnor2_1 _332_ (.Y(_048_),
    .A(net45),
    .B(_089_));
 sg13g2_o21ai_1 _333_ (.B1(_055_),
    .Y(_090_),
    .A1(_056_),
    .A2(_088_));
 sg13g2_and2_1 _334_ (.A(_089_),
    .B(_090_),
    .X(_047_));
 sg13g2_nor2_1 _335_ (.A(net141),
    .B(_088_),
    .Y(_091_));
 sg13g2_a21oi_1 _336_ (.A1(_056_),
    .A2(_088_),
    .Y(_046_),
    .B1(net142));
 sg13g2_nor2_2 _337_ (.A(_078_),
    .B(_082_),
    .Y(_092_));
 sg13g2_mux2_1 _338_ (.A0(net105),
    .A1(net4),
    .S(_092_),
    .X(_010_));
 sg13g2_mux2_1 _339_ (.A0(net98),
    .A1(net5),
    .S(_092_),
    .X(_011_));
 sg13g2_mux2_1 _340_ (.A0(net113),
    .A1(net6),
    .S(_092_),
    .X(_012_));
 sg13g2_mux2_1 _341_ (.A0(net103),
    .A1(net7),
    .S(_092_),
    .X(_013_));
 sg13g2_nor4_2 _342_ (.A(net45),
    .B(\wr_reg[1] ),
    .C(\wr_reg[0] ),
    .Y(_093_),
    .D(net34));
 sg13g2_mux2_1 _343_ (.A0(net96),
    .A1(net4),
    .S(_093_),
    .X(_014_));
 sg13g2_mux2_1 _344_ (.A0(net89),
    .A1(net5),
    .S(_093_),
    .X(_015_));
 sg13g2_mux2_1 _345_ (.A0(net92),
    .A1(net6),
    .S(_093_),
    .X(_016_));
 sg13g2_mux2_1 _346_ (.A0(net91),
    .A1(net7),
    .S(_093_),
    .X(_017_));
 sg13g2_nor3_2 _347_ (.A(net148),
    .B(net34),
    .C(_081_),
    .Y(_094_));
 sg13g2_mux2_1 _348_ (.A0(net97),
    .A1(net4),
    .S(_094_),
    .X(_018_));
 sg13g2_mux2_1 _349_ (.A0(net94),
    .A1(net5),
    .S(_094_),
    .X(_019_));
 sg13g2_mux2_1 _350_ (.A0(net90),
    .A1(net6),
    .S(_094_),
    .X(_020_));
 sg13g2_mux2_1 _351_ (.A0(net112),
    .A1(net7),
    .S(_094_),
    .X(_021_));
 sg13g2_nor4_2 _352_ (.A(net45),
    .B(\wr_reg[1] ),
    .C(\wr_next[0] ),
    .Y(_095_),
    .D(net34));
 sg13g2_nand2_1 _353_ (.Y(_096_),
    .A(net4),
    .B(_095_));
 sg13g2_o21ai_1 _354_ (.B1(_096_),
    .Y(_022_),
    .A1(_057_),
    .A2(_095_));
 sg13g2_nand2_1 _355_ (.Y(_097_),
    .A(net5),
    .B(_095_));
 sg13g2_o21ai_1 _356_ (.B1(_097_),
    .Y(_023_),
    .A1(_058_),
    .A2(_095_));
 sg13g2_nand2_1 _357_ (.Y(_098_),
    .A(net6),
    .B(_095_));
 sg13g2_o21ai_1 _358_ (.B1(_098_),
    .Y(_024_),
    .A1(_059_),
    .A2(_095_));
 sg13g2_nand2_1 _359_ (.Y(_099_),
    .A(net7),
    .B(_095_));
 sg13g2_o21ai_1 _360_ (.B1(_099_),
    .Y(_025_),
    .A1(_060_),
    .A2(_095_));
 sg13g2_nor4_2 _361_ (.A(_054_),
    .B(\wr_reg[1] ),
    .C(net148),
    .Y(_100_),
    .D(net34));
 sg13g2_mux2_1 _362_ (.A0(net100),
    .A1(net4),
    .S(_100_),
    .X(_026_));
 sg13g2_mux2_1 _363_ (.A0(net117),
    .A1(net5),
    .S(_100_),
    .X(_027_));
 sg13g2_mux2_1 _364_ (.A0(net118),
    .A1(net6),
    .S(_100_),
    .X(_028_));
 sg13g2_mux2_1 _365_ (.A0(net123),
    .A1(net7),
    .S(_100_),
    .X(_029_));
 sg13g2_nor4_2 _366_ (.A(_054_),
    .B(\wr_reg[1] ),
    .C(\wr_reg[0] ),
    .Y(_101_),
    .D(net34));
 sg13g2_mux2_1 _367_ (.A0(net109),
    .A1(net4),
    .S(_101_),
    .X(_030_));
 sg13g2_mux2_1 _368_ (.A0(net107),
    .A1(net5),
    .S(_101_),
    .X(_031_));
 sg13g2_mux2_1 _369_ (.A0(net93),
    .A1(net6),
    .S(_101_),
    .X(_032_));
 sg13g2_mux2_1 _370_ (.A0(net95),
    .A1(net7),
    .S(_101_),
    .X(_033_));
 sg13g2_nand2_1 _371_ (.Y(_102_),
    .A(net125),
    .B(_066_));
 sg13g2_nor2b_1 _372_ (.A(net100),
    .B_N(net43),
    .Y(_103_));
 sg13g2_nor2_1 _373_ (.A(net42),
    .B(net109),
    .Y(_104_));
 sg13g2_nor3_1 _374_ (.A(net37),
    .B(_103_),
    .C(_104_),
    .Y(_105_));
 sg13g2_nor2b_1 _375_ (.A(\regarray[7][0] ),
    .B_N(net41),
    .Y(_106_));
 sg13g2_o21ai_1 _376_ (.B1(net38),
    .Y(_107_),
    .A1(net41),
    .A2(\regarray[6][0] ));
 sg13g2_o21ai_1 _377_ (.B1(\rd_reg[2] ),
    .Y(_108_),
    .A1(_106_),
    .A2(_107_));
 sg13g2_or2_1 _378_ (.X(_109_),
    .B(\regarray[0][0] ),
    .A(net43));
 sg13g2_a21oi_1 _379_ (.A1(net43),
    .A2(_057_),
    .Y(_110_),
    .B1(net37));
 sg13g2_mux2_1 _380_ (.A0(\regarray[2][0] ),
    .A1(\regarray[3][0] ),
    .S(net43),
    .X(_111_));
 sg13g2_a221oi_1 _381_ (.B2(net37),
    .C1(\rd_reg[2] ),
    .B1(_111_),
    .A1(_109_),
    .Y(_112_),
    .A2(_110_));
 sg13g2_o21ai_1 _382_ (.B1(_065_),
    .Y(_113_),
    .A1(_105_),
    .A2(_108_));
 sg13g2_o21ai_1 _383_ (.B1(_102_),
    .Y(_034_),
    .A1(_112_),
    .A2(_113_));
 sg13g2_nand2_1 _384_ (.Y(_114_),
    .A(net121),
    .B(_066_));
 sg13g2_nor2b_1 _385_ (.A(\regarray[5][1] ),
    .B_N(net42),
    .Y(_115_));
 sg13g2_dfrbp_1 _386_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net75),
    .D(net106),
    .Q_N(_192_),
    .Q(\regarray[6][0] ));
 sg13g2_dfrbp_1 _387_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net32),
    .D(net99),
    .Q_N(_191_),
    .Q(\regarray[6][1] ));
 sg13g2_dfrbp_1 _388_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net31),
    .D(net114),
    .Q_N(_190_),
    .Q(\regarray[6][2] ));
 sg13g2_dfrbp_1 _389_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net30),
    .D(net104),
    .Q_N(_189_),
    .Q(\regarray[6][3] ));
 sg13g2_dfrbp_1 _390_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net29),
    .D(_014_),
    .Q_N(_188_),
    .Q(\regarray[0][0] ));
 sg13g2_dfrbp_1 _391_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net28),
    .D(_015_),
    .Q_N(_187_),
    .Q(\regarray[0][1] ));
 sg13g2_dfrbp_1 _392_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net27),
    .D(_016_),
    .Q_N(_186_),
    .Q(\regarray[0][2] ));
 sg13g2_dfrbp_1 _393_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net26),
    .D(_017_),
    .Q_N(_185_),
    .Q(\regarray[0][3] ));
 sg13g2_dfrbp_1 _394_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net74),
    .D(_018_),
    .Q_N(_184_),
    .Q(\regarray[7][0] ));
 sg13g2_dfrbp_1 _395_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net73),
    .D(_019_),
    .Q_N(_183_),
    .Q(\regarray[7][1] ));
 sg13g2_dfrbp_1 _396_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net72),
    .D(_020_),
    .Q_N(_182_),
    .Q(\regarray[7][2] ));
 sg13g2_dfrbp_1 _397_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net71),
    .D(_021_),
    .Q_N(_181_),
    .Q(\regarray[7][3] ));
 sg13g2_dfrbp_1 _398_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net70),
    .D(net111),
    .Q_N(_180_),
    .Q(\regarray[1][0] ));
 sg13g2_dfrbp_1 _399_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net69),
    .D(net102),
    .Q_N(_179_),
    .Q(\regarray[1][1] ));
 sg13g2_dfrbp_1 _400_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net68),
    .D(net130),
    .Q_N(_178_),
    .Q(\regarray[1][2] ));
 sg13g2_dfrbp_1 _401_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net67),
    .D(net128),
    .Q_N(_177_),
    .Q(\regarray[1][3] ));
 sg13g2_dfrbp_1 _402_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net66),
    .D(_026_),
    .Q_N(_176_),
    .Q(\regarray[5][0] ));
 sg13g2_dfrbp_1 _403_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net65),
    .D(_027_),
    .Q_N(_175_),
    .Q(\regarray[5][1] ));
 sg13g2_dfrbp_1 _404_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net64),
    .D(net119),
    .Q_N(_174_),
    .Q(\regarray[5][2] ));
 sg13g2_dfrbp_1 _405_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net63),
    .D(net124),
    .Q_N(_173_),
    .Q(\regarray[5][3] ));
 sg13g2_dfrbp_1 _406_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net62),
    .D(_030_),
    .Q_N(_172_),
    .Q(\regarray[4][0] ));
 sg13g2_dfrbp_1 _407_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net61),
    .D(_031_),
    .Q_N(_171_),
    .Q(\regarray[4][1] ));
 sg13g2_dfrbp_1 _408_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net60),
    .D(_032_),
    .Q_N(_170_),
    .Q(\regarray[4][2] ));
 sg13g2_dfrbp_1 _409_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net59),
    .D(_033_),
    .Q_N(_169_),
    .Q(\regarray[4][3] ));
 sg13g2_dfrbp_1 _410_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net58),
    .D(net126),
    .Q_N(_168_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _411_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net57),
    .D(net122),
    .Q_N(_167_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _412_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net56),
    .D(net132),
    .Q_N(_166_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _413_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net55),
    .D(net134),
    .Q_N(_165_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _414_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net54),
    .D(_038_),
    .Q_N(_164_),
    .Q(\regarray[3][0] ));
 sg13g2_dfrbp_1 _415_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net53),
    .D(_039_),
    .Q_N(_163_),
    .Q(\regarray[3][1] ));
 sg13g2_dfrbp_1 _416_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net52),
    .D(_040_),
    .Q_N(_162_),
    .Q(\regarray[3][2] ));
 sg13g2_dfrbp_1 _417_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net51),
    .D(_041_),
    .Q_N(_161_),
    .Q(\regarray[3][3] ));
 sg13g2_dfrbp_1 _418_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net50),
    .D(_042_),
    .Q_N(_160_),
    .Q(\regarray[2][0] ));
 sg13g2_dfrbp_1 _419_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net49),
    .D(_043_),
    .Q_N(_159_),
    .Q(\regarray[2][1] ));
 sg13g2_dfrbp_1 _420_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net48),
    .D(_044_),
    .Q_N(_158_),
    .Q(\regarray[2][2] ));
 sg13g2_dfrbp_1 _421_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net47),
    .D(_045_),
    .Q_N(_157_),
    .Q(\regarray[2][3] ));
 sg13g2_dfrbp_1 _422_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(_002_),
    .D(net143),
    .Q_N(\wr_next[0] ),
    .Q(\wr_reg[0] ));
 sg13g2_dfrbp_1 _423_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(_003_),
    .D(_047_),
    .Q_N(_156_),
    .Q(\wr_reg[1] ));
 sg13g2_dfrbp_1 _424_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(_004_),
    .D(net145),
    .Q_N(_155_),
    .Q(\wr_reg[2] ));
 sg13g2_dfrbp_1 _425_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(_005_),
    .D(net81),
    .Q_N(\rd_next[0] ),
    .Q(\rd_reg[0] ));
 sg13g2_dfrbp_1 _426_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(_006_),
    .D(_050_),
    .Q_N(_154_),
    .Q(\rd_reg[1] ));
 sg13g2_dfrbp_1 _427_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(_007_),
    .D(net140),
    .Q_N(_153_),
    .Q(\rd_reg[2] ));
 sg13g2_dfrbp_1 _428_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(_008_),
    .D(net84),
    .Q_N(_000_),
    .Q(full));
 sg13g2_dfrbp_1 _429_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(_009_),
    .D(net137),
    .Q_N(empty),
    .Q(_001_));
 sg13g2_dfrbp_1 _430_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net76),
    .D(net78),
    .Q_N(_193_),
    .Q(dffr2));
 sg13g2_dfrbp_1 _431_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net77),
    .D(net3),
    .Q_N(_194_),
    .Q(dffr1));
 sg13g2_dfrbp_1 _432_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net46),
    .D(net79),
    .Q_N(_195_),
    .Q(dffw2));
 sg13g2_dfrbp_1 _433_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net33),
    .D(net2),
    .Q_N(_152_),
    .Q(dffw1));
 sg13g2_tiehi _392__27 (.L_HI(net27));
 sg13g2_tiehi _391__28 (.L_HI(net28));
 sg13g2_tiehi _390__29 (.L_HI(net29));
 sg13g2_tiehi _389__30 (.L_HI(net30));
 sg13g2_tiehi _388__31 (.L_HI(net31));
 sg13g2_tiehi _387__32 (.L_HI(net32));
 sg13g2_tiehi _433__33 (.L_HI(net33));
 sg13g2_tiehi _432__34 (.L_HI(net46));
 sg13g2_tiehi _421__35 (.L_HI(net47));
 sg13g2_tiehi _420__36 (.L_HI(net48));
 sg13g2_tiehi _419__37 (.L_HI(net49));
 sg13g2_tiehi _418__38 (.L_HI(net50));
 sg13g2_tiehi _417__39 (.L_HI(net51));
 sg13g2_tiehi _416__40 (.L_HI(net52));
 sg13g2_tiehi _415__41 (.L_HI(net53));
 sg13g2_tiehi _414__42 (.L_HI(net54));
 sg13g2_tiehi _413__43 (.L_HI(net55));
 sg13g2_tiehi _412__44 (.L_HI(net56));
 sg13g2_tiehi _411__45 (.L_HI(net57));
 sg13g2_tiehi _410__46 (.L_HI(net58));
 sg13g2_tiehi _409__47 (.L_HI(net59));
 sg13g2_tiehi _408__48 (.L_HI(net60));
 sg13g2_tiehi _407__49 (.L_HI(net61));
 sg13g2_tiehi _406__50 (.L_HI(net62));
 sg13g2_tiehi _405__51 (.L_HI(net63));
 sg13g2_tiehi _404__52 (.L_HI(net64));
 sg13g2_tiehi _403__53 (.L_HI(net65));
 sg13g2_tiehi _402__54 (.L_HI(net66));
 sg13g2_tiehi _401__55 (.L_HI(net67));
 sg13g2_tiehi _400__56 (.L_HI(net68));
 sg13g2_tiehi _399__57 (.L_HI(net69));
 sg13g2_tiehi _398__58 (.L_HI(net70));
 sg13g2_tiehi _397__59 (.L_HI(net71));
 sg13g2_tiehi _396__60 (.L_HI(net72));
 sg13g2_tiehi _395__61 (.L_HI(net73));
 sg13g2_tiehi _394__62 (.L_HI(net74));
 sg13g2_tiehi _386__63 (.L_HI(net75));
 sg13g2_tiehi _430__64 (.L_HI(net76));
 sg13g2_tiehi _431__65 (.L_HI(net77));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_monishvr_fifo_9 (.L_LO(net9));
 sg13g2_tielo tt_um_monishvr_fifo_10 (.L_LO(net10));
 sg13g2_tielo tt_um_monishvr_fifo_11 (.L_LO(net11));
 sg13g2_tielo tt_um_monishvr_fifo_12 (.L_LO(net12));
 sg13g2_tielo tt_um_monishvr_fifo_13 (.L_LO(net13));
 sg13g2_tielo tt_um_monishvr_fifo_14 (.L_LO(net14));
 sg13g2_tielo tt_um_monishvr_fifo_15 (.L_LO(net15));
 sg13g2_tielo tt_um_monishvr_fifo_16 (.L_LO(net16));
 sg13g2_tielo tt_um_monishvr_fifo_17 (.L_LO(net17));
 sg13g2_tielo tt_um_monishvr_fifo_18 (.L_LO(net18));
 sg13g2_tielo tt_um_monishvr_fifo_19 (.L_LO(net19));
 sg13g2_tielo tt_um_monishvr_fifo_20 (.L_LO(net20));
 sg13g2_tielo tt_um_monishvr_fifo_21 (.L_LO(net21));
 sg13g2_tielo tt_um_monishvr_fifo_22 (.L_LO(net22));
 sg13g2_tielo tt_um_monishvr_fifo_23 (.L_LO(net23));
 sg13g2_tielo tt_um_monishvr_fifo_24 (.L_LO(net24));
 sg13g2_tielo tt_um_monishvr_fifo_25 (.L_LO(net25));
 sg13g2_tiehi _393__26 (.L_HI(net26));
 sg13g2_buf_1 _492_ (.A(full),
    .X(uo_out[0]));
 sg13g2_buf_1 _493_ (.A(empty),
    .X(uo_out[1]));
 sg13g2_buf_4 fanout34 (.X(net34),
    .A(_078_));
 sg13g2_buf_2 fanout35 (.A(\rd_reg[2] ),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(net38),
    .X(net36));
 sg13g2_buf_4 fanout37 (.X(net37),
    .A(net38));
 sg13g2_buf_2 fanout38 (.A(\rd_reg[1] ),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(net41),
    .X(net39));
 sg13g2_buf_1 fanout40 (.A(net41),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(net44),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(net43),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(net44),
    .X(net43));
 sg13g2_buf_1 fanout44 (.A(\rd_reg[0] ),
    .X(net44));
 sg13g2_buf_4 fanout45 (.X(net45),
    .A(net144));
 sg13g2_buf_4 input1 (.X(net1),
    .A(rst_n));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[4]));
 sg13g2_buf_4 input5 (.X(net5),
    .A(ui_in[5]));
 sg13g2_buf_4 input6 (.X(net6),
    .A(ui_in[6]));
 sg13g2_buf_4 input7 (.X(net7),
    .A(ui_in[7]));
 sg13g2_tielo tt_um_monishvr_fifo_8 (.L_LO(net8));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(dffr1),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold2 (.A(dffw1),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold3 (.A(\rd_next[0] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold4 (.A(_049_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold5 (.A(full),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold6 (.A(_083_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold7 (.A(_052_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold8 (.A(\regarray[2][0] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold9 (.A(\regarray[2][1] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold10 (.A(\regarray[2][2] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold11 (.A(\regarray[2][3] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold12 (.A(\regarray[0][1] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold13 (.A(\regarray[7][2] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold14 (.A(\regarray[0][3] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold15 (.A(\regarray[0][2] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold16 (.A(\regarray[4][2] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold17 (.A(\regarray[7][1] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold18 (.A(\regarray[4][3] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold19 (.A(\regarray[0][0] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold20 (.A(\regarray[7][0] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold21 (.A(\regarray[6][1] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold22 (.A(_011_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold23 (.A(\regarray[5][0] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold24 (.A(\regarray[1][1] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold25 (.A(_023_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold26 (.A(\regarray[6][3] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold27 (.A(_013_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold28 (.A(\regarray[6][0] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold29 (.A(_010_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold30 (.A(\regarray[4][1] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold31 (.A(\regarray[3][1] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold32 (.A(\regarray[4][0] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold33 (.A(\regarray[1][0] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold34 (.A(_022_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold35 (.A(\regarray[7][3] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold36 (.A(\regarray[6][2] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold37 (.A(_012_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold38 (.A(\regarray[3][0] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold39 (.A(\regarray[3][3] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold40 (.A(\regarray[5][1] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold41 (.A(\regarray[5][2] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold42 (.A(_028_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold43 (.A(\regarray[3][2] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold44 (.A(uo_out[3]),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold45 (.A(_035_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold46 (.A(\regarray[5][3] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold47 (.A(_029_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold48 (.A(uo_out[2]),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold49 (.A(_034_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold50 (.A(\regarray[1][3] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold51 (.A(_025_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold52 (.A(\regarray[1][2] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold53 (.A(_024_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold54 (.A(uo_out[4]),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold55 (.A(_036_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold56 (.A(uo_out[5]),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold57 (.A(_037_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold58 (.A(_001_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold59 (.A(_080_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold60 (.A(_053_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold61 (.A(\rd_reg[2] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold62 (.A(_086_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold63 (.A(_051_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold64 (.A(\wr_next[0] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold65 (.A(_091_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold66 (.A(_046_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold67 (.A(\wr_reg[2] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold68 (.A(_048_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold69 (.A(dffr2),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold70 (.A(_084_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold71 (.A(\wr_next[0] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold72 (.A(\wr_next[0] ),
    .X(net149));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_4 FILLER_20_175 ();
 sg13g2_fill_2 FILLER_20_179 ();
 sg13g2_decap_8 FILLER_20_190 ();
 sg13g2_decap_8 FILLER_20_197 ();
 sg13g2_decap_8 FILLER_20_204 ();
 sg13g2_decap_8 FILLER_20_211 ();
 sg13g2_decap_8 FILLER_20_218 ();
 sg13g2_decap_8 FILLER_20_225 ();
 sg13g2_decap_8 FILLER_20_232 ();
 sg13g2_decap_8 FILLER_20_239 ();
 sg13g2_decap_8 FILLER_20_246 ();
 sg13g2_decap_8 FILLER_20_253 ();
 sg13g2_decap_8 FILLER_20_260 ();
 sg13g2_decap_8 FILLER_20_267 ();
 sg13g2_decap_8 FILLER_20_274 ();
 sg13g2_decap_8 FILLER_20_281 ();
 sg13g2_decap_8 FILLER_20_288 ();
 sg13g2_decap_8 FILLER_20_295 ();
 sg13g2_decap_8 FILLER_20_302 ();
 sg13g2_decap_8 FILLER_20_309 ();
 sg13g2_decap_8 FILLER_20_316 ();
 sg13g2_decap_8 FILLER_20_323 ();
 sg13g2_decap_8 FILLER_20_330 ();
 sg13g2_decap_8 FILLER_20_337 ();
 sg13g2_decap_8 FILLER_20_344 ();
 sg13g2_decap_8 FILLER_20_351 ();
 sg13g2_decap_8 FILLER_20_358 ();
 sg13g2_decap_8 FILLER_20_365 ();
 sg13g2_decap_8 FILLER_20_372 ();
 sg13g2_decap_8 FILLER_20_379 ();
 sg13g2_decap_8 FILLER_20_386 ();
 sg13g2_decap_8 FILLER_20_393 ();
 sg13g2_decap_8 FILLER_20_400 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_4 FILLER_21_112 ();
 sg13g2_fill_1 FILLER_21_126 ();
 sg13g2_fill_1 FILLER_21_136 ();
 sg13g2_fill_1 FILLER_21_160 ();
 sg13g2_decap_8 FILLER_21_191 ();
 sg13g2_fill_2 FILLER_21_198 ();
 sg13g2_fill_1 FILLER_21_200 ();
 sg13g2_decap_8 FILLER_21_205 ();
 sg13g2_fill_2 FILLER_21_212 ();
 sg13g2_fill_1 FILLER_21_214 ();
 sg13g2_fill_2 FILLER_21_250 ();
 sg13g2_decap_8 FILLER_21_256 ();
 sg13g2_decap_8 FILLER_21_263 ();
 sg13g2_decap_8 FILLER_21_270 ();
 sg13g2_decap_8 FILLER_21_277 ();
 sg13g2_decap_8 FILLER_21_284 ();
 sg13g2_decap_8 FILLER_21_291 ();
 sg13g2_decap_8 FILLER_21_298 ();
 sg13g2_decap_8 FILLER_21_305 ();
 sg13g2_decap_8 FILLER_21_312 ();
 sg13g2_decap_8 FILLER_21_319 ();
 sg13g2_decap_8 FILLER_21_326 ();
 sg13g2_decap_8 FILLER_21_333 ();
 sg13g2_decap_8 FILLER_21_340 ();
 sg13g2_decap_8 FILLER_21_347 ();
 sg13g2_decap_8 FILLER_21_354 ();
 sg13g2_decap_8 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_decap_8 FILLER_21_375 ();
 sg13g2_decap_8 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_21_389 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_fill_2 FILLER_22_105 ();
 sg13g2_fill_1 FILLER_22_107 ();
 sg13g2_decap_8 FILLER_22_134 ();
 sg13g2_fill_1 FILLER_22_230 ();
 sg13g2_decap_4 FILLER_22_276 ();
 sg13g2_fill_2 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_313 ();
 sg13g2_decap_8 FILLER_22_320 ();
 sg13g2_decap_8 FILLER_22_327 ();
 sg13g2_decap_8 FILLER_22_334 ();
 sg13g2_decap_8 FILLER_22_341 ();
 sg13g2_decap_8 FILLER_22_348 ();
 sg13g2_decap_8 FILLER_22_355 ();
 sg13g2_decap_8 FILLER_22_362 ();
 sg13g2_decap_8 FILLER_22_369 ();
 sg13g2_decap_8 FILLER_22_376 ();
 sg13g2_decap_8 FILLER_22_383 ();
 sg13g2_decap_8 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_fill_1 FILLER_23_105 ();
 sg13g2_fill_2 FILLER_23_110 ();
 sg13g2_fill_1 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_127 ();
 sg13g2_fill_1 FILLER_23_134 ();
 sg13g2_fill_2 FILLER_23_155 ();
 sg13g2_fill_1 FILLER_23_179 ();
 sg13g2_fill_2 FILLER_23_206 ();
 sg13g2_fill_2 FILLER_23_218 ();
 sg13g2_fill_1 FILLER_23_220 ();
 sg13g2_fill_1 FILLER_23_257 ();
 sg13g2_decap_8 FILLER_23_339 ();
 sg13g2_decap_8 FILLER_23_346 ();
 sg13g2_decap_8 FILLER_23_353 ();
 sg13g2_decap_8 FILLER_23_360 ();
 sg13g2_decap_8 FILLER_23_367 ();
 sg13g2_decap_8 FILLER_23_374 ();
 sg13g2_decap_8 FILLER_23_381 ();
 sg13g2_decap_8 FILLER_23_388 ();
 sg13g2_decap_8 FILLER_23_395 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_4 FILLER_24_91 ();
 sg13g2_fill_2 FILLER_24_147 ();
 sg13g2_fill_1 FILLER_24_149 ();
 sg13g2_fill_2 FILLER_24_189 ();
 sg13g2_fill_2 FILLER_24_217 ();
 sg13g2_fill_1 FILLER_24_219 ();
 sg13g2_fill_2 FILLER_24_251 ();
 sg13g2_fill_2 FILLER_24_281 ();
 sg13g2_fill_1 FILLER_24_283 ();
 sg13g2_decap_4 FILLER_24_294 ();
 sg13g2_fill_1 FILLER_24_306 ();
 sg13g2_decap_8 FILLER_24_339 ();
 sg13g2_decap_8 FILLER_24_346 ();
 sg13g2_decap_8 FILLER_24_353 ();
 sg13g2_decap_8 FILLER_24_360 ();
 sg13g2_decap_8 FILLER_24_367 ();
 sg13g2_decap_8 FILLER_24_374 ();
 sg13g2_decap_8 FILLER_24_381 ();
 sg13g2_decap_8 FILLER_24_388 ();
 sg13g2_decap_8 FILLER_24_395 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_fill_2 FILLER_25_112 ();
 sg13g2_fill_1 FILLER_25_114 ();
 sg13g2_fill_2 FILLER_25_128 ();
 sg13g2_fill_1 FILLER_25_130 ();
 sg13g2_fill_2 FILLER_25_155 ();
 sg13g2_fill_1 FILLER_25_157 ();
 sg13g2_decap_4 FILLER_25_206 ();
 sg13g2_fill_1 FILLER_25_210 ();
 sg13g2_fill_2 FILLER_25_246 ();
 sg13g2_fill_2 FILLER_25_289 ();
 sg13g2_fill_2 FILLER_25_317 ();
 sg13g2_decap_8 FILLER_25_345 ();
 sg13g2_decap_8 FILLER_25_352 ();
 sg13g2_decap_8 FILLER_25_359 ();
 sg13g2_decap_8 FILLER_25_366 ();
 sg13g2_decap_8 FILLER_25_373 ();
 sg13g2_decap_8 FILLER_25_380 ();
 sg13g2_decap_8 FILLER_25_387 ();
 sg13g2_decap_8 FILLER_25_394 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_fill_1 FILLER_26_98 ();
 sg13g2_decap_4 FILLER_26_152 ();
 sg13g2_fill_1 FILLER_26_166 ();
 sg13g2_fill_1 FILLER_26_217 ();
 sg13g2_fill_2 FILLER_26_239 ();
 sg13g2_fill_2 FILLER_26_251 ();
 sg13g2_decap_8 FILLER_26_295 ();
 sg13g2_fill_2 FILLER_26_325 ();
 sg13g2_fill_1 FILLER_26_327 ();
 sg13g2_decap_8 FILLER_26_345 ();
 sg13g2_decap_8 FILLER_26_352 ();
 sg13g2_decap_8 FILLER_26_359 ();
 sg13g2_decap_8 FILLER_26_366 ();
 sg13g2_decap_8 FILLER_26_373 ();
 sg13g2_decap_8 FILLER_26_380 ();
 sg13g2_decap_8 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_4 FILLER_27_91 ();
 sg13g2_fill_1 FILLER_27_131 ();
 sg13g2_fill_2 FILLER_27_150 ();
 sg13g2_fill_1 FILLER_27_152 ();
 sg13g2_fill_1 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_208 ();
 sg13g2_fill_2 FILLER_27_215 ();
 sg13g2_decap_8 FILLER_27_220 ();
 sg13g2_fill_2 FILLER_27_251 ();
 sg13g2_fill_1 FILLER_27_265 ();
 sg13g2_fill_1 FILLER_27_279 ();
 sg13g2_decap_8 FILLER_27_290 ();
 sg13g2_decap_4 FILLER_27_297 ();
 sg13g2_fill_1 FILLER_27_306 ();
 sg13g2_decap_8 FILLER_27_346 ();
 sg13g2_decap_8 FILLER_27_353 ();
 sg13g2_decap_8 FILLER_27_360 ();
 sg13g2_decap_8 FILLER_27_367 ();
 sg13g2_decap_8 FILLER_27_374 ();
 sg13g2_decap_8 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_27_388 ();
 sg13g2_decap_8 FILLER_27_395 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_fill_1 FILLER_28_132 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_fill_2 FILLER_28_161 ();
 sg13g2_fill_1 FILLER_28_163 ();
 sg13g2_fill_1 FILLER_28_168 ();
 sg13g2_fill_1 FILLER_28_183 ();
 sg13g2_decap_4 FILLER_28_197 ();
 sg13g2_fill_1 FILLER_28_201 ();
 sg13g2_decap_8 FILLER_28_206 ();
 sg13g2_fill_2 FILLER_28_218 ();
 sg13g2_fill_1 FILLER_28_220 ();
 sg13g2_fill_2 FILLER_28_226 ();
 sg13g2_fill_1 FILLER_28_258 ();
 sg13g2_fill_1 FILLER_28_267 ();
 sg13g2_decap_4 FILLER_28_283 ();
 sg13g2_decap_8 FILLER_28_347 ();
 sg13g2_decap_8 FILLER_28_354 ();
 sg13g2_decap_8 FILLER_28_361 ();
 sg13g2_decap_8 FILLER_28_368 ();
 sg13g2_decap_8 FILLER_28_375 ();
 sg13g2_decap_8 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_396 ();
 sg13g2_decap_4 FILLER_28_403 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_fill_1 FILLER_29_91 ();
 sg13g2_fill_2 FILLER_29_149 ();
 sg13g2_fill_2 FILLER_29_227 ();
 sg13g2_fill_1 FILLER_29_229 ();
 sg13g2_fill_2 FILLER_29_235 ();
 sg13g2_fill_1 FILLER_29_277 ();
 sg13g2_fill_1 FILLER_29_298 ();
 sg13g2_fill_2 FILLER_29_326 ();
 sg13g2_decap_8 FILLER_29_350 ();
 sg13g2_decap_8 FILLER_29_357 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_4 FILLER_30_98 ();
 sg13g2_fill_1 FILLER_30_115 ();
 sg13g2_fill_1 FILLER_30_135 ();
 sg13g2_fill_2 FILLER_30_160 ();
 sg13g2_fill_1 FILLER_30_176 ();
 sg13g2_fill_2 FILLER_30_191 ();
 sg13g2_fill_2 FILLER_30_232 ();
 sg13g2_fill_1 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_294 ();
 sg13g2_decap_8 FILLER_30_340 ();
 sg13g2_decap_8 FILLER_30_347 ();
 sg13g2_decap_8 FILLER_30_354 ();
 sg13g2_decap_8 FILLER_30_361 ();
 sg13g2_decap_8 FILLER_30_368 ();
 sg13g2_decap_8 FILLER_30_375 ();
 sg13g2_decap_8 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_30_389 ();
 sg13g2_decap_8 FILLER_30_396 ();
 sg13g2_decap_4 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_4 FILLER_31_91 ();
 sg13g2_fill_2 FILLER_31_95 ();
 sg13g2_decap_4 FILLER_31_138 ();
 sg13g2_fill_2 FILLER_31_184 ();
 sg13g2_fill_2 FILLER_31_235 ();
 sg13g2_fill_1 FILLER_31_280 ();
 sg13g2_fill_1 FILLER_31_309 ();
 sg13g2_decap_8 FILLER_31_336 ();
 sg13g2_decap_8 FILLER_31_343 ();
 sg13g2_decap_8 FILLER_31_350 ();
 sg13g2_decap_8 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_371 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_fill_2 FILLER_32_105 ();
 sg13g2_fill_1 FILLER_32_107 ();
 sg13g2_fill_1 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_188 ();
 sg13g2_fill_1 FILLER_32_199 ();
 sg13g2_fill_1 FILLER_32_213 ();
 sg13g2_fill_1 FILLER_32_274 ();
 sg13g2_fill_1 FILLER_32_280 ();
 sg13g2_fill_2 FILLER_32_298 ();
 sg13g2_fill_1 FILLER_32_300 ();
 sg13g2_decap_8 FILLER_32_327 ();
 sg13g2_decap_8 FILLER_32_334 ();
 sg13g2_decap_8 FILLER_32_341 ();
 sg13g2_decap_8 FILLER_32_348 ();
 sg13g2_decap_8 FILLER_32_355 ();
 sg13g2_decap_8 FILLER_32_362 ();
 sg13g2_decap_8 FILLER_32_369 ();
 sg13g2_decap_8 FILLER_32_376 ();
 sg13g2_decap_8 FILLER_32_383 ();
 sg13g2_decap_8 FILLER_32_390 ();
 sg13g2_decap_8 FILLER_32_397 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_4 FILLER_33_105 ();
 sg13g2_fill_1 FILLER_33_109 ();
 sg13g2_fill_2 FILLER_33_145 ();
 sg13g2_fill_2 FILLER_33_165 ();
 sg13g2_fill_2 FILLER_33_180 ();
 sg13g2_fill_1 FILLER_33_182 ();
 sg13g2_fill_2 FILLER_33_197 ();
 sg13g2_fill_2 FILLER_33_264 ();
 sg13g2_fill_1 FILLER_33_318 ();
 sg13g2_decap_8 FILLER_33_328 ();
 sg13g2_decap_8 FILLER_33_335 ();
 sg13g2_decap_8 FILLER_33_342 ();
 sg13g2_decap_8 FILLER_33_349 ();
 sg13g2_decap_8 FILLER_33_356 ();
 sg13g2_decap_8 FILLER_33_363 ();
 sg13g2_decap_8 FILLER_33_370 ();
 sg13g2_decap_8 FILLER_33_377 ();
 sg13g2_decap_8 FILLER_33_384 ();
 sg13g2_decap_8 FILLER_33_391 ();
 sg13g2_decap_8 FILLER_33_398 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_4 FILLER_34_128 ();
 sg13g2_fill_1 FILLER_34_132 ();
 sg13g2_decap_4 FILLER_34_138 ();
 sg13g2_decap_4 FILLER_34_172 ();
 sg13g2_fill_2 FILLER_34_220 ();
 sg13g2_fill_2 FILLER_34_253 ();
 sg13g2_fill_2 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_321 ();
 sg13g2_decap_8 FILLER_34_328 ();
 sg13g2_decap_8 FILLER_34_335 ();
 sg13g2_decap_8 FILLER_34_342 ();
 sg13g2_decap_8 FILLER_34_349 ();
 sg13g2_decap_8 FILLER_34_356 ();
 sg13g2_decap_8 FILLER_34_363 ();
 sg13g2_decap_8 FILLER_34_370 ();
 sg13g2_decap_8 FILLER_34_377 ();
 sg13g2_decap_8 FILLER_34_384 ();
 sg13g2_decap_8 FILLER_34_391 ();
 sg13g2_decap_8 FILLER_34_398 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_fill_2 FILLER_35_133 ();
 sg13g2_fill_1 FILLER_35_135 ();
 sg13g2_decap_8 FILLER_35_141 ();
 sg13g2_decap_4 FILLER_35_148 ();
 sg13g2_decap_4 FILLER_35_160 ();
 sg13g2_fill_1 FILLER_35_164 ();
 sg13g2_decap_8 FILLER_35_174 ();
 sg13g2_decap_4 FILLER_35_181 ();
 sg13g2_fill_2 FILLER_35_185 ();
 sg13g2_decap_8 FILLER_35_191 ();
 sg13g2_decap_8 FILLER_35_198 ();
 sg13g2_decap_4 FILLER_35_205 ();
 sg13g2_fill_1 FILLER_35_209 ();
 sg13g2_decap_4 FILLER_35_214 ();
 sg13g2_decap_8 FILLER_35_222 ();
 sg13g2_decap_4 FILLER_35_229 ();
 sg13g2_fill_2 FILLER_35_233 ();
 sg13g2_fill_2 FILLER_35_266 ();
 sg13g2_fill_1 FILLER_35_268 ();
 sg13g2_decap_8 FILLER_35_302 ();
 sg13g2_decap_8 FILLER_35_309 ();
 sg13g2_decap_8 FILLER_35_316 ();
 sg13g2_decap_8 FILLER_35_323 ();
 sg13g2_decap_8 FILLER_35_330 ();
 sg13g2_decap_8 FILLER_35_337 ();
 sg13g2_decap_8 FILLER_35_344 ();
 sg13g2_decap_8 FILLER_35_351 ();
 sg13g2_decap_8 FILLER_35_358 ();
 sg13g2_decap_8 FILLER_35_365 ();
 sg13g2_decap_8 FILLER_35_372 ();
 sg13g2_decap_8 FILLER_35_379 ();
 sg13g2_decap_8 FILLER_35_386 ();
 sg13g2_decap_8 FILLER_35_393 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_fill_2 FILLER_36_264 ();
 sg13g2_fill_1 FILLER_36_266 ();
 sg13g2_decap_8 FILLER_36_292 ();
 sg13g2_decap_8 FILLER_36_299 ();
 sg13g2_decap_8 FILLER_36_306 ();
 sg13g2_decap_8 FILLER_36_313 ();
 sg13g2_decap_8 FILLER_36_320 ();
 sg13g2_decap_8 FILLER_36_327 ();
 sg13g2_decap_8 FILLER_36_334 ();
 sg13g2_decap_8 FILLER_36_341 ();
 sg13g2_decap_8 FILLER_36_348 ();
 sg13g2_decap_8 FILLER_36_355 ();
 sg13g2_decap_8 FILLER_36_362 ();
 sg13g2_decap_8 FILLER_36_369 ();
 sg13g2_decap_8 FILLER_36_376 ();
 sg13g2_decap_8 FILLER_36_383 ();
 sg13g2_decap_8 FILLER_36_390 ();
 sg13g2_decap_8 FILLER_36_397 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_4 FILLER_37_231 ();
 sg13g2_fill_1 FILLER_37_235 ();
 sg13g2_decap_8 FILLER_37_297 ();
 sg13g2_decap_8 FILLER_37_304 ();
 sg13g2_decap_8 FILLER_37_311 ();
 sg13g2_decap_8 FILLER_37_318 ();
 sg13g2_decap_8 FILLER_37_325 ();
 sg13g2_decap_8 FILLER_37_332 ();
 sg13g2_decap_8 FILLER_37_339 ();
 sg13g2_decap_8 FILLER_37_346 ();
 sg13g2_decap_8 FILLER_37_353 ();
 sg13g2_decap_8 FILLER_37_360 ();
 sg13g2_decap_8 FILLER_37_367 ();
 sg13g2_decap_8 FILLER_37_374 ();
 sg13g2_decap_8 FILLER_37_381 ();
 sg13g2_decap_8 FILLER_37_388 ();
 sg13g2_decap_8 FILLER_37_395 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_4 FILLER_38_180 ();
 sg13g2_decap_4 FILLER_38_188 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_decap_8 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_fill_2 FILLER_38_245 ();
 sg13g2_decap_4 FILLER_38_256 ();
 sg13g2_fill_2 FILLER_38_260 ();
 sg13g2_decap_8 FILLER_38_282 ();
 sg13g2_decap_8 FILLER_38_289 ();
 sg13g2_decap_8 FILLER_38_296 ();
 sg13g2_decap_8 FILLER_38_303 ();
 sg13g2_fill_2 FILLER_38_310 ();
 sg13g2_decap_4 FILLER_38_348 ();
 sg13g2_decap_8 FILLER_38_356 ();
 sg13g2_decap_8 FILLER_38_363 ();
 sg13g2_decap_4 FILLER_38_370 ();
 sg13g2_fill_2 FILLER_38_374 ();
 sg13g2_decap_8 FILLER_38_384 ();
 sg13g2_decap_8 FILLER_38_391 ();
 sg13g2_decap_8 FILLER_38_398 ();
 sg13g2_decap_4 FILLER_38_405 ();
 assign uio_oe[0] = net8;
 assign uio_oe[1] = net9;
 assign uio_oe[2] = net10;
 assign uio_oe[3] = net11;
 assign uio_oe[4] = net12;
 assign uio_oe[5] = net13;
 assign uio_oe[6] = net14;
 assign uio_oe[7] = net15;
 assign uio_out[0] = net16;
 assign uio_out[1] = net17;
 assign uio_out[2] = net18;
 assign uio_out[3] = net19;
 assign uio_out[4] = net20;
 assign uio_out[5] = net21;
 assign uio_out[6] = net22;
 assign uio_out[7] = net23;
 assign uo_out[6] = net24;
 assign uo_out[7] = net25;
endmodule

module tt_um_underserved (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire clknet_leaf_0_clk;
 wire \cpu.alu.add_cy_r ;
 wire \cpu.alu.cmp_r ;
 wire \cpu.bne_or_bge ;
 wire \cpu.branch_op ;
 wire \cpu.bufreg.c_r ;
 wire \cpu.bufreg.data[0] ;
 wire \cpu.bufreg.data[10] ;
 wire \cpu.bufreg.data[11] ;
 wire \cpu.bufreg.data[12] ;
 wire \cpu.bufreg.data[13] ;
 wire \cpu.bufreg.data[14] ;
 wire \cpu.bufreg.data[15] ;
 wire \cpu.bufreg.data[16] ;
 wire \cpu.bufreg.data[17] ;
 wire \cpu.bufreg.data[18] ;
 wire \cpu.bufreg.data[19] ;
 wire \cpu.bufreg.data[1] ;
 wire \cpu.bufreg.data[20] ;
 wire \cpu.bufreg.data[21] ;
 wire \cpu.bufreg.data[22] ;
 wire \cpu.bufreg.data[23] ;
 wire \cpu.bufreg.data[24] ;
 wire \cpu.bufreg.data[25] ;
 wire \cpu.bufreg.data[26] ;
 wire \cpu.bufreg.data[27] ;
 wire \cpu.bufreg.data[28] ;
 wire \cpu.bufreg.data[29] ;
 wire \cpu.bufreg.data[2] ;
 wire \cpu.bufreg.data[30] ;
 wire \cpu.bufreg.data[31] ;
 wire \cpu.bufreg.data[3] ;
 wire \cpu.bufreg.data[4] ;
 wire \cpu.bufreg.data[5] ;
 wire \cpu.bufreg.data[6] ;
 wire \cpu.bufreg.data[7] ;
 wire \cpu.bufreg.data[8] ;
 wire \cpu.bufreg.data[9] ;
 wire \cpu.bufreg.i_sh_signed ;
 wire \cpu.bufreg2.dat[0] ;
 wire \cpu.bufreg2.dat[10] ;
 wire \cpu.bufreg2.dat[11] ;
 wire \cpu.bufreg2.dat[12] ;
 wire \cpu.bufreg2.dat[13] ;
 wire \cpu.bufreg2.dat[14] ;
 wire \cpu.bufreg2.dat[15] ;
 wire \cpu.bufreg2.dat[16] ;
 wire \cpu.bufreg2.dat[17] ;
 wire \cpu.bufreg2.dat[18] ;
 wire \cpu.bufreg2.dat[19] ;
 wire \cpu.bufreg2.dat[1] ;
 wire \cpu.bufreg2.dat[20] ;
 wire \cpu.bufreg2.dat[21] ;
 wire \cpu.bufreg2.dat[22] ;
 wire \cpu.bufreg2.dat[23] ;
 wire \cpu.bufreg2.dat[24] ;
 wire \cpu.bufreg2.dat[25] ;
 wire \cpu.bufreg2.dat[26] ;
 wire \cpu.bufreg2.dat[27] ;
 wire \cpu.bufreg2.dat[28] ;
 wire \cpu.bufreg2.dat[29] ;
 wire \cpu.bufreg2.dat[2] ;
 wire \cpu.bufreg2.dat[30] ;
 wire \cpu.bufreg2.dat[31] ;
 wire \cpu.bufreg2.dat[3] ;
 wire \cpu.bufreg2.dat[4] ;
 wire \cpu.bufreg2.dat[5] ;
 wire \cpu.bufreg2.dat[6] ;
 wire \cpu.bufreg2.dat[7] ;
 wire \cpu.bufreg2.dat[8] ;
 wire \cpu.bufreg2.dat[9] ;
 wire \cpu.bufreg2.i_dat[0] ;
 wire \cpu.bufreg2.i_dat[10] ;
 wire \cpu.bufreg2.i_dat[11] ;
 wire \cpu.bufreg2.i_dat[12] ;
 wire \cpu.bufreg2.i_dat[13] ;
 wire \cpu.bufreg2.i_dat[14] ;
 wire \cpu.bufreg2.i_dat[15] ;
 wire \cpu.bufreg2.i_dat[16] ;
 wire \cpu.bufreg2.i_dat[17] ;
 wire \cpu.bufreg2.i_dat[18] ;
 wire \cpu.bufreg2.i_dat[19] ;
 wire \cpu.bufreg2.i_dat[1] ;
 wire \cpu.bufreg2.i_dat[20] ;
 wire \cpu.bufreg2.i_dat[21] ;
 wire \cpu.bufreg2.i_dat[22] ;
 wire \cpu.bufreg2.i_dat[23] ;
 wire \cpu.bufreg2.i_dat[24] ;
 wire \cpu.bufreg2.i_dat[25] ;
 wire \cpu.bufreg2.i_dat[26] ;
 wire \cpu.bufreg2.i_dat[27] ;
 wire \cpu.bufreg2.i_dat[28] ;
 wire \cpu.bufreg2.i_dat[29] ;
 wire \cpu.bufreg2.i_dat[2] ;
 wire \cpu.bufreg2.i_dat[30] ;
 wire \cpu.bufreg2.i_dat[31] ;
 wire \cpu.bufreg2.i_dat[3] ;
 wire \cpu.bufreg2.i_dat[4] ;
 wire \cpu.bufreg2.i_dat[5] ;
 wire \cpu.bufreg2.i_dat[6] ;
 wire \cpu.bufreg2.i_dat[7] ;
 wire \cpu.bufreg2.i_dat[8] ;
 wire \cpu.bufreg2.i_dat[9] ;
 wire \cpu.bufreg2.i_op_b_sel ;
 wire \cpu.csr_d_sel ;
 wire \cpu.csr_imm ;
 wire \cpu.ctrl.i_jump ;
 wire \cpu.ctrl.o_ibus_adr[0] ;
 wire \cpu.ctrl.o_ibus_adr[10] ;
 wire \cpu.ctrl.o_ibus_adr[11] ;
 wire \cpu.ctrl.o_ibus_adr[12] ;
 wire \cpu.ctrl.o_ibus_adr[13] ;
 wire \cpu.ctrl.o_ibus_adr[14] ;
 wire \cpu.ctrl.o_ibus_adr[15] ;
 wire \cpu.ctrl.o_ibus_adr[16] ;
 wire \cpu.ctrl.o_ibus_adr[17] ;
 wire \cpu.ctrl.o_ibus_adr[18] ;
 wire \cpu.ctrl.o_ibus_adr[19] ;
 wire \cpu.ctrl.o_ibus_adr[1] ;
 wire \cpu.ctrl.o_ibus_adr[20] ;
 wire \cpu.ctrl.o_ibus_adr[21] ;
 wire \cpu.ctrl.o_ibus_adr[22] ;
 wire \cpu.ctrl.o_ibus_adr[23] ;
 wire \cpu.ctrl.o_ibus_adr[24] ;
 wire \cpu.ctrl.o_ibus_adr[25] ;
 wire \cpu.ctrl.o_ibus_adr[26] ;
 wire \cpu.ctrl.o_ibus_adr[27] ;
 wire \cpu.ctrl.o_ibus_adr[28] ;
 wire \cpu.ctrl.o_ibus_adr[29] ;
 wire \cpu.ctrl.o_ibus_adr[2] ;
 wire \cpu.ctrl.o_ibus_adr[30] ;
 wire \cpu.ctrl.o_ibus_adr[31] ;
 wire \cpu.ctrl.o_ibus_adr[3] ;
 wire \cpu.ctrl.o_ibus_adr[4] ;
 wire \cpu.ctrl.o_ibus_adr[5] ;
 wire \cpu.ctrl.o_ibus_adr[6] ;
 wire \cpu.ctrl.o_ibus_adr[7] ;
 wire \cpu.ctrl.o_ibus_adr[8] ;
 wire \cpu.ctrl.o_ibus_adr[9] ;
 wire \cpu.ctrl.pc_plus_4_cy_r ;
 wire \cpu.ctrl.pc_plus_offset_cy_r ;
 wire \cpu.decode.co_ebreak ;
 wire \cpu.decode.co_mem_word ;
 wire \cpu.decode.opcode[0] ;
 wire \cpu.decode.opcode[1] ;
 wire \cpu.decode.opcode[2] ;
 wire \cpu.immdec.imm11_7[0] ;
 wire \cpu.immdec.imm11_7[1] ;
 wire \cpu.immdec.imm11_7[2] ;
 wire \cpu.immdec.imm11_7[3] ;
 wire \cpu.immdec.imm11_7[4] ;
 wire \cpu.immdec.imm19_12_20[0] ;
 wire \cpu.immdec.imm19_12_20[1] ;
 wire \cpu.immdec.imm19_12_20[2] ;
 wire \cpu.immdec.imm19_12_20[3] ;
 wire \cpu.immdec.imm19_12_20[5] ;
 wire \cpu.immdec.imm19_12_20[6] ;
 wire \cpu.immdec.imm19_12_20[7] ;
 wire \cpu.immdec.imm19_12_20[8] ;
 wire \cpu.immdec.imm24_20[0] ;
 wire \cpu.immdec.imm24_20[1] ;
 wire \cpu.immdec.imm24_20[2] ;
 wire \cpu.immdec.imm24_20[3] ;
 wire \cpu.immdec.imm24_20[4] ;
 wire \cpu.immdec.imm30_25[0] ;
 wire \cpu.immdec.imm30_25[1] ;
 wire \cpu.immdec.imm30_25[2] ;
 wire \cpu.immdec.imm30_25[3] ;
 wire \cpu.immdec.imm30_25[4] ;
 wire \cpu.immdec.imm30_25[5] ;
 wire \cpu.immdec.imm31 ;
 wire \cpu.immdec.imm7 ;
 wire \cpu.mem_bytecnt[0] ;
 wire \cpu.mem_bytecnt[1] ;
 wire \cpu.mem_if.signbit ;
 wire \cpu.state.cnt_r[0] ;
 wire \cpu.state.cnt_r[1] ;
 wire \cpu.state.cnt_r[2] ;
 wire \cpu.state.cnt_r[3] ;
 wire \cpu.state.ibus_cyc ;
 wire \cpu.state.init_done ;
 wire \cpu.state.o_cnt[2] ;
 wire \cpu.state.stage_two_req ;
 wire \dut.buffer[0] ;
 wire \dut.buffer[10] ;
 wire \dut.buffer[11] ;
 wire \dut.buffer[12] ;
 wire \dut.buffer[13] ;
 wire \dut.buffer[14] ;
 wire \dut.buffer[15] ;
 wire \dut.buffer[16] ;
 wire \dut.buffer[17] ;
 wire \dut.buffer[18] ;
 wire \dut.buffer[19] ;
 wire \dut.buffer[1] ;
 wire \dut.buffer[20] ;
 wire \dut.buffer[21] ;
 wire \dut.buffer[22] ;
 wire \dut.buffer[23] ;
 wire \dut.buffer[2] ;
 wire \dut.buffer[3] ;
 wire \dut.buffer[4] ;
 wire \dut.buffer[5] ;
 wire \dut.buffer[6] ;
 wire \dut.buffer[7] ;
 wire \dut.buffer[8] ;
 wire \dut.buffer[9] ;
 wire \dut.din_data[0] ;
 wire \dut.din_data[1] ;
 wire \dut.din_data[2] ;
 wire \dut.din_data[3] ;
 wire \dut.din_data[4] ;
 wire \dut.din_data[5] ;
 wire \dut.din_data[6] ;
 wire \dut.din_data[7] ;
 wire \dut.din_rd ;
 wire \dut.din_tag[0] ;
 wire \dut.din_tag[1] ;
 wire \dut.din_tag[2] ;
 wire \dut.din_valid ;
 wire \dut.dout_data[0] ;
 wire \dut.dout_data[1] ;
 wire \dut.dout_data[2] ;
 wire \dut.dout_data[3] ;
 wire \dut.dout_data[4] ;
 wire \dut.dout_data[5] ;
 wire \dut.dout_data[6] ;
 wire \dut.dout_data[7] ;
 wire \dut.dout_tag[0] ;
 wire \dut.dout_tag[1] ;
 wire \dut.dout_tag[2] ;
 wire \dut.flash_clk ;
 wire \dut.flash_csb ;
 wire \dut.flash_io0_do ;
 wire \dut.rd_addr[0] ;
 wire \dut.rd_addr[10] ;
 wire \dut.rd_addr[11] ;
 wire \dut.rd_addr[12] ;
 wire \dut.rd_addr[13] ;
 wire \dut.rd_addr[14] ;
 wire \dut.rd_addr[15] ;
 wire \dut.rd_addr[16] ;
 wire \dut.rd_addr[17] ;
 wire \dut.rd_addr[18] ;
 wire \dut.rd_addr[19] ;
 wire \dut.rd_addr[1] ;
 wire \dut.rd_addr[20] ;
 wire \dut.rd_addr[21] ;
 wire \dut.rd_addr[22] ;
 wire \dut.rd_addr[23] ;
 wire \dut.rd_addr[2] ;
 wire \dut.rd_addr[3] ;
 wire \dut.rd_addr[4] ;
 wire \dut.rd_addr[5] ;
 wire \dut.rd_addr[6] ;
 wire \dut.rd_addr[7] ;
 wire \dut.rd_addr[8] ;
 wire \dut.rd_addr[9] ;
 wire \dut.rd_inc ;
 wire \dut.rd_valid ;
 wire \dut.rd_wait ;
 wire \dut.softreset ;
 wire \dut.state[0] ;
 wire \dut.state[10] ;
 wire \dut.state[11] ;
 wire \dut.state[12] ;
 wire \dut.state[1] ;
 wire \dut.state[2] ;
 wire \dut.state[3] ;
 wire \dut.state[4] ;
 wire \dut.state[5] ;
 wire \dut.state[6] ;
 wire \dut.state[7] ;
 wire \dut.state[8] ;
 wire \dut.state[9] ;
 wire \dut.xfer.count[0] ;
 wire \dut.xfer.count[1] ;
 wire \dut.xfer.count[2] ;
 wire \dut.xfer.count[3] ;
 wire \dut.xfer.dummy_count[0] ;
 wire \dut.xfer.dummy_count[1] ;
 wire \dut.xfer.dummy_count[2] ;
 wire \dut.xfer.dummy_count[3] ;
 wire \dut.xfer.fetch ;
 wire \dut.xfer.next_obuffer[1] ;
 wire \dut.xfer.next_obuffer[2] ;
 wire \dut.xfer.next_obuffer[3] ;
 wire \dut.xfer.next_obuffer[4] ;
 wire \dut.xfer.next_obuffer[5] ;
 wire \dut.xfer.next_obuffer[6] ;
 wire \dut.xfer.next_obuffer[7] ;
 wire \dut.xfer.obuffer[7] ;
 wire \dut.xfer.resetn ;
 wire \dut.xfer.xfer_tag[0] ;
 wire \dut.xfer.xfer_tag[1] ;
 wire \dut.xfer.xfer_tag[2] ;
 wire \gpio.o_wb_ack ;
 wire \rf_shift_reg.cnt[0] ;
 wire \rf_shift_reg.cnt[1] ;
 wire \rf_shift_reg.cnt[2] ;
 wire \rf_shift_reg.cnt[3] ;
 wire \rf_shift_reg.cnt[4] ;
 wire \rf_shift_reg.rd_active ;
 wire \rf_shift_reg.rdata[1] ;
 wire \rf_shift_reg.rdata[2] ;
 wire \rf_shift_reg.rdata[3] ;
 wire \rf_shift_reg.rdata[4] ;
 wire \rf_shift_reg.rdata[5] ;
 wire \rf_shift_reg.rreq_2r ;
 wire \rf_shift_reg.rreq_r ;
 wire \rf_shift_reg.x[1][10] ;
 wire \rf_shift_reg.x[1][11] ;
 wire \rf_shift_reg.x[1][12] ;
 wire \rf_shift_reg.x[1][13] ;
 wire \rf_shift_reg.x[1][14] ;
 wire \rf_shift_reg.x[1][15] ;
 wire \rf_shift_reg.x[1][16] ;
 wire \rf_shift_reg.x[1][17] ;
 wire \rf_shift_reg.x[1][18] ;
 wire \rf_shift_reg.x[1][19] ;
 wire \rf_shift_reg.x[1][1] ;
 wire \rf_shift_reg.x[1][20] ;
 wire \rf_shift_reg.x[1][21] ;
 wire \rf_shift_reg.x[1][22] ;
 wire \rf_shift_reg.x[1][23] ;
 wire \rf_shift_reg.x[1][24] ;
 wire \rf_shift_reg.x[1][25] ;
 wire \rf_shift_reg.x[1][26] ;
 wire \rf_shift_reg.x[1][27] ;
 wire \rf_shift_reg.x[1][28] ;
 wire \rf_shift_reg.x[1][29] ;
 wire \rf_shift_reg.x[1][2] ;
 wire \rf_shift_reg.x[1][30] ;
 wire \rf_shift_reg.x[1][31] ;
 wire \rf_shift_reg.x[1][3] ;
 wire \rf_shift_reg.x[1][4] ;
 wire \rf_shift_reg.x[1][5] ;
 wire \rf_shift_reg.x[1][6] ;
 wire \rf_shift_reg.x[1][7] ;
 wire \rf_shift_reg.x[1][8] ;
 wire \rf_shift_reg.x[1][9] ;
 wire \rf_shift_reg.x[2][10] ;
 wire \rf_shift_reg.x[2][11] ;
 wire \rf_shift_reg.x[2][12] ;
 wire \rf_shift_reg.x[2][13] ;
 wire \rf_shift_reg.x[2][14] ;
 wire \rf_shift_reg.x[2][15] ;
 wire \rf_shift_reg.x[2][16] ;
 wire \rf_shift_reg.x[2][17] ;
 wire \rf_shift_reg.x[2][18] ;
 wire \rf_shift_reg.x[2][19] ;
 wire \rf_shift_reg.x[2][1] ;
 wire \rf_shift_reg.x[2][20] ;
 wire \rf_shift_reg.x[2][21] ;
 wire \rf_shift_reg.x[2][22] ;
 wire \rf_shift_reg.x[2][23] ;
 wire \rf_shift_reg.x[2][24] ;
 wire \rf_shift_reg.x[2][25] ;
 wire \rf_shift_reg.x[2][26] ;
 wire \rf_shift_reg.x[2][27] ;
 wire \rf_shift_reg.x[2][28] ;
 wire \rf_shift_reg.x[2][29] ;
 wire \rf_shift_reg.x[2][2] ;
 wire \rf_shift_reg.x[2][30] ;
 wire \rf_shift_reg.x[2][31] ;
 wire \rf_shift_reg.x[2][3] ;
 wire \rf_shift_reg.x[2][4] ;
 wire \rf_shift_reg.x[2][5] ;
 wire \rf_shift_reg.x[2][6] ;
 wire \rf_shift_reg.x[2][7] ;
 wire \rf_shift_reg.x[2][8] ;
 wire \rf_shift_reg.x[2][9] ;
 wire \rf_shift_reg.x[3][10] ;
 wire \rf_shift_reg.x[3][11] ;
 wire \rf_shift_reg.x[3][12] ;
 wire \rf_shift_reg.x[3][13] ;
 wire \rf_shift_reg.x[3][14] ;
 wire \rf_shift_reg.x[3][15] ;
 wire \rf_shift_reg.x[3][16] ;
 wire \rf_shift_reg.x[3][17] ;
 wire \rf_shift_reg.x[3][18] ;
 wire \rf_shift_reg.x[3][19] ;
 wire \rf_shift_reg.x[3][1] ;
 wire \rf_shift_reg.x[3][20] ;
 wire \rf_shift_reg.x[3][21] ;
 wire \rf_shift_reg.x[3][22] ;
 wire \rf_shift_reg.x[3][23] ;
 wire \rf_shift_reg.x[3][24] ;
 wire \rf_shift_reg.x[3][25] ;
 wire \rf_shift_reg.x[3][26] ;
 wire \rf_shift_reg.x[3][27] ;
 wire \rf_shift_reg.x[3][28] ;
 wire \rf_shift_reg.x[3][29] ;
 wire \rf_shift_reg.x[3][2] ;
 wire \rf_shift_reg.x[3][30] ;
 wire \rf_shift_reg.x[3][31] ;
 wire \rf_shift_reg.x[3][3] ;
 wire \rf_shift_reg.x[3][4] ;
 wire \rf_shift_reg.x[3][5] ;
 wire \rf_shift_reg.x[3][6] ;
 wire \rf_shift_reg.x[3][7] ;
 wire \rf_shift_reg.x[3][8] ;
 wire \rf_shift_reg.x[3][9] ;
 wire \rf_shift_reg.x[4][10] ;
 wire \rf_shift_reg.x[4][11] ;
 wire \rf_shift_reg.x[4][12] ;
 wire \rf_shift_reg.x[4][13] ;
 wire \rf_shift_reg.x[4][14] ;
 wire \rf_shift_reg.x[4][15] ;
 wire \rf_shift_reg.x[4][16] ;
 wire \rf_shift_reg.x[4][17] ;
 wire \rf_shift_reg.x[4][18] ;
 wire \rf_shift_reg.x[4][19] ;
 wire \rf_shift_reg.x[4][1] ;
 wire \rf_shift_reg.x[4][20] ;
 wire \rf_shift_reg.x[4][21] ;
 wire \rf_shift_reg.x[4][22] ;
 wire \rf_shift_reg.x[4][23] ;
 wire \rf_shift_reg.x[4][24] ;
 wire \rf_shift_reg.x[4][25] ;
 wire \rf_shift_reg.x[4][26] ;
 wire \rf_shift_reg.x[4][27] ;
 wire \rf_shift_reg.x[4][28] ;
 wire \rf_shift_reg.x[4][29] ;
 wire \rf_shift_reg.x[4][2] ;
 wire \rf_shift_reg.x[4][30] ;
 wire \rf_shift_reg.x[4][31] ;
 wire \rf_shift_reg.x[4][3] ;
 wire \rf_shift_reg.x[4][4] ;
 wire \rf_shift_reg.x[4][5] ;
 wire \rf_shift_reg.x[4][6] ;
 wire \rf_shift_reg.x[4][7] ;
 wire \rf_shift_reg.x[4][8] ;
 wire \rf_shift_reg.x[4][9] ;
 wire \rf_shift_reg.x[5][10] ;
 wire \rf_shift_reg.x[5][11] ;
 wire \rf_shift_reg.x[5][12] ;
 wire \rf_shift_reg.x[5][13] ;
 wire \rf_shift_reg.x[5][14] ;
 wire \rf_shift_reg.x[5][15] ;
 wire \rf_shift_reg.x[5][16] ;
 wire \rf_shift_reg.x[5][17] ;
 wire \rf_shift_reg.x[5][18] ;
 wire \rf_shift_reg.x[5][19] ;
 wire \rf_shift_reg.x[5][1] ;
 wire \rf_shift_reg.x[5][20] ;
 wire \rf_shift_reg.x[5][21] ;
 wire \rf_shift_reg.x[5][22] ;
 wire \rf_shift_reg.x[5][23] ;
 wire \rf_shift_reg.x[5][24] ;
 wire \rf_shift_reg.x[5][25] ;
 wire \rf_shift_reg.x[5][26] ;
 wire \rf_shift_reg.x[5][27] ;
 wire \rf_shift_reg.x[5][28] ;
 wire \rf_shift_reg.x[5][29] ;
 wire \rf_shift_reg.x[5][2] ;
 wire \rf_shift_reg.x[5][30] ;
 wire \rf_shift_reg.x[5][31] ;
 wire \rf_shift_reg.x[5][3] ;
 wire \rf_shift_reg.x[5][4] ;
 wire \rf_shift_reg.x[5][5] ;
 wire \rf_shift_reg.x[5][6] ;
 wire \rf_shift_reg.x[5][7] ;
 wire \rf_shift_reg.x[5][8] ;
 wire \rf_shift_reg.x[5][9] ;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net1;
 wire net2;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;

 sg13g2_inv_1 _2317_ (.Y(_0542_),
    .A(net804));
 sg13g2_inv_1 _2318_ (.Y(_0543_),
    .A(net765));
 sg13g2_inv_1 _2319_ (.Y(_0544_),
    .A(net688));
 sg13g2_inv_1 _2320_ (.Y(_0545_),
    .A(net1220));
 sg13g2_inv_1 _2321_ (.Y(_0546_),
    .A(net1259));
 sg13g2_inv_1 _2322_ (.Y(_0547_),
    .A(\dut.xfer.count[3] ));
 sg13g2_inv_1 _2323_ (.Y(_0548_),
    .A(net567));
 sg13g2_inv_1 _2324_ (.Y(_0549_),
    .A(net1128));
 sg13g2_inv_1 _2325_ (.Y(_0550_),
    .A(net1203));
 sg13g2_inv_2 _2326_ (.Y(_0465_),
    .A(net585));
 sg13g2_inv_1 _2327_ (.Y(_0551_),
    .A(net1226));
 sg13g2_inv_1 _2328_ (.Y(_0552_),
    .A(net1244));
 sg13g2_inv_1 _2329_ (.Y(_0553_),
    .A(net1200));
 sg13g2_inv_1 _2330_ (.Y(_0554_),
    .A(net1213));
 sg13g2_inv_1 _2331_ (.Y(_0555_),
    .A(net1205));
 sg13g2_inv_1 _2332_ (.Y(_0556_),
    .A(net1138));
 sg13g2_inv_1 _2333_ (.Y(_0557_),
    .A(net636));
 sg13g2_inv_1 _2334_ (.Y(_0558_),
    .A(net794));
 sg13g2_inv_1 _2335_ (.Y(_0559_),
    .A(\dut.state[4] ));
 sg13g2_inv_1 _2336_ (.Y(_0560_),
    .A(\dut.state[6] ));
 sg13g2_inv_1 _2337_ (.Y(_0561_),
    .A(\dut.state[5] ));
 sg13g2_inv_1 _2338_ (.Y(_0562_),
    .A(\dut.state[9] ));
 sg13g2_inv_1 _2339_ (.Y(_0563_),
    .A(net571));
 sg13g2_inv_1 _2340_ (.Y(_0564_),
    .A(_0020_));
 sg13g2_inv_1 _2341_ (.Y(_0565_),
    .A(_0021_));
 sg13g2_inv_2 _2342_ (.Y(_0566_),
    .A(_0026_));
 sg13g2_inv_1 _2343_ (.Y(_0567_),
    .A(_0029_));
 sg13g2_inv_1 _2344_ (.Y(_0568_),
    .A(_0088_));
 sg13g2_inv_1 _2345_ (.Y(_0569_),
    .A(net720));
 sg13g2_inv_1 _2346_ (.Y(_0570_),
    .A(\dut.state[11] ));
 sg13g2_inv_1 _2347_ (.Y(_0571_),
    .A(net1098));
 sg13g2_inv_1 _2348_ (.Y(_0572_),
    .A(net854));
 sg13g2_inv_1 _2349_ (.Y(_0573_),
    .A(net1215));
 sg13g2_inv_1 _2350_ (.Y(_0574_),
    .A(net1327));
 sg13g2_inv_1 _2351_ (.Y(_0575_),
    .A(net1304));
 sg13g2_inv_1 _2352_ (.Y(_0576_),
    .A(_0090_));
 sg13g2_inv_1 _2353_ (.Y(_0577_),
    .A(_0089_));
 sg13g2_inv_1 _2354_ (.Y(_0578_),
    .A(_0091_));
 sg13g2_inv_1 _2355_ (.Y(_0579_),
    .A(net1276));
 sg13g2_inv_1 _2356_ (.Y(_0580_),
    .A(_0092_));
 sg13g2_inv_1 _2357_ (.Y(_0581_),
    .A(net1209));
 sg13g2_inv_2 _2358_ (.Y(_0582_),
    .A(\cpu.bufreg.data[0] ));
 sg13g2_inv_1 _2359_ (.Y(_0583_),
    .A(\cpu.immdec.imm24_20[0] ));
 sg13g2_inv_1 _2360_ (.Y(_0584_),
    .A(\rf_shift_reg.rdata[1] ));
 sg13g2_inv_1 _2361_ (.Y(_0585_),
    .A(\rf_shift_reg.rdata[3] ));
 sg13g2_inv_1 _2362_ (.Y(_0586_),
    .A(\rf_shift_reg.rdata[4] ));
 sg13g2_inv_2 _2363_ (.Y(_0587_),
    .A(\rf_shift_reg.rdata[5] ));
 sg13g2_inv_1 _2364_ (.Y(_0588_),
    .A(\cpu.alu.add_cy_r ));
 sg13g2_inv_1 _2365_ (.Y(_0589_),
    .A(\cpu.immdec.imm24_20[1] ));
 sg13g2_inv_1 _2366_ (.Y(_0590_),
    .A(net1248));
 sg13g2_inv_1 _2367_ (.Y(_0591_),
    .A(net1189));
 sg13g2_inv_1 _2368_ (.Y(_0592_),
    .A(net1272));
 sg13g2_inv_2 _2369_ (.Y(_0593_),
    .A(_0018_));
 sg13g2_inv_1 _2370_ (.Y(_0594_),
    .A(_0019_));
 sg13g2_inv_1 _2371_ (.Y(_0595_),
    .A(net1257));
 sg13g2_inv_1 _2372_ (.Y(_0596_),
    .A(net1198));
 sg13g2_inv_1 _2373_ (.Y(_0597_),
    .A(\cpu.bufreg2.dat[9] ));
 sg13g2_inv_1 _2374_ (.Y(_0598_),
    .A(net1228));
 sg13g2_inv_1 _2375_ (.Y(_0599_),
    .A(net1084));
 sg13g2_inv_1 _2376_ (.Y(_0600_),
    .A(net929));
 sg13g2_inv_1 _2377_ (.Y(_0601_),
    .A(net1196));
 sg13g2_inv_1 _2378_ (.Y(_0602_),
    .A(net1155));
 sg13g2_inv_1 _2379_ (.Y(_0603_),
    .A(net1069));
 sg13g2_inv_1 _2380_ (.Y(_0604_),
    .A(net1143));
 sg13g2_inv_1 _2381_ (.Y(_0605_),
    .A(net1176));
 sg13g2_inv_1 _2382_ (.Y(_0606_),
    .A(net1110));
 sg13g2_inv_1 _2383_ (.Y(_0607_),
    .A(net1283));
 sg13g2_inv_1 _2384_ (.Y(_0608_),
    .A(net1172));
 sg13g2_inv_1 _2385_ (.Y(_0609_),
    .A(net1267));
 sg13g2_inv_1 _2386_ (.Y(_0610_),
    .A(net1167));
 sg13g2_inv_1 _2387_ (.Y(_0611_),
    .A(net1202));
 sg13g2_inv_1 _2388_ (.Y(_0612_),
    .A(net1193));
 sg13g2_inv_1 _2389_ (.Y(_0613_),
    .A(net881));
 sg13g2_inv_1 _2390_ (.Y(_0614_),
    .A(net1188));
 sg13g2_inv_1 _2391_ (.Y(_0615_),
    .A(net1265));
 sg13g2_nor2_2 _2392_ (.A(_0465_),
    .B(net1156),
    .Y(_0616_));
 sg13g2_nand2b_2 _2393_ (.Y(_0617_),
    .B(net586),
    .A_N(net1156));
 sg13g2_and2_2 _2394_ (.A(net585),
    .B(net557),
    .X(_0618_));
 sg13g2_nand2_1 _2395_ (.Y(_0619_),
    .A(net580),
    .B(net555));
 sg13g2_nor3_1 _2396_ (.A(net819),
    .B(\cpu.state.cnt_r[0] ),
    .C(net771),
    .Y(_0620_));
 sg13g2_nor2b_1 _2397_ (.A(\cpu.state.cnt_r[3] ),
    .B_N(_0620_),
    .Y(_0621_));
 sg13g2_nand2_1 _2398_ (.Y(_0622_),
    .A(\cpu.state.init_done ),
    .B(net549));
 sg13g2_nor3_2 _2399_ (.A(net569),
    .B(net572),
    .C(_0622_),
    .Y(_0623_));
 sg13g2_a21oi_2 _2400_ (.B1(_0618_),
    .Y(_0624_),
    .A2(_0623_),
    .A1(_0020_));
 sg13g2_a21o_2 _2401_ (.A2(_0623_),
    .A1(_0020_),
    .B1(_0618_),
    .X(_0625_));
 sg13g2_mux2_2 _2402_ (.A0(_0058_),
    .A1(_0057_),
    .S(net551),
    .X(_0626_));
 sg13g2_xor2_1 _2403_ (.B(_0626_),
    .A(_0056_),
    .X(_0627_));
 sg13g2_nand3_1 _2404_ (.B(net752),
    .C(net557),
    .A(net585),
    .Y(_0628_));
 sg13g2_xor2_1 _2405_ (.B(_0628_),
    .A(\dut.rd_addr[1] ),
    .X(_0629_));
 sg13g2_nand3_1 _2406_ (.B(net557),
    .C(\cpu.ctrl.o_ibus_adr[0] ),
    .A(net585),
    .Y(_0630_));
 sg13g2_xor2_1 _2407_ (.B(_0630_),
    .A(\dut.rd_addr[0] ),
    .X(_0631_));
 sg13g2_nand2_2 _2408_ (.Y(_0632_),
    .A(_0629_),
    .B(_0631_));
 sg13g2_and3_1 _2409_ (.X(_0633_),
    .A(net580),
    .B(net555),
    .C(_0064_));
 sg13g2_a21oi_2 _2410_ (.B1(_0633_),
    .Y(_0634_),
    .A2(net551),
    .A1(_0063_));
 sg13g2_xnor2_1 _2411_ (.Y(_0635_),
    .A(_0062_),
    .B(_0634_));
 sg13g2_mux2_1 _2412_ (.A0(_0061_),
    .A1(_0060_),
    .S(net551),
    .X(_0636_));
 sg13g2_inv_1 _2413_ (.Y(_0637_),
    .A(_0636_));
 sg13g2_xor2_1 _2414_ (.B(_0636_),
    .A(_0059_),
    .X(_0638_));
 sg13g2_nor4_1 _2415_ (.A(_0627_),
    .B(_0632_),
    .C(_0635_),
    .D(_0638_),
    .Y(_0639_));
 sg13g2_and3_1 _2416_ (.X(_0640_),
    .A(net580),
    .B(net555),
    .C(_0085_));
 sg13g2_a21oi_2 _2417_ (.B1(_0640_),
    .Y(_0641_),
    .A2(net552),
    .A1(_0084_));
 sg13g2_xnor2_1 _2418_ (.Y(_0642_),
    .A(_0083_),
    .B(_0641_));
 sg13g2_and3_1 _2419_ (.X(_0643_),
    .A(net580),
    .B(net555),
    .C(_0070_));
 sg13g2_a21oi_2 _2420_ (.B1(_0643_),
    .Y(_0644_),
    .A2(net551),
    .A1(_0069_));
 sg13g2_xnor2_1 _2421_ (.Y(_0645_),
    .A(_0068_),
    .B(_0644_));
 sg13g2_mux2_2 _2422_ (.A0(_0067_),
    .A1(_0066_),
    .S(net551),
    .X(_0646_));
 sg13g2_inv_1 _2423_ (.Y(_0647_),
    .A(_0646_));
 sg13g2_xor2_1 _2424_ (.B(_0646_),
    .A(_0065_),
    .X(_0648_));
 sg13g2_mux2_2 _2425_ (.A0(_0037_),
    .A1(_0036_),
    .S(net553),
    .X(_0649_));
 sg13g2_xor2_1 _2426_ (.B(_0649_),
    .A(_0035_),
    .X(_0650_));
 sg13g2_nor4_1 _2427_ (.A(_0642_),
    .B(_0645_),
    .C(_0648_),
    .D(_0650_),
    .Y(_0651_));
 sg13g2_nand2_1 _2428_ (.Y(_0652_),
    .A(_0639_),
    .B(_0651_));
 sg13g2_mux2_2 _2429_ (.A0(_0025_),
    .A1(_0024_),
    .S(net554),
    .X(_0653_));
 sg13g2_nor2_1 _2430_ (.A(net568),
    .B(_0653_),
    .Y(_0654_));
 sg13g2_xor2_1 _2431_ (.B(_0653_),
    .A(net568),
    .X(_0655_));
 sg13g2_mux2_2 _2432_ (.A0(_0031_),
    .A1(_0030_),
    .S(net553),
    .X(_0656_));
 sg13g2_xnor2_1 _2433_ (.Y(_0657_),
    .A(_0029_),
    .B(_0656_));
 sg13g2_and3_1 _2434_ (.X(_0658_),
    .A(net585),
    .B(net557),
    .C(_0023_));
 sg13g2_a21oi_2 _2435_ (.B1(_0658_),
    .Y(_0659_),
    .A2(net554),
    .A1(_0022_));
 sg13g2_a21o_2 _2436_ (.A2(net553),
    .A1(_0022_),
    .B1(_0658_),
    .X(_0660_));
 sg13g2_a21oi_1 _2437_ (.A1(_0021_),
    .A2(_0659_),
    .Y(_0661_),
    .B1(_0546_));
 sg13g2_and3_1 _2438_ (.X(_0662_),
    .A(net581),
    .B(\cpu.state.ibus_cyc ),
    .C(_0034_));
 sg13g2_a21oi_2 _2439_ (.B1(_0662_),
    .Y(_0663_),
    .A2(net553),
    .A1(_0033_));
 sg13g2_a21o_2 _2440_ (.A2(net553),
    .A1(_0033_),
    .B1(_0662_),
    .X(_0664_));
 sg13g2_a22oi_1 _2441_ (.Y(_0665_),
    .B1(_0663_),
    .B2(_0032_),
    .A2(_0660_),
    .A1(_0565_));
 sg13g2_and4_1 _2442_ (.A(_0655_),
    .B(_0657_),
    .C(_0661_),
    .D(_0665_),
    .X(_0666_));
 sg13g2_a21o_1 _2443_ (.A2(net556),
    .A1(net581),
    .B1(_0045_),
    .X(_0667_));
 sg13g2_nand3b_1 _2444_ (.B(net556),
    .C(net581),
    .Y(_0668_),
    .A_N(_0046_));
 sg13g2_nand2_1 _2445_ (.Y(_0669_),
    .A(_0667_),
    .B(_0668_));
 sg13g2_and3_1 _2446_ (.X(_0670_),
    .A(_0044_),
    .B(_0667_),
    .C(_0668_));
 sg13g2_a21oi_1 _2447_ (.A1(_0667_),
    .A2(_0668_),
    .Y(_0671_),
    .B1(_0044_));
 sg13g2_nor2_1 _2448_ (.A(_0670_),
    .B(_0671_),
    .Y(_0672_));
 sg13g2_a21o_1 _2449_ (.A2(net556),
    .A1(net581),
    .B1(_0048_),
    .X(_0673_));
 sg13g2_nand3b_1 _2450_ (.B(net555),
    .C(net580),
    .Y(_0674_),
    .A_N(_0049_));
 sg13g2_nand2_2 _2451_ (.Y(_0675_),
    .A(_0673_),
    .B(_0674_));
 sg13g2_and3_1 _2452_ (.X(_0676_),
    .A(_0047_),
    .B(_0673_),
    .C(_0674_));
 sg13g2_a21oi_2 _2453_ (.B1(_0047_),
    .Y(_0677_),
    .A2(_0674_),
    .A1(_0673_));
 sg13g2_nor2_1 _2454_ (.A(_0676_),
    .B(_0677_),
    .Y(_0678_));
 sg13g2_nor2_1 _2455_ (.A(_0032_),
    .B(_0663_),
    .Y(_0679_));
 sg13g2_mux2_2 _2456_ (.A0(_0028_),
    .A1(_0027_),
    .S(net553),
    .X(_0680_));
 sg13g2_and2_1 _2457_ (.A(_0566_),
    .B(_0680_),
    .X(_0681_));
 sg13g2_or2_1 _2458_ (.X(_0682_),
    .B(_0680_),
    .A(_0566_));
 sg13g2_xnor2_1 _2459_ (.Y(_0683_),
    .A(_0566_),
    .B(_0680_));
 sg13g2_nor4_1 _2460_ (.A(_0672_),
    .B(_0678_),
    .C(_0679_),
    .D(_0683_),
    .Y(_0684_));
 sg13g2_mux2_2 _2461_ (.A0(_0073_),
    .A1(_0072_),
    .S(net552),
    .X(_0685_));
 sg13g2_xor2_1 _2462_ (.B(_0685_),
    .A(_0071_),
    .X(_0686_));
 sg13g2_and3_1 _2463_ (.X(_0687_),
    .A(net581),
    .B(net557),
    .C(_0040_));
 sg13g2_a21oi_2 _2464_ (.B1(_0687_),
    .Y(_0688_),
    .A2(net553),
    .A1(_0039_));
 sg13g2_xnor2_1 _2465_ (.Y(_0689_),
    .A(_0038_),
    .B(_0688_));
 sg13g2_and3_1 _2466_ (.X(_0690_),
    .A(net580),
    .B(net555),
    .C(_0055_));
 sg13g2_a21oi_2 _2467_ (.B1(_0690_),
    .Y(_0691_),
    .A2(net551),
    .A1(_0054_));
 sg13g2_xnor2_1 _2468_ (.Y(_0692_),
    .A(_0053_),
    .B(_0691_));
 sg13g2_and3_1 _2469_ (.X(_0693_),
    .A(net580),
    .B(net555),
    .C(_0052_));
 sg13g2_a21oi_2 _2470_ (.B1(_0693_),
    .Y(_0694_),
    .A2(net551),
    .A1(_0051_));
 sg13g2_xnor2_1 _2471_ (.Y(_0695_),
    .A(_0050_),
    .B(_0694_));
 sg13g2_nor4_1 _2472_ (.A(_0686_),
    .B(_0689_),
    .C(_0692_),
    .D(_0695_),
    .Y(_0696_));
 sg13g2_mux2_2 _2473_ (.A0(_0076_),
    .A1(_0075_),
    .S(net552),
    .X(_0697_));
 sg13g2_xor2_1 _2474_ (.B(_0697_),
    .A(_0074_),
    .X(_0698_));
 sg13g2_and2_1 _2475_ (.A(_0082_),
    .B(_0618_),
    .X(_0699_));
 sg13g2_a21oi_1 _2476_ (.A1(_0081_),
    .A2(net552),
    .Y(_0700_),
    .B1(_0699_));
 sg13g2_mux2_1 _2477_ (.A0(_0082_),
    .A1(_0081_),
    .S(net552),
    .X(_0701_));
 sg13g2_xor2_1 _2478_ (.B(_0701_),
    .A(_0080_),
    .X(_0702_));
 sg13g2_and3_1 _2479_ (.X(_0703_),
    .A(net580),
    .B(net555),
    .C(_0079_));
 sg13g2_a21oi_2 _2480_ (.B1(_0703_),
    .Y(_0704_),
    .A2(net551),
    .A1(_0078_));
 sg13g2_xnor2_1 _2481_ (.Y(_0705_),
    .A(_0077_),
    .B(_0704_));
 sg13g2_and3_1 _2482_ (.X(_0706_),
    .A(net581),
    .B(net556),
    .C(_0043_));
 sg13g2_a21oi_2 _2483_ (.B1(_0706_),
    .Y(_0707_),
    .A2(net553),
    .A1(_0042_));
 sg13g2_xnor2_1 _2484_ (.Y(_0708_),
    .A(_0041_),
    .B(_0707_));
 sg13g2_nor4_1 _2485_ (.A(_0698_),
    .B(_0702_),
    .C(_0705_),
    .D(_0708_),
    .Y(_0709_));
 sg13g2_nand4_1 _2486_ (.B(_0684_),
    .C(_0696_),
    .A(_0666_),
    .Y(_0710_),
    .D(_0709_));
 sg13g2_nor3_2 _2487_ (.A(_0624_),
    .B(_0652_),
    .C(_0710_),
    .Y(_0711_));
 sg13g2_o21ai_1 _2488_ (.B1(\dut.rd_valid ),
    .Y(_0712_),
    .A1(_0567_),
    .A2(_0656_));
 sg13g2_xnor2_1 _2489_ (.Y(_0713_),
    .A(_0021_),
    .B(_0659_));
 sg13g2_nor4_1 _2490_ (.A(_0648_),
    .B(_0698_),
    .C(_0705_),
    .D(_0712_),
    .Y(_0714_));
 sg13g2_nor3_1 _2491_ (.A(_0650_),
    .B(_0654_),
    .C(_0679_),
    .Y(_0715_));
 sg13g2_a22oi_1 _2492_ (.Y(_0716_),
    .B1(_0663_),
    .B2(_0032_),
    .A2(_0653_),
    .A1(net568));
 sg13g2_a22oi_1 _2493_ (.Y(_0717_),
    .B1(_0688_),
    .B2(_0038_),
    .A2(_0656_),
    .A1(_0567_));
 sg13g2_nand4_1 _2494_ (.B(_0715_),
    .C(_0716_),
    .A(_0714_),
    .Y(_0718_),
    .D(_0717_));
 sg13g2_o21ai_1 _2495_ (.B1(_0682_),
    .Y(_0719_),
    .A1(_0038_),
    .A2(_0688_));
 sg13g2_or4_1 _2496_ (.A(_0642_),
    .B(_0681_),
    .C(_0702_),
    .D(_0719_),
    .X(_0720_));
 sg13g2_nor4_1 _2497_ (.A(_0627_),
    .B(_0645_),
    .C(_0686_),
    .D(_0713_),
    .Y(_0721_));
 sg13g2_nor4_1 _2498_ (.A(_0632_),
    .B(_0635_),
    .C(_0692_),
    .D(_0708_),
    .Y(_0722_));
 sg13g2_nor4_1 _2499_ (.A(_0638_),
    .B(_0672_),
    .C(_0678_),
    .D(_0695_),
    .Y(_0723_));
 sg13g2_nand3_1 _2500_ (.B(_0722_),
    .C(_0723_),
    .A(_0721_),
    .Y(_0724_));
 sg13g2_nor4_2 _2501_ (.A(_0624_),
    .B(_0718_),
    .C(_0720_),
    .Y(_0725_),
    .D(_0724_));
 sg13g2_o21ai_1 _2502_ (.B1(_0625_),
    .Y(_0726_),
    .A1(_0652_),
    .A2(_0710_));
 sg13g2_inv_1 _2503_ (.Y(_0727_),
    .A(_0726_));
 sg13g2_or2_1 _2504_ (.X(_0728_),
    .B(_0726_),
    .A(_0546_));
 sg13g2_nand2_1 _2505_ (.Y(_0729_),
    .A(\dut.rd_addr[2] ),
    .B(net568));
 sg13g2_and4_1 _2506_ (.A(\dut.rd_addr[2] ),
    .B(net568),
    .C(\dut.rd_addr[4] ),
    .D(\dut.rd_addr[5] ),
    .X(_0730_));
 sg13g2_nand4_1 _2507_ (.B(\dut.rd_addr[3] ),
    .C(\dut.rd_addr[4] ),
    .A(\dut.rd_addr[2] ),
    .Y(_0731_),
    .D(\dut.rd_addr[5] ));
 sg13g2_and2_1 _2508_ (.A(\dut.rd_addr[6] ),
    .B(\dut.rd_addr[7] ),
    .X(_0732_));
 sg13g2_nand2_2 _2509_ (.Y(_0733_),
    .A(\dut.rd_addr[6] ),
    .B(\dut.rd_addr[7] ));
 sg13g2_nor2_1 _2510_ (.A(_0731_),
    .B(_0733_),
    .Y(_0734_));
 sg13g2_and2_1 _2511_ (.A(\dut.rd_addr[8] ),
    .B(\dut.rd_addr[9] ),
    .X(_0735_));
 sg13g2_nand2_1 _2512_ (.Y(_0736_),
    .A(\dut.rd_addr[8] ),
    .B(\dut.rd_addr[9] ));
 sg13g2_nor3_1 _2513_ (.A(_0731_),
    .B(_0733_),
    .C(_0736_),
    .Y(_0737_));
 sg13g2_nand2_1 _2514_ (.Y(_0738_),
    .A(_0734_),
    .B(_0735_));
 sg13g2_and2_1 _2515_ (.A(\dut.rd_addr[10] ),
    .B(\dut.rd_addr[11] ),
    .X(_0739_));
 sg13g2_and4_2 _2516_ (.A(_0730_),
    .B(_0732_),
    .C(_0735_),
    .D(_0739_),
    .X(_0740_));
 sg13g2_nand4_1 _2517_ (.B(_0732_),
    .C(_0735_),
    .A(_0730_),
    .Y(_0741_),
    .D(_0739_));
 sg13g2_and2_1 _2518_ (.A(\dut.rd_addr[12] ),
    .B(\dut.rd_addr[13] ),
    .X(_0742_));
 sg13g2_nand2_1 _2519_ (.Y(_0743_),
    .A(\dut.rd_addr[12] ),
    .B(\dut.rd_addr[13] ));
 sg13g2_nand2_1 _2520_ (.Y(_0744_),
    .A(_0740_),
    .B(_0742_));
 sg13g2_nand2_1 _2521_ (.Y(_0745_),
    .A(\dut.rd_addr[14] ),
    .B(\dut.rd_addr[15] ));
 sg13g2_nor3_2 _2522_ (.A(_0741_),
    .B(_0743_),
    .C(_0745_),
    .Y(_0746_));
 sg13g2_nand2_1 _2523_ (.Y(_0747_),
    .A(\dut.rd_addr[16] ),
    .B(\dut.rd_addr[17] ));
 sg13g2_or4_2 _2524_ (.A(_0741_),
    .B(_0743_),
    .C(_0745_),
    .D(_0747_),
    .X(_0748_));
 sg13g2_nand2_2 _2525_ (.Y(_0749_),
    .A(\dut.rd_addr[18] ),
    .B(\dut.rd_addr[19] ));
 sg13g2_nor2_1 _2526_ (.A(_0748_),
    .B(_0749_),
    .Y(_0750_));
 sg13g2_nand2_1 _2527_ (.Y(_0751_),
    .A(\dut.rd_addr[20] ),
    .B(\dut.rd_addr[21] ));
 sg13g2_nor3_2 _2528_ (.A(_0748_),
    .B(_0749_),
    .C(_0751_),
    .Y(_0752_));
 sg13g2_nand3_1 _2529_ (.B(\dut.rd_addr[23] ),
    .C(_0752_),
    .A(\dut.rd_addr[22] ),
    .Y(_0753_));
 sg13g2_nand2b_1 _2530_ (.Y(_0754_),
    .B(_0752_),
    .A_N(_0702_));
 sg13g2_nor3_2 _2531_ (.A(_0074_),
    .B(_0748_),
    .C(_0749_),
    .Y(_0755_));
 sg13g2_nor2b_2 _2532_ (.A(_0062_),
    .B_N(_0746_),
    .Y(_0756_));
 sg13g2_xnor2_1 _2533_ (.Y(_0757_),
    .A(_0648_),
    .B(_0756_));
 sg13g2_nor3_2 _2534_ (.A(_0038_),
    .B(_0731_),
    .C(_0733_),
    .Y(_0758_));
 sg13g2_xor2_1 _2535_ (.B(_0758_),
    .A(_0708_),
    .X(_0759_));
 sg13g2_nor2_2 _2536_ (.A(_0050_),
    .B(_0741_),
    .Y(_0760_));
 sg13g2_nor2_1 _2537_ (.A(_0032_),
    .B(_0731_),
    .Y(_0761_));
 sg13g2_xor2_1 _2538_ (.B(_0761_),
    .A(_0035_),
    .X(_0762_));
 sg13g2_xnor2_1 _2539_ (.Y(_0763_),
    .A(_0650_),
    .B(_0761_));
 sg13g2_xor2_1 _2540_ (.B(_0734_),
    .A(_0038_),
    .X(_0764_));
 sg13g2_xnor2_1 _2541_ (.Y(_0765_),
    .A(_0688_),
    .B(_0764_));
 sg13g2_nor4_2 _2542_ (.A(_0080_),
    .B(_0748_),
    .C(_0749_),
    .Y(_0766_),
    .D(_0751_));
 sg13g2_nor2b_1 _2543_ (.A(_0766_),
    .B_N(_0642_),
    .Y(_0767_));
 sg13g2_o21ai_1 _2544_ (.B1(_0752_),
    .Y(_0768_),
    .A1(_0080_),
    .A2(_0642_));
 sg13g2_a21o_1 _2545_ (.A2(_0768_),
    .A1(_0702_),
    .B1(_0767_),
    .X(_0769_));
 sg13g2_xnor2_1 _2546_ (.Y(_0770_),
    .A(_0645_),
    .B(_0748_));
 sg13g2_nor2_2 _2547_ (.A(_0068_),
    .B(_0748_),
    .Y(_0771_));
 sg13g2_xnor2_1 _2548_ (.Y(_0772_),
    .A(_0686_),
    .B(_0771_));
 sg13g2_nor4_2 _2549_ (.A(_0044_),
    .B(_0731_),
    .C(_0733_),
    .Y(_0773_),
    .D(_0736_));
 sg13g2_nor3_1 _2550_ (.A(_0676_),
    .B(_0677_),
    .C(_0773_),
    .Y(_0774_));
 sg13g2_a21oi_1 _2551_ (.A1(_0672_),
    .A2(_0738_),
    .Y(_0775_),
    .B1(_0774_));
 sg13g2_nand3b_1 _2552_ (.B(_0740_),
    .C(_0742_),
    .Y(_0776_),
    .A_N(_0056_));
 sg13g2_nor2_1 _2553_ (.A(_0638_),
    .B(_0776_),
    .Y(_0777_));
 sg13g2_xnor2_1 _2554_ (.Y(_0778_),
    .A(_0695_),
    .B(_0740_));
 sg13g2_xnor2_1 _2555_ (.Y(_0779_),
    .A(_0032_),
    .B(_0731_));
 sg13g2_xnor2_1 _2556_ (.Y(_0780_),
    .A(_0664_),
    .B(_0779_));
 sg13g2_xnor2_1 _2557_ (.Y(_0781_),
    .A(\dut.rd_addr[2] ),
    .B(_0659_));
 sg13g2_xor2_1 _2558_ (.B(net568),
    .A(\dut.rd_addr[2] ),
    .X(_0782_));
 sg13g2_xnor2_1 _2559_ (.Y(_0783_),
    .A(_0653_),
    .B(_0782_));
 sg13g2_nand3b_1 _2560_ (.B(net568),
    .C(\dut.rd_addr[2] ),
    .Y(_0784_),
    .A_N(_0026_));
 sg13g2_xnor2_1 _2561_ (.Y(_0785_),
    .A(_0029_),
    .B(_0784_));
 sg13g2_xnor2_1 _2562_ (.Y(_0786_),
    .A(_0566_),
    .B(_0729_));
 sg13g2_xnor2_1 _2563_ (.Y(_0787_),
    .A(_0680_),
    .B(_0786_));
 sg13g2_and2_1 _2564_ (.A(_0638_),
    .B(_0776_),
    .X(_0788_));
 sg13g2_xnor2_1 _2565_ (.Y(_0789_),
    .A(_0698_),
    .B(_0750_));
 sg13g2_xor2_1 _2566_ (.B(_0746_),
    .A(_0635_),
    .X(_0790_));
 sg13g2_xnor2_1 _2567_ (.Y(_0791_),
    .A(_0656_),
    .B(_0785_));
 sg13g2_xnor2_1 _2568_ (.Y(_0792_),
    .A(_0627_),
    .B(_0744_));
 sg13g2_xnor2_1 _2569_ (.Y(_0793_),
    .A(_0705_),
    .B(_0755_));
 sg13g2_nand4_1 _2570_ (.B(_0754_),
    .C(_0772_),
    .A(_0753_),
    .Y(_0794_),
    .D(_0793_));
 sg13g2_nor2_1 _2571_ (.A(_0770_),
    .B(_0790_),
    .Y(_0795_));
 sg13g2_o21ai_1 _2572_ (.B1(_0737_),
    .Y(_0796_),
    .A1(_0670_),
    .A2(_0671_));
 sg13g2_o21ai_1 _2573_ (.B1(_0773_),
    .Y(_0797_),
    .A1(_0676_),
    .A2(_0677_));
 sg13g2_nand4_1 _2574_ (.B(_0791_),
    .C(_0796_),
    .A(_0780_),
    .Y(_0798_),
    .D(_0797_));
 sg13g2_xor2_1 _2575_ (.B(_0760_),
    .A(_0692_),
    .X(_0799_));
 sg13g2_nor4_1 _2576_ (.A(_0777_),
    .B(_0788_),
    .C(_0798_),
    .D(_0799_),
    .Y(_0800_));
 sg13g2_nor3_1 _2577_ (.A(_0759_),
    .B(_0765_),
    .C(_0792_),
    .Y(_0801_));
 sg13g2_nor4_1 _2578_ (.A(_0632_),
    .B(_0781_),
    .C(_0783_),
    .D(_0787_),
    .Y(_0802_));
 sg13g2_and4_1 _2579_ (.A(_0763_),
    .B(_0775_),
    .C(_0778_),
    .D(_0802_),
    .X(_0803_));
 sg13g2_nand4_1 _2580_ (.B(_0800_),
    .C(_0801_),
    .A(_0795_),
    .Y(_0804_),
    .D(_0803_));
 sg13g2_nand2_1 _2581_ (.Y(_0805_),
    .A(_0757_),
    .B(_0789_));
 sg13g2_nor4_2 _2582_ (.A(_0769_),
    .B(_0794_),
    .C(_0804_),
    .Y(_0806_),
    .D(_0805_));
 sg13g2_nor2_1 _2583_ (.A(_0728_),
    .B(_0806_),
    .Y(_0807_));
 sg13g2_o21ai_1 _2584_ (.B1(_0616_),
    .Y(_0808_),
    .A1(_0728_),
    .A2(_0806_));
 sg13g2_nor4_2 _2585_ (.A(\dut.xfer.count[3] ),
    .B(\dut.xfer.count[2] ),
    .C(\dut.xfer.count[1] ),
    .Y(_0809_),
    .D(\dut.xfer.count[0] ));
 sg13g2_or2_1 _2586_ (.X(_0810_),
    .B(_0809_),
    .A(\dut.xfer.count[0] ));
 sg13g2_nor3_1 _2587_ (.A(\dut.xfer.count[1] ),
    .B(\dut.xfer.count[0] ),
    .C(_0809_),
    .Y(_0811_));
 sg13g2_nor4_2 _2588_ (.A(\dut.xfer.count[1] ),
    .B(\dut.xfer.count[0] ),
    .C(_0568_),
    .Y(_0812_),
    .D(_0809_));
 sg13g2_a21oi_1 _2589_ (.A1(net567),
    .A2(_0812_),
    .Y(_0813_),
    .B1(_0547_));
 sg13g2_nand3_1 _2590_ (.B(net567),
    .C(_0812_),
    .A(_0547_),
    .Y(_0814_));
 sg13g2_nor4_2 _2591_ (.A(net1241),
    .B(net1274),
    .C(\dut.xfer.dummy_count[1] ),
    .Y(_0815_),
    .D(\dut.xfer.dummy_count[0] ));
 sg13g2_or4_2 _2592_ (.A(\dut.xfer.dummy_count[3] ),
    .B(\dut.xfer.dummy_count[2] ),
    .C(\dut.xfer.dummy_count[1] ),
    .D(\dut.xfer.dummy_count[0] ),
    .X(_0816_));
 sg13g2_nand3b_1 _2593_ (.B(_0814_),
    .C(_0815_),
    .Y(_0817_),
    .A_N(_0813_));
 sg13g2_inv_1 _2594_ (.Y(_0818_),
    .A(_0817_));
 sg13g2_xnor2_1 _2595_ (.Y(_0819_),
    .A(_0088_),
    .B(_0811_));
 sg13g2_mux2_1 _2596_ (.A0(net809),
    .A1(_0819_),
    .S(\dut.flash_clk ),
    .X(_0820_));
 sg13g2_nor2_1 _2597_ (.A(\dut.flash_clk ),
    .B(net778),
    .Y(_0821_));
 sg13g2_a21oi_1 _2598_ (.A1(\dut.flash_clk ),
    .A2(_0810_),
    .Y(_0822_),
    .B1(_0821_));
 sg13g2_nor4_2 _2599_ (.A(net746),
    .B(_0817_),
    .C(_0820_),
    .Y(_0823_),
    .D(_0822_));
 sg13g2_nor2_1 _2600_ (.A(\dut.xfer.fetch ),
    .B(net1311),
    .Y(_0824_));
 sg13g2_and2_2 _2601_ (.A(_0823_),
    .B(net1312),
    .X(_0825_));
 sg13g2_or2_1 _2602_ (.X(_0826_),
    .B(_0825_),
    .A(_0808_));
 sg13g2_and3_1 _2603_ (.X(_0827_),
    .A(\dut.xfer.resetn ),
    .B(\dut.din_valid ),
    .C(_0823_));
 sg13g2_nand3_1 _2604_ (.B(\dut.din_valid ),
    .C(_0823_),
    .A(net558),
    .Y(_0828_));
 sg13g2_nor2_1 _2605_ (.A(_0808_),
    .B(net533),
    .Y(_0829_));
 sg13g2_nand2_1 _2606_ (.Y(_0830_),
    .A(net794),
    .B(net441));
 sg13g2_o21ai_1 _2607_ (.B1(_0830_),
    .Y(_0010_),
    .A1(_0569_),
    .A2(_0826_));
 sg13g2_nand3b_1 _2608_ (.B(net533),
    .C(_0616_),
    .Y(_0831_),
    .A_N(_0807_));
 sg13g2_nand2_1 _2609_ (.Y(_0832_),
    .A(net578),
    .B(_0727_));
 sg13g2_nand3_1 _2610_ (.B(_0727_),
    .C(net441),
    .A(net1191),
    .Y(_0833_));
 sg13g2_o21ai_1 _2611_ (.B1(_0833_),
    .Y(_0009_),
    .A1(_0560_),
    .A2(_0831_));
 sg13g2_o21ai_1 _2612_ (.B1(_0616_),
    .Y(_0001_),
    .A1(_0558_),
    .A2(_0831_));
 sg13g2_nand2_1 _2613_ (.Y(_0834_),
    .A(net1178),
    .B(_0829_));
 sg13g2_o21ai_1 _2614_ (.B1(_0834_),
    .Y(_0003_),
    .A1(_0570_),
    .A2(_0831_));
 sg13g2_nand2_1 _2615_ (.Y(_0835_),
    .A(net1184),
    .B(net441));
 sg13g2_o21ai_1 _2616_ (.B1(_0835_),
    .Y(_0002_),
    .A1(_0571_),
    .A2(_0826_));
 sg13g2_nand2_1 _2617_ (.Y(_0836_),
    .A(\dut.state[9] ),
    .B(_0726_));
 sg13g2_nand3_1 _2618_ (.B(_0616_),
    .C(_0726_),
    .A(net578),
    .Y(_0837_));
 sg13g2_o21ai_1 _2619_ (.B1(_0837_),
    .Y(_0838_),
    .A1(_0831_),
    .A2(_0832_));
 sg13g2_a21o_1 _2620_ (.A2(net441),
    .A1(net1271),
    .B1(_0838_),
    .X(_0012_));
 sg13g2_nor2b_1 _2621_ (.A(_0808_),
    .B_N(_0825_),
    .Y(_0839_));
 sg13g2_nand2_1 _2622_ (.Y(_0840_),
    .A(net1098),
    .B(_0839_));
 sg13g2_o21ai_1 _2623_ (.B1(_0616_),
    .Y(_0841_),
    .A1(net1271),
    .A2(_0807_));
 sg13g2_nor2_1 _2624_ (.A(_0807_),
    .B(net532),
    .Y(_0842_));
 sg13g2_o21ai_1 _2625_ (.B1(_0840_),
    .Y(_0005_),
    .A1(_0841_),
    .A2(_0842_));
 sg13g2_nand2_1 _2626_ (.Y(_0843_),
    .A(net1232),
    .B(net532));
 sg13g2_nand2_1 _2627_ (.Y(_0844_),
    .A(net579),
    .B(net441));
 sg13g2_o21ai_1 _2628_ (.B1(_0844_),
    .Y(_0004_),
    .A1(_0808_),
    .A2(_0843_));
 sg13g2_o21ai_1 _2629_ (.B1(net1246),
    .Y(_0845_),
    .A1(_0573_),
    .A2(_0625_));
 sg13g2_inv_1 _2630_ (.Y(_0846_),
    .A(_0845_));
 sg13g2_nor2_1 _2631_ (.A(net1299),
    .B(net1232),
    .Y(_0847_));
 sg13g2_nand2_1 _2632_ (.Y(_0848_),
    .A(_0845_),
    .B(_0847_));
 sg13g2_nand2_1 _2633_ (.Y(_0849_),
    .A(_0829_),
    .B(_0848_));
 sg13g2_o21ai_1 _2634_ (.B1(_0849_),
    .Y(_0011_),
    .A1(_0572_),
    .A2(_0831_));
 sg13g2_nand2_1 _2635_ (.Y(_0850_),
    .A(net854),
    .B(net441));
 sg13g2_o21ai_1 _2636_ (.B1(_0850_),
    .Y(_0008_),
    .A1(_0561_),
    .A2(_0831_));
 sg13g2_nand2_1 _2637_ (.Y(_0851_),
    .A(net720),
    .B(_0839_));
 sg13g2_o21ai_1 _2638_ (.B1(_0851_),
    .Y(_0007_),
    .A1(_0559_),
    .A2(_0831_));
 sg13g2_nand3_1 _2639_ (.B(\dut.state[3] ),
    .C(_0624_),
    .A(net1215),
    .Y(_0852_));
 sg13g2_or2_1 _2640_ (.X(_0853_),
    .B(_0852_),
    .A(_0617_));
 sg13g2_o21ai_1 _2641_ (.B1(_0853_),
    .Y(_0854_),
    .A1(_0831_),
    .A2(_0845_));
 sg13g2_a21o_1 _2642_ (.A2(net441),
    .A1(net1237),
    .B1(_0854_),
    .X(_0006_));
 sg13g2_nor2_1 _2643_ (.A(net577),
    .B(\cpu.bne_or_bge ),
    .Y(_0855_));
 sg13g2_nand2_1 _2644_ (.Y(_0856_),
    .A(_0090_),
    .B(_0855_));
 sg13g2_a21oi_1 _2645_ (.A1(net1335),
    .A2(net1248),
    .Y(_0857_),
    .B1(_0856_));
 sg13g2_a22oi_1 _2646_ (.Y(_0858_),
    .B1(_0587_),
    .B2(\cpu.immdec.imm19_12_20[6] ),
    .A2(\cpu.immdec.imm19_12_20[5] ),
    .A1(_0585_));
 sg13g2_nand2b_1 _2647_ (.Y(_0859_),
    .B(\cpu.csr_imm ),
    .A_N(_0858_));
 sg13g2_a21oi_1 _2648_ (.A1(\cpu.csr_imm ),
    .A2(\rf_shift_reg.rdata[1] ),
    .Y(_0860_),
    .B1(\cpu.immdec.imm19_12_20[5] ));
 sg13g2_nor2_1 _2649_ (.A(\cpu.csr_imm ),
    .B(\rf_shift_reg.rdata[2] ),
    .Y(_0861_));
 sg13g2_nor3_1 _2650_ (.A(\cpu.immdec.imm19_12_20[6] ),
    .B(_0860_),
    .C(_0861_),
    .Y(_0862_));
 sg13g2_o21ai_1 _2651_ (.B1(\cpu.immdec.imm19_12_20[6] ),
    .Y(_0863_),
    .A1(\cpu.csr_imm ),
    .A2(\rf_shift_reg.rdata[4] ));
 sg13g2_nor2_1 _2652_ (.A(\cpu.immdec.imm19_12_20[5] ),
    .B(_0863_),
    .Y(_0864_));
 sg13g2_o21ai_1 _2653_ (.B1(_0859_),
    .Y(_0865_),
    .A1(_0862_),
    .A2(_0864_));
 sg13g2_nor2_1 _2654_ (.A(_0588_),
    .B(_0865_),
    .Y(_0866_));
 sg13g2_xnor2_1 _2655_ (.Y(_0867_),
    .A(_0588_),
    .B(_0865_));
 sg13g2_o21ai_1 _2656_ (.B1(\cpu.immdec.imm24_20[2] ),
    .Y(_0868_),
    .A1(\cpu.immdec.imm24_20[0] ),
    .A2(\rf_shift_reg.rdata[4] ));
 sg13g2_a21oi_1 _2657_ (.A1(\cpu.immdec.imm24_20[0] ),
    .A2(_0587_),
    .Y(_0869_),
    .B1(_0868_));
 sg13g2_nor3_1 _2658_ (.A(_0583_),
    .B(_0584_),
    .C(\cpu.immdec.imm24_20[2] ),
    .Y(_0870_));
 sg13g2_o21ai_1 _2659_ (.B1(_0589_),
    .Y(_0871_),
    .A1(_0869_),
    .A2(_0870_));
 sg13g2_nor2_1 _2660_ (.A(\cpu.immdec.imm24_20[0] ),
    .B(\rf_shift_reg.rdata[2] ),
    .Y(_0872_));
 sg13g2_nor3_1 _2661_ (.A(_0589_),
    .B(\cpu.immdec.imm24_20[2] ),
    .C(_0872_),
    .Y(_0873_));
 sg13g2_o21ai_1 _2662_ (.B1(_0873_),
    .Y(_0874_),
    .A1(_0583_),
    .A2(\rf_shift_reg.rdata[3] ));
 sg13g2_and3_1 _2663_ (.X(_0875_),
    .A(\cpu.bufreg2.i_op_b_sel ),
    .B(_0871_),
    .C(_0874_));
 sg13g2_nand3_1 _2664_ (.B(_0871_),
    .C(_0874_),
    .A(net571),
    .Y(_0876_));
 sg13g2_nand3_1 _2665_ (.B(\cpu.state.o_cnt[2] ),
    .C(net1292),
    .A(net1211),
    .Y(_0877_));
 sg13g2_or2_2 _2666_ (.X(_0878_),
    .B(_0877_),
    .A(_0574_));
 sg13g2_inv_1 _2667_ (.Y(_0879_),
    .A(_0878_));
 sg13g2_nand2_1 _2668_ (.Y(_0880_),
    .A(net570),
    .B(net573));
 sg13g2_or2_1 _2669_ (.X(_0881_),
    .B(_0880_),
    .A(_0017_));
 sg13g2_o21ai_1 _2670_ (.B1(net995),
    .Y(_0882_),
    .A1(_0017_),
    .A2(_0880_));
 sg13g2_nor2_2 _2671_ (.A(net575),
    .B(\cpu.decode.opcode[1] ),
    .Y(_0883_));
 sg13g2_nor2b_1 _2672_ (.A(net573),
    .B_N(net571),
    .Y(_0884_));
 sg13g2_nor2_1 _2673_ (.A(net572),
    .B(net574),
    .Y(_0885_));
 sg13g2_and3_1 _2674_ (.X(_0886_),
    .A(\cpu.immdec.imm11_7[0] ),
    .B(_0883_),
    .C(_0884_));
 sg13g2_a21oi_1 _2675_ (.A1(_0883_),
    .A2(_0884_),
    .Y(_0887_),
    .B1(_0583_));
 sg13g2_o21ai_1 _2676_ (.B1(_0878_),
    .Y(_0888_),
    .A1(_0886_),
    .A2(_0887_));
 sg13g2_or2_1 _2677_ (.X(_0889_),
    .B(_0882_),
    .A(_0878_));
 sg13g2_and2_1 _2678_ (.A(_0888_),
    .B(_0889_),
    .X(_0890_));
 sg13g2_and3_1 _2679_ (.X(_0891_),
    .A(_0563_),
    .B(_0888_),
    .C(_0889_));
 sg13g2_nand3_1 _2680_ (.B(_0888_),
    .C(_0889_),
    .A(_0563_),
    .Y(_0892_));
 sg13g2_nor3_1 _2681_ (.A(_0857_),
    .B(_0875_),
    .C(_0891_),
    .Y(_0893_));
 sg13g2_a221oi_1 _2682_ (.B2(_0892_),
    .C1(_0856_),
    .B1(_0876_),
    .A1(net571),
    .Y(_0894_),
    .A2(\cpu.bufreg.i_sh_signed ));
 sg13g2_nor3_2 _2683_ (.A(_0867_),
    .B(_0893_),
    .C(_0894_),
    .Y(_0895_));
 sg13g2_nor3_1 _2684_ (.A(net550),
    .B(_0866_),
    .C(_0895_),
    .Y(_0896_));
 sg13g2_a21oi_1 _2685_ (.A1(net550),
    .A2(net1336),
    .Y(_0013_),
    .B1(_0896_));
 sg13g2_and2_1 _2686_ (.A(net577),
    .B(net576),
    .X(_0897_));
 sg13g2_nor4_1 _2687_ (.A(net574),
    .B(_0576_),
    .C(_0855_),
    .D(_0897_),
    .Y(_0898_));
 sg13g2_nand2b_1 _2688_ (.Y(_0899_),
    .B(net572),
    .A_N(_0898_));
 sg13g2_nand2_2 _2689_ (.Y(_0900_),
    .A(net1320),
    .B(_0899_));
 sg13g2_nand2b_2 _2690_ (.Y(_0901_),
    .B(_0900_),
    .A_N(net549));
 sg13g2_nand2_1 _2691_ (.Y(_0902_),
    .A(\cpu.ctrl.o_ibus_adr[0] ),
    .B(net1129));
 sg13g2_nor3_2 _2692_ (.A(\cpu.state.o_cnt[2] ),
    .B(\cpu.mem_bytecnt[0] ),
    .C(\cpu.mem_bytecnt[1] ),
    .Y(_0903_));
 sg13g2_xor2_1 _2693_ (.B(net1129),
    .A(\cpu.ctrl.o_ibus_adr[0] ),
    .X(_0904_));
 sg13g2_nand3_1 _2694_ (.B(_0903_),
    .C(_0904_),
    .A(net771),
    .Y(_0905_));
 sg13g2_a21oi_1 _2695_ (.A1(net1130),
    .A2(_0905_),
    .Y(_0015_),
    .B1(_0901_));
 sg13g2_nand2_1 _2696_ (.Y(_0906_),
    .A(_0092_),
    .B(_0883_));
 sg13g2_nand3_1 _2697_ (.B(net573),
    .C(\cpu.decode.co_ebreak ),
    .A(net570),
    .Y(_0907_));
 sg13g2_nand2_1 _2698_ (.Y(_0908_),
    .A(net575),
    .B(\cpu.decode.opcode[1] ));
 sg13g2_or2_1 _2699_ (.X(_0909_),
    .B(net570),
    .A(net571));
 sg13g2_nand4_1 _2700_ (.B(_0907_),
    .C(_0908_),
    .A(_0906_),
    .Y(_0910_),
    .D(_0909_));
 sg13g2_nand3_1 _2701_ (.B(net1229),
    .C(_0910_),
    .A(\cpu.ctrl.o_ibus_adr[0] ),
    .Y(_0911_));
 sg13g2_a21o_1 _2702_ (.A2(_0910_),
    .A1(\cpu.ctrl.o_ibus_adr[0] ),
    .B1(\cpu.ctrl.pc_plus_offset_cy_r ),
    .X(_0912_));
 sg13g2_and2_1 _2703_ (.A(_0911_),
    .B(_0912_),
    .X(_0913_));
 sg13g2_nor2b_1 _2704_ (.A(net569),
    .B_N(net572),
    .Y(_0914_));
 sg13g2_and2_1 _2705_ (.A(net574),
    .B(_0914_),
    .X(_0915_));
 sg13g2_nand2_1 _2706_ (.Y(_0916_),
    .A(net574),
    .B(_0914_));
 sg13g2_a21oi_1 _2707_ (.A1(\cpu.state.o_cnt[2] ),
    .A2(\cpu.mem_bytecnt[0] ),
    .Y(_0917_),
    .B1(\cpu.mem_bytecnt[1] ));
 sg13g2_nand2b_2 _2708_ (.Y(_0918_),
    .B(net572),
    .A_N(net577));
 sg13g2_o21ai_1 _2709_ (.B1(\cpu.state.init_done ),
    .Y(_0919_),
    .A1(net576),
    .A2(\cpu.bufreg2.dat[5] ));
 sg13g2_nor3_1 _2710_ (.A(\cpu.state.stage_two_req ),
    .B(_0918_),
    .C(_0919_),
    .Y(_0920_));
 sg13g2_a21oi_1 _2711_ (.A1(_0090_),
    .A2(_0577_),
    .Y(_0921_),
    .B1(net549));
 sg13g2_a21oi_1 _2712_ (.A1(_0899_),
    .A2(_0921_),
    .Y(_0922_),
    .B1(_0920_));
 sg13g2_nor3_1 _2713_ (.A(_0890_),
    .B(_0916_),
    .C(_0917_),
    .Y(_0923_));
 sg13g2_nor3_1 _2714_ (.A(_0582_),
    .B(_0915_),
    .C(net546),
    .Y(_0924_));
 sg13g2_o21ai_1 _2715_ (.B1(_0913_),
    .Y(_0925_),
    .A1(_0923_),
    .A2(_0924_));
 sg13g2_a21oi_1 _2716_ (.A1(net1230),
    .A2(_0925_),
    .Y(_0016_),
    .B1(_0901_));
 sg13g2_nand2b_1 _2717_ (.Y(_0926_),
    .B(net575),
    .A_N(\cpu.decode.opcode[1] ));
 sg13g2_a21oi_1 _2718_ (.A1(net569),
    .A2(_0926_),
    .Y(_0927_),
    .B1(_0865_));
 sg13g2_nand2_1 _2719_ (.Y(_0928_),
    .A(net978),
    .B(_0927_));
 sg13g2_nand2_1 _2720_ (.Y(_0929_),
    .A(\cpu.state.cnt_r[0] ),
    .B(_0903_));
 sg13g2_nor2b_1 _2721_ (.A(_0883_),
    .B_N(_0908_),
    .Y(_0930_));
 sg13g2_nor3_1 _2722_ (.A(_0090_),
    .B(_0929_),
    .C(_0930_),
    .Y(_0931_));
 sg13g2_or3_1 _2723_ (.A(net572),
    .B(_0890_),
    .C(_0931_),
    .X(_0932_));
 sg13g2_xnor2_1 _2724_ (.Y(_0933_),
    .A(net978),
    .B(_0927_));
 sg13g2_or2_1 _2725_ (.X(_0934_),
    .B(_0933_),
    .A(_0932_));
 sg13g2_a21oi_1 _2726_ (.A1(_0928_),
    .A2(_0934_),
    .Y(_0014_),
    .B1(net545));
 sg13g2_nand2_2 _2727_ (.Y(_0935_),
    .A(net1278),
    .B(net532));
 sg13g2_nor2_1 _2728_ (.A(_0808_),
    .B(_0935_),
    .Y(_0000_));
 sg13g2_and2_1 _2729_ (.A(\dut.xfer.obuffer[7] ),
    .B(_0815_),
    .X(\dut.flash_io0_do ));
 sg13g2_and2_1 _2730_ (.A(\rf_shift_reg.cnt[2] ),
    .B(net826),
    .X(_0936_));
 sg13g2_nand4_1 _2731_ (.B(\rf_shift_reg.cnt[3] ),
    .C(\rf_shift_reg.cnt[0] ),
    .A(net1138),
    .Y(_0937_),
    .D(_0936_));
 sg13g2_a21oi_1 _2732_ (.A1(\rf_shift_reg.rd_active ),
    .A2(_0937_),
    .Y(_0938_),
    .B1(net1140));
 sg13g2_nor2_1 _2733_ (.A(_0465_),
    .B(net1141),
    .Y(_0094_));
 sg13g2_nand2_2 _2734_ (.Y(_0939_),
    .A(_0618_),
    .B(_0711_));
 sg13g2_inv_1 _2735_ (.Y(_0095_),
    .A(_0939_));
 sg13g2_nor2_1 _2736_ (.A(\cpu.immdec.imm11_7[0] ),
    .B(\cpu.immdec.imm11_7[4] ),
    .Y(_0940_));
 sg13g2_nor3_1 _2737_ (.A(\cpu.immdec.imm11_7[0] ),
    .B(\cpu.immdec.imm11_7[1] ),
    .C(\cpu.immdec.imm11_7[4] ),
    .Y(_0941_));
 sg13g2_nor2_2 _2738_ (.A(net1072),
    .B(\cpu.immdec.imm11_7[2] ),
    .Y(_0942_));
 sg13g2_and2_1 _2739_ (.A(net569),
    .B(net574),
    .X(_0943_));
 sg13g2_a221oi_1 _2740_ (.B2(_0563_),
    .C1(net573),
    .B1(_0091_),
    .A1(net570),
    .Y(_0944_),
    .A2(net574));
 sg13g2_a21oi_1 _2741_ (.A1(_0941_),
    .A2(_0942_),
    .Y(_0945_),
    .B1(_0944_));
 sg13g2_nor2b_2 _2742_ (.A(_0901_),
    .B_N(_0945_),
    .Y(_0946_));
 sg13g2_nor2_1 _2743_ (.A(\rf_shift_reg.rd_active ),
    .B(_0946_),
    .Y(_0947_));
 sg13g2_mux2_1 _2744_ (.A0(net646),
    .A1(\rf_shift_reg.rdata[1] ),
    .S(net517),
    .X(_0096_));
 sg13g2_mux2_1 _2745_ (.A0(net1028),
    .A1(net646),
    .S(net518),
    .X(_0097_));
 sg13g2_mux2_1 _2746_ (.A0(\rf_shift_reg.x[1][3] ),
    .A1(net1028),
    .S(net518),
    .X(_0098_));
 sg13g2_mux2_1 _2747_ (.A0(net640),
    .A1(\rf_shift_reg.x[1][3] ),
    .S(net518),
    .X(_0099_));
 sg13g2_mux2_1 _2748_ (.A0(net1077),
    .A1(net640),
    .S(net518),
    .X(_0100_));
 sg13g2_mux2_1 _2749_ (.A0(net925),
    .A1(\rf_shift_reg.x[1][5] ),
    .S(net518),
    .X(_0101_));
 sg13g2_mux2_1 _2750_ (.A0(net886),
    .A1(\rf_shift_reg.x[1][6] ),
    .S(net518),
    .X(_0102_));
 sg13g2_mux2_1 _2751_ (.A0(net1151),
    .A1(net886),
    .S(net515),
    .X(_0103_));
 sg13g2_mux2_1 _2752_ (.A0(net1013),
    .A1(\rf_shift_reg.x[1][8] ),
    .S(net515),
    .X(_0104_));
 sg13g2_mux2_1 _2753_ (.A0(net1063),
    .A1(net1013),
    .S(net515),
    .X(_0105_));
 sg13g2_mux2_1 _2754_ (.A0(net914),
    .A1(\rf_shift_reg.x[1][10] ),
    .S(net515),
    .X(_0106_));
 sg13g2_mux2_1 _2755_ (.A0(net1121),
    .A1(net914),
    .S(net515),
    .X(_0107_));
 sg13g2_mux2_1 _2756_ (.A0(net1064),
    .A1(\rf_shift_reg.x[1][12] ),
    .S(net507),
    .X(_0108_));
 sg13g2_mux2_1 _2757_ (.A0(net867),
    .A1(\rf_shift_reg.x[1][13] ),
    .S(net507),
    .X(_0109_));
 sg13g2_mux2_1 _2758_ (.A0(net1086),
    .A1(net867),
    .S(net507),
    .X(_0110_));
 sg13g2_mux2_1 _2759_ (.A0(net949),
    .A1(\rf_shift_reg.x[1][15] ),
    .S(net507),
    .X(_0111_));
 sg13g2_mux2_1 _2760_ (.A0(net1035),
    .A1(net949),
    .S(net507),
    .X(_0112_));
 sg13g2_mux2_1 _2761_ (.A0(net957),
    .A1(\rf_shift_reg.x[1][17] ),
    .S(net507),
    .X(_0113_));
 sg13g2_mux2_1 _2762_ (.A0(net975),
    .A1(net957),
    .S(net507),
    .X(_0114_));
 sg13g2_mux2_1 _2763_ (.A0(net1004),
    .A1(net975),
    .S(net507),
    .X(_0115_));
 sg13g2_mux2_1 _2764_ (.A0(net1123),
    .A1(net1004),
    .S(net508),
    .X(_0116_));
 sg13g2_mux2_1 _2765_ (.A0(net910),
    .A1(\rf_shift_reg.x[1][21] ),
    .S(net515),
    .X(_0117_));
 sg13g2_mux2_1 _2766_ (.A0(net792),
    .A1(\rf_shift_reg.x[1][22] ),
    .S(net515),
    .X(_0118_));
 sg13g2_mux2_1 _2767_ (.A0(net1003),
    .A1(net792),
    .S(net515),
    .X(_0119_));
 sg13g2_mux2_1 _2768_ (.A0(net904),
    .A1(\rf_shift_reg.x[1][24] ),
    .S(net516),
    .X(_0120_));
 sg13g2_mux2_1 _2769_ (.A0(net1106),
    .A1(net904),
    .S(net516),
    .X(_0121_));
 sg13g2_mux2_1 _2770_ (.A0(net916),
    .A1(\rf_shift_reg.x[1][26] ),
    .S(net517),
    .X(_0122_));
 sg13g2_mux2_1 _2771_ (.A0(net1124),
    .A1(net916),
    .S(net517),
    .X(_0123_));
 sg13g2_mux2_1 _2772_ (.A0(net642),
    .A1(\rf_shift_reg.x[1][28] ),
    .S(net517),
    .X(_0124_));
 sg13g2_mux2_1 _2773_ (.A0(net962),
    .A1(net642),
    .S(net517),
    .X(_0125_));
 sg13g2_mux2_1 _2774_ (.A0(net852),
    .A1(\rf_shift_reg.x[1][30] ),
    .S(net513),
    .X(_0126_));
 sg13g2_o21ai_1 _2775_ (.B1(_0867_),
    .Y(_0948_),
    .A1(_0893_),
    .A2(_0894_));
 sg13g2_nand2b_1 _2776_ (.Y(_0949_),
    .B(_0948_),
    .A_N(_0895_));
 sg13g2_nand2_1 _2777_ (.Y(_0950_),
    .A(_0017_),
    .B(_0855_));
 sg13g2_nor3_1 _2778_ (.A(_0865_),
    .B(_0875_),
    .C(_0891_),
    .Y(_0951_));
 sg13g2_o21ai_1 _2779_ (.B1(_0865_),
    .Y(_0952_),
    .A1(_0875_),
    .A2(_0891_));
 sg13g2_nor2b_1 _2780_ (.A(_0951_),
    .B_N(_0952_),
    .Y(_0953_));
 sg13g2_nor2b_1 _2781_ (.A(\cpu.bne_or_bge ),
    .B_N(net576),
    .Y(_0954_));
 sg13g2_nor2b_1 _2782_ (.A(net576),
    .B_N(net577),
    .Y(_0955_));
 sg13g2_nand4_1 _2783_ (.B(\cpu.alu.cmp_r ),
    .C(_0903_),
    .A(\cpu.state.cnt_r[0] ),
    .Y(_0956_),
    .D(_0955_));
 sg13g2_o21ai_1 _2784_ (.B1(_0956_),
    .Y(_0957_),
    .A1(_0582_),
    .A2(net545));
 sg13g2_a221oi_1 _2785_ (.B2(_0954_),
    .C1(_0957_),
    .B1(_0953_),
    .A1(_0897_),
    .Y(_0958_),
    .A2(_0951_));
 sg13g2_o21ai_1 _2786_ (.B1(_0958_),
    .Y(_0959_),
    .A1(_0949_),
    .A2(_0950_));
 sg13g2_nor2b_1 _2787_ (.A(net574),
    .B_N(_0914_),
    .Y(_0960_));
 sg13g2_or3_1 _2788_ (.A(_0913_),
    .B(_0923_),
    .C(_0924_),
    .X(_0961_));
 sg13g2_nand3_1 _2789_ (.B(_0929_),
    .C(_0961_),
    .A(_0925_),
    .Y(_0962_));
 sg13g2_mux4_1 _2790_ (.S0(_0582_),
    .A0(\cpu.bufreg2.dat[24] ),
    .A1(\cpu.bufreg2.dat[16] ),
    .A2(\cpu.bufreg2.dat[8] ),
    .A3(_0593_),
    .S1(_0591_),
    .X(_0963_));
 sg13g2_a21oi_1 _2791_ (.A1(\cpu.mem_bytecnt[0] ),
    .A2(_0575_),
    .Y(_0964_),
    .B1(\cpu.mem_bytecnt[1] ));
 sg13g2_nor2_1 _2792_ (.A(\cpu.decode.co_mem_word ),
    .B(_0964_),
    .Y(_0965_));
 sg13g2_o21ai_1 _2793_ (.B1(_0963_),
    .Y(_0966_),
    .A1(net577),
    .A2(_0964_));
 sg13g2_nand2_1 _2794_ (.Y(_0967_),
    .A(net799),
    .B(_0965_));
 sg13g2_nand2_1 _2795_ (.Y(_0413_),
    .A(_0966_),
    .B(net800));
 sg13g2_o21ai_1 _2796_ (.B1(_0966_),
    .Y(_0968_),
    .A1(\cpu.csr_d_sel ),
    .A2(_0967_));
 sg13g2_a21o_1 _2797_ (.A2(_0903_),
    .A1(\cpu.state.cnt_r[2] ),
    .B1(_0904_),
    .X(_0969_));
 sg13g2_and2_1 _2798_ (.A(_0905_),
    .B(_0969_),
    .X(_0970_));
 sg13g2_a22oi_1 _2799_ (.Y(_0971_),
    .B1(_0970_),
    .B2(_0943_),
    .A2(_0968_),
    .A1(_0885_));
 sg13g2_o21ai_1 _2800_ (.B1(_0971_),
    .Y(_0972_),
    .A1(_0916_),
    .A2(_0962_));
 sg13g2_a21o_2 _2801_ (.A2(_0960_),
    .A1(_0959_),
    .B1(_0972_),
    .X(_0973_));
 sg13g2_inv_1 _2802_ (.Y(_0974_),
    .A(_0973_));
 sg13g2_nor2b_1 _2803_ (.A(\cpu.immdec.imm11_7[4] ),
    .B_N(\cpu.immdec.imm11_7[0] ),
    .Y(_0975_));
 sg13g2_nor2b_1 _2804_ (.A(\cpu.immdec.imm11_7[1] ),
    .B_N(_0975_),
    .Y(_0976_));
 sg13g2_nand3_1 _2805_ (.B(_0946_),
    .C(_0976_),
    .A(net1073),
    .Y(_0977_));
 sg13g2_nor2b_1 _2806_ (.A(net514),
    .B_N(\rf_shift_reg.rdata[1] ),
    .Y(_0978_));
 sg13g2_a22oi_1 _2807_ (.Y(_0979_),
    .B1(_0977_),
    .B2(_0978_),
    .A2(net512),
    .A1(net852));
 sg13g2_o21ai_1 _2808_ (.B1(_0979_),
    .Y(_0127_),
    .A1(_0974_),
    .A2(net1074));
 sg13g2_o21ai_1 _2809_ (.B1(net582),
    .Y(_0980_),
    .A1(\rf_shift_reg.rd_active ),
    .A2(\rf_shift_reg.cnt[0] ));
 sg13g2_a21oi_1 _2810_ (.A1(\rf_shift_reg.rd_active ),
    .A2(_0557_),
    .Y(_0128_),
    .B1(_0980_));
 sg13g2_a21oi_1 _2811_ (.A1(\rf_shift_reg.rd_active ),
    .A2(\rf_shift_reg.cnt[0] ),
    .Y(_0981_),
    .B1(net826));
 sg13g2_nand3_1 _2812_ (.B(net826),
    .C(\rf_shift_reg.cnt[0] ),
    .A(\rf_shift_reg.rd_active ),
    .Y(_0982_));
 sg13g2_nand2_1 _2813_ (.Y(_0983_),
    .A(net582),
    .B(_0982_));
 sg13g2_nor2_1 _2814_ (.A(net827),
    .B(_0983_),
    .Y(_0129_));
 sg13g2_nand2b_1 _2815_ (.Y(_0984_),
    .B(_0982_),
    .A_N(net1308));
 sg13g2_nand3_1 _2816_ (.B(\rf_shift_reg.cnt[0] ),
    .C(_0936_),
    .A(\rf_shift_reg.rd_active ),
    .Y(_0985_));
 sg13g2_and3_1 _2817_ (.X(_0130_),
    .A(net582),
    .B(net1309),
    .C(_0985_));
 sg13g2_nand2b_1 _2818_ (.Y(_0986_),
    .B(_0985_),
    .A_N(net1321));
 sg13g2_nand4_1 _2819_ (.B(net1321),
    .C(\rf_shift_reg.cnt[0] ),
    .A(\rf_shift_reg.rd_active ),
    .Y(_0987_),
    .D(_0936_));
 sg13g2_and3_1 _2820_ (.X(_0131_),
    .A(net583),
    .B(net1322),
    .C(_0987_));
 sg13g2_o21ai_1 _2821_ (.B1(net582),
    .Y(_0988_),
    .A1(_0556_),
    .A2(_0987_));
 sg13g2_a21oi_1 _2822_ (.A1(_0556_),
    .A2(_0987_),
    .Y(_0132_),
    .B1(_0988_));
 sg13g2_mux2_1 _2823_ (.A0(net663),
    .A1(\rf_shift_reg.rdata[2] ),
    .S(net510),
    .X(_0133_));
 sg13g2_mux2_1 _2824_ (.A0(net1169),
    .A1(net663),
    .S(net510),
    .X(_0134_));
 sg13g2_mux2_1 _2825_ (.A0(net1007),
    .A1(\rf_shift_reg.x[2][2] ),
    .S(net500),
    .X(_0135_));
 sg13g2_mux2_1 _2826_ (.A0(net817),
    .A1(\rf_shift_reg.x[2][3] ),
    .S(net497),
    .X(_0136_));
 sg13g2_mux2_1 _2827_ (.A0(net1181),
    .A1(net817),
    .S(net498),
    .X(_0137_));
 sg13g2_mux2_1 _2828_ (.A0(net1018),
    .A1(\rf_shift_reg.x[2][5] ),
    .S(net498),
    .X(_0138_));
 sg13g2_mux2_1 _2829_ (.A0(net1087),
    .A1(net1018),
    .S(net498),
    .X(_0139_));
 sg13g2_mux2_1 _2830_ (.A0(net1157),
    .A1(net1087),
    .S(net495),
    .X(_0140_));
 sg13g2_mux2_1 _2831_ (.A0(net933),
    .A1(\rf_shift_reg.x[2][8] ),
    .S(net495),
    .X(_0141_));
 sg13g2_mux2_1 _2832_ (.A0(net1127),
    .A1(net933),
    .S(net495),
    .X(_0142_));
 sg13g2_mux2_1 _2833_ (.A0(net1194),
    .A1(net1127),
    .S(net495),
    .X(_0143_));
 sg13g2_mux2_1 _2834_ (.A0(net981),
    .A1(\rf_shift_reg.x[2][11] ),
    .S(net495),
    .X(_0144_));
 sg13g2_mux2_1 _2835_ (.A0(net999),
    .A1(net981),
    .S(net495),
    .X(_0145_));
 sg13g2_mux2_1 _2836_ (.A0(net1095),
    .A1(net999),
    .S(net495),
    .X(_0146_));
 sg13g2_mux2_1 _2837_ (.A0(net979),
    .A1(\rf_shift_reg.x[2][14] ),
    .S(net495),
    .X(_0147_));
 sg13g2_mux2_1 _2838_ (.A0(net863),
    .A1(\rf_shift_reg.x[2][15] ),
    .S(net494),
    .X(_0148_));
 sg13g2_mux2_1 _2839_ (.A0(net959),
    .A1(net863),
    .S(net494),
    .X(_0149_));
 sg13g2_mux2_1 _2840_ (.A0(net974),
    .A1(net959),
    .S(net494),
    .X(_0150_));
 sg13g2_mux2_1 _2841_ (.A0(net994),
    .A1(net974),
    .S(net491),
    .X(_0151_));
 sg13g2_mux2_1 _2842_ (.A0(net912),
    .A1(\rf_shift_reg.x[2][19] ),
    .S(net491),
    .X(_0152_));
 sg13g2_mux2_1 _2843_ (.A0(net1093),
    .A1(net912),
    .S(net491),
    .X(_0153_));
 sg13g2_mux2_1 _2844_ (.A0(net1160),
    .A1(net1093),
    .S(net491),
    .X(_0154_));
 sg13g2_mux2_1 _2845_ (.A0(net890),
    .A1(\rf_shift_reg.x[2][22] ),
    .S(net497),
    .X(_0155_));
 sg13g2_mux2_1 _2846_ (.A0(net893),
    .A1(net890),
    .S(net497),
    .X(_0156_));
 sg13g2_mux2_1 _2847_ (.A0(net1108),
    .A1(net893),
    .S(net497),
    .X(_0157_));
 sg13g2_mux2_1 _2848_ (.A0(net1024),
    .A1(\rf_shift_reg.x[2][25] ),
    .S(net497),
    .X(_0158_));
 sg13g2_mux2_1 _2849_ (.A0(net1020),
    .A1(\rf_shift_reg.x[2][26] ),
    .S(net497),
    .X(_0159_));
 sg13g2_mux2_1 _2850_ (.A0(net1080),
    .A1(net1020),
    .S(net500),
    .X(_0160_));
 sg13g2_mux2_1 _2851_ (.A0(net830),
    .A1(\rf_shift_reg.x[2][28] ),
    .S(net500),
    .X(_0161_));
 sg13g2_mux2_1 _2852_ (.A0(net682),
    .A1(net830),
    .S(net500),
    .X(_0162_));
 sg13g2_nand2_1 _2853_ (.Y(_0989_),
    .A(net682),
    .B(net501));
 sg13g2_o21ai_1 _2854_ (.B1(_0989_),
    .Y(_0163_),
    .A1(_0615_),
    .A2(net502));
 sg13g2_nand4_1 _2855_ (.B(_0940_),
    .C(_0942_),
    .A(net1185),
    .Y(_0990_),
    .D(_0946_));
 sg13g2_nand2b_1 _2856_ (.Y(_0991_),
    .B(_0973_),
    .A_N(_0990_));
 sg13g2_a21oi_1 _2857_ (.A1(\rf_shift_reg.rdata[2] ),
    .A2(_0990_),
    .Y(_0992_),
    .B1(net513));
 sg13g2_a22oi_1 _2858_ (.Y(_0164_),
    .B1(_0991_),
    .B2(_0992_),
    .A2(net513),
    .A1(_0615_));
 sg13g2_nor2_1 _2859_ (.A(net644),
    .B(net512),
    .Y(_0993_));
 sg13g2_a21oi_1 _2860_ (.A1(_0585_),
    .A2(net512),
    .Y(_0165_),
    .B1(_0993_));
 sg13g2_mux2_1 _2861_ (.A0(net1031),
    .A1(net644),
    .S(net512),
    .X(_0166_));
 sg13g2_mux2_1 _2862_ (.A0(net1112),
    .A1(net1031),
    .S(net512),
    .X(_0167_));
 sg13g2_mux2_1 _2863_ (.A0(net1122),
    .A1(net1112),
    .S(net511),
    .X(_0168_));
 sg13g2_mux2_1 _2864_ (.A0(net1088),
    .A1(\rf_shift_reg.x[3][4] ),
    .S(net511),
    .X(_0169_));
 sg13g2_mux2_1 _2865_ (.A0(net953),
    .A1(\rf_shift_reg.x[3][5] ),
    .S(net511),
    .X(_0170_));
 sg13g2_mux2_1 _2866_ (.A0(net1039),
    .A1(net953),
    .S(net511),
    .X(_0171_));
 sg13g2_mux2_1 _2867_ (.A0(net1045),
    .A1(net1039),
    .S(net505),
    .X(_0172_));
 sg13g2_mux2_1 _2868_ (.A0(net992),
    .A1(\rf_shift_reg.x[3][8] ),
    .S(net505),
    .X(_0173_));
 sg13g2_mux2_1 _2869_ (.A0(net1038),
    .A1(net992),
    .S(net505),
    .X(_0174_));
 sg13g2_mux2_1 _2870_ (.A0(net968),
    .A1(\rf_shift_reg.x[3][10] ),
    .S(net506),
    .X(_0175_));
 sg13g2_mux2_1 _2871_ (.A0(net1105),
    .A1(net968),
    .S(net506),
    .X(_0176_));
 sg13g2_mux2_1 _2872_ (.A0(net1090),
    .A1(\rf_shift_reg.x[3][12] ),
    .S(net504),
    .X(_0177_));
 sg13g2_mux2_1 _2873_ (.A0(net882),
    .A1(\rf_shift_reg.x[3][13] ),
    .S(net503),
    .X(_0178_));
 sg13g2_mux2_1 _2874_ (.A0(net1115),
    .A1(net882),
    .S(net504),
    .X(_0179_));
 sg13g2_mux2_1 _2875_ (.A0(net1000),
    .A1(\rf_shift_reg.x[3][15] ),
    .S(net504),
    .X(_0180_));
 sg13g2_mux2_1 _2876_ (.A0(net1027),
    .A1(net1000),
    .S(net503),
    .X(_0181_));
 sg13g2_mux2_1 _2877_ (.A0(net738),
    .A1(\rf_shift_reg.x[3][17] ),
    .S(net503),
    .X(_0182_));
 sg13g2_mux2_1 _2878_ (.A0(net1071),
    .A1(net738),
    .S(net503),
    .X(_0183_));
 sg13g2_mux2_1 _2879_ (.A0(net726),
    .A1(\rf_shift_reg.x[3][19] ),
    .S(net503),
    .X(_0184_));
 sg13g2_mux2_1 _2880_ (.A0(net1113),
    .A1(net726),
    .S(net505),
    .X(_0185_));
 sg13g2_mux2_1 _2881_ (.A0(net802),
    .A1(\rf_shift_reg.x[3][21] ),
    .S(net505),
    .X(_0186_));
 sg13g2_mux2_1 _2882_ (.A0(net973),
    .A1(net802),
    .S(net505),
    .X(_0187_));
 sg13g2_mux2_1 _2883_ (.A0(net1136),
    .A1(net973),
    .S(net505),
    .X(_0188_));
 sg13g2_mux2_1 _2884_ (.A0(net1150),
    .A1(net1136),
    .S(net505),
    .X(_0189_));
 sg13g2_mux2_1 _2885_ (.A0(net790),
    .A1(\rf_shift_reg.x[3][25] ),
    .S(net510),
    .X(_0190_));
 sg13g2_mux2_1 _2886_ (.A0(net1050),
    .A1(net790),
    .S(net510),
    .X(_0191_));
 sg13g2_mux2_1 _2887_ (.A0(net1079),
    .A1(net1050),
    .S(net510),
    .X(_0192_));
 sg13g2_mux2_1 _2888_ (.A0(net703),
    .A1(\rf_shift_reg.x[3][28] ),
    .S(net511),
    .X(_0193_));
 sg13g2_mux2_1 _2889_ (.A0(net1162),
    .A1(net703),
    .S(net512),
    .X(_0194_));
 sg13g2_mux2_1 _2890_ (.A0(net678),
    .A1(\rf_shift_reg.x[3][30] ),
    .S(net512),
    .X(_0195_));
 sg13g2_nand4_1 _2891_ (.B(net1073),
    .C(_0946_),
    .A(net1185),
    .Y(_0994_),
    .D(_0975_));
 sg13g2_nor2_1 _2892_ (.A(_0585_),
    .B(net512),
    .Y(_0995_));
 sg13g2_a22oi_1 _2893_ (.Y(_0996_),
    .B1(_0994_),
    .B2(_0995_),
    .A2(net513),
    .A1(net678));
 sg13g2_o21ai_1 _2894_ (.B1(_0996_),
    .Y(_0196_),
    .A1(_0974_),
    .A2(net1186));
 sg13g2_nor2_1 _2895_ (.A(net652),
    .B(net501),
    .Y(_0997_));
 sg13g2_a21oi_1 _2896_ (.A1(_0586_),
    .A2(net513),
    .Y(_0197_),
    .B1(_0997_));
 sg13g2_mux2_1 _2897_ (.A0(net946),
    .A1(net652),
    .S(net501),
    .X(_0198_));
 sg13g2_mux2_1 _2898_ (.A0(net1133),
    .A1(net946),
    .S(net501),
    .X(_0199_));
 sg13g2_mux2_1 _2899_ (.A0(net1146),
    .A1(net1133),
    .S(net500),
    .X(_0200_));
 sg13g2_mux2_1 _2900_ (.A0(net1066),
    .A1(\rf_shift_reg.x[4][4] ),
    .S(net500),
    .X(_0201_));
 sg13g2_mux2_1 _2901_ (.A0(net1040),
    .A1(\rf_shift_reg.x[4][5] ),
    .S(net500),
    .X(_0202_));
 sg13g2_mux2_1 _2902_ (.A0(net935),
    .A1(\rf_shift_reg.x[4][6] ),
    .S(net502),
    .X(_0203_));
 sg13g2_mux2_1 _2903_ (.A0(net859),
    .A1(\rf_shift_reg.x[4][7] ),
    .S(net493),
    .X(_0204_));
 sg13g2_mux2_1 _2904_ (.A0(net892),
    .A1(net859),
    .S(net493),
    .X(_0205_));
 sg13g2_mux2_1 _2905_ (.A0(net1030),
    .A1(net892),
    .S(net493),
    .X(_0206_));
 sg13g2_mux2_1 _2906_ (.A0(net1107),
    .A1(net1030),
    .S(net493),
    .X(_0207_));
 sg13g2_mux2_1 _2907_ (.A0(net955),
    .A1(\rf_shift_reg.x[4][11] ),
    .S(net493),
    .X(_0208_));
 sg13g2_mux2_1 _2908_ (.A0(net1002),
    .A1(net955),
    .S(net493),
    .X(_0209_));
 sg13g2_mux2_1 _2909_ (.A0(net1165),
    .A1(net1002),
    .S(net492),
    .X(_0210_));
 sg13g2_mux2_1 _2910_ (.A0(net985),
    .A1(\rf_shift_reg.x[4][14] ),
    .S(net491),
    .X(_0211_));
 sg13g2_mux2_1 _2911_ (.A0(net964),
    .A1(\rf_shift_reg.x[4][15] ),
    .S(net491),
    .X(_0212_));
 sg13g2_mux2_1 _2912_ (.A0(net1109),
    .A1(net964),
    .S(net491),
    .X(_0213_));
 sg13g2_mux2_1 _2913_ (.A0(net865),
    .A1(\rf_shift_reg.x[4][17] ),
    .S(net491),
    .X(_0214_));
 sg13g2_mux2_1 _2914_ (.A0(net1094),
    .A1(net865),
    .S(net492),
    .X(_0215_));
 sg13g2_mux2_1 _2915_ (.A0(net676),
    .A1(\rf_shift_reg.x[4][19] ),
    .S(net492),
    .X(_0216_));
 sg13g2_mux2_1 _2916_ (.A0(net1076),
    .A1(net676),
    .S(net492),
    .X(_0217_));
 sg13g2_mux2_1 _2917_ (.A0(net750),
    .A1(\rf_shift_reg.x[4][21] ),
    .S(net492),
    .X(_0218_));
 sg13g2_mux2_1 _2918_ (.A0(net1180),
    .A1(net750),
    .S(net492),
    .X(_0219_));
 sg13g2_mux2_1 _2919_ (.A0(net832),
    .A1(\rf_shift_reg.x[4][23] ),
    .S(net492),
    .X(_0220_));
 sg13g2_mux2_1 _2920_ (.A0(net1166),
    .A1(net832),
    .S(net492),
    .X(_0221_));
 sg13g2_mux2_1 _2921_ (.A0(net997),
    .A1(\rf_shift_reg.x[4][25] ),
    .S(net502),
    .X(_0222_));
 sg13g2_mux2_1 _2922_ (.A0(net902),
    .A1(\rf_shift_reg.x[4][26] ),
    .S(net502),
    .X(_0223_));
 sg13g2_mux2_1 _2923_ (.A0(net1092),
    .A1(net902),
    .S(net502),
    .X(_0224_));
 sg13g2_mux2_1 _2924_ (.A0(net1154),
    .A1(net1092),
    .S(net502),
    .X(_0225_));
 sg13g2_mux2_1 _2925_ (.A0(net960),
    .A1(\rf_shift_reg.x[4][29] ),
    .S(net500),
    .X(_0226_));
 sg13g2_mux2_1 _2926_ (.A0(net730),
    .A1(net960),
    .S(net501),
    .X(_0227_));
 sg13g2_nand2_1 _2927_ (.Y(_0998_),
    .A(net730),
    .B(net501));
 sg13g2_nor2b_1 _2928_ (.A(\cpu.immdec.imm11_7[3] ),
    .B_N(\cpu.immdec.imm11_7[2] ),
    .Y(_0999_));
 sg13g2_nand3_1 _2929_ (.B(_0946_),
    .C(_0999_),
    .A(_0941_),
    .Y(_1000_));
 sg13g2_a21oi_1 _2930_ (.A1(_0586_),
    .A2(_1000_),
    .Y(_1001_),
    .B1(net501));
 sg13g2_o21ai_1 _2931_ (.B1(_1001_),
    .Y(_1002_),
    .A1(_0973_),
    .A2(_1000_));
 sg13g2_nand2_1 _2932_ (.Y(_0228_),
    .A(_0998_),
    .B(_1002_));
 sg13g2_nor2_1 _2933_ (.A(net667),
    .B(net517),
    .Y(_1003_));
 sg13g2_a21oi_1 _2934_ (.A1(_0587_),
    .A2(net517),
    .Y(_0229_),
    .B1(_1003_));
 sg13g2_mux2_1 _2935_ (.A0(net963),
    .A1(net667),
    .S(net517),
    .X(_0230_));
 sg13g2_mux2_1 _2936_ (.A0(net944),
    .A1(\rf_shift_reg.x[5][2] ),
    .S(net516),
    .X(_0231_));
 sg13g2_mux2_1 _2937_ (.A0(net923),
    .A1(\rf_shift_reg.x[5][3] ),
    .S(net516),
    .X(_0232_));
 sg13g2_mux2_1 _2938_ (.A0(net1023),
    .A1(net923),
    .S(net516),
    .X(_0233_));
 sg13g2_mux2_1 _2939_ (.A0(net1145),
    .A1(net1023),
    .S(net508),
    .X(_0234_));
 sg13g2_mux2_1 _2940_ (.A0(net966),
    .A1(\rf_shift_reg.x[5][6] ),
    .S(net508),
    .X(_0235_));
 sg13g2_mux2_1 _2941_ (.A0(net908),
    .A1(\rf_shift_reg.x[5][7] ),
    .S(net508),
    .X(_0236_));
 sg13g2_mux2_1 _2942_ (.A0(net847),
    .A1(\rf_shift_reg.x[5][8] ),
    .S(net509),
    .X(_0237_));
 sg13g2_mux2_1 _2943_ (.A0(net1132),
    .A1(net847),
    .S(net509),
    .X(_0238_));
 sg13g2_mux2_1 _2944_ (.A0(net1147),
    .A1(net1132),
    .S(net509),
    .X(_0239_));
 sg13g2_mux2_1 _2945_ (.A0(net856),
    .A1(\rf_shift_reg.x[5][11] ),
    .S(net509),
    .X(_0240_));
 sg13g2_mux2_1 _2946_ (.A0(net1044),
    .A1(net856),
    .S(net509),
    .X(_0241_));
 sg13g2_mux2_1 _2947_ (.A0(net1142),
    .A1(net1044),
    .S(net509),
    .X(_0242_));
 sg13g2_mux2_1 _2948_ (.A0(net951),
    .A1(\rf_shift_reg.x[5][14] ),
    .S(net509),
    .X(_0243_));
 sg13g2_mux2_1 _2949_ (.A0(net1134),
    .A1(net951),
    .S(net504),
    .X(_0244_));
 sg13g2_mux2_1 _2950_ (.A0(net1053),
    .A1(\rf_shift_reg.x[5][16] ),
    .S(net504),
    .X(_0245_));
 sg13g2_mux2_1 _2951_ (.A0(net1036),
    .A1(\rf_shift_reg.x[5][17] ),
    .S(net504),
    .X(_0246_));
 sg13g2_mux2_1 _2952_ (.A0(net1005),
    .A1(\rf_shift_reg.x[5][18] ),
    .S(net503),
    .X(_0247_));
 sg13g2_mux2_1 _2953_ (.A0(net811),
    .A1(\rf_shift_reg.x[5][19] ),
    .S(net503),
    .X(_0248_));
 sg13g2_mux2_1 _2954_ (.A0(net991),
    .A1(net811),
    .S(net503),
    .X(_0249_));
 sg13g2_mux2_1 _2955_ (.A0(net896),
    .A1(\rf_shift_reg.x[5][21] ),
    .S(net496),
    .X(_0250_));
 sg13g2_mux2_1 _2956_ (.A0(net1068),
    .A1(net896),
    .S(net496),
    .X(_0251_));
 sg13g2_mux2_1 _2957_ (.A0(net942),
    .A1(\rf_shift_reg.x[5][23] ),
    .S(net496),
    .X(_0252_));
 sg13g2_mux2_1 _2958_ (.A0(net948),
    .A1(net942),
    .S(net496),
    .X(_0253_));
 sg13g2_mux2_1 _2959_ (.A0(net871),
    .A1(\rf_shift_reg.x[5][25] ),
    .S(net498),
    .X(_0254_));
 sg13g2_mux2_1 _2960_ (.A0(net970),
    .A1(net871),
    .S(net497),
    .X(_0255_));
 sg13g2_mux2_1 _2961_ (.A0(net1135),
    .A1(net970),
    .S(net497),
    .X(_0256_));
 sg13g2_mux2_1 _2962_ (.A0(net1171),
    .A1(net1135),
    .S(net510),
    .X(_0257_));
 sg13g2_mux2_1 _2963_ (.A0(net918),
    .A1(\rf_shift_reg.x[5][29] ),
    .S(net510),
    .X(_0258_));
 sg13g2_mux2_1 _2964_ (.A0(net669),
    .A1(net918),
    .S(net510),
    .X(_0259_));
 sg13g2_nand2_1 _2965_ (.Y(_1004_),
    .A(net669),
    .B(net513));
 sg13g2_nand3_1 _2966_ (.B(_0976_),
    .C(_0999_),
    .A(_0946_),
    .Y(_1005_));
 sg13g2_a21oi_1 _2967_ (.A1(_0587_),
    .A2(_1005_),
    .Y(_1006_),
    .B1(net513));
 sg13g2_o21ai_1 _2968_ (.B1(_1006_),
    .Y(_1007_),
    .A1(_0973_),
    .A2(_1005_));
 sg13g2_nand2_1 _2969_ (.Y(_0260_),
    .A(_1004_),
    .B(_1007_));
 sg13g2_and4_1 _2970_ (.A(net585),
    .B(_0564_),
    .C(net638),
    .D(_0623_),
    .X(_0261_));
 sg13g2_nor2_1 _2971_ (.A(_0809_),
    .B(_0816_),
    .Y(_1008_));
 sg13g2_a22oi_1 _2972_ (.Y(_1009_),
    .B1(_0822_),
    .B2(_1008_),
    .A2(_0816_),
    .A1(net778));
 sg13g2_nor3_1 _2973_ (.A(net744),
    .B(net537),
    .C(net779),
    .Y(_0262_));
 sg13g2_nor3_1 _2974_ (.A(_0548_),
    .B(_0810_),
    .C(_0816_),
    .Y(_1010_));
 sg13g2_xnor2_1 _2975_ (.Y(_1011_),
    .A(net746),
    .B(_1010_));
 sg13g2_nor3_1 _2976_ (.A(net744),
    .B(net537),
    .C(_1011_),
    .Y(_0263_));
 sg13g2_a22oi_1 _2977_ (.Y(_1012_),
    .B1(_0820_),
    .B2(_1008_),
    .A2(_0816_),
    .A1(net809));
 sg13g2_nor3_1 _2978_ (.A(net744),
    .B(net537),
    .C(net810),
    .Y(_0264_));
 sg13g2_and2_1 _2979_ (.A(net583),
    .B(net635),
    .X(_0265_));
 sg13g2_nand2_2 _2980_ (.Y(_1013_),
    .A(net571),
    .B(_0623_));
 sg13g2_o21ai_1 _2981_ (.B1(net586),
    .Y(_1014_),
    .A1(\cpu.bufreg2.dat[0] ),
    .A2(net540));
 sg13g2_a21oi_1 _2982_ (.A1(_0555_),
    .A2(_1013_),
    .Y(_0266_),
    .B1(_1014_));
 sg13g2_o21ai_1 _2983_ (.B1(net586),
    .Y(_1015_),
    .A1(\cpu.bufreg2.dat[1] ),
    .A2(net540));
 sg13g2_a21oi_1 _2984_ (.A1(_0554_),
    .A2(_1013_),
    .Y(_0267_),
    .B1(_1015_));
 sg13g2_o21ai_1 _2985_ (.B1(net586),
    .Y(_1016_),
    .A1(\cpu.bufreg2.dat[2] ),
    .A2(net540));
 sg13g2_a21oi_1 _2986_ (.A1(_0553_),
    .A2(net540),
    .Y(_0268_),
    .B1(_1016_));
 sg13g2_o21ai_1 _2987_ (.B1(net586),
    .Y(_1017_),
    .A1(\cpu.bufreg2.dat[3] ),
    .A2(net540));
 sg13g2_a21oi_1 _2988_ (.A1(_0552_),
    .A2(net540),
    .Y(_0269_),
    .B1(_1017_));
 sg13g2_o21ai_1 _2989_ (.B1(net586),
    .Y(_1018_),
    .A1(\cpu.bufreg2.dat[4] ),
    .A2(net540));
 sg13g2_a21oi_1 _2990_ (.A1(_0551_),
    .A2(net540),
    .Y(_0270_),
    .B1(_1018_));
 sg13g2_nor2b_2 _2991_ (.A(net550),
    .B_N(_0944_),
    .Y(_1019_));
 sg13g2_and2_1 _2992_ (.A(_0618_),
    .B(_0725_),
    .X(_1020_));
 sg13g2_inv_2 _2993_ (.Y(_1021_),
    .A(net487));
 sg13g2_nand3_1 _2994_ (.B(_1019_),
    .C(_1021_),
    .A(net1185),
    .Y(_1022_));
 sg13g2_nor2_2 _2995_ (.A(_1019_),
    .B(net486),
    .Y(_1023_));
 sg13g2_nand2_1 _2996_ (.Y(_1024_),
    .A(net1307),
    .B(_1023_));
 sg13g2_nand2_2 _2997_ (.Y(_1025_),
    .A(net1234),
    .B(net482));
 sg13g2_nand3_1 _2998_ (.B(_1024_),
    .C(_1025_),
    .A(_1022_),
    .Y(_0271_));
 sg13g2_and3_1 _2999_ (.X(_1026_),
    .A(net1288),
    .B(_1019_),
    .C(_1021_));
 sg13g2_a221oi_1 _3000_ (.B2(net1185),
    .C1(_1026_),
    .B1(_1023_),
    .A1(net1334),
    .Y(_1027_),
    .A2(net486));
 sg13g2_inv_1 _3001_ (.Y(_0272_),
    .A(_1027_));
 sg13g2_and3_1 _3002_ (.X(_1028_),
    .A(net1072),
    .B(_1019_),
    .C(_1021_));
 sg13g2_a221oi_1 _3003_ (.B2(net1288),
    .C1(_1028_),
    .B1(_1023_),
    .A1(net1057),
    .Y(_1029_),
    .A2(net488));
 sg13g2_inv_1 _3004_ (.Y(_0273_),
    .A(_1029_));
 sg13g2_and3_1 _3005_ (.X(_1030_),
    .A(net1276),
    .B(_1019_),
    .C(_1021_));
 sg13g2_a221oi_1 _3006_ (.B2(net1072),
    .C1(_1030_),
    .B1(_1023_),
    .A1(net851),
    .Y(_1031_),
    .A2(net486));
 sg13g2_inv_1 _3007_ (.Y(_0274_),
    .A(_1031_));
 sg13g2_nand2_1 _3008_ (.Y(_1032_),
    .A(net1252),
    .B(_0939_));
 sg13g2_a21oi_1 _3009_ (.A1(net789),
    .A2(_0095_),
    .Y(_1033_),
    .B1(_1023_));
 sg13g2_a22oi_1 _3010_ (.Y(_0275_),
    .B1(_1032_),
    .B2(_1033_),
    .A2(_1023_),
    .A1(_0579_));
 sg13g2_nor2_1 _3011_ (.A(_0465_),
    .B(_0901_),
    .Y(_1034_));
 sg13g2_and2_1 _3012_ (.A(net582),
    .B(_0901_),
    .X(_1035_));
 sg13g2_a22oi_1 _3013_ (.Y(_1036_),
    .B1(net524),
    .B2(net1251),
    .A2(net530),
    .A1(net752));
 sg13g2_inv_1 _3014_ (.Y(_0276_),
    .A(_1036_));
 sg13g2_a22oi_1 _3015_ (.Y(_1037_),
    .B1(net525),
    .B2(net752),
    .A2(net530),
    .A1(net661));
 sg13g2_inv_1 _3016_ (.Y(_0277_),
    .A(_1037_));
 sg13g2_a22oi_1 _3017_ (.Y(_1038_),
    .B1(net525),
    .B2(net661),
    .A2(net529),
    .A1(\cpu.ctrl.o_ibus_adr[3] ));
 sg13g2_inv_1 _3018_ (.Y(_0278_),
    .A(net662));
 sg13g2_a22oi_1 _3019_ (.Y(_1039_),
    .B1(net525),
    .B2(net735),
    .A2(net529),
    .A1(net656));
 sg13g2_inv_1 _3020_ (.Y(_0279_),
    .A(_1039_));
 sg13g2_a22oi_1 _3021_ (.Y(_1040_),
    .B1(net525),
    .B2(net656),
    .A2(net530),
    .A1(\cpu.ctrl.o_ibus_adr[5] ));
 sg13g2_inv_1 _3022_ (.Y(_0280_),
    .A(net657));
 sg13g2_a22oi_1 _3023_ (.Y(_1041_),
    .B1(net526),
    .B2(net724),
    .A2(net529),
    .A1(net684));
 sg13g2_inv_1 _3024_ (.Y(_0281_),
    .A(_1041_));
 sg13g2_a22oi_1 _3025_ (.Y(_1042_),
    .B1(net526),
    .B2(net684),
    .A2(net529),
    .A1(\cpu.ctrl.o_ibus_adr[7] ));
 sg13g2_inv_1 _3026_ (.Y(_0282_),
    .A(net685));
 sg13g2_a22oi_1 _3027_ (.Y(_1043_),
    .B1(net526),
    .B2(net686),
    .A2(net529),
    .A1(\cpu.ctrl.o_ibus_adr[8] ));
 sg13g2_inv_1 _3028_ (.Y(_0283_),
    .A(net687));
 sg13g2_a22oi_1 _3029_ (.Y(_1044_),
    .B1(net526),
    .B2(net692),
    .A2(net528),
    .A1(\cpu.ctrl.o_ibus_adr[9] ));
 sg13g2_inv_1 _3030_ (.Y(_0284_),
    .A(net693));
 sg13g2_a22oi_1 _3031_ (.Y(_1045_),
    .B1(net523),
    .B2(net712),
    .A2(net531),
    .A1(net707));
 sg13g2_inv_1 _3032_ (.Y(_0285_),
    .A(_1045_));
 sg13g2_a22oi_1 _3033_ (.Y(_1046_),
    .B1(net523),
    .B2(net707),
    .A2(net528),
    .A1(\cpu.ctrl.o_ibus_adr[11] ));
 sg13g2_inv_1 _3034_ (.Y(_0286_),
    .A(net708));
 sg13g2_a22oi_1 _3035_ (.Y(_1047_),
    .B1(net523),
    .B2(net723),
    .A2(net528),
    .A1(net671));
 sg13g2_inv_1 _3036_ (.Y(_0287_),
    .A(_1047_));
 sg13g2_a22oi_1 _3037_ (.Y(_1048_),
    .B1(net522),
    .B2(net671),
    .A2(net527),
    .A1(net650));
 sg13g2_inv_1 _3038_ (.Y(_0288_),
    .A(_1048_));
 sg13g2_a22oi_1 _3039_ (.Y(_1049_),
    .B1(net522),
    .B2(net650),
    .A2(net527),
    .A1(\cpu.ctrl.o_ibus_adr[14] ));
 sg13g2_inv_1 _3040_ (.Y(_0289_),
    .A(net651));
 sg13g2_a22oi_1 _3041_ (.Y(_1050_),
    .B1(net522),
    .B2(net660),
    .A2(net527),
    .A1(net648));
 sg13g2_inv_1 _3042_ (.Y(_0290_),
    .A(_1050_));
 sg13g2_a22oi_1 _3043_ (.Y(_1051_),
    .B1(net522),
    .B2(net648),
    .A2(net527),
    .A1(\cpu.ctrl.o_ibus_adr[16] ));
 sg13g2_inv_1 _3044_ (.Y(_0291_),
    .A(net649));
 sg13g2_a22oi_1 _3045_ (.Y(_1052_),
    .B1(net522),
    .B2(net711),
    .A2(net527),
    .A1(net665));
 sg13g2_inv_1 _3046_ (.Y(_0292_),
    .A(_1052_));
 sg13g2_a22oi_1 _3047_ (.Y(_1053_),
    .B1(net522),
    .B2(net665),
    .A2(net527),
    .A1(\cpu.ctrl.o_ibus_adr[18] ));
 sg13g2_inv_1 _3048_ (.Y(_0293_),
    .A(net666));
 sg13g2_a22oi_1 _3049_ (.Y(_1054_),
    .B1(net522),
    .B2(net734),
    .A2(net528),
    .A1(net674));
 sg13g2_inv_1 _3050_ (.Y(_0294_),
    .A(_1054_));
 sg13g2_a22oi_1 _3051_ (.Y(_1055_),
    .B1(net523),
    .B2(net674),
    .A2(net527),
    .A1(\cpu.ctrl.o_ibus_adr[20] ));
 sg13g2_inv_1 _3052_ (.Y(_0295_),
    .A(net675));
 sg13g2_a22oi_1 _3053_ (.Y(_1056_),
    .B1(net523),
    .B2(net702),
    .A2(net528),
    .A1(net680));
 sg13g2_inv_1 _3054_ (.Y(_0296_),
    .A(_1056_));
 sg13g2_a22oi_1 _3055_ (.Y(_1057_),
    .B1(net523),
    .B2(net680),
    .A2(net528),
    .A1(\cpu.ctrl.o_ibus_adr[22] ));
 sg13g2_inv_1 _3056_ (.Y(_0297_),
    .A(net681));
 sg13g2_a22oi_1 _3057_ (.Y(_1058_),
    .B1(net522),
    .B2(net718),
    .A2(net527),
    .A1(\cpu.ctrl.o_ibus_adr[23] ));
 sg13g2_inv_1 _3058_ (.Y(_0298_),
    .A(net719));
 sg13g2_a22oi_1 _3059_ (.Y(_1059_),
    .B1(net523),
    .B2(net732),
    .A2(net528),
    .A1(\cpu.ctrl.o_ibus_adr[24] ));
 sg13g2_inv_1 _3060_ (.Y(_0299_),
    .A(net733));
 sg13g2_a22oi_1 _3061_ (.Y(_1060_),
    .B1(net526),
    .B2(net858),
    .A2(net529),
    .A1(net700));
 sg13g2_inv_1 _3062_ (.Y(_0300_),
    .A(_1060_));
 sg13g2_a22oi_1 _3063_ (.Y(_1061_),
    .B1(net526),
    .B2(net700),
    .A2(net529),
    .A1(\cpu.ctrl.o_ibus_adr[26] ));
 sg13g2_inv_1 _3064_ (.Y(_0301_),
    .A(net701));
 sg13g2_a22oi_1 _3065_ (.Y(_1062_),
    .B1(net524),
    .B2(net777),
    .A2(net529),
    .A1(net722));
 sg13g2_inv_1 _3066_ (.Y(_0302_),
    .A(_1062_));
 sg13g2_a22oi_1 _3067_ (.Y(_1063_),
    .B1(net524),
    .B2(net722),
    .A2(net531),
    .A1(net717));
 sg13g2_inv_1 _3068_ (.Y(_0303_),
    .A(_1063_));
 sg13g2_a22oi_1 _3069_ (.Y(_1064_),
    .B1(net524),
    .B2(net717),
    .A2(net530),
    .A1(net694));
 sg13g2_inv_1 _3070_ (.Y(_0304_),
    .A(_1064_));
 sg13g2_a22oi_1 _3071_ (.Y(_1065_),
    .B1(net524),
    .B2(net694),
    .A2(net530),
    .A1(\cpu.ctrl.o_ibus_adr[30] ));
 sg13g2_inv_1 _3072_ (.Y(_0305_),
    .A(net695));
 sg13g2_a22oi_1 _3073_ (.Y(_1066_),
    .B1(net524),
    .B2(net728),
    .A2(net530),
    .A1(\cpu.ctrl.o_ibus_adr[31] ));
 sg13g2_inv_1 _3074_ (.Y(_0306_),
    .A(net729));
 sg13g2_o21ai_1 _3075_ (.B1(net530),
    .Y(_1067_),
    .A1(\cpu.ctrl.i_jump ),
    .A2(_0970_));
 sg13g2_a21oi_1 _3076_ (.A1(\cpu.ctrl.i_jump ),
    .A2(_0962_),
    .Y(_1068_),
    .B1(_1067_));
 sg13g2_a21o_1 _3077_ (.A2(net524),
    .A1(net1059),
    .B1(_1068_),
    .X(_0307_));
 sg13g2_mux2_1 _3078_ (.A0(net1158),
    .A1(\cpu.bufreg.data[2] ),
    .S(net544),
    .X(_0308_));
 sg13g2_mux2_1 _3079_ (.A0(net1148),
    .A1(\cpu.bufreg.data[3] ),
    .S(net544),
    .X(_0309_));
 sg13g2_mux2_1 _3080_ (.A0(net1152),
    .A1(net1148),
    .S(net546),
    .X(_0310_));
 sg13g2_mux2_1 _3081_ (.A0(net875),
    .A1(\cpu.bufreg.data[5] ),
    .S(net544),
    .X(_0311_));
 sg13g2_mux2_1 _3082_ (.A0(net1026),
    .A1(net875),
    .S(net544),
    .X(_0312_));
 sg13g2_mux2_1 _3083_ (.A0(net1137),
    .A1(net1026),
    .S(net543),
    .X(_0313_));
 sg13g2_mux2_1 _3084_ (.A0(net1117),
    .A1(\cpu.bufreg.data[8] ),
    .S(net543),
    .X(_0314_));
 sg13g2_mux2_1 _3085_ (.A0(net1048),
    .A1(\cpu.bufreg.data[9] ),
    .S(net543),
    .X(_0315_));
 sg13g2_mux2_1 _3086_ (.A0(net1061),
    .A1(net1048),
    .S(net543),
    .X(_0316_));
 sg13g2_mux2_1 _3087_ (.A0(net713),
    .A1(\cpu.bufreg.data[11] ),
    .S(net543),
    .X(_0317_));
 sg13g2_mux2_1 _3088_ (.A0(net920),
    .A1(net713),
    .S(net541),
    .X(_0318_));
 sg13g2_mux2_1 _3089_ (.A0(net1043),
    .A1(net920),
    .S(net542),
    .X(_0319_));
 sg13g2_mux2_1 _3090_ (.A0(net940),
    .A1(\cpu.bufreg.data[14] ),
    .S(net541),
    .X(_0320_));
 sg13g2_mux2_1 _3091_ (.A0(net1042),
    .A1(net940),
    .S(net541),
    .X(_0321_));
 sg13g2_mux2_1 _3092_ (.A0(net1047),
    .A1(net1042),
    .S(net541),
    .X(_0322_));
 sg13g2_mux2_1 _3093_ (.A0(net1062),
    .A1(net1047),
    .S(net541),
    .X(_0323_));
 sg13g2_mux2_1 _3094_ (.A0(net1011),
    .A1(\cpu.bufreg.data[18] ),
    .S(net541),
    .X(_0324_));
 sg13g2_mux2_1 _3095_ (.A0(net1161),
    .A1(net1011),
    .S(net542),
    .X(_0325_));
 sg13g2_mux2_1 _3096_ (.A0(net976),
    .A1(\cpu.bufreg.data[20] ),
    .S(net542),
    .X(_0326_));
 sg13g2_mux2_1 _3097_ (.A0(net1170),
    .A1(net976),
    .S(net541),
    .X(_0327_));
 sg13g2_mux2_1 _3098_ (.A0(net1163),
    .A1(\cpu.bufreg.data[22] ),
    .S(net541),
    .X(_0328_));
 sg13g2_mux2_1 _3099_ (.A0(net888),
    .A1(\cpu.bufreg.data[23] ),
    .S(net543),
    .X(_0329_));
 sg13g2_mux2_1 _3100_ (.A0(net1182),
    .A1(net888),
    .S(net543),
    .X(_0330_));
 sg13g2_mux2_1 _3101_ (.A0(net931),
    .A1(\cpu.bufreg.data[25] ),
    .S(net544),
    .X(_0331_));
 sg13g2_mux2_1 _3102_ (.A0(net1102),
    .A1(net931),
    .S(net544),
    .X(_0332_));
 sg13g2_mux2_1 _3103_ (.A0(net1126),
    .A1(net1102),
    .S(net544),
    .X(_0333_));
 sg13g2_mux2_1 _3104_ (.A0(net939),
    .A1(net1126),
    .S(net544),
    .X(_0334_));
 sg13g2_mux2_1 _3105_ (.A0(net658),
    .A1(net939),
    .S(net545),
    .X(_0335_));
 sg13g2_nand2_1 _3106_ (.Y(_1069_),
    .A(net658),
    .B(net545));
 sg13g2_o21ai_1 _3107_ (.B1(_1069_),
    .Y(_0336_),
    .A1(_0607_),
    .A2(net545));
 sg13g2_a21oi_1 _3108_ (.A1(_0932_),
    .A2(_0933_),
    .Y(_1070_),
    .B1(_0900_));
 sg13g2_nand2_1 _3109_ (.Y(_1071_),
    .A(_0934_),
    .B(_1070_));
 sg13g2_nor2_1 _3110_ (.A(_0590_),
    .B(_0607_),
    .Y(_1072_));
 sg13g2_a21oi_1 _3111_ (.A1(_0900_),
    .A2(_1072_),
    .Y(_1073_),
    .B1(net545));
 sg13g2_a22oi_1 _3112_ (.Y(_0337_),
    .B1(_1071_),
    .B2(_1073_),
    .A2(net545),
    .A1(_0607_));
 sg13g2_nor2_1 _3113_ (.A(net577),
    .B(net576),
    .Y(_1074_));
 sg13g2_nand2b_1 _3114_ (.Y(_1075_),
    .B(_0929_),
    .A_N(\cpu.alu.cmp_r ));
 sg13g2_o21ai_1 _3115_ (.B1(\cpu.decode.co_mem_word ),
    .Y(_1076_),
    .A1(\cpu.bne_or_bge ),
    .A2(net576));
 sg13g2_nand3b_1 _3116_ (.B(_0952_),
    .C(_1076_),
    .Y(_1077_),
    .A_N(_0951_));
 sg13g2_nand3_1 _3117_ (.B(_1074_),
    .C(_1075_),
    .A(_0949_),
    .Y(_1078_));
 sg13g2_or3_1 _3118_ (.A(_0866_),
    .B(_0895_),
    .C(_1077_),
    .X(_1079_));
 sg13g2_o21ai_1 _3119_ (.B1(_1077_),
    .Y(_1080_),
    .A1(_0866_),
    .A2(_0895_));
 sg13g2_nand3b_1 _3120_ (.B(_1079_),
    .C(_1080_),
    .Y(_1081_),
    .A_N(_1074_));
 sg13g2_a21oi_1 _3121_ (.A1(_1078_),
    .A2(_1081_),
    .Y(_1082_),
    .B1(net549));
 sg13g2_a21o_1 _3122_ (.A2(net549),
    .A1(net1183),
    .B1(_1082_),
    .X(_0338_));
 sg13g2_nand2_1 _3123_ (.Y(_1083_),
    .A(net1236),
    .B(net484));
 sg13g2_o21ai_1 _3124_ (.B1(_1083_),
    .Y(_0339_),
    .A1(_0590_),
    .A2(net483));
 sg13g2_mux2_1 _3125_ (.A0(net995),
    .A1(\cpu.bufreg2.i_dat[31] ),
    .S(net482),
    .X(_0340_));
 sg13g2_nand2b_1 _3126_ (.Y(_1084_),
    .B(net573),
    .A_N(net575));
 sg13g2_o21ai_1 _3127_ (.B1(_1084_),
    .Y(_1085_),
    .A1(net573),
    .A2(\cpu.decode.opcode[1] ));
 sg13g2_a21oi_1 _3128_ (.A1(_0881_),
    .A2(_1085_),
    .Y(_1086_),
    .B1(net550));
 sg13g2_nor2b_1 _3129_ (.A(net548),
    .B_N(\cpu.immdec.imm19_12_20[0] ),
    .Y(_1087_));
 sg13g2_a21oi_1 _3130_ (.A1(net1280),
    .A2(net548),
    .Y(_1088_),
    .B1(_1087_));
 sg13g2_nand2_2 _3131_ (.Y(_1089_),
    .A(net1285),
    .B(net490));
 sg13g2_o21ai_1 _3132_ (.B1(_1089_),
    .Y(_0341_),
    .A1(net489),
    .A2(net1281));
 sg13g2_nor2b_1 _3133_ (.A(net548),
    .B_N(net1280),
    .Y(_1090_));
 sg13g2_a21oi_1 _3134_ (.A1(\cpu.immdec.imm19_12_20[2] ),
    .A2(net548),
    .Y(_1091_),
    .B1(_1090_));
 sg13g2_nand2_1 _3135_ (.Y(_1092_),
    .A(net1286),
    .B(net489));
 sg13g2_o21ai_1 _3136_ (.B1(_1092_),
    .Y(_0342_),
    .A1(net488),
    .A2(_1091_));
 sg13g2_nor2b_1 _3137_ (.A(net547),
    .B_N(\cpu.immdec.imm19_12_20[2] ),
    .Y(_1093_));
 sg13g2_a21oi_1 _3138_ (.A1(net1174),
    .A2(net547),
    .Y(_1094_),
    .B1(_1093_));
 sg13g2_nand2_1 _3139_ (.Y(_1095_),
    .A(net1239),
    .B(net487));
 sg13g2_o21ai_1 _3140_ (.B1(_1095_),
    .Y(_0343_),
    .A1(net487),
    .A2(_1094_));
 sg13g2_nor2b_1 _3141_ (.A(net548),
    .B_N(net1174),
    .Y(_1096_));
 sg13g2_a21oi_1 _3142_ (.A1(\cpu.csr_imm ),
    .A2(net547),
    .Y(_1097_),
    .B1(_1096_));
 sg13g2_nand2_1 _3143_ (.Y(_1098_),
    .A(net829),
    .B(net489));
 sg13g2_o21ai_1 _3144_ (.B1(_1098_),
    .Y(_0344_),
    .A1(net489),
    .A2(net1175));
 sg13g2_nand2_1 _3145_ (.Y(_1099_),
    .A(net1254),
    .B(net547));
 sg13g2_nor2_2 _3146_ (.A(net488),
    .B(net547),
    .Y(_1100_));
 sg13g2_a22oi_1 _3147_ (.Y(_1101_),
    .B1(_1100_),
    .B2(\cpu.csr_imm ),
    .A2(net487),
    .A1(net772));
 sg13g2_o21ai_1 _3148_ (.B1(_1101_),
    .Y(_0345_),
    .A1(net487),
    .A2(_1099_));
 sg13g2_and3_1 _3149_ (.X(_1102_),
    .A(\cpu.immdec.imm19_12_20[6] ),
    .B(_1021_),
    .C(net547));
 sg13g2_a221oi_1 _3150_ (.B2(net1254),
    .C1(_1102_),
    .B1(_1100_),
    .A1(net1305),
    .Y(_1103_),
    .A2(net487));
 sg13g2_inv_1 _3151_ (.Y(_0346_),
    .A(net1306));
 sg13g2_and3_1 _3152_ (.X(_1104_),
    .A(\cpu.immdec.imm19_12_20[7] ),
    .B(_1021_),
    .C(net547));
 sg13g2_a221oi_1 _3153_ (.B2(\cpu.immdec.imm19_12_20[6] ),
    .C1(_1104_),
    .B1(_1100_),
    .A1(net1297),
    .Y(_1105_),
    .A2(net487));
 sg13g2_inv_1 _3154_ (.Y(_0347_),
    .A(net1298));
 sg13g2_nand2_1 _3155_ (.Y(_1106_),
    .A(net869),
    .B(net547));
 sg13g2_a22oi_1 _3156_ (.Y(_1107_),
    .B1(_1100_),
    .B2(\cpu.immdec.imm19_12_20[7] ),
    .A2(net488),
    .A1(\cpu.bufreg2.i_dat[18] ));
 sg13g2_o21ai_1 _3157_ (.B1(_1107_),
    .Y(_0348_),
    .A1(net487),
    .A2(_1106_));
 sg13g2_o21ai_1 _3158_ (.B1(_1086_),
    .Y(_1108_),
    .A1(net570),
    .A2(\cpu.immdec.imm24_20[0] ));
 sg13g2_a21oi_1 _3159_ (.A1(net569),
    .A2(_0882_),
    .Y(_1109_),
    .B1(_1108_));
 sg13g2_mux2_1 _3160_ (.A0(_1109_),
    .A1(net1116),
    .S(net489),
    .X(_1110_));
 sg13g2_a21o_1 _3161_ (.A2(_1100_),
    .A1(net869),
    .B1(_1110_),
    .X(_0349_));
 sg13g2_nor2_1 _3162_ (.A(net550),
    .B(_0882_),
    .Y(_1111_));
 sg13g2_a21oi_1 _3163_ (.A1(\cpu.immdec.imm7 ),
    .A2(net550),
    .Y(_1112_),
    .B1(_1111_));
 sg13g2_o21ai_1 _3164_ (.B1(_1025_),
    .Y(_0350_),
    .A1(net482),
    .A2(_1112_));
 sg13g2_nor2b_1 _3165_ (.A(net482),
    .B_N(net575),
    .Y(_1113_));
 sg13g2_nor2_1 _3166_ (.A(_0580_),
    .B(_0909_),
    .Y(_1114_));
 sg13g2_a22oi_1 _3167_ (.Y(_1115_),
    .B1(_1113_),
    .B2(_1114_),
    .A2(_0939_),
    .A1(net549));
 sg13g2_mux2_1 _3168_ (.A0(net824),
    .A1(\cpu.bufreg2.i_dat[25] ),
    .S(net490),
    .X(_1116_));
 sg13g2_mux2_1 _3169_ (.A0(net1252),
    .A1(_1116_),
    .S(_1115_),
    .X(_0351_));
 sg13g2_mux2_1 _3170_ (.A0(net797),
    .A1(\cpu.bufreg2.i_dat[26] ),
    .S(net490),
    .X(_1117_));
 sg13g2_mux2_1 _3171_ (.A0(net824),
    .A1(_1117_),
    .S(_1115_),
    .X(_0352_));
 sg13g2_mux2_1 _3172_ (.A0(net773),
    .A1(\cpu.bufreg2.i_dat[27] ),
    .S(net490),
    .X(_1118_));
 sg13g2_mux2_1 _3173_ (.A0(net797),
    .A1(_1118_),
    .S(_1115_),
    .X(_0353_));
 sg13g2_mux2_1 _3174_ (.A0(\cpu.immdec.imm30_25[4] ),
    .A1(\cpu.bufreg2.i_dat[28] ),
    .S(net484),
    .X(_1119_));
 sg13g2_mux2_1 _3175_ (.A0(net773),
    .A1(_1119_),
    .S(_1115_),
    .X(_0354_));
 sg13g2_mux2_1 _3176_ (.A0(net795),
    .A1(\cpu.bufreg2.i_dat[29] ),
    .S(net484),
    .X(_1120_));
 sg13g2_mux2_1 _3177_ (.A0(net807),
    .A1(_1120_),
    .S(_1115_),
    .X(_0355_));
 sg13g2_nor2b_1 _3178_ (.A(net575),
    .B_N(net569),
    .Y(_1121_));
 sg13g2_a21oi_1 _3179_ (.A1(net573),
    .A2(net574),
    .Y(_1122_),
    .B1(\cpu.decode.opcode[1] ));
 sg13g2_nor2_1 _3180_ (.A(\cpu.immdec.imm19_12_20[0] ),
    .B(_1122_),
    .Y(_1123_));
 sg13g2_or2_1 _3181_ (.X(_1124_),
    .B(_1123_),
    .A(_1121_));
 sg13g2_a21oi_1 _3182_ (.A1(_0882_),
    .A2(_1122_),
    .Y(_1125_),
    .B1(_1124_));
 sg13g2_a21oi_1 _3183_ (.A1(\cpu.immdec.imm7 ),
    .A2(_1121_),
    .Y(_1126_),
    .B1(_1125_));
 sg13g2_o21ai_1 _3184_ (.B1(_1083_),
    .Y(_1127_),
    .A1(net482),
    .A2(_1126_));
 sg13g2_mux2_1 _3185_ (.A0(net795),
    .A1(_1127_),
    .S(_1115_),
    .X(_0356_));
 sg13g2_nor2_1 _3186_ (.A(_0020_),
    .B(_0578_),
    .Y(_1128_));
 sg13g2_a21oi_2 _3187_ (.B1(net550),
    .Y(_1129_),
    .A2(_1128_),
    .A1(_0880_));
 sg13g2_nor2_1 _3188_ (.A(_0583_),
    .B(_1129_),
    .Y(_1130_));
 sg13g2_a21oi_1 _3189_ (.A1(net1217),
    .A2(_1129_),
    .Y(_1131_),
    .B1(_1130_));
 sg13g2_o21ai_1 _3190_ (.B1(_1089_),
    .Y(_0357_),
    .A1(net486),
    .A2(_1131_));
 sg13g2_nand2_1 _3191_ (.Y(_1132_),
    .A(\cpu.immdec.imm24_20[2] ),
    .B(_1129_));
 sg13g2_nor2_2 _3192_ (.A(net485),
    .B(_1129_),
    .Y(_1133_));
 sg13g2_a22oi_1 _3193_ (.Y(_1134_),
    .B1(_1133_),
    .B2(net1217),
    .A2(net485),
    .A1(\cpu.bufreg2.i_dat[21] ));
 sg13g2_o21ai_1 _3194_ (.B1(net1218),
    .Y(_0358_),
    .A1(net486),
    .A2(_1132_));
 sg13g2_and3_1 _3195_ (.X(_1135_),
    .A(\cpu.immdec.imm24_20[3] ),
    .B(_1021_),
    .C(_1129_));
 sg13g2_a221oi_1 _3196_ (.B2(\cpu.immdec.imm24_20[2] ),
    .C1(_1135_),
    .B1(_1133_),
    .A1(net1332),
    .Y(_1136_),
    .A2(net485));
 sg13g2_inv_1 _3197_ (.Y(_0359_),
    .A(net1333));
 sg13g2_nand2_1 _3198_ (.Y(_1137_),
    .A(net1051),
    .B(_1129_));
 sg13g2_a22oi_1 _3199_ (.Y(_1138_),
    .B1(_1133_),
    .B2(\cpu.immdec.imm24_20[3] ),
    .A2(net485),
    .A1(\cpu.bufreg2.i_dat[23] ));
 sg13g2_o21ai_1 _3200_ (.B1(_1138_),
    .Y(_0360_),
    .A1(net485),
    .A2(_1137_));
 sg13g2_nor2_1 _3201_ (.A(_1032_),
    .B(_1133_),
    .Y(_1139_));
 sg13g2_a221oi_1 _3202_ (.B2(net1051),
    .C1(_1139_),
    .B1(_1133_),
    .A1(net1277),
    .Y(_1140_),
    .A2(net485));
 sg13g2_inv_1 _3203_ (.Y(_0361_),
    .A(_1140_));
 sg13g2_o21ai_1 _3204_ (.B1(_1089_),
    .Y(_0362_),
    .A1(_0581_),
    .A2(net485));
 sg13g2_o21ai_1 _3205_ (.B1(_1092_),
    .Y(_0363_),
    .A1(_0575_),
    .A2(net482));
 sg13g2_mux2_1 _3206_ (.A0(net577),
    .A1(net1239),
    .S(net485),
    .X(_0364_));
 sg13g2_mux2_1 _3207_ (.A0(net576),
    .A1(net829),
    .S(net482),
    .X(_0365_));
 sg13g2_a21o_1 _3208_ (.A2(net482),
    .A1(net1313),
    .B1(_1113_),
    .X(_0366_));
 sg13g2_mux2_1 _3209_ (.A0(\cpu.decode.opcode[1] ),
    .A1(net1302),
    .S(net484),
    .X(_0367_));
 sg13g2_mux2_1 _3210_ (.A0(net572),
    .A1(net1295),
    .S(net483),
    .X(_0368_));
 sg13g2_nor2_1 _3211_ (.A(net571),
    .B(net483),
    .Y(_1141_));
 sg13g2_a21oi_1 _3212_ (.A1(_0595_),
    .A2(net483),
    .Y(_0369_),
    .B1(_1141_));
 sg13g2_mux2_1 _3213_ (.A0(net569),
    .A1(net1268),
    .S(net483),
    .X(_0370_));
 sg13g2_and2_1 _3214_ (.A(_0563_),
    .B(_0623_),
    .X(_1142_));
 sg13g2_a22oi_1 _3215_ (.Y(_1143_),
    .B1(_0711_),
    .B2(_1142_),
    .A2(_0594_),
    .A1(net571));
 sg13g2_o21ai_1 _3216_ (.B1(\cpu.mem_bytecnt[0] ),
    .Y(_1144_),
    .A1(\cpu.mem_bytecnt[1] ),
    .A2(\cpu.bufreg.data[1] ));
 sg13g2_a21oi_1 _3217_ (.A1(\cpu.mem_bytecnt[1] ),
    .A2(\cpu.bufreg.data[1] ),
    .Y(_1145_),
    .B1(net549));
 sg13g2_o21ai_1 _3218_ (.B1(_1145_),
    .Y(_1146_),
    .A1(_0582_),
    .A2(_1144_));
 sg13g2_and3_1 _3219_ (.X(_1147_),
    .A(_0918_),
    .B(net472),
    .C(_1146_));
 sg13g2_nand2b_2 _3220_ (.Y(_1148_),
    .B(_0900_),
    .A_N(_0918_));
 sg13g2_nand2_1 _3221_ (.Y(_1149_),
    .A(\cpu.bufreg2.dat[1] ),
    .B(_1148_));
 sg13g2_o21ai_1 _3222_ (.B1(_1149_),
    .Y(_1150_),
    .A1(_0593_),
    .A2(_1148_));
 sg13g2_mux2_1 _3223_ (.A0(\cpu.bufreg2.i_dat[0] ),
    .A1(_1150_),
    .S(net472),
    .X(_1151_));
 sg13g2_mux2_1 _3224_ (.A0(_1151_),
    .A1(net1323),
    .S(net461),
    .X(_0371_));
 sg13g2_xor2_1 _3225_ (.B(\cpu.bufreg2.dat[0] ),
    .A(\cpu.bufreg2.dat[1] ),
    .X(_1152_));
 sg13g2_nor2_1 _3226_ (.A(\cpu.bufreg2.i_dat[1] ),
    .B(net471),
    .Y(_1153_));
 sg13g2_o21ai_1 _3227_ (.B1(net471),
    .Y(_1154_),
    .A1(_1148_),
    .A2(_1152_));
 sg13g2_a21oi_1 _3228_ (.A1(net1317),
    .A2(net539),
    .Y(_1155_),
    .B1(_1154_));
 sg13g2_nor3_1 _3229_ (.A(net460),
    .B(_1153_),
    .C(_1155_),
    .Y(_1156_));
 sg13g2_a21o_1 _3230_ (.A2(net460),
    .A1(net1325),
    .B1(_1156_),
    .X(_0372_));
 sg13g2_nor3_2 _3231_ (.A(\cpu.bufreg2.dat[2] ),
    .B(\cpu.bufreg2.dat[1] ),
    .C(\cpu.bufreg2.dat[0] ),
    .Y(_1157_));
 sg13g2_o21ai_1 _3232_ (.B1(\cpu.bufreg2.dat[2] ),
    .Y(_1158_),
    .A1(\cpu.bufreg2.dat[1] ),
    .A2(\cpu.bufreg2.dat[0] ));
 sg13g2_nor2b_1 _3233_ (.A(_1157_),
    .B_N(_1158_),
    .Y(_1159_));
 sg13g2_nor2_1 _3234_ (.A(net1313),
    .B(net471),
    .Y(_1160_));
 sg13g2_o21ai_1 _3235_ (.B1(net471),
    .Y(_1161_),
    .A1(net539),
    .A2(_1159_));
 sg13g2_a21oi_1 _3236_ (.A1(net1300),
    .A2(net539),
    .Y(_1162_),
    .B1(_1161_));
 sg13g2_nor3_1 _3237_ (.A(net460),
    .B(_1160_),
    .C(_1162_),
    .Y(_1163_));
 sg13g2_a21o_1 _3238_ (.A2(net460),
    .A1(net1317),
    .B1(_1163_),
    .X(_0373_));
 sg13g2_nor2b_1 _3239_ (.A(\cpu.bufreg2.dat[3] ),
    .B_N(_1157_),
    .Y(_1164_));
 sg13g2_xnor2_1 _3240_ (.Y(_1165_),
    .A(\cpu.bufreg2.dat[3] ),
    .B(_1157_));
 sg13g2_nor2_1 _3241_ (.A(\cpu.bufreg2.i_dat[3] ),
    .B(net471),
    .Y(_1166_));
 sg13g2_o21ai_1 _3242_ (.B1(net471),
    .Y(_1167_),
    .A1(net539),
    .A2(_1165_));
 sg13g2_a21oi_1 _3243_ (.A1(\cpu.bufreg2.dat[4] ),
    .A2(net539),
    .Y(_1168_),
    .B1(_1167_));
 sg13g2_nor3_1 _3244_ (.A(net460),
    .B(_1166_),
    .C(_1168_),
    .Y(_1169_));
 sg13g2_a21o_1 _3245_ (.A2(net460),
    .A1(net1300),
    .B1(_1169_),
    .X(_0374_));
 sg13g2_nor2b_1 _3246_ (.A(\cpu.bufreg2.dat[4] ),
    .B_N(_1164_),
    .Y(_1170_));
 sg13g2_xnor2_1 _3247_ (.Y(_1171_),
    .A(\cpu.bufreg2.dat[4] ),
    .B(_1164_));
 sg13g2_nor2_1 _3248_ (.A(net1295),
    .B(net471),
    .Y(_1172_));
 sg13g2_o21ai_1 _3249_ (.B1(net471),
    .Y(_1173_),
    .A1(net539),
    .A2(_1171_));
 sg13g2_a21oi_1 _3250_ (.A1(net1279),
    .A2(net539),
    .Y(_1174_),
    .B1(_1173_));
 sg13g2_nor3_1 _3251_ (.A(net460),
    .B(_1172_),
    .C(_1174_),
    .Y(_1175_));
 sg13g2_a21o_1 _3252_ (.A2(net460),
    .A1(net1318),
    .B1(_1175_),
    .X(_0375_));
 sg13g2_o21ai_1 _3253_ (.B1(net696),
    .Y(_1176_),
    .A1(_0878_),
    .A2(_0918_));
 sg13g2_xnor2_1 _3254_ (.Y(_1177_),
    .A(\cpu.bufreg2.dat[5] ),
    .B(_1170_));
 sg13g2_mux2_1 _3255_ (.A0(_1177_),
    .A1(_1176_),
    .S(net539),
    .X(_1178_));
 sg13g2_mux2_1 _3256_ (.A0(_0595_),
    .A1(_1178_),
    .S(net472),
    .X(_1179_));
 sg13g2_nand2_1 _3257_ (.Y(_1180_),
    .A(net1279),
    .B(net461));
 sg13g2_o21ai_1 _3258_ (.B1(_1180_),
    .Y(_0376_),
    .A1(net461),
    .A2(_1179_));
 sg13g2_nand2_1 _3259_ (.Y(_1181_),
    .A(net696),
    .B(net461));
 sg13g2_nand2_1 _3260_ (.Y(_1182_),
    .A(_0596_),
    .B(net472));
 sg13g2_o21ai_1 _3261_ (.B1(_1182_),
    .Y(_1183_),
    .A1(\cpu.bufreg2.i_dat[6] ),
    .A2(net472));
 sg13g2_o21ai_1 _3262_ (.B1(_1181_),
    .Y(_0377_),
    .A1(net461),
    .A2(_1183_));
 sg13g2_nand2b_1 _3263_ (.Y(_1184_),
    .B(\cpu.bufreg2.i_dat[7] ),
    .A_N(net472));
 sg13g2_a21oi_1 _3264_ (.A1(\cpu.bufreg2.dat[8] ),
    .A2(net472),
    .Y(_1185_),
    .B1(net462));
 sg13g2_a22oi_1 _3265_ (.Y(_0378_),
    .B1(_1184_),
    .B2(_1185_),
    .A2(net461),
    .A1(_0596_));
 sg13g2_nand2_1 _3266_ (.Y(_1186_),
    .A(net1207),
    .B(net469));
 sg13g2_nand2_1 _3267_ (.Y(_1187_),
    .A(_0597_),
    .B(net479));
 sg13g2_o21ai_1 _3268_ (.B1(_1187_),
    .Y(_1188_),
    .A1(\cpu.bufreg2.i_dat[8] ),
    .A2(net476));
 sg13g2_o21ai_1 _3269_ (.B1(_1186_),
    .Y(_0379_),
    .A1(net469),
    .A2(_1188_));
 sg13g2_nand2b_1 _3270_ (.Y(_1189_),
    .B(net1057),
    .A_N(net479));
 sg13g2_a21oi_1 _3271_ (.A1(net813),
    .A2(net477),
    .Y(_1190_),
    .B1(net466));
 sg13g2_a22oi_1 _3272_ (.Y(_0380_),
    .B1(_1189_),
    .B2(_1190_),
    .A2(net467),
    .A1(_0597_));
 sg13g2_nand2_1 _3273_ (.Y(_1191_),
    .A(net813),
    .B(net465));
 sg13g2_nand2_1 _3274_ (.Y(_1192_),
    .A(_0598_),
    .B(net477));
 sg13g2_o21ai_1 _3275_ (.B1(_1192_),
    .Y(_1193_),
    .A1(\cpu.bufreg2.i_dat[10] ),
    .A2(net477));
 sg13g2_o21ai_1 _3276_ (.B1(_1191_),
    .Y(_0381_),
    .A1(net465),
    .A2(_1193_));
 sg13g2_nand2b_1 _3277_ (.Y(_1194_),
    .B(net789),
    .A_N(net477));
 sg13g2_a21oi_1 _3278_ (.A1(net786),
    .A2(net478),
    .Y(_1195_),
    .B1(net465));
 sg13g2_a22oi_1 _3279_ (.Y(_0382_),
    .B1(_1194_),
    .B2(_1195_),
    .A2(net466),
    .A1(_0598_));
 sg13g2_nand2_1 _3280_ (.Y(_1196_),
    .A(net786),
    .B(net465));
 sg13g2_nand2_1 _3281_ (.Y(_1197_),
    .A(_0599_),
    .B(net478));
 sg13g2_o21ai_1 _3282_ (.B1(_1197_),
    .Y(_1198_),
    .A1(\cpu.bufreg2.i_dat[12] ),
    .A2(net478));
 sg13g2_o21ai_1 _3283_ (.B1(_1196_),
    .Y(_0383_),
    .A1(net466),
    .A2(_1198_));
 sg13g2_nand2b_1 _3284_ (.Y(_1199_),
    .B(\cpu.bufreg2.i_dat[13] ),
    .A_N(net479));
 sg13g2_a21oi_1 _3285_ (.A1(net698),
    .A2(net478),
    .Y(_1200_),
    .B1(net466));
 sg13g2_a22oi_1 _3286_ (.Y(_0384_),
    .B1(_1199_),
    .B2(_1200_),
    .A2(net466),
    .A1(_0599_));
 sg13g2_nand2_1 _3287_ (.Y(_1201_),
    .A(net698),
    .B(net466));
 sg13g2_nand2_1 _3288_ (.Y(_1202_),
    .A(_0600_),
    .B(net477));
 sg13g2_o21ai_1 _3289_ (.B1(_1202_),
    .Y(_1203_),
    .A1(\cpu.bufreg2.i_dat[14] ),
    .A2(net479));
 sg13g2_o21ai_1 _3290_ (.B1(_1201_),
    .Y(_0385_),
    .A1(net466),
    .A2(_1203_));
 sg13g2_nand2b_1 _3291_ (.Y(_1204_),
    .B(net772),
    .A_N(net477));
 sg13g2_a21oi_1 _3292_ (.A1(\cpu.bufreg2.dat[16] ),
    .A2(net478),
    .Y(_1205_),
    .B1(net465));
 sg13g2_a22oi_1 _3293_ (.Y(_0386_),
    .B1(_1204_),
    .B2(_1205_),
    .A2(net465),
    .A1(_0600_));
 sg13g2_nand2_1 _3294_ (.Y(_1206_),
    .A(net1242),
    .B(net465));
 sg13g2_nand2_1 _3295_ (.Y(_1207_),
    .A(_0601_),
    .B(net477));
 sg13g2_o21ai_1 _3296_ (.B1(_1207_),
    .Y(_1208_),
    .A1(\cpu.bufreg2.i_dat[16] ),
    .A2(net477));
 sg13g2_o21ai_1 _3297_ (.B1(_1206_),
    .Y(_0387_),
    .A1(net465),
    .A2(_1208_));
 sg13g2_nand2b_1 _3298_ (.Y(_1209_),
    .B(\cpu.bufreg2.i_dat[17] ),
    .A_N(net478));
 sg13g2_a21oi_1 _3299_ (.A1(net672),
    .A2(net478),
    .Y(_1210_),
    .B1(net467));
 sg13g2_a22oi_1 _3300_ (.Y(_0388_),
    .B1(_1209_),
    .B2(_1210_),
    .A2(net467),
    .A1(_0601_));
 sg13g2_nand2_1 _3301_ (.Y(_1211_),
    .A(net672),
    .B(net468));
 sg13g2_nand2_1 _3302_ (.Y(_1212_),
    .A(_0602_),
    .B(net480));
 sg13g2_o21ai_1 _3303_ (.B1(_1212_),
    .Y(_1213_),
    .A1(\cpu.bufreg2.i_dat[18] ),
    .A2(net480));
 sg13g2_o21ai_1 _3304_ (.B1(_1211_),
    .Y(_0389_),
    .A1(net468),
    .A2(_1213_));
 sg13g2_nand2b_1 _3305_ (.Y(_1214_),
    .B(net1116),
    .A_N(net480));
 sg13g2_a21oi_1 _3306_ (.A1(net705),
    .A2(net480),
    .Y(_1215_),
    .B1(net468));
 sg13g2_a22oi_1 _3307_ (.Y(_0390_),
    .B1(_1214_),
    .B2(_1215_),
    .A2(net468),
    .A1(_0602_));
 sg13g2_nand2_1 _3308_ (.Y(_1216_),
    .A(net705),
    .B(net468));
 sg13g2_nand2_1 _3309_ (.Y(_1217_),
    .A(_0603_),
    .B(net480));
 sg13g2_o21ai_1 _3310_ (.B1(_1217_),
    .Y(_1218_),
    .A1(\cpu.bufreg2.i_dat[20] ),
    .A2(net480));
 sg13g2_o21ai_1 _3311_ (.B1(_1216_),
    .Y(_0391_),
    .A1(net468),
    .A2(_1218_));
 sg13g2_nand2b_1 _3312_ (.Y(_1219_),
    .B(\cpu.bufreg2.i_dat[21] ),
    .A_N(net475));
 sg13g2_a21oi_1 _3313_ (.A1(net784),
    .A2(net475),
    .Y(_1220_),
    .B1(net463));
 sg13g2_a22oi_1 _3314_ (.Y(_0392_),
    .B1(_1219_),
    .B2(_1220_),
    .A2(net464),
    .A1(_0603_));
 sg13g2_nand2_1 _3315_ (.Y(_1221_),
    .A(net784),
    .B(net463));
 sg13g2_nand2b_1 _3316_ (.Y(_1222_),
    .B(net474),
    .A_N(net757));
 sg13g2_o21ai_1 _3317_ (.B1(_1222_),
    .Y(_1223_),
    .A1(\cpu.bufreg2.i_dat[22] ),
    .A2(net474));
 sg13g2_o21ai_1 _3318_ (.B1(_1221_),
    .Y(_0393_),
    .A1(net464),
    .A2(_1223_));
 sg13g2_nor2b_1 _3319_ (.A(net476),
    .B_N(\cpu.bufreg2.i_dat[23] ),
    .Y(_1224_));
 sg13g2_a21oi_1 _3320_ (.A1(\cpu.bufreg2.dat[24] ),
    .A2(net476),
    .Y(_1225_),
    .B1(_1224_));
 sg13g2_nand2_1 _3321_ (.Y(_1226_),
    .A(net757),
    .B(net464));
 sg13g2_o21ai_1 _3322_ (.B1(_1226_),
    .Y(_0394_),
    .A1(net464),
    .A2(_1225_));
 sg13g2_nand2b_1 _3323_ (.Y(_1227_),
    .B(\cpu.bufreg2.i_dat[24] ),
    .A_N(net474));
 sg13g2_a21oi_1 _3324_ (.A1(net690),
    .A2(net475),
    .Y(_1228_),
    .B1(net463));
 sg13g2_a22oi_1 _3325_ (.Y(_0395_),
    .B1(_1227_),
    .B2(_1228_),
    .A2(net463),
    .A1(_0592_));
 sg13g2_nand2_1 _3326_ (.Y(_1229_),
    .A(net690),
    .B(net464));
 sg13g2_nand2_1 _3327_ (.Y(_1230_),
    .A(_0604_),
    .B(net474));
 sg13g2_o21ai_1 _3328_ (.B1(_1230_),
    .Y(_1231_),
    .A1(\cpu.bufreg2.i_dat[25] ),
    .A2(net474));
 sg13g2_o21ai_1 _3329_ (.B1(_1229_),
    .Y(_0396_),
    .A1(net463),
    .A2(_1231_));
 sg13g2_nand2b_1 _3330_ (.Y(_1232_),
    .B(\cpu.bufreg2.i_dat[26] ),
    .A_N(net474));
 sg13g2_a21oi_1 _3331_ (.A1(net780),
    .A2(net475),
    .Y(_1233_),
    .B1(net463));
 sg13g2_a22oi_1 _3332_ (.Y(_0397_),
    .B1(_1232_),
    .B2(_1233_),
    .A2(net463),
    .A1(_0604_));
 sg13g2_nand2_1 _3333_ (.Y(_1234_),
    .A(net780),
    .B(net463));
 sg13g2_nand2_1 _3334_ (.Y(_1235_),
    .A(_0605_),
    .B(net474));
 sg13g2_o21ai_1 _3335_ (.B1(_1235_),
    .Y(_1236_),
    .A1(\cpu.bufreg2.i_dat[27] ),
    .A2(net474));
 sg13g2_o21ai_1 _3336_ (.B1(_1234_),
    .Y(_0398_),
    .A1(net464),
    .A2(_1236_));
 sg13g2_nand2b_1 _3337_ (.Y(_1237_),
    .B(\cpu.bufreg2.i_dat[28] ),
    .A_N(net473));
 sg13g2_a21oi_1 _3338_ (.A1(net775),
    .A2(net473),
    .Y(_1238_),
    .B1(net462));
 sg13g2_a22oi_1 _3339_ (.Y(_0399_),
    .B1(_1237_),
    .B2(_1238_),
    .A2(net462),
    .A1(_0605_));
 sg13g2_nand2_1 _3340_ (.Y(_1239_),
    .A(net775),
    .B(net470));
 sg13g2_nand2_1 _3341_ (.Y(_1240_),
    .A(_0606_),
    .B(net473));
 sg13g2_o21ai_1 _3342_ (.B1(_1240_),
    .Y(_1241_),
    .A1(\cpu.bufreg2.i_dat[29] ),
    .A2(net473));
 sg13g2_o21ai_1 _3343_ (.B1(_1239_),
    .Y(_0400_),
    .A1(net462),
    .A2(_1241_));
 sg13g2_nand2b_1 _3344_ (.Y(_1242_),
    .B(\cpu.bufreg2.i_dat[30] ),
    .A_N(net473));
 sg13g2_a21oi_1 _3345_ (.A1(net759),
    .A2(net473),
    .Y(_1243_),
    .B1(net462));
 sg13g2_a22oi_1 _3346_ (.Y(_0401_),
    .B1(_1242_),
    .B2(_1243_),
    .A2(net462),
    .A1(_0606_));
 sg13g2_nand2_1 _3347_ (.Y(_1244_),
    .A(net759),
    .B(net462));
 sg13g2_o21ai_1 _3348_ (.B1(net481),
    .Y(_1245_),
    .A1(_0875_),
    .A2(_0891_));
 sg13g2_o21ai_1 _3349_ (.B1(_1245_),
    .Y(_1246_),
    .A1(\cpu.bufreg2.i_dat[31] ),
    .A2(net481));
 sg13g2_o21ai_1 _3350_ (.B1(_1244_),
    .Y(_0402_),
    .A1(net462),
    .A2(_1246_));
 sg13g2_nor3_1 _3351_ (.A(_0465_),
    .B(_0878_),
    .C(_0900_),
    .Y(_0403_));
 sg13g2_nand2_2 _3352_ (.Y(_1247_),
    .A(net584),
    .B(_0878_));
 sg13g2_nand3_1 _3353_ (.B(net584),
    .C(_0878_),
    .A(net1222),
    .Y(_1248_));
 sg13g2_nand2b_1 _3354_ (.Y(_0404_),
    .B(_1248_),
    .A_N(_0403_));
 sg13g2_a21oi_1 _3355_ (.A1(net1140),
    .A2(net1250),
    .Y(_1249_),
    .B1(net1211));
 sg13g2_a21o_1 _3356_ (.A2(_1178_),
    .A1(net576),
    .B1(_0918_),
    .X(_1250_));
 sg13g2_nand3_1 _3357_ (.B(_0017_),
    .C(\cpu.bufreg.i_sh_signed ),
    .A(_0564_),
    .Y(_1251_));
 sg13g2_nand2b_1 _3358_ (.Y(_1252_),
    .B(_1251_),
    .A_N(net577));
 sg13g2_a21oi_1 _3359_ (.A1(net572),
    .A2(_1252_),
    .Y(_1253_),
    .B1(net569));
 sg13g2_nand3_1 _3360_ (.B(_1250_),
    .C(_1253_),
    .A(net472),
    .Y(_1254_));
 sg13g2_nand4_1 _3361_ (.B(net584),
    .C(net549),
    .A(net1222),
    .Y(_1255_),
    .D(_1254_));
 sg13g2_o21ai_1 _3362_ (.B1(_1255_),
    .Y(_0405_),
    .A1(_1247_),
    .A2(_1249_));
 sg13g2_and2_1 _3363_ (.A(net582),
    .B(net1249),
    .X(_0406_));
 sg13g2_and2_1 _3364_ (.A(net582),
    .B(net819),
    .X(_0407_));
 sg13g2_and2_1 _3365_ (.A(net582),
    .B(net771),
    .X(_0408_));
 sg13g2_nand3_1 _3366_ (.B(net584),
    .C(_0878_),
    .A(net1103),
    .Y(_1256_));
 sg13g2_and3_1 _3367_ (.X(_1257_),
    .A(\cpu.bne_or_bge ),
    .B(_1078_),
    .C(_1081_));
 sg13g2_a21oi_1 _3368_ (.A1(_1078_),
    .A2(_1081_),
    .Y(_1258_),
    .B1(\cpu.bne_or_bge ));
 sg13g2_nor3_1 _3369_ (.A(_0578_),
    .B(_1257_),
    .C(_1258_),
    .Y(_1259_));
 sg13g2_nand2_1 _3370_ (.Y(_1260_),
    .A(_0576_),
    .B(_0403_));
 sg13g2_o21ai_1 _3371_ (.B1(_1256_),
    .Y(_0409_),
    .A1(_1259_),
    .A2(_1260_));
 sg13g2_o21ai_1 _3372_ (.B1(net583),
    .Y(_1261_),
    .A1(net1211),
    .A2(\cpu.state.o_cnt[2] ));
 sg13g2_a21oi_1 _3373_ (.A1(net1211),
    .A2(\cpu.state.o_cnt[2] ),
    .Y(_0410_),
    .B1(_1261_));
 sg13g2_a21oi_1 _3374_ (.A1(net1211),
    .A2(\cpu.state.o_cnt[2] ),
    .Y(_1262_),
    .B1(net1292));
 sg13g2_nand2_1 _3375_ (.Y(_1263_),
    .A(net583),
    .B(_0877_));
 sg13g2_nor2_1 _3376_ (.A(net1293),
    .B(_1263_),
    .Y(_0411_));
 sg13g2_a21oi_1 _3377_ (.A1(_0574_),
    .A2(_0877_),
    .Y(_0412_),
    .B1(_1247_));
 sg13g2_o21ai_1 _3378_ (.B1(\dut.xfer.resetn ),
    .Y(_1264_),
    .A1(net634),
    .A2(net536));
 sg13g2_a21oi_1 _3379_ (.A1(_0544_),
    .A2(net536),
    .Y(_0414_),
    .B1(_1264_));
 sg13g2_o21ai_1 _3380_ (.B1(net558),
    .Y(_1265_),
    .A1(net633),
    .A2(net536));
 sg13g2_a21oi_1 _3381_ (.A1(_0543_),
    .A2(net536),
    .Y(_0415_),
    .B1(_1265_));
 sg13g2_o21ai_1 _3382_ (.B1(net558),
    .Y(_1266_),
    .A1(net632),
    .A2(net536));
 sg13g2_a21oi_1 _3383_ (.A1(_0542_),
    .A2(net536),
    .Y(_0416_),
    .B1(_1266_));
 sg13g2_nand2_1 _3384_ (.Y(_1267_),
    .A(_0809_),
    .B(_0815_));
 sg13g2_o21ai_1 _3385_ (.B1(_0815_),
    .Y(_1268_),
    .A1(_0087_),
    .A2(_0809_));
 sg13g2_o21ai_1 _3386_ (.B1(net558),
    .Y(_1269_),
    .A1(net536),
    .A2(_1268_));
 sg13g2_nor2_1 _3387_ (.A(_0816_),
    .B(_1269_),
    .Y(_1270_));
 sg13g2_nor2_1 _3388_ (.A(_0608_),
    .B(net533),
    .Y(_1271_));
 sg13g2_a21oi_1 _3389_ (.A1(net861),
    .A2(net533),
    .Y(_1272_),
    .B1(_1271_));
 sg13g2_nor2_1 _3390_ (.A(net1082),
    .B(net459),
    .Y(_1273_));
 sg13g2_a21oi_1 _3391_ (.A1(net459),
    .A2(_1272_),
    .Y(_0417_),
    .B1(_1273_));
 sg13g2_and2_1 _3392_ (.A(\dut.xfer.next_obuffer[2] ),
    .B(_0828_),
    .X(_1274_));
 sg13g2_a21oi_1 _3393_ (.A1(\dut.din_data[2] ),
    .A2(net535),
    .Y(_1275_),
    .B1(_1274_));
 sg13g2_nor2_1 _3394_ (.A(net987),
    .B(net459),
    .Y(_1276_));
 sg13g2_a21oi_1 _3395_ (.A1(net459),
    .A2(_1275_),
    .Y(_0418_),
    .B1(_1276_));
 sg13g2_and2_1 _3396_ (.A(\dut.xfer.next_obuffer[3] ),
    .B(_0828_),
    .X(_1277_));
 sg13g2_a21oi_1 _3397_ (.A1(\dut.din_data[3] ),
    .A2(net534),
    .Y(_1278_),
    .B1(_1277_));
 sg13g2_nor2_1 _3398_ (.A(net822),
    .B(net458),
    .Y(_1279_));
 sg13g2_a21oi_1 _3399_ (.A1(net458),
    .A2(_1278_),
    .Y(_0419_),
    .B1(_1279_));
 sg13g2_and2_1 _3400_ (.A(net822),
    .B(net532),
    .X(_1280_));
 sg13g2_a21oi_1 _3401_ (.A1(\dut.din_data[4] ),
    .A2(net534),
    .Y(_1281_),
    .B1(_1280_));
 sg13g2_nor2_1 _3402_ (.A(net1055),
    .B(net458),
    .Y(_1282_));
 sg13g2_a21oi_1 _3403_ (.A1(net458),
    .A2(_1281_),
    .Y(_0420_),
    .B1(_1282_));
 sg13g2_and2_1 _3404_ (.A(\dut.xfer.next_obuffer[5] ),
    .B(net532),
    .X(_1283_));
 sg13g2_a21oi_1 _3405_ (.A1(\dut.din_data[5] ),
    .A2(net534),
    .Y(_1284_),
    .B1(_1283_));
 sg13g2_nor2_1 _3406_ (.A(net879),
    .B(net458),
    .Y(_1285_));
 sg13g2_a21oi_1 _3407_ (.A1(net458),
    .A2(_1284_),
    .Y(_0421_),
    .B1(_1285_));
 sg13g2_and2_1 _3408_ (.A(net879),
    .B(net532),
    .X(_1286_));
 sg13g2_a21oi_1 _3409_ (.A1(net881),
    .A2(net534),
    .Y(_1287_),
    .B1(_1286_));
 sg13g2_nor2_1 _3410_ (.A(net1078),
    .B(net458),
    .Y(_1288_));
 sg13g2_a21oi_1 _3411_ (.A1(net458),
    .A2(_1287_),
    .Y(_0422_),
    .B1(_1288_));
 sg13g2_and2_1 _3412_ (.A(\dut.xfer.next_obuffer[7] ),
    .B(net532),
    .X(_1289_));
 sg13g2_a21oi_1 _3413_ (.A1(\dut.din_data[7] ),
    .A2(net534),
    .Y(_1290_),
    .B1(_1289_));
 sg13g2_nor2_1 _3414_ (.A(net877),
    .B(net459),
    .Y(_1291_));
 sg13g2_a21oi_1 _3415_ (.A1(net459),
    .A2(_1290_),
    .Y(_0423_),
    .B1(_1291_));
 sg13g2_o21ai_1 _3416_ (.B1(net861),
    .Y(_1292_),
    .A1(_0816_),
    .A2(_1269_));
 sg13g2_o21ai_1 _3417_ (.B1(_1292_),
    .Y(_0424_),
    .A1(_0550_),
    .A2(net533));
 sg13g2_nor2_1 _3418_ (.A(\dut.dout_tag[0] ),
    .B(net1022),
    .Y(_1293_));
 sg13g2_nand3_1 _3419_ (.B(_0825_),
    .C(_1293_),
    .A(\dut.dout_tag[2] ),
    .Y(_1294_));
 sg13g2_or2_1 _3420_ (.X(_1295_),
    .B(_1294_),
    .A(_0617_));
 sg13g2_nor2_1 _3421_ (.A(net566),
    .B(_0660_),
    .Y(_1296_));
 sg13g2_a21oi_1 _3422_ (.A1(net566),
    .A2(_0021_),
    .Y(_1297_),
    .B1(_1296_));
 sg13g2_nand2_1 _3423_ (.Y(_1298_),
    .A(net1315),
    .B(net450));
 sg13g2_o21ai_1 _3424_ (.B1(_1298_),
    .Y(_0425_),
    .A1(net450),
    .A2(_1297_));
 sg13g2_nor2_1 _3425_ (.A(net566),
    .B(_0653_),
    .Y(_1299_));
 sg13g2_a21oi_1 _3426_ (.A1(net566),
    .A2(_0782_),
    .Y(_1300_),
    .B1(_1299_));
 sg13g2_nand2_1 _3427_ (.Y(_1301_),
    .A(net568),
    .B(net450));
 sg13g2_o21ai_1 _3428_ (.B1(_1301_),
    .Y(_0426_),
    .A1(net450),
    .A2(_1300_));
 sg13g2_nand2_1 _3429_ (.Y(_1302_),
    .A(net884),
    .B(net449));
 sg13g2_nor2_1 _3430_ (.A(net565),
    .B(_0680_),
    .Y(_1303_));
 sg13g2_a21oi_1 _3431_ (.A1(net566),
    .A2(_0786_),
    .Y(_1304_),
    .B1(_1303_));
 sg13g2_o21ai_1 _3432_ (.B1(_1302_),
    .Y(_0427_),
    .A1(net449),
    .A2(_1304_));
 sg13g2_nand2_1 _3433_ (.Y(_1305_),
    .A(net921),
    .B(net449));
 sg13g2_mux2_1 _3434_ (.A0(_0656_),
    .A1(_0785_),
    .S(net565),
    .X(_1306_));
 sg13g2_o21ai_1 _3435_ (.B1(_1305_),
    .Y(_0428_),
    .A1(net449),
    .A2(_1306_));
 sg13g2_nand2_1 _3436_ (.Y(_1307_),
    .A(net565),
    .B(_0779_));
 sg13g2_o21ai_1 _3437_ (.B1(_1307_),
    .Y(_1308_),
    .A1(net565),
    .A2(_0663_));
 sg13g2_nand2_1 _3438_ (.Y(_1309_),
    .A(net1119),
    .B(net449));
 sg13g2_o21ai_1 _3439_ (.B1(_1309_),
    .Y(_0429_),
    .A1(net449),
    .A2(_1308_));
 sg13g2_mux2_1 _3440_ (.A0(_0649_),
    .A1(_0762_),
    .S(net565),
    .X(_1310_));
 sg13g2_nand2_1 _3441_ (.Y(_1311_),
    .A(net971),
    .B(net449));
 sg13g2_o21ai_1 _3442_ (.B1(_1311_),
    .Y(_0430_),
    .A1(net449),
    .A2(_1310_));
 sg13g2_nand2_1 _3443_ (.Y(_1312_),
    .A(net564),
    .B(_0764_));
 sg13g2_o21ai_1 _3444_ (.B1(_1312_),
    .Y(_1313_),
    .A1(net564),
    .A2(_0688_));
 sg13g2_nand2_1 _3445_ (.Y(_1314_),
    .A(net839),
    .B(net448));
 sg13g2_o21ai_1 _3446_ (.B1(_1314_),
    .Y(_0431_),
    .A1(net448),
    .A2(_1313_));
 sg13g2_xor2_1 _3447_ (.B(_0758_),
    .A(_0041_),
    .X(_1315_));
 sg13g2_nand2_1 _3448_ (.Y(_1316_),
    .A(net564),
    .B(_1315_));
 sg13g2_o21ai_1 _3449_ (.B1(_1316_),
    .Y(_1317_),
    .A1(net564),
    .A2(_0707_));
 sg13g2_nand2_1 _3450_ (.Y(_1318_),
    .A(net845),
    .B(net448));
 sg13g2_o21ai_1 _3451_ (.B1(_1318_),
    .Y(_0432_),
    .A1(net448),
    .A2(_1317_));
 sg13g2_nor2b_1 _3452_ (.A(_0737_),
    .B_N(_0044_),
    .Y(_1319_));
 sg13g2_o21ai_1 _3453_ (.B1(net564),
    .Y(_1320_),
    .A1(_0773_),
    .A2(_1319_));
 sg13g2_o21ai_1 _3454_ (.B1(_1320_),
    .Y(_1321_),
    .A1(net564),
    .A2(_0669_));
 sg13g2_nand2_1 _3455_ (.Y(_1322_),
    .A(net725),
    .B(net448));
 sg13g2_o21ai_1 _3456_ (.B1(_1322_),
    .Y(_0433_),
    .A1(net457),
    .A2(_1321_));
 sg13g2_xor2_1 _3457_ (.B(_0773_),
    .A(_0047_),
    .X(_1323_));
 sg13g2_nand2_1 _3458_ (.Y(_1324_),
    .A(net564),
    .B(_1323_));
 sg13g2_o21ai_1 _3459_ (.B1(_1324_),
    .Y(_1325_),
    .A1(net564),
    .A2(_0675_));
 sg13g2_nand2_1 _3460_ (.Y(_1326_),
    .A(net740),
    .B(net448));
 sg13g2_o21ai_1 _3461_ (.B1(_1326_),
    .Y(_0434_),
    .A1(net448),
    .A2(_1325_));
 sg13g2_and2_1 _3462_ (.A(_0050_),
    .B(_0741_),
    .X(_1327_));
 sg13g2_o21ai_1 _3463_ (.B1(net560),
    .Y(_1328_),
    .A1(_0760_),
    .A2(_1327_));
 sg13g2_o21ai_1 _3464_ (.B1(_1328_),
    .Y(_1329_),
    .A1(net560),
    .A2(_0694_));
 sg13g2_nand2_1 _3465_ (.Y(_1330_),
    .A(net767),
    .B(net447));
 sg13g2_o21ai_1 _3466_ (.B1(_1330_),
    .Y(_0435_),
    .A1(net447),
    .A2(_1329_));
 sg13g2_xor2_1 _3467_ (.B(_0760_),
    .A(_0053_),
    .X(_1331_));
 sg13g2_nand2_1 _3468_ (.Y(_1332_),
    .A(net560),
    .B(_1331_));
 sg13g2_o21ai_1 _3469_ (.B1(_1332_),
    .Y(_1333_),
    .A1(net560),
    .A2(_0691_));
 sg13g2_nand2_1 _3470_ (.Y(_1334_),
    .A(net898),
    .B(net444));
 sg13g2_o21ai_1 _3471_ (.B1(_1334_),
    .Y(_0436_),
    .A1(net444),
    .A2(_1333_));
 sg13g2_nand2_1 _3472_ (.Y(_1335_),
    .A(_0056_),
    .B(_0744_));
 sg13g2_nand3_1 _3473_ (.B(_0776_),
    .C(_1335_),
    .A(net559),
    .Y(_1336_));
 sg13g2_o21ai_1 _3474_ (.B1(_1336_),
    .Y(_1337_),
    .A1(net559),
    .A2(_0626_));
 sg13g2_mux2_1 _3475_ (.A0(_1337_),
    .A1(net1224),
    .S(net447),
    .X(_0437_));
 sg13g2_nor2_1 _3476_ (.A(net559),
    .B(_0636_),
    .Y(_1338_));
 sg13g2_xor2_1 _3477_ (.B(_0776_),
    .A(_0059_),
    .X(_1339_));
 sg13g2_a21oi_1 _3478_ (.A1(net559),
    .A2(_1339_),
    .Y(_1340_),
    .B1(_1338_));
 sg13g2_nand2_1 _3479_ (.Y(_1341_),
    .A(net709),
    .B(net444));
 sg13g2_o21ai_1 _3480_ (.B1(_1341_),
    .Y(_0438_),
    .A1(net444),
    .A2(_1340_));
 sg13g2_nand2_1 _3481_ (.Y(_1342_),
    .A(net769),
    .B(net444));
 sg13g2_nor2b_1 _3482_ (.A(_0746_),
    .B_N(_0062_),
    .Y(_1343_));
 sg13g2_o21ai_1 _3483_ (.B1(net559),
    .Y(_1344_),
    .A1(_0756_),
    .A2(_1343_));
 sg13g2_o21ai_1 _3484_ (.B1(_1344_),
    .Y(_1345_),
    .A1(net559),
    .A2(_0634_));
 sg13g2_o21ai_1 _3485_ (.B1(_1342_),
    .Y(_0439_),
    .A1(net444),
    .A2(_1345_));
 sg13g2_nor2_1 _3486_ (.A(net559),
    .B(_0646_),
    .Y(_1346_));
 sg13g2_xnor2_1 _3487_ (.Y(_1347_),
    .A(_0065_),
    .B(_0756_));
 sg13g2_a21oi_1 _3488_ (.A1(net559),
    .A2(_1347_),
    .Y(_1348_),
    .B1(_1346_));
 sg13g2_nand2_1 _3489_ (.Y(_1349_),
    .A(net755),
    .B(net444));
 sg13g2_o21ai_1 _3490_ (.B1(_1349_),
    .Y(_0440_),
    .A1(net444),
    .A2(_1348_));
 sg13g2_and2_1 _3491_ (.A(_0068_),
    .B(_0748_),
    .X(_1350_));
 sg13g2_o21ai_1 _3492_ (.B1(net561),
    .Y(_1351_),
    .A1(_0771_),
    .A2(_1350_));
 sg13g2_o21ai_1 _3493_ (.B1(_1351_),
    .Y(_1352_),
    .A1(net561),
    .A2(_0644_));
 sg13g2_nand2_1 _3494_ (.Y(_1353_),
    .A(net841),
    .B(net445));
 sg13g2_o21ai_1 _3495_ (.B1(_1353_),
    .Y(_0441_),
    .A1(net445),
    .A2(_1352_));
 sg13g2_xnor2_1 _3496_ (.Y(_1354_),
    .A(_0071_),
    .B(_0771_));
 sg13g2_nor2_1 _3497_ (.A(net561),
    .B(_0685_),
    .Y(_1355_));
 sg13g2_a21oi_1 _3498_ (.A1(net561),
    .A2(_1354_),
    .Y(_1356_),
    .B1(_1355_));
 sg13g2_nand2_1 _3499_ (.Y(_1357_),
    .A(net843),
    .B(net445));
 sg13g2_o21ai_1 _3500_ (.B1(_1357_),
    .Y(_0442_),
    .A1(net445),
    .A2(_1356_));
 sg13g2_xor2_1 _3501_ (.B(_0750_),
    .A(_0074_),
    .X(_1358_));
 sg13g2_mux2_1 _3502_ (.A0(_0697_),
    .A1(_1358_),
    .S(net561),
    .X(_1359_));
 sg13g2_nand2_1 _3503_ (.Y(_1360_),
    .A(net849),
    .B(net446));
 sg13g2_o21ai_1 _3504_ (.B1(_1360_),
    .Y(_0443_),
    .A1(net445),
    .A2(_1359_));
 sg13g2_nand2_1 _3505_ (.Y(_1361_),
    .A(net742),
    .B(net445));
 sg13g2_xnor2_1 _3506_ (.Y(_1362_),
    .A(_0077_),
    .B(_0755_));
 sg13g2_nor2b_1 _3507_ (.A(net561),
    .B_N(_0704_),
    .Y(_1363_));
 sg13g2_a21oi_1 _3508_ (.A1(net561),
    .A2(_1362_),
    .Y(_1364_),
    .B1(_1363_));
 sg13g2_o21ai_1 _3509_ (.B1(_1361_),
    .Y(_0444_),
    .A1(net445),
    .A2(_1364_));
 sg13g2_nor2b_1 _3510_ (.A(_0752_),
    .B_N(_0080_),
    .Y(_1365_));
 sg13g2_o21ai_1 _3511_ (.B1(net562),
    .Y(_1366_),
    .A1(_0766_),
    .A2(_1365_));
 sg13g2_o21ai_1 _3512_ (.B1(_1366_),
    .Y(_1367_),
    .A1(net562),
    .A2(_0700_));
 sg13g2_nand2_1 _3513_ (.Y(_1368_),
    .A(net815),
    .B(net446));
 sg13g2_o21ai_1 _3514_ (.B1(_1368_),
    .Y(_0445_),
    .A1(net446),
    .A2(_1367_));
 sg13g2_xor2_1 _3515_ (.B(_0766_),
    .A(_0083_),
    .X(_1369_));
 sg13g2_nand2_1 _3516_ (.Y(_1370_),
    .A(net715),
    .B(net446));
 sg13g2_nand2_1 _3517_ (.Y(_1371_),
    .A(net562),
    .B(_1369_));
 sg13g2_o21ai_1 _3518_ (.B1(_1371_),
    .Y(_1372_),
    .A1(net562),
    .A2(_0641_));
 sg13g2_o21ai_1 _3519_ (.B1(_1370_),
    .Y(_0446_),
    .A1(net446),
    .A2(_1372_));
 sg13g2_o21ai_1 _3520_ (.B1(_0903_),
    .Y(_1373_),
    .A1(\cpu.state.cnt_r[1] ),
    .A2(\cpu.state.cnt_r[0] ));
 sg13g2_mux2_1 _3521_ (.A0(_1373_),
    .A1(net545),
    .S(_0900_),
    .X(_1374_));
 sg13g2_nor2_1 _3522_ (.A(net1189),
    .B(_1374_),
    .Y(_1375_));
 sg13g2_a21oi_1 _3523_ (.A1(_0582_),
    .A2(_1374_),
    .Y(_0447_),
    .B1(_1375_));
 sg13g2_a21oi_1 _3524_ (.A1(net1289),
    .A2(_0900_),
    .Y(_1376_),
    .B1(_1374_));
 sg13g2_a22oi_1 _3525_ (.Y(_0448_),
    .B1(net1290),
    .B2(_1071_),
    .A2(_1374_),
    .A1(_0591_));
 sg13g2_a21oi_1 _3526_ (.A1(_0549_),
    .A2(net558),
    .Y(_0449_),
    .B1(net537));
 sg13g2_o21ai_1 _3527_ (.B1(_1267_),
    .Y(_1377_),
    .A1(net567),
    .A2(\dut.flash_csb ));
 sg13g2_o21ai_1 _3528_ (.B1(_1377_),
    .Y(_1378_),
    .A1(net567),
    .A2(_1267_));
 sg13g2_nor3_1 _3529_ (.A(net744),
    .B(net536),
    .C(_1378_),
    .Y(_0450_));
 sg13g2_o21ai_1 _3530_ (.B1(net558),
    .Y(_1379_),
    .A1(net1329),
    .A2(_0815_));
 sg13g2_o21ai_1 _3531_ (.B1(net533),
    .Y(_0451_),
    .A1(_0818_),
    .A2(net1330));
 sg13g2_a21oi_2 _3532_ (.B1(net537),
    .Y(_1380_),
    .A2(_0816_),
    .A1(net558));
 sg13g2_nand2b_1 _3533_ (.Y(_1381_),
    .B(net567),
    .A_N(\dut.xfer.dummy_count[0] ));
 sg13g2_nand2_1 _3534_ (.Y(_1382_),
    .A(\dut.xfer.dummy_count[0] ),
    .B(_0548_));
 sg13g2_a21o_1 _3535_ (.A2(_1382_),
    .A1(_1381_),
    .B1(net534),
    .X(_1383_));
 sg13g2_nand3_1 _3536_ (.B(net1203),
    .C(net535),
    .A(net1220),
    .Y(_1384_));
 sg13g2_a21oi_1 _3537_ (.A1(_1383_),
    .A2(_1384_),
    .Y(_0452_),
    .B1(_1380_));
 sg13g2_xnor2_1 _3538_ (.Y(_1385_),
    .A(net1247),
    .B(_1381_));
 sg13g2_nand2_1 _3539_ (.Y(_1386_),
    .A(net533),
    .B(_1385_));
 sg13g2_nand3_1 _3540_ (.B(net1172),
    .C(net535),
    .A(net1220),
    .Y(_1387_));
 sg13g2_a21oi_1 _3541_ (.A1(_1386_),
    .A2(_1387_),
    .Y(_0453_),
    .B1(_1380_));
 sg13g2_or3_1 _3542_ (.A(\dut.xfer.dummy_count[2] ),
    .B(\dut.xfer.dummy_count[1] ),
    .C(_1381_),
    .X(_1388_));
 sg13g2_o21ai_1 _3543_ (.B1(net1274),
    .Y(_1389_),
    .A1(\dut.xfer.dummy_count[1] ),
    .A2(_1381_));
 sg13g2_a21o_1 _3544_ (.A2(_1389_),
    .A1(_1388_),
    .B1(net534),
    .X(_1390_));
 sg13g2_nand3_1 _3545_ (.B(net1267),
    .C(net535),
    .A(net1220),
    .Y(_1391_));
 sg13g2_a21oi_1 _3546_ (.A1(net1275),
    .A2(_1391_),
    .Y(_0454_),
    .B1(_1380_));
 sg13g2_a22oi_1 _3547_ (.Y(_1392_),
    .B1(_1388_),
    .B2(net1241),
    .A2(_0815_),
    .A1(net567));
 sg13g2_or2_1 _3548_ (.X(_1393_),
    .B(_1392_),
    .A(net534));
 sg13g2_nand3_1 _3549_ (.B(net1167),
    .C(net535),
    .A(net1220),
    .Y(_1394_));
 sg13g2_a21oi_1 _3550_ (.A1(_1393_),
    .A2(_1394_),
    .Y(_0455_),
    .B1(_1380_));
 sg13g2_and3_2 _3551_ (.X(_1395_),
    .A(\dut.xfer.resetn ),
    .B(_0087_),
    .C(_1008_));
 sg13g2_mux2_1 _3552_ (.A0(net801),
    .A1(net1),
    .S(_1395_),
    .X(_0456_));
 sg13g2_mux2_1 _3553_ (.A0(net947),
    .A1(net801),
    .S(_1395_),
    .X(_0457_));
 sg13g2_mux2_1 _3554_ (.A0(net1114),
    .A1(net947),
    .S(_1395_),
    .X(_0458_));
 sg13g2_mux2_1 _3555_ (.A0(net1081),
    .A1(net1114),
    .S(_1395_),
    .X(_0459_));
 sg13g2_mux2_1 _3556_ (.A0(net788),
    .A1(net1081),
    .S(_1395_),
    .X(_0460_));
 sg13g2_mux2_1 _3557_ (.A0(net749),
    .A1(net788),
    .S(_1395_),
    .X(_0461_));
 sg13g2_mux2_1 _3558_ (.A0(net1125),
    .A1(net749),
    .S(_1395_),
    .X(_0462_));
 sg13g2_mux2_1 _3559_ (.A0(net1015),
    .A1(net1125),
    .S(_1395_),
    .X(_0463_));
 sg13g2_nand2b_1 _3560_ (.Y(_0464_),
    .B(net558),
    .A_N(_0823_));
 sg13g2_nand2b_1 _3561_ (.Y(_1396_),
    .B(net445),
    .A_N(net561));
 sg13g2_and2_1 _3562_ (.A(_0841_),
    .B(_1396_),
    .X(_0466_));
 sg13g2_nor2_2 _3563_ (.A(net566),
    .B(net450),
    .Y(_1397_));
 sg13g2_a221oi_1 _3564_ (.B2(_0573_),
    .C1(_1397_),
    .B1(net450),
    .A1(_0616_),
    .Y(_0467_),
    .A2(_0625_));
 sg13g2_a21oi_1 _3565_ (.A1(_0546_),
    .A2(_1294_),
    .Y(_0468_),
    .B1(_0808_));
 sg13g2_nand2b_1 _3566_ (.Y(_1398_),
    .B(\dut.dout_tag[0] ),
    .A_N(\dut.dout_tag[2] ));
 sg13g2_nand3_1 _3567_ (.B(_0616_),
    .C(_0825_),
    .A(\dut.dout_tag[1] ),
    .Y(_1399_));
 sg13g2_or2_2 _3568_ (.X(_1400_),
    .B(_1399_),
    .A(_1398_));
 sg13g2_mux2_1 _3569_ (.A0(net801),
    .A1(net906),
    .S(_1400_),
    .X(_0469_));
 sg13g2_mux2_1 _3570_ (.A0(net947),
    .A1(net937),
    .S(_1400_),
    .X(_0470_));
 sg13g2_mux2_1 _3571_ (.A0(\dut.dout_data[2] ),
    .A1(net983),
    .S(_1400_),
    .X(_0471_));
 sg13g2_mux2_1 _3572_ (.A0(net1081),
    .A1(net1153),
    .S(_1400_),
    .X(_0472_));
 sg13g2_mux2_1 _3573_ (.A0(net788),
    .A1(net900),
    .S(_1400_),
    .X(_0473_));
 sg13g2_mux2_1 _3574_ (.A0(net749),
    .A1(net1100),
    .S(_1400_),
    .X(_0474_));
 sg13g2_mux2_1 _3575_ (.A0(net1125),
    .A1(net1096),
    .S(_1400_),
    .X(_0475_));
 sg13g2_mux2_1 _3576_ (.A0(net1015),
    .A1(net1009),
    .S(_1400_),
    .X(_0476_));
 sg13g2_nand2_1 _3577_ (.Y(_1401_),
    .A(net1278),
    .B(net441));
 sg13g2_o21ai_1 _3578_ (.B1(_1401_),
    .Y(_0477_),
    .A1(_0545_),
    .A2(_0808_));
 sg13g2_nand2_1 _3579_ (.Y(_1402_),
    .A(_0569_),
    .B(_0571_));
 sg13g2_a21oi_1 _3580_ (.A1(_0825_),
    .A2(_1402_),
    .Y(_0478_),
    .B1(_0808_));
 sg13g2_mux2_1 _3581_ (.A0(net873),
    .A1(\cpu.bufreg2.i_dat[0] ),
    .S(net451),
    .X(_0479_));
 sg13g2_mux2_1 _3582_ (.A0(net1016),
    .A1(\cpu.bufreg2.i_dat[1] ),
    .S(net451),
    .X(_0480_));
 sg13g2_mux2_1 _3583_ (.A0(net835),
    .A1(\cpu.bufreg2.i_dat[2] ),
    .S(net452),
    .X(_0481_));
 sg13g2_mux2_1 _3584_ (.A0(net837),
    .A1(\cpu.bufreg2.i_dat[3] ),
    .S(net452),
    .X(_0482_));
 sg13g2_mux2_1 _3585_ (.A0(net989),
    .A1(\cpu.bufreg2.i_dat[4] ),
    .S(net451),
    .X(_0483_));
 sg13g2_nor2_1 _3586_ (.A(net736),
    .B(net451),
    .Y(_1403_));
 sg13g2_a21oi_1 _3587_ (.A1(_0595_),
    .A2(net451),
    .Y(_0484_),
    .B1(_1403_));
 sg13g2_mux2_1 _3588_ (.A0(net1033),
    .A1(\cpu.bufreg2.i_dat[6] ),
    .S(net452),
    .X(_0485_));
 sg13g2_mux2_1 _3589_ (.A0(net927),
    .A1(\cpu.bufreg2.i_dat[7] ),
    .S(net452),
    .X(_0486_));
 sg13g2_mux2_1 _3590_ (.A0(net654),
    .A1(\cpu.bufreg2.i_dat[8] ),
    .S(net454),
    .X(_0487_));
 sg13g2_mux2_1 _3591_ (.A0(net894),
    .A1(\cpu.bufreg2.i_dat[9] ),
    .S(net456),
    .X(_0488_));
 sg13g2_mux2_1 _3592_ (.A0(net782),
    .A1(net851),
    .S(net455),
    .X(_0489_));
 sg13g2_mux2_1 _3593_ (.A0(net753),
    .A1(net789),
    .S(net454),
    .X(_0490_));
 sg13g2_mux2_1 _3594_ (.A0(net763),
    .A1(\cpu.bufreg2.i_dat[12] ),
    .S(net455),
    .X(_0491_));
 sg13g2_mux2_1 _3595_ (.A0(net747),
    .A1(\cpu.bufreg2.i_dat[13] ),
    .S(net453),
    .X(_0492_));
 sg13g2_mux2_1 _3596_ (.A0(net820),
    .A1(net829),
    .S(net453),
    .X(_0493_));
 sg13g2_mux2_1 _3597_ (.A0(net761),
    .A1(net772),
    .S(net455),
    .X(_0494_));
 sg13g2_mux2_1 _3598_ (.A0(net906),
    .A1(\cpu.bufreg2.i_dat[16] ),
    .S(net456),
    .X(_0495_));
 sg13g2_mux2_1 _3599_ (.A0(net937),
    .A1(\cpu.bufreg2.i_dat[17] ),
    .S(net455),
    .X(_0496_));
 sg13g2_mux2_1 _3600_ (.A0(net983),
    .A1(net1046),
    .S(net455),
    .X(_0497_));
 sg13g2_mux2_1 _3601_ (.A0(net1153),
    .A1(net1116),
    .S(net455),
    .X(_0498_));
 sg13g2_mux2_1 _3602_ (.A0(net900),
    .A1(\cpu.bufreg2.i_dat[20] ),
    .S(net454),
    .X(_0499_));
 sg13g2_mux2_1 _3603_ (.A0(net1100),
    .A1(\cpu.bufreg2.i_dat[21] ),
    .S(net454),
    .X(_0500_));
 sg13g2_mux2_1 _3604_ (.A0(net1096),
    .A1(\cpu.bufreg2.i_dat[22] ),
    .S(net453),
    .X(_0501_));
 sg13g2_mux2_1 _3605_ (.A0(net1009),
    .A1(\cpu.bufreg2.i_dat[23] ),
    .S(net454),
    .X(_0502_));
 sg13g2_mux2_1 _3606_ (.A0(net801),
    .A1(net1277),
    .S(net454),
    .X(_0503_));
 sg13g2_mux2_1 _3607_ (.A0(net947),
    .A1(net1256),
    .S(net454),
    .X(_0504_));
 sg13g2_mux2_1 _3608_ (.A0(net1114),
    .A1(net1270),
    .S(net454),
    .X(_0505_));
 sg13g2_mux2_1 _3609_ (.A0(net1081),
    .A1(net1263),
    .S(net452),
    .X(_0506_));
 sg13g2_mux2_1 _3610_ (.A0(net788),
    .A1(net1264),
    .S(net452),
    .X(_0507_));
 sg13g2_mux2_1 _3611_ (.A0(net749),
    .A1(net1261),
    .S(net452),
    .X(_0508_));
 sg13g2_mux2_1 _3612_ (.A0(net1125),
    .A1(net1236),
    .S(net452),
    .X(_0509_));
 sg13g2_mux2_1 _3613_ (.A0(net1015),
    .A1(net1262),
    .S(net453),
    .X(_0510_));
 sg13g2_o21ai_1 _3614_ (.B1(net524),
    .Y(_1404_),
    .A1(_0879_),
    .A2(net483));
 sg13g2_o21ai_1 _3615_ (.B1(_1404_),
    .Y(_1405_),
    .A1(net557),
    .A2(_1247_));
 sg13g2_inv_1 _3616_ (.Y(_0511_),
    .A(_1405_));
 sg13g2_nor3_1 _3617_ (.A(\dut.state[0] ),
    .B(\dut.state[1] ),
    .C(\dut.state[12] ),
    .Y(_1406_));
 sg13g2_and3_1 _3618_ (.X(_1407_),
    .A(_0570_),
    .B(_0572_),
    .C(_1406_));
 sg13g2_nor4_1 _3619_ (.A(\dut.state[4] ),
    .B(\dut.state[2] ),
    .C(\dut.state[6] ),
    .D(\dut.state[5] ),
    .Y(_1408_));
 sg13g2_and2_1 _3620_ (.A(_0562_),
    .B(_1408_),
    .X(_1409_));
 sg13g2_nand3b_1 _3621_ (.B(_1407_),
    .C(_1409_),
    .Y(_1410_),
    .A_N(net1246));
 sg13g2_nand3_1 _3622_ (.B(_0852_),
    .C(_1410_),
    .A(_0836_),
    .Y(_1411_));
 sg13g2_and2_1 _3623_ (.A(_0544_),
    .B(_1411_),
    .X(_1412_));
 sg13g2_nor3_1 _3624_ (.A(net1237),
    .B(net854),
    .C(_1411_),
    .Y(_1413_));
 sg13g2_nor3_1 _3625_ (.A(_0617_),
    .B(_1412_),
    .C(_1413_),
    .Y(_0512_));
 sg13g2_nor3_1 _3626_ (.A(net1178),
    .B(net1237),
    .C(_1411_),
    .Y(_1414_));
 sg13g2_a21oi_1 _3627_ (.A1(_0543_),
    .A2(_1411_),
    .Y(_1415_),
    .B1(_0617_));
 sg13g2_nor2b_1 _3628_ (.A(_1414_),
    .B_N(_1415_),
    .Y(_0513_));
 sg13g2_a22oi_1 _3629_ (.Y(_1416_),
    .B1(_1411_),
    .B2(net804),
    .A2(_0846_),
    .A1(_0836_));
 sg13g2_nor2_1 _3630_ (.A(_0617_),
    .B(net805),
    .Y(_0514_));
 sg13g2_nor3_1 _3631_ (.A(\dut.dout_tag[1] ),
    .B(_0617_),
    .C(_1398_),
    .Y(_1417_));
 sg13g2_nand2_2 _3632_ (.Y(_1418_),
    .A(_0825_),
    .B(_1417_));
 sg13g2_mux2_1 _3633_ (.A0(net801),
    .A1(net873),
    .S(_1418_),
    .X(_0515_));
 sg13g2_mux2_1 _3634_ (.A0(net947),
    .A1(net1016),
    .S(_1418_),
    .X(_0516_));
 sg13g2_mux2_1 _3635_ (.A0(net1114),
    .A1(net835),
    .S(_1418_),
    .X(_0517_));
 sg13g2_mux2_1 _3636_ (.A0(net1081),
    .A1(net837),
    .S(_1418_),
    .X(_0518_));
 sg13g2_mux2_1 _3637_ (.A0(net788),
    .A1(net989),
    .S(_1418_),
    .X(_0519_));
 sg13g2_mux2_1 _3638_ (.A0(net749),
    .A1(net736),
    .S(_1418_),
    .X(_0520_));
 sg13g2_mux2_1 _3639_ (.A0(net1125),
    .A1(net1033),
    .S(_1418_),
    .X(_0521_));
 sg13g2_mux2_1 _3640_ (.A0(net1015),
    .A1(net927),
    .S(_1418_),
    .X(_0522_));
 sg13g2_nor2_1 _3641_ (.A(net1032),
    .B(_1397_),
    .Y(_1419_));
 sg13g2_a21oi_1 _3642_ (.A1(_0630_),
    .A2(_1397_),
    .Y(_0523_),
    .B1(_1419_));
 sg13g2_nor2_1 _3643_ (.A(net1195),
    .B(_1397_),
    .Y(_1420_));
 sg13g2_a21oi_1 _3644_ (.A1(_0628_),
    .A2(_1397_),
    .Y(_0524_),
    .B1(_1420_));
 sg13g2_nor3_2 _3645_ (.A(\dut.dout_tag[0] ),
    .B(\dut.dout_tag[2] ),
    .C(_1399_),
    .Y(_1421_));
 sg13g2_mux2_1 _3646_ (.A0(net654),
    .A1(net801),
    .S(_1421_),
    .X(_0525_));
 sg13g2_mux2_1 _3647_ (.A0(net894),
    .A1(net947),
    .S(_1421_),
    .X(_0526_));
 sg13g2_mux2_1 _3648_ (.A0(net782),
    .A1(\dut.dout_data[2] ),
    .S(_1421_),
    .X(_0527_));
 sg13g2_mux2_1 _3649_ (.A0(net753),
    .A1(\dut.dout_data[3] ),
    .S(_1421_),
    .X(_0528_));
 sg13g2_mux2_1 _3650_ (.A0(net763),
    .A1(net788),
    .S(_1421_),
    .X(_0529_));
 sg13g2_mux2_1 _3651_ (.A0(net747),
    .A1(net749),
    .S(_1421_),
    .X(_0530_));
 sg13g2_mux2_1 _3652_ (.A0(net820),
    .A1(\dut.dout_data[6] ),
    .S(_1421_),
    .X(_0531_));
 sg13g2_mux2_1 _3653_ (.A0(net761),
    .A1(\dut.dout_data[7] ),
    .S(_1421_),
    .X(_0532_));
 sg13g2_nand4_1 _3654_ (.B(_0845_),
    .C(_1407_),
    .A(_0726_),
    .Y(_1422_),
    .D(_1408_));
 sg13g2_and4_1 _3655_ (.A(_0616_),
    .B(net532),
    .C(_1410_),
    .D(_1422_),
    .X(_0533_));
 sg13g2_a21oi_1 _3656_ (.A1(_1406_),
    .A2(_1409_),
    .Y(_1423_),
    .B1(_0617_));
 sg13g2_nand2_1 _3657_ (.Y(_1424_),
    .A(_0836_),
    .B(_1423_));
 sg13g2_nor2b_2 _3658_ (.A(net443),
    .B_N(_0935_),
    .Y(_1425_));
 sg13g2_and2_1 _3659_ (.A(_0847_),
    .B(_1409_),
    .X(_1426_));
 sg13g2_or2_2 _3660_ (.X(_1427_),
    .B(_1426_),
    .A(\dut.state[4] ));
 sg13g2_a221oi_1 _3661_ (.B2(net578),
    .C1(_1427_),
    .B1(_0641_),
    .A1(net579),
    .Y(_1428_),
    .A2(_0637_));
 sg13g2_o21ai_1 _3662_ (.B1(_1428_),
    .Y(_1429_),
    .A1(_0649_),
    .A2(net521));
 sg13g2_inv_1 _3663_ (.Y(_1430_),
    .A(_1429_));
 sg13g2_a22oi_1 _3664_ (.Y(_0534_),
    .B1(_1425_),
    .B2(_1430_),
    .A2(net442),
    .A1(_0614_));
 sg13g2_nand2_1 _3665_ (.Y(_1431_),
    .A(net578),
    .B(_0700_));
 sg13g2_o21ai_1 _3666_ (.B1(_1431_),
    .Y(_1432_),
    .A1(_0560_),
    .A2(_0626_));
 sg13g2_o21ai_1 _3667_ (.B1(_0935_),
    .Y(_1433_),
    .A1(_0664_),
    .A2(net521));
 sg13g2_nor4_1 _3668_ (.A(net443),
    .B(_1426_),
    .C(_1432_),
    .D(_1433_),
    .Y(_1434_));
 sg13g2_a21oi_1 _3669_ (.A1(_0613_),
    .A2(net442),
    .Y(_0535_),
    .B1(_1434_));
 sg13g2_a221oi_1 _3670_ (.B2(net578),
    .C1(_1427_),
    .B1(_0704_),
    .A1(net579),
    .Y(_1435_),
    .A2(_0691_));
 sg13g2_o21ai_1 _3671_ (.B1(_1435_),
    .Y(_1436_),
    .A1(_0656_),
    .A2(net521));
 sg13g2_inv_1 _3672_ (.Y(_1437_),
    .A(_1436_));
 sg13g2_a22oi_1 _3673_ (.Y(_0536_),
    .B1(_1425_),
    .B2(_1437_),
    .A2(net442),
    .A1(_0612_));
 sg13g2_nor2_1 _3674_ (.A(_0680_),
    .B(net521),
    .Y(_1438_));
 sg13g2_nand2_1 _3675_ (.Y(_1439_),
    .A(net579),
    .B(_0694_));
 sg13g2_o21ai_1 _3676_ (.B1(_1439_),
    .Y(_1440_),
    .A1(_0562_),
    .A2(_0697_));
 sg13g2_nor3_2 _3677_ (.A(_1426_),
    .B(_1438_),
    .C(_1440_),
    .Y(_1441_));
 sg13g2_a22oi_1 _3678_ (.Y(_0537_),
    .B1(_1425_),
    .B2(_1441_),
    .A2(net442),
    .A1(_0611_));
 sg13g2_nor2_1 _3679_ (.A(_0653_),
    .B(net521),
    .Y(_1442_));
 sg13g2_a21oi_1 _3680_ (.A1(net579),
    .A2(_0675_),
    .Y(_1443_),
    .B1(\dut.state[1] ));
 sg13g2_o21ai_1 _3681_ (.B1(_1443_),
    .Y(_1444_),
    .A1(_0562_),
    .A2(_0685_));
 sg13g2_nor4_2 _3682_ (.A(net442),
    .B(_1427_),
    .C(_1442_),
    .Y(_1445_),
    .D(_1444_));
 sg13g2_a21oi_1 _3683_ (.A1(_0610_),
    .A2(net443),
    .Y(_0538_),
    .B1(_1445_));
 sg13g2_a221oi_1 _3684_ (.B2(net579),
    .C1(_1426_),
    .B1(_0669_),
    .A1(net578),
    .Y(_1446_),
    .A2(_0644_));
 sg13g2_o21ai_1 _3685_ (.B1(_1446_),
    .Y(_1447_),
    .A1(_0660_),
    .A2(net521));
 sg13g2_inv_1 _3686_ (.Y(_1448_),
    .A(_1447_));
 sg13g2_a22oi_1 _3687_ (.Y(_0539_),
    .B1(_1425_),
    .B2(_1448_),
    .A2(net442),
    .A1(_0609_));
 sg13g2_nor2_1 _3688_ (.A(_0628_),
    .B(net521),
    .Y(_1449_));
 sg13g2_nor2_1 _3689_ (.A(\dut.state[2] ),
    .B(_1427_),
    .Y(_1450_));
 sg13g2_a22oi_1 _3690_ (.Y(_1451_),
    .B1(_0707_),
    .B2(net579),
    .A2(_0647_),
    .A1(net578));
 sg13g2_nand3_1 _3691_ (.B(_1450_),
    .C(_1451_),
    .A(_0935_),
    .Y(_1452_));
 sg13g2_nor3_2 _3692_ (.A(net442),
    .B(_1449_),
    .C(_1452_),
    .Y(_1453_));
 sg13g2_a21oi_1 _3693_ (.A1(_0608_),
    .A2(net443),
    .Y(_0540_),
    .B1(_1453_));
 sg13g2_nor2_1 _3694_ (.A(_0630_),
    .B(net521),
    .Y(_1454_));
 sg13g2_a22oi_1 _3695_ (.Y(_1455_),
    .B1(_0688_),
    .B2(net579),
    .A2(_0634_),
    .A1(net578));
 sg13g2_nand3_1 _3696_ (.B(_1450_),
    .C(_1455_),
    .A(_0935_),
    .Y(_1456_));
 sg13g2_nor3_1 _3697_ (.A(net442),
    .B(_1454_),
    .C(_1456_),
    .Y(_1457_));
 sg13g2_a21oi_1 _3698_ (.A1(_0550_),
    .A2(net443),
    .Y(_0541_),
    .B1(_1457_));
 sg13g2_dfrbp_1 _3699_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net189),
    .D(_0094_),
    .Q_N(_1829_),
    .Q(\rf_shift_reg.rd_active ));
 sg13g2_dfrbp_1 _3700_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net419),
    .D(_0095_),
    .Q_N(_1828_),
    .Q(\rf_shift_reg.rreq_r ));
 sg13g2_dfrbp_1 _3701_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net418),
    .D(net647),
    .Q_N(_1827_),
    .Q(\rf_shift_reg.rdata[1] ));
 sg13g2_dfrbp_1 _3702_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net417),
    .D(_0097_),
    .Q_N(_1826_),
    .Q(\rf_shift_reg.x[1][1] ));
 sg13g2_dfrbp_1 _3703_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net416),
    .D(net1029),
    .Q_N(_1825_),
    .Q(\rf_shift_reg.x[1][2] ));
 sg13g2_dfrbp_1 _3704_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net415),
    .D(net641),
    .Q_N(_1824_),
    .Q(\rf_shift_reg.x[1][3] ));
 sg13g2_dfrbp_1 _3705_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net414),
    .D(_0100_),
    .Q_N(_1823_),
    .Q(\rf_shift_reg.x[1][4] ));
 sg13g2_dfrbp_1 _3706_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net413),
    .D(net926),
    .Q_N(_1822_),
    .Q(\rf_shift_reg.x[1][5] ));
 sg13g2_dfrbp_1 _3707_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net412),
    .D(net887),
    .Q_N(_1821_),
    .Q(\rf_shift_reg.x[1][6] ));
 sg13g2_dfrbp_1 _3708_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net411),
    .D(_0103_),
    .Q_N(_1820_),
    .Q(\rf_shift_reg.x[1][7] ));
 sg13g2_dfrbp_1 _3709_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net410),
    .D(net1014),
    .Q_N(_1819_),
    .Q(\rf_shift_reg.x[1][8] ));
 sg13g2_dfrbp_1 _3710_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net409),
    .D(_0105_),
    .Q_N(_1818_),
    .Q(\rf_shift_reg.x[1][9] ));
 sg13g2_dfrbp_1 _3711_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net408),
    .D(net915),
    .Q_N(_1817_),
    .Q(\rf_shift_reg.x[1][10] ));
 sg13g2_dfrbp_1 _3712_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net407),
    .D(_0107_),
    .Q_N(_1816_),
    .Q(\rf_shift_reg.x[1][11] ));
 sg13g2_dfrbp_1 _3713_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net406),
    .D(net1065),
    .Q_N(_1815_),
    .Q(\rf_shift_reg.x[1][12] ));
 sg13g2_dfrbp_1 _3714_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net405),
    .D(net868),
    .Q_N(_1814_),
    .Q(\rf_shift_reg.x[1][13] ));
 sg13g2_dfrbp_1 _3715_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net404),
    .D(_0110_),
    .Q_N(_1813_),
    .Q(\rf_shift_reg.x[1][14] ));
 sg13g2_dfrbp_1 _3716_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net403),
    .D(net950),
    .Q_N(_1812_),
    .Q(\rf_shift_reg.x[1][15] ));
 sg13g2_dfrbp_1 _3717_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net402),
    .D(_0112_),
    .Q_N(_1811_),
    .Q(\rf_shift_reg.x[1][16] ));
 sg13g2_dfrbp_1 _3718_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net401),
    .D(net958),
    .Q_N(_1810_),
    .Q(\rf_shift_reg.x[1][17] ));
 sg13g2_dfrbp_1 _3719_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net400),
    .D(_0114_),
    .Q_N(_1809_),
    .Q(\rf_shift_reg.x[1][18] ));
 sg13g2_dfrbp_1 _3720_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net396),
    .D(_0115_),
    .Q_N(_1808_),
    .Q(\rf_shift_reg.x[1][19] ));
 sg13g2_dfrbp_1 _3721_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net395),
    .D(_0116_),
    .Q_N(_1807_),
    .Q(\rf_shift_reg.x[1][20] ));
 sg13g2_dfrbp_1 _3722_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net394),
    .D(net911),
    .Q_N(_1806_),
    .Q(\rf_shift_reg.x[1][21] ));
 sg13g2_dfrbp_1 _3723_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net393),
    .D(net793),
    .Q_N(_1805_),
    .Q(\rf_shift_reg.x[1][22] ));
 sg13g2_dfrbp_1 _3724_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net392),
    .D(_0119_),
    .Q_N(_1804_),
    .Q(\rf_shift_reg.x[1][23] ));
 sg13g2_dfrbp_1 _3725_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net391),
    .D(net905),
    .Q_N(_1803_),
    .Q(\rf_shift_reg.x[1][24] ));
 sg13g2_dfrbp_1 _3726_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net390),
    .D(_0121_),
    .Q_N(_1802_),
    .Q(\rf_shift_reg.x[1][25] ));
 sg13g2_dfrbp_1 _3727_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net389),
    .D(net917),
    .Q_N(_1801_),
    .Q(\rf_shift_reg.x[1][26] ));
 sg13g2_dfrbp_1 _3728_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net388),
    .D(_0123_),
    .Q_N(_1800_),
    .Q(\rf_shift_reg.x[1][27] ));
 sg13g2_dfrbp_1 _3729_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net387),
    .D(net643),
    .Q_N(_1799_),
    .Q(\rf_shift_reg.x[1][28] ));
 sg13g2_dfrbp_1 _3730_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net386),
    .D(_0125_),
    .Q_N(_1798_),
    .Q(\rf_shift_reg.x[1][29] ));
 sg13g2_dfrbp_1 _3731_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net385),
    .D(net853),
    .Q_N(_1797_),
    .Q(\rf_shift_reg.x[1][30] ));
 sg13g2_dfrbp_1 _3732_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net384),
    .D(net1075),
    .Q_N(_1796_),
    .Q(\rf_shift_reg.x[1][31] ));
 sg13g2_dfrbp_1 _3733_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net383),
    .D(net637),
    .Q_N(_0093_),
    .Q(\rf_shift_reg.cnt[0] ));
 sg13g2_dfrbp_1 _3734_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net381),
    .D(net828),
    .Q_N(_1795_),
    .Q(\rf_shift_reg.cnt[1] ));
 sg13g2_dfrbp_1 _3735_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net379),
    .D(net1310),
    .Q_N(_1794_),
    .Q(\rf_shift_reg.cnt[2] ));
 sg13g2_dfrbp_1 _3736_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net377),
    .D(_0131_),
    .Q_N(_1793_),
    .Q(\rf_shift_reg.cnt[3] ));
 sg13g2_dfrbp_1 _3737_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net375),
    .D(net1139),
    .Q_N(_1792_),
    .Q(\rf_shift_reg.cnt[4] ));
 sg13g2_dfrbp_1 _3738_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net373),
    .D(net664),
    .Q_N(_1791_),
    .Q(\rf_shift_reg.rdata[2] ));
 sg13g2_dfrbp_1 _3739_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net372),
    .D(_0134_),
    .Q_N(_1790_),
    .Q(\rf_shift_reg.x[2][1] ));
 sg13g2_dfrbp_1 _3740_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net371),
    .D(net1008),
    .Q_N(_1789_),
    .Q(\rf_shift_reg.x[2][2] ));
 sg13g2_dfrbp_1 _3741_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net370),
    .D(net818),
    .Q_N(_1788_),
    .Q(\rf_shift_reg.x[2][3] ));
 sg13g2_dfrbp_1 _3742_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net369),
    .D(_0137_),
    .Q_N(_1787_),
    .Q(\rf_shift_reg.x[2][4] ));
 sg13g2_dfrbp_1 _3743_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net368),
    .D(net1019),
    .Q_N(_1786_),
    .Q(\rf_shift_reg.x[2][5] ));
 sg13g2_dfrbp_1 _3744_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net367),
    .D(_0139_),
    .Q_N(_1785_),
    .Q(\rf_shift_reg.x[2][6] ));
 sg13g2_dfrbp_1 _3745_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net366),
    .D(_0140_),
    .Q_N(_1784_),
    .Q(\rf_shift_reg.x[2][7] ));
 sg13g2_dfrbp_1 _3746_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net365),
    .D(net934),
    .Q_N(_1783_),
    .Q(\rf_shift_reg.x[2][8] ));
 sg13g2_dfrbp_1 _3747_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net364),
    .D(_0142_),
    .Q_N(_1782_),
    .Q(\rf_shift_reg.x[2][9] ));
 sg13g2_dfrbp_1 _3748_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net363),
    .D(_0143_),
    .Q_N(_1781_),
    .Q(\rf_shift_reg.x[2][10] ));
 sg13g2_dfrbp_1 _3749_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net362),
    .D(net982),
    .Q_N(_1780_),
    .Q(\rf_shift_reg.x[2][11] ));
 sg13g2_dfrbp_1 _3750_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net361),
    .D(_0145_),
    .Q_N(_1779_),
    .Q(\rf_shift_reg.x[2][12] ));
 sg13g2_dfrbp_1 _3751_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net360),
    .D(_0146_),
    .Q_N(_1778_),
    .Q(\rf_shift_reg.x[2][13] ));
 sg13g2_dfrbp_1 _3752_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net359),
    .D(net980),
    .Q_N(_1777_),
    .Q(\rf_shift_reg.x[2][14] ));
 sg13g2_dfrbp_1 _3753_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net358),
    .D(net864),
    .Q_N(_1776_),
    .Q(\rf_shift_reg.x[2][15] ));
 sg13g2_dfrbp_1 _3754_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net357),
    .D(_0149_),
    .Q_N(_1775_),
    .Q(\rf_shift_reg.x[2][16] ));
 sg13g2_dfrbp_1 _3755_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net356),
    .D(_0150_),
    .Q_N(_1774_),
    .Q(\rf_shift_reg.x[2][17] ));
 sg13g2_dfrbp_1 _3756_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net355),
    .D(_0151_),
    .Q_N(_1773_),
    .Q(\rf_shift_reg.x[2][18] ));
 sg13g2_dfrbp_1 _3757_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net354),
    .D(net913),
    .Q_N(_1772_),
    .Q(\rf_shift_reg.x[2][19] ));
 sg13g2_dfrbp_1 _3758_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net353),
    .D(_0153_),
    .Q_N(_1771_),
    .Q(\rf_shift_reg.x[2][20] ));
 sg13g2_dfrbp_1 _3759_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net352),
    .D(_0154_),
    .Q_N(_1770_),
    .Q(\rf_shift_reg.x[2][21] ));
 sg13g2_dfrbp_1 _3760_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net351),
    .D(net891),
    .Q_N(_1769_),
    .Q(\rf_shift_reg.x[2][22] ));
 sg13g2_dfrbp_1 _3761_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net350),
    .D(_0156_),
    .Q_N(_1768_),
    .Q(\rf_shift_reg.x[2][23] ));
 sg13g2_dfrbp_1 _3762_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net349),
    .D(_0157_),
    .Q_N(_1767_),
    .Q(\rf_shift_reg.x[2][24] ));
 sg13g2_dfrbp_1 _3763_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net348),
    .D(net1025),
    .Q_N(_1766_),
    .Q(\rf_shift_reg.x[2][25] ));
 sg13g2_dfrbp_1 _3764_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net347),
    .D(net1021),
    .Q_N(_1765_),
    .Q(\rf_shift_reg.x[2][26] ));
 sg13g2_dfrbp_1 _3765_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net346),
    .D(_0160_),
    .Q_N(_1764_),
    .Q(\rf_shift_reg.x[2][27] ));
 sg13g2_dfrbp_1 _3766_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net345),
    .D(net831),
    .Q_N(_1763_),
    .Q(\rf_shift_reg.x[2][28] ));
 sg13g2_dfrbp_1 _3767_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net344),
    .D(_0162_),
    .Q_N(_1762_),
    .Q(\rf_shift_reg.x[2][29] ));
 sg13g2_dfrbp_1 _3768_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net343),
    .D(net683),
    .Q_N(_1761_),
    .Q(\rf_shift_reg.x[2][30] ));
 sg13g2_dfrbp_1 _3769_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net342),
    .D(net1266),
    .Q_N(_1760_),
    .Q(\rf_shift_reg.x[2][31] ));
 sg13g2_dfrbp_1 _3770_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net341),
    .D(net645),
    .Q_N(_1759_),
    .Q(\rf_shift_reg.rdata[3] ));
 sg13g2_dfrbp_1 _3771_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net340),
    .D(_0166_),
    .Q_N(_1758_),
    .Q(\rf_shift_reg.x[3][1] ));
 sg13g2_dfrbp_1 _3772_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net339),
    .D(_0167_),
    .Q_N(_1757_),
    .Q(\rf_shift_reg.x[3][2] ));
 sg13g2_dfrbp_1 _3773_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net338),
    .D(_0168_),
    .Q_N(_1756_),
    .Q(\rf_shift_reg.x[3][3] ));
 sg13g2_dfrbp_1 _3774_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net337),
    .D(net1089),
    .Q_N(_1755_),
    .Q(\rf_shift_reg.x[3][4] ));
 sg13g2_dfrbp_1 _3775_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net336),
    .D(net954),
    .Q_N(_1754_),
    .Q(\rf_shift_reg.x[3][5] ));
 sg13g2_dfrbp_1 _3776_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net335),
    .D(_0171_),
    .Q_N(_1753_),
    .Q(\rf_shift_reg.x[3][6] ));
 sg13g2_dfrbp_1 _3777_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net334),
    .D(_0172_),
    .Q_N(_1752_),
    .Q(\rf_shift_reg.x[3][7] ));
 sg13g2_dfrbp_1 _3778_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net333),
    .D(net993),
    .Q_N(_1751_),
    .Q(\rf_shift_reg.x[3][8] ));
 sg13g2_dfrbp_1 _3779_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net332),
    .D(_0174_),
    .Q_N(_1750_),
    .Q(\rf_shift_reg.x[3][9] ));
 sg13g2_dfrbp_1 _3780_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net331),
    .D(net969),
    .Q_N(_1749_),
    .Q(\rf_shift_reg.x[3][10] ));
 sg13g2_dfrbp_1 _3781_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net330),
    .D(_0176_),
    .Q_N(_1748_),
    .Q(\rf_shift_reg.x[3][11] ));
 sg13g2_dfrbp_1 _3782_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net329),
    .D(net1091),
    .Q_N(_1747_),
    .Q(\rf_shift_reg.x[3][12] ));
 sg13g2_dfrbp_1 _3783_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net328),
    .D(net883),
    .Q_N(_1746_),
    .Q(\rf_shift_reg.x[3][13] ));
 sg13g2_dfrbp_1 _3784_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net327),
    .D(_0179_),
    .Q_N(_1745_),
    .Q(\rf_shift_reg.x[3][14] ));
 sg13g2_dfrbp_1 _3785_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net326),
    .D(net1001),
    .Q_N(_1744_),
    .Q(\rf_shift_reg.x[3][15] ));
 sg13g2_dfrbp_1 _3786_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net325),
    .D(_0181_),
    .Q_N(_1743_),
    .Q(\rf_shift_reg.x[3][16] ));
 sg13g2_dfrbp_1 _3787_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net324),
    .D(net739),
    .Q_N(_1742_),
    .Q(\rf_shift_reg.x[3][17] ));
 sg13g2_dfrbp_1 _3788_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net323),
    .D(_0183_),
    .Q_N(_1741_),
    .Q(\rf_shift_reg.x[3][18] ));
 sg13g2_dfrbp_1 _3789_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net322),
    .D(net727),
    .Q_N(_1740_),
    .Q(\rf_shift_reg.x[3][19] ));
 sg13g2_dfrbp_1 _3790_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net321),
    .D(_0185_),
    .Q_N(_1739_),
    .Q(\rf_shift_reg.x[3][20] ));
 sg13g2_dfrbp_1 _3791_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net320),
    .D(net803),
    .Q_N(_1738_),
    .Q(\rf_shift_reg.x[3][21] ));
 sg13g2_dfrbp_1 _3792_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net319),
    .D(_0187_),
    .Q_N(_1737_),
    .Q(\rf_shift_reg.x[3][22] ));
 sg13g2_dfrbp_1 _3793_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net318),
    .D(_0188_),
    .Q_N(_1736_),
    .Q(\rf_shift_reg.x[3][23] ));
 sg13g2_dfrbp_1 _3794_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net317),
    .D(_0189_),
    .Q_N(_1735_),
    .Q(\rf_shift_reg.x[3][24] ));
 sg13g2_dfrbp_1 _3795_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net316),
    .D(net791),
    .Q_N(_1734_),
    .Q(\rf_shift_reg.x[3][25] ));
 sg13g2_dfrbp_1 _3796_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net315),
    .D(_0191_),
    .Q_N(_1733_),
    .Q(\rf_shift_reg.x[3][26] ));
 sg13g2_dfrbp_1 _3797_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net314),
    .D(_0192_),
    .Q_N(_1732_),
    .Q(\rf_shift_reg.x[3][27] ));
 sg13g2_dfrbp_1 _3798_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net313),
    .D(net704),
    .Q_N(_1731_),
    .Q(\rf_shift_reg.x[3][28] ));
 sg13g2_dfrbp_1 _3799_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net312),
    .D(_0194_),
    .Q_N(_1730_),
    .Q(\rf_shift_reg.x[3][29] ));
 sg13g2_dfrbp_1 _3800_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net311),
    .D(net679),
    .Q_N(_1729_),
    .Q(\rf_shift_reg.x[3][30] ));
 sg13g2_dfrbp_1 _3801_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net310),
    .D(net1187),
    .Q_N(_1728_),
    .Q(\rf_shift_reg.x[3][31] ));
 sg13g2_dfrbp_1 _3802_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net309),
    .D(net653),
    .Q_N(_1727_),
    .Q(\rf_shift_reg.rdata[4] ));
 sg13g2_dfrbp_1 _3803_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net308),
    .D(_0198_),
    .Q_N(_1726_),
    .Q(\rf_shift_reg.x[4][1] ));
 sg13g2_dfrbp_1 _3804_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net307),
    .D(_0199_),
    .Q_N(_1725_),
    .Q(\rf_shift_reg.x[4][2] ));
 sg13g2_dfrbp_1 _3805_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net306),
    .D(_0200_),
    .Q_N(_1724_),
    .Q(\rf_shift_reg.x[4][3] ));
 sg13g2_dfrbp_1 _3806_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net305),
    .D(net1067),
    .Q_N(_1723_),
    .Q(\rf_shift_reg.x[4][4] ));
 sg13g2_dfrbp_1 _3807_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net304),
    .D(net1041),
    .Q_N(_1722_),
    .Q(\rf_shift_reg.x[4][5] ));
 sg13g2_dfrbp_1 _3808_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net303),
    .D(net936),
    .Q_N(_1721_),
    .Q(\rf_shift_reg.x[4][6] ));
 sg13g2_dfrbp_1 _3809_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net302),
    .D(net860),
    .Q_N(_1720_),
    .Q(\rf_shift_reg.x[4][7] ));
 sg13g2_dfrbp_1 _3810_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net301),
    .D(_0205_),
    .Q_N(_1719_),
    .Q(\rf_shift_reg.x[4][8] ));
 sg13g2_dfrbp_1 _3811_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net300),
    .D(_0206_),
    .Q_N(_1718_),
    .Q(\rf_shift_reg.x[4][9] ));
 sg13g2_dfrbp_1 _3812_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net299),
    .D(_0207_),
    .Q_N(_1717_),
    .Q(\rf_shift_reg.x[4][10] ));
 sg13g2_dfrbp_1 _3813_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net298),
    .D(net956),
    .Q_N(_1716_),
    .Q(\rf_shift_reg.x[4][11] ));
 sg13g2_dfrbp_1 _3814_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net297),
    .D(_0209_),
    .Q_N(_1715_),
    .Q(\rf_shift_reg.x[4][12] ));
 sg13g2_dfrbp_1 _3815_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net296),
    .D(_0210_),
    .Q_N(_1714_),
    .Q(\rf_shift_reg.x[4][13] ));
 sg13g2_dfrbp_1 _3816_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net295),
    .D(net986),
    .Q_N(_1713_),
    .Q(\rf_shift_reg.x[4][14] ));
 sg13g2_dfrbp_1 _3817_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net294),
    .D(net965),
    .Q_N(_1712_),
    .Q(\rf_shift_reg.x[4][15] ));
 sg13g2_dfrbp_1 _3818_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net293),
    .D(_0213_),
    .Q_N(_1711_),
    .Q(\rf_shift_reg.x[4][16] ));
 sg13g2_dfrbp_1 _3819_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net292),
    .D(net866),
    .Q_N(_1710_),
    .Q(\rf_shift_reg.x[4][17] ));
 sg13g2_dfrbp_1 _3820_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net291),
    .D(_0215_),
    .Q_N(_1709_),
    .Q(\rf_shift_reg.x[4][18] ));
 sg13g2_dfrbp_1 _3821_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net290),
    .D(net677),
    .Q_N(_1708_),
    .Q(\rf_shift_reg.x[4][19] ));
 sg13g2_dfrbp_1 _3822_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net289),
    .D(_0217_),
    .Q_N(_1707_),
    .Q(\rf_shift_reg.x[4][20] ));
 sg13g2_dfrbp_1 _3823_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net288),
    .D(net751),
    .Q_N(_1706_),
    .Q(\rf_shift_reg.x[4][21] ));
 sg13g2_dfrbp_1 _3824_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net287),
    .D(_0219_),
    .Q_N(_1705_),
    .Q(\rf_shift_reg.x[4][22] ));
 sg13g2_dfrbp_1 _3825_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net286),
    .D(net833),
    .Q_N(_1704_),
    .Q(\rf_shift_reg.x[4][23] ));
 sg13g2_dfrbp_1 _3826_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net285),
    .D(_0221_),
    .Q_N(_1703_),
    .Q(\rf_shift_reg.x[4][24] ));
 sg13g2_dfrbp_1 _3827_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net284),
    .D(net998),
    .Q_N(_1702_),
    .Q(\rf_shift_reg.x[4][25] ));
 sg13g2_dfrbp_1 _3828_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net283),
    .D(net903),
    .Q_N(_1701_),
    .Q(\rf_shift_reg.x[4][26] ));
 sg13g2_dfrbp_1 _3829_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net282),
    .D(_0224_),
    .Q_N(_1700_),
    .Q(\rf_shift_reg.x[4][27] ));
 sg13g2_dfrbp_1 _3830_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net281),
    .D(_0225_),
    .Q_N(_1699_),
    .Q(\rf_shift_reg.x[4][28] ));
 sg13g2_dfrbp_1 _3831_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net280),
    .D(net961),
    .Q_N(_1698_),
    .Q(\rf_shift_reg.x[4][29] ));
 sg13g2_dfrbp_1 _3832_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net279),
    .D(_0227_),
    .Q_N(_1697_),
    .Q(\rf_shift_reg.x[4][30] ));
 sg13g2_dfrbp_1 _3833_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net277),
    .D(net731),
    .Q_N(_1696_),
    .Q(\rf_shift_reg.x[4][31] ));
 sg13g2_dfrbp_1 _3834_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net276),
    .D(net668),
    .Q_N(_1695_),
    .Q(\rf_shift_reg.rdata[5] ));
 sg13g2_dfrbp_1 _3835_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net275),
    .D(_0230_),
    .Q_N(_1694_),
    .Q(\rf_shift_reg.x[5][1] ));
 sg13g2_dfrbp_1 _3836_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net274),
    .D(net945),
    .Q_N(_1693_),
    .Q(\rf_shift_reg.x[5][2] ));
 sg13g2_dfrbp_1 _3837_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net273),
    .D(net924),
    .Q_N(_1692_),
    .Q(\rf_shift_reg.x[5][3] ));
 sg13g2_dfrbp_1 _3838_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net272),
    .D(_0233_),
    .Q_N(_1691_),
    .Q(\rf_shift_reg.x[5][4] ));
 sg13g2_dfrbp_1 _3839_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net271),
    .D(_0234_),
    .Q_N(_1690_),
    .Q(\rf_shift_reg.x[5][5] ));
 sg13g2_dfrbp_1 _3840_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net270),
    .D(net967),
    .Q_N(_1689_),
    .Q(\rf_shift_reg.x[5][6] ));
 sg13g2_dfrbp_1 _3841_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net269),
    .D(net909),
    .Q_N(_1688_),
    .Q(\rf_shift_reg.x[5][7] ));
 sg13g2_dfrbp_1 _3842_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net268),
    .D(net848),
    .Q_N(_1687_),
    .Q(\rf_shift_reg.x[5][8] ));
 sg13g2_dfrbp_1 _3843_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net267),
    .D(_0238_),
    .Q_N(_1686_),
    .Q(\rf_shift_reg.x[5][9] ));
 sg13g2_dfrbp_1 _3844_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net266),
    .D(_0239_),
    .Q_N(_1685_),
    .Q(\rf_shift_reg.x[5][10] ));
 sg13g2_dfrbp_1 _3845_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net265),
    .D(net857),
    .Q_N(_1684_),
    .Q(\rf_shift_reg.x[5][11] ));
 sg13g2_dfrbp_1 _3846_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net264),
    .D(_0241_),
    .Q_N(_1683_),
    .Q(\rf_shift_reg.x[5][12] ));
 sg13g2_dfrbp_1 _3847_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net263),
    .D(_0242_),
    .Q_N(_1682_),
    .Q(\rf_shift_reg.x[5][13] ));
 sg13g2_dfrbp_1 _3848_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net262),
    .D(net952),
    .Q_N(_1681_),
    .Q(\rf_shift_reg.x[5][14] ));
 sg13g2_dfrbp_1 _3849_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net261),
    .D(_0244_),
    .Q_N(_1680_),
    .Q(\rf_shift_reg.x[5][15] ));
 sg13g2_dfrbp_1 _3850_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net260),
    .D(net1054),
    .Q_N(_1679_),
    .Q(\rf_shift_reg.x[5][16] ));
 sg13g2_dfrbp_1 _3851_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net259),
    .D(net1037),
    .Q_N(_1678_),
    .Q(\rf_shift_reg.x[5][17] ));
 sg13g2_dfrbp_1 _3852_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net258),
    .D(net1006),
    .Q_N(_1677_),
    .Q(\rf_shift_reg.x[5][18] ));
 sg13g2_dfrbp_1 _3853_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net257),
    .D(net812),
    .Q_N(_1676_),
    .Q(\rf_shift_reg.x[5][19] ));
 sg13g2_dfrbp_1 _3854_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net256),
    .D(_0249_),
    .Q_N(_1675_),
    .Q(\rf_shift_reg.x[5][20] ));
 sg13g2_dfrbp_1 _3855_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net255),
    .D(net897),
    .Q_N(_1674_),
    .Q(\rf_shift_reg.x[5][21] ));
 sg13g2_dfrbp_1 _3856_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net254),
    .D(_0251_),
    .Q_N(_1673_),
    .Q(\rf_shift_reg.x[5][22] ));
 sg13g2_dfrbp_1 _3857_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net253),
    .D(net943),
    .Q_N(_1672_),
    .Q(\rf_shift_reg.x[5][23] ));
 sg13g2_dfrbp_1 _3858_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net252),
    .D(_0253_),
    .Q_N(_1671_),
    .Q(\rf_shift_reg.x[5][24] ));
 sg13g2_dfrbp_1 _3859_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net251),
    .D(net872),
    .Q_N(_1670_),
    .Q(\rf_shift_reg.x[5][25] ));
 sg13g2_dfrbp_1 _3860_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net250),
    .D(_0255_),
    .Q_N(_1669_),
    .Q(\rf_shift_reg.x[5][26] ));
 sg13g2_dfrbp_1 _3861_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net249),
    .D(_0256_),
    .Q_N(_1668_),
    .Q(\rf_shift_reg.x[5][27] ));
 sg13g2_dfrbp_1 _3862_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net248),
    .D(_0257_),
    .Q_N(_1667_),
    .Q(\rf_shift_reg.x[5][28] ));
 sg13g2_dfrbp_1 _3863_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net245),
    .D(net919),
    .Q_N(_1666_),
    .Q(\rf_shift_reg.x[5][29] ));
 sg13g2_dfrbp_1 _3864_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net244),
    .D(_0259_),
    .Q_N(_1665_),
    .Q(\rf_shift_reg.x[5][30] ));
 sg13g2_dfrbp_1 _3865_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net243),
    .D(net670),
    .Q_N(_1664_),
    .Q(\rf_shift_reg.x[5][31] ));
 sg13g2_dfrbp_1 _3866_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net242),
    .D(net639),
    .Q_N(_0019_),
    .Q(\gpio.o_wb_ack ));
 sg13g2_dfrbp_1 _3867_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net241),
    .D(_0262_),
    .Q_N(_1663_),
    .Q(\dut.xfer.count[0] ));
 sg13g2_dfrbp_1 _3868_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net239),
    .D(_0263_),
    .Q_N(_1662_),
    .Q(\dut.xfer.count[1] ));
 sg13g2_dfrbp_1 _3869_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net190),
    .D(_0264_),
    .Q_N(_0088_),
    .Q(\dut.xfer.count[2] ));
 sg13g2_dfrbp_1 _3870_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net191),
    .D(_0001_),
    .Q_N(_1830_),
    .Q(\dut.state[0] ));
 sg13g2_dfrbp_1 _3871_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net192),
    .D(_0000_),
    .Q_N(_1831_),
    .Q(\dut.state[1] ));
 sg13g2_dfrbp_1 _3872_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net193),
    .D(net1099),
    .Q_N(_1832_),
    .Q(\dut.state[2] ));
 sg13g2_dfrbp_1 _3873_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net194),
    .D(net1238),
    .Q_N(_1833_),
    .Q(\dut.state[3] ));
 sg13g2_dfrbp_1 _3874_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net195),
    .D(net721),
    .Q_N(_1834_),
    .Q(\dut.state[4] ));
 sg13g2_dfrbp_1 _3875_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net196),
    .D(net855),
    .Q_N(_1835_),
    .Q(\dut.state[5] ));
 sg13g2_dfrbp_1 _3876_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net197),
    .D(net1192),
    .Q_N(_1836_),
    .Q(\dut.state[6] ));
 sg13g2_dfrbp_1 _3877_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net198),
    .D(_0010_),
    .Q_N(_1837_),
    .Q(\dut.state[7] ));
 sg13g2_dfrbp_1 _3878_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net199),
    .D(_0011_),
    .Q_N(_1838_),
    .Q(\dut.state[8] ));
 sg13g2_dfrbp_1 _3879_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net200),
    .D(_0012_),
    .Q_N(_1839_),
    .Q(\dut.state[9] ));
 sg13g2_dfrbp_1 _3880_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net201),
    .D(_0002_),
    .Q_N(_1840_),
    .Q(\dut.state[10] ));
 sg13g2_dfrbp_1 _3881_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net213),
    .D(net1179),
    .Q_N(_1841_),
    .Q(\dut.state[11] ));
 sg13g2_dfrbp_1 _3882_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net237),
    .D(net1233),
    .Q_N(_1661_),
    .Q(\dut.state[12] ));
 sg13g2_dfrbp_1 _3883_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net235),
    .D(_0265_),
    .Q_N(_1660_),
    .Q(\rf_shift_reg.rreq_2r ));
 sg13g2_dfrbp_1 _3884_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net234),
    .D(net1206),
    .Q_N(_1659_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _3885_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net232),
    .D(net1214),
    .Q_N(_1658_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _3886_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net230),
    .D(net1201),
    .Q_N(_1657_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _3887_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net228),
    .D(net1245),
    .Q_N(_1656_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _3888_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net226),
    .D(net1227),
    .Q_N(_1655_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _3889_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net224),
    .D(_0271_),
    .Q_N(_1654_),
    .Q(\cpu.immdec.imm11_7[0] ));
 sg13g2_dfrbp_1 _3890_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net223),
    .D(_0272_),
    .Q_N(_1653_),
    .Q(\cpu.immdec.imm11_7[1] ));
 sg13g2_dfrbp_1 _3891_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net222),
    .D(_0273_),
    .Q_N(_1652_),
    .Q(\cpu.immdec.imm11_7[2] ));
 sg13g2_dfrbp_1 _3892_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net221),
    .D(_0274_),
    .Q_N(_1651_),
    .Q(\cpu.immdec.imm11_7[3] ));
 sg13g2_dfrbp_1 _3893_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net246),
    .D(_0275_),
    .Q_N(_1842_),
    .Q(\cpu.immdec.imm11_7[4] ));
 sg13g2_dfrbp_1 _3894_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net220),
    .D(net1337),
    .Q_N(_1650_),
    .Q(\cpu.alu.add_cy_r ));
 sg13g2_dfrbp_1 _3895_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net219),
    .D(_0276_),
    .Q_N(_1649_),
    .Q(\cpu.ctrl.o_ibus_adr[0] ));
 sg13g2_dfrbp_1 _3896_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net217),
    .D(_0277_),
    .Q_N(_1648_),
    .Q(\cpu.ctrl.o_ibus_adr[1] ));
 sg13g2_dfrbp_1 _3897_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net215),
    .D(_0278_),
    .Q_N(_0023_),
    .Q(\cpu.ctrl.o_ibus_adr[2] ));
 sg13g2_dfrbp_1 _3898_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net212),
    .D(_0279_),
    .Q_N(_0025_),
    .Q(\cpu.ctrl.o_ibus_adr[3] ));
 sg13g2_dfrbp_1 _3899_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net210),
    .D(_0280_),
    .Q_N(_0028_),
    .Q(\cpu.ctrl.o_ibus_adr[4] ));
 sg13g2_dfrbp_1 _3900_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net208),
    .D(_0281_),
    .Q_N(_0031_),
    .Q(\cpu.ctrl.o_ibus_adr[5] ));
 sg13g2_dfrbp_1 _3901_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net206),
    .D(_0282_),
    .Q_N(_0034_),
    .Q(\cpu.ctrl.o_ibus_adr[6] ));
 sg13g2_dfrbp_1 _3902_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net204),
    .D(_0283_),
    .Q_N(_0037_),
    .Q(\cpu.ctrl.o_ibus_adr[7] ));
 sg13g2_dfrbp_1 _3903_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net202),
    .D(_0284_),
    .Q_N(_0040_),
    .Q(\cpu.ctrl.o_ibus_adr[8] ));
 sg13g2_dfrbp_1 _3904_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net187),
    .D(_0285_),
    .Q_N(_0043_),
    .Q(\cpu.ctrl.o_ibus_adr[9] ));
 sg13g2_dfrbp_1 _3905_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net185),
    .D(_0286_),
    .Q_N(_0046_),
    .Q(\cpu.ctrl.o_ibus_adr[10] ));
 sg13g2_dfrbp_1 _3906_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net183),
    .D(_0287_),
    .Q_N(_0049_),
    .Q(\cpu.ctrl.o_ibus_adr[11] ));
 sg13g2_dfrbp_1 _3907_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net181),
    .D(_0288_),
    .Q_N(_0052_),
    .Q(\cpu.ctrl.o_ibus_adr[12] ));
 sg13g2_dfrbp_1 _3908_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net179),
    .D(_0289_),
    .Q_N(_0055_),
    .Q(\cpu.ctrl.o_ibus_adr[13] ));
 sg13g2_dfrbp_1 _3909_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net177),
    .D(_0290_),
    .Q_N(_0058_),
    .Q(\cpu.ctrl.o_ibus_adr[14] ));
 sg13g2_dfrbp_1 _3910_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net175),
    .D(_0291_),
    .Q_N(_0061_),
    .Q(\cpu.ctrl.o_ibus_adr[15] ));
 sg13g2_dfrbp_1 _3911_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net173),
    .D(_0292_),
    .Q_N(_0064_),
    .Q(\cpu.ctrl.o_ibus_adr[16] ));
 sg13g2_dfrbp_1 _3912_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net171),
    .D(_0293_),
    .Q_N(_0067_),
    .Q(\cpu.ctrl.o_ibus_adr[17] ));
 sg13g2_dfrbp_1 _3913_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net169),
    .D(_0294_),
    .Q_N(_0070_),
    .Q(\cpu.ctrl.o_ibus_adr[18] ));
 sg13g2_dfrbp_1 _3914_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net167),
    .D(_0295_),
    .Q_N(_0073_),
    .Q(\cpu.ctrl.o_ibus_adr[19] ));
 sg13g2_dfrbp_1 _3915_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net165),
    .D(_0296_),
    .Q_N(_0076_),
    .Q(\cpu.ctrl.o_ibus_adr[20] ));
 sg13g2_dfrbp_1 _3916_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net163),
    .D(_0297_),
    .Q_N(_0079_),
    .Q(\cpu.ctrl.o_ibus_adr[21] ));
 sg13g2_dfrbp_1 _3917_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net161),
    .D(_0298_),
    .Q_N(_0082_),
    .Q(\cpu.ctrl.o_ibus_adr[22] ));
 sg13g2_dfrbp_1 _3918_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net159),
    .D(_0299_),
    .Q_N(_0085_),
    .Q(\cpu.ctrl.o_ibus_adr[23] ));
 sg13g2_dfrbp_1 _3919_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net157),
    .D(_0300_),
    .Q_N(_1647_),
    .Q(\cpu.ctrl.o_ibus_adr[24] ));
 sg13g2_dfrbp_1 _3920_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net155),
    .D(_0301_),
    .Q_N(_1646_),
    .Q(\cpu.ctrl.o_ibus_adr[25] ));
 sg13g2_dfrbp_1 _3921_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net153),
    .D(_0302_),
    .Q_N(_1645_),
    .Q(\cpu.ctrl.o_ibus_adr[26] ));
 sg13g2_dfrbp_1 _3922_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net151),
    .D(_0303_),
    .Q_N(_1644_),
    .Q(\cpu.ctrl.o_ibus_adr[27] ));
 sg13g2_dfrbp_1 _3923_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net149),
    .D(_0304_),
    .Q_N(_1643_),
    .Q(\cpu.ctrl.o_ibus_adr[28] ));
 sg13g2_dfrbp_1 _3924_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net147),
    .D(_0305_),
    .Q_N(_1642_),
    .Q(\cpu.ctrl.o_ibus_adr[29] ));
 sg13g2_dfrbp_1 _3925_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net145),
    .D(_0306_),
    .Q_N(_1641_),
    .Q(\cpu.ctrl.o_ibus_adr[30] ));
 sg13g2_dfrbp_1 _3926_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net247),
    .D(net1060),
    .Q_N(_1843_),
    .Q(\cpu.ctrl.o_ibus_adr[31] ));
 sg13g2_dfrbp_1 _3927_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net278),
    .D(net1131),
    .Q_N(_1844_),
    .Q(\cpu.ctrl.pc_plus_4_cy_r ));
 sg13g2_dfrbp_1 _3928_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net143),
    .D(net1231),
    .Q_N(_1640_),
    .Q(\cpu.ctrl.pc_plus_offset_cy_r ));
 sg13g2_dfrbp_1 _3929_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net141),
    .D(net1159),
    .Q_N(_0022_),
    .Q(\cpu.bufreg.data[2] ));
 sg13g2_dfrbp_1 _3930_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net140),
    .D(net1149),
    .Q_N(_0024_),
    .Q(\cpu.bufreg.data[3] ));
 sg13g2_dfrbp_1 _3931_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net139),
    .D(_0310_),
    .Q_N(_0027_),
    .Q(\cpu.bufreg.data[4] ));
 sg13g2_dfrbp_1 _3932_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net138),
    .D(net876),
    .Q_N(_0030_),
    .Q(\cpu.bufreg.data[5] ));
 sg13g2_dfrbp_1 _3933_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net137),
    .D(_0312_),
    .Q_N(_0033_),
    .Q(\cpu.bufreg.data[6] ));
 sg13g2_dfrbp_1 _3934_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net136),
    .D(_0313_),
    .Q_N(_0036_),
    .Q(\cpu.bufreg.data[7] ));
 sg13g2_dfrbp_1 _3935_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net135),
    .D(net1118),
    .Q_N(_0039_),
    .Q(\cpu.bufreg.data[8] ));
 sg13g2_dfrbp_1 _3936_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net134),
    .D(net1049),
    .Q_N(_0042_),
    .Q(\cpu.bufreg.data[9] ));
 sg13g2_dfrbp_1 _3937_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net133),
    .D(_0316_),
    .Q_N(_0045_),
    .Q(\cpu.bufreg.data[10] ));
 sg13g2_dfrbp_1 _3938_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net132),
    .D(net714),
    .Q_N(_0048_),
    .Q(\cpu.bufreg.data[11] ));
 sg13g2_dfrbp_1 _3939_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net131),
    .D(_0318_),
    .Q_N(_0051_),
    .Q(\cpu.bufreg.data[12] ));
 sg13g2_dfrbp_1 _3940_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net130),
    .D(_0319_),
    .Q_N(_0054_),
    .Q(\cpu.bufreg.data[13] ));
 sg13g2_dfrbp_1 _3941_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net129),
    .D(net941),
    .Q_N(_0057_),
    .Q(\cpu.bufreg.data[14] ));
 sg13g2_dfrbp_1 _3942_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net128),
    .D(_0321_),
    .Q_N(_0060_),
    .Q(\cpu.bufreg.data[15] ));
 sg13g2_dfrbp_1 _3943_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net127),
    .D(_0322_),
    .Q_N(_0063_),
    .Q(\cpu.bufreg.data[16] ));
 sg13g2_dfrbp_1 _3944_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net126),
    .D(_0323_),
    .Q_N(_0066_),
    .Q(\cpu.bufreg.data[17] ));
 sg13g2_dfrbp_1 _3945_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net125),
    .D(net1012),
    .Q_N(_0069_),
    .Q(\cpu.bufreg.data[18] ));
 sg13g2_dfrbp_1 _3946_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net124),
    .D(_0325_),
    .Q_N(_0072_),
    .Q(\cpu.bufreg.data[19] ));
 sg13g2_dfrbp_1 _3947_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net123),
    .D(net977),
    .Q_N(_0075_),
    .Q(\cpu.bufreg.data[20] ));
 sg13g2_dfrbp_1 _3948_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net122),
    .D(_0327_),
    .Q_N(_0078_),
    .Q(\cpu.bufreg.data[21] ));
 sg13g2_dfrbp_1 _3949_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net121),
    .D(net1164),
    .Q_N(_0081_),
    .Q(\cpu.bufreg.data[22] ));
 sg13g2_dfrbp_1 _3950_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net120),
    .D(net889),
    .Q_N(_0084_),
    .Q(\cpu.bufreg.data[23] ));
 sg13g2_dfrbp_1 _3951_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net119),
    .D(_0330_),
    .Q_N(_1639_),
    .Q(\cpu.bufreg.data[24] ));
 sg13g2_dfrbp_1 _3952_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net118),
    .D(net932),
    .Q_N(_1638_),
    .Q(\cpu.bufreg.data[25] ));
 sg13g2_dfrbp_1 _3953_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net117),
    .D(_0332_),
    .Q_N(_1637_),
    .Q(\cpu.bufreg.data[26] ));
 sg13g2_dfrbp_1 _3954_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net116),
    .D(_0333_),
    .Q_N(_1636_),
    .Q(\cpu.bufreg.data[27] ));
 sg13g2_dfrbp_1 _3955_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net115),
    .D(_0334_),
    .Q_N(_1635_),
    .Q(\cpu.bufreg.data[28] ));
 sg13g2_dfrbp_1 _3956_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net114),
    .D(_0335_),
    .Q_N(_1634_),
    .Q(\cpu.bufreg.data[29] ));
 sg13g2_dfrbp_1 _3957_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net113),
    .D(net659),
    .Q_N(_1633_),
    .Q(\cpu.bufreg.data[30] ));
 sg13g2_dfrbp_1 _3958_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net397),
    .D(net1284),
    .Q_N(_1845_),
    .Q(\cpu.bufreg.data[31] ));
 sg13g2_dfrbp_1 _3959_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net112),
    .D(_0014_),
    .Q_N(_1632_),
    .Q(\cpu.bufreg.c_r ));
 sg13g2_dfrbp_1 _3960_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net111),
    .D(_0338_),
    .Q_N(_1631_),
    .Q(\cpu.alu.cmp_r ));
 sg13g2_dfrbp_1 _3961_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net110),
    .D(_0339_),
    .Q_N(_1630_),
    .Q(\cpu.bufreg.i_sh_signed ));
 sg13g2_dfrbp_1 _3962_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net109),
    .D(net996),
    .Q_N(_1629_),
    .Q(\cpu.immdec.imm31 ));
 sg13g2_dfrbp_1 _3963_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net108),
    .D(net1282),
    .Q_N(_1628_),
    .Q(\cpu.immdec.imm19_12_20[0] ));
 sg13g2_dfrbp_1 _3964_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net107),
    .D(net1287),
    .Q_N(_1627_),
    .Q(\cpu.immdec.imm19_12_20[1] ));
 sg13g2_dfrbp_1 _3965_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net106),
    .D(net1240),
    .Q_N(_1626_),
    .Q(\cpu.immdec.imm19_12_20[2] ));
 sg13g2_dfrbp_1 _3966_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net105),
    .D(_0344_),
    .Q_N(_1625_),
    .Q(\cpu.immdec.imm19_12_20[3] ));
 sg13g2_dfrbp_1 _3967_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net104),
    .D(net1255),
    .Q_N(_1624_),
    .Q(\cpu.csr_imm ));
 sg13g2_dfrbp_1 _3968_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net103),
    .D(_0346_),
    .Q_N(_1623_),
    .Q(\cpu.immdec.imm19_12_20[5] ));
 sg13g2_dfrbp_1 _3969_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net102),
    .D(_0347_),
    .Q_N(_1622_),
    .Q(\cpu.immdec.imm19_12_20[6] ));
 sg13g2_dfrbp_1 _3970_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net101),
    .D(net870),
    .Q_N(_1621_),
    .Q(\cpu.immdec.imm19_12_20[7] ));
 sg13g2_dfrbp_1 _3971_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net100),
    .D(_0349_),
    .Q_N(_1620_),
    .Q(\cpu.immdec.imm19_12_20[8] ));
 sg13g2_dfrbp_1 _3972_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net99),
    .D(net1235),
    .Q_N(_1619_),
    .Q(\cpu.immdec.imm7 ));
 sg13g2_dfrbp_1 _3973_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net98),
    .D(net1253),
    .Q_N(_1618_),
    .Q(\cpu.immdec.imm30_25[0] ));
 sg13g2_dfrbp_1 _3974_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net97),
    .D(net825),
    .Q_N(_1617_),
    .Q(\cpu.immdec.imm30_25[1] ));
 sg13g2_dfrbp_1 _3975_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net96),
    .D(net798),
    .Q_N(_1616_),
    .Q(\cpu.immdec.imm30_25[2] ));
 sg13g2_dfrbp_1 _3976_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net95),
    .D(net774),
    .Q_N(_1615_),
    .Q(\cpu.immdec.imm30_25[3] ));
 sg13g2_dfrbp_1 _3977_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net94),
    .D(net808),
    .Q_N(_1614_),
    .Q(\cpu.immdec.imm30_25[4] ));
 sg13g2_dfrbp_1 _3978_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net93),
    .D(net796),
    .Q_N(_1613_),
    .Q(\cpu.immdec.imm30_25[5] ));
 sg13g2_dfrbp_1 _3979_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net92),
    .D(_0357_),
    .Q_N(_1612_),
    .Q(\cpu.immdec.imm24_20[0] ));
 sg13g2_dfrbp_1 _3980_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net91),
    .D(net1219),
    .Q_N(_1611_),
    .Q(\cpu.immdec.imm24_20[1] ));
 sg13g2_dfrbp_1 _3981_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net90),
    .D(_0359_),
    .Q_N(_1610_),
    .Q(\cpu.immdec.imm24_20[2] ));
 sg13g2_dfrbp_1 _3982_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net89),
    .D(net1052),
    .Q_N(_1609_),
    .Q(\cpu.immdec.imm24_20[3] ));
 sg13g2_dfrbp_1 _3983_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net88),
    .D(_0361_),
    .Q_N(_1608_),
    .Q(\cpu.immdec.imm24_20[4] ));
 sg13g2_dfrbp_1 _3984_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net87),
    .D(net1210),
    .Q_N(_1607_),
    .Q(\cpu.decode.co_ebreak ));
 sg13g2_dfrbp_1 _3985_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net86),
    .D(_0363_),
    .Q_N(_1606_),
    .Q(\cpu.bne_or_bge ));
 sg13g2_dfrbp_1 _3986_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net85),
    .D(_0364_),
    .Q_N(_1605_),
    .Q(\cpu.decode.co_mem_word ));
 sg13g2_dfrbp_1 _3987_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net84),
    .D(_0365_),
    .Q_N(_0017_),
    .Q(\cpu.csr_d_sel ));
 sg13g2_dfrbp_1 _3988_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net83),
    .D(net1314),
    .Q_N(_0091_),
    .Q(\cpu.decode.opcode[0] ));
 sg13g2_dfrbp_1 _3989_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net82),
    .D(net1303),
    .Q_N(_1604_),
    .Q(\cpu.decode.opcode[1] ));
 sg13g2_dfrbp_1 _3990_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net81),
    .D(net1296),
    .Q_N(_0092_),
    .Q(\cpu.decode.opcode[2] ));
 sg13g2_dfrbp_1 _3991_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net80),
    .D(net1258),
    .Q_N(_0020_),
    .Q(\cpu.bufreg2.i_op_b_sel ));
 sg13g2_dfrbp_1 _3992_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net79),
    .D(net1269),
    .Q_N(_0090_),
    .Q(\cpu.branch_op ));
 sg13g2_dfrbp_1 _3993_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net78),
    .D(net1324),
    .Q_N(_0018_),
    .Q(\cpu.bufreg2.dat[0] ));
 sg13g2_dfrbp_1 _3994_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net77),
    .D(net1326),
    .Q_N(_1603_),
    .Q(\cpu.bufreg2.dat[1] ));
 sg13g2_dfrbp_1 _3995_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net76),
    .D(_0373_),
    .Q_N(_1602_),
    .Q(\cpu.bufreg2.dat[2] ));
 sg13g2_dfrbp_1 _3996_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net75),
    .D(net1301),
    .Q_N(_1601_),
    .Q(\cpu.bufreg2.dat[3] ));
 sg13g2_dfrbp_1 _3997_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net74),
    .D(_0375_),
    .Q_N(_1600_),
    .Q(\cpu.bufreg2.dat[4] ));
 sg13g2_dfrbp_1 _3998_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net73),
    .D(_0376_),
    .Q_N(_1599_),
    .Q(\cpu.bufreg2.dat[5] ));
 sg13g2_dfrbp_1 _3999_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net72),
    .D(net697),
    .Q_N(_1598_),
    .Q(\cpu.bufreg2.dat[6] ));
 sg13g2_dfrbp_1 _4000_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net71),
    .D(net1199),
    .Q_N(_1597_),
    .Q(\cpu.bufreg2.dat[7] ));
 sg13g2_dfrbp_1 _4001_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net70),
    .D(net1208),
    .Q_N(_1596_),
    .Q(\cpu.bufreg2.dat[8] ));
 sg13g2_dfrbp_1 _4002_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net69),
    .D(net1058),
    .Q_N(_1595_),
    .Q(\cpu.bufreg2.dat[9] ));
 sg13g2_dfrbp_1 _4003_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net68),
    .D(net814),
    .Q_N(_1594_),
    .Q(\cpu.bufreg2.dat[10] ));
 sg13g2_dfrbp_1 _4004_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net67),
    .D(_0382_),
    .Q_N(_1593_),
    .Q(\cpu.bufreg2.dat[11] ));
 sg13g2_dfrbp_1 _4005_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net66),
    .D(net787),
    .Q_N(_1592_),
    .Q(\cpu.bufreg2.dat[12] ));
 sg13g2_dfrbp_1 _4006_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net65),
    .D(net1085),
    .Q_N(_1591_),
    .Q(\cpu.bufreg2.dat[13] ));
 sg13g2_dfrbp_1 _4007_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net64),
    .D(net699),
    .Q_N(_1590_),
    .Q(\cpu.bufreg2.dat[14] ));
 sg13g2_dfrbp_1 _4008_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net63),
    .D(net930),
    .Q_N(_1589_),
    .Q(\cpu.bufreg2.dat[15] ));
 sg13g2_dfrbp_1 _4009_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net62),
    .D(net1243),
    .Q_N(_1588_),
    .Q(\cpu.bufreg2.dat[16] ));
 sg13g2_dfrbp_1 _4010_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net61),
    .D(net1197),
    .Q_N(_1587_),
    .Q(\cpu.bufreg2.dat[17] ));
 sg13g2_dfrbp_1 _4011_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net60),
    .D(net673),
    .Q_N(_1586_),
    .Q(\cpu.bufreg2.dat[18] ));
 sg13g2_dfrbp_1 _4012_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net59),
    .D(_0390_),
    .Q_N(_1585_),
    .Q(\cpu.bufreg2.dat[19] ));
 sg13g2_dfrbp_1 _4013_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net58),
    .D(net706),
    .Q_N(_1584_),
    .Q(\cpu.bufreg2.dat[20] ));
 sg13g2_dfrbp_1 _4014_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net57),
    .D(net1070),
    .Q_N(_1583_),
    .Q(\cpu.bufreg2.dat[21] ));
 sg13g2_dfrbp_1 _4015_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net56),
    .D(net785),
    .Q_N(_1582_),
    .Q(\cpu.bufreg2.dat[22] ));
 sg13g2_dfrbp_1 _4016_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net55),
    .D(net758),
    .Q_N(_1581_),
    .Q(\cpu.bufreg2.dat[23] ));
 sg13g2_dfrbp_1 _4017_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net54),
    .D(net1273),
    .Q_N(_1580_),
    .Q(\cpu.bufreg2.dat[24] ));
 sg13g2_dfrbp_1 _4018_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net53),
    .D(net691),
    .Q_N(_1579_),
    .Q(\cpu.bufreg2.dat[25] ));
 sg13g2_dfrbp_1 _4019_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net52),
    .D(net1144),
    .Q_N(_1578_),
    .Q(\cpu.bufreg2.dat[26] ));
 sg13g2_dfrbp_1 _4020_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net51),
    .D(net781),
    .Q_N(_1577_),
    .Q(\cpu.bufreg2.dat[27] ));
 sg13g2_dfrbp_1 _4021_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net50),
    .D(net1177),
    .Q_N(_1576_),
    .Q(\cpu.bufreg2.dat[28] ));
 sg13g2_dfrbp_1 _4022_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net49),
    .D(net776),
    .Q_N(_1575_),
    .Q(\cpu.bufreg2.dat[29] ));
 sg13g2_dfrbp_1 _4023_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net48),
    .D(net1111),
    .Q_N(_1574_),
    .Q(\cpu.bufreg2.dat[30] ));
 sg13g2_dfrbp_1 _4024_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net47),
    .D(net760),
    .Q_N(_1573_),
    .Q(\cpu.bufreg2.dat[31] ));
 sg13g2_dfrbp_1 _4025_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net46),
    .D(_0403_),
    .Q_N(_1572_),
    .Q(\cpu.state.stage_two_req ));
 sg13g2_dfrbp_1 _4026_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net45),
    .D(net1223),
    .Q_N(_0089_),
    .Q(\cpu.state.init_done ));
 sg13g2_dfrbp_1 _4027_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net43),
    .D(_0405_),
    .Q_N(_1571_),
    .Q(\cpu.state.cnt_r[0] ));
 sg13g2_dfrbp_1 _4028_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net42),
    .D(_0406_),
    .Q_N(_1570_),
    .Q(\cpu.state.cnt_r[1] ));
 sg13g2_dfrbp_1 _4029_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net41),
    .D(_0407_),
    .Q_N(_1569_),
    .Q(\cpu.state.cnt_r[2] ));
 sg13g2_dfrbp_1 _4030_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net40),
    .D(_0408_),
    .Q_N(_1568_),
    .Q(\cpu.state.cnt_r[3] ));
 sg13g2_dfrbp_1 _4031_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net39),
    .D(net1104),
    .Q_N(_1567_),
    .Q(\cpu.ctrl.i_jump ));
 sg13g2_dfrbp_1 _4032_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net37),
    .D(net1212),
    .Q_N(_1566_),
    .Q(\cpu.state.o_cnt[2] ));
 sg13g2_dfrbp_1 _4033_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net36),
    .D(net1294),
    .Q_N(_1565_),
    .Q(\cpu.mem_bytecnt[0] ));
 sg13g2_dfrbp_1 _4034_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net35),
    .D(net1328),
    .Q_N(_1564_),
    .Q(\cpu.mem_bytecnt[1] ));
 sg13g2_dfrbp_1 _4035_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net34),
    .D(_0413_),
    .Q_N(_1563_),
    .Q(\cpu.mem_if.signbit ));
 sg13g2_dfrbp_1 _4036_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net33),
    .D(net689),
    .Q_N(_1562_),
    .Q(\dut.xfer.xfer_tag[0] ));
 sg13g2_dfrbp_1 _4037_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net31),
    .D(net766),
    .Q_N(_1561_),
    .Q(\dut.xfer.xfer_tag[1] ));
 sg13g2_dfrbp_1 _4038_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net29),
    .D(_0416_),
    .Q_N(_1560_),
    .Q(\dut.xfer.xfer_tag[2] ));
 sg13g2_dfrbp_1 _4039_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net27),
    .D(net1083),
    .Q_N(_1559_),
    .Q(\dut.xfer.next_obuffer[2] ));
 sg13g2_dfrbp_1 _4040_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net26),
    .D(net988),
    .Q_N(_1558_),
    .Q(\dut.xfer.next_obuffer[3] ));
 sg13g2_dfrbp_1 _4041_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net25),
    .D(net823),
    .Q_N(_1557_),
    .Q(\dut.xfer.next_obuffer[4] ));
 sg13g2_dfrbp_1 _4042_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net24),
    .D(net1056),
    .Q_N(_1556_),
    .Q(\dut.xfer.next_obuffer[5] ));
 sg13g2_dfrbp_1 _4043_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net23),
    .D(net880),
    .Q_N(_1555_),
    .Q(\dut.xfer.next_obuffer[6] ));
 sg13g2_dfrbp_1 _4044_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net22),
    .D(_0422_),
    .Q_N(_1554_),
    .Q(\dut.xfer.next_obuffer[7] ));
 sg13g2_dfrbp_1 _4045_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net21),
    .D(net878),
    .Q_N(_1553_),
    .Q(\dut.xfer.obuffer[7] ));
 sg13g2_dfrbp_1 _4046_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net20),
    .D(net862),
    .Q_N(_1552_),
    .Q(\dut.xfer.next_obuffer[1] ));
 sg13g2_dfrbp_1 _4047_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net18),
    .D(net1316),
    .Q_N(_0021_),
    .Q(\dut.rd_addr[2] ));
 sg13g2_dfrbp_1 _4048_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net631),
    .D(net1340),
    .Q_N(_1551_),
    .Q(\dut.rd_addr[3] ));
 sg13g2_dfrbp_1 _4049_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net630),
    .D(net885),
    .Q_N(_0026_),
    .Q(\dut.rd_addr[4] ));
 sg13g2_dfrbp_1 _4050_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net629),
    .D(net922),
    .Q_N(_0029_),
    .Q(\dut.rd_addr[5] ));
 sg13g2_dfrbp_1 _4051_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net628),
    .D(net1120),
    .Q_N(_0032_),
    .Q(\dut.rd_addr[6] ));
 sg13g2_dfrbp_1 _4052_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net627),
    .D(net972),
    .Q_N(_0035_),
    .Q(\dut.rd_addr[7] ));
 sg13g2_dfrbp_1 _4053_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net626),
    .D(net840),
    .Q_N(_0038_),
    .Q(\dut.rd_addr[8] ));
 sg13g2_dfrbp_1 _4054_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net625),
    .D(net846),
    .Q_N(_0041_),
    .Q(\dut.rd_addr[9] ));
 sg13g2_dfrbp_1 _4055_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net624),
    .D(_0433_),
    .Q_N(_0044_),
    .Q(\dut.rd_addr[10] ));
 sg13g2_dfrbp_1 _4056_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net623),
    .D(net741),
    .Q_N(_0047_),
    .Q(\dut.rd_addr[11] ));
 sg13g2_dfrbp_1 _4057_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net622),
    .D(net768),
    .Q_N(_0050_),
    .Q(\dut.rd_addr[12] ));
 sg13g2_dfrbp_1 _4058_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net621),
    .D(net899),
    .Q_N(_0053_),
    .Q(\dut.rd_addr[13] ));
 sg13g2_dfrbp_1 _4059_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net620),
    .D(net1225),
    .Q_N(_0056_),
    .Q(\dut.rd_addr[14] ));
 sg13g2_dfrbp_1 _4060_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net619),
    .D(net710),
    .Q_N(_0059_),
    .Q(\dut.rd_addr[15] ));
 sg13g2_dfrbp_1 _4061_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net618),
    .D(net770),
    .Q_N(_0062_),
    .Q(\dut.rd_addr[16] ));
 sg13g2_dfrbp_1 _4062_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net617),
    .D(net756),
    .Q_N(_0065_),
    .Q(\dut.rd_addr[17] ));
 sg13g2_dfrbp_1 _4063_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net616),
    .D(net842),
    .Q_N(_0068_),
    .Q(\dut.rd_addr[18] ));
 sg13g2_dfrbp_1 _4064_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net615),
    .D(net844),
    .Q_N(_0071_),
    .Q(\dut.rd_addr[19] ));
 sg13g2_dfrbp_1 _4065_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net614),
    .D(net850),
    .Q_N(_0074_),
    .Q(\dut.rd_addr[20] ));
 sg13g2_dfrbp_1 _4066_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net613),
    .D(net743),
    .Q_N(_0077_),
    .Q(\dut.rd_addr[21] ));
 sg13g2_dfrbp_1 _4067_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net612),
    .D(net816),
    .Q_N(_0080_),
    .Q(\dut.rd_addr[22] ));
 sg13g2_dfrbp_1 _4068_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net611),
    .D(net716),
    .Q_N(_0083_),
    .Q(\dut.rd_addr[23] ));
 sg13g2_dfrbp_1 _4069_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net610),
    .D(net1190),
    .Q_N(_1550_),
    .Q(\cpu.bufreg.data[0] ));
 sg13g2_dfrbp_1 _4070_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net609),
    .D(net1291),
    .Q_N(_1549_),
    .Q(\cpu.bufreg.data[1] ));
 sg13g2_dfrbp_1 _4071_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net608),
    .D(_0449_),
    .Q_N(_1548_),
    .Q(\dut.flash_csb ));
 sg13g2_dfrbp_1 _4072_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net606),
    .D(net745),
    .Q_N(_0087_),
    .Q(\dut.flash_clk ));
 sg13g2_dfrbp_1 _4073_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net604),
    .D(net1331),
    .Q_N(_1547_),
    .Q(\dut.xfer.count[3] ));
 sg13g2_dfrbp_1 _4074_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net602),
    .D(net1221),
    .Q_N(_1546_),
    .Q(\dut.xfer.dummy_count[0] ));
 sg13g2_dfrbp_1 _4075_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net600),
    .D(_0453_),
    .Q_N(_1545_),
    .Q(\dut.xfer.dummy_count[1] ));
 sg13g2_dfrbp_1 _4076_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net598),
    .D(_0454_),
    .Q_N(_1544_),
    .Q(\dut.xfer.dummy_count[2] ));
 sg13g2_dfrbp_1 _4077_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net398),
    .D(_0455_),
    .Q_N(_1846_),
    .Q(\dut.xfer.dummy_count[3] ));
 sg13g2_dfrbp_1 _4078_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net399),
    .D(net634),
    .Q_N(_1847_),
    .Q(\dut.dout_tag[0] ));
 sg13g2_dfrbp_1 _4079_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net595),
    .D(net633),
    .Q_N(_1848_),
    .Q(\dut.dout_tag[1] ));
 sg13g2_dfrbp_1 _4080_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net596),
    .D(net632),
    .Q_N(_1543_),
    .Q(\dut.dout_tag[2] ));
 sg13g2_dfrbp_1 _4081_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net594),
    .D(_0456_),
    .Q_N(_1542_),
    .Q(\dut.dout_data[0] ));
 sg13g2_dfrbp_1 _4082_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net593),
    .D(_0457_),
    .Q_N(_1541_),
    .Q(\dut.dout_data[1] ));
 sg13g2_dfrbp_1 _4083_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net592),
    .D(_0458_),
    .Q_N(_1540_),
    .Q(\dut.dout_data[2] ));
 sg13g2_dfrbp_1 _4084_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net591),
    .D(_0459_),
    .Q_N(_1539_),
    .Q(\dut.dout_data[3] ));
 sg13g2_dfrbp_1 _4085_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net590),
    .D(_0460_),
    .Q_N(_1538_),
    .Q(\dut.dout_data[4] ));
 sg13g2_dfrbp_1 _4086_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net589),
    .D(_0461_),
    .Q_N(_1537_),
    .Q(\dut.dout_data[5] ));
 sg13g2_dfrbp_1 _4087_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net588),
    .D(_0462_),
    .Q_N(_1536_),
    .Q(\dut.dout_data[6] ));
 sg13g2_dfrbp_1 _4088_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net587),
    .D(_0463_),
    .Q_N(_1535_),
    .Q(\dut.dout_data[7] ));
 sg13g2_dfrbp_1 _4089_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net440),
    .D(_0464_),
    .Q_N(_1534_),
    .Q(\dut.xfer.fetch ));
 sg13g2_dfrbp_1 _4090_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net439),
    .D(_0465_),
    .Q_N(_1533_),
    .Q(\dut.softreset ));
 sg13g2_dfrbp_1 _4091_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net438),
    .D(_0466_),
    .Q_N(_1532_),
    .Q(\dut.rd_inc ));
 sg13g2_dfrbp_1 _4092_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net436),
    .D(net1216),
    .Q_N(_1531_),
    .Q(\dut.rd_wait ));
 sg13g2_dfrbp_1 _4093_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net434),
    .D(net1260),
    .Q_N(_1530_),
    .Q(\dut.rd_valid ));
 sg13g2_dfrbp_1 _4094_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net432),
    .D(_0469_),
    .Q_N(_1529_),
    .Q(\dut.buffer[16] ));
 sg13g2_dfrbp_1 _4095_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net431),
    .D(_0470_),
    .Q_N(_1528_),
    .Q(\dut.buffer[17] ));
 sg13g2_dfrbp_1 _4096_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net430),
    .D(net984),
    .Q_N(_1527_),
    .Q(\dut.buffer[18] ));
 sg13g2_dfrbp_1 _4097_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net429),
    .D(_0472_),
    .Q_N(_1526_),
    .Q(\dut.buffer[19] ));
 sg13g2_dfrbp_1 _4098_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net428),
    .D(_0473_),
    .Q_N(_1525_),
    .Q(\dut.buffer[20] ));
 sg13g2_dfrbp_1 _4099_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net427),
    .D(_0474_),
    .Q_N(_1524_),
    .Q(\dut.buffer[21] ));
 sg13g2_dfrbp_1 _4100_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net426),
    .D(_0475_),
    .Q_N(_1523_),
    .Q(\dut.buffer[22] ));
 sg13g2_dfrbp_1 _4101_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net425),
    .D(_0476_),
    .Q_N(_1522_),
    .Q(\dut.buffer[23] ));
 sg13g2_dfrbp_1 _4102_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net424),
    .D(_0477_),
    .Q_N(_1521_),
    .Q(\dut.din_rd ));
 sg13g2_dfrbp_1 _4103_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net422),
    .D(_0478_),
    .Q_N(_0086_),
    .Q(\dut.xfer.resetn ));
 sg13g2_dfrbp_1 _4104_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net421),
    .D(net874),
    .Q_N(_1520_),
    .Q(\cpu.bufreg2.i_dat[0] ));
 sg13g2_dfrbp_1 _4105_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net420),
    .D(net1017),
    .Q_N(_1519_),
    .Q(\cpu.bufreg2.i_dat[1] ));
 sg13g2_dfrbp_1 _4106_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net382),
    .D(net836),
    .Q_N(_1518_),
    .Q(\cpu.bufreg2.i_dat[2] ));
 sg13g2_dfrbp_1 _4107_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net380),
    .D(net838),
    .Q_N(_1517_),
    .Q(\cpu.bufreg2.i_dat[3] ));
 sg13g2_dfrbp_1 _4108_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net378),
    .D(net990),
    .Q_N(_1516_),
    .Q(\cpu.bufreg2.i_dat[4] ));
 sg13g2_dfrbp_1 _4109_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net376),
    .D(net737),
    .Q_N(_1515_),
    .Q(\cpu.bufreg2.i_dat[5] ));
 sg13g2_dfrbp_1 _4110_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net374),
    .D(net1034),
    .Q_N(_1514_),
    .Q(\cpu.bufreg2.i_dat[6] ));
 sg13g2_dfrbp_1 _4111_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net240),
    .D(net928),
    .Q_N(_1513_),
    .Q(\cpu.bufreg2.i_dat[7] ));
 sg13g2_dfrbp_1 _4112_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net238),
    .D(net655),
    .Q_N(_1512_),
    .Q(\cpu.bufreg2.i_dat[8] ));
 sg13g2_dfrbp_1 _4113_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net236),
    .D(net895),
    .Q_N(_1511_),
    .Q(\cpu.bufreg2.i_dat[9] ));
 sg13g2_dfrbp_1 _4114_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net233),
    .D(_0489_),
    .Q_N(_1510_),
    .Q(\cpu.bufreg2.i_dat[10] ));
 sg13g2_dfrbp_1 _4115_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net231),
    .D(_0490_),
    .Q_N(_1509_),
    .Q(\cpu.bufreg2.i_dat[11] ));
 sg13g2_dfrbp_1 _4116_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net229),
    .D(net764),
    .Q_N(_1508_),
    .Q(\cpu.bufreg2.i_dat[12] ));
 sg13g2_dfrbp_1 _4117_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net227),
    .D(net748),
    .Q_N(_1507_),
    .Q(\cpu.bufreg2.i_dat[13] ));
 sg13g2_dfrbp_1 _4118_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net225),
    .D(_0493_),
    .Q_N(_1506_),
    .Q(\cpu.bufreg2.i_dat[14] ));
 sg13g2_dfrbp_1 _4119_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net218),
    .D(_0494_),
    .Q_N(_1505_),
    .Q(\cpu.bufreg2.i_dat[15] ));
 sg13g2_dfrbp_1 _4120_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net216),
    .D(net907),
    .Q_N(_1504_),
    .Q(\cpu.bufreg2.i_dat[16] ));
 sg13g2_dfrbp_1 _4121_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net214),
    .D(net938),
    .Q_N(_1503_),
    .Q(\cpu.bufreg2.i_dat[17] ));
 sg13g2_dfrbp_1 _4122_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net211),
    .D(_0497_),
    .Q_N(_1502_),
    .Q(\cpu.bufreg2.i_dat[18] ));
 sg13g2_dfrbp_1 _4123_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net209),
    .D(_0498_),
    .Q_N(_1501_),
    .Q(\cpu.bufreg2.i_dat[19] ));
 sg13g2_dfrbp_1 _4124_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net207),
    .D(net901),
    .Q_N(_1500_),
    .Q(\cpu.bufreg2.i_dat[20] ));
 sg13g2_dfrbp_1 _4125_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net205),
    .D(net1101),
    .Q_N(_1499_),
    .Q(\cpu.bufreg2.i_dat[21] ));
 sg13g2_dfrbp_1 _4126_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net203),
    .D(net1097),
    .Q_N(_1498_),
    .Q(\cpu.bufreg2.i_dat[22] ));
 sg13g2_dfrbp_1 _4127_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net188),
    .D(net1010),
    .Q_N(_1497_),
    .Q(\cpu.bufreg2.i_dat[23] ));
 sg13g2_dfrbp_1 _4128_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net186),
    .D(_0503_),
    .Q_N(_1496_),
    .Q(\cpu.bufreg2.i_dat[24] ));
 sg13g2_dfrbp_1 _4129_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net184),
    .D(_0504_),
    .Q_N(_1495_),
    .Q(\cpu.bufreg2.i_dat[25] ));
 sg13g2_dfrbp_1 _4130_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net182),
    .D(_0505_),
    .Q_N(_1494_),
    .Q(\cpu.bufreg2.i_dat[26] ));
 sg13g2_dfrbp_1 _4131_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net180),
    .D(_0506_),
    .Q_N(_1493_),
    .Q(\cpu.bufreg2.i_dat[27] ));
 sg13g2_dfrbp_1 _4132_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net178),
    .D(_0507_),
    .Q_N(_1492_),
    .Q(\cpu.bufreg2.i_dat[28] ));
 sg13g2_dfrbp_1 _4133_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net176),
    .D(_0508_),
    .Q_N(_1491_),
    .Q(\cpu.bufreg2.i_dat[29] ));
 sg13g2_dfrbp_1 _4134_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net174),
    .D(_0509_),
    .Q_N(_1490_),
    .Q(\cpu.bufreg2.i_dat[30] ));
 sg13g2_dfrbp_1 _4135_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net172),
    .D(_0510_),
    .Q_N(_1489_),
    .Q(\cpu.bufreg2.i_dat[31] ));
 sg13g2_dfrbp_1 _4136_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net170),
    .D(_0511_),
    .Q_N(_1488_),
    .Q(\cpu.state.ibus_cyc ));
 sg13g2_dfrbp_1 _4137_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net168),
    .D(_0512_),
    .Q_N(_1487_),
    .Q(\dut.din_tag[0] ));
 sg13g2_dfrbp_1 _4138_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net164),
    .D(_0513_),
    .Q_N(_1486_),
    .Q(\dut.din_tag[1] ));
 sg13g2_dfrbp_1 _4139_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net160),
    .D(net806),
    .Q_N(_1485_),
    .Q(\dut.din_tag[2] ));
 sg13g2_dfrbp_1 _4140_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net156),
    .D(_0515_),
    .Q_N(_1484_),
    .Q(\dut.buffer[0] ));
 sg13g2_dfrbp_1 _4141_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net154),
    .D(_0516_),
    .Q_N(_1483_),
    .Q(\dut.buffer[1] ));
 sg13g2_dfrbp_1 _4142_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net152),
    .D(_0517_),
    .Q_N(_1482_),
    .Q(\dut.buffer[2] ));
 sg13g2_dfrbp_1 _4143_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net150),
    .D(_0518_),
    .Q_N(_1481_),
    .Q(\dut.buffer[3] ));
 sg13g2_dfrbp_1 _4144_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net148),
    .D(_0519_),
    .Q_N(_1480_),
    .Q(\dut.buffer[4] ));
 sg13g2_dfrbp_1 _4145_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net146),
    .D(_0520_),
    .Q_N(_1479_),
    .Q(\dut.buffer[5] ));
 sg13g2_dfrbp_1 _4146_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net144),
    .D(_0521_),
    .Q_N(_1478_),
    .Q(\dut.buffer[6] ));
 sg13g2_dfrbp_1 _4147_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net142),
    .D(_0522_),
    .Q_N(_1477_),
    .Q(\dut.buffer[7] ));
 sg13g2_dfrbp_1 _4148_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net44),
    .D(_0523_),
    .Q_N(_1476_),
    .Q(\dut.rd_addr[0] ));
 sg13g2_dfrbp_1 _4149_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net38),
    .D(_0524_),
    .Q_N(_1475_),
    .Q(\dut.rd_addr[1] ));
 sg13g2_dfrbp_1 _4150_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net32),
    .D(_0525_),
    .Q_N(_1474_),
    .Q(\dut.buffer[8] ));
 sg13g2_dfrbp_1 _4151_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net30),
    .D(_0526_),
    .Q_N(_1473_),
    .Q(\dut.buffer[9] ));
 sg13g2_dfrbp_1 _4152_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net28),
    .D(net783),
    .Q_N(_1472_),
    .Q(\dut.buffer[10] ));
 sg13g2_dfrbp_1 _4153_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net19),
    .D(net754),
    .Q_N(_1471_),
    .Q(\dut.buffer[11] ));
 sg13g2_dfrbp_1 _4154_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net607),
    .D(_0529_),
    .Q_N(_1470_),
    .Q(\dut.buffer[12] ));
 sg13g2_dfrbp_1 _4155_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net605),
    .D(_0530_),
    .Q_N(_1469_),
    .Q(\dut.buffer[13] ));
 sg13g2_dfrbp_1 _4156_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net603),
    .D(net821),
    .Q_N(_1468_),
    .Q(\dut.buffer[14] ));
 sg13g2_dfrbp_1 _4157_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net601),
    .D(net762),
    .Q_N(_1467_),
    .Q(\dut.buffer[15] ));
 sg13g2_dfrbp_1 _4158_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net599),
    .D(_0533_),
    .Q_N(_1466_),
    .Q(\dut.din_valid ));
 sg13g2_dfrbp_1 _4159_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net597),
    .D(_0534_),
    .Q_N(_1465_),
    .Q(\dut.din_data[7] ));
 sg13g2_dfrbp_1 _4160_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net437),
    .D(_0535_),
    .Q_N(_1464_),
    .Q(\dut.din_data[6] ));
 sg13g2_dfrbp_1 _4161_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net433),
    .D(_0536_),
    .Q_N(_1463_),
    .Q(\dut.din_data[5] ));
 sg13g2_dfrbp_1 _4162_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net166),
    .D(_0537_),
    .Q_N(_1462_),
    .Q(\dut.din_data[4] ));
 sg13g2_dfrbp_1 _4163_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net158),
    .D(net1168),
    .Q_N(_1461_),
    .Q(\dut.din_data[3] ));
 sg13g2_dfrbp_1 _4164_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net435),
    .D(_0539_),
    .Q_N(_1460_),
    .Q(\dut.din_data[2] ));
 sg13g2_dfrbp_1 _4165_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net162),
    .D(net1173),
    .Q_N(_1459_),
    .Q(\dut.din_data[1] ));
 sg13g2_dfrbp_1 _4166_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net423),
    .D(net1204),
    .Q_N(_1458_),
    .Q(\dut.din_data[0] ));
 sg13g2_tiehi _4153__19 (.L_HI(net19));
 sg13g2_tiehi _4046__20 (.L_HI(net20));
 sg13g2_tiehi _4045__21 (.L_HI(net21));
 sg13g2_tiehi _4044__22 (.L_HI(net22));
 sg13g2_tiehi _4043__23 (.L_HI(net23));
 sg13g2_tiehi _4042__24 (.L_HI(net24));
 sg13g2_tiehi _4041__25 (.L_HI(net25));
 sg13g2_tiehi _4040__26 (.L_HI(net26));
 sg13g2_tiehi _4039__27 (.L_HI(net27));
 sg13g2_tiehi _4152__28 (.L_HI(net28));
 sg13g2_tiehi _4038__29 (.L_HI(net29));
 sg13g2_tiehi _4151__30 (.L_HI(net30));
 sg13g2_tiehi _4037__31 (.L_HI(net31));
 sg13g2_tiehi _4150__32 (.L_HI(net32));
 sg13g2_tiehi _4036__33 (.L_HI(net33));
 sg13g2_tiehi _4035__34 (.L_HI(net34));
 sg13g2_tiehi _4034__35 (.L_HI(net35));
 sg13g2_tiehi _4033__36 (.L_HI(net36));
 sg13g2_tiehi _4032__37 (.L_HI(net37));
 sg13g2_tiehi _4149__38 (.L_HI(net38));
 sg13g2_tiehi _4031__39 (.L_HI(net39));
 sg13g2_tiehi _4030__40 (.L_HI(net40));
 sg13g2_tiehi _4029__41 (.L_HI(net41));
 sg13g2_tiehi _4028__42 (.L_HI(net42));
 sg13g2_tiehi _4027__43 (.L_HI(net43));
 sg13g2_tiehi _4148__44 (.L_HI(net44));
 sg13g2_tiehi _4026__45 (.L_HI(net45));
 sg13g2_tiehi _4025__46 (.L_HI(net46));
 sg13g2_tiehi _4024__47 (.L_HI(net47));
 sg13g2_tiehi _4023__48 (.L_HI(net48));
 sg13g2_tiehi _4022__49 (.L_HI(net49));
 sg13g2_tiehi _4021__50 (.L_HI(net50));
 sg13g2_tiehi _4020__51 (.L_HI(net51));
 sg13g2_tiehi _4019__52 (.L_HI(net52));
 sg13g2_tiehi _4018__53 (.L_HI(net53));
 sg13g2_tiehi _4017__54 (.L_HI(net54));
 sg13g2_tiehi _4016__55 (.L_HI(net55));
 sg13g2_tiehi _4015__56 (.L_HI(net56));
 sg13g2_tiehi _4014__57 (.L_HI(net57));
 sg13g2_tiehi _4013__58 (.L_HI(net58));
 sg13g2_tiehi _4012__59 (.L_HI(net59));
 sg13g2_tiehi _4011__60 (.L_HI(net60));
 sg13g2_tiehi _4010__61 (.L_HI(net61));
 sg13g2_tiehi _4009__62 (.L_HI(net62));
 sg13g2_tiehi _4008__63 (.L_HI(net63));
 sg13g2_tiehi _4007__64 (.L_HI(net64));
 sg13g2_tiehi _4006__65 (.L_HI(net65));
 sg13g2_tiehi _4005__66 (.L_HI(net66));
 sg13g2_tiehi _4004__67 (.L_HI(net67));
 sg13g2_tiehi _4003__68 (.L_HI(net68));
 sg13g2_tiehi _4002__69 (.L_HI(net69));
 sg13g2_tiehi _4001__70 (.L_HI(net70));
 sg13g2_tiehi _4000__71 (.L_HI(net71));
 sg13g2_tiehi _3999__72 (.L_HI(net72));
 sg13g2_tiehi _3998__73 (.L_HI(net73));
 sg13g2_tiehi _3997__74 (.L_HI(net74));
 sg13g2_tiehi _3996__75 (.L_HI(net75));
 sg13g2_tiehi _3995__76 (.L_HI(net76));
 sg13g2_tiehi _3994__77 (.L_HI(net77));
 sg13g2_tiehi _3993__78 (.L_HI(net78));
 sg13g2_tiehi _3992__79 (.L_HI(net79));
 sg13g2_tiehi _3991__80 (.L_HI(net80));
 sg13g2_tiehi _3990__81 (.L_HI(net81));
 sg13g2_tiehi _3989__82 (.L_HI(net82));
 sg13g2_tiehi _3988__83 (.L_HI(net83));
 sg13g2_tiehi _3987__84 (.L_HI(net84));
 sg13g2_tiehi _3986__85 (.L_HI(net85));
 sg13g2_tiehi _3985__86 (.L_HI(net86));
 sg13g2_tiehi _3984__87 (.L_HI(net87));
 sg13g2_tiehi _3983__88 (.L_HI(net88));
 sg13g2_tiehi _3982__89 (.L_HI(net89));
 sg13g2_tiehi _3981__90 (.L_HI(net90));
 sg13g2_tiehi _3980__91 (.L_HI(net91));
 sg13g2_tiehi _3979__92 (.L_HI(net92));
 sg13g2_tiehi _3978__93 (.L_HI(net93));
 sg13g2_tiehi _3977__94 (.L_HI(net94));
 sg13g2_tiehi _3976__95 (.L_HI(net95));
 sg13g2_tiehi _3975__96 (.L_HI(net96));
 sg13g2_tiehi _3974__97 (.L_HI(net97));
 sg13g2_tiehi _3973__98 (.L_HI(net98));
 sg13g2_tiehi _3972__99 (.L_HI(net99));
 sg13g2_tiehi _3971__100 (.L_HI(net100));
 sg13g2_tiehi _3970__101 (.L_HI(net101));
 sg13g2_tiehi _3969__102 (.L_HI(net102));
 sg13g2_tiehi _3968__103 (.L_HI(net103));
 sg13g2_tiehi _3967__104 (.L_HI(net104));
 sg13g2_tiehi _3966__105 (.L_HI(net105));
 sg13g2_tiehi _3965__106 (.L_HI(net106));
 sg13g2_tiehi _3964__107 (.L_HI(net107));
 sg13g2_tiehi _3963__108 (.L_HI(net108));
 sg13g2_tiehi _3962__109 (.L_HI(net109));
 sg13g2_tiehi _3961__110 (.L_HI(net110));
 sg13g2_tiehi _3960__111 (.L_HI(net111));
 sg13g2_tiehi _3959__112 (.L_HI(net112));
 sg13g2_tiehi _3957__113 (.L_HI(net113));
 sg13g2_tiehi _3956__114 (.L_HI(net114));
 sg13g2_tiehi _3955__115 (.L_HI(net115));
 sg13g2_tiehi _3954__116 (.L_HI(net116));
 sg13g2_tiehi _3953__117 (.L_HI(net117));
 sg13g2_tiehi _3952__118 (.L_HI(net118));
 sg13g2_tiehi _3951__119 (.L_HI(net119));
 sg13g2_tiehi _3950__120 (.L_HI(net120));
 sg13g2_tiehi _3949__121 (.L_HI(net121));
 sg13g2_tiehi _3948__122 (.L_HI(net122));
 sg13g2_tiehi _3947__123 (.L_HI(net123));
 sg13g2_tiehi _3946__124 (.L_HI(net124));
 sg13g2_tiehi _3945__125 (.L_HI(net125));
 sg13g2_tiehi _3944__126 (.L_HI(net126));
 sg13g2_tiehi _3943__127 (.L_HI(net127));
 sg13g2_tiehi _3942__128 (.L_HI(net128));
 sg13g2_tiehi _3941__129 (.L_HI(net129));
 sg13g2_tiehi _3940__130 (.L_HI(net130));
 sg13g2_tiehi _3939__131 (.L_HI(net131));
 sg13g2_tiehi _3938__132 (.L_HI(net132));
 sg13g2_tiehi _3937__133 (.L_HI(net133));
 sg13g2_tiehi _3936__134 (.L_HI(net134));
 sg13g2_tiehi _3935__135 (.L_HI(net135));
 sg13g2_tiehi _3934__136 (.L_HI(net136));
 sg13g2_tiehi _3933__137 (.L_HI(net137));
 sg13g2_tiehi _3932__138 (.L_HI(net138));
 sg13g2_tiehi _3931__139 (.L_HI(net139));
 sg13g2_tiehi _3930__140 (.L_HI(net140));
 sg13g2_tiehi _3929__141 (.L_HI(net141));
 sg13g2_tiehi _4147__142 (.L_HI(net142));
 sg13g2_tiehi _3928__143 (.L_HI(net143));
 sg13g2_tiehi _4146__144 (.L_HI(net144));
 sg13g2_tiehi _3925__145 (.L_HI(net145));
 sg13g2_tiehi _4145__146 (.L_HI(net146));
 sg13g2_tiehi _3924__147 (.L_HI(net147));
 sg13g2_tiehi _4144__148 (.L_HI(net148));
 sg13g2_tiehi _3923__149 (.L_HI(net149));
 sg13g2_tiehi _4143__150 (.L_HI(net150));
 sg13g2_tiehi _3922__151 (.L_HI(net151));
 sg13g2_tiehi _4142__152 (.L_HI(net152));
 sg13g2_tiehi _3921__153 (.L_HI(net153));
 sg13g2_tiehi _4141__154 (.L_HI(net154));
 sg13g2_tiehi _3920__155 (.L_HI(net155));
 sg13g2_tiehi _4140__156 (.L_HI(net156));
 sg13g2_tiehi _3919__157 (.L_HI(net157));
 sg13g2_tiehi _4163__158 (.L_HI(net158));
 sg13g2_tiehi _3918__159 (.L_HI(net159));
 sg13g2_tiehi _4139__160 (.L_HI(net160));
 sg13g2_tiehi _3917__161 (.L_HI(net161));
 sg13g2_tiehi _4165__162 (.L_HI(net162));
 sg13g2_tiehi _3916__163 (.L_HI(net163));
 sg13g2_tiehi _4138__164 (.L_HI(net164));
 sg13g2_tiehi _3915__165 (.L_HI(net165));
 sg13g2_tiehi _4162__166 (.L_HI(net166));
 sg13g2_tiehi _3914__167 (.L_HI(net167));
 sg13g2_tiehi _4137__168 (.L_HI(net168));
 sg13g2_tiehi _3913__169 (.L_HI(net169));
 sg13g2_tiehi _4136__170 (.L_HI(net170));
 sg13g2_tiehi _3912__171 (.L_HI(net171));
 sg13g2_tiehi _4135__172 (.L_HI(net172));
 sg13g2_tiehi _3911__173 (.L_HI(net173));
 sg13g2_tiehi _4134__174 (.L_HI(net174));
 sg13g2_tiehi _3910__175 (.L_HI(net175));
 sg13g2_tiehi _4133__176 (.L_HI(net176));
 sg13g2_tiehi _3909__177 (.L_HI(net177));
 sg13g2_tiehi _4132__178 (.L_HI(net178));
 sg13g2_tiehi _3908__179 (.L_HI(net179));
 sg13g2_tiehi _4131__180 (.L_HI(net180));
 sg13g2_tiehi _3907__181 (.L_HI(net181));
 sg13g2_tiehi _4130__182 (.L_HI(net182));
 sg13g2_tiehi _3906__183 (.L_HI(net183));
 sg13g2_tiehi _4129__184 (.L_HI(net184));
 sg13g2_tiehi _3905__185 (.L_HI(net185));
 sg13g2_tiehi _4128__186 (.L_HI(net186));
 sg13g2_tiehi _3904__187 (.L_HI(net187));
 sg13g2_tiehi _4127__188 (.L_HI(net188));
 sg13g2_tiehi _3699__189 (.L_HI(net189));
 sg13g2_tiehi _3869__190 (.L_HI(net190));
 sg13g2_tiehi _3870__191 (.L_HI(net191));
 sg13g2_tiehi _3871__192 (.L_HI(net192));
 sg13g2_tiehi _3872__193 (.L_HI(net193));
 sg13g2_tiehi _3873__194 (.L_HI(net194));
 sg13g2_tiehi _3874__195 (.L_HI(net195));
 sg13g2_tiehi _3875__196 (.L_HI(net196));
 sg13g2_tiehi _3876__197 (.L_HI(net197));
 sg13g2_tiehi _3877__198 (.L_HI(net198));
 sg13g2_tiehi _3878__199 (.L_HI(net199));
 sg13g2_tiehi _3879__200 (.L_HI(net200));
 sg13g2_tiehi _3880__201 (.L_HI(net201));
 sg13g2_tiehi _3903__202 (.L_HI(net202));
 sg13g2_tiehi _4126__203 (.L_HI(net203));
 sg13g2_tiehi _3902__204 (.L_HI(net204));
 sg13g2_tiehi _4125__205 (.L_HI(net205));
 sg13g2_tiehi _3901__206 (.L_HI(net206));
 sg13g2_tiehi _4124__207 (.L_HI(net207));
 sg13g2_tiehi _3900__208 (.L_HI(net208));
 sg13g2_tiehi _4123__209 (.L_HI(net209));
 sg13g2_tiehi _3899__210 (.L_HI(net210));
 sg13g2_tiehi _4122__211 (.L_HI(net211));
 sg13g2_tiehi _3898__212 (.L_HI(net212));
 sg13g2_tiehi _3881__213 (.L_HI(net213));
 sg13g2_tiehi _4121__214 (.L_HI(net214));
 sg13g2_tiehi _3897__215 (.L_HI(net215));
 sg13g2_tiehi _4120__216 (.L_HI(net216));
 sg13g2_tiehi _3896__217 (.L_HI(net217));
 sg13g2_tiehi _4119__218 (.L_HI(net218));
 sg13g2_tiehi _3895__219 (.L_HI(net219));
 sg13g2_tiehi _3894__220 (.L_HI(net220));
 sg13g2_tiehi _3892__221 (.L_HI(net221));
 sg13g2_tiehi _3891__222 (.L_HI(net222));
 sg13g2_tiehi _3890__223 (.L_HI(net223));
 sg13g2_tiehi _3889__224 (.L_HI(net224));
 sg13g2_tiehi _4118__225 (.L_HI(net225));
 sg13g2_tiehi _3888__226 (.L_HI(net226));
 sg13g2_tiehi _4117__227 (.L_HI(net227));
 sg13g2_tiehi _3887__228 (.L_HI(net228));
 sg13g2_tiehi _4116__229 (.L_HI(net229));
 sg13g2_tiehi _3886__230 (.L_HI(net230));
 sg13g2_tiehi _4115__231 (.L_HI(net231));
 sg13g2_tiehi _3885__232 (.L_HI(net232));
 sg13g2_tiehi _4114__233 (.L_HI(net233));
 sg13g2_tiehi _3884__234 (.L_HI(net234));
 sg13g2_tiehi _3883__235 (.L_HI(net235));
 sg13g2_tiehi _4113__236 (.L_HI(net236));
 sg13g2_tiehi _3882__237 (.L_HI(net237));
 sg13g2_tiehi _4112__238 (.L_HI(net238));
 sg13g2_tiehi _3868__239 (.L_HI(net239));
 sg13g2_tiehi _4111__240 (.L_HI(net240));
 sg13g2_tiehi _3867__241 (.L_HI(net241));
 sg13g2_tiehi _3866__242 (.L_HI(net242));
 sg13g2_tiehi _3865__243 (.L_HI(net243));
 sg13g2_tiehi _3864__244 (.L_HI(net244));
 sg13g2_tiehi _3863__245 (.L_HI(net245));
 sg13g2_tiehi _3893__246 (.L_HI(net246));
 sg13g2_tiehi _3926__247 (.L_HI(net247));
 sg13g2_tiehi _3862__248 (.L_HI(net248));
 sg13g2_tiehi _3861__249 (.L_HI(net249));
 sg13g2_tiehi _3860__250 (.L_HI(net250));
 sg13g2_tiehi _3859__251 (.L_HI(net251));
 sg13g2_tiehi _3858__252 (.L_HI(net252));
 sg13g2_tiehi _3857__253 (.L_HI(net253));
 sg13g2_tiehi _3856__254 (.L_HI(net254));
 sg13g2_tiehi _3855__255 (.L_HI(net255));
 sg13g2_tiehi _3854__256 (.L_HI(net256));
 sg13g2_tiehi _3853__257 (.L_HI(net257));
 sg13g2_tiehi _3852__258 (.L_HI(net258));
 sg13g2_tiehi _3851__259 (.L_HI(net259));
 sg13g2_tiehi _3850__260 (.L_HI(net260));
 sg13g2_tiehi _3849__261 (.L_HI(net261));
 sg13g2_tiehi _3848__262 (.L_HI(net262));
 sg13g2_tiehi _3847__263 (.L_HI(net263));
 sg13g2_tiehi _3846__264 (.L_HI(net264));
 sg13g2_tiehi _3845__265 (.L_HI(net265));
 sg13g2_tiehi _3844__266 (.L_HI(net266));
 sg13g2_tiehi _3843__267 (.L_HI(net267));
 sg13g2_tiehi _3842__268 (.L_HI(net268));
 sg13g2_tiehi _3841__269 (.L_HI(net269));
 sg13g2_tiehi _3840__270 (.L_HI(net270));
 sg13g2_tiehi _3839__271 (.L_HI(net271));
 sg13g2_tiehi _3838__272 (.L_HI(net272));
 sg13g2_tiehi _3837__273 (.L_HI(net273));
 sg13g2_tiehi _3836__274 (.L_HI(net274));
 sg13g2_tiehi _3835__275 (.L_HI(net275));
 sg13g2_tiehi _3834__276 (.L_HI(net276));
 sg13g2_tiehi _3833__277 (.L_HI(net277));
 sg13g2_tiehi _3927__278 (.L_HI(net278));
 sg13g2_tiehi _3832__279 (.L_HI(net279));
 sg13g2_tiehi _3831__280 (.L_HI(net280));
 sg13g2_tiehi _3830__281 (.L_HI(net281));
 sg13g2_tiehi _3829__282 (.L_HI(net282));
 sg13g2_tiehi _3828__283 (.L_HI(net283));
 sg13g2_tiehi _3827__284 (.L_HI(net284));
 sg13g2_tiehi _3826__285 (.L_HI(net285));
 sg13g2_tiehi _3825__286 (.L_HI(net286));
 sg13g2_tiehi _3824__287 (.L_HI(net287));
 sg13g2_tiehi _3823__288 (.L_HI(net288));
 sg13g2_tiehi _3822__289 (.L_HI(net289));
 sg13g2_tiehi _3821__290 (.L_HI(net290));
 sg13g2_tiehi _3820__291 (.L_HI(net291));
 sg13g2_tiehi _3819__292 (.L_HI(net292));
 sg13g2_tiehi _3818__293 (.L_HI(net293));
 sg13g2_tiehi _3817__294 (.L_HI(net294));
 sg13g2_tiehi _3816__295 (.L_HI(net295));
 sg13g2_tiehi _3815__296 (.L_HI(net296));
 sg13g2_tiehi _3814__297 (.L_HI(net297));
 sg13g2_tiehi _3813__298 (.L_HI(net298));
 sg13g2_tiehi _3812__299 (.L_HI(net299));
 sg13g2_tiehi _3811__300 (.L_HI(net300));
 sg13g2_tiehi _3810__301 (.L_HI(net301));
 sg13g2_tiehi _3809__302 (.L_HI(net302));
 sg13g2_tiehi _3808__303 (.L_HI(net303));
 sg13g2_tiehi _3807__304 (.L_HI(net304));
 sg13g2_tiehi _3806__305 (.L_HI(net305));
 sg13g2_tiehi _3805__306 (.L_HI(net306));
 sg13g2_tiehi _3804__307 (.L_HI(net307));
 sg13g2_tiehi _3803__308 (.L_HI(net308));
 sg13g2_tiehi _3802__309 (.L_HI(net309));
 sg13g2_tiehi _3801__310 (.L_HI(net310));
 sg13g2_tiehi _3800__311 (.L_HI(net311));
 sg13g2_tiehi _3799__312 (.L_HI(net312));
 sg13g2_tiehi _3798__313 (.L_HI(net313));
 sg13g2_tiehi _3797__314 (.L_HI(net314));
 sg13g2_tiehi _3796__315 (.L_HI(net315));
 sg13g2_tiehi _3795__316 (.L_HI(net316));
 sg13g2_tiehi _3794__317 (.L_HI(net317));
 sg13g2_tiehi _3793__318 (.L_HI(net318));
 sg13g2_tiehi _3792__319 (.L_HI(net319));
 sg13g2_tiehi _3791__320 (.L_HI(net320));
 sg13g2_tiehi _3790__321 (.L_HI(net321));
 sg13g2_tiehi _3789__322 (.L_HI(net322));
 sg13g2_tiehi _3788__323 (.L_HI(net323));
 sg13g2_tiehi _3787__324 (.L_HI(net324));
 sg13g2_tiehi _3786__325 (.L_HI(net325));
 sg13g2_tiehi _3785__326 (.L_HI(net326));
 sg13g2_tiehi _3784__327 (.L_HI(net327));
 sg13g2_tiehi _3783__328 (.L_HI(net328));
 sg13g2_tiehi _3782__329 (.L_HI(net329));
 sg13g2_tiehi _3781__330 (.L_HI(net330));
 sg13g2_tiehi _3780__331 (.L_HI(net331));
 sg13g2_tiehi _3779__332 (.L_HI(net332));
 sg13g2_tiehi _3778__333 (.L_HI(net333));
 sg13g2_tiehi _3777__334 (.L_HI(net334));
 sg13g2_tiehi _3776__335 (.L_HI(net335));
 sg13g2_tiehi _3775__336 (.L_HI(net336));
 sg13g2_tiehi _3774__337 (.L_HI(net337));
 sg13g2_tiehi _3773__338 (.L_HI(net338));
 sg13g2_tiehi _3772__339 (.L_HI(net339));
 sg13g2_tiehi _3771__340 (.L_HI(net340));
 sg13g2_tiehi _3770__341 (.L_HI(net341));
 sg13g2_tiehi _3769__342 (.L_HI(net342));
 sg13g2_tiehi _3768__343 (.L_HI(net343));
 sg13g2_tiehi _3767__344 (.L_HI(net344));
 sg13g2_tiehi _3766__345 (.L_HI(net345));
 sg13g2_tiehi _3765__346 (.L_HI(net346));
 sg13g2_tiehi _3764__347 (.L_HI(net347));
 sg13g2_tiehi _3763__348 (.L_HI(net348));
 sg13g2_tiehi _3762__349 (.L_HI(net349));
 sg13g2_tiehi _3761__350 (.L_HI(net350));
 sg13g2_tiehi _3760__351 (.L_HI(net351));
 sg13g2_tiehi _3759__352 (.L_HI(net352));
 sg13g2_tiehi _3758__353 (.L_HI(net353));
 sg13g2_tiehi _3757__354 (.L_HI(net354));
 sg13g2_tiehi _3756__355 (.L_HI(net355));
 sg13g2_tiehi _3755__356 (.L_HI(net356));
 sg13g2_tiehi _3754__357 (.L_HI(net357));
 sg13g2_tiehi _3753__358 (.L_HI(net358));
 sg13g2_tiehi _3752__359 (.L_HI(net359));
 sg13g2_tiehi _3751__360 (.L_HI(net360));
 sg13g2_tiehi _3750__361 (.L_HI(net361));
 sg13g2_tiehi _3749__362 (.L_HI(net362));
 sg13g2_tiehi _3748__363 (.L_HI(net363));
 sg13g2_tiehi _3747__364 (.L_HI(net364));
 sg13g2_tiehi _3746__365 (.L_HI(net365));
 sg13g2_tiehi _3745__366 (.L_HI(net366));
 sg13g2_tiehi _3744__367 (.L_HI(net367));
 sg13g2_tiehi _3743__368 (.L_HI(net368));
 sg13g2_tiehi _3742__369 (.L_HI(net369));
 sg13g2_tiehi _3741__370 (.L_HI(net370));
 sg13g2_tiehi _3740__371 (.L_HI(net371));
 sg13g2_tiehi _3739__372 (.L_HI(net372));
 sg13g2_tiehi _3738__373 (.L_HI(net373));
 sg13g2_tiehi _4110__374 (.L_HI(net374));
 sg13g2_tiehi _3737__375 (.L_HI(net375));
 sg13g2_tiehi _4109__376 (.L_HI(net376));
 sg13g2_tiehi _3736__377 (.L_HI(net377));
 sg13g2_tiehi _4108__378 (.L_HI(net378));
 sg13g2_tiehi _3735__379 (.L_HI(net379));
 sg13g2_tiehi _4107__380 (.L_HI(net380));
 sg13g2_tiehi _3734__381 (.L_HI(net381));
 sg13g2_tiehi _4106__382 (.L_HI(net382));
 sg13g2_tiehi _3733__383 (.L_HI(net383));
 sg13g2_tiehi _3732__384 (.L_HI(net384));
 sg13g2_tiehi _3731__385 (.L_HI(net385));
 sg13g2_tiehi _3730__386 (.L_HI(net386));
 sg13g2_tiehi _3729__387 (.L_HI(net387));
 sg13g2_tiehi _3728__388 (.L_HI(net388));
 sg13g2_tiehi _3727__389 (.L_HI(net389));
 sg13g2_tiehi _3726__390 (.L_HI(net390));
 sg13g2_tiehi _3725__391 (.L_HI(net391));
 sg13g2_tiehi _3724__392 (.L_HI(net392));
 sg13g2_tiehi _3723__393 (.L_HI(net393));
 sg13g2_tiehi _3722__394 (.L_HI(net394));
 sg13g2_tiehi _3721__395 (.L_HI(net395));
 sg13g2_tiehi _3720__396 (.L_HI(net396));
 sg13g2_tiehi _3958__397 (.L_HI(net397));
 sg13g2_tiehi _4077__398 (.L_HI(net398));
 sg13g2_tiehi _4078__399 (.L_HI(net399));
 sg13g2_tiehi _3719__400 (.L_HI(net400));
 sg13g2_tiehi _3718__401 (.L_HI(net401));
 sg13g2_tiehi _3717__402 (.L_HI(net402));
 sg13g2_tiehi _3716__403 (.L_HI(net403));
 sg13g2_tiehi _3715__404 (.L_HI(net404));
 sg13g2_tiehi _3714__405 (.L_HI(net405));
 sg13g2_tiehi _3713__406 (.L_HI(net406));
 sg13g2_tiehi _3712__407 (.L_HI(net407));
 sg13g2_tiehi _3711__408 (.L_HI(net408));
 sg13g2_tiehi _3710__409 (.L_HI(net409));
 sg13g2_tiehi _3709__410 (.L_HI(net410));
 sg13g2_tiehi _3708__411 (.L_HI(net411));
 sg13g2_tiehi _3707__412 (.L_HI(net412));
 sg13g2_tiehi _3706__413 (.L_HI(net413));
 sg13g2_tiehi _3705__414 (.L_HI(net414));
 sg13g2_tiehi _3704__415 (.L_HI(net415));
 sg13g2_tiehi _3703__416 (.L_HI(net416));
 sg13g2_tiehi _3702__417 (.L_HI(net417));
 sg13g2_tiehi _3701__418 (.L_HI(net418));
 sg13g2_tiehi _3700__419 (.L_HI(net419));
 sg13g2_tiehi _4105__420 (.L_HI(net420));
 sg13g2_tiehi _4104__421 (.L_HI(net421));
 sg13g2_tiehi _4103__422 (.L_HI(net422));
 sg13g2_tiehi _4166__423 (.L_HI(net423));
 sg13g2_tiehi _4102__424 (.L_HI(net424));
 sg13g2_tiehi _4101__425 (.L_HI(net425));
 sg13g2_tiehi _4100__426 (.L_HI(net426));
 sg13g2_tiehi _4099__427 (.L_HI(net427));
 sg13g2_tiehi _4098__428 (.L_HI(net428));
 sg13g2_tiehi _4097__429 (.L_HI(net429));
 sg13g2_tiehi _4096__430 (.L_HI(net430));
 sg13g2_tiehi _4095__431 (.L_HI(net431));
 sg13g2_tiehi _4094__432 (.L_HI(net432));
 sg13g2_tiehi _4161__433 (.L_HI(net433));
 sg13g2_tiehi _4093__434 (.L_HI(net434));
 sg13g2_tiehi _4164__435 (.L_HI(net435));
 sg13g2_tiehi _4092__436 (.L_HI(net436));
 sg13g2_tiehi _4160__437 (.L_HI(net437));
 sg13g2_tiehi _4091__438 (.L_HI(net438));
 sg13g2_tiehi _4090__439 (.L_HI(net439));
 sg13g2_tiehi _4089__440 (.L_HI(net440));
 sg13g2_tiehi _4088__441 (.L_HI(net587));
 sg13g2_tiehi _4087__442 (.L_HI(net588));
 sg13g2_tiehi _4086__443 (.L_HI(net589));
 sg13g2_tiehi _4085__444 (.L_HI(net590));
 sg13g2_tiehi _4084__445 (.L_HI(net591));
 sg13g2_tiehi _4083__446 (.L_HI(net592));
 sg13g2_tiehi _4082__447 (.L_HI(net593));
 sg13g2_tiehi _4081__448 (.L_HI(net594));
 sg13g2_tiehi _4079__449 (.L_HI(net595));
 sg13g2_tiehi _4080__450 (.L_HI(net596));
 sg13g2_tiehi _4159__451 (.L_HI(net597));
 sg13g2_tiehi _4076__452 (.L_HI(net598));
 sg13g2_tiehi _4158__453 (.L_HI(net599));
 sg13g2_tiehi _4075__454 (.L_HI(net600));
 sg13g2_tiehi _4157__455 (.L_HI(net601));
 sg13g2_tiehi _4074__456 (.L_HI(net602));
 sg13g2_tiehi _4156__457 (.L_HI(net603));
 sg13g2_tiehi _4073__458 (.L_HI(net604));
 sg13g2_tiehi _4155__459 (.L_HI(net605));
 sg13g2_tiehi _4072__460 (.L_HI(net606));
 sg13g2_tiehi _4154__461 (.L_HI(net607));
 sg13g2_tiehi _4071__462 (.L_HI(net608));
 sg13g2_tiehi _4070__463 (.L_HI(net609));
 sg13g2_tiehi _4069__464 (.L_HI(net610));
 sg13g2_tiehi _4068__465 (.L_HI(net611));
 sg13g2_tiehi _4067__466 (.L_HI(net612));
 sg13g2_tiehi _4066__467 (.L_HI(net613));
 sg13g2_tiehi _4065__468 (.L_HI(net614));
 sg13g2_tiehi _4064__469 (.L_HI(net615));
 sg13g2_tiehi _4063__470 (.L_HI(net616));
 sg13g2_tiehi _4062__471 (.L_HI(net617));
 sg13g2_tiehi _4061__472 (.L_HI(net618));
 sg13g2_tiehi _4060__473 (.L_HI(net619));
 sg13g2_tiehi _4059__474 (.L_HI(net620));
 sg13g2_tiehi _4058__475 (.L_HI(net621));
 sg13g2_tiehi _4057__476 (.L_HI(net622));
 sg13g2_tiehi _4056__477 (.L_HI(net623));
 sg13g2_tiehi _4055__478 (.L_HI(net624));
 sg13g2_tiehi _4054__479 (.L_HI(net625));
 sg13g2_tiehi _4053__480 (.L_HI(net626));
 sg13g2_tiehi _4052__481 (.L_HI(net627));
 sg13g2_tiehi _4051__482 (.L_HI(net628));
 sg13g2_tiehi _4050__483 (.L_HI(net629));
 sg13g2_tiehi _4049__484 (.L_HI(net630));
 sg13g2_tiehi _4048__485 (.L_HI(net631));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_underserved_3 (.L_LO(net3));
 sg13g2_tielo tt_um_underserved_4 (.L_LO(net4));
 sg13g2_tielo tt_um_underserved_5 (.L_LO(net5));
 sg13g2_tielo tt_um_underserved_6 (.L_LO(net6));
 sg13g2_tielo tt_um_underserved_7 (.L_LO(net7));
 sg13g2_tielo tt_um_underserved_8 (.L_LO(net8));
 sg13g2_tielo tt_um_underserved_9 (.L_LO(net9));
 sg13g2_tielo tt_um_underserved_10 (.L_LO(net10));
 sg13g2_tielo tt_um_underserved_11 (.L_LO(net11));
 sg13g2_tielo tt_um_underserved_12 (.L_LO(net12));
 sg13g2_tielo tt_um_underserved_13 (.L_LO(net13));
 sg13g2_tielo tt_um_underserved_14 (.L_LO(net14));
 sg13g2_tielo tt_um_underserved_15 (.L_LO(net15));
 sg13g2_tielo tt_um_underserved_16 (.L_LO(net16));
 sg13g2_tielo tt_um_underserved_17 (.L_LO(net17));
 sg13g2_tiehi _4047__18 (.L_HI(net18));
 sg13g2_buf_1 _4651_ (.A(net567),
    .X(uo_out[5]));
 sg13g2_buf_1 _4652_ (.A(\dut.flash_csb ),
    .X(uo_out[6]));
 sg13g2_buf_1 _4653_ (.A(\dut.flash_io0_do ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout441 (.A(_0829_),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(net443),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_1424_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(net447),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(net446),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(net447),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(net448),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(net457),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(net451),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(net451),
    .X(net450));
 sg13g2_buf_4 fanout451 (.X(net451),
    .A(net457));
 sg13g2_buf_4 fanout452 (.X(net452),
    .A(net457));
 sg13g2_buf_2 fanout453 (.A(net457),
    .X(net453));
 sg13g2_buf_4 fanout454 (.X(net454),
    .A(net456));
 sg13g2_buf_2 fanout455 (.A(net456),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(net457),
    .X(net456));
 sg13g2_buf_4 fanout457 (.X(net457),
    .A(_1295_));
 sg13g2_buf_2 fanout458 (.A(_1270_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(_1270_),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(net461),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(net470),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(net470),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(net464),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(net469),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(net466),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(net467),
    .X(net466));
 sg13g2_buf_1 fanout467 (.A(net468),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(net469),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(net470),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_1147_),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(net473),
    .X(net471));
 sg13g2_buf_4 fanout472 (.X(net472),
    .A(net473));
 sg13g2_buf_2 fanout473 (.A(net481),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(net476),
    .X(net474));
 sg13g2_buf_1 fanout475 (.A(net476),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(net481),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(net478),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(net479),
    .X(net478));
 sg13g2_buf_1 fanout479 (.A(net480),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(net481),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_1143_),
    .X(net481));
 sg13g2_buf_4 fanout482 (.X(net482),
    .A(net483));
 sg13g2_buf_4 fanout483 (.X(net483),
    .A(net484));
 sg13g2_buf_2 fanout484 (.A(_1020_),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(net486),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(net490),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(net488),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(net489),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(net490),
    .X(net489));
 sg13g2_buf_4 fanout490 (.X(net490),
    .A(_1020_));
 sg13g2_buf_4 fanout491 (.X(net491),
    .A(net494));
 sg13g2_buf_4 fanout492 (.X(net492),
    .A(net494));
 sg13g2_buf_2 fanout493 (.A(net494),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(net520),
    .X(net494));
 sg13g2_buf_4 fanout495 (.X(net495),
    .A(net499));
 sg13g2_buf_2 fanout496 (.A(net499),
    .X(net496));
 sg13g2_buf_4 fanout497 (.X(net497),
    .A(net499));
 sg13g2_buf_2 fanout498 (.A(net499),
    .X(net498));
 sg13g2_buf_1 fanout499 (.A(net520),
    .X(net499));
 sg13g2_buf_4 fanout500 (.X(net500),
    .A(net501));
 sg13g2_buf_2 fanout501 (.A(net502),
    .X(net501));
 sg13g2_buf_4 fanout502 (.X(net502),
    .A(net520));
 sg13g2_buf_4 fanout503 (.X(net503),
    .A(net506));
 sg13g2_buf_2 fanout504 (.A(net506),
    .X(net504));
 sg13g2_buf_4 fanout505 (.X(net505),
    .A(net506));
 sg13g2_buf_2 fanout506 (.A(net520),
    .X(net506));
 sg13g2_buf_4 fanout507 (.X(net507),
    .A(net508));
 sg13g2_buf_2 fanout508 (.A(net509),
    .X(net508));
 sg13g2_buf_4 fanout509 (.X(net509),
    .A(net520));
 sg13g2_buf_4 fanout510 (.X(net510),
    .A(net514));
 sg13g2_buf_2 fanout511 (.A(net514),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(net513),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(net514),
    .X(net513));
 sg13g2_buf_1 fanout514 (.A(net519),
    .X(net514));
 sg13g2_buf_4 fanout515 (.X(net515),
    .A(net516));
 sg13g2_buf_2 fanout516 (.A(net519),
    .X(net516));
 sg13g2_buf_4 fanout517 (.X(net517),
    .A(net519));
 sg13g2_buf_2 fanout518 (.A(net519),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(net520),
    .X(net519));
 sg13g2_buf_4 fanout520 (.X(net520),
    .A(_0947_));
 sg13g2_buf_2 fanout521 (.A(_0843_),
    .X(net521));
 sg13g2_buf_4 fanout522 (.X(net522),
    .A(net523));
 sg13g2_buf_4 fanout523 (.X(net523),
    .A(_1035_));
 sg13g2_buf_4 fanout524 (.X(net524),
    .A(net526));
 sg13g2_buf_1 fanout525 (.A(net526),
    .X(net525));
 sg13g2_buf_4 fanout526 (.X(net526),
    .A(_1035_));
 sg13g2_buf_2 fanout527 (.A(net528),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(net531),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(net530),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(net531),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(_1034_),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(net533),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(_0828_),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(net538),
    .X(net534));
 sg13g2_buf_1 fanout535 (.A(net538),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(net538),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(net538),
    .X(net537));
 sg13g2_buf_1 fanout538 (.A(_0827_),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(_1148_),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(_1013_),
    .X(net540));
 sg13g2_buf_4 fanout541 (.X(net541),
    .A(net542));
 sg13g2_buf_2 fanout542 (.A(net543),
    .X(net542));
 sg13g2_buf_4 fanout543 (.X(net543),
    .A(_0922_));
 sg13g2_buf_4 fanout544 (.X(net544),
    .A(net546));
 sg13g2_buf_2 fanout545 (.A(net546),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_0922_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(net548),
    .X(net547));
 sg13g2_buf_1 fanout548 (.A(_1086_),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(_0621_),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(_0621_),
    .X(net550));
 sg13g2_buf_4 fanout551 (.X(net551),
    .A(net552));
 sg13g2_buf_4 fanout552 (.X(net552),
    .A(net554));
 sg13g2_buf_4 fanout553 (.X(net553),
    .A(net554));
 sg13g2_buf_2 fanout554 (.A(_0619_),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(net557),
    .X(net555));
 sg13g2_buf_1 fanout556 (.A(net557),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(net1341),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(net834),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(net563),
    .X(net559));
 sg13g2_buf_1 fanout560 (.A(net563),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(net563),
    .X(net561));
 sg13g2_buf_1 fanout562 (.A(net563),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(\dut.rd_inc ),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(net566),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(net566),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(\dut.rd_inc ),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(\dut.flash_clk ),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(net1339),
    .X(net568));
 sg13g2_buf_4 fanout569 (.X(net569),
    .A(\cpu.branch_op ));
 sg13g2_buf_1 fanout570 (.A(\cpu.branch_op ),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(\cpu.bufreg2.i_op_b_sel ),
    .X(net571));
 sg13g2_buf_4 fanout572 (.X(net572),
    .A(\cpu.decode.opcode[2] ));
 sg13g2_buf_2 fanout573 (.A(\cpu.decode.opcode[2] ),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(\cpu.decode.opcode[0] ),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(\cpu.decode.opcode[0] ),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(net1319),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(net1338),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(\dut.state[9] ),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(\dut.state[6] ),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(rst_n),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(rst_n),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(net584),
    .X(net582));
 sg13g2_buf_1 fanout583 (.A(net584),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(net585),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(net586),
    .X(net585));
 sg13g2_buf_4 fanout586 (.X(net586),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[7]),
    .X(net1));
 sg13g2_tielo tt_um_underserved_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_4_7_0_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_4_11_0_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_4_15_0_clk));
 sg13g2_inv_8 clkload3 (.A(clknet_leaf_59_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_leaf_60_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_leaf_20_clk));
 sg13g2_inv_4 clkload6 (.A(clknet_leaf_32_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_36_clk));
 sg13g2_inv_8 clkload8 (.A(clknet_leaf_28_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\dut.xfer.xfer_tag[2] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold2 (.A(\dut.xfer.xfer_tag[1] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold3 (.A(\dut.xfer.xfer_tag[0] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold4 (.A(\rf_shift_reg.rreq_r ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0093_),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0128_),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0019_),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0261_),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold9 (.A(\rf_shift_reg.x[1][4] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0099_),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold11 (.A(\rf_shift_reg.x[1][29] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0124_),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold13 (.A(\rf_shift_reg.x[3][1] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0165_),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold15 (.A(\rf_shift_reg.x[1][1] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0096_),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold17 (.A(\cpu.ctrl.o_ibus_adr[15] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold18 (.A(_1051_),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold19 (.A(\cpu.ctrl.o_ibus_adr[13] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold20 (.A(_1049_),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold21 (.A(\rf_shift_reg.x[4][1] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0197_),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold23 (.A(\dut.buffer[8] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0487_),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold25 (.A(\cpu.ctrl.o_ibus_adr[4] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold26 (.A(_1040_),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold27 (.A(\cpu.bufreg.data[30] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0336_),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold29 (.A(\cpu.ctrl.o_ibus_adr[14] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold30 (.A(\cpu.ctrl.o_ibus_adr[2] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold31 (.A(_1038_),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold32 (.A(\rf_shift_reg.x[2][1] ),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0133_),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold34 (.A(\cpu.ctrl.o_ibus_adr[17] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold35 (.A(_1053_),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold36 (.A(\rf_shift_reg.x[5][1] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0229_),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold38 (.A(\rf_shift_reg.x[5][31] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0260_),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold40 (.A(\cpu.ctrl.o_ibus_adr[12] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold41 (.A(\cpu.bufreg2.dat[18] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0389_),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold43 (.A(\cpu.ctrl.o_ibus_adr[19] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold44 (.A(_1055_),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold45 (.A(\rf_shift_reg.x[4][20] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0216_),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold47 (.A(\rf_shift_reg.x[3][31] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0195_),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold49 (.A(\cpu.ctrl.o_ibus_adr[21] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold50 (.A(_1057_),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold51 (.A(\rf_shift_reg.x[2][30] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0163_),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold53 (.A(\cpu.ctrl.o_ibus_adr[6] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold54 (.A(_1042_),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold55 (.A(\cpu.ctrl.o_ibus_adr[7] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold56 (.A(_1043_),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold57 (.A(\dut.din_tag[0] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0414_),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold59 (.A(\cpu.bufreg2.dat[25] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0396_),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold61 (.A(\cpu.ctrl.o_ibus_adr[8] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold62 (.A(_1044_),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold63 (.A(\cpu.ctrl.o_ibus_adr[29] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold64 (.A(_1065_),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold65 (.A(\cpu.bufreg2.dat[6] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0377_),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold67 (.A(\cpu.bufreg2.dat[14] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0385_),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold69 (.A(\cpu.ctrl.o_ibus_adr[25] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold70 (.A(_1061_),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold71 (.A(\cpu.ctrl.o_ibus_adr[20] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold72 (.A(\rf_shift_reg.x[3][29] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0193_),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold74 (.A(\cpu.bufreg2.dat[20] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0391_),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold76 (.A(\cpu.ctrl.o_ibus_adr[10] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold77 (.A(_1046_),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold78 (.A(\dut.rd_addr[15] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0438_),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold80 (.A(\cpu.ctrl.o_ibus_adr[16] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold81 (.A(\cpu.ctrl.o_ibus_adr[9] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold82 (.A(\cpu.bufreg.data[12] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0317_),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold84 (.A(\dut.rd_addr[23] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0446_),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold86 (.A(\cpu.ctrl.o_ibus_adr[28] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold87 (.A(\cpu.ctrl.o_ibus_adr[22] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold88 (.A(_1058_),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold89 (.A(\dut.state[7] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0007_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold91 (.A(\cpu.ctrl.o_ibus_adr[27] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold92 (.A(\cpu.ctrl.o_ibus_adr[11] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold93 (.A(\cpu.ctrl.o_ibus_adr[5] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold94 (.A(\dut.rd_addr[10] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold95 (.A(\rf_shift_reg.x[3][20] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0184_),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold97 (.A(\cpu.ctrl.o_ibus_adr[30] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold98 (.A(_1066_),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold99 (.A(\rf_shift_reg.x[4][31] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0228_),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold101 (.A(\cpu.ctrl.o_ibus_adr[23] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold102 (.A(_1059_),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold103 (.A(\cpu.ctrl.o_ibus_adr[18] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold104 (.A(\cpu.ctrl.o_ibus_adr[3] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold105 (.A(\dut.buffer[5] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0484_),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold107 (.A(\rf_shift_reg.x[3][18] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0182_),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold109 (.A(\dut.rd_addr[11] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0434_),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold111 (.A(\dut.rd_addr[21] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0444_),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0086_),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0450_),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold115 (.A(\dut.xfer.count[1] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold116 (.A(\dut.buffer[13] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0492_),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold118 (.A(\dut.dout_data[5] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold119 (.A(\rf_shift_reg.x[4][22] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0218_),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold121 (.A(\cpu.ctrl.o_ibus_adr[1] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold122 (.A(\dut.buffer[11] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0528_),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold124 (.A(\dut.rd_addr[17] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0440_),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold126 (.A(\cpu.bufreg2.dat[23] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0394_),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold128 (.A(\cpu.bufreg2.dat[31] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0402_),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold130 (.A(\dut.buffer[15] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0532_),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold132 (.A(\dut.buffer[12] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0491_),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold134 (.A(\dut.din_tag[1] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0415_),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold136 (.A(\dut.rd_addr[12] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0435_),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold138 (.A(\dut.rd_addr[16] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0439_),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold140 (.A(\cpu.state.cnt_r[2] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold141 (.A(\cpu.bufreg2.i_dat[15] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold142 (.A(\cpu.immdec.imm30_25[3] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0354_),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold144 (.A(\cpu.bufreg2.dat[29] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0400_),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold146 (.A(\cpu.ctrl.o_ibus_adr[26] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold147 (.A(\dut.xfer.count[0] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold148 (.A(_1009_),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold149 (.A(\cpu.bufreg2.dat[27] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0398_),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold151 (.A(\dut.buffer[10] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0527_),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold153 (.A(\cpu.bufreg2.dat[22] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0393_),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold155 (.A(\cpu.bufreg2.dat[12] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0383_),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold157 (.A(\dut.dout_data[4] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold158 (.A(\cpu.bufreg2.i_dat[11] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold159 (.A(\rf_shift_reg.x[3][26] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0190_),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold161 (.A(\rf_shift_reg.x[1][23] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0118_),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold163 (.A(\dut.state[0] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold164 (.A(\cpu.immdec.imm30_25[5] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0356_),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold166 (.A(\cpu.immdec.imm30_25[2] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0353_),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold168 (.A(\cpu.mem_if.signbit ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0967_),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold170 (.A(\dut.dout_data[0] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold171 (.A(\rf_shift_reg.x[3][22] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0186_),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold173 (.A(\dut.din_tag[2] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold174 (.A(_1416_),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0514_),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold176 (.A(\cpu.immdec.imm30_25[4] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0355_),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold178 (.A(\dut.xfer.count[2] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold179 (.A(_1012_),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold180 (.A(\rf_shift_reg.x[5][20] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0248_),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold182 (.A(\cpu.bufreg2.dat[10] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0381_),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold184 (.A(\dut.rd_addr[22] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0445_),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold186 (.A(\rf_shift_reg.x[2][4] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0136_),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold188 (.A(\cpu.state.cnt_r[1] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold189 (.A(\dut.buffer[14] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0531_),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold191 (.A(\dut.xfer.next_obuffer[4] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0419_),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold193 (.A(\cpu.immdec.imm30_25[1] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0352_),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold195 (.A(\rf_shift_reg.cnt[1] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0981_),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0129_),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold198 (.A(\cpu.bufreg2.i_dat[14] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold199 (.A(\rf_shift_reg.x[2][29] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0161_),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold201 (.A(\rf_shift_reg.x[4][24] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0220_),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold203 (.A(\dut.xfer.resetn ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold204 (.A(\dut.buffer[2] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0481_),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold206 (.A(\dut.buffer[3] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0482_),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold208 (.A(\dut.rd_addr[8] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0431_),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold210 (.A(\dut.rd_addr[18] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0441_),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold212 (.A(\dut.rd_addr[19] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0442_),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold214 (.A(\dut.rd_addr[9] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0432_),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold216 (.A(\rf_shift_reg.x[5][9] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0237_),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold218 (.A(\dut.rd_addr[20] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0443_),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold220 (.A(\cpu.bufreg2.i_dat[10] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold221 (.A(\rf_shift_reg.x[1][31] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0126_),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold223 (.A(\dut.state[8] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0008_),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold225 (.A(\rf_shift_reg.x[5][12] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0240_),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold227 (.A(\cpu.ctrl.o_ibus_adr[24] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold228 (.A(\rf_shift_reg.x[4][8] ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0204_),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold230 (.A(\dut.xfer.next_obuffer[1] ),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0424_),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold232 (.A(\rf_shift_reg.x[2][16] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0148_),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold234 (.A(\rf_shift_reg.x[4][18] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0214_),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold236 (.A(\rf_shift_reg.x[1][14] ),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0109_),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold238 (.A(\cpu.immdec.imm19_12_20[8] ),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0348_),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold240 (.A(\rf_shift_reg.x[5][26] ),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0254_),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold242 (.A(\dut.buffer[0] ),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0479_),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold244 (.A(\cpu.bufreg.data[6] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0311_),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold246 (.A(\dut.xfer.obuffer[7] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0423_),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold248 (.A(\dut.xfer.next_obuffer[6] ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0421_),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold250 (.A(\dut.din_data[6] ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold251 (.A(\rf_shift_reg.x[3][14] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0178_),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold253 (.A(\dut.rd_addr[4] ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0427_),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold255 (.A(\rf_shift_reg.x[1][7] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0102_),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold257 (.A(\cpu.bufreg.data[24] ),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0329_),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold259 (.A(\rf_shift_reg.x[2][23] ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0155_),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold261 (.A(\rf_shift_reg.x[4][9] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold262 (.A(\rf_shift_reg.x[2][24] ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold263 (.A(\dut.buffer[9] ),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0488_),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold265 (.A(\rf_shift_reg.x[5][22] ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0250_),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold267 (.A(\dut.rd_addr[13] ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0436_),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold269 (.A(\dut.buffer[20] ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0499_),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold271 (.A(\rf_shift_reg.x[4][27] ),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold272 (.A(_0223_),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold273 (.A(\rf_shift_reg.x[1][25] ),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0120_),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold275 (.A(\dut.buffer[16] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0495_),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold277 (.A(\rf_shift_reg.x[5][8] ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0236_),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold279 (.A(\rf_shift_reg.x[1][22] ),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0117_),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold281 (.A(\rf_shift_reg.x[2][20] ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0152_),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold283 (.A(\rf_shift_reg.x[1][11] ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold284 (.A(_0106_),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold285 (.A(\rf_shift_reg.x[1][27] ),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0122_),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold287 (.A(\rf_shift_reg.x[5][30] ),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0258_),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold289 (.A(\cpu.bufreg.data[13] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold290 (.A(\dut.rd_addr[5] ),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0428_),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold292 (.A(\rf_shift_reg.x[5][4] ),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0232_),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold294 (.A(\rf_shift_reg.x[1][6] ),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0101_),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold296 (.A(\dut.buffer[7] ),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold297 (.A(_0486_),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold298 (.A(\cpu.bufreg2.dat[15] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold299 (.A(_0386_),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold300 (.A(\cpu.bufreg.data[26] ),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0331_),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold302 (.A(\rf_shift_reg.x[2][9] ),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0141_),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold304 (.A(\rf_shift_reg.x[4][7] ),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0203_),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold306 (.A(\dut.buffer[17] ),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold307 (.A(_0496_),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold308 (.A(\cpu.bufreg.data[29] ),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold309 (.A(\cpu.bufreg.data[15] ),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold310 (.A(_0320_),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold311 (.A(\rf_shift_reg.x[5][24] ),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0252_),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold313 (.A(\rf_shift_reg.x[5][3] ),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0231_),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold315 (.A(\rf_shift_reg.x[4][2] ),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold316 (.A(\dut.dout_data[1] ),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold317 (.A(\rf_shift_reg.x[5][25] ),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold318 (.A(\rf_shift_reg.x[1][16] ),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold319 (.A(_0111_),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold320 (.A(\rf_shift_reg.x[5][15] ),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold321 (.A(_0243_),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold322 (.A(\rf_shift_reg.x[3][6] ),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0170_),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold324 (.A(\rf_shift_reg.x[4][12] ),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold325 (.A(_0208_),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold326 (.A(\rf_shift_reg.x[1][18] ),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold327 (.A(_0113_),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold328 (.A(\rf_shift_reg.x[2][17] ),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold329 (.A(\rf_shift_reg.x[4][30] ),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold330 (.A(_0226_),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold331 (.A(\rf_shift_reg.x[1][30] ),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold332 (.A(\rf_shift_reg.x[5][2] ),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold333 (.A(\rf_shift_reg.x[4][16] ),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold334 (.A(_0212_),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold335 (.A(\rf_shift_reg.x[5][7] ),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold336 (.A(_0235_),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold337 (.A(\rf_shift_reg.x[3][11] ),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold338 (.A(_0175_),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold339 (.A(\rf_shift_reg.x[5][27] ),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold340 (.A(\dut.rd_addr[7] ),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold341 (.A(_0430_),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold342 (.A(\rf_shift_reg.x[3][23] ),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold343 (.A(\rf_shift_reg.x[2][18] ),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold344 (.A(\rf_shift_reg.x[1][19] ),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold345 (.A(\cpu.bufreg.data[21] ),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold346 (.A(_0326_),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold347 (.A(\cpu.bufreg.c_r ),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold348 (.A(\rf_shift_reg.x[2][15] ),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold349 (.A(_0147_),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold350 (.A(\rf_shift_reg.x[2][12] ),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0144_),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold352 (.A(\dut.buffer[18] ),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold353 (.A(_0471_),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold354 (.A(\rf_shift_reg.x[4][15] ),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0211_),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold356 (.A(\dut.xfer.next_obuffer[3] ),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0418_),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold358 (.A(\dut.buffer[4] ),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0483_),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold360 (.A(\rf_shift_reg.x[5][21] ),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold361 (.A(\rf_shift_reg.x[3][9] ),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0173_),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold363 (.A(\rf_shift_reg.x[2][19] ),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold364 (.A(\cpu.immdec.imm31 ),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold365 (.A(_0340_),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold366 (.A(\rf_shift_reg.x[4][26] ),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0222_),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold368 (.A(\rf_shift_reg.x[2][13] ),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold369 (.A(\rf_shift_reg.x[3][16] ),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0180_),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold371 (.A(\rf_shift_reg.x[4][13] ),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold372 (.A(\rf_shift_reg.x[1][24] ),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold373 (.A(\rf_shift_reg.x[1][20] ),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold374 (.A(\rf_shift_reg.x[5][19] ),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold375 (.A(_0247_),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold376 (.A(\rf_shift_reg.x[2][3] ),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold377 (.A(_0135_),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold378 (.A(\dut.buffer[23] ),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold379 (.A(_0502_),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold380 (.A(\cpu.bufreg.data[19] ),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold381 (.A(_0324_),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold382 (.A(\rf_shift_reg.x[1][9] ),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold383 (.A(_0104_),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold384 (.A(\dut.dout_data[7] ),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold385 (.A(\dut.buffer[1] ),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold386 (.A(_0480_),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold387 (.A(\rf_shift_reg.x[2][6] ),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold388 (.A(_0138_),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold389 (.A(\rf_shift_reg.x[2][27] ),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold390 (.A(_0159_),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold391 (.A(\dut.dout_tag[1] ),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold392 (.A(\rf_shift_reg.x[5][5] ),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold393 (.A(\rf_shift_reg.x[2][26] ),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold394 (.A(_0158_),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold395 (.A(\cpu.bufreg.data[7] ),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold396 (.A(\rf_shift_reg.x[3][17] ),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold397 (.A(\rf_shift_reg.x[1][2] ),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold398 (.A(_0098_),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold399 (.A(\rf_shift_reg.x[4][10] ),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold400 (.A(\rf_shift_reg.x[3][2] ),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold401 (.A(\dut.rd_addr[0] ),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold402 (.A(\dut.buffer[6] ),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold403 (.A(_0485_),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold404 (.A(\rf_shift_reg.x[1][17] ),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold405 (.A(\rf_shift_reg.x[5][18] ),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold406 (.A(_0246_),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold407 (.A(\rf_shift_reg.x[3][10] ),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold408 (.A(\rf_shift_reg.x[3][7] ),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold409 (.A(\rf_shift_reg.x[4][6] ),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold410 (.A(_0202_),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold411 (.A(\cpu.bufreg.data[16] ),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold412 (.A(\cpu.bufreg.data[14] ),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold413 (.A(\rf_shift_reg.x[5][13] ),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold414 (.A(\rf_shift_reg.x[3][8] ),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold415 (.A(\cpu.bufreg2.i_dat[18] ),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold416 (.A(\cpu.bufreg.data[17] ),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold417 (.A(\cpu.bufreg.data[10] ),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold418 (.A(_0315_),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold419 (.A(\rf_shift_reg.x[3][27] ),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold420 (.A(\cpu.immdec.imm24_20[4] ),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold421 (.A(_0360_),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold422 (.A(\rf_shift_reg.x[5][17] ),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0245_),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold424 (.A(\dut.xfer.next_obuffer[5] ),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold425 (.A(_0420_),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold426 (.A(\cpu.bufreg2.i_dat[9] ),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold427 (.A(_0380_),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold428 (.A(\cpu.ctrl.o_ibus_adr[31] ),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold429 (.A(_0307_),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold430 (.A(\cpu.bufreg.data[11] ),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold431 (.A(\cpu.bufreg.data[18] ),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold432 (.A(\rf_shift_reg.x[1][10] ),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold433 (.A(\rf_shift_reg.x[1][13] ),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold434 (.A(_0108_),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold435 (.A(\rf_shift_reg.x[4][5] ),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold436 (.A(_0201_),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold437 (.A(\rf_shift_reg.x[5][23] ),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold438 (.A(\cpu.bufreg2.dat[21] ),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold439 (.A(_0392_),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold440 (.A(\rf_shift_reg.x[3][19] ),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold441 (.A(\cpu.immdec.imm11_7[3] ),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold442 (.A(_0942_),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold443 (.A(_0977_),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold444 (.A(_0127_),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold445 (.A(\rf_shift_reg.x[4][21] ),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold446 (.A(\rf_shift_reg.x[1][5] ),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold447 (.A(\dut.xfer.next_obuffer[7] ),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold448 (.A(\rf_shift_reg.x[3][28] ),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold449 (.A(\rf_shift_reg.x[2][28] ),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold450 (.A(\dut.dout_data[3] ),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold451 (.A(\dut.xfer.next_obuffer[2] ),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold452 (.A(_0417_),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold453 (.A(\cpu.bufreg2.dat[13] ),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold454 (.A(_0384_),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold455 (.A(\rf_shift_reg.x[1][15] ),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold456 (.A(\rf_shift_reg.x[2][7] ),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold457 (.A(\rf_shift_reg.x[3][5] ),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold458 (.A(_0169_),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold459 (.A(\rf_shift_reg.x[3][13] ),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold460 (.A(_0177_),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold461 (.A(\rf_shift_reg.x[4][28] ),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold462 (.A(\rf_shift_reg.x[2][21] ),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold463 (.A(\rf_shift_reg.x[4][19] ),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold464 (.A(\rf_shift_reg.x[2][14] ),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold465 (.A(\dut.buffer[22] ),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold466 (.A(_0501_),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold467 (.A(\dut.state[10] ),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold468 (.A(_0005_),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold469 (.A(\dut.buffer[21] ),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold470 (.A(_0500_),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold471 (.A(\cpu.bufreg.data[27] ),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold472 (.A(\cpu.ctrl.i_jump ),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold473 (.A(_0409_),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold474 (.A(\rf_shift_reg.x[3][12] ),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold475 (.A(\rf_shift_reg.x[1][26] ),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold476 (.A(\rf_shift_reg.x[4][11] ),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold477 (.A(\rf_shift_reg.x[2][25] ),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold478 (.A(\rf_shift_reg.x[4][17] ),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold479 (.A(\cpu.bufreg2.dat[30] ),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold480 (.A(_0401_),
    .X(net1111));
 sg13g2_dlygate4sd3_1 hold481 (.A(\rf_shift_reg.x[3][3] ),
    .X(net1112));
 sg13g2_dlygate4sd3_1 hold482 (.A(\rf_shift_reg.x[3][21] ),
    .X(net1113));
 sg13g2_dlygate4sd3_1 hold483 (.A(\dut.dout_data[2] ),
    .X(net1114));
 sg13g2_dlygate4sd3_1 hold484 (.A(\rf_shift_reg.x[3][15] ),
    .X(net1115));
 sg13g2_dlygate4sd3_1 hold485 (.A(\cpu.bufreg2.i_dat[19] ),
    .X(net1116));
 sg13g2_dlygate4sd3_1 hold486 (.A(\cpu.bufreg.data[9] ),
    .X(net1117));
 sg13g2_dlygate4sd3_1 hold487 (.A(_0314_),
    .X(net1118));
 sg13g2_dlygate4sd3_1 hold488 (.A(\dut.rd_addr[6] ),
    .X(net1119));
 sg13g2_dlygate4sd3_1 hold489 (.A(_0429_),
    .X(net1120));
 sg13g2_dlygate4sd3_1 hold490 (.A(\rf_shift_reg.x[1][12] ),
    .X(net1121));
 sg13g2_dlygate4sd3_1 hold491 (.A(\rf_shift_reg.x[3][4] ),
    .X(net1122));
 sg13g2_dlygate4sd3_1 hold492 (.A(\rf_shift_reg.x[1][21] ),
    .X(net1123));
 sg13g2_dlygate4sd3_1 hold493 (.A(\rf_shift_reg.x[1][28] ),
    .X(net1124));
 sg13g2_dlygate4sd3_1 hold494 (.A(\dut.dout_data[6] ),
    .X(net1125));
 sg13g2_dlygate4sd3_1 hold495 (.A(\cpu.bufreg.data[28] ),
    .X(net1126));
 sg13g2_dlygate4sd3_1 hold496 (.A(\rf_shift_reg.x[2][10] ),
    .X(net1127));
 sg13g2_dlygate4sd3_1 hold497 (.A(\dut.flash_csb ),
    .X(net1128));
 sg13g2_dlygate4sd3_1 hold498 (.A(\cpu.ctrl.pc_plus_4_cy_r ),
    .X(net1129));
 sg13g2_dlygate4sd3_1 hold499 (.A(_0902_),
    .X(net1130));
 sg13g2_dlygate4sd3_1 hold500 (.A(_0015_),
    .X(net1131));
 sg13g2_dlygate4sd3_1 hold501 (.A(\rf_shift_reg.x[5][10] ),
    .X(net1132));
 sg13g2_dlygate4sd3_1 hold502 (.A(\rf_shift_reg.x[4][3] ),
    .X(net1133));
 sg13g2_dlygate4sd3_1 hold503 (.A(\rf_shift_reg.x[5][16] ),
    .X(net1134));
 sg13g2_dlygate4sd3_1 hold504 (.A(\rf_shift_reg.x[5][28] ),
    .X(net1135));
 sg13g2_dlygate4sd3_1 hold505 (.A(\rf_shift_reg.x[3][24] ),
    .X(net1136));
 sg13g2_dlygate4sd3_1 hold506 (.A(\cpu.bufreg.data[8] ),
    .X(net1137));
 sg13g2_dlygate4sd3_1 hold507 (.A(\rf_shift_reg.cnt[4] ),
    .X(net1138));
 sg13g2_dlygate4sd3_1 hold508 (.A(_0132_),
    .X(net1139));
 sg13g2_dlygate4sd3_1 hold509 (.A(\rf_shift_reg.rreq_2r ),
    .X(net1140));
 sg13g2_dlygate4sd3_1 hold510 (.A(_0938_),
    .X(net1141));
 sg13g2_dlygate4sd3_1 hold511 (.A(\rf_shift_reg.x[5][14] ),
    .X(net1142));
 sg13g2_dlygate4sd3_1 hold512 (.A(\cpu.bufreg2.dat[26] ),
    .X(net1143));
 sg13g2_dlygate4sd3_1 hold513 (.A(_0397_),
    .X(net1144));
 sg13g2_dlygate4sd3_1 hold514 (.A(\rf_shift_reg.x[5][6] ),
    .X(net1145));
 sg13g2_dlygate4sd3_1 hold515 (.A(\rf_shift_reg.x[4][4] ),
    .X(net1146));
 sg13g2_dlygate4sd3_1 hold516 (.A(\rf_shift_reg.x[5][11] ),
    .X(net1147));
 sg13g2_dlygate4sd3_1 hold517 (.A(\cpu.bufreg.data[4] ),
    .X(net1148));
 sg13g2_dlygate4sd3_1 hold518 (.A(_0309_),
    .X(net1149));
 sg13g2_dlygate4sd3_1 hold519 (.A(\rf_shift_reg.x[3][25] ),
    .X(net1150));
 sg13g2_dlygate4sd3_1 hold520 (.A(\rf_shift_reg.x[1][8] ),
    .X(net1151));
 sg13g2_dlygate4sd3_1 hold521 (.A(\cpu.bufreg.data[5] ),
    .X(net1152));
 sg13g2_dlygate4sd3_1 hold522 (.A(\dut.buffer[19] ),
    .X(net1153));
 sg13g2_dlygate4sd3_1 hold523 (.A(\rf_shift_reg.x[4][29] ),
    .X(net1154));
 sg13g2_dlygate4sd3_1 hold524 (.A(\cpu.bufreg2.dat[19] ),
    .X(net1155));
 sg13g2_dlygate4sd3_1 hold525 (.A(\dut.softreset ),
    .X(net1156));
 sg13g2_dlygate4sd3_1 hold526 (.A(\rf_shift_reg.x[2][8] ),
    .X(net1157));
 sg13g2_dlygate4sd3_1 hold527 (.A(\cpu.bufreg.data[3] ),
    .X(net1158));
 sg13g2_dlygate4sd3_1 hold528 (.A(_0308_),
    .X(net1159));
 sg13g2_dlygate4sd3_1 hold529 (.A(\rf_shift_reg.x[2][22] ),
    .X(net1160));
 sg13g2_dlygate4sd3_1 hold530 (.A(\cpu.bufreg.data[20] ),
    .X(net1161));
 sg13g2_dlygate4sd3_1 hold531 (.A(\rf_shift_reg.x[3][30] ),
    .X(net1162));
 sg13g2_dlygate4sd3_1 hold532 (.A(\cpu.bufreg.data[23] ),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold533 (.A(_0328_),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold534 (.A(\rf_shift_reg.x[4][14] ),
    .X(net1165));
 sg13g2_dlygate4sd3_1 hold535 (.A(\rf_shift_reg.x[4][25] ),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold536 (.A(\dut.din_data[3] ),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold537 (.A(_0538_),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold538 (.A(\rf_shift_reg.x[2][2] ),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold539 (.A(\cpu.bufreg.data[22] ),
    .X(net1170));
 sg13g2_dlygate4sd3_1 hold540 (.A(\rf_shift_reg.x[5][29] ),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold541 (.A(\dut.din_data[1] ),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold542 (.A(_0540_),
    .X(net1173));
 sg13g2_dlygate4sd3_1 hold543 (.A(\cpu.immdec.imm19_12_20[3] ),
    .X(net1174));
 sg13g2_dlygate4sd3_1 hold544 (.A(_1097_),
    .X(net1175));
 sg13g2_dlygate4sd3_1 hold545 (.A(\cpu.bufreg2.dat[28] ),
    .X(net1176));
 sg13g2_dlygate4sd3_1 hold546 (.A(_0399_),
    .X(net1177));
 sg13g2_dlygate4sd3_1 hold547 (.A(\dut.state[5] ),
    .X(net1178));
 sg13g2_dlygate4sd3_1 hold548 (.A(_0003_),
    .X(net1179));
 sg13g2_dlygate4sd3_1 hold549 (.A(\rf_shift_reg.x[4][23] ),
    .X(net1180));
 sg13g2_dlygate4sd3_1 hold550 (.A(\rf_shift_reg.x[2][5] ),
    .X(net1181));
 sg13g2_dlygate4sd3_1 hold551 (.A(\cpu.bufreg.data[25] ),
    .X(net1182));
 sg13g2_dlygate4sd3_1 hold552 (.A(\cpu.alu.cmp_r ),
    .X(net1183));
 sg13g2_dlygate4sd3_1 hold553 (.A(\dut.state[4] ),
    .X(net1184));
 sg13g2_dlygate4sd3_1 hold554 (.A(\cpu.immdec.imm11_7[1] ),
    .X(net1185));
 sg13g2_dlygate4sd3_1 hold555 (.A(_0994_),
    .X(net1186));
 sg13g2_dlygate4sd3_1 hold556 (.A(_0196_),
    .X(net1187));
 sg13g2_dlygate4sd3_1 hold557 (.A(\dut.din_data[7] ),
    .X(net1188));
 sg13g2_dlygate4sd3_1 hold558 (.A(\cpu.bufreg.data[1] ),
    .X(net1189));
 sg13g2_dlygate4sd3_1 hold559 (.A(_0447_),
    .X(net1190));
 sg13g2_dlygate4sd3_1 hold560 (.A(\dut.state[9] ),
    .X(net1191));
 sg13g2_dlygate4sd3_1 hold561 (.A(_0009_),
    .X(net1192));
 sg13g2_dlygate4sd3_1 hold562 (.A(\dut.din_data[5] ),
    .X(net1193));
 sg13g2_dlygate4sd3_1 hold563 (.A(\rf_shift_reg.x[2][11] ),
    .X(net1194));
 sg13g2_dlygate4sd3_1 hold564 (.A(\dut.rd_addr[1] ),
    .X(net1195));
 sg13g2_dlygate4sd3_1 hold565 (.A(\cpu.bufreg2.dat[17] ),
    .X(net1196));
 sg13g2_dlygate4sd3_1 hold566 (.A(_0388_),
    .X(net1197));
 sg13g2_dlygate4sd3_1 hold567 (.A(\cpu.bufreg2.dat[7] ),
    .X(net1198));
 sg13g2_dlygate4sd3_1 hold568 (.A(_0378_),
    .X(net1199));
 sg13g2_dlygate4sd3_1 hold569 (.A(uo_out[2]),
    .X(net1200));
 sg13g2_dlygate4sd3_1 hold570 (.A(_0268_),
    .X(net1201));
 sg13g2_dlygate4sd3_1 hold571 (.A(\dut.din_data[4] ),
    .X(net1202));
 sg13g2_dlygate4sd3_1 hold572 (.A(\dut.din_data[0] ),
    .X(net1203));
 sg13g2_dlygate4sd3_1 hold573 (.A(_0541_),
    .X(net1204));
 sg13g2_dlygate4sd3_1 hold574 (.A(uo_out[0]),
    .X(net1205));
 sg13g2_dlygate4sd3_1 hold575 (.A(_0266_),
    .X(net1206));
 sg13g2_dlygate4sd3_1 hold576 (.A(\cpu.bufreg2.dat[8] ),
    .X(net1207));
 sg13g2_dlygate4sd3_1 hold577 (.A(_0379_),
    .X(net1208));
 sg13g2_dlygate4sd3_1 hold578 (.A(\cpu.decode.co_ebreak ),
    .X(net1209));
 sg13g2_dlygate4sd3_1 hold579 (.A(_0362_),
    .X(net1210));
 sg13g2_dlygate4sd3_1 hold580 (.A(\cpu.state.cnt_r[3] ),
    .X(net1211));
 sg13g2_dlygate4sd3_1 hold581 (.A(_0410_),
    .X(net1212));
 sg13g2_dlygate4sd3_1 hold582 (.A(uo_out[1]),
    .X(net1213));
 sg13g2_dlygate4sd3_1 hold583 (.A(_0267_),
    .X(net1214));
 sg13g2_dlygate4sd3_1 hold584 (.A(\dut.rd_wait ),
    .X(net1215));
 sg13g2_dlygate4sd3_1 hold585 (.A(_0467_),
    .X(net1216));
 sg13g2_dlygate4sd3_1 hold586 (.A(\cpu.immdec.imm24_20[1] ),
    .X(net1217));
 sg13g2_dlygate4sd3_1 hold587 (.A(_1134_),
    .X(net1218));
 sg13g2_dlygate4sd3_1 hold588 (.A(_0358_),
    .X(net1219));
 sg13g2_dlygate4sd3_1 hold589 (.A(\dut.din_rd ),
    .X(net1220));
 sg13g2_dlygate4sd3_1 hold590 (.A(_0452_),
    .X(net1221));
 sg13g2_dlygate4sd3_1 hold591 (.A(\cpu.state.init_done ),
    .X(net1222));
 sg13g2_dlygate4sd3_1 hold592 (.A(_0404_),
    .X(net1223));
 sg13g2_dlygate4sd3_1 hold593 (.A(\dut.rd_addr[14] ),
    .X(net1224));
 sg13g2_dlygate4sd3_1 hold594 (.A(_0437_),
    .X(net1225));
 sg13g2_dlygate4sd3_1 hold595 (.A(uo_out[4]),
    .X(net1226));
 sg13g2_dlygate4sd3_1 hold596 (.A(_0270_),
    .X(net1227));
 sg13g2_dlygate4sd3_1 hold597 (.A(\cpu.bufreg2.dat[11] ),
    .X(net1228));
 sg13g2_dlygate4sd3_1 hold598 (.A(\cpu.ctrl.pc_plus_offset_cy_r ),
    .X(net1229));
 sg13g2_dlygate4sd3_1 hold599 (.A(_0911_),
    .X(net1230));
 sg13g2_dlygate4sd3_1 hold600 (.A(_0016_),
    .X(net1231));
 sg13g2_dlygate4sd3_1 hold601 (.A(\dut.state[12] ),
    .X(net1232));
 sg13g2_dlygate4sd3_1 hold602 (.A(_0004_),
    .X(net1233));
 sg13g2_dlygate4sd3_1 hold603 (.A(\cpu.bufreg2.i_dat[7] ),
    .X(net1234));
 sg13g2_dlygate4sd3_1 hold604 (.A(_0350_),
    .X(net1235));
 sg13g2_dlygate4sd3_1 hold605 (.A(\cpu.bufreg2.i_dat[30] ),
    .X(net1236));
 sg13g2_dlygate4sd3_1 hold606 (.A(\dut.state[11] ),
    .X(net1237));
 sg13g2_dlygate4sd3_1 hold607 (.A(_0006_),
    .X(net1238));
 sg13g2_dlygate4sd3_1 hold608 (.A(\cpu.bufreg2.i_dat[13] ),
    .X(net1239));
 sg13g2_dlygate4sd3_1 hold609 (.A(_0343_),
    .X(net1240));
 sg13g2_dlygate4sd3_1 hold610 (.A(\dut.xfer.dummy_count[3] ),
    .X(net1241));
 sg13g2_dlygate4sd3_1 hold611 (.A(\cpu.bufreg2.dat[16] ),
    .X(net1242));
 sg13g2_dlygate4sd3_1 hold612 (.A(_0387_),
    .X(net1243));
 sg13g2_dlygate4sd3_1 hold613 (.A(uo_out[3]),
    .X(net1244));
 sg13g2_dlygate4sd3_1 hold614 (.A(_0269_),
    .X(net1245));
 sg13g2_dlygate4sd3_1 hold615 (.A(\dut.state[3] ),
    .X(net1246));
 sg13g2_dlygate4sd3_1 hold616 (.A(\dut.xfer.dummy_count[1] ),
    .X(net1247));
 sg13g2_dlygate4sd3_1 hold617 (.A(\cpu.bufreg.i_sh_signed ),
    .X(net1248));
 sg13g2_dlygate4sd3_1 hold618 (.A(\cpu.state.cnt_r[0] ),
    .X(net1249));
 sg13g2_dlygate4sd3_1 hold619 (.A(_0620_),
    .X(net1250));
 sg13g2_dlygate4sd3_1 hold620 (.A(\cpu.ctrl.o_ibus_adr[0] ),
    .X(net1251));
 sg13g2_dlygate4sd3_1 hold621 (.A(\cpu.immdec.imm30_25[0] ),
    .X(net1252));
 sg13g2_dlygate4sd3_1 hold622 (.A(_0351_),
    .X(net1253));
 sg13g2_dlygate4sd3_1 hold623 (.A(\cpu.immdec.imm19_12_20[5] ),
    .X(net1254));
 sg13g2_dlygate4sd3_1 hold624 (.A(_0345_),
    .X(net1255));
 sg13g2_dlygate4sd3_1 hold625 (.A(\cpu.bufreg2.i_dat[25] ),
    .X(net1256));
 sg13g2_dlygate4sd3_1 hold626 (.A(\cpu.bufreg2.i_dat[5] ),
    .X(net1257));
 sg13g2_dlygate4sd3_1 hold627 (.A(_0369_),
    .X(net1258));
 sg13g2_dlygate4sd3_1 hold628 (.A(\dut.rd_valid ),
    .X(net1259));
 sg13g2_dlygate4sd3_1 hold629 (.A(_0468_),
    .X(net1260));
 sg13g2_dlygate4sd3_1 hold630 (.A(\cpu.bufreg2.i_dat[29] ),
    .X(net1261));
 sg13g2_dlygate4sd3_1 hold631 (.A(\cpu.bufreg2.i_dat[31] ),
    .X(net1262));
 sg13g2_dlygate4sd3_1 hold632 (.A(\cpu.bufreg2.i_dat[27] ),
    .X(net1263));
 sg13g2_dlygate4sd3_1 hold633 (.A(\cpu.bufreg2.i_dat[28] ),
    .X(net1264));
 sg13g2_dlygate4sd3_1 hold634 (.A(\rf_shift_reg.x[2][31] ),
    .X(net1265));
 sg13g2_dlygate4sd3_1 hold635 (.A(_0164_),
    .X(net1266));
 sg13g2_dlygate4sd3_1 hold636 (.A(\dut.din_data[2] ),
    .X(net1267));
 sg13g2_dlygate4sd3_1 hold637 (.A(\cpu.bufreg2.i_dat[6] ),
    .X(net1268));
 sg13g2_dlygate4sd3_1 hold638 (.A(_0370_),
    .X(net1269));
 sg13g2_dlygate4sd3_1 hold639 (.A(\cpu.bufreg2.i_dat[26] ),
    .X(net1270));
 sg13g2_dlygate4sd3_1 hold640 (.A(\dut.state[2] ),
    .X(net1271));
 sg13g2_dlygate4sd3_1 hold641 (.A(\cpu.bufreg2.dat[24] ),
    .X(net1272));
 sg13g2_dlygate4sd3_1 hold642 (.A(_0395_),
    .X(net1273));
 sg13g2_dlygate4sd3_1 hold643 (.A(\dut.xfer.dummy_count[2] ),
    .X(net1274));
 sg13g2_dlygate4sd3_1 hold644 (.A(_1390_),
    .X(net1275));
 sg13g2_dlygate4sd3_1 hold645 (.A(\cpu.immdec.imm11_7[4] ),
    .X(net1276));
 sg13g2_dlygate4sd3_1 hold646 (.A(\cpu.bufreg2.i_dat[24] ),
    .X(net1277));
 sg13g2_dlygate4sd3_1 hold647 (.A(\dut.state[1] ),
    .X(net1278));
 sg13g2_dlygate4sd3_1 hold648 (.A(\cpu.bufreg2.dat[5] ),
    .X(net1279));
 sg13g2_dlygate4sd3_1 hold649 (.A(\cpu.immdec.imm19_12_20[1] ),
    .X(net1280));
 sg13g2_dlygate4sd3_1 hold650 (.A(_1088_),
    .X(net1281));
 sg13g2_dlygate4sd3_1 hold651 (.A(_0341_),
    .X(net1282));
 sg13g2_dlygate4sd3_1 hold652 (.A(\cpu.bufreg.data[31] ),
    .X(net1283));
 sg13g2_dlygate4sd3_1 hold653 (.A(_0337_),
    .X(net1284));
 sg13g2_dlygate4sd3_1 hold654 (.A(\cpu.bufreg2.i_dat[20] ),
    .X(net1285));
 sg13g2_dlygate4sd3_1 hold655 (.A(\cpu.bufreg2.i_dat[12] ),
    .X(net1286));
 sg13g2_dlygate4sd3_1 hold656 (.A(_0342_),
    .X(net1287));
 sg13g2_dlygate4sd3_1 hold657 (.A(\cpu.immdec.imm11_7[2] ),
    .X(net1288));
 sg13g2_dlygate4sd3_1 hold658 (.A(\cpu.bufreg.data[2] ),
    .X(net1289));
 sg13g2_dlygate4sd3_1 hold659 (.A(_1376_),
    .X(net1290));
 sg13g2_dlygate4sd3_1 hold660 (.A(_0448_),
    .X(net1291));
 sg13g2_dlygate4sd3_1 hold661 (.A(\cpu.mem_bytecnt[0] ),
    .X(net1292));
 sg13g2_dlygate4sd3_1 hold662 (.A(_1262_),
    .X(net1293));
 sg13g2_dlygate4sd3_1 hold663 (.A(_0411_),
    .X(net1294));
 sg13g2_dlygate4sd3_1 hold664 (.A(\cpu.bufreg2.i_dat[4] ),
    .X(net1295));
 sg13g2_dlygate4sd3_1 hold665 (.A(_0368_),
    .X(net1296));
 sg13g2_dlygate4sd3_1 hold666 (.A(\cpu.bufreg2.i_dat[17] ),
    .X(net1297));
 sg13g2_dlygate4sd3_1 hold667 (.A(_1105_),
    .X(net1298));
 sg13g2_dlygate4sd3_1 hold668 (.A(\dut.state[1] ),
    .X(net1299));
 sg13g2_dlygate4sd3_1 hold669 (.A(\cpu.bufreg2.dat[3] ),
    .X(net1300));
 sg13g2_dlygate4sd3_1 hold670 (.A(_0374_),
    .X(net1301));
 sg13g2_dlygate4sd3_1 hold671 (.A(\cpu.bufreg2.i_dat[3] ),
    .X(net1302));
 sg13g2_dlygate4sd3_1 hold672 (.A(_0367_),
    .X(net1303));
 sg13g2_dlygate4sd3_1 hold673 (.A(\cpu.bne_or_bge ),
    .X(net1304));
 sg13g2_dlygate4sd3_1 hold674 (.A(\cpu.bufreg2.i_dat[16] ),
    .X(net1305));
 sg13g2_dlygate4sd3_1 hold675 (.A(_1103_),
    .X(net1306));
 sg13g2_dlygate4sd3_1 hold676 (.A(\cpu.immdec.imm11_7[0] ),
    .X(net1307));
 sg13g2_dlygate4sd3_1 hold677 (.A(\rf_shift_reg.cnt[2] ),
    .X(net1308));
 sg13g2_dlygate4sd3_1 hold678 (.A(_0984_),
    .X(net1309));
 sg13g2_dlygate4sd3_1 hold679 (.A(_0130_),
    .X(net1310));
 sg13g2_dlygate4sd3_1 hold680 (.A(_0086_),
    .X(net1311));
 sg13g2_dlygate4sd3_1 hold681 (.A(_0824_),
    .X(net1312));
 sg13g2_dlygate4sd3_1 hold682 (.A(\cpu.bufreg2.i_dat[2] ),
    .X(net1313));
 sg13g2_dlygate4sd3_1 hold683 (.A(_0366_),
    .X(net1314));
 sg13g2_dlygate4sd3_1 hold684 (.A(\dut.rd_addr[2] ),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold685 (.A(_0425_),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold686 (.A(\cpu.bufreg2.dat[2] ),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold687 (.A(\cpu.bufreg2.dat[4] ),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold688 (.A(\cpu.csr_d_sel ),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold689 (.A(_0089_),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold690 (.A(\rf_shift_reg.cnt[3] ),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold691 (.A(_0986_),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold692 (.A(\cpu.bufreg2.dat[0] ),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold693 (.A(_0371_),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold694 (.A(\cpu.bufreg2.dat[1] ),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold695 (.A(_0372_),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold696 (.A(\cpu.mem_bytecnt[1] ),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold697 (.A(_0412_),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold698 (.A(\dut.xfer.count[3] ),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold699 (.A(_1379_),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold700 (.A(_0451_),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold701 (.A(\cpu.bufreg2.i_dat[22] ),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold702 (.A(_1136_),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold703 (.A(\cpu.bufreg2.i_dat[8] ),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold704 (.A(\cpu.bufreg2.i_op_b_sel ),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold705 (.A(_0857_),
    .X(net1336));
 sg13g2_dlygate4sd3_1 hold706 (.A(_0013_),
    .X(net1337));
 sg13g2_dlygate4sd3_1 hold707 (.A(\cpu.decode.co_mem_word ),
    .X(net1338));
 sg13g2_dlygate4sd3_1 hold708 (.A(\dut.rd_addr[3] ),
    .X(net1339));
 sg13g2_dlygate4sd3_1 hold709 (.A(_0426_),
    .X(net1340));
 sg13g2_dlygate4sd3_1 hold710 (.A(\cpu.state.ibus_cyc ),
    .X(net1341));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_decap_8 FILLER_13_588 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_decap_8 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_637 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_8 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_decap_8 FILLER_13_798 ();
 sg13g2_decap_8 FILLER_13_805 ();
 sg13g2_decap_8 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_833 ();
 sg13g2_decap_8 FILLER_13_840 ();
 sg13g2_decap_8 FILLER_13_847 ();
 sg13g2_decap_8 FILLER_13_854 ();
 sg13g2_fill_1 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_8 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_511 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_574 ();
 sg13g2_decap_8 FILLER_14_581 ();
 sg13g2_decap_8 FILLER_14_588 ();
 sg13g2_decap_8 FILLER_14_595 ();
 sg13g2_decap_8 FILLER_14_602 ();
 sg13g2_decap_8 FILLER_14_609 ();
 sg13g2_decap_8 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_623 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_decap_8 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_decap_8 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_658 ();
 sg13g2_decap_8 FILLER_14_665 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_decap_8 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_decap_8 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_14_840 ();
 sg13g2_decap_8 FILLER_14_847 ();
 sg13g2_decap_8 FILLER_14_854 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_434 ();
 sg13g2_decap_8 FILLER_15_441 ();
 sg13g2_decap_8 FILLER_15_448 ();
 sg13g2_decap_8 FILLER_15_455 ();
 sg13g2_decap_8 FILLER_15_462 ();
 sg13g2_decap_8 FILLER_15_469 ();
 sg13g2_decap_8 FILLER_15_476 ();
 sg13g2_decap_8 FILLER_15_483 ();
 sg13g2_decap_8 FILLER_15_490 ();
 sg13g2_decap_8 FILLER_15_497 ();
 sg13g2_decap_8 FILLER_15_504 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_518 ();
 sg13g2_decap_8 FILLER_15_525 ();
 sg13g2_decap_8 FILLER_15_532 ();
 sg13g2_decap_8 FILLER_15_539 ();
 sg13g2_decap_8 FILLER_15_546 ();
 sg13g2_decap_8 FILLER_15_553 ();
 sg13g2_decap_8 FILLER_15_560 ();
 sg13g2_decap_8 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_574 ();
 sg13g2_decap_8 FILLER_15_581 ();
 sg13g2_decap_8 FILLER_15_588 ();
 sg13g2_decap_8 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_602 ();
 sg13g2_decap_8 FILLER_15_609 ();
 sg13g2_decap_8 FILLER_15_616 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_8 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_644 ();
 sg13g2_decap_8 FILLER_15_651 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_decap_8 FILLER_15_665 ();
 sg13g2_decap_8 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_679 ();
 sg13g2_decap_8 FILLER_15_686 ();
 sg13g2_decap_8 FILLER_15_693 ();
 sg13g2_decap_8 FILLER_15_700 ();
 sg13g2_decap_8 FILLER_15_707 ();
 sg13g2_decap_8 FILLER_15_714 ();
 sg13g2_decap_8 FILLER_15_721 ();
 sg13g2_decap_8 FILLER_15_728 ();
 sg13g2_decap_8 FILLER_15_735 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_decap_8 FILLER_15_749 ();
 sg13g2_decap_8 FILLER_15_756 ();
 sg13g2_decap_8 FILLER_15_763 ();
 sg13g2_decap_8 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_777 ();
 sg13g2_decap_8 FILLER_15_784 ();
 sg13g2_decap_8 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_798 ();
 sg13g2_decap_8 FILLER_15_805 ();
 sg13g2_decap_8 FILLER_15_812 ();
 sg13g2_decap_8 FILLER_15_819 ();
 sg13g2_decap_8 FILLER_15_826 ();
 sg13g2_decap_8 FILLER_15_833 ();
 sg13g2_decap_8 FILLER_15_840 ();
 sg13g2_decap_8 FILLER_15_847 ();
 sg13g2_decap_8 FILLER_15_854 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_8 FILLER_16_455 ();
 sg13g2_decap_8 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_469 ();
 sg13g2_decap_8 FILLER_16_476 ();
 sg13g2_decap_8 FILLER_16_483 ();
 sg13g2_decap_8 FILLER_16_490 ();
 sg13g2_decap_8 FILLER_16_497 ();
 sg13g2_decap_8 FILLER_16_504 ();
 sg13g2_decap_8 FILLER_16_511 ();
 sg13g2_decap_8 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_525 ();
 sg13g2_decap_8 FILLER_16_532 ();
 sg13g2_decap_8 FILLER_16_539 ();
 sg13g2_decap_8 FILLER_16_546 ();
 sg13g2_decap_8 FILLER_16_553 ();
 sg13g2_decap_8 FILLER_16_560 ();
 sg13g2_decap_8 FILLER_16_567 ();
 sg13g2_decap_8 FILLER_16_574 ();
 sg13g2_decap_8 FILLER_16_581 ();
 sg13g2_decap_8 FILLER_16_588 ();
 sg13g2_decap_8 FILLER_16_595 ();
 sg13g2_decap_8 FILLER_16_602 ();
 sg13g2_decap_8 FILLER_16_609 ();
 sg13g2_decap_8 FILLER_16_616 ();
 sg13g2_decap_8 FILLER_16_623 ();
 sg13g2_decap_8 FILLER_16_630 ();
 sg13g2_decap_8 FILLER_16_637 ();
 sg13g2_decap_8 FILLER_16_644 ();
 sg13g2_decap_8 FILLER_16_651 ();
 sg13g2_decap_8 FILLER_16_658 ();
 sg13g2_decap_8 FILLER_16_665 ();
 sg13g2_decap_8 FILLER_16_672 ();
 sg13g2_decap_8 FILLER_16_679 ();
 sg13g2_decap_8 FILLER_16_686 ();
 sg13g2_decap_8 FILLER_16_693 ();
 sg13g2_decap_8 FILLER_16_700 ();
 sg13g2_decap_8 FILLER_16_707 ();
 sg13g2_decap_8 FILLER_16_714 ();
 sg13g2_decap_8 FILLER_16_721 ();
 sg13g2_decap_8 FILLER_16_728 ();
 sg13g2_decap_8 FILLER_16_735 ();
 sg13g2_decap_8 FILLER_16_742 ();
 sg13g2_decap_8 FILLER_16_749 ();
 sg13g2_decap_8 FILLER_16_756 ();
 sg13g2_decap_8 FILLER_16_763 ();
 sg13g2_decap_8 FILLER_16_770 ();
 sg13g2_decap_8 FILLER_16_777 ();
 sg13g2_decap_8 FILLER_16_784 ();
 sg13g2_decap_8 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_798 ();
 sg13g2_decap_8 FILLER_16_805 ();
 sg13g2_decap_8 FILLER_16_812 ();
 sg13g2_decap_8 FILLER_16_819 ();
 sg13g2_decap_8 FILLER_16_826 ();
 sg13g2_decap_8 FILLER_16_833 ();
 sg13g2_decap_8 FILLER_16_840 ();
 sg13g2_decap_8 FILLER_16_847 ();
 sg13g2_decap_8 FILLER_16_854 ();
 sg13g2_fill_1 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_427 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_448 ();
 sg13g2_decap_8 FILLER_17_455 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_497 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_fill_1 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_decap_8 FILLER_18_427 ();
 sg13g2_decap_8 FILLER_18_434 ();
 sg13g2_decap_8 FILLER_18_441 ();
 sg13g2_decap_8 FILLER_18_448 ();
 sg13g2_decap_8 FILLER_18_455 ();
 sg13g2_decap_8 FILLER_18_462 ();
 sg13g2_decap_8 FILLER_18_469 ();
 sg13g2_decap_8 FILLER_18_476 ();
 sg13g2_decap_8 FILLER_18_483 ();
 sg13g2_decap_8 FILLER_18_490 ();
 sg13g2_decap_8 FILLER_18_497 ();
 sg13g2_decap_8 FILLER_18_504 ();
 sg13g2_decap_8 FILLER_18_511 ();
 sg13g2_decap_8 FILLER_18_518 ();
 sg13g2_decap_8 FILLER_18_525 ();
 sg13g2_decap_8 FILLER_18_532 ();
 sg13g2_decap_8 FILLER_18_539 ();
 sg13g2_decap_8 FILLER_18_546 ();
 sg13g2_decap_8 FILLER_18_553 ();
 sg13g2_decap_8 FILLER_18_560 ();
 sg13g2_decap_8 FILLER_18_567 ();
 sg13g2_decap_8 FILLER_18_574 ();
 sg13g2_decap_8 FILLER_18_581 ();
 sg13g2_decap_8 FILLER_18_588 ();
 sg13g2_decap_8 FILLER_18_595 ();
 sg13g2_decap_8 FILLER_18_602 ();
 sg13g2_decap_8 FILLER_18_609 ();
 sg13g2_decap_8 FILLER_18_616 ();
 sg13g2_decap_8 FILLER_18_623 ();
 sg13g2_decap_8 FILLER_18_630 ();
 sg13g2_decap_8 FILLER_18_637 ();
 sg13g2_decap_8 FILLER_18_644 ();
 sg13g2_decap_8 FILLER_18_651 ();
 sg13g2_decap_8 FILLER_18_658 ();
 sg13g2_decap_8 FILLER_18_665 ();
 sg13g2_decap_8 FILLER_18_672 ();
 sg13g2_decap_8 FILLER_18_679 ();
 sg13g2_decap_8 FILLER_18_686 ();
 sg13g2_decap_8 FILLER_18_693 ();
 sg13g2_decap_8 FILLER_18_700 ();
 sg13g2_decap_8 FILLER_18_707 ();
 sg13g2_decap_8 FILLER_18_714 ();
 sg13g2_decap_8 FILLER_18_721 ();
 sg13g2_decap_8 FILLER_18_728 ();
 sg13g2_decap_8 FILLER_18_735 ();
 sg13g2_decap_8 FILLER_18_742 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_decap_8 FILLER_18_756 ();
 sg13g2_decap_8 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_770 ();
 sg13g2_decap_8 FILLER_18_777 ();
 sg13g2_decap_8 FILLER_18_784 ();
 sg13g2_decap_8 FILLER_18_791 ();
 sg13g2_decap_8 FILLER_18_798 ();
 sg13g2_decap_8 FILLER_18_805 ();
 sg13g2_decap_8 FILLER_18_812 ();
 sg13g2_decap_8 FILLER_18_819 ();
 sg13g2_decap_8 FILLER_18_826 ();
 sg13g2_decap_8 FILLER_18_833 ();
 sg13g2_decap_8 FILLER_18_840 ();
 sg13g2_decap_8 FILLER_18_847 ();
 sg13g2_decap_8 FILLER_18_854 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_decap_8 FILLER_19_427 ();
 sg13g2_decap_8 FILLER_19_434 ();
 sg13g2_decap_8 FILLER_19_441 ();
 sg13g2_decap_8 FILLER_19_448 ();
 sg13g2_decap_8 FILLER_19_455 ();
 sg13g2_decap_8 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_490 ();
 sg13g2_decap_8 FILLER_19_497 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_532 ();
 sg13g2_decap_8 FILLER_19_539 ();
 sg13g2_decap_8 FILLER_19_546 ();
 sg13g2_decap_8 FILLER_19_553 ();
 sg13g2_decap_8 FILLER_19_560 ();
 sg13g2_decap_8 FILLER_19_567 ();
 sg13g2_decap_8 FILLER_19_574 ();
 sg13g2_decap_8 FILLER_19_581 ();
 sg13g2_decap_8 FILLER_19_588 ();
 sg13g2_decap_8 FILLER_19_595 ();
 sg13g2_decap_8 FILLER_19_602 ();
 sg13g2_decap_8 FILLER_19_609 ();
 sg13g2_decap_8 FILLER_19_616 ();
 sg13g2_decap_8 FILLER_19_623 ();
 sg13g2_decap_8 FILLER_19_630 ();
 sg13g2_decap_8 FILLER_19_637 ();
 sg13g2_decap_8 FILLER_19_644 ();
 sg13g2_decap_8 FILLER_19_651 ();
 sg13g2_decap_8 FILLER_19_658 ();
 sg13g2_decap_8 FILLER_19_665 ();
 sg13g2_decap_8 FILLER_19_672 ();
 sg13g2_decap_8 FILLER_19_679 ();
 sg13g2_decap_8 FILLER_19_686 ();
 sg13g2_decap_8 FILLER_19_693 ();
 sg13g2_decap_8 FILLER_19_700 ();
 sg13g2_decap_8 FILLER_19_707 ();
 sg13g2_decap_8 FILLER_19_714 ();
 sg13g2_decap_8 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_784 ();
 sg13g2_decap_8 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_798 ();
 sg13g2_decap_8 FILLER_19_805 ();
 sg13g2_decap_8 FILLER_19_812 ();
 sg13g2_decap_8 FILLER_19_819 ();
 sg13g2_decap_8 FILLER_19_826 ();
 sg13g2_decap_8 FILLER_19_833 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_decap_8 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_854 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_decap_8 FILLER_20_427 ();
 sg13g2_decap_8 FILLER_20_434 ();
 sg13g2_decap_8 FILLER_20_441 ();
 sg13g2_decap_8 FILLER_20_448 ();
 sg13g2_decap_8 FILLER_20_455 ();
 sg13g2_decap_8 FILLER_20_462 ();
 sg13g2_decap_8 FILLER_20_469 ();
 sg13g2_decap_8 FILLER_20_476 ();
 sg13g2_decap_8 FILLER_20_483 ();
 sg13g2_decap_8 FILLER_20_490 ();
 sg13g2_decap_8 FILLER_20_497 ();
 sg13g2_decap_8 FILLER_20_504 ();
 sg13g2_decap_8 FILLER_20_511 ();
 sg13g2_decap_8 FILLER_20_518 ();
 sg13g2_decap_8 FILLER_20_525 ();
 sg13g2_decap_8 FILLER_20_532 ();
 sg13g2_decap_8 FILLER_20_539 ();
 sg13g2_decap_8 FILLER_20_546 ();
 sg13g2_decap_8 FILLER_20_553 ();
 sg13g2_decap_8 FILLER_20_560 ();
 sg13g2_decap_8 FILLER_20_567 ();
 sg13g2_decap_8 FILLER_20_574 ();
 sg13g2_decap_8 FILLER_20_581 ();
 sg13g2_decap_8 FILLER_20_588 ();
 sg13g2_decap_8 FILLER_20_595 ();
 sg13g2_decap_8 FILLER_20_602 ();
 sg13g2_decap_8 FILLER_20_609 ();
 sg13g2_decap_8 FILLER_20_616 ();
 sg13g2_decap_8 FILLER_20_623 ();
 sg13g2_decap_8 FILLER_20_630 ();
 sg13g2_decap_8 FILLER_20_637 ();
 sg13g2_decap_8 FILLER_20_644 ();
 sg13g2_decap_8 FILLER_20_651 ();
 sg13g2_decap_8 FILLER_20_658 ();
 sg13g2_decap_8 FILLER_20_665 ();
 sg13g2_decap_8 FILLER_20_672 ();
 sg13g2_decap_8 FILLER_20_679 ();
 sg13g2_decap_8 FILLER_20_686 ();
 sg13g2_decap_8 FILLER_20_693 ();
 sg13g2_decap_8 FILLER_20_700 ();
 sg13g2_decap_8 FILLER_20_707 ();
 sg13g2_decap_8 FILLER_20_714 ();
 sg13g2_decap_8 FILLER_20_721 ();
 sg13g2_decap_8 FILLER_20_728 ();
 sg13g2_decap_8 FILLER_20_735 ();
 sg13g2_decap_8 FILLER_20_742 ();
 sg13g2_decap_8 FILLER_20_749 ();
 sg13g2_decap_8 FILLER_20_756 ();
 sg13g2_decap_8 FILLER_20_763 ();
 sg13g2_decap_8 FILLER_20_770 ();
 sg13g2_decap_8 FILLER_20_777 ();
 sg13g2_decap_8 FILLER_20_784 ();
 sg13g2_decap_8 FILLER_20_791 ();
 sg13g2_decap_8 FILLER_20_798 ();
 sg13g2_decap_8 FILLER_20_805 ();
 sg13g2_decap_8 FILLER_20_812 ();
 sg13g2_decap_8 FILLER_20_819 ();
 sg13g2_decap_8 FILLER_20_826 ();
 sg13g2_decap_8 FILLER_20_833 ();
 sg13g2_decap_8 FILLER_20_840 ();
 sg13g2_decap_8 FILLER_20_847 ();
 sg13g2_decap_8 FILLER_20_854 ();
 sg13g2_fill_1 FILLER_20_861 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_decap_8 FILLER_21_427 ();
 sg13g2_decap_8 FILLER_21_434 ();
 sg13g2_decap_8 FILLER_21_441 ();
 sg13g2_decap_8 FILLER_21_448 ();
 sg13g2_decap_8 FILLER_21_455 ();
 sg13g2_decap_8 FILLER_21_462 ();
 sg13g2_decap_8 FILLER_21_469 ();
 sg13g2_decap_8 FILLER_21_476 ();
 sg13g2_decap_8 FILLER_21_483 ();
 sg13g2_decap_8 FILLER_21_490 ();
 sg13g2_decap_8 FILLER_21_497 ();
 sg13g2_decap_8 FILLER_21_504 ();
 sg13g2_decap_8 FILLER_21_511 ();
 sg13g2_decap_8 FILLER_21_518 ();
 sg13g2_decap_8 FILLER_21_525 ();
 sg13g2_decap_8 FILLER_21_532 ();
 sg13g2_decap_8 FILLER_21_539 ();
 sg13g2_decap_8 FILLER_21_546 ();
 sg13g2_decap_8 FILLER_21_553 ();
 sg13g2_decap_8 FILLER_21_560 ();
 sg13g2_decap_8 FILLER_21_567 ();
 sg13g2_decap_8 FILLER_21_574 ();
 sg13g2_decap_8 FILLER_21_581 ();
 sg13g2_decap_8 FILLER_21_588 ();
 sg13g2_decap_8 FILLER_21_595 ();
 sg13g2_decap_8 FILLER_21_602 ();
 sg13g2_decap_8 FILLER_21_609 ();
 sg13g2_decap_8 FILLER_21_616 ();
 sg13g2_decap_8 FILLER_21_623 ();
 sg13g2_decap_8 FILLER_21_630 ();
 sg13g2_decap_8 FILLER_21_637 ();
 sg13g2_decap_8 FILLER_21_644 ();
 sg13g2_decap_8 FILLER_21_651 ();
 sg13g2_decap_8 FILLER_21_658 ();
 sg13g2_decap_8 FILLER_21_665 ();
 sg13g2_decap_8 FILLER_21_672 ();
 sg13g2_decap_8 FILLER_21_679 ();
 sg13g2_decap_8 FILLER_21_686 ();
 sg13g2_decap_8 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_700 ();
 sg13g2_decap_8 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_714 ();
 sg13g2_decap_8 FILLER_21_721 ();
 sg13g2_decap_8 FILLER_21_728 ();
 sg13g2_decap_8 FILLER_21_735 ();
 sg13g2_decap_8 FILLER_21_742 ();
 sg13g2_decap_8 FILLER_21_749 ();
 sg13g2_decap_8 FILLER_21_756 ();
 sg13g2_decap_8 FILLER_21_763 ();
 sg13g2_decap_8 FILLER_21_770 ();
 sg13g2_decap_8 FILLER_21_777 ();
 sg13g2_decap_8 FILLER_21_784 ();
 sg13g2_decap_8 FILLER_21_791 ();
 sg13g2_decap_8 FILLER_21_798 ();
 sg13g2_decap_8 FILLER_21_805 ();
 sg13g2_decap_8 FILLER_21_812 ();
 sg13g2_decap_8 FILLER_21_819 ();
 sg13g2_decap_8 FILLER_21_826 ();
 sg13g2_decap_8 FILLER_21_833 ();
 sg13g2_decap_8 FILLER_21_840 ();
 sg13g2_decap_8 FILLER_21_847 ();
 sg13g2_decap_8 FILLER_21_854 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_22_406 ();
 sg13g2_decap_8 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_decap_8 FILLER_22_427 ();
 sg13g2_decap_8 FILLER_22_434 ();
 sg13g2_decap_8 FILLER_22_441 ();
 sg13g2_decap_8 FILLER_22_448 ();
 sg13g2_decap_8 FILLER_22_455 ();
 sg13g2_decap_8 FILLER_22_462 ();
 sg13g2_decap_8 FILLER_22_469 ();
 sg13g2_decap_8 FILLER_22_476 ();
 sg13g2_decap_8 FILLER_22_483 ();
 sg13g2_decap_8 FILLER_22_490 ();
 sg13g2_decap_8 FILLER_22_497 ();
 sg13g2_decap_8 FILLER_22_504 ();
 sg13g2_decap_8 FILLER_22_511 ();
 sg13g2_decap_8 FILLER_22_518 ();
 sg13g2_decap_8 FILLER_22_525 ();
 sg13g2_decap_8 FILLER_22_532 ();
 sg13g2_decap_8 FILLER_22_539 ();
 sg13g2_decap_8 FILLER_22_546 ();
 sg13g2_decap_8 FILLER_22_553 ();
 sg13g2_decap_8 FILLER_22_560 ();
 sg13g2_decap_8 FILLER_22_567 ();
 sg13g2_decap_8 FILLER_22_574 ();
 sg13g2_decap_8 FILLER_22_581 ();
 sg13g2_decap_8 FILLER_22_588 ();
 sg13g2_decap_8 FILLER_22_595 ();
 sg13g2_decap_8 FILLER_22_602 ();
 sg13g2_decap_8 FILLER_22_609 ();
 sg13g2_decap_8 FILLER_22_616 ();
 sg13g2_decap_8 FILLER_22_623 ();
 sg13g2_decap_8 FILLER_22_630 ();
 sg13g2_decap_8 FILLER_22_637 ();
 sg13g2_decap_8 FILLER_22_644 ();
 sg13g2_decap_8 FILLER_22_651 ();
 sg13g2_decap_8 FILLER_22_658 ();
 sg13g2_decap_8 FILLER_22_665 ();
 sg13g2_decap_8 FILLER_22_672 ();
 sg13g2_decap_8 FILLER_22_679 ();
 sg13g2_decap_8 FILLER_22_686 ();
 sg13g2_decap_8 FILLER_22_693 ();
 sg13g2_decap_8 FILLER_22_700 ();
 sg13g2_decap_8 FILLER_22_707 ();
 sg13g2_decap_8 FILLER_22_714 ();
 sg13g2_decap_8 FILLER_22_721 ();
 sg13g2_decap_8 FILLER_22_728 ();
 sg13g2_decap_8 FILLER_22_735 ();
 sg13g2_decap_8 FILLER_22_742 ();
 sg13g2_decap_8 FILLER_22_749 ();
 sg13g2_decap_8 FILLER_22_756 ();
 sg13g2_decap_8 FILLER_22_763 ();
 sg13g2_decap_8 FILLER_22_770 ();
 sg13g2_decap_8 FILLER_22_777 ();
 sg13g2_decap_8 FILLER_22_784 ();
 sg13g2_decap_8 FILLER_22_791 ();
 sg13g2_decap_8 FILLER_22_798 ();
 sg13g2_decap_8 FILLER_22_805 ();
 sg13g2_decap_8 FILLER_22_812 ();
 sg13g2_decap_8 FILLER_22_819 ();
 sg13g2_decap_8 FILLER_22_826 ();
 sg13g2_decap_8 FILLER_22_833 ();
 sg13g2_decap_8 FILLER_22_840 ();
 sg13g2_decap_8 FILLER_22_847 ();
 sg13g2_decap_8 FILLER_22_854 ();
 sg13g2_fill_1 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_decap_8 FILLER_23_406 ();
 sg13g2_decap_8 FILLER_23_413 ();
 sg13g2_decap_8 FILLER_23_420 ();
 sg13g2_decap_8 FILLER_23_427 ();
 sg13g2_decap_8 FILLER_23_434 ();
 sg13g2_decap_8 FILLER_23_441 ();
 sg13g2_decap_8 FILLER_23_448 ();
 sg13g2_decap_8 FILLER_23_455 ();
 sg13g2_decap_8 FILLER_23_462 ();
 sg13g2_decap_8 FILLER_23_469 ();
 sg13g2_decap_8 FILLER_23_476 ();
 sg13g2_decap_8 FILLER_23_483 ();
 sg13g2_decap_8 FILLER_23_490 ();
 sg13g2_decap_8 FILLER_23_497 ();
 sg13g2_decap_8 FILLER_23_504 ();
 sg13g2_decap_8 FILLER_23_511 ();
 sg13g2_decap_8 FILLER_23_518 ();
 sg13g2_decap_8 FILLER_23_525 ();
 sg13g2_decap_8 FILLER_23_532 ();
 sg13g2_decap_8 FILLER_23_539 ();
 sg13g2_decap_8 FILLER_23_546 ();
 sg13g2_decap_8 FILLER_23_553 ();
 sg13g2_decap_8 FILLER_23_560 ();
 sg13g2_decap_8 FILLER_23_567 ();
 sg13g2_decap_8 FILLER_23_574 ();
 sg13g2_decap_8 FILLER_23_581 ();
 sg13g2_decap_8 FILLER_23_588 ();
 sg13g2_decap_8 FILLER_23_595 ();
 sg13g2_decap_8 FILLER_23_602 ();
 sg13g2_decap_8 FILLER_23_609 ();
 sg13g2_decap_8 FILLER_23_616 ();
 sg13g2_decap_8 FILLER_23_623 ();
 sg13g2_decap_8 FILLER_23_630 ();
 sg13g2_decap_8 FILLER_23_637 ();
 sg13g2_decap_8 FILLER_23_644 ();
 sg13g2_decap_8 FILLER_23_651 ();
 sg13g2_decap_8 FILLER_23_658 ();
 sg13g2_decap_8 FILLER_23_665 ();
 sg13g2_decap_8 FILLER_23_672 ();
 sg13g2_decap_8 FILLER_23_679 ();
 sg13g2_decap_8 FILLER_23_686 ();
 sg13g2_decap_8 FILLER_23_693 ();
 sg13g2_decap_8 FILLER_23_700 ();
 sg13g2_decap_8 FILLER_23_707 ();
 sg13g2_decap_8 FILLER_23_714 ();
 sg13g2_decap_8 FILLER_23_721 ();
 sg13g2_decap_8 FILLER_23_728 ();
 sg13g2_decap_8 FILLER_23_735 ();
 sg13g2_decap_8 FILLER_23_742 ();
 sg13g2_decap_8 FILLER_23_749 ();
 sg13g2_decap_8 FILLER_23_756 ();
 sg13g2_decap_8 FILLER_23_763 ();
 sg13g2_decap_8 FILLER_23_770 ();
 sg13g2_decap_8 FILLER_23_777 ();
 sg13g2_decap_8 FILLER_23_784 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_798 ();
 sg13g2_decap_8 FILLER_23_805 ();
 sg13g2_decap_8 FILLER_23_812 ();
 sg13g2_decap_8 FILLER_23_819 ();
 sg13g2_decap_8 FILLER_23_826 ();
 sg13g2_decap_8 FILLER_23_833 ();
 sg13g2_decap_8 FILLER_23_840 ();
 sg13g2_decap_8 FILLER_23_847 ();
 sg13g2_decap_8 FILLER_23_854 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_decap_8 FILLER_24_406 ();
 sg13g2_decap_8 FILLER_24_413 ();
 sg13g2_decap_8 FILLER_24_420 ();
 sg13g2_decap_8 FILLER_24_427 ();
 sg13g2_decap_8 FILLER_24_434 ();
 sg13g2_decap_8 FILLER_24_441 ();
 sg13g2_decap_8 FILLER_24_448 ();
 sg13g2_decap_8 FILLER_24_455 ();
 sg13g2_decap_8 FILLER_24_462 ();
 sg13g2_decap_8 FILLER_24_469 ();
 sg13g2_decap_8 FILLER_24_476 ();
 sg13g2_decap_8 FILLER_24_483 ();
 sg13g2_decap_8 FILLER_24_490 ();
 sg13g2_decap_8 FILLER_24_497 ();
 sg13g2_decap_8 FILLER_24_504 ();
 sg13g2_decap_8 FILLER_24_511 ();
 sg13g2_decap_8 FILLER_24_518 ();
 sg13g2_decap_8 FILLER_24_525 ();
 sg13g2_decap_8 FILLER_24_532 ();
 sg13g2_decap_8 FILLER_24_539 ();
 sg13g2_decap_8 FILLER_24_546 ();
 sg13g2_decap_8 FILLER_24_553 ();
 sg13g2_decap_8 FILLER_24_560 ();
 sg13g2_decap_8 FILLER_24_567 ();
 sg13g2_decap_8 FILLER_24_574 ();
 sg13g2_decap_8 FILLER_24_581 ();
 sg13g2_decap_8 FILLER_24_588 ();
 sg13g2_decap_8 FILLER_24_595 ();
 sg13g2_decap_8 FILLER_24_602 ();
 sg13g2_decap_8 FILLER_24_609 ();
 sg13g2_decap_8 FILLER_24_616 ();
 sg13g2_decap_8 FILLER_24_623 ();
 sg13g2_decap_8 FILLER_24_630 ();
 sg13g2_decap_8 FILLER_24_637 ();
 sg13g2_decap_8 FILLER_24_644 ();
 sg13g2_decap_8 FILLER_24_651 ();
 sg13g2_decap_8 FILLER_24_658 ();
 sg13g2_decap_8 FILLER_24_665 ();
 sg13g2_decap_8 FILLER_24_672 ();
 sg13g2_decap_8 FILLER_24_679 ();
 sg13g2_decap_8 FILLER_24_686 ();
 sg13g2_decap_8 FILLER_24_693 ();
 sg13g2_decap_8 FILLER_24_700 ();
 sg13g2_decap_8 FILLER_24_707 ();
 sg13g2_decap_8 FILLER_24_714 ();
 sg13g2_decap_8 FILLER_24_721 ();
 sg13g2_decap_8 FILLER_24_728 ();
 sg13g2_decap_8 FILLER_24_735 ();
 sg13g2_decap_8 FILLER_24_742 ();
 sg13g2_decap_8 FILLER_24_749 ();
 sg13g2_decap_8 FILLER_24_756 ();
 sg13g2_decap_8 FILLER_24_763 ();
 sg13g2_decap_8 FILLER_24_770 ();
 sg13g2_decap_8 FILLER_24_777 ();
 sg13g2_decap_8 FILLER_24_784 ();
 sg13g2_decap_8 FILLER_24_791 ();
 sg13g2_decap_8 FILLER_24_798 ();
 sg13g2_decap_8 FILLER_24_805 ();
 sg13g2_decap_8 FILLER_24_812 ();
 sg13g2_decap_8 FILLER_24_819 ();
 sg13g2_decap_8 FILLER_24_826 ();
 sg13g2_decap_8 FILLER_24_833 ();
 sg13g2_decap_8 FILLER_24_840 ();
 sg13g2_decap_8 FILLER_24_847 ();
 sg13g2_decap_8 FILLER_24_854 ();
 sg13g2_fill_1 FILLER_24_861 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_decap_8 FILLER_25_406 ();
 sg13g2_decap_8 FILLER_25_413 ();
 sg13g2_decap_8 FILLER_25_420 ();
 sg13g2_decap_8 FILLER_25_427 ();
 sg13g2_decap_8 FILLER_25_434 ();
 sg13g2_decap_8 FILLER_25_441 ();
 sg13g2_decap_8 FILLER_25_448 ();
 sg13g2_decap_8 FILLER_25_455 ();
 sg13g2_decap_8 FILLER_25_462 ();
 sg13g2_decap_8 FILLER_25_469 ();
 sg13g2_decap_8 FILLER_25_476 ();
 sg13g2_decap_8 FILLER_25_483 ();
 sg13g2_decap_8 FILLER_25_490 ();
 sg13g2_decap_8 FILLER_25_497 ();
 sg13g2_decap_8 FILLER_25_504 ();
 sg13g2_decap_8 FILLER_25_511 ();
 sg13g2_decap_8 FILLER_25_518 ();
 sg13g2_decap_8 FILLER_25_525 ();
 sg13g2_decap_8 FILLER_25_532 ();
 sg13g2_decap_8 FILLER_25_539 ();
 sg13g2_decap_8 FILLER_25_546 ();
 sg13g2_decap_8 FILLER_25_553 ();
 sg13g2_decap_8 FILLER_25_560 ();
 sg13g2_decap_8 FILLER_25_567 ();
 sg13g2_decap_8 FILLER_25_574 ();
 sg13g2_decap_8 FILLER_25_581 ();
 sg13g2_decap_8 FILLER_25_588 ();
 sg13g2_decap_8 FILLER_25_595 ();
 sg13g2_decap_8 FILLER_25_602 ();
 sg13g2_decap_8 FILLER_25_609 ();
 sg13g2_decap_8 FILLER_25_616 ();
 sg13g2_decap_8 FILLER_25_623 ();
 sg13g2_decap_8 FILLER_25_630 ();
 sg13g2_decap_8 FILLER_25_637 ();
 sg13g2_decap_8 FILLER_25_644 ();
 sg13g2_decap_8 FILLER_25_651 ();
 sg13g2_decap_8 FILLER_25_658 ();
 sg13g2_decap_8 FILLER_25_665 ();
 sg13g2_decap_8 FILLER_25_672 ();
 sg13g2_decap_8 FILLER_25_679 ();
 sg13g2_decap_8 FILLER_25_686 ();
 sg13g2_decap_8 FILLER_25_693 ();
 sg13g2_decap_8 FILLER_25_700 ();
 sg13g2_decap_8 FILLER_25_707 ();
 sg13g2_decap_8 FILLER_25_714 ();
 sg13g2_decap_8 FILLER_25_721 ();
 sg13g2_decap_8 FILLER_25_728 ();
 sg13g2_decap_8 FILLER_25_735 ();
 sg13g2_decap_8 FILLER_25_742 ();
 sg13g2_decap_8 FILLER_25_749 ();
 sg13g2_decap_8 FILLER_25_756 ();
 sg13g2_decap_8 FILLER_25_763 ();
 sg13g2_decap_8 FILLER_25_770 ();
 sg13g2_decap_8 FILLER_25_777 ();
 sg13g2_decap_8 FILLER_25_784 ();
 sg13g2_decap_8 FILLER_25_791 ();
 sg13g2_decap_8 FILLER_25_798 ();
 sg13g2_decap_8 FILLER_25_805 ();
 sg13g2_decap_8 FILLER_25_812 ();
 sg13g2_decap_8 FILLER_25_819 ();
 sg13g2_decap_8 FILLER_25_826 ();
 sg13g2_decap_8 FILLER_25_833 ();
 sg13g2_decap_8 FILLER_25_840 ();
 sg13g2_decap_8 FILLER_25_847 ();
 sg13g2_decap_8 FILLER_25_854 ();
 sg13g2_fill_1 FILLER_25_861 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_decap_8 FILLER_26_406 ();
 sg13g2_decap_8 FILLER_26_413 ();
 sg13g2_decap_8 FILLER_26_420 ();
 sg13g2_decap_8 FILLER_26_427 ();
 sg13g2_decap_8 FILLER_26_434 ();
 sg13g2_decap_8 FILLER_26_441 ();
 sg13g2_decap_8 FILLER_26_448 ();
 sg13g2_decap_8 FILLER_26_455 ();
 sg13g2_decap_8 FILLER_26_462 ();
 sg13g2_decap_8 FILLER_26_469 ();
 sg13g2_decap_8 FILLER_26_476 ();
 sg13g2_decap_8 FILLER_26_483 ();
 sg13g2_decap_8 FILLER_26_490 ();
 sg13g2_decap_8 FILLER_26_497 ();
 sg13g2_decap_8 FILLER_26_504 ();
 sg13g2_decap_8 FILLER_26_511 ();
 sg13g2_decap_8 FILLER_26_518 ();
 sg13g2_decap_8 FILLER_26_525 ();
 sg13g2_decap_8 FILLER_26_532 ();
 sg13g2_decap_8 FILLER_26_539 ();
 sg13g2_decap_8 FILLER_26_546 ();
 sg13g2_decap_8 FILLER_26_553 ();
 sg13g2_decap_8 FILLER_26_560 ();
 sg13g2_decap_8 FILLER_26_567 ();
 sg13g2_decap_8 FILLER_26_574 ();
 sg13g2_decap_8 FILLER_26_581 ();
 sg13g2_decap_8 FILLER_26_588 ();
 sg13g2_decap_8 FILLER_26_595 ();
 sg13g2_decap_8 FILLER_26_602 ();
 sg13g2_decap_8 FILLER_26_609 ();
 sg13g2_decap_8 FILLER_26_616 ();
 sg13g2_decap_8 FILLER_26_623 ();
 sg13g2_decap_8 FILLER_26_630 ();
 sg13g2_decap_8 FILLER_26_637 ();
 sg13g2_decap_8 FILLER_26_644 ();
 sg13g2_decap_8 FILLER_26_651 ();
 sg13g2_decap_8 FILLER_26_658 ();
 sg13g2_decap_8 FILLER_26_665 ();
 sg13g2_decap_8 FILLER_26_672 ();
 sg13g2_decap_8 FILLER_26_679 ();
 sg13g2_decap_8 FILLER_26_686 ();
 sg13g2_decap_8 FILLER_26_693 ();
 sg13g2_decap_8 FILLER_26_700 ();
 sg13g2_decap_8 FILLER_26_707 ();
 sg13g2_decap_8 FILLER_26_714 ();
 sg13g2_decap_8 FILLER_26_721 ();
 sg13g2_decap_8 FILLER_26_728 ();
 sg13g2_decap_8 FILLER_26_735 ();
 sg13g2_decap_8 FILLER_26_742 ();
 sg13g2_decap_8 FILLER_26_749 ();
 sg13g2_decap_8 FILLER_26_756 ();
 sg13g2_decap_8 FILLER_26_763 ();
 sg13g2_decap_8 FILLER_26_770 ();
 sg13g2_decap_8 FILLER_26_777 ();
 sg13g2_decap_8 FILLER_26_784 ();
 sg13g2_decap_8 FILLER_26_791 ();
 sg13g2_decap_8 FILLER_26_798 ();
 sg13g2_decap_8 FILLER_26_805 ();
 sg13g2_decap_8 FILLER_26_812 ();
 sg13g2_decap_8 FILLER_26_819 ();
 sg13g2_decap_8 FILLER_26_826 ();
 sg13g2_decap_8 FILLER_26_833 ();
 sg13g2_decap_8 FILLER_26_840 ();
 sg13g2_decap_8 FILLER_26_847 ();
 sg13g2_decap_8 FILLER_26_854 ();
 sg13g2_fill_1 FILLER_26_861 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_decap_8 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_294 ();
 sg13g2_decap_8 FILLER_27_301 ();
 sg13g2_decap_8 FILLER_27_308 ();
 sg13g2_decap_8 FILLER_27_315 ();
 sg13g2_decap_8 FILLER_27_322 ();
 sg13g2_decap_8 FILLER_27_329 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_decap_8 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_decap_8 FILLER_27_406 ();
 sg13g2_decap_8 FILLER_27_413 ();
 sg13g2_decap_8 FILLER_27_420 ();
 sg13g2_decap_8 FILLER_27_427 ();
 sg13g2_decap_8 FILLER_27_434 ();
 sg13g2_decap_8 FILLER_27_441 ();
 sg13g2_decap_8 FILLER_27_448 ();
 sg13g2_decap_8 FILLER_27_455 ();
 sg13g2_decap_8 FILLER_27_462 ();
 sg13g2_decap_8 FILLER_27_469 ();
 sg13g2_decap_8 FILLER_27_476 ();
 sg13g2_decap_8 FILLER_27_483 ();
 sg13g2_decap_8 FILLER_27_490 ();
 sg13g2_decap_8 FILLER_27_497 ();
 sg13g2_decap_8 FILLER_27_504 ();
 sg13g2_decap_8 FILLER_27_511 ();
 sg13g2_decap_8 FILLER_27_518 ();
 sg13g2_decap_8 FILLER_27_525 ();
 sg13g2_decap_8 FILLER_27_532 ();
 sg13g2_decap_8 FILLER_27_539 ();
 sg13g2_decap_8 FILLER_27_546 ();
 sg13g2_decap_8 FILLER_27_553 ();
 sg13g2_decap_8 FILLER_27_560 ();
 sg13g2_decap_8 FILLER_27_567 ();
 sg13g2_decap_8 FILLER_27_574 ();
 sg13g2_decap_8 FILLER_27_581 ();
 sg13g2_decap_8 FILLER_27_588 ();
 sg13g2_decap_8 FILLER_27_599 ();
 sg13g2_decap_8 FILLER_27_606 ();
 sg13g2_decap_8 FILLER_27_613 ();
 sg13g2_decap_8 FILLER_27_620 ();
 sg13g2_decap_8 FILLER_27_627 ();
 sg13g2_decap_4 FILLER_27_634 ();
 sg13g2_decap_8 FILLER_27_651 ();
 sg13g2_decap_8 FILLER_27_658 ();
 sg13g2_decap_8 FILLER_27_665 ();
 sg13g2_decap_8 FILLER_27_672 ();
 sg13g2_decap_8 FILLER_27_679 ();
 sg13g2_decap_8 FILLER_27_686 ();
 sg13g2_decap_8 FILLER_27_693 ();
 sg13g2_decap_8 FILLER_27_700 ();
 sg13g2_decap_8 FILLER_27_707 ();
 sg13g2_decap_8 FILLER_27_714 ();
 sg13g2_decap_8 FILLER_27_721 ();
 sg13g2_decap_8 FILLER_27_728 ();
 sg13g2_decap_8 FILLER_27_735 ();
 sg13g2_decap_8 FILLER_27_742 ();
 sg13g2_decap_8 FILLER_27_749 ();
 sg13g2_decap_8 FILLER_27_756 ();
 sg13g2_decap_8 FILLER_27_763 ();
 sg13g2_decap_8 FILLER_27_770 ();
 sg13g2_decap_8 FILLER_27_777 ();
 sg13g2_decap_8 FILLER_27_784 ();
 sg13g2_decap_8 FILLER_27_791 ();
 sg13g2_decap_8 FILLER_27_798 ();
 sg13g2_decap_8 FILLER_27_805 ();
 sg13g2_decap_8 FILLER_27_812 ();
 sg13g2_decap_8 FILLER_27_819 ();
 sg13g2_decap_8 FILLER_27_826 ();
 sg13g2_decap_8 FILLER_27_833 ();
 sg13g2_decap_8 FILLER_27_840 ();
 sg13g2_decap_8 FILLER_27_847 ();
 sg13g2_decap_8 FILLER_27_854 ();
 sg13g2_fill_1 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_8 FILLER_28_245 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_decap_8 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_266 ();
 sg13g2_decap_8 FILLER_28_273 ();
 sg13g2_decap_8 FILLER_28_280 ();
 sg13g2_decap_8 FILLER_28_287 ();
 sg13g2_decap_8 FILLER_28_294 ();
 sg13g2_decap_8 FILLER_28_301 ();
 sg13g2_decap_8 FILLER_28_308 ();
 sg13g2_decap_8 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_322 ();
 sg13g2_decap_8 FILLER_28_329 ();
 sg13g2_decap_8 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_343 ();
 sg13g2_decap_8 FILLER_28_350 ();
 sg13g2_decap_8 FILLER_28_357 ();
 sg13g2_decap_8 FILLER_28_364 ();
 sg13g2_decap_8 FILLER_28_371 ();
 sg13g2_decap_8 FILLER_28_378 ();
 sg13g2_decap_8 FILLER_28_385 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_decap_8 FILLER_28_406 ();
 sg13g2_decap_4 FILLER_28_413 ();
 sg13g2_fill_1 FILLER_28_417 ();
 sg13g2_decap_8 FILLER_28_428 ();
 sg13g2_decap_4 FILLER_28_435 ();
 sg13g2_fill_2 FILLER_28_439 ();
 sg13g2_decap_8 FILLER_28_460 ();
 sg13g2_fill_1 FILLER_28_467 ();
 sg13g2_decap_8 FILLER_28_477 ();
 sg13g2_decap_8 FILLER_28_484 ();
 sg13g2_decap_8 FILLER_28_491 ();
 sg13g2_decap_8 FILLER_28_498 ();
 sg13g2_decap_8 FILLER_28_505 ();
 sg13g2_decap_8 FILLER_28_512 ();
 sg13g2_decap_8 FILLER_28_519 ();
 sg13g2_decap_8 FILLER_28_526 ();
 sg13g2_decap_8 FILLER_28_533 ();
 sg13g2_decap_4 FILLER_28_540 ();
 sg13g2_fill_1 FILLER_28_544 ();
 sg13g2_decap_8 FILLER_28_554 ();
 sg13g2_decap_8 FILLER_28_561 ();
 sg13g2_decap_8 FILLER_28_568 ();
 sg13g2_decap_4 FILLER_28_575 ();
 sg13g2_fill_1 FILLER_28_579 ();
 sg13g2_fill_2 FILLER_28_599 ();
 sg13g2_fill_1 FILLER_28_601 ();
 sg13g2_fill_2 FILLER_28_625 ();
 sg13g2_fill_2 FILLER_28_646 ();
 sg13g2_fill_1 FILLER_28_648 ();
 sg13g2_fill_1 FILLER_28_668 ();
 sg13g2_fill_1 FILLER_28_691 ();
 sg13g2_decap_8 FILLER_28_696 ();
 sg13g2_fill_2 FILLER_28_703 ();
 sg13g2_decap_8 FILLER_28_714 ();
 sg13g2_decap_8 FILLER_28_721 ();
 sg13g2_decap_8 FILLER_28_728 ();
 sg13g2_decap_8 FILLER_28_735 ();
 sg13g2_decap_8 FILLER_28_742 ();
 sg13g2_decap_8 FILLER_28_749 ();
 sg13g2_decap_8 FILLER_28_756 ();
 sg13g2_decap_8 FILLER_28_763 ();
 sg13g2_decap_8 FILLER_28_770 ();
 sg13g2_decap_8 FILLER_28_777 ();
 sg13g2_decap_8 FILLER_28_784 ();
 sg13g2_decap_8 FILLER_28_791 ();
 sg13g2_decap_8 FILLER_28_798 ();
 sg13g2_decap_8 FILLER_28_805 ();
 sg13g2_decap_8 FILLER_28_812 ();
 sg13g2_decap_8 FILLER_28_819 ();
 sg13g2_decap_8 FILLER_28_826 ();
 sg13g2_decap_8 FILLER_28_833 ();
 sg13g2_decap_8 FILLER_28_840 ();
 sg13g2_decap_8 FILLER_28_847 ();
 sg13g2_decap_8 FILLER_28_854 ();
 sg13g2_fill_1 FILLER_28_861 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_231 ();
 sg13g2_decap_8 FILLER_29_238 ();
 sg13g2_decap_8 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_252 ();
 sg13g2_decap_8 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_decap_8 FILLER_29_280 ();
 sg13g2_decap_8 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_29_294 ();
 sg13g2_decap_8 FILLER_29_301 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_decap_8 FILLER_29_322 ();
 sg13g2_decap_8 FILLER_29_329 ();
 sg13g2_decap_8 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_343 ();
 sg13g2_decap_8 FILLER_29_350 ();
 sg13g2_decap_8 FILLER_29_357 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_4 FILLER_29_399 ();
 sg13g2_fill_2 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_418 ();
 sg13g2_decap_8 FILLER_29_472 ();
 sg13g2_decap_8 FILLER_29_498 ();
 sg13g2_decap_8 FILLER_29_505 ();
 sg13g2_decap_4 FILLER_29_512 ();
 sg13g2_fill_1 FILLER_29_516 ();
 sg13g2_fill_2 FILLER_29_525 ();
 sg13g2_fill_1 FILLER_29_527 ();
 sg13g2_decap_8 FILLER_29_727 ();
 sg13g2_decap_8 FILLER_29_734 ();
 sg13g2_decap_8 FILLER_29_741 ();
 sg13g2_decap_8 FILLER_29_748 ();
 sg13g2_decap_8 FILLER_29_755 ();
 sg13g2_decap_8 FILLER_29_762 ();
 sg13g2_decap_8 FILLER_29_769 ();
 sg13g2_decap_8 FILLER_29_776 ();
 sg13g2_decap_8 FILLER_29_783 ();
 sg13g2_decap_8 FILLER_29_790 ();
 sg13g2_decap_8 FILLER_29_797 ();
 sg13g2_decap_8 FILLER_29_804 ();
 sg13g2_decap_8 FILLER_29_811 ();
 sg13g2_decap_8 FILLER_29_818 ();
 sg13g2_decap_8 FILLER_29_825 ();
 sg13g2_decap_8 FILLER_29_832 ();
 sg13g2_decap_8 FILLER_29_839 ();
 sg13g2_decap_8 FILLER_29_846 ();
 sg13g2_decap_8 FILLER_29_853 ();
 sg13g2_fill_2 FILLER_29_860 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_decap_4 FILLER_30_252 ();
 sg13g2_fill_2 FILLER_30_256 ();
 sg13g2_decap_8 FILLER_30_267 ();
 sg13g2_decap_8 FILLER_30_274 ();
 sg13g2_decap_8 FILLER_30_281 ();
 sg13g2_decap_8 FILLER_30_288 ();
 sg13g2_decap_8 FILLER_30_295 ();
 sg13g2_decap_8 FILLER_30_302 ();
 sg13g2_decap_8 FILLER_30_309 ();
 sg13g2_decap_8 FILLER_30_316 ();
 sg13g2_decap_8 FILLER_30_323 ();
 sg13g2_decap_4 FILLER_30_330 ();
 sg13g2_fill_2 FILLER_30_334 ();
 sg13g2_decap_8 FILLER_30_354 ();
 sg13g2_decap_8 FILLER_30_361 ();
 sg13g2_decap_8 FILLER_30_368 ();
 sg13g2_decap_8 FILLER_30_375 ();
 sg13g2_decap_8 FILLER_30_382 ();
 sg13g2_decap_4 FILLER_30_389 ();
 sg13g2_fill_1 FILLER_30_393 ();
 sg13g2_fill_1 FILLER_30_457 ();
 sg13g2_decap_4 FILLER_30_507 ();
 sg13g2_decap_4 FILLER_30_537 ();
 sg13g2_fill_2 FILLER_30_586 ();
 sg13g2_fill_1 FILLER_30_629 ();
 sg13g2_fill_2 FILLER_30_649 ();
 sg13g2_fill_1 FILLER_30_651 ();
 sg13g2_fill_2 FILLER_30_707 ();
 sg13g2_fill_1 FILLER_30_709 ();
 sg13g2_decap_8 FILLER_30_736 ();
 sg13g2_decap_8 FILLER_30_743 ();
 sg13g2_decap_8 FILLER_30_750 ();
 sg13g2_decap_8 FILLER_30_757 ();
 sg13g2_decap_8 FILLER_30_764 ();
 sg13g2_decap_8 FILLER_30_771 ();
 sg13g2_decap_8 FILLER_30_778 ();
 sg13g2_decap_8 FILLER_30_785 ();
 sg13g2_decap_8 FILLER_30_792 ();
 sg13g2_decap_8 FILLER_30_799 ();
 sg13g2_decap_8 FILLER_30_806 ();
 sg13g2_decap_8 FILLER_30_813 ();
 sg13g2_decap_8 FILLER_30_820 ();
 sg13g2_decap_8 FILLER_30_827 ();
 sg13g2_decap_8 FILLER_30_834 ();
 sg13g2_decap_8 FILLER_30_841 ();
 sg13g2_decap_8 FILLER_30_848 ();
 sg13g2_decap_8 FILLER_30_855 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_4 FILLER_31_238 ();
 sg13g2_fill_1 FILLER_31_242 ();
 sg13g2_decap_8 FILLER_31_247 ();
 sg13g2_fill_1 FILLER_31_254 ();
 sg13g2_decap_8 FILLER_31_278 ();
 sg13g2_decap_8 FILLER_31_285 ();
 sg13g2_decap_8 FILLER_31_292 ();
 sg13g2_decap_8 FILLER_31_299 ();
 sg13g2_decap_8 FILLER_31_306 ();
 sg13g2_decap_8 FILLER_31_313 ();
 sg13g2_decap_8 FILLER_31_320 ();
 sg13g2_fill_2 FILLER_31_327 ();
 sg13g2_fill_1 FILLER_31_447 ();
 sg13g2_fill_2 FILLER_31_467 ();
 sg13g2_fill_1 FILLER_31_469 ();
 sg13g2_decap_4 FILLER_31_562 ();
 sg13g2_fill_1 FILLER_31_566 ();
 sg13g2_fill_2 FILLER_31_575 ();
 sg13g2_fill_1 FILLER_31_577 ();
 sg13g2_decap_4 FILLER_31_692 ();
 sg13g2_decap_4 FILLER_31_746 ();
 sg13g2_decap_8 FILLER_31_773 ();
 sg13g2_decap_8 FILLER_31_780 ();
 sg13g2_decap_8 FILLER_31_787 ();
 sg13g2_decap_8 FILLER_31_794 ();
 sg13g2_decap_8 FILLER_31_801 ();
 sg13g2_decap_8 FILLER_31_808 ();
 sg13g2_decap_8 FILLER_31_815 ();
 sg13g2_decap_8 FILLER_31_822 ();
 sg13g2_decap_8 FILLER_31_829 ();
 sg13g2_decap_8 FILLER_31_836 ();
 sg13g2_decap_8 FILLER_31_843 ();
 sg13g2_decap_8 FILLER_31_850 ();
 sg13g2_decap_4 FILLER_31_857 ();
 sg13g2_fill_1 FILLER_31_861 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_fill_1 FILLER_32_231 ();
 sg13g2_fill_2 FILLER_32_258 ();
 sg13g2_fill_1 FILLER_32_260 ();
 sg13g2_decap_8 FILLER_32_296 ();
 sg13g2_fill_2 FILLER_32_303 ();
 sg13g2_decap_4 FILLER_32_313 ();
 sg13g2_fill_2 FILLER_32_317 ();
 sg13g2_fill_1 FILLER_32_352 ();
 sg13g2_fill_1 FILLER_32_363 ();
 sg13g2_fill_1 FILLER_32_387 ();
 sg13g2_decap_4 FILLER_32_424 ();
 sg13g2_fill_2 FILLER_32_490 ();
 sg13g2_fill_1 FILLER_32_518 ();
 sg13g2_fill_2 FILLER_32_609 ();
 sg13g2_fill_1 FILLER_32_611 ();
 sg13g2_fill_1 FILLER_32_634 ();
 sg13g2_fill_2 FILLER_32_675 ();
 sg13g2_fill_1 FILLER_32_757 ();
 sg13g2_decap_8 FILLER_32_784 ();
 sg13g2_decap_8 FILLER_32_791 ();
 sg13g2_decap_8 FILLER_32_798 ();
 sg13g2_decap_8 FILLER_32_805 ();
 sg13g2_decap_8 FILLER_32_812 ();
 sg13g2_decap_8 FILLER_32_819 ();
 sg13g2_decap_8 FILLER_32_826 ();
 sg13g2_decap_8 FILLER_32_833 ();
 sg13g2_decap_8 FILLER_32_840 ();
 sg13g2_decap_8 FILLER_32_847 ();
 sg13g2_decap_8 FILLER_32_854 ();
 sg13g2_fill_1 FILLER_32_861 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_fill_2 FILLER_33_224 ();
 sg13g2_fill_2 FILLER_33_267 ();
 sg13g2_fill_2 FILLER_33_305 ();
 sg13g2_fill_1 FILLER_33_333 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_decap_4 FILLER_33_416 ();
 sg13g2_fill_2 FILLER_33_466 ();
 sg13g2_fill_1 FILLER_33_468 ();
 sg13g2_decap_4 FILLER_33_473 ();
 sg13g2_fill_2 FILLER_33_507 ();
 sg13g2_fill_1 FILLER_33_509 ();
 sg13g2_fill_2 FILLER_33_518 ();
 sg13g2_fill_1 FILLER_33_520 ();
 sg13g2_decap_8 FILLER_33_557 ();
 sg13g2_decap_4 FILLER_33_564 ();
 sg13g2_fill_1 FILLER_33_568 ();
 sg13g2_fill_2 FILLER_33_592 ();
 sg13g2_fill_1 FILLER_33_594 ();
 sg13g2_fill_1 FILLER_33_635 ();
 sg13g2_fill_1 FILLER_33_645 ();
 sg13g2_fill_2 FILLER_33_682 ();
 sg13g2_fill_2 FILLER_33_717 ();
 sg13g2_fill_1 FILLER_33_719 ();
 sg13g2_decap_8 FILLER_33_743 ();
 sg13g2_fill_1 FILLER_33_750 ();
 sg13g2_decap_8 FILLER_33_796 ();
 sg13g2_decap_8 FILLER_33_803 ();
 sg13g2_decap_8 FILLER_33_810 ();
 sg13g2_decap_8 FILLER_33_817 ();
 sg13g2_decap_8 FILLER_33_824 ();
 sg13g2_decap_8 FILLER_33_831 ();
 sg13g2_decap_8 FILLER_33_838 ();
 sg13g2_decap_8 FILLER_33_845 ();
 sg13g2_decap_8 FILLER_33_852 ();
 sg13g2_fill_2 FILLER_33_859 ();
 sg13g2_fill_1 FILLER_33_861 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_fill_2 FILLER_34_224 ();
 sg13g2_fill_2 FILLER_34_294 ();
 sg13g2_fill_1 FILLER_34_317 ();
 sg13g2_fill_2 FILLER_34_336 ();
 sg13g2_fill_1 FILLER_34_338 ();
 sg13g2_fill_2 FILLER_34_376 ();
 sg13g2_fill_1 FILLER_34_486 ();
 sg13g2_fill_2 FILLER_34_507 ();
 sg13g2_decap_8 FILLER_34_559 ();
 sg13g2_fill_1 FILLER_34_566 ();
 sg13g2_fill_2 FILLER_34_624 ();
 sg13g2_decap_4 FILLER_34_679 ();
 sg13g2_fill_2 FILLER_34_683 ();
 sg13g2_fill_1 FILLER_34_689 ();
 sg13g2_decap_4 FILLER_34_742 ();
 sg13g2_decap_8 FILLER_34_787 ();
 sg13g2_decap_8 FILLER_34_794 ();
 sg13g2_decap_8 FILLER_34_801 ();
 sg13g2_decap_8 FILLER_34_808 ();
 sg13g2_decap_8 FILLER_34_815 ();
 sg13g2_decap_8 FILLER_34_822 ();
 sg13g2_decap_8 FILLER_34_829 ();
 sg13g2_decap_8 FILLER_34_836 ();
 sg13g2_decap_8 FILLER_34_843 ();
 sg13g2_decap_8 FILLER_34_850 ();
 sg13g2_decap_4 FILLER_34_857 ();
 sg13g2_fill_1 FILLER_34_861 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_fill_2 FILLER_35_224 ();
 sg13g2_decap_4 FILLER_35_284 ();
 sg13g2_fill_1 FILLER_35_314 ();
 sg13g2_fill_1 FILLER_35_330 ();
 sg13g2_fill_1 FILLER_35_363 ();
 sg13g2_decap_8 FILLER_35_387 ();
 sg13g2_decap_4 FILLER_35_394 ();
 sg13g2_fill_1 FILLER_35_398 ();
 sg13g2_fill_2 FILLER_35_417 ();
 sg13g2_fill_1 FILLER_35_432 ();
 sg13g2_fill_2 FILLER_35_452 ();
 sg13g2_fill_2 FILLER_35_517 ();
 sg13g2_fill_1 FILLER_35_623 ();
 sg13g2_fill_2 FILLER_35_643 ();
 sg13g2_fill_1 FILLER_35_645 ();
 sg13g2_fill_1 FILLER_35_672 ();
 sg13g2_decap_8 FILLER_35_782 ();
 sg13g2_decap_8 FILLER_35_789 ();
 sg13g2_decap_8 FILLER_35_796 ();
 sg13g2_decap_8 FILLER_35_803 ();
 sg13g2_decap_8 FILLER_35_810 ();
 sg13g2_decap_8 FILLER_35_817 ();
 sg13g2_decap_8 FILLER_35_824 ();
 sg13g2_decap_8 FILLER_35_831 ();
 sg13g2_decap_8 FILLER_35_838 ();
 sg13g2_decap_8 FILLER_35_845 ();
 sg13g2_decap_8 FILLER_35_852 ();
 sg13g2_fill_2 FILLER_35_859 ();
 sg13g2_fill_1 FILLER_35_861 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_fill_2 FILLER_36_224 ();
 sg13g2_fill_1 FILLER_36_226 ();
 sg13g2_decap_4 FILLER_36_287 ();
 sg13g2_fill_2 FILLER_36_313 ();
 sg13g2_fill_2 FILLER_36_437 ();
 sg13g2_fill_1 FILLER_36_439 ();
 sg13g2_fill_2 FILLER_36_464 ();
 sg13g2_fill_2 FILLER_36_475 ();
 sg13g2_fill_2 FILLER_36_490 ();
 sg13g2_fill_1 FILLER_36_531 ();
 sg13g2_fill_2 FILLER_36_555 ();
 sg13g2_decap_4 FILLER_36_570 ();
 sg13g2_fill_1 FILLER_36_574 ();
 sg13g2_fill_2 FILLER_36_579 ();
 sg13g2_fill_1 FILLER_36_581 ();
 sg13g2_fill_2 FILLER_36_708 ();
 sg13g2_fill_1 FILLER_36_710 ();
 sg13g2_fill_2 FILLER_36_724 ();
 sg13g2_fill_1 FILLER_36_726 ();
 sg13g2_decap_4 FILLER_36_746 ();
 sg13g2_decap_8 FILLER_36_786 ();
 sg13g2_decap_8 FILLER_36_793 ();
 sg13g2_decap_8 FILLER_36_800 ();
 sg13g2_decap_8 FILLER_36_807 ();
 sg13g2_decap_8 FILLER_36_814 ();
 sg13g2_decap_8 FILLER_36_821 ();
 sg13g2_decap_8 FILLER_36_828 ();
 sg13g2_decap_8 FILLER_36_835 ();
 sg13g2_decap_8 FILLER_36_842 ();
 sg13g2_decap_8 FILLER_36_849 ();
 sg13g2_decap_4 FILLER_36_856 ();
 sg13g2_fill_2 FILLER_36_860 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_66 ();
 sg13g2_decap_8 FILLER_37_73 ();
 sg13g2_decap_8 FILLER_37_80 ();
 sg13g2_fill_2 FILLER_37_87 ();
 sg13g2_fill_1 FILLER_37_89 ();
 sg13g2_fill_2 FILLER_37_93 ();
 sg13g2_decap_8 FILLER_37_99 ();
 sg13g2_decap_8 FILLER_37_109 ();
 sg13g2_decap_8 FILLER_37_116 ();
 sg13g2_fill_2 FILLER_37_123 ();
 sg13g2_fill_2 FILLER_37_128 ();
 sg13g2_decap_8 FILLER_37_136 ();
 sg13g2_decap_8 FILLER_37_143 ();
 sg13g2_decap_8 FILLER_37_150 ();
 sg13g2_decap_8 FILLER_37_157 ();
 sg13g2_decap_8 FILLER_37_164 ();
 sg13g2_decap_8 FILLER_37_171 ();
 sg13g2_decap_8 FILLER_37_178 ();
 sg13g2_decap_8 FILLER_37_185 ();
 sg13g2_decap_8 FILLER_37_192 ();
 sg13g2_decap_8 FILLER_37_199 ();
 sg13g2_decap_8 FILLER_37_206 ();
 sg13g2_decap_8 FILLER_37_213 ();
 sg13g2_fill_2 FILLER_37_220 ();
 sg13g2_fill_1 FILLER_37_222 ();
 sg13g2_decap_4 FILLER_37_259 ();
 sg13g2_fill_2 FILLER_37_298 ();
 sg13g2_fill_1 FILLER_37_300 ();
 sg13g2_fill_2 FILLER_37_315 ();
 sg13g2_fill_1 FILLER_37_317 ();
 sg13g2_decap_8 FILLER_37_331 ();
 sg13g2_decap_4 FILLER_37_338 ();
 sg13g2_fill_1 FILLER_37_342 ();
 sg13g2_fill_2 FILLER_37_352 ();
 sg13g2_fill_1 FILLER_37_354 ();
 sg13g2_fill_2 FILLER_37_381 ();
 sg13g2_fill_2 FILLER_37_413 ();
 sg13g2_decap_4 FILLER_37_419 ();
 sg13g2_fill_1 FILLER_37_423 ();
 sg13g2_fill_1 FILLER_37_454 ();
 sg13g2_fill_1 FILLER_37_485 ();
 sg13g2_fill_1 FILLER_37_536 ();
 sg13g2_fill_1 FILLER_37_563 ();
 sg13g2_fill_1 FILLER_37_675 ();
 sg13g2_decap_8 FILLER_37_787 ();
 sg13g2_decap_8 FILLER_37_794 ();
 sg13g2_decap_8 FILLER_37_801 ();
 sg13g2_decap_8 FILLER_37_808 ();
 sg13g2_decap_8 FILLER_37_815 ();
 sg13g2_decap_8 FILLER_37_822 ();
 sg13g2_decap_8 FILLER_37_829 ();
 sg13g2_decap_8 FILLER_37_836 ();
 sg13g2_decap_8 FILLER_37_843 ();
 sg13g2_decap_8 FILLER_37_850 ();
 sg13g2_decap_4 FILLER_37_857 ();
 sg13g2_fill_1 FILLER_37_861 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_38 ();
 sg13g2_fill_2 FILLER_38_45 ();
 sg13g2_fill_1 FILLER_38_47 ();
 sg13g2_fill_2 FILLER_38_81 ();
 sg13g2_fill_1 FILLER_38_83 ();
 sg13g2_fill_2 FILLER_38_108 ();
 sg13g2_fill_1 FILLER_38_136 ();
 sg13g2_decap_8 FILLER_38_143 ();
 sg13g2_decap_8 FILLER_38_150 ();
 sg13g2_decap_8 FILLER_38_157 ();
 sg13g2_decap_8 FILLER_38_164 ();
 sg13g2_decap_8 FILLER_38_171 ();
 sg13g2_decap_8 FILLER_38_178 ();
 sg13g2_decap_8 FILLER_38_185 ();
 sg13g2_decap_8 FILLER_38_192 ();
 sg13g2_decap_8 FILLER_38_199 ();
 sg13g2_decap_8 FILLER_38_206 ();
 sg13g2_decap_8 FILLER_38_213 ();
 sg13g2_decap_8 FILLER_38_220 ();
 sg13g2_fill_2 FILLER_38_227 ();
 sg13g2_fill_1 FILLER_38_229 ();
 sg13g2_fill_1 FILLER_38_266 ();
 sg13g2_fill_2 FILLER_38_355 ();
 sg13g2_fill_2 FILLER_38_431 ();
 sg13g2_fill_1 FILLER_38_433 ();
 sg13g2_fill_1 FILLER_38_443 ();
 sg13g2_fill_1 FILLER_38_454 ();
 sg13g2_fill_2 FILLER_38_465 ();
 sg13g2_fill_1 FILLER_38_515 ();
 sg13g2_decap_4 FILLER_38_562 ();
 sg13g2_fill_1 FILLER_38_628 ();
 sg13g2_fill_2 FILLER_38_653 ();
 sg13g2_fill_2 FILLER_38_668 ();
 sg13g2_fill_1 FILLER_38_670 ();
 sg13g2_fill_1 FILLER_38_720 ();
 sg13g2_decap_8 FILLER_38_787 ();
 sg13g2_decap_8 FILLER_38_794 ();
 sg13g2_decap_8 FILLER_38_801 ();
 sg13g2_decap_8 FILLER_38_808 ();
 sg13g2_decap_8 FILLER_38_815 ();
 sg13g2_decap_8 FILLER_38_822 ();
 sg13g2_decap_8 FILLER_38_829 ();
 sg13g2_decap_8 FILLER_38_836 ();
 sg13g2_decap_8 FILLER_38_843 ();
 sg13g2_decap_8 FILLER_38_850 ();
 sg13g2_decap_4 FILLER_38_857 ();
 sg13g2_fill_1 FILLER_38_861 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_fill_2 FILLER_39_28 ();
 sg13g2_fill_1 FILLER_39_30 ();
 sg13g2_fill_1 FILLER_39_57 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_196 ();
 sg13g2_fill_1 FILLER_39_203 ();
 sg13g2_decap_4 FILLER_39_214 ();
 sg13g2_fill_2 FILLER_39_218 ();
 sg13g2_decap_4 FILLER_39_286 ();
 sg13g2_decap_4 FILLER_39_300 ();
 sg13g2_fill_2 FILLER_39_304 ();
 sg13g2_fill_2 FILLER_39_315 ();
 sg13g2_decap_8 FILLER_39_321 ();
 sg13g2_decap_8 FILLER_39_328 ();
 sg13g2_fill_2 FILLER_39_366 ();
 sg13g2_fill_1 FILLER_39_387 ();
 sg13g2_fill_2 FILLER_39_482 ();
 sg13g2_fill_1 FILLER_39_484 ();
 sg13g2_fill_2 FILLER_39_521 ();
 sg13g2_fill_1 FILLER_39_523 ();
 sg13g2_fill_2 FILLER_39_584 ();
 sg13g2_fill_1 FILLER_39_586 ();
 sg13g2_fill_2 FILLER_39_601 ();
 sg13g2_fill_2 FILLER_39_639 ();
 sg13g2_fill_1 FILLER_39_641 ();
 sg13g2_fill_2 FILLER_39_672 ();
 sg13g2_fill_1 FILLER_39_674 ();
 sg13g2_fill_1 FILLER_39_705 ();
 sg13g2_fill_2 FILLER_39_741 ();
 sg13g2_fill_1 FILLER_39_743 ();
 sg13g2_fill_2 FILLER_39_748 ();
 sg13g2_fill_1 FILLER_39_750 ();
 sg13g2_decap_8 FILLER_39_779 ();
 sg13g2_decap_8 FILLER_39_786 ();
 sg13g2_decap_8 FILLER_39_793 ();
 sg13g2_decap_8 FILLER_39_800 ();
 sg13g2_decap_8 FILLER_39_807 ();
 sg13g2_decap_8 FILLER_39_814 ();
 sg13g2_decap_8 FILLER_39_821 ();
 sg13g2_decap_8 FILLER_39_828 ();
 sg13g2_decap_8 FILLER_39_835 ();
 sg13g2_decap_8 FILLER_39_842 ();
 sg13g2_decap_8 FILLER_39_849 ();
 sg13g2_decap_4 FILLER_39_856 ();
 sg13g2_fill_2 FILLER_39_860 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_fill_2 FILLER_40_28 ();
 sg13g2_fill_1 FILLER_40_30 ();
 sg13g2_decap_4 FILLER_40_35 ();
 sg13g2_fill_1 FILLER_40_71 ();
 sg13g2_fill_2 FILLER_40_95 ();
 sg13g2_decap_4 FILLER_40_101 ();
 sg13g2_fill_1 FILLER_40_105 ();
 sg13g2_fill_1 FILLER_40_129 ();
 sg13g2_fill_1 FILLER_40_165 ();
 sg13g2_fill_2 FILLER_40_172 ();
 sg13g2_fill_1 FILLER_40_174 ();
 sg13g2_decap_4 FILLER_40_178 ();
 sg13g2_decap_8 FILLER_40_191 ();
 sg13g2_fill_2 FILLER_40_198 ();
 sg13g2_fill_1 FILLER_40_200 ();
 sg13g2_decap_8 FILLER_40_283 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_40_413 ();
 sg13g2_decap_4 FILLER_40_429 ();
 sg13g2_fill_2 FILLER_40_455 ();
 sg13g2_fill_2 FILLER_40_511 ();
 sg13g2_fill_1 FILLER_40_513 ();
 sg13g2_fill_1 FILLER_40_522 ();
 sg13g2_fill_1 FILLER_40_578 ();
 sg13g2_fill_1 FILLER_40_588 ();
 sg13g2_fill_2 FILLER_40_629 ();
 sg13g2_fill_1 FILLER_40_631 ();
 sg13g2_decap_8 FILLER_40_662 ();
 sg13g2_fill_1 FILLER_40_669 ();
 sg13g2_fill_2 FILLER_40_706 ();
 sg13g2_fill_1 FILLER_40_708 ();
 sg13g2_fill_1 FILLER_40_727 ();
 sg13g2_decap_8 FILLER_40_785 ();
 sg13g2_decap_8 FILLER_40_792 ();
 sg13g2_decap_8 FILLER_40_799 ();
 sg13g2_decap_8 FILLER_40_806 ();
 sg13g2_decap_8 FILLER_40_813 ();
 sg13g2_decap_8 FILLER_40_820 ();
 sg13g2_decap_8 FILLER_40_827 ();
 sg13g2_decap_8 FILLER_40_834 ();
 sg13g2_decap_8 FILLER_40_841 ();
 sg13g2_decap_8 FILLER_40_848 ();
 sg13g2_decap_8 FILLER_40_855 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_7 ();
 sg13g2_fill_1 FILLER_41_9 ();
 sg13g2_fill_2 FILLER_41_138 ();
 sg13g2_fill_2 FILLER_41_166 ();
 sg13g2_fill_2 FILLER_41_200 ();
 sg13g2_fill_1 FILLER_41_202 ();
 sg13g2_fill_2 FILLER_41_212 ();
 sg13g2_fill_2 FILLER_41_241 ();
 sg13g2_fill_1 FILLER_41_251 ();
 sg13g2_fill_1 FILLER_41_291 ();
 sg13g2_fill_1 FILLER_41_295 ();
 sg13g2_fill_2 FILLER_41_312 ();
 sg13g2_fill_1 FILLER_41_343 ();
 sg13g2_fill_2 FILLER_41_367 ();
 sg13g2_decap_8 FILLER_41_379 ();
 sg13g2_fill_2 FILLER_41_462 ();
 sg13g2_fill_2 FILLER_41_542 ();
 sg13g2_fill_1 FILLER_41_544 ();
 sg13g2_fill_2 FILLER_41_594 ();
 sg13g2_fill_1 FILLER_41_596 ();
 sg13g2_decap_8 FILLER_41_619 ();
 sg13g2_fill_2 FILLER_41_626 ();
 sg13g2_fill_1 FILLER_41_655 ();
 sg13g2_fill_2 FILLER_41_661 ();
 sg13g2_fill_1 FILLER_41_699 ();
 sg13g2_fill_2 FILLER_41_745 ();
 sg13g2_fill_1 FILLER_41_747 ();
 sg13g2_decap_8 FILLER_41_793 ();
 sg13g2_decap_8 FILLER_41_800 ();
 sg13g2_decap_8 FILLER_41_807 ();
 sg13g2_decap_8 FILLER_41_814 ();
 sg13g2_decap_8 FILLER_41_821 ();
 sg13g2_decap_8 FILLER_41_828 ();
 sg13g2_decap_8 FILLER_41_835 ();
 sg13g2_decap_8 FILLER_41_842 ();
 sg13g2_decap_8 FILLER_41_849 ();
 sg13g2_decap_4 FILLER_41_856 ();
 sg13g2_fill_2 FILLER_41_860 ();
 sg13g2_fill_1 FILLER_42_83 ();
 sg13g2_fill_2 FILLER_42_101 ();
 sg13g2_fill_1 FILLER_42_113 ();
 sg13g2_fill_1 FILLER_42_127 ();
 sg13g2_fill_1 FILLER_42_146 ();
 sg13g2_fill_1 FILLER_42_177 ();
 sg13g2_decap_8 FILLER_42_424 ();
 sg13g2_fill_2 FILLER_42_431 ();
 sg13g2_fill_1 FILLER_42_433 ();
 sg13g2_fill_1 FILLER_42_477 ();
 sg13g2_fill_2 FILLER_42_487 ();
 sg13g2_fill_2 FILLER_42_498 ();
 sg13g2_fill_2 FILLER_42_519 ();
 sg13g2_fill_1 FILLER_42_521 ();
 sg13g2_fill_2 FILLER_42_532 ();
 sg13g2_fill_1 FILLER_42_534 ();
 sg13g2_fill_2 FILLER_42_579 ();
 sg13g2_fill_2 FILLER_42_710 ();
 sg13g2_fill_1 FILLER_42_712 ();
 sg13g2_fill_2 FILLER_42_749 ();
 sg13g2_decap_8 FILLER_42_787 ();
 sg13g2_decap_8 FILLER_42_794 ();
 sg13g2_decap_8 FILLER_42_801 ();
 sg13g2_decap_8 FILLER_42_808 ();
 sg13g2_decap_8 FILLER_42_815 ();
 sg13g2_decap_8 FILLER_42_822 ();
 sg13g2_decap_8 FILLER_42_829 ();
 sg13g2_decap_8 FILLER_42_836 ();
 sg13g2_decap_8 FILLER_42_843 ();
 sg13g2_decap_8 FILLER_42_850 ();
 sg13g2_decap_4 FILLER_42_857 ();
 sg13g2_fill_1 FILLER_42_861 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_fill_1 FILLER_43_14 ();
 sg13g2_fill_2 FILLER_43_51 ();
 sg13g2_fill_2 FILLER_43_77 ();
 sg13g2_fill_1 FILLER_43_117 ();
 sg13g2_decap_4 FILLER_43_137 ();
 sg13g2_fill_2 FILLER_43_141 ();
 sg13g2_fill_2 FILLER_43_151 ();
 sg13g2_fill_2 FILLER_43_209 ();
 sg13g2_fill_1 FILLER_43_218 ();
 sg13g2_fill_2 FILLER_43_256 ();
 sg13g2_fill_1 FILLER_43_264 ();
 sg13g2_fill_1 FILLER_43_274 ();
 sg13g2_fill_2 FILLER_43_316 ();
 sg13g2_fill_2 FILLER_43_330 ();
 sg13g2_fill_1 FILLER_43_358 ();
 sg13g2_fill_2 FILLER_43_404 ();
 sg13g2_fill_1 FILLER_43_406 ();
 sg13g2_fill_1 FILLER_43_425 ();
 sg13g2_fill_2 FILLER_43_492 ();
 sg13g2_decap_4 FILLER_43_520 ();
 sg13g2_decap_4 FILLER_43_554 ();
 sg13g2_fill_1 FILLER_43_558 ();
 sg13g2_fill_1 FILLER_43_569 ();
 sg13g2_fill_1 FILLER_43_623 ();
 sg13g2_fill_1 FILLER_43_634 ();
 sg13g2_fill_2 FILLER_43_671 ();
 sg13g2_fill_2 FILLER_43_745 ();
 sg13g2_decap_8 FILLER_43_783 ();
 sg13g2_decap_8 FILLER_43_790 ();
 sg13g2_decap_8 FILLER_43_797 ();
 sg13g2_decap_8 FILLER_43_804 ();
 sg13g2_decap_8 FILLER_43_811 ();
 sg13g2_decap_8 FILLER_43_818 ();
 sg13g2_decap_8 FILLER_43_825 ();
 sg13g2_decap_8 FILLER_43_832 ();
 sg13g2_decap_8 FILLER_43_839 ();
 sg13g2_decap_8 FILLER_43_846 ();
 sg13g2_decap_8 FILLER_43_853 ();
 sg13g2_fill_2 FILLER_43_860 ();
 sg13g2_decap_4 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_34 ();
 sg13g2_fill_2 FILLER_44_51 ();
 sg13g2_fill_1 FILLER_44_154 ();
 sg13g2_fill_2 FILLER_44_164 ();
 sg13g2_fill_2 FILLER_44_182 ();
 sg13g2_decap_4 FILLER_44_205 ();
 sg13g2_fill_2 FILLER_44_209 ();
 sg13g2_fill_1 FILLER_44_234 ();
 sg13g2_fill_2 FILLER_44_274 ();
 sg13g2_fill_1 FILLER_44_313 ();
 sg13g2_decap_4 FILLER_44_327 ();
 sg13g2_fill_1 FILLER_44_331 ();
 sg13g2_fill_2 FILLER_44_515 ();
 sg13g2_decap_4 FILLER_44_539 ();
 sg13g2_fill_2 FILLER_44_543 ();
 sg13g2_decap_4 FILLER_44_616 ();
 sg13g2_fill_2 FILLER_44_620 ();
 sg13g2_fill_1 FILLER_44_657 ();
 sg13g2_decap_8 FILLER_44_784 ();
 sg13g2_decap_8 FILLER_44_791 ();
 sg13g2_decap_8 FILLER_44_798 ();
 sg13g2_decap_8 FILLER_44_805 ();
 sg13g2_decap_8 FILLER_44_812 ();
 sg13g2_decap_8 FILLER_44_819 ();
 sg13g2_decap_8 FILLER_44_826 ();
 sg13g2_decap_8 FILLER_44_833 ();
 sg13g2_decap_8 FILLER_44_840 ();
 sg13g2_decap_8 FILLER_44_847 ();
 sg13g2_decap_8 FILLER_44_854 ();
 sg13g2_fill_1 FILLER_44_861 ();
 sg13g2_fill_1 FILLER_45_83 ();
 sg13g2_fill_2 FILLER_45_110 ();
 sg13g2_fill_1 FILLER_45_112 ();
 sg13g2_fill_1 FILLER_45_134 ();
 sg13g2_fill_1 FILLER_45_215 ();
 sg13g2_fill_2 FILLER_45_331 ();
 sg13g2_fill_1 FILLER_45_357 ();
 sg13g2_fill_2 FILLER_45_376 ();
 sg13g2_fill_1 FILLER_45_458 ();
 sg13g2_fill_1 FILLER_45_480 ();
 sg13g2_fill_2 FILLER_45_507 ();
 sg13g2_fill_1 FILLER_45_509 ();
 sg13g2_fill_1 FILLER_45_696 ();
 sg13g2_fill_2 FILLER_45_732 ();
 sg13g2_fill_1 FILLER_45_734 ();
 sg13g2_decap_8 FILLER_45_758 ();
 sg13g2_fill_1 FILLER_45_765 ();
 sg13g2_decap_8 FILLER_45_779 ();
 sg13g2_decap_8 FILLER_45_786 ();
 sg13g2_decap_8 FILLER_45_793 ();
 sg13g2_decap_8 FILLER_45_800 ();
 sg13g2_decap_8 FILLER_45_807 ();
 sg13g2_decap_8 FILLER_45_814 ();
 sg13g2_decap_8 FILLER_45_821 ();
 sg13g2_decap_8 FILLER_45_828 ();
 sg13g2_decap_8 FILLER_45_835 ();
 sg13g2_decap_8 FILLER_45_842 ();
 sg13g2_decap_8 FILLER_45_849 ();
 sg13g2_decap_4 FILLER_45_856 ();
 sg13g2_fill_2 FILLER_45_860 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_4 FILLER_46_7 ();
 sg13g2_fill_2 FILLER_46_15 ();
 sg13g2_fill_1 FILLER_46_17 ();
 sg13g2_fill_2 FILLER_46_38 ();
 sg13g2_fill_1 FILLER_46_40 ();
 sg13g2_fill_1 FILLER_46_86 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_4 FILLER_46_112 ();
 sg13g2_fill_1 FILLER_46_116 ();
 sg13g2_fill_2 FILLER_46_161 ();
 sg13g2_decap_4 FILLER_46_176 ();
 sg13g2_fill_1 FILLER_46_197 ();
 sg13g2_decap_4 FILLER_46_228 ();
 sg13g2_fill_2 FILLER_46_232 ();
 sg13g2_fill_2 FILLER_46_265 ();
 sg13g2_decap_4 FILLER_46_290 ();
 sg13g2_fill_2 FILLER_46_342 ();
 sg13g2_fill_1 FILLER_46_349 ();
 sg13g2_decap_4 FILLER_46_385 ();
 sg13g2_fill_1 FILLER_46_389 ();
 sg13g2_decap_4 FILLER_46_421 ();
 sg13g2_fill_1 FILLER_46_436 ();
 sg13g2_fill_1 FILLER_46_466 ();
 sg13g2_fill_1 FILLER_46_474 ();
 sg13g2_fill_1 FILLER_46_523 ();
 sg13g2_fill_2 FILLER_46_541 ();
 sg13g2_fill_1 FILLER_46_543 ();
 sg13g2_fill_2 FILLER_46_565 ();
 sg13g2_fill_1 FILLER_46_579 ();
 sg13g2_decap_4 FILLER_46_584 ();
 sg13g2_fill_1 FILLER_46_588 ();
 sg13g2_fill_2 FILLER_46_619 ();
 sg13g2_fill_2 FILLER_46_656 ();
 sg13g2_fill_2 FILLER_46_723 ();
 sg13g2_fill_1 FILLER_46_733 ();
 sg13g2_fill_1 FILLER_46_738 ();
 sg13g2_decap_8 FILLER_46_775 ();
 sg13g2_decap_8 FILLER_46_782 ();
 sg13g2_decap_8 FILLER_46_789 ();
 sg13g2_decap_8 FILLER_46_796 ();
 sg13g2_decap_8 FILLER_46_803 ();
 sg13g2_decap_8 FILLER_46_810 ();
 sg13g2_decap_8 FILLER_46_817 ();
 sg13g2_decap_8 FILLER_46_824 ();
 sg13g2_decap_8 FILLER_46_831 ();
 sg13g2_decap_8 FILLER_46_838 ();
 sg13g2_decap_8 FILLER_46_845 ();
 sg13g2_decap_8 FILLER_46_852 ();
 sg13g2_fill_2 FILLER_46_859 ();
 sg13g2_fill_1 FILLER_46_861 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_decap_4 FILLER_47_83 ();
 sg13g2_fill_2 FILLER_47_87 ();
 sg13g2_decap_4 FILLER_47_115 ();
 sg13g2_fill_1 FILLER_47_119 ();
 sg13g2_fill_1 FILLER_47_125 ();
 sg13g2_decap_8 FILLER_47_135 ();
 sg13g2_decap_4 FILLER_47_142 ();
 sg13g2_decap_8 FILLER_47_150 ();
 sg13g2_decap_4 FILLER_47_157 ();
 sg13g2_fill_1 FILLER_47_177 ();
 sg13g2_decap_4 FILLER_47_187 ();
 sg13g2_fill_1 FILLER_47_191 ();
 sg13g2_decap_8 FILLER_47_263 ();
 sg13g2_fill_1 FILLER_47_277 ();
 sg13g2_fill_2 FILLER_47_304 ();
 sg13g2_fill_1 FILLER_47_324 ();
 sg13g2_fill_2 FILLER_47_351 ();
 sg13g2_fill_1 FILLER_47_353 ();
 sg13g2_decap_4 FILLER_47_384 ();
 sg13g2_fill_1 FILLER_47_388 ();
 sg13g2_fill_1 FILLER_47_397 ();
 sg13g2_fill_2 FILLER_47_411 ();
 sg13g2_fill_1 FILLER_47_608 ();
 sg13g2_fill_2 FILLER_47_627 ();
 sg13g2_fill_2 FILLER_47_643 ();
 sg13g2_decap_4 FILLER_47_710 ();
 sg13g2_fill_1 FILLER_47_759 ();
 sg13g2_decap_8 FILLER_47_778 ();
 sg13g2_decap_8 FILLER_47_785 ();
 sg13g2_decap_8 FILLER_47_792 ();
 sg13g2_decap_8 FILLER_47_799 ();
 sg13g2_decap_8 FILLER_47_806 ();
 sg13g2_decap_8 FILLER_47_813 ();
 sg13g2_decap_8 FILLER_47_820 ();
 sg13g2_decap_8 FILLER_47_827 ();
 sg13g2_decap_8 FILLER_47_834 ();
 sg13g2_decap_8 FILLER_47_841 ();
 sg13g2_decap_8 FILLER_47_848 ();
 sg13g2_decap_8 FILLER_47_855 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_4 FILLER_48_7 ();
 sg13g2_fill_1 FILLER_48_11 ();
 sg13g2_fill_2 FILLER_48_16 ();
 sg13g2_fill_2 FILLER_48_45 ();
 sg13g2_fill_1 FILLER_48_47 ();
 sg13g2_fill_1 FILLER_48_62 ();
 sg13g2_decap_4 FILLER_48_98 ();
 sg13g2_fill_1 FILLER_48_106 ();
 sg13g2_decap_4 FILLER_48_119 ();
 sg13g2_fill_2 FILLER_48_123 ();
 sg13g2_fill_1 FILLER_48_196 ();
 sg13g2_fill_2 FILLER_48_212 ();
 sg13g2_fill_1 FILLER_48_235 ();
 sg13g2_decap_4 FILLER_48_245 ();
 sg13g2_fill_2 FILLER_48_256 ();
 sg13g2_fill_1 FILLER_48_258 ();
 sg13g2_fill_2 FILLER_48_270 ();
 sg13g2_fill_1 FILLER_48_272 ();
 sg13g2_decap_4 FILLER_48_281 ();
 sg13g2_fill_2 FILLER_48_321 ();
 sg13g2_fill_1 FILLER_48_377 ();
 sg13g2_decap_4 FILLER_48_407 ();
 sg13g2_fill_2 FILLER_48_416 ();
 sg13g2_fill_2 FILLER_48_432 ();
 sg13g2_fill_1 FILLER_48_470 ();
 sg13g2_fill_2 FILLER_48_527 ();
 sg13g2_fill_2 FILLER_48_534 ();
 sg13g2_fill_2 FILLER_48_596 ();
 sg13g2_fill_1 FILLER_48_598 ();
 sg13g2_fill_2 FILLER_48_648 ();
 sg13g2_fill_1 FILLER_48_650 ();
 sg13g2_fill_1 FILLER_48_667 ();
 sg13g2_fill_2 FILLER_48_672 ();
 sg13g2_fill_1 FILLER_48_674 ();
 sg13g2_decap_8 FILLER_48_711 ();
 sg13g2_decap_4 FILLER_48_718 ();
 sg13g2_decap_8 FILLER_48_771 ();
 sg13g2_decap_8 FILLER_48_778 ();
 sg13g2_decap_8 FILLER_48_785 ();
 sg13g2_decap_8 FILLER_48_792 ();
 sg13g2_decap_8 FILLER_48_799 ();
 sg13g2_decap_8 FILLER_48_806 ();
 sg13g2_decap_8 FILLER_48_813 ();
 sg13g2_decap_8 FILLER_48_820 ();
 sg13g2_decap_8 FILLER_48_827 ();
 sg13g2_decap_8 FILLER_48_834 ();
 sg13g2_decap_8 FILLER_48_841 ();
 sg13g2_decap_8 FILLER_48_848 ();
 sg13g2_decap_8 FILLER_48_855 ();
 sg13g2_fill_2 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_58 ();
 sg13g2_fill_1 FILLER_49_80 ();
 sg13g2_fill_2 FILLER_49_95 ();
 sg13g2_fill_1 FILLER_49_97 ();
 sg13g2_fill_1 FILLER_49_123 ();
 sg13g2_fill_2 FILLER_49_134 ();
 sg13g2_fill_1 FILLER_49_136 ();
 sg13g2_fill_2 FILLER_49_155 ();
 sg13g2_fill_2 FILLER_49_179 ();
 sg13g2_fill_1 FILLER_49_181 ();
 sg13g2_decap_4 FILLER_49_242 ();
 sg13g2_fill_2 FILLER_49_246 ();
 sg13g2_decap_8 FILLER_49_279 ();
 sg13g2_fill_2 FILLER_49_286 ();
 sg13g2_fill_2 FILLER_49_310 ();
 sg13g2_fill_1 FILLER_49_386 ();
 sg13g2_fill_2 FILLER_49_425 ();
 sg13g2_fill_2 FILLER_49_436 ();
 sg13g2_fill_1 FILLER_49_463 ();
 sg13g2_fill_2 FILLER_49_473 ();
 sg13g2_fill_2 FILLER_49_502 ();
 sg13g2_fill_1 FILLER_49_504 ();
 sg13g2_decap_4 FILLER_49_640 ();
 sg13g2_fill_2 FILLER_49_657 ();
 sg13g2_fill_1 FILLER_49_659 ();
 sg13g2_fill_1 FILLER_49_683 ();
 sg13g2_fill_2 FILLER_49_693 ();
 sg13g2_fill_1 FILLER_49_735 ();
 sg13g2_decap_8 FILLER_49_768 ();
 sg13g2_decap_8 FILLER_49_775 ();
 sg13g2_decap_8 FILLER_49_782 ();
 sg13g2_decap_8 FILLER_49_789 ();
 sg13g2_decap_8 FILLER_49_796 ();
 sg13g2_decap_8 FILLER_49_803 ();
 sg13g2_decap_8 FILLER_49_810 ();
 sg13g2_decap_8 FILLER_49_817 ();
 sg13g2_decap_8 FILLER_49_824 ();
 sg13g2_decap_8 FILLER_49_831 ();
 sg13g2_decap_8 FILLER_49_838 ();
 sg13g2_decap_8 FILLER_49_845 ();
 sg13g2_decap_8 FILLER_49_852 ();
 sg13g2_fill_2 FILLER_49_859 ();
 sg13g2_fill_1 FILLER_49_861 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_29 ();
 sg13g2_fill_1 FILLER_50_31 ();
 sg13g2_fill_2 FILLER_50_46 ();
 sg13g2_fill_1 FILLER_50_66 ();
 sg13g2_fill_2 FILLER_50_81 ();
 sg13g2_fill_1 FILLER_50_83 ();
 sg13g2_fill_2 FILLER_50_125 ();
 sg13g2_fill_1 FILLER_50_148 ();
 sg13g2_fill_2 FILLER_50_196 ();
 sg13g2_decap_4 FILLER_50_202 ();
 sg13g2_fill_2 FILLER_50_206 ();
 sg13g2_decap_4 FILLER_50_220 ();
 sg13g2_fill_2 FILLER_50_224 ();
 sg13g2_fill_2 FILLER_50_235 ();
 sg13g2_fill_1 FILLER_50_237 ();
 sg13g2_decap_4 FILLER_50_251 ();
 sg13g2_fill_1 FILLER_50_255 ();
 sg13g2_decap_4 FILLER_50_288 ();
 sg13g2_fill_2 FILLER_50_292 ();
 sg13g2_fill_2 FILLER_50_340 ();
 sg13g2_decap_8 FILLER_50_351 ();
 sg13g2_fill_2 FILLER_50_367 ();
 sg13g2_fill_1 FILLER_50_378 ();
 sg13g2_fill_1 FILLER_50_406 ();
 sg13g2_fill_1 FILLER_50_422 ();
 sg13g2_fill_2 FILLER_50_454 ();
 sg13g2_fill_1 FILLER_50_602 ();
 sg13g2_fill_2 FILLER_50_705 ();
 sg13g2_decap_8 FILLER_50_773 ();
 sg13g2_decap_8 FILLER_50_780 ();
 sg13g2_decap_8 FILLER_50_787 ();
 sg13g2_decap_8 FILLER_50_794 ();
 sg13g2_decap_8 FILLER_50_801 ();
 sg13g2_decap_8 FILLER_50_808 ();
 sg13g2_decap_8 FILLER_50_815 ();
 sg13g2_decap_8 FILLER_50_822 ();
 sg13g2_decap_8 FILLER_50_829 ();
 sg13g2_decap_8 FILLER_50_836 ();
 sg13g2_decap_8 FILLER_50_843 ();
 sg13g2_decap_8 FILLER_50_850 ();
 sg13g2_decap_4 FILLER_50_857 ();
 sg13g2_fill_1 FILLER_50_861 ();
 sg13g2_decap_4 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_4 ();
 sg13g2_fill_2 FILLER_51_102 ();
 sg13g2_fill_1 FILLER_51_104 ();
 sg13g2_fill_2 FILLER_51_159 ();
 sg13g2_fill_2 FILLER_51_175 ();
 sg13g2_fill_2 FILLER_51_200 ();
 sg13g2_decap_4 FILLER_51_219 ();
 sg13g2_fill_1 FILLER_51_259 ();
 sg13g2_fill_1 FILLER_51_312 ();
 sg13g2_decap_4 FILLER_51_329 ();
 sg13g2_fill_1 FILLER_51_333 ();
 sg13g2_decap_4 FILLER_51_342 ();
 sg13g2_fill_1 FILLER_51_346 ();
 sg13g2_fill_2 FILLER_51_387 ();
 sg13g2_fill_2 FILLER_51_474 ();
 sg13g2_fill_1 FILLER_51_493 ();
 sg13g2_decap_4 FILLER_51_511 ();
 sg13g2_fill_1 FILLER_51_515 ();
 sg13g2_fill_1 FILLER_51_527 ();
 sg13g2_fill_2 FILLER_51_548 ();
 sg13g2_fill_1 FILLER_51_550 ();
 sg13g2_fill_1 FILLER_51_580 ();
 sg13g2_decap_4 FILLER_51_656 ();
 sg13g2_fill_2 FILLER_51_660 ();
 sg13g2_decap_8 FILLER_51_738 ();
 sg13g2_fill_2 FILLER_51_745 ();
 sg13g2_decap_8 FILLER_51_756 ();
 sg13g2_decap_8 FILLER_51_763 ();
 sg13g2_decap_8 FILLER_51_770 ();
 sg13g2_decap_8 FILLER_51_777 ();
 sg13g2_decap_8 FILLER_51_784 ();
 sg13g2_decap_8 FILLER_51_791 ();
 sg13g2_decap_8 FILLER_51_798 ();
 sg13g2_decap_8 FILLER_51_805 ();
 sg13g2_decap_8 FILLER_51_812 ();
 sg13g2_decap_8 FILLER_51_819 ();
 sg13g2_decap_8 FILLER_51_826 ();
 sg13g2_decap_8 FILLER_51_833 ();
 sg13g2_decap_8 FILLER_51_840 ();
 sg13g2_decap_8 FILLER_51_847 ();
 sg13g2_decap_8 FILLER_51_854 ();
 sg13g2_fill_1 FILLER_51_861 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_7 ();
 sg13g2_fill_2 FILLER_52_34 ();
 sg13g2_fill_1 FILLER_52_36 ();
 sg13g2_fill_1 FILLER_52_50 ();
 sg13g2_fill_2 FILLER_52_56 ();
 sg13g2_fill_1 FILLER_52_58 ();
 sg13g2_decap_4 FILLER_52_67 ();
 sg13g2_fill_2 FILLER_52_71 ();
 sg13g2_decap_8 FILLER_52_146 ();
 sg13g2_fill_1 FILLER_52_153 ();
 sg13g2_fill_1 FILLER_52_167 ();
 sg13g2_fill_2 FILLER_52_176 ();
 sg13g2_fill_1 FILLER_52_178 ();
 sg13g2_fill_1 FILLER_52_183 ();
 sg13g2_decap_4 FILLER_52_222 ();
 sg13g2_decap_4 FILLER_52_250 ();
 sg13g2_fill_1 FILLER_52_254 ();
 sg13g2_decap_4 FILLER_52_334 ();
 sg13g2_fill_1 FILLER_52_347 ();
 sg13g2_decap_8 FILLER_52_352 ();
 sg13g2_fill_2 FILLER_52_359 ();
 sg13g2_fill_1 FILLER_52_361 ();
 sg13g2_fill_2 FILLER_52_372 ();
 sg13g2_fill_2 FILLER_52_417 ();
 sg13g2_fill_2 FILLER_52_428 ();
 sg13g2_fill_1 FILLER_52_430 ();
 sg13g2_fill_2 FILLER_52_436 ();
 sg13g2_fill_1 FILLER_52_438 ();
 sg13g2_fill_1 FILLER_52_467 ();
 sg13g2_fill_1 FILLER_52_494 ();
 sg13g2_fill_1 FILLER_52_521 ();
 sg13g2_fill_1 FILLER_52_540 ();
 sg13g2_fill_2 FILLER_52_550 ();
 sg13g2_fill_1 FILLER_52_581 ();
 sg13g2_decap_8 FILLER_52_664 ();
 sg13g2_decap_4 FILLER_52_671 ();
 sg13g2_fill_2 FILLER_52_675 ();
 sg13g2_decap_4 FILLER_52_688 ();
 sg13g2_fill_1 FILLER_52_692 ();
 sg13g2_decap_8 FILLER_52_702 ();
 sg13g2_decap_8 FILLER_52_709 ();
 sg13g2_decap_8 FILLER_52_716 ();
 sg13g2_decap_8 FILLER_52_723 ();
 sg13g2_decap_8 FILLER_52_730 ();
 sg13g2_decap_8 FILLER_52_737 ();
 sg13g2_decap_8 FILLER_52_744 ();
 sg13g2_decap_8 FILLER_52_751 ();
 sg13g2_decap_8 FILLER_52_758 ();
 sg13g2_decap_8 FILLER_52_765 ();
 sg13g2_decap_8 FILLER_52_772 ();
 sg13g2_decap_8 FILLER_52_779 ();
 sg13g2_decap_8 FILLER_52_786 ();
 sg13g2_decap_8 FILLER_52_793 ();
 sg13g2_decap_8 FILLER_52_800 ();
 sg13g2_decap_8 FILLER_52_807 ();
 sg13g2_decap_8 FILLER_52_814 ();
 sg13g2_decap_8 FILLER_52_821 ();
 sg13g2_decap_8 FILLER_52_828 ();
 sg13g2_decap_8 FILLER_52_835 ();
 sg13g2_decap_8 FILLER_52_842 ();
 sg13g2_decap_8 FILLER_52_849 ();
 sg13g2_decap_4 FILLER_52_856 ();
 sg13g2_fill_2 FILLER_52_860 ();
 sg13g2_fill_1 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_32 ();
 sg13g2_fill_1 FILLER_53_58 ();
 sg13g2_decap_4 FILLER_53_67 ();
 sg13g2_fill_2 FILLER_53_79 ();
 sg13g2_fill_1 FILLER_53_89 ();
 sg13g2_fill_2 FILLER_53_98 ();
 sg13g2_fill_1 FILLER_53_100 ();
 sg13g2_fill_2 FILLER_53_110 ();
 sg13g2_fill_1 FILLER_53_112 ();
 sg13g2_fill_2 FILLER_53_121 ();
 sg13g2_decap_8 FILLER_53_140 ();
 sg13g2_fill_1 FILLER_53_147 ();
 sg13g2_fill_1 FILLER_53_160 ();
 sg13g2_fill_2 FILLER_53_167 ();
 sg13g2_fill_1 FILLER_53_169 ();
 sg13g2_fill_2 FILLER_53_187 ();
 sg13g2_fill_1 FILLER_53_189 ();
 sg13g2_fill_1 FILLER_53_207 ();
 sg13g2_fill_2 FILLER_53_212 ();
 sg13g2_decap_4 FILLER_53_220 ();
 sg13g2_decap_4 FILLER_53_228 ();
 sg13g2_fill_2 FILLER_53_232 ();
 sg13g2_fill_1 FILLER_53_239 ();
 sg13g2_decap_8 FILLER_53_255 ();
 sg13g2_decap_4 FILLER_53_262 ();
 sg13g2_fill_2 FILLER_53_266 ();
 sg13g2_fill_1 FILLER_53_276 ();
 sg13g2_fill_2 FILLER_53_312 ();
 sg13g2_fill_1 FILLER_53_329 ();
 sg13g2_fill_1 FILLER_53_334 ();
 sg13g2_fill_1 FILLER_53_387 ();
 sg13g2_fill_2 FILLER_53_402 ();
 sg13g2_fill_1 FILLER_53_431 ();
 sg13g2_decap_4 FILLER_53_456 ();
 sg13g2_fill_2 FILLER_53_460 ();
 sg13g2_fill_1 FILLER_53_496 ();
 sg13g2_decap_4 FILLER_53_523 ();
 sg13g2_decap_4 FILLER_53_531 ();
 sg13g2_fill_1 FILLER_53_535 ();
 sg13g2_fill_1 FILLER_53_566 ();
 sg13g2_fill_2 FILLER_53_611 ();
 sg13g2_fill_1 FILLER_53_613 ();
 sg13g2_decap_8 FILLER_53_627 ();
 sg13g2_decap_4 FILLER_53_634 ();
 sg13g2_fill_2 FILLER_53_638 ();
 sg13g2_decap_8 FILLER_53_653 ();
 sg13g2_decap_8 FILLER_53_660 ();
 sg13g2_decap_8 FILLER_53_667 ();
 sg13g2_decap_8 FILLER_53_674 ();
 sg13g2_decap_8 FILLER_53_681 ();
 sg13g2_decap_8 FILLER_53_688 ();
 sg13g2_decap_8 FILLER_53_695 ();
 sg13g2_decap_8 FILLER_53_702 ();
 sg13g2_decap_8 FILLER_53_709 ();
 sg13g2_decap_8 FILLER_53_716 ();
 sg13g2_decap_8 FILLER_53_723 ();
 sg13g2_decap_8 FILLER_53_730 ();
 sg13g2_decap_8 FILLER_53_737 ();
 sg13g2_decap_8 FILLER_53_744 ();
 sg13g2_decap_8 FILLER_53_751 ();
 sg13g2_decap_8 FILLER_53_758 ();
 sg13g2_decap_8 FILLER_53_765 ();
 sg13g2_decap_8 FILLER_53_772 ();
 sg13g2_decap_8 FILLER_53_779 ();
 sg13g2_decap_8 FILLER_53_786 ();
 sg13g2_decap_8 FILLER_53_793 ();
 sg13g2_decap_8 FILLER_53_800 ();
 sg13g2_decap_8 FILLER_53_807 ();
 sg13g2_decap_8 FILLER_53_814 ();
 sg13g2_decap_8 FILLER_53_821 ();
 sg13g2_decap_8 FILLER_53_828 ();
 sg13g2_decap_8 FILLER_53_835 ();
 sg13g2_decap_8 FILLER_53_842 ();
 sg13g2_decap_8 FILLER_53_849 ();
 sg13g2_decap_4 FILLER_53_856 ();
 sg13g2_fill_2 FILLER_53_860 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_decap_4 FILLER_54_60 ();
 sg13g2_fill_1 FILLER_54_64 ();
 sg13g2_fill_2 FILLER_54_73 ();
 sg13g2_fill_1 FILLER_54_75 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_fill_1 FILLER_54_119 ();
 sg13g2_decap_8 FILLER_54_124 ();
 sg13g2_fill_2 FILLER_54_137 ();
 sg13g2_decap_8 FILLER_54_164 ();
 sg13g2_decap_8 FILLER_54_176 ();
 sg13g2_decap_8 FILLER_54_183 ();
 sg13g2_fill_2 FILLER_54_190 ();
 sg13g2_decap_8 FILLER_54_200 ();
 sg13g2_fill_1 FILLER_54_215 ();
 sg13g2_fill_2 FILLER_54_224 ();
 sg13g2_decap_4 FILLER_54_265 ();
 sg13g2_fill_1 FILLER_54_269 ();
 sg13g2_fill_2 FILLER_54_278 ();
 sg13g2_fill_1 FILLER_54_280 ();
 sg13g2_fill_1 FILLER_54_285 ();
 sg13g2_decap_8 FILLER_54_312 ();
 sg13g2_fill_1 FILLER_54_371 ();
 sg13g2_fill_2 FILLER_54_390 ();
 sg13g2_fill_2 FILLER_54_410 ();
 sg13g2_fill_1 FILLER_54_417 ();
 sg13g2_fill_2 FILLER_54_441 ();
 sg13g2_decap_8 FILLER_54_448 ();
 sg13g2_decap_8 FILLER_54_455 ();
 sg13g2_fill_1 FILLER_54_462 ();
 sg13g2_decap_4 FILLER_54_486 ();
 sg13g2_fill_1 FILLER_54_490 ();
 sg13g2_fill_2 FILLER_54_505 ();
 sg13g2_decap_4 FILLER_54_545 ();
 sg13g2_fill_1 FILLER_54_549 ();
 sg13g2_fill_1 FILLER_54_561 ();
 sg13g2_decap_8 FILLER_54_565 ();
 sg13g2_fill_1 FILLER_54_572 ();
 sg13g2_fill_2 FILLER_54_591 ();
 sg13g2_fill_1 FILLER_54_597 ();
 sg13g2_decap_8 FILLER_54_624 ();
 sg13g2_decap_8 FILLER_54_631 ();
 sg13g2_decap_8 FILLER_54_638 ();
 sg13g2_decap_8 FILLER_54_645 ();
 sg13g2_decap_8 FILLER_54_652 ();
 sg13g2_decap_8 FILLER_54_659 ();
 sg13g2_decap_8 FILLER_54_666 ();
 sg13g2_decap_8 FILLER_54_673 ();
 sg13g2_decap_8 FILLER_54_680 ();
 sg13g2_decap_8 FILLER_54_687 ();
 sg13g2_decap_8 FILLER_54_694 ();
 sg13g2_decap_8 FILLER_54_701 ();
 sg13g2_decap_8 FILLER_54_708 ();
 sg13g2_decap_8 FILLER_54_715 ();
 sg13g2_decap_8 FILLER_54_722 ();
 sg13g2_decap_8 FILLER_54_729 ();
 sg13g2_decap_8 FILLER_54_736 ();
 sg13g2_decap_8 FILLER_54_743 ();
 sg13g2_decap_8 FILLER_54_750 ();
 sg13g2_decap_8 FILLER_54_757 ();
 sg13g2_decap_8 FILLER_54_764 ();
 sg13g2_decap_8 FILLER_54_771 ();
 sg13g2_decap_8 FILLER_54_778 ();
 sg13g2_decap_8 FILLER_54_785 ();
 sg13g2_decap_8 FILLER_54_792 ();
 sg13g2_decap_8 FILLER_54_799 ();
 sg13g2_decap_8 FILLER_54_806 ();
 sg13g2_decap_8 FILLER_54_813 ();
 sg13g2_decap_8 FILLER_54_820 ();
 sg13g2_decap_8 FILLER_54_827 ();
 sg13g2_decap_8 FILLER_54_834 ();
 sg13g2_decap_8 FILLER_54_841 ();
 sg13g2_decap_8 FILLER_54_848 ();
 sg13g2_decap_8 FILLER_54_855 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_7 ();
 sg13g2_fill_2 FILLER_55_40 ();
 sg13g2_fill_2 FILLER_55_50 ();
 sg13g2_fill_1 FILLER_55_52 ();
 sg13g2_fill_1 FILLER_55_65 ();
 sg13g2_fill_2 FILLER_55_81 ();
 sg13g2_fill_1 FILLER_55_95 ();
 sg13g2_decap_8 FILLER_55_104 ();
 sg13g2_fill_2 FILLER_55_111 ();
 sg13g2_fill_2 FILLER_55_119 ();
 sg13g2_fill_1 FILLER_55_121 ();
 sg13g2_decap_8 FILLER_55_130 ();
 sg13g2_decap_4 FILLER_55_137 ();
 sg13g2_fill_2 FILLER_55_141 ();
 sg13g2_decap_8 FILLER_55_159 ();
 sg13g2_fill_1 FILLER_55_196 ();
 sg13g2_decap_4 FILLER_55_209 ();
 sg13g2_fill_1 FILLER_55_213 ();
 sg13g2_fill_2 FILLER_55_237 ();
 sg13g2_fill_1 FILLER_55_244 ();
 sg13g2_fill_1 FILLER_55_275 ();
 sg13g2_decap_8 FILLER_55_284 ();
 sg13g2_decap_4 FILLER_55_291 ();
 sg13g2_fill_2 FILLER_55_332 ();
 sg13g2_fill_1 FILLER_55_348 ();
 sg13g2_fill_2 FILLER_55_369 ();
 sg13g2_fill_2 FILLER_55_401 ();
 sg13g2_fill_2 FILLER_55_438 ();
 sg13g2_fill_1 FILLER_55_440 ();
 sg13g2_decap_4 FILLER_55_462 ();
 sg13g2_fill_1 FILLER_55_490 ();
 sg13g2_decap_4 FILLER_55_509 ();
 sg13g2_fill_1 FILLER_55_529 ();
 sg13g2_fill_1 FILLER_55_559 ();
 sg13g2_decap_8 FILLER_55_604 ();
 sg13g2_fill_2 FILLER_55_611 ();
 sg13g2_fill_1 FILLER_55_613 ();
 sg13g2_decap_4 FILLER_55_617 ();
 sg13g2_fill_1 FILLER_55_621 ();
 sg13g2_decap_8 FILLER_55_626 ();
 sg13g2_fill_1 FILLER_55_633 ();
 sg13g2_decap_8 FILLER_55_641 ();
 sg13g2_decap_8 FILLER_55_648 ();
 sg13g2_decap_8 FILLER_55_655 ();
 sg13g2_decap_8 FILLER_55_662 ();
 sg13g2_decap_8 FILLER_55_669 ();
 sg13g2_decap_8 FILLER_55_676 ();
 sg13g2_decap_8 FILLER_55_683 ();
 sg13g2_decap_8 FILLER_55_690 ();
 sg13g2_decap_8 FILLER_55_697 ();
 sg13g2_decap_8 FILLER_55_704 ();
 sg13g2_decap_8 FILLER_55_711 ();
 sg13g2_decap_8 FILLER_55_718 ();
 sg13g2_decap_8 FILLER_55_725 ();
 sg13g2_decap_8 FILLER_55_732 ();
 sg13g2_decap_8 FILLER_55_739 ();
 sg13g2_decap_8 FILLER_55_746 ();
 sg13g2_decap_8 FILLER_55_753 ();
 sg13g2_decap_8 FILLER_55_760 ();
 sg13g2_decap_8 FILLER_55_767 ();
 sg13g2_decap_8 FILLER_55_774 ();
 sg13g2_decap_8 FILLER_55_781 ();
 sg13g2_decap_8 FILLER_55_788 ();
 sg13g2_decap_8 FILLER_55_795 ();
 sg13g2_decap_8 FILLER_55_802 ();
 sg13g2_decap_8 FILLER_55_809 ();
 sg13g2_decap_8 FILLER_55_816 ();
 sg13g2_decap_8 FILLER_55_823 ();
 sg13g2_decap_8 FILLER_55_830 ();
 sg13g2_decap_8 FILLER_55_837 ();
 sg13g2_decap_8 FILLER_55_844 ();
 sg13g2_decap_8 FILLER_55_851 ();
 sg13g2_decap_4 FILLER_55_858 ();
 sg13g2_fill_2 FILLER_56_26 ();
 sg13g2_fill_1 FILLER_56_28 ();
 sg13g2_decap_4 FILLER_56_79 ();
 sg13g2_decap_4 FILLER_56_129 ();
 sg13g2_decap_8 FILLER_56_174 ();
 sg13g2_fill_2 FILLER_56_181 ();
 sg13g2_fill_1 FILLER_56_189 ();
 sg13g2_decap_8 FILLER_56_199 ();
 sg13g2_decap_4 FILLER_56_206 ();
 sg13g2_fill_2 FILLER_56_227 ();
 sg13g2_fill_2 FILLER_56_308 ();
 sg13g2_decap_4 FILLER_56_410 ();
 sg13g2_fill_1 FILLER_56_414 ();
 sg13g2_decap_8 FILLER_56_424 ();
 sg13g2_fill_2 FILLER_56_431 ();
 sg13g2_fill_1 FILLER_56_433 ();
 sg13g2_decap_4 FILLER_56_440 ();
 sg13g2_fill_2 FILLER_56_457 ();
 sg13g2_fill_2 FILLER_56_464 ();
 sg13g2_fill_1 FILLER_56_466 ();
 sg13g2_fill_1 FILLER_56_477 ();
 sg13g2_fill_1 FILLER_56_490 ();
 sg13g2_decap_4 FILLER_56_500 ();
 sg13g2_fill_1 FILLER_56_504 ();
 sg13g2_decap_4 FILLER_56_546 ();
 sg13g2_fill_2 FILLER_56_550 ();
 sg13g2_fill_2 FILLER_56_562 ();
 sg13g2_fill_1 FILLER_56_564 ();
 sg13g2_fill_1 FILLER_56_585 ();
 sg13g2_fill_1 FILLER_56_590 ();
 sg13g2_decap_8 FILLER_56_663 ();
 sg13g2_decap_8 FILLER_56_670 ();
 sg13g2_decap_8 FILLER_56_677 ();
 sg13g2_decap_8 FILLER_56_684 ();
 sg13g2_decap_8 FILLER_56_691 ();
 sg13g2_decap_8 FILLER_56_698 ();
 sg13g2_decap_8 FILLER_56_705 ();
 sg13g2_decap_8 FILLER_56_712 ();
 sg13g2_decap_8 FILLER_56_719 ();
 sg13g2_decap_8 FILLER_56_726 ();
 sg13g2_decap_8 FILLER_56_733 ();
 sg13g2_decap_8 FILLER_56_740 ();
 sg13g2_decap_8 FILLER_56_747 ();
 sg13g2_decap_8 FILLER_56_754 ();
 sg13g2_decap_8 FILLER_56_761 ();
 sg13g2_decap_8 FILLER_56_768 ();
 sg13g2_decap_8 FILLER_56_775 ();
 sg13g2_decap_8 FILLER_56_782 ();
 sg13g2_decap_8 FILLER_56_789 ();
 sg13g2_decap_8 FILLER_56_796 ();
 sg13g2_decap_8 FILLER_56_803 ();
 sg13g2_decap_8 FILLER_56_810 ();
 sg13g2_decap_8 FILLER_56_817 ();
 sg13g2_decap_8 FILLER_56_824 ();
 sg13g2_decap_8 FILLER_56_831 ();
 sg13g2_decap_8 FILLER_56_838 ();
 sg13g2_decap_8 FILLER_56_845 ();
 sg13g2_decap_8 FILLER_56_852 ();
 sg13g2_fill_2 FILLER_56_859 ();
 sg13g2_fill_1 FILLER_56_861 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_20 ();
 sg13g2_fill_1 FILLER_57_22 ();
 sg13g2_fill_1 FILLER_57_42 ();
 sg13g2_fill_2 FILLER_57_55 ();
 sg13g2_fill_1 FILLER_57_57 ();
 sg13g2_decap_4 FILLER_57_67 ();
 sg13g2_fill_2 FILLER_57_86 ();
 sg13g2_fill_1 FILLER_57_97 ();
 sg13g2_fill_2 FILLER_57_115 ();
 sg13g2_fill_1 FILLER_57_117 ();
 sg13g2_fill_1 FILLER_57_123 ();
 sg13g2_decap_8 FILLER_57_129 ();
 sg13g2_decap_4 FILLER_57_136 ();
 sg13g2_fill_1 FILLER_57_140 ();
 sg13g2_decap_4 FILLER_57_152 ();
 sg13g2_fill_2 FILLER_57_156 ();
 sg13g2_fill_1 FILLER_57_173 ();
 sg13g2_decap_8 FILLER_57_198 ();
 sg13g2_fill_1 FILLER_57_205 ();
 sg13g2_fill_2 FILLER_57_214 ();
 sg13g2_fill_1 FILLER_57_239 ();
 sg13g2_fill_1 FILLER_57_289 ();
 sg13g2_fill_2 FILLER_57_316 ();
 sg13g2_fill_1 FILLER_57_318 ();
 sg13g2_fill_1 FILLER_57_345 ();
 sg13g2_fill_1 FILLER_57_371 ();
 sg13g2_fill_1 FILLER_57_398 ();
 sg13g2_fill_1 FILLER_57_433 ();
 sg13g2_decap_8 FILLER_57_452 ();
 sg13g2_decap_4 FILLER_57_464 ();
 sg13g2_fill_1 FILLER_57_476 ();
 sg13g2_fill_2 FILLER_57_487 ();
 sg13g2_decap_8 FILLER_57_547 ();
 sg13g2_fill_2 FILLER_57_554 ();
 sg13g2_decap_8 FILLER_57_571 ();
 sg13g2_decap_4 FILLER_57_578 ();
 sg13g2_fill_2 FILLER_57_585 ();
 sg13g2_decap_4 FILLER_57_606 ();
 sg13g2_fill_2 FILLER_57_610 ();
 sg13g2_fill_1 FILLER_57_645 ();
 sg13g2_decap_8 FILLER_57_663 ();
 sg13g2_decap_8 FILLER_57_670 ();
 sg13g2_decap_8 FILLER_57_677 ();
 sg13g2_decap_8 FILLER_57_684 ();
 sg13g2_decap_8 FILLER_57_691 ();
 sg13g2_decap_8 FILLER_57_698 ();
 sg13g2_decap_8 FILLER_57_705 ();
 sg13g2_decap_8 FILLER_57_712 ();
 sg13g2_decap_8 FILLER_57_719 ();
 sg13g2_decap_8 FILLER_57_726 ();
 sg13g2_decap_8 FILLER_57_733 ();
 sg13g2_decap_8 FILLER_57_740 ();
 sg13g2_decap_8 FILLER_57_747 ();
 sg13g2_decap_8 FILLER_57_754 ();
 sg13g2_decap_8 FILLER_57_761 ();
 sg13g2_decap_8 FILLER_57_768 ();
 sg13g2_decap_8 FILLER_57_775 ();
 sg13g2_decap_8 FILLER_57_782 ();
 sg13g2_decap_8 FILLER_57_789 ();
 sg13g2_decap_8 FILLER_57_796 ();
 sg13g2_decap_8 FILLER_57_803 ();
 sg13g2_decap_8 FILLER_57_810 ();
 sg13g2_decap_8 FILLER_57_817 ();
 sg13g2_decap_8 FILLER_57_824 ();
 sg13g2_decap_8 FILLER_57_831 ();
 sg13g2_decap_8 FILLER_57_838 ();
 sg13g2_decap_8 FILLER_57_845 ();
 sg13g2_decap_8 FILLER_57_852 ();
 sg13g2_fill_2 FILLER_57_859 ();
 sg13g2_fill_1 FILLER_57_861 ();
 sg13g2_decap_4 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_4 ();
 sg13g2_decap_4 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_138 ();
 sg13g2_decap_4 FILLER_58_145 ();
 sg13g2_decap_8 FILLER_58_170 ();
 sg13g2_decap_4 FILLER_58_177 ();
 sg13g2_fill_1 FILLER_58_181 ();
 sg13g2_decap_4 FILLER_58_191 ();
 sg13g2_fill_2 FILLER_58_195 ();
 sg13g2_fill_2 FILLER_58_205 ();
 sg13g2_fill_1 FILLER_58_207 ();
 sg13g2_fill_2 FILLER_58_222 ();
 sg13g2_fill_1 FILLER_58_269 ();
 sg13g2_fill_2 FILLER_58_275 ();
 sg13g2_fill_1 FILLER_58_290 ();
 sg13g2_fill_1 FILLER_58_297 ();
 sg13g2_fill_1 FILLER_58_363 ();
 sg13g2_decap_4 FILLER_58_413 ();
 sg13g2_decap_4 FILLER_58_431 ();
 sg13g2_fill_2 FILLER_58_435 ();
 sg13g2_fill_2 FILLER_58_440 ();
 sg13g2_decap_8 FILLER_58_446 ();
 sg13g2_fill_2 FILLER_58_489 ();
 sg13g2_fill_1 FILLER_58_496 ();
 sg13g2_fill_1 FILLER_58_536 ();
 sg13g2_fill_2 FILLER_58_542 ();
 sg13g2_fill_1 FILLER_58_544 ();
 sg13g2_fill_2 FILLER_58_552 ();
 sg13g2_fill_1 FILLER_58_572 ();
 sg13g2_decap_4 FILLER_58_599 ();
 sg13g2_fill_2 FILLER_58_603 ();
 sg13g2_fill_1 FILLER_58_620 ();
 sg13g2_decap_8 FILLER_58_664 ();
 sg13g2_decap_8 FILLER_58_671 ();
 sg13g2_decap_8 FILLER_58_678 ();
 sg13g2_decap_8 FILLER_58_685 ();
 sg13g2_decap_8 FILLER_58_692 ();
 sg13g2_decap_8 FILLER_58_699 ();
 sg13g2_decap_8 FILLER_58_706 ();
 sg13g2_decap_8 FILLER_58_713 ();
 sg13g2_decap_8 FILLER_58_720 ();
 sg13g2_decap_8 FILLER_58_727 ();
 sg13g2_decap_8 FILLER_58_734 ();
 sg13g2_decap_8 FILLER_58_741 ();
 sg13g2_decap_8 FILLER_58_748 ();
 sg13g2_decap_8 FILLER_58_755 ();
 sg13g2_decap_8 FILLER_58_762 ();
 sg13g2_decap_8 FILLER_58_769 ();
 sg13g2_decap_8 FILLER_58_776 ();
 sg13g2_decap_8 FILLER_58_783 ();
 sg13g2_decap_8 FILLER_58_790 ();
 sg13g2_decap_8 FILLER_58_797 ();
 sg13g2_decap_8 FILLER_58_804 ();
 sg13g2_decap_8 FILLER_58_811 ();
 sg13g2_decap_8 FILLER_58_818 ();
 sg13g2_decap_8 FILLER_58_825 ();
 sg13g2_decap_8 FILLER_58_832 ();
 sg13g2_decap_8 FILLER_58_839 ();
 sg13g2_decap_8 FILLER_58_846 ();
 sg13g2_decap_8 FILLER_58_853 ();
 sg13g2_fill_2 FILLER_58_860 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_fill_2 FILLER_59_14 ();
 sg13g2_fill_1 FILLER_59_25 ();
 sg13g2_decap_4 FILLER_59_44 ();
 sg13g2_fill_2 FILLER_59_48 ();
 sg13g2_fill_2 FILLER_59_55 ();
 sg13g2_fill_1 FILLER_59_61 ();
 sg13g2_fill_1 FILLER_59_67 ();
 sg13g2_fill_1 FILLER_59_86 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_102 ();
 sg13g2_fill_2 FILLER_59_109 ();
 sg13g2_fill_1 FILLER_59_111 ();
 sg13g2_decap_4 FILLER_59_126 ();
 sg13g2_fill_2 FILLER_59_135 ();
 sg13g2_fill_1 FILLER_59_137 ();
 sg13g2_decap_8 FILLER_59_173 ();
 sg13g2_decap_4 FILLER_59_180 ();
 sg13g2_fill_1 FILLER_59_184 ();
 sg13g2_fill_1 FILLER_59_190 ();
 sg13g2_fill_2 FILLER_59_219 ();
 sg13g2_fill_1 FILLER_59_221 ();
 sg13g2_fill_2 FILLER_59_278 ();
 sg13g2_fill_2 FILLER_59_288 ();
 sg13g2_fill_1 FILLER_59_290 ();
 sg13g2_fill_2 FILLER_59_297 ();
 sg13g2_fill_1 FILLER_59_299 ();
 sg13g2_fill_2 FILLER_59_357 ();
 sg13g2_fill_1 FILLER_59_374 ();
 sg13g2_fill_2 FILLER_59_396 ();
 sg13g2_fill_1 FILLER_59_398 ();
 sg13g2_fill_2 FILLER_59_451 ();
 sg13g2_fill_1 FILLER_59_453 ();
 sg13g2_decap_8 FILLER_59_489 ();
 sg13g2_fill_1 FILLER_59_496 ();
 sg13g2_fill_2 FILLER_59_501 ();
 sg13g2_decap_4 FILLER_59_513 ();
 sg13g2_fill_2 FILLER_59_526 ();
 sg13g2_decap_4 FILLER_59_563 ();
 sg13g2_fill_2 FILLER_59_567 ();
 sg13g2_fill_2 FILLER_59_591 ();
 sg13g2_fill_1 FILLER_59_593 ();
 sg13g2_decap_8 FILLER_59_666 ();
 sg13g2_decap_8 FILLER_59_673 ();
 sg13g2_decap_8 FILLER_59_680 ();
 sg13g2_decap_8 FILLER_59_687 ();
 sg13g2_decap_8 FILLER_59_694 ();
 sg13g2_decap_8 FILLER_59_701 ();
 sg13g2_decap_8 FILLER_59_708 ();
 sg13g2_decap_8 FILLER_59_715 ();
 sg13g2_decap_8 FILLER_59_722 ();
 sg13g2_decap_8 FILLER_59_729 ();
 sg13g2_decap_8 FILLER_59_736 ();
 sg13g2_decap_8 FILLER_59_743 ();
 sg13g2_decap_8 FILLER_59_750 ();
 sg13g2_decap_8 FILLER_59_757 ();
 sg13g2_decap_8 FILLER_59_764 ();
 sg13g2_decap_8 FILLER_59_771 ();
 sg13g2_decap_8 FILLER_59_778 ();
 sg13g2_decap_8 FILLER_59_785 ();
 sg13g2_decap_8 FILLER_59_792 ();
 sg13g2_decap_8 FILLER_59_799 ();
 sg13g2_decap_8 FILLER_59_806 ();
 sg13g2_decap_8 FILLER_59_813 ();
 sg13g2_decap_8 FILLER_59_820 ();
 sg13g2_decap_8 FILLER_59_827 ();
 sg13g2_decap_8 FILLER_59_834 ();
 sg13g2_decap_8 FILLER_59_841 ();
 sg13g2_decap_8 FILLER_59_848 ();
 sg13g2_decap_8 FILLER_59_855 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_fill_1 FILLER_60_64 ();
 sg13g2_fill_2 FILLER_60_73 ();
 sg13g2_fill_1 FILLER_60_75 ();
 sg13g2_fill_2 FILLER_60_85 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_decap_4 FILLER_60_105 ();
 sg13g2_fill_2 FILLER_60_121 ();
 sg13g2_decap_4 FILLER_60_134 ();
 sg13g2_decap_4 FILLER_60_161 ();
 sg13g2_fill_2 FILLER_60_165 ();
 sg13g2_fill_2 FILLER_60_213 ();
 sg13g2_fill_2 FILLER_60_298 ();
 sg13g2_fill_1 FILLER_60_300 ();
 sg13g2_fill_2 FILLER_60_305 ();
 sg13g2_fill_1 FILLER_60_307 ();
 sg13g2_fill_1 FILLER_60_341 ();
 sg13g2_fill_2 FILLER_60_357 ();
 sg13g2_fill_2 FILLER_60_385 ();
 sg13g2_fill_1 FILLER_60_387 ();
 sg13g2_decap_8 FILLER_60_434 ();
 sg13g2_fill_2 FILLER_60_441 ();
 sg13g2_fill_1 FILLER_60_443 ();
 sg13g2_fill_2 FILLER_60_454 ();
 sg13g2_fill_1 FILLER_60_456 ();
 sg13g2_fill_2 FILLER_60_462 ();
 sg13g2_fill_2 FILLER_60_588 ();
 sg13g2_fill_1 FILLER_60_590 ();
 sg13g2_fill_1 FILLER_60_596 ();
 sg13g2_fill_2 FILLER_60_639 ();
 sg13g2_fill_1 FILLER_60_641 ();
 sg13g2_decap_8 FILLER_60_669 ();
 sg13g2_decap_8 FILLER_60_676 ();
 sg13g2_decap_8 FILLER_60_683 ();
 sg13g2_decap_8 FILLER_60_690 ();
 sg13g2_decap_8 FILLER_60_697 ();
 sg13g2_decap_8 FILLER_60_704 ();
 sg13g2_decap_8 FILLER_60_711 ();
 sg13g2_decap_8 FILLER_60_718 ();
 sg13g2_decap_8 FILLER_60_725 ();
 sg13g2_decap_8 FILLER_60_732 ();
 sg13g2_decap_8 FILLER_60_739 ();
 sg13g2_decap_8 FILLER_60_746 ();
 sg13g2_decap_8 FILLER_60_753 ();
 sg13g2_decap_8 FILLER_60_760 ();
 sg13g2_decap_8 FILLER_60_767 ();
 sg13g2_decap_8 FILLER_60_774 ();
 sg13g2_decap_8 FILLER_60_781 ();
 sg13g2_decap_8 FILLER_60_788 ();
 sg13g2_decap_8 FILLER_60_795 ();
 sg13g2_decap_8 FILLER_60_802 ();
 sg13g2_decap_8 FILLER_60_809 ();
 sg13g2_decap_8 FILLER_60_816 ();
 sg13g2_decap_8 FILLER_60_823 ();
 sg13g2_decap_8 FILLER_60_830 ();
 sg13g2_decap_8 FILLER_60_837 ();
 sg13g2_decap_8 FILLER_60_844 ();
 sg13g2_decap_8 FILLER_60_851 ();
 sg13g2_decap_4 FILLER_60_858 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_4 FILLER_61_7 ();
 sg13g2_fill_2 FILLER_61_11 ();
 sg13g2_fill_2 FILLER_61_39 ();
 sg13g2_fill_1 FILLER_61_59 ();
 sg13g2_fill_2 FILLER_61_65 ();
 sg13g2_fill_1 FILLER_61_67 ();
 sg13g2_decap_4 FILLER_61_171 ();
 sg13g2_fill_1 FILLER_61_175 ();
 sg13g2_fill_2 FILLER_61_211 ();
 sg13g2_fill_1 FILLER_61_213 ();
 sg13g2_fill_2 FILLER_61_264 ();
 sg13g2_fill_1 FILLER_61_266 ();
 sg13g2_fill_2 FILLER_61_280 ();
 sg13g2_fill_1 FILLER_61_282 ();
 sg13g2_decap_4 FILLER_61_287 ();
 sg13g2_fill_1 FILLER_61_317 ();
 sg13g2_decap_4 FILLER_61_328 ();
 sg13g2_decap_4 FILLER_61_346 ();
 sg13g2_fill_2 FILLER_61_376 ();
 sg13g2_decap_4 FILLER_61_408 ();
 sg13g2_fill_2 FILLER_61_432 ();
 sg13g2_fill_1 FILLER_61_434 ();
 sg13g2_fill_2 FILLER_61_445 ();
 sg13g2_fill_1 FILLER_61_447 ();
 sg13g2_fill_2 FILLER_61_468 ();
 sg13g2_decap_8 FILLER_61_485 ();
 sg13g2_decap_4 FILLER_61_492 ();
 sg13g2_fill_2 FILLER_61_496 ();
 sg13g2_fill_2 FILLER_61_528 ();
 sg13g2_fill_1 FILLER_61_536 ();
 sg13g2_fill_1 FILLER_61_625 ();
 sg13g2_decap_8 FILLER_61_666 ();
 sg13g2_decap_8 FILLER_61_673 ();
 sg13g2_decap_8 FILLER_61_680 ();
 sg13g2_decap_8 FILLER_61_687 ();
 sg13g2_decap_8 FILLER_61_694 ();
 sg13g2_decap_8 FILLER_61_701 ();
 sg13g2_decap_8 FILLER_61_708 ();
 sg13g2_decap_8 FILLER_61_715 ();
 sg13g2_decap_8 FILLER_61_722 ();
 sg13g2_decap_8 FILLER_61_729 ();
 sg13g2_decap_8 FILLER_61_736 ();
 sg13g2_decap_8 FILLER_61_743 ();
 sg13g2_decap_8 FILLER_61_750 ();
 sg13g2_decap_8 FILLER_61_757 ();
 sg13g2_decap_8 FILLER_61_764 ();
 sg13g2_decap_8 FILLER_61_771 ();
 sg13g2_decap_8 FILLER_61_778 ();
 sg13g2_decap_8 FILLER_61_785 ();
 sg13g2_decap_8 FILLER_61_792 ();
 sg13g2_decap_8 FILLER_61_799 ();
 sg13g2_decap_8 FILLER_61_806 ();
 sg13g2_decap_8 FILLER_61_813 ();
 sg13g2_decap_8 FILLER_61_820 ();
 sg13g2_decap_8 FILLER_61_827 ();
 sg13g2_decap_8 FILLER_61_834 ();
 sg13g2_decap_8 FILLER_61_841 ();
 sg13g2_decap_8 FILLER_61_848 ();
 sg13g2_decap_8 FILLER_61_855 ();
 sg13g2_fill_1 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_55 ();
 sg13g2_fill_1 FILLER_62_66 ();
 sg13g2_fill_2 FILLER_62_81 ();
 sg13g2_fill_1 FILLER_62_83 ();
 sg13g2_fill_2 FILLER_62_104 ();
 sg13g2_fill_1 FILLER_62_116 ();
 sg13g2_fill_1 FILLER_62_123 ();
 sg13g2_fill_1 FILLER_62_168 ();
 sg13g2_fill_2 FILLER_62_226 ();
 sg13g2_fill_1 FILLER_62_228 ();
 sg13g2_fill_1 FILLER_62_249 ();
 sg13g2_fill_2 FILLER_62_258 ();
 sg13g2_fill_1 FILLER_62_260 ();
 sg13g2_fill_2 FILLER_62_299 ();
 sg13g2_fill_1 FILLER_62_301 ();
 sg13g2_fill_1 FILLER_62_306 ();
 sg13g2_fill_2 FILLER_62_325 ();
 sg13g2_fill_1 FILLER_62_327 ();
 sg13g2_decap_8 FILLER_62_372 ();
 sg13g2_decap_8 FILLER_62_397 ();
 sg13g2_fill_1 FILLER_62_404 ();
 sg13g2_fill_2 FILLER_62_438 ();
 sg13g2_fill_2 FILLER_62_464 ();
 sg13g2_fill_2 FILLER_62_476 ();
 sg13g2_fill_1 FILLER_62_478 ();
 sg13g2_fill_1 FILLER_62_483 ();
 sg13g2_fill_2 FILLER_62_493 ();
 sg13g2_fill_1 FILLER_62_495 ();
 sg13g2_fill_2 FILLER_62_499 ();
 sg13g2_fill_2 FILLER_62_519 ();
 sg13g2_fill_2 FILLER_62_600 ();
 sg13g2_fill_1 FILLER_62_650 ();
 sg13g2_fill_1 FILLER_62_663 ();
 sg13g2_decap_8 FILLER_62_676 ();
 sg13g2_decap_8 FILLER_62_683 ();
 sg13g2_decap_8 FILLER_62_690 ();
 sg13g2_decap_8 FILLER_62_697 ();
 sg13g2_decap_8 FILLER_62_704 ();
 sg13g2_decap_8 FILLER_62_711 ();
 sg13g2_decap_8 FILLER_62_718 ();
 sg13g2_decap_8 FILLER_62_725 ();
 sg13g2_decap_8 FILLER_62_732 ();
 sg13g2_decap_8 FILLER_62_739 ();
 sg13g2_decap_8 FILLER_62_746 ();
 sg13g2_decap_8 FILLER_62_753 ();
 sg13g2_decap_8 FILLER_62_760 ();
 sg13g2_decap_8 FILLER_62_767 ();
 sg13g2_decap_8 FILLER_62_774 ();
 sg13g2_decap_8 FILLER_62_781 ();
 sg13g2_decap_8 FILLER_62_788 ();
 sg13g2_decap_8 FILLER_62_795 ();
 sg13g2_decap_8 FILLER_62_802 ();
 sg13g2_decap_8 FILLER_62_809 ();
 sg13g2_decap_8 FILLER_62_816 ();
 sg13g2_decap_8 FILLER_62_823 ();
 sg13g2_decap_8 FILLER_62_830 ();
 sg13g2_decap_8 FILLER_62_837 ();
 sg13g2_decap_8 FILLER_62_844 ();
 sg13g2_decap_8 FILLER_62_851 ();
 sg13g2_decap_4 FILLER_62_858 ();
 sg13g2_fill_1 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_36 ();
 sg13g2_fill_1 FILLER_63_62 ();
 sg13g2_fill_2 FILLER_63_89 ();
 sg13g2_fill_1 FILLER_63_91 ();
 sg13g2_fill_2 FILLER_63_183 ();
 sg13g2_decap_8 FILLER_63_252 ();
 sg13g2_decap_4 FILLER_63_259 ();
 sg13g2_decap_4 FILLER_63_281 ();
 sg13g2_fill_1 FILLER_63_325 ();
 sg13g2_fill_1 FILLER_63_348 ();
 sg13g2_decap_4 FILLER_63_407 ();
 sg13g2_fill_1 FILLER_63_411 ();
 sg13g2_decap_4 FILLER_63_431 ();
 sg13g2_fill_1 FILLER_63_435 ();
 sg13g2_fill_2 FILLER_63_466 ();
 sg13g2_fill_1 FILLER_63_529 ();
 sg13g2_decap_8 FILLER_63_581 ();
 sg13g2_fill_2 FILLER_63_588 ();
 sg13g2_fill_2 FILLER_63_607 ();
 sg13g2_decap_8 FILLER_63_694 ();
 sg13g2_decap_8 FILLER_63_701 ();
 sg13g2_decap_8 FILLER_63_708 ();
 sg13g2_decap_8 FILLER_63_715 ();
 sg13g2_decap_8 FILLER_63_722 ();
 sg13g2_decap_8 FILLER_63_729 ();
 sg13g2_decap_8 FILLER_63_736 ();
 sg13g2_decap_8 FILLER_63_743 ();
 sg13g2_decap_8 FILLER_63_750 ();
 sg13g2_decap_8 FILLER_63_757 ();
 sg13g2_decap_8 FILLER_63_764 ();
 sg13g2_decap_8 FILLER_63_771 ();
 sg13g2_decap_8 FILLER_63_778 ();
 sg13g2_decap_8 FILLER_63_785 ();
 sg13g2_decap_8 FILLER_63_792 ();
 sg13g2_decap_8 FILLER_63_799 ();
 sg13g2_decap_8 FILLER_63_806 ();
 sg13g2_decap_8 FILLER_63_813 ();
 sg13g2_decap_8 FILLER_63_820 ();
 sg13g2_decap_8 FILLER_63_827 ();
 sg13g2_decap_8 FILLER_63_834 ();
 sg13g2_decap_8 FILLER_63_841 ();
 sg13g2_decap_8 FILLER_63_848 ();
 sg13g2_decap_8 FILLER_63_855 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_7 ();
 sg13g2_fill_1 FILLER_64_9 ();
 sg13g2_fill_1 FILLER_64_73 ();
 sg13g2_fill_2 FILLER_64_78 ();
 sg13g2_fill_1 FILLER_64_80 ();
 sg13g2_fill_1 FILLER_64_110 ();
 sg13g2_fill_2 FILLER_64_128 ();
 sg13g2_fill_2 FILLER_64_155 ();
 sg13g2_fill_1 FILLER_64_221 ();
 sg13g2_fill_2 FILLER_64_243 ();
 sg13g2_fill_1 FILLER_64_245 ();
 sg13g2_fill_2 FILLER_64_255 ();
 sg13g2_decap_8 FILLER_64_314 ();
 sg13g2_fill_2 FILLER_64_321 ();
 sg13g2_fill_1 FILLER_64_323 ();
 sg13g2_fill_2 FILLER_64_359 ();
 sg13g2_fill_1 FILLER_64_361 ();
 sg13g2_decap_8 FILLER_64_439 ();
 sg13g2_fill_1 FILLER_64_446 ();
 sg13g2_decap_4 FILLER_64_451 ();
 sg13g2_fill_1 FILLER_64_455 ();
 sg13g2_fill_2 FILLER_64_511 ();
 sg13g2_fill_1 FILLER_64_513 ();
 sg13g2_fill_2 FILLER_64_547 ();
 sg13g2_fill_2 FILLER_64_558 ();
 sg13g2_fill_1 FILLER_64_560 ();
 sg13g2_fill_2 FILLER_64_669 ();
 sg13g2_fill_1 FILLER_64_671 ();
 sg13g2_decap_8 FILLER_64_698 ();
 sg13g2_decap_8 FILLER_64_705 ();
 sg13g2_decap_8 FILLER_64_712 ();
 sg13g2_decap_8 FILLER_64_719 ();
 sg13g2_decap_8 FILLER_64_726 ();
 sg13g2_decap_8 FILLER_64_733 ();
 sg13g2_decap_8 FILLER_64_740 ();
 sg13g2_decap_8 FILLER_64_747 ();
 sg13g2_decap_8 FILLER_64_754 ();
 sg13g2_decap_8 FILLER_64_761 ();
 sg13g2_decap_8 FILLER_64_768 ();
 sg13g2_decap_8 FILLER_64_775 ();
 sg13g2_decap_8 FILLER_64_782 ();
 sg13g2_decap_8 FILLER_64_789 ();
 sg13g2_decap_8 FILLER_64_796 ();
 sg13g2_decap_8 FILLER_64_803 ();
 sg13g2_decap_8 FILLER_64_810 ();
 sg13g2_decap_8 FILLER_64_817 ();
 sg13g2_decap_8 FILLER_64_824 ();
 sg13g2_decap_8 FILLER_64_831 ();
 sg13g2_decap_8 FILLER_64_838 ();
 sg13g2_decap_8 FILLER_64_845 ();
 sg13g2_decap_8 FILLER_64_852 ();
 sg13g2_fill_2 FILLER_64_859 ();
 sg13g2_fill_1 FILLER_64_861 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_fill_2 FILLER_65_7 ();
 sg13g2_fill_1 FILLER_65_9 ();
 sg13g2_fill_2 FILLER_65_23 ();
 sg13g2_fill_2 FILLER_65_96 ();
 sg13g2_fill_1 FILLER_65_129 ();
 sg13g2_fill_2 FILLER_65_223 ();
 sg13g2_fill_2 FILLER_65_269 ();
 sg13g2_fill_1 FILLER_65_271 ();
 sg13g2_decap_8 FILLER_65_276 ();
 sg13g2_fill_2 FILLER_65_296 ();
 sg13g2_fill_1 FILLER_65_298 ();
 sg13g2_fill_1 FILLER_65_380 ();
 sg13g2_fill_1 FILLER_65_391 ();
 sg13g2_fill_2 FILLER_65_414 ();
 sg13g2_fill_1 FILLER_65_416 ();
 sg13g2_decap_8 FILLER_65_421 ();
 sg13g2_decap_8 FILLER_65_428 ();
 sg13g2_fill_1 FILLER_65_435 ();
 sg13g2_fill_1 FILLER_65_462 ();
 sg13g2_fill_1 FILLER_65_515 ();
 sg13g2_fill_1 FILLER_65_546 ();
 sg13g2_fill_2 FILLER_65_596 ();
 sg13g2_fill_1 FILLER_65_598 ();
 sg13g2_fill_1 FILLER_65_658 ();
 sg13g2_decap_8 FILLER_65_698 ();
 sg13g2_decap_8 FILLER_65_705 ();
 sg13g2_decap_8 FILLER_65_712 ();
 sg13g2_decap_8 FILLER_65_719 ();
 sg13g2_decap_8 FILLER_65_726 ();
 sg13g2_decap_8 FILLER_65_733 ();
 sg13g2_decap_8 FILLER_65_740 ();
 sg13g2_decap_8 FILLER_65_747 ();
 sg13g2_decap_8 FILLER_65_754 ();
 sg13g2_decap_8 FILLER_65_761 ();
 sg13g2_decap_8 FILLER_65_768 ();
 sg13g2_decap_8 FILLER_65_775 ();
 sg13g2_decap_8 FILLER_65_782 ();
 sg13g2_decap_8 FILLER_65_789 ();
 sg13g2_decap_8 FILLER_65_796 ();
 sg13g2_decap_8 FILLER_65_803 ();
 sg13g2_decap_8 FILLER_65_810 ();
 sg13g2_decap_8 FILLER_65_817 ();
 sg13g2_decap_8 FILLER_65_824 ();
 sg13g2_decap_8 FILLER_65_831 ();
 sg13g2_decap_8 FILLER_65_838 ();
 sg13g2_decap_8 FILLER_65_845 ();
 sg13g2_decap_8 FILLER_65_852 ();
 sg13g2_fill_2 FILLER_65_859 ();
 sg13g2_fill_1 FILLER_65_861 ();
 sg13g2_fill_2 FILLER_66_70 ();
 sg13g2_fill_1 FILLER_66_72 ();
 sg13g2_fill_1 FILLER_66_90 ();
 sg13g2_fill_2 FILLER_66_130 ();
 sg13g2_decap_8 FILLER_66_200 ();
 sg13g2_fill_1 FILLER_66_207 ();
 sg13g2_decap_4 FILLER_66_221 ();
 sg13g2_fill_2 FILLER_66_225 ();
 sg13g2_decap_8 FILLER_66_235 ();
 sg13g2_fill_2 FILLER_66_242 ();
 sg13g2_fill_2 FILLER_66_248 ();
 sg13g2_fill_2 FILLER_66_286 ();
 sg13g2_fill_1 FILLER_66_288 ();
 sg13g2_fill_1 FILLER_66_305 ();
 sg13g2_fill_2 FILLER_66_334 ();
 sg13g2_fill_2 FILLER_66_353 ();
 sg13g2_fill_1 FILLER_66_355 ();
 sg13g2_fill_2 FILLER_66_374 ();
 sg13g2_fill_1 FILLER_66_376 ();
 sg13g2_decap_4 FILLER_66_469 ();
 sg13g2_fill_1 FILLER_66_473 ();
 sg13g2_decap_4 FILLER_66_488 ();
 sg13g2_fill_2 FILLER_66_505 ();
 sg13g2_fill_1 FILLER_66_507 ();
 sg13g2_fill_2 FILLER_66_574 ();
 sg13g2_fill_1 FILLER_66_576 ();
 sg13g2_fill_2 FILLER_66_617 ();
 sg13g2_fill_1 FILLER_66_619 ();
 sg13g2_fill_2 FILLER_66_633 ();
 sg13g2_fill_1 FILLER_66_635 ();
 sg13g2_fill_1 FILLER_66_656 ();
 sg13g2_fill_2 FILLER_66_666 ();
 sg13g2_decap_8 FILLER_66_703 ();
 sg13g2_decap_8 FILLER_66_710 ();
 sg13g2_decap_8 FILLER_66_717 ();
 sg13g2_decap_8 FILLER_66_724 ();
 sg13g2_decap_8 FILLER_66_731 ();
 sg13g2_decap_8 FILLER_66_738 ();
 sg13g2_decap_8 FILLER_66_745 ();
 sg13g2_decap_8 FILLER_66_752 ();
 sg13g2_decap_8 FILLER_66_759 ();
 sg13g2_decap_8 FILLER_66_766 ();
 sg13g2_decap_8 FILLER_66_773 ();
 sg13g2_decap_8 FILLER_66_780 ();
 sg13g2_decap_8 FILLER_66_787 ();
 sg13g2_decap_8 FILLER_66_794 ();
 sg13g2_decap_8 FILLER_66_801 ();
 sg13g2_decap_8 FILLER_66_808 ();
 sg13g2_decap_8 FILLER_66_815 ();
 sg13g2_decap_8 FILLER_66_822 ();
 sg13g2_decap_8 FILLER_66_829 ();
 sg13g2_decap_8 FILLER_66_836 ();
 sg13g2_decap_8 FILLER_66_843 ();
 sg13g2_decap_8 FILLER_66_850 ();
 sg13g2_decap_4 FILLER_66_857 ();
 sg13g2_fill_1 FILLER_66_861 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_4 FILLER_67_7 ();
 sg13g2_fill_1 FILLER_67_15 ();
 sg13g2_fill_2 FILLER_67_35 ();
 sg13g2_fill_1 FILLER_67_37 ();
 sg13g2_fill_2 FILLER_67_55 ();
 sg13g2_fill_1 FILLER_67_57 ();
 sg13g2_fill_1 FILLER_67_84 ();
 sg13g2_fill_2 FILLER_67_227 ();
 sg13g2_fill_1 FILLER_67_234 ();
 sg13g2_decap_8 FILLER_67_246 ();
 sg13g2_fill_2 FILLER_67_253 ();
 sg13g2_decap_4 FILLER_67_265 ();
 sg13g2_decap_4 FILLER_67_311 ();
 sg13g2_fill_1 FILLER_67_406 ();
 sg13g2_fill_1 FILLER_67_416 ();
 sg13g2_fill_1 FILLER_67_462 ();
 sg13g2_fill_2 FILLER_67_499 ();
 sg13g2_fill_1 FILLER_67_510 ();
 sg13g2_fill_2 FILLER_67_525 ();
 sg13g2_fill_1 FILLER_67_573 ();
 sg13g2_fill_2 FILLER_67_610 ();
 sg13g2_fill_1 FILLER_67_612 ();
 sg13g2_fill_2 FILLER_67_618 ();
 sg13g2_fill_1 FILLER_67_620 ();
 sg13g2_fill_2 FILLER_67_646 ();
 sg13g2_fill_1 FILLER_67_648 ();
 sg13g2_decap_8 FILLER_67_698 ();
 sg13g2_decap_8 FILLER_67_705 ();
 sg13g2_decap_8 FILLER_67_712 ();
 sg13g2_decap_8 FILLER_67_719 ();
 sg13g2_decap_8 FILLER_67_726 ();
 sg13g2_decap_8 FILLER_67_733 ();
 sg13g2_decap_8 FILLER_67_740 ();
 sg13g2_decap_8 FILLER_67_747 ();
 sg13g2_decap_8 FILLER_67_754 ();
 sg13g2_decap_8 FILLER_67_761 ();
 sg13g2_decap_8 FILLER_67_768 ();
 sg13g2_decap_8 FILLER_67_775 ();
 sg13g2_decap_8 FILLER_67_782 ();
 sg13g2_decap_8 FILLER_67_789 ();
 sg13g2_decap_8 FILLER_67_796 ();
 sg13g2_decap_8 FILLER_67_803 ();
 sg13g2_decap_8 FILLER_67_810 ();
 sg13g2_decap_8 FILLER_67_817 ();
 sg13g2_decap_8 FILLER_67_824 ();
 sg13g2_decap_8 FILLER_67_831 ();
 sg13g2_decap_8 FILLER_67_838 ();
 sg13g2_decap_8 FILLER_67_845 ();
 sg13g2_decap_8 FILLER_67_852 ();
 sg13g2_fill_2 FILLER_67_859 ();
 sg13g2_fill_1 FILLER_67_861 ();
 sg13g2_fill_1 FILLER_68_26 ();
 sg13g2_fill_2 FILLER_68_50 ();
 sg13g2_fill_1 FILLER_68_66 ();
 sg13g2_fill_2 FILLER_68_173 ();
 sg13g2_fill_1 FILLER_68_210 ();
 sg13g2_decap_4 FILLER_68_253 ();
 sg13g2_fill_1 FILLER_68_257 ();
 sg13g2_fill_2 FILLER_68_295 ();
 sg13g2_fill_1 FILLER_68_297 ();
 sg13g2_fill_1 FILLER_68_320 ();
 sg13g2_fill_1 FILLER_68_331 ();
 sg13g2_fill_2 FILLER_68_342 ();
 sg13g2_fill_1 FILLER_68_344 ();
 sg13g2_fill_2 FILLER_68_354 ();
 sg13g2_fill_2 FILLER_68_399 ();
 sg13g2_fill_1 FILLER_68_401 ();
 sg13g2_fill_2 FILLER_68_432 ();
 sg13g2_fill_1 FILLER_68_457 ();
 sg13g2_fill_2 FILLER_68_503 ();
 sg13g2_fill_1 FILLER_68_505 ();
 sg13g2_fill_1 FILLER_68_529 ();
 sg13g2_fill_2 FILLER_68_581 ();
 sg13g2_fill_1 FILLER_68_610 ();
 sg13g2_fill_2 FILLER_68_693 ();
 sg13g2_fill_1 FILLER_68_695 ();
 sg13g2_decap_8 FILLER_68_705 ();
 sg13g2_decap_8 FILLER_68_712 ();
 sg13g2_decap_8 FILLER_68_719 ();
 sg13g2_decap_8 FILLER_68_726 ();
 sg13g2_decap_8 FILLER_68_733 ();
 sg13g2_decap_8 FILLER_68_740 ();
 sg13g2_decap_8 FILLER_68_747 ();
 sg13g2_decap_8 FILLER_68_754 ();
 sg13g2_decap_8 FILLER_68_761 ();
 sg13g2_decap_8 FILLER_68_768 ();
 sg13g2_decap_8 FILLER_68_775 ();
 sg13g2_decap_8 FILLER_68_782 ();
 sg13g2_decap_8 FILLER_68_789 ();
 sg13g2_decap_8 FILLER_68_796 ();
 sg13g2_decap_8 FILLER_68_803 ();
 sg13g2_decap_8 FILLER_68_810 ();
 sg13g2_decap_8 FILLER_68_817 ();
 sg13g2_decap_8 FILLER_68_824 ();
 sg13g2_decap_8 FILLER_68_831 ();
 sg13g2_decap_8 FILLER_68_838 ();
 sg13g2_decap_8 FILLER_68_845 ();
 sg13g2_decap_8 FILLER_68_852 ();
 sg13g2_fill_2 FILLER_68_859 ();
 sg13g2_fill_1 FILLER_68_861 ();
 sg13g2_fill_2 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_2 ();
 sg13g2_fill_1 FILLER_69_21 ();
 sg13g2_fill_2 FILLER_69_92 ();
 sg13g2_fill_2 FILLER_69_99 ();
 sg13g2_fill_1 FILLER_69_110 ();
 sg13g2_decap_4 FILLER_69_123 ();
 sg13g2_fill_1 FILLER_69_127 ();
 sg13g2_fill_2 FILLER_69_132 ();
 sg13g2_decap_4 FILLER_69_138 ();
 sg13g2_fill_1 FILLER_69_210 ();
 sg13g2_decap_4 FILLER_69_237 ();
 sg13g2_fill_1 FILLER_69_241 ();
 sg13g2_fill_2 FILLER_69_294 ();
 sg13g2_fill_2 FILLER_69_318 ();
 sg13g2_fill_1 FILLER_69_320 ();
 sg13g2_fill_1 FILLER_69_367 ();
 sg13g2_fill_2 FILLER_69_415 ();
 sg13g2_fill_1 FILLER_69_417 ();
 sg13g2_fill_2 FILLER_69_427 ();
 sg13g2_fill_2 FILLER_69_467 ();
 sg13g2_fill_2 FILLER_69_514 ();
 sg13g2_decap_8 FILLER_69_587 ();
 sg13g2_fill_1 FILLER_69_624 ();
 sg13g2_fill_2 FILLER_69_656 ();
 sg13g2_fill_1 FILLER_69_658 ();
 sg13g2_fill_2 FILLER_69_664 ();
 sg13g2_decap_8 FILLER_69_679 ();
 sg13g2_decap_8 FILLER_69_686 ();
 sg13g2_decap_8 FILLER_69_693 ();
 sg13g2_decap_8 FILLER_69_700 ();
 sg13g2_decap_8 FILLER_69_707 ();
 sg13g2_decap_8 FILLER_69_714 ();
 sg13g2_decap_8 FILLER_69_721 ();
 sg13g2_decap_8 FILLER_69_728 ();
 sg13g2_decap_8 FILLER_69_735 ();
 sg13g2_decap_8 FILLER_69_742 ();
 sg13g2_decap_8 FILLER_69_749 ();
 sg13g2_decap_8 FILLER_69_756 ();
 sg13g2_decap_8 FILLER_69_763 ();
 sg13g2_decap_8 FILLER_69_770 ();
 sg13g2_decap_8 FILLER_69_777 ();
 sg13g2_decap_8 FILLER_69_784 ();
 sg13g2_decap_8 FILLER_69_791 ();
 sg13g2_decap_8 FILLER_69_798 ();
 sg13g2_decap_8 FILLER_69_805 ();
 sg13g2_decap_8 FILLER_69_812 ();
 sg13g2_decap_8 FILLER_69_819 ();
 sg13g2_decap_8 FILLER_69_826 ();
 sg13g2_decap_8 FILLER_69_833 ();
 sg13g2_decap_8 FILLER_69_840 ();
 sg13g2_decap_8 FILLER_69_847 ();
 sg13g2_decap_8 FILLER_69_854 ();
 sg13g2_fill_1 FILLER_69_861 ();
 sg13g2_fill_1 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_27 ();
 sg13g2_fill_1 FILLER_70_29 ();
 sg13g2_fill_2 FILLER_70_57 ();
 sg13g2_fill_2 FILLER_70_80 ();
 sg13g2_decap_4 FILLER_70_112 ();
 sg13g2_fill_1 FILLER_70_116 ();
 sg13g2_fill_2 FILLER_70_143 ();
 sg13g2_fill_1 FILLER_70_145 ();
 sg13g2_fill_2 FILLER_70_155 ();
 sg13g2_fill_1 FILLER_70_161 ();
 sg13g2_decap_8 FILLER_70_166 ();
 sg13g2_fill_2 FILLER_70_230 ();
 sg13g2_fill_1 FILLER_70_232 ();
 sg13g2_fill_2 FILLER_70_240 ();
 sg13g2_fill_2 FILLER_70_304 ();
 sg13g2_fill_2 FILLER_70_311 ();
 sg13g2_fill_2 FILLER_70_318 ();
 sg13g2_fill_1 FILLER_70_320 ();
 sg13g2_fill_2 FILLER_70_339 ();
 sg13g2_fill_1 FILLER_70_350 ();
 sg13g2_fill_1 FILLER_70_395 ();
 sg13g2_decap_8 FILLER_70_441 ();
 sg13g2_fill_2 FILLER_70_448 ();
 sg13g2_fill_2 FILLER_70_455 ();
 sg13g2_fill_2 FILLER_70_493 ();
 sg13g2_fill_1 FILLER_70_495 ();
 sg13g2_fill_2 FILLER_70_561 ();
 sg13g2_fill_1 FILLER_70_567 ();
 sg13g2_fill_2 FILLER_70_576 ();
 sg13g2_fill_1 FILLER_70_619 ();
 sg13g2_fill_1 FILLER_70_624 ();
 sg13g2_fill_1 FILLER_70_660 ();
 sg13g2_decap_8 FILLER_70_674 ();
 sg13g2_decap_8 FILLER_70_681 ();
 sg13g2_decap_8 FILLER_70_688 ();
 sg13g2_decap_8 FILLER_70_695 ();
 sg13g2_decap_8 FILLER_70_702 ();
 sg13g2_decap_8 FILLER_70_709 ();
 sg13g2_decap_8 FILLER_70_716 ();
 sg13g2_decap_8 FILLER_70_723 ();
 sg13g2_decap_8 FILLER_70_730 ();
 sg13g2_decap_8 FILLER_70_737 ();
 sg13g2_decap_8 FILLER_70_744 ();
 sg13g2_decap_8 FILLER_70_751 ();
 sg13g2_decap_8 FILLER_70_758 ();
 sg13g2_decap_8 FILLER_70_765 ();
 sg13g2_decap_8 FILLER_70_772 ();
 sg13g2_decap_8 FILLER_70_779 ();
 sg13g2_decap_8 FILLER_70_786 ();
 sg13g2_decap_8 FILLER_70_793 ();
 sg13g2_decap_8 FILLER_70_800 ();
 sg13g2_decap_8 FILLER_70_807 ();
 sg13g2_decap_8 FILLER_70_814 ();
 sg13g2_decap_8 FILLER_70_821 ();
 sg13g2_decap_8 FILLER_70_828 ();
 sg13g2_decap_8 FILLER_70_835 ();
 sg13g2_decap_8 FILLER_70_842 ();
 sg13g2_decap_8 FILLER_70_849 ();
 sg13g2_decap_4 FILLER_70_856 ();
 sg13g2_fill_2 FILLER_70_860 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_33 ();
 sg13g2_fill_2 FILLER_71_45 ();
 sg13g2_fill_2 FILLER_71_133 ();
 sg13g2_fill_1 FILLER_71_135 ();
 sg13g2_decap_4 FILLER_71_192 ();
 sg13g2_fill_1 FILLER_71_209 ();
 sg13g2_fill_2 FILLER_71_219 ();
 sg13g2_fill_1 FILLER_71_221 ();
 sg13g2_fill_1 FILLER_71_248 ();
 sg13g2_fill_1 FILLER_71_275 ();
 sg13g2_fill_1 FILLER_71_329 ();
 sg13g2_fill_2 FILLER_71_339 ();
 sg13g2_fill_1 FILLER_71_377 ();
 sg13g2_fill_1 FILLER_71_403 ();
 sg13g2_fill_2 FILLER_71_418 ();
 sg13g2_fill_1 FILLER_71_456 ();
 sg13g2_fill_1 FILLER_71_461 ();
 sg13g2_fill_2 FILLER_71_473 ();
 sg13g2_fill_2 FILLER_71_494 ();
 sg13g2_fill_1 FILLER_71_505 ();
 sg13g2_fill_1 FILLER_71_520 ();
 sg13g2_fill_2 FILLER_71_557 ();
 sg13g2_fill_1 FILLER_71_559 ();
 sg13g2_decap_8 FILLER_71_665 ();
 sg13g2_decap_8 FILLER_71_672 ();
 sg13g2_decap_8 FILLER_71_679 ();
 sg13g2_decap_8 FILLER_71_686 ();
 sg13g2_decap_8 FILLER_71_693 ();
 sg13g2_decap_8 FILLER_71_700 ();
 sg13g2_decap_8 FILLER_71_707 ();
 sg13g2_decap_8 FILLER_71_714 ();
 sg13g2_decap_8 FILLER_71_721 ();
 sg13g2_decap_8 FILLER_71_728 ();
 sg13g2_decap_8 FILLER_71_735 ();
 sg13g2_decap_8 FILLER_71_742 ();
 sg13g2_decap_8 FILLER_71_749 ();
 sg13g2_decap_8 FILLER_71_756 ();
 sg13g2_decap_8 FILLER_71_763 ();
 sg13g2_decap_8 FILLER_71_770 ();
 sg13g2_decap_8 FILLER_71_777 ();
 sg13g2_decap_8 FILLER_71_784 ();
 sg13g2_decap_8 FILLER_71_791 ();
 sg13g2_decap_8 FILLER_71_798 ();
 sg13g2_decap_8 FILLER_71_805 ();
 sg13g2_decap_8 FILLER_71_812 ();
 sg13g2_decap_8 FILLER_71_819 ();
 sg13g2_decap_8 FILLER_71_826 ();
 sg13g2_decap_8 FILLER_71_833 ();
 sg13g2_decap_8 FILLER_71_840 ();
 sg13g2_decap_8 FILLER_71_847 ();
 sg13g2_decap_8 FILLER_71_854 ();
 sg13g2_fill_1 FILLER_71_861 ();
 sg13g2_fill_2 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_32 ();
 sg13g2_fill_2 FILLER_72_43 ();
 sg13g2_fill_1 FILLER_72_55 ();
 sg13g2_fill_1 FILLER_72_78 ();
 sg13g2_fill_2 FILLER_72_116 ();
 sg13g2_fill_1 FILLER_72_122 ();
 sg13g2_fill_2 FILLER_72_132 ();
 sg13g2_fill_1 FILLER_72_146 ();
 sg13g2_fill_1 FILLER_72_156 ();
 sg13g2_fill_2 FILLER_72_198 ();
 sg13g2_fill_1 FILLER_72_200 ();
 sg13g2_fill_1 FILLER_72_239 ();
 sg13g2_fill_1 FILLER_72_258 ();
 sg13g2_fill_1 FILLER_72_346 ();
 sg13g2_fill_1 FILLER_72_370 ();
 sg13g2_fill_2 FILLER_72_399 ();
 sg13g2_fill_1 FILLER_72_401 ();
 sg13g2_fill_1 FILLER_72_440 ();
 sg13g2_fill_1 FILLER_72_445 ();
 sg13g2_fill_2 FILLER_72_503 ();
 sg13g2_fill_1 FILLER_72_505 ();
 sg13g2_fill_1 FILLER_72_558 ();
 sg13g2_fill_2 FILLER_72_623 ();
 sg13g2_decap_8 FILLER_72_651 ();
 sg13g2_decap_8 FILLER_72_658 ();
 sg13g2_decap_8 FILLER_72_665 ();
 sg13g2_decap_8 FILLER_72_672 ();
 sg13g2_decap_8 FILLER_72_679 ();
 sg13g2_decap_8 FILLER_72_686 ();
 sg13g2_decap_8 FILLER_72_693 ();
 sg13g2_decap_8 FILLER_72_700 ();
 sg13g2_decap_8 FILLER_72_707 ();
 sg13g2_decap_8 FILLER_72_714 ();
 sg13g2_decap_8 FILLER_72_721 ();
 sg13g2_decap_8 FILLER_72_728 ();
 sg13g2_decap_8 FILLER_72_735 ();
 sg13g2_decap_8 FILLER_72_742 ();
 sg13g2_decap_8 FILLER_72_749 ();
 sg13g2_decap_8 FILLER_72_756 ();
 sg13g2_decap_8 FILLER_72_763 ();
 sg13g2_decap_8 FILLER_72_770 ();
 sg13g2_decap_8 FILLER_72_777 ();
 sg13g2_decap_8 FILLER_72_784 ();
 sg13g2_decap_8 FILLER_72_791 ();
 sg13g2_decap_8 FILLER_72_798 ();
 sg13g2_decap_8 FILLER_72_805 ();
 sg13g2_decap_8 FILLER_72_812 ();
 sg13g2_decap_8 FILLER_72_819 ();
 sg13g2_decap_8 FILLER_72_826 ();
 sg13g2_decap_8 FILLER_72_833 ();
 sg13g2_decap_8 FILLER_72_840 ();
 sg13g2_decap_8 FILLER_72_847 ();
 sg13g2_decap_8 FILLER_72_854 ();
 sg13g2_fill_1 FILLER_72_861 ();
 sg13g2_decap_4 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_30 ();
 sg13g2_fill_1 FILLER_73_32 ();
 sg13g2_fill_2 FILLER_73_61 ();
 sg13g2_fill_1 FILLER_73_63 ();
 sg13g2_fill_2 FILLER_73_82 ();
 sg13g2_fill_1 FILLER_73_84 ();
 sg13g2_fill_1 FILLER_73_139 ();
 sg13g2_fill_2 FILLER_73_149 ();
 sg13g2_fill_1 FILLER_73_151 ();
 sg13g2_fill_1 FILLER_73_156 ();
 sg13g2_fill_2 FILLER_73_187 ();
 sg13g2_fill_1 FILLER_73_189 ();
 sg13g2_fill_2 FILLER_73_207 ();
 sg13g2_fill_1 FILLER_73_209 ();
 sg13g2_fill_2 FILLER_73_236 ();
 sg13g2_fill_1 FILLER_73_267 ();
 sg13g2_fill_1 FILLER_73_282 ();
 sg13g2_fill_2 FILLER_73_321 ();
 sg13g2_fill_1 FILLER_73_336 ();
 sg13g2_fill_2 FILLER_73_429 ();
 sg13g2_fill_2 FILLER_73_443 ();
 sg13g2_fill_2 FILLER_73_487 ();
 sg13g2_fill_2 FILLER_73_548 ();
 sg13g2_fill_2 FILLER_73_568 ();
 sg13g2_fill_1 FILLER_73_578 ();
 sg13g2_decap_8 FILLER_73_647 ();
 sg13g2_decap_8 FILLER_73_654 ();
 sg13g2_decap_8 FILLER_73_661 ();
 sg13g2_decap_8 FILLER_73_668 ();
 sg13g2_decap_8 FILLER_73_675 ();
 sg13g2_decap_8 FILLER_73_682 ();
 sg13g2_decap_8 FILLER_73_689 ();
 sg13g2_decap_8 FILLER_73_696 ();
 sg13g2_decap_8 FILLER_73_703 ();
 sg13g2_decap_8 FILLER_73_710 ();
 sg13g2_decap_8 FILLER_73_717 ();
 sg13g2_decap_8 FILLER_73_724 ();
 sg13g2_decap_8 FILLER_73_731 ();
 sg13g2_decap_8 FILLER_73_738 ();
 sg13g2_decap_8 FILLER_73_745 ();
 sg13g2_decap_8 FILLER_73_752 ();
 sg13g2_decap_8 FILLER_73_759 ();
 sg13g2_decap_8 FILLER_73_766 ();
 sg13g2_decap_8 FILLER_73_773 ();
 sg13g2_decap_8 FILLER_73_780 ();
 sg13g2_decap_8 FILLER_73_787 ();
 sg13g2_decap_8 FILLER_73_794 ();
 sg13g2_decap_8 FILLER_73_801 ();
 sg13g2_decap_8 FILLER_73_808 ();
 sg13g2_decap_8 FILLER_73_815 ();
 sg13g2_decap_8 FILLER_73_822 ();
 sg13g2_decap_8 FILLER_73_829 ();
 sg13g2_decap_8 FILLER_73_836 ();
 sg13g2_decap_8 FILLER_73_843 ();
 sg13g2_decap_8 FILLER_73_850 ();
 sg13g2_decap_4 FILLER_73_857 ();
 sg13g2_fill_1 FILLER_73_861 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_7 ();
 sg13g2_fill_2 FILLER_74_35 ();
 sg13g2_fill_1 FILLER_74_37 ();
 sg13g2_fill_1 FILLER_74_52 ();
 sg13g2_fill_2 FILLER_74_98 ();
 sg13g2_fill_1 FILLER_74_104 ();
 sg13g2_fill_2 FILLER_74_114 ();
 sg13g2_fill_2 FILLER_74_152 ();
 sg13g2_decap_8 FILLER_74_206 ();
 sg13g2_fill_2 FILLER_74_213 ();
 sg13g2_fill_2 FILLER_74_271 ();
 sg13g2_fill_2 FILLER_74_349 ();
 sg13g2_fill_2 FILLER_74_355 ();
 sg13g2_fill_1 FILLER_74_374 ();
 sg13g2_fill_2 FILLER_74_398 ();
 sg13g2_fill_1 FILLER_74_444 ();
 sg13g2_fill_2 FILLER_74_471 ();
 sg13g2_fill_1 FILLER_74_473 ();
 sg13g2_fill_2 FILLER_74_500 ();
 sg13g2_fill_1 FILLER_74_502 ();
 sg13g2_fill_2 FILLER_74_544 ();
 sg13g2_fill_2 FILLER_74_582 ();
 sg13g2_fill_1 FILLER_74_601 ();
 sg13g2_fill_2 FILLER_74_616 ();
 sg13g2_decap_4 FILLER_74_636 ();
 sg13g2_fill_1 FILLER_74_640 ();
 sg13g2_decap_8 FILLER_74_650 ();
 sg13g2_decap_8 FILLER_74_657 ();
 sg13g2_decap_8 FILLER_74_664 ();
 sg13g2_decap_8 FILLER_74_671 ();
 sg13g2_decap_8 FILLER_74_678 ();
 sg13g2_decap_8 FILLER_74_685 ();
 sg13g2_decap_8 FILLER_74_692 ();
 sg13g2_decap_8 FILLER_74_699 ();
 sg13g2_decap_8 FILLER_74_706 ();
 sg13g2_decap_8 FILLER_74_713 ();
 sg13g2_decap_8 FILLER_74_720 ();
 sg13g2_decap_8 FILLER_74_727 ();
 sg13g2_decap_8 FILLER_74_734 ();
 sg13g2_decap_8 FILLER_74_741 ();
 sg13g2_decap_8 FILLER_74_748 ();
 sg13g2_decap_8 FILLER_74_755 ();
 sg13g2_decap_8 FILLER_74_762 ();
 sg13g2_decap_8 FILLER_74_769 ();
 sg13g2_decap_8 FILLER_74_776 ();
 sg13g2_decap_8 FILLER_74_783 ();
 sg13g2_decap_8 FILLER_74_790 ();
 sg13g2_decap_8 FILLER_74_797 ();
 sg13g2_decap_8 FILLER_74_804 ();
 sg13g2_decap_8 FILLER_74_811 ();
 sg13g2_decap_8 FILLER_74_818 ();
 sg13g2_decap_8 FILLER_74_825 ();
 sg13g2_decap_8 FILLER_74_832 ();
 sg13g2_decap_8 FILLER_74_839 ();
 sg13g2_decap_8 FILLER_74_846 ();
 sg13g2_decap_8 FILLER_74_853 ();
 sg13g2_fill_2 FILLER_74_860 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_fill_2 FILLER_75_14 ();
 sg13g2_fill_2 FILLER_75_61 ();
 sg13g2_fill_1 FILLER_75_63 ();
 sg13g2_fill_2 FILLER_75_118 ();
 sg13g2_fill_1 FILLER_75_120 ();
 sg13g2_fill_2 FILLER_75_142 ();
 sg13g2_fill_1 FILLER_75_144 ();
 sg13g2_decap_8 FILLER_75_212 ();
 sg13g2_fill_1 FILLER_75_219 ();
 sg13g2_fill_2 FILLER_75_252 ();
 sg13g2_fill_1 FILLER_75_293 ();
 sg13g2_fill_2 FILLER_75_302 ();
 sg13g2_fill_1 FILLER_75_345 ();
 sg13g2_fill_2 FILLER_75_435 ();
 sg13g2_fill_1 FILLER_75_437 ();
 sg13g2_fill_2 FILLER_75_537 ();
 sg13g2_decap_8 FILLER_75_620 ();
 sg13g2_decap_8 FILLER_75_627 ();
 sg13g2_decap_8 FILLER_75_634 ();
 sg13g2_decap_8 FILLER_75_641 ();
 sg13g2_decap_8 FILLER_75_648 ();
 sg13g2_decap_8 FILLER_75_655 ();
 sg13g2_decap_8 FILLER_75_662 ();
 sg13g2_decap_8 FILLER_75_669 ();
 sg13g2_decap_8 FILLER_75_676 ();
 sg13g2_decap_8 FILLER_75_683 ();
 sg13g2_decap_8 FILLER_75_690 ();
 sg13g2_decap_8 FILLER_75_697 ();
 sg13g2_decap_8 FILLER_75_704 ();
 sg13g2_decap_8 FILLER_75_711 ();
 sg13g2_decap_8 FILLER_75_718 ();
 sg13g2_decap_8 FILLER_75_725 ();
 sg13g2_decap_8 FILLER_75_732 ();
 sg13g2_decap_8 FILLER_75_739 ();
 sg13g2_decap_8 FILLER_75_746 ();
 sg13g2_decap_8 FILLER_75_753 ();
 sg13g2_decap_8 FILLER_75_760 ();
 sg13g2_decap_8 FILLER_75_767 ();
 sg13g2_decap_8 FILLER_75_774 ();
 sg13g2_decap_8 FILLER_75_781 ();
 sg13g2_decap_8 FILLER_75_788 ();
 sg13g2_decap_8 FILLER_75_795 ();
 sg13g2_decap_8 FILLER_75_802 ();
 sg13g2_decap_8 FILLER_75_809 ();
 sg13g2_decap_8 FILLER_75_816 ();
 sg13g2_decap_8 FILLER_75_823 ();
 sg13g2_decap_8 FILLER_75_830 ();
 sg13g2_decap_8 FILLER_75_837 ();
 sg13g2_decap_8 FILLER_75_844 ();
 sg13g2_decap_8 FILLER_75_851 ();
 sg13g2_decap_4 FILLER_75_858 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_fill_1 FILLER_76_103 ();
 sg13g2_fill_1 FILLER_76_138 ();
 sg13g2_fill_1 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_207 ();
 sg13g2_decap_8 FILLER_76_214 ();
 sg13g2_fill_2 FILLER_76_221 ();
 sg13g2_decap_8 FILLER_76_249 ();
 sg13g2_decap_8 FILLER_76_256 ();
 sg13g2_fill_1 FILLER_76_263 ();
 sg13g2_decap_4 FILLER_76_295 ();
 sg13g2_fill_1 FILLER_76_299 ();
 sg13g2_decap_4 FILLER_76_330 ();
 sg13g2_fill_1 FILLER_76_334 ();
 sg13g2_fill_1 FILLER_76_370 ();
 sg13g2_fill_2 FILLER_76_407 ();
 sg13g2_decap_4 FILLER_76_454 ();
 sg13g2_fill_1 FILLER_76_531 ();
 sg13g2_fill_2 FILLER_76_558 ();
 sg13g2_decap_8 FILLER_76_590 ();
 sg13g2_decap_8 FILLER_76_623 ();
 sg13g2_decap_8 FILLER_76_630 ();
 sg13g2_decap_8 FILLER_76_637 ();
 sg13g2_decap_8 FILLER_76_644 ();
 sg13g2_decap_8 FILLER_76_651 ();
 sg13g2_decap_8 FILLER_76_658 ();
 sg13g2_decap_8 FILLER_76_665 ();
 sg13g2_decap_8 FILLER_76_672 ();
 sg13g2_decap_8 FILLER_76_679 ();
 sg13g2_decap_8 FILLER_76_686 ();
 sg13g2_decap_8 FILLER_76_693 ();
 sg13g2_decap_8 FILLER_76_700 ();
 sg13g2_decap_8 FILLER_76_707 ();
 sg13g2_decap_8 FILLER_76_714 ();
 sg13g2_decap_8 FILLER_76_721 ();
 sg13g2_decap_8 FILLER_76_728 ();
 sg13g2_decap_8 FILLER_76_735 ();
 sg13g2_decap_8 FILLER_76_742 ();
 sg13g2_decap_8 FILLER_76_749 ();
 sg13g2_decap_8 FILLER_76_756 ();
 sg13g2_decap_8 FILLER_76_763 ();
 sg13g2_decap_8 FILLER_76_770 ();
 sg13g2_decap_8 FILLER_76_777 ();
 sg13g2_decap_8 FILLER_76_784 ();
 sg13g2_decap_8 FILLER_76_791 ();
 sg13g2_decap_8 FILLER_76_798 ();
 sg13g2_decap_8 FILLER_76_805 ();
 sg13g2_decap_8 FILLER_76_812 ();
 sg13g2_decap_8 FILLER_76_819 ();
 sg13g2_decap_8 FILLER_76_826 ();
 sg13g2_decap_8 FILLER_76_833 ();
 sg13g2_decap_8 FILLER_76_840 ();
 sg13g2_decap_8 FILLER_76_847 ();
 sg13g2_decap_8 FILLER_76_854 ();
 sg13g2_fill_1 FILLER_76_861 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_fill_2 FILLER_77_44 ();
 sg13g2_fill_1 FILLER_77_72 ();
 sg13g2_decap_4 FILLER_77_91 ();
 sg13g2_fill_1 FILLER_77_124 ();
 sg13g2_fill_1 FILLER_77_161 ();
 sg13g2_fill_2 FILLER_77_188 ();
 sg13g2_fill_1 FILLER_77_190 ();
 sg13g2_decap_8 FILLER_77_204 ();
 sg13g2_decap_8 FILLER_77_211 ();
 sg13g2_decap_8 FILLER_77_218 ();
 sg13g2_decap_8 FILLER_77_225 ();
 sg13g2_decap_8 FILLER_77_232 ();
 sg13g2_decap_8 FILLER_77_239 ();
 sg13g2_decap_8 FILLER_77_246 ();
 sg13g2_fill_2 FILLER_77_273 ();
 sg13g2_decap_4 FILLER_77_301 ();
 sg13g2_fill_2 FILLER_77_305 ();
 sg13g2_fill_1 FILLER_77_342 ();
 sg13g2_fill_2 FILLER_77_380 ();
 sg13g2_fill_1 FILLER_77_382 ();
 sg13g2_decap_8 FILLER_77_402 ();
 sg13g2_fill_1 FILLER_77_409 ();
 sg13g2_fill_1 FILLER_77_423 ();
 sg13g2_fill_1 FILLER_77_439 ();
 sg13g2_fill_1 FILLER_77_529 ();
 sg13g2_fill_1 FILLER_77_549 ();
 sg13g2_fill_1 FILLER_77_586 ();
 sg13g2_decap_8 FILLER_77_629 ();
 sg13g2_decap_8 FILLER_77_636 ();
 sg13g2_decap_8 FILLER_77_643 ();
 sg13g2_decap_8 FILLER_77_650 ();
 sg13g2_decap_8 FILLER_77_657 ();
 sg13g2_decap_8 FILLER_77_664 ();
 sg13g2_decap_8 FILLER_77_671 ();
 sg13g2_decap_8 FILLER_77_678 ();
 sg13g2_decap_8 FILLER_77_685 ();
 sg13g2_decap_8 FILLER_77_692 ();
 sg13g2_decap_8 FILLER_77_699 ();
 sg13g2_decap_8 FILLER_77_706 ();
 sg13g2_decap_8 FILLER_77_713 ();
 sg13g2_decap_8 FILLER_77_720 ();
 sg13g2_decap_8 FILLER_77_727 ();
 sg13g2_decap_8 FILLER_77_734 ();
 sg13g2_decap_8 FILLER_77_741 ();
 sg13g2_decap_8 FILLER_77_748 ();
 sg13g2_decap_8 FILLER_77_755 ();
 sg13g2_decap_8 FILLER_77_762 ();
 sg13g2_decap_8 FILLER_77_769 ();
 sg13g2_decap_8 FILLER_77_776 ();
 sg13g2_decap_8 FILLER_77_783 ();
 sg13g2_decap_8 FILLER_77_790 ();
 sg13g2_decap_8 FILLER_77_797 ();
 sg13g2_decap_8 FILLER_77_804 ();
 sg13g2_decap_8 FILLER_77_811 ();
 sg13g2_decap_8 FILLER_77_818 ();
 sg13g2_decap_8 FILLER_77_825 ();
 sg13g2_decap_8 FILLER_77_832 ();
 sg13g2_decap_8 FILLER_77_839 ();
 sg13g2_decap_8 FILLER_77_846 ();
 sg13g2_decap_8 FILLER_77_853 ();
 sg13g2_fill_2 FILLER_77_860 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_4 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_43 ();
 sg13g2_fill_2 FILLER_78_50 ();
 sg13g2_fill_1 FILLER_78_52 ();
 sg13g2_decap_8 FILLER_78_89 ();
 sg13g2_decap_8 FILLER_78_96 ();
 sg13g2_fill_2 FILLER_78_103 ();
 sg13g2_fill_1 FILLER_78_105 ();
 sg13g2_fill_2 FILLER_78_122 ();
 sg13g2_fill_2 FILLER_78_128 ();
 sg13g2_fill_1 FILLER_78_130 ();
 sg13g2_fill_1 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_145 ();
 sg13g2_decap_4 FILLER_78_152 ();
 sg13g2_fill_1 FILLER_78_156 ();
 sg13g2_decap_8 FILLER_78_162 ();
 sg13g2_decap_4 FILLER_78_169 ();
 sg13g2_decap_8 FILLER_78_186 ();
 sg13g2_decap_8 FILLER_78_193 ();
 sg13g2_decap_8 FILLER_78_200 ();
 sg13g2_decap_8 FILLER_78_207 ();
 sg13g2_decap_8 FILLER_78_214 ();
 sg13g2_decap_8 FILLER_78_221 ();
 sg13g2_decap_8 FILLER_78_228 ();
 sg13g2_decap_8 FILLER_78_235 ();
 sg13g2_decap_8 FILLER_78_242 ();
 sg13g2_decap_8 FILLER_78_249 ();
 sg13g2_decap_8 FILLER_78_256 ();
 sg13g2_decap_8 FILLER_78_263 ();
 sg13g2_decap_4 FILLER_78_270 ();
 sg13g2_fill_1 FILLER_78_274 ();
 sg13g2_decap_8 FILLER_78_279 ();
 sg13g2_decap_8 FILLER_78_290 ();
 sg13g2_decap_4 FILLER_78_297 ();
 sg13g2_fill_2 FILLER_78_301 ();
 sg13g2_decap_4 FILLER_78_313 ();
 sg13g2_fill_1 FILLER_78_317 ();
 sg13g2_fill_1 FILLER_78_384 ();
 sg13g2_fill_2 FILLER_78_394 ();
 sg13g2_decap_4 FILLER_78_442 ();
 sg13g2_fill_1 FILLER_78_446 ();
 sg13g2_fill_2 FILLER_78_457 ();
 sg13g2_fill_1 FILLER_78_459 ();
 sg13g2_fill_2 FILLER_78_477 ();
 sg13g2_fill_2 FILLER_78_497 ();
 sg13g2_fill_1 FILLER_78_499 ();
 sg13g2_fill_2 FILLER_78_536 ();
 sg13g2_fill_1 FILLER_78_577 ();
 sg13g2_decap_8 FILLER_78_619 ();
 sg13g2_decap_8 FILLER_78_626 ();
 sg13g2_decap_8 FILLER_78_633 ();
 sg13g2_decap_8 FILLER_78_640 ();
 sg13g2_decap_8 FILLER_78_647 ();
 sg13g2_decap_8 FILLER_78_654 ();
 sg13g2_decap_8 FILLER_78_661 ();
 sg13g2_decap_8 FILLER_78_668 ();
 sg13g2_decap_8 FILLER_78_675 ();
 sg13g2_decap_8 FILLER_78_682 ();
 sg13g2_decap_8 FILLER_78_689 ();
 sg13g2_decap_8 FILLER_78_696 ();
 sg13g2_decap_8 FILLER_78_703 ();
 sg13g2_decap_8 FILLER_78_710 ();
 sg13g2_decap_8 FILLER_78_717 ();
 sg13g2_decap_8 FILLER_78_724 ();
 sg13g2_decap_8 FILLER_78_731 ();
 sg13g2_decap_8 FILLER_78_738 ();
 sg13g2_decap_8 FILLER_78_745 ();
 sg13g2_decap_8 FILLER_78_752 ();
 sg13g2_decap_8 FILLER_78_759 ();
 sg13g2_decap_8 FILLER_78_766 ();
 sg13g2_decap_8 FILLER_78_773 ();
 sg13g2_decap_8 FILLER_78_780 ();
 sg13g2_decap_8 FILLER_78_787 ();
 sg13g2_decap_8 FILLER_78_794 ();
 sg13g2_decap_8 FILLER_78_801 ();
 sg13g2_decap_8 FILLER_78_808 ();
 sg13g2_decap_8 FILLER_78_815 ();
 sg13g2_decap_8 FILLER_78_822 ();
 sg13g2_decap_8 FILLER_78_829 ();
 sg13g2_decap_8 FILLER_78_836 ();
 sg13g2_decap_8 FILLER_78_843 ();
 sg13g2_decap_8 FILLER_78_850 ();
 sg13g2_decap_4 FILLER_78_857 ();
 sg13g2_fill_1 FILLER_78_861 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_fill_1 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_61 ();
 sg13g2_decap_4 FILLER_79_68 ();
 sg13g2_fill_2 FILLER_79_72 ();
 sg13g2_decap_8 FILLER_79_78 ();
 sg13g2_decap_8 FILLER_79_85 ();
 sg13g2_decap_8 FILLER_79_92 ();
 sg13g2_decap_8 FILLER_79_99 ();
 sg13g2_decap_8 FILLER_79_106 ();
 sg13g2_decap_8 FILLER_79_113 ();
 sg13g2_decap_8 FILLER_79_120 ();
 sg13g2_decap_8 FILLER_79_127 ();
 sg13g2_decap_8 FILLER_79_134 ();
 sg13g2_decap_8 FILLER_79_141 ();
 sg13g2_decap_8 FILLER_79_148 ();
 sg13g2_decap_8 FILLER_79_155 ();
 sg13g2_decap_8 FILLER_79_162 ();
 sg13g2_decap_8 FILLER_79_169 ();
 sg13g2_decap_8 FILLER_79_176 ();
 sg13g2_decap_8 FILLER_79_183 ();
 sg13g2_decap_8 FILLER_79_190 ();
 sg13g2_decap_8 FILLER_79_197 ();
 sg13g2_decap_8 FILLER_79_204 ();
 sg13g2_decap_8 FILLER_79_211 ();
 sg13g2_decap_8 FILLER_79_218 ();
 sg13g2_decap_8 FILLER_79_225 ();
 sg13g2_decap_8 FILLER_79_232 ();
 sg13g2_decap_8 FILLER_79_239 ();
 sg13g2_decap_8 FILLER_79_246 ();
 sg13g2_decap_8 FILLER_79_253 ();
 sg13g2_decap_8 FILLER_79_260 ();
 sg13g2_decap_8 FILLER_79_267 ();
 sg13g2_decap_8 FILLER_79_274 ();
 sg13g2_decap_8 FILLER_79_281 ();
 sg13g2_decap_8 FILLER_79_288 ();
 sg13g2_decap_8 FILLER_79_295 ();
 sg13g2_decap_8 FILLER_79_302 ();
 sg13g2_decap_8 FILLER_79_309 ();
 sg13g2_decap_8 FILLER_79_316 ();
 sg13g2_decap_8 FILLER_79_323 ();
 sg13g2_decap_8 FILLER_79_330 ();
 sg13g2_decap_8 FILLER_79_337 ();
 sg13g2_fill_1 FILLER_79_344 ();
 sg13g2_decap_8 FILLER_79_349 ();
 sg13g2_decap_8 FILLER_79_356 ();
 sg13g2_decap_4 FILLER_79_363 ();
 sg13g2_fill_1 FILLER_79_367 ();
 sg13g2_decap_8 FILLER_79_372 ();
 sg13g2_decap_8 FILLER_79_379 ();
 sg13g2_decap_8 FILLER_79_386 ();
 sg13g2_fill_1 FILLER_79_393 ();
 sg13g2_fill_1 FILLER_79_422 ();
 sg13g2_decap_4 FILLER_79_449 ();
 sg13g2_decap_4 FILLER_79_479 ();
 sg13g2_decap_8 FILLER_79_531 ();
 sg13g2_decap_4 FILLER_79_538 ();
 sg13g2_decap_8 FILLER_79_560 ();
 sg13g2_fill_2 FILLER_79_567 ();
 sg13g2_fill_1 FILLER_79_569 ();
 sg13g2_decap_8 FILLER_79_579 ();
 sg13g2_decap_8 FILLER_79_586 ();
 sg13g2_decap_4 FILLER_79_593 ();
 sg13g2_fill_2 FILLER_79_597 ();
 sg13g2_decap_8 FILLER_79_603 ();
 sg13g2_decap_8 FILLER_79_610 ();
 sg13g2_decap_8 FILLER_79_617 ();
 sg13g2_decap_8 FILLER_79_624 ();
 sg13g2_decap_8 FILLER_79_631 ();
 sg13g2_decap_8 FILLER_79_638 ();
 sg13g2_decap_8 FILLER_79_645 ();
 sg13g2_decap_8 FILLER_79_652 ();
 sg13g2_decap_8 FILLER_79_659 ();
 sg13g2_decap_8 FILLER_79_666 ();
 sg13g2_decap_8 FILLER_79_673 ();
 sg13g2_decap_8 FILLER_79_680 ();
 sg13g2_decap_8 FILLER_79_687 ();
 sg13g2_decap_8 FILLER_79_694 ();
 sg13g2_decap_8 FILLER_79_701 ();
 sg13g2_decap_8 FILLER_79_708 ();
 sg13g2_decap_8 FILLER_79_715 ();
 sg13g2_decap_8 FILLER_79_722 ();
 sg13g2_decap_8 FILLER_79_729 ();
 sg13g2_decap_8 FILLER_79_736 ();
 sg13g2_decap_8 FILLER_79_743 ();
 sg13g2_decap_8 FILLER_79_750 ();
 sg13g2_decap_8 FILLER_79_757 ();
 sg13g2_decap_8 FILLER_79_764 ();
 sg13g2_decap_8 FILLER_79_771 ();
 sg13g2_decap_8 FILLER_79_778 ();
 sg13g2_decap_8 FILLER_79_785 ();
 sg13g2_decap_8 FILLER_79_792 ();
 sg13g2_decap_8 FILLER_79_799 ();
 sg13g2_decap_8 FILLER_79_806 ();
 sg13g2_decap_8 FILLER_79_813 ();
 sg13g2_decap_8 FILLER_79_820 ();
 sg13g2_decap_8 FILLER_79_827 ();
 sg13g2_decap_8 FILLER_79_834 ();
 sg13g2_decap_8 FILLER_79_841 ();
 sg13g2_decap_8 FILLER_79_848 ();
 sg13g2_decap_8 FILLER_79_855 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_208 ();
 sg13g2_decap_8 FILLER_80_215 ();
 sg13g2_decap_8 FILLER_80_222 ();
 sg13g2_decap_8 FILLER_80_229 ();
 sg13g2_decap_8 FILLER_80_236 ();
 sg13g2_decap_8 FILLER_80_243 ();
 sg13g2_decap_8 FILLER_80_250 ();
 sg13g2_decap_8 FILLER_80_257 ();
 sg13g2_decap_8 FILLER_80_264 ();
 sg13g2_decap_8 FILLER_80_271 ();
 sg13g2_decap_8 FILLER_80_278 ();
 sg13g2_decap_8 FILLER_80_285 ();
 sg13g2_decap_8 FILLER_80_292 ();
 sg13g2_decap_8 FILLER_80_299 ();
 sg13g2_decap_4 FILLER_80_306 ();
 sg13g2_fill_2 FILLER_80_310 ();
 sg13g2_decap_8 FILLER_80_316 ();
 sg13g2_decap_8 FILLER_80_323 ();
 sg13g2_decap_8 FILLER_80_330 ();
 sg13g2_decap_8 FILLER_80_337 ();
 sg13g2_decap_8 FILLER_80_344 ();
 sg13g2_decap_8 FILLER_80_351 ();
 sg13g2_decap_8 FILLER_80_358 ();
 sg13g2_decap_8 FILLER_80_365 ();
 sg13g2_decap_8 FILLER_80_372 ();
 sg13g2_decap_8 FILLER_80_379 ();
 sg13g2_decap_8 FILLER_80_386 ();
 sg13g2_fill_2 FILLER_80_393 ();
 sg13g2_fill_1 FILLER_80_395 ();
 sg13g2_fill_1 FILLER_80_405 ();
 sg13g2_decap_8 FILLER_80_410 ();
 sg13g2_decap_8 FILLER_80_417 ();
 sg13g2_fill_2 FILLER_80_424 ();
 sg13g2_fill_1 FILLER_80_426 ();
 sg13g2_decap_8 FILLER_80_449 ();
 sg13g2_decap_8 FILLER_80_456 ();
 sg13g2_fill_2 FILLER_80_463 ();
 sg13g2_decap_8 FILLER_80_474 ();
 sg13g2_decap_8 FILLER_80_481 ();
 sg13g2_decap_4 FILLER_80_488 ();
 sg13g2_fill_2 FILLER_80_492 ();
 sg13g2_decap_8 FILLER_80_498 ();
 sg13g2_decap_8 FILLER_80_505 ();
 sg13g2_decap_8 FILLER_80_512 ();
 sg13g2_decap_8 FILLER_80_519 ();
 sg13g2_decap_8 FILLER_80_526 ();
 sg13g2_decap_8 FILLER_80_533 ();
 sg13g2_decap_8 FILLER_80_540 ();
 sg13g2_fill_2 FILLER_80_547 ();
 sg13g2_decap_8 FILLER_80_553 ();
 sg13g2_decap_8 FILLER_80_560 ();
 sg13g2_decap_8 FILLER_80_567 ();
 sg13g2_decap_8 FILLER_80_574 ();
 sg13g2_decap_8 FILLER_80_581 ();
 sg13g2_decap_8 FILLER_80_588 ();
 sg13g2_decap_8 FILLER_80_595 ();
 sg13g2_decap_8 FILLER_80_602 ();
 sg13g2_decap_8 FILLER_80_609 ();
 sg13g2_decap_8 FILLER_80_616 ();
 sg13g2_decap_8 FILLER_80_623 ();
 sg13g2_decap_8 FILLER_80_630 ();
 sg13g2_decap_8 FILLER_80_637 ();
 sg13g2_decap_8 FILLER_80_644 ();
 sg13g2_decap_8 FILLER_80_651 ();
 sg13g2_decap_8 FILLER_80_658 ();
 sg13g2_decap_8 FILLER_80_665 ();
 sg13g2_decap_8 FILLER_80_672 ();
 sg13g2_decap_8 FILLER_80_679 ();
 sg13g2_decap_8 FILLER_80_686 ();
 sg13g2_decap_8 FILLER_80_693 ();
 sg13g2_decap_8 FILLER_80_700 ();
 sg13g2_decap_8 FILLER_80_707 ();
 sg13g2_decap_8 FILLER_80_714 ();
 sg13g2_decap_8 FILLER_80_721 ();
 sg13g2_decap_8 FILLER_80_728 ();
 sg13g2_decap_8 FILLER_80_735 ();
 sg13g2_decap_8 FILLER_80_742 ();
 sg13g2_decap_8 FILLER_80_749 ();
 sg13g2_decap_8 FILLER_80_756 ();
 sg13g2_decap_8 FILLER_80_763 ();
 sg13g2_decap_8 FILLER_80_770 ();
 sg13g2_decap_8 FILLER_80_777 ();
 sg13g2_decap_8 FILLER_80_784 ();
 sg13g2_decap_8 FILLER_80_791 ();
 sg13g2_decap_8 FILLER_80_798 ();
 sg13g2_decap_8 FILLER_80_805 ();
 sg13g2_decap_8 FILLER_80_812 ();
 sg13g2_decap_8 FILLER_80_819 ();
 sg13g2_decap_8 FILLER_80_826 ();
 sg13g2_decap_8 FILLER_80_833 ();
 sg13g2_decap_8 FILLER_80_840 ();
 sg13g2_decap_8 FILLER_80_847 ();
 sg13g2_decap_8 FILLER_80_854 ();
 sg13g2_fill_1 FILLER_80_861 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
endmodule

module tt_um_moody_mimosa (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire \actions.clk ;
 wire \actions.development_stage[0] ;
 wire \actions.development_stage[1] ;
 wire \actions.is_asleep ;
 wire \actions.next_action[0] ;
 wire \actions.next_action[1] ;
 wire \actions.next_action[2] ;
 wire \actions.next_action[4] ;
 wire \actions.next_action[5] ;
 wire \actions.next_action[6] ;
 wire \actions.next_action[7] ;
 wire \actions.vital_energy_level[0] ;
 wire \actions.vital_energy_level[1] ;
 wire \counter_.count[0] ;
 wire \counter_.count[1] ;
 wire \counter_.count[2] ;
 wire \counter_.count[3] ;
 wire \development_stage_sys.dev_stage_reg.cry ;
 wire \development_stage_sys.dev_stage_reg.is_ill ;
 wire \development_stage_sys.development_stage_level[0] ;
 wire \development_stage_sys.development_stage_level[1] ;
 wire \development_stage_sys.development_stage_level[2] ;
 wire \development_stage_sys.development_stage_level[3] ;
 wire \development_stage_sys.development_stage_level[4] ;
 wire \development_stage_sys.development_stage_level[5] ;
 wire \development_stage_sys.development_stage_level[6] ;
 wire \emotions.CORT[0] ;
 wire \emotions.CORT[1] ;
 wire \emotions.DOP[0] ;
 wire \emotions.DOP[1] ;
 wire \emotions.GABA[0] ;
 wire \emotions.GABA[1] ;
 wire \emotions.NE[0] ;
 wire \emotions.NE[1] ;
 wire \emotions.SER[0] ;
 wire \emotions.SER[1] ;
 wire \heartbeat_divider.counter[0] ;
 wire \heartbeat_divider.counter[10] ;
 wire \heartbeat_divider.counter[11] ;
 wire \heartbeat_divider.counter[12] ;
 wire \heartbeat_divider.counter[1] ;
 wire \heartbeat_divider.counter[2] ;
 wire \heartbeat_divider.counter[3] ;
 wire \heartbeat_divider.counter[4] ;
 wire \heartbeat_divider.counter[5] ;
 wire \heartbeat_divider.counter[6] ;
 wire \heartbeat_divider.counter[7] ;
 wire \heartbeat_divider.counter[8] ;
 wire \heartbeat_divider.counter[9] ;
 wire \illness_sys.illness[0] ;
 wire \illness_sys.illness[1] ;
 wire \illness_sys.illness[2] ;
 wire \illness_sys.illness[3] ;
 wire \illness_sys.illness[4] ;
 wire \illness_sys.illness[5] ;
 wire \illness_sys.illness[6] ;
 wire \illness_sys.illness[7] ;
 wire \illness_sys.illness[8] ;
 wire \neurotransmitter.cortisol_system.cortisol[0] ;
 wire \neurotransmitter.cortisol_system.cortisol[1] ;
 wire \neurotransmitter.cortisol_system.cortisol[2] ;
 wire \neurotransmitter.cortisol_system.cortisol[3] ;
 wire \neurotransmitter.cortisol_system.cortisol[4] ;
 wire \neurotransmitter.cortisol_system.cortisol_regulator.CORT[0] ;
 wire \neurotransmitter.cortisol_system.cortisol_regulator.CORT[1] ;
 wire \neurotransmitter.cortisol_system.cortisol_regulator.DOP[0] ;
 wire \neurotransmitter.cortisol_system.cortisol_regulator.DOP[1] ;
 wire \neurotransmitter.cortisol_system.cortisol_regulator.GABA[0] ;
 wire \neurotransmitter.cortisol_system.cortisol_regulator.GABA[1] ;
 wire \neurotransmitter.cortisol_system.cortisol_regulator.NE[0] ;
 wire \neurotransmitter.cortisol_system.cortisol_regulator.NE[1] ;
 wire \neurotransmitter.cortisol_system.cortisol_regulator.SER[0] ;
 wire \neurotransmitter.cortisol_system.cortisol_regulator.SER[1] ;
 wire \neurotransmitter.cortisol_system.cortisol_regulator.babble ;
 wire \neurotransmitter.cortisol_system.cortisol_regulator.eat ;
 wire \neurotransmitter.cortisol_system.cortisol_regulator.idle ;
 wire \neurotransmitter.cortisol_system.cortisol_regulator.kick_legs ;
 wire \neurotransmitter.cortisol_system.cortisol_regulator.play ;
 wire \neurotransmitter.cortisol_system.cortisol_regulator.smile ;
 wire \neurotransmitter.dopamine_system.dopamine[0] ;
 wire \neurotransmitter.dopamine_system.dopamine[1] ;
 wire \neurotransmitter.dopamine_system.dopamine[2] ;
 wire \neurotransmitter.dopamine_system.dopamine[3] ;
 wire \neurotransmitter.dopamine_system.dopamine[4] ;
 wire \neurotransmitter.gaba_system.gaba[0] ;
 wire \neurotransmitter.gaba_system.gaba[1] ;
 wire \neurotransmitter.gaba_system.gaba[2] ;
 wire \neurotransmitter.gaba_system.gaba[3] ;
 wire \neurotransmitter.gaba_system.gaba[4] ;
 wire \neurotransmitter.norepinephrine_system.norepinephrine[0] ;
 wire \neurotransmitter.norepinephrine_system.norepinephrine[1] ;
 wire \neurotransmitter.norepinephrine_system.norepinephrine[2] ;
 wire \neurotransmitter.norepinephrine_system.norepinephrine[3] ;
 wire \neurotransmitter.serotonin_system.serotonin[0] ;
 wire \neurotransmitter.serotonin_system.serotonin[1] ;
 wire \neurotransmitter.serotonin_system.serotonin[2] ;
 wire \neurotransmitter.serotonin_system.serotonin[3] ;
 wire \neurotransmitter.serotonin_system.serotonin[4] ;
 wire \nourishment.glucose[0] ;
 wire \nourishment.glucose[1] ;
 wire \nourishment.glucose[2] ;
 wire \nourishment.glucose[3] ;
 wire \nourishment.glucose[4] ;
 wire \nourishment.glucose[5] ;
 wire \nourishment.glucose[6] ;
 wire \nourishment.glucose[7] ;
 wire \speech_planner_.variant_bit ;
 wire spi_cs;
 wire spi_mosi;
 wire spi_sck;
 wire \talking.address_reg[10] ;
 wire \talking.address_reg[11] ;
 wire \talking.address_reg[12] ;
 wire \talking.address_reg[13] ;
 wire \talking.address_reg[14] ;
 wire \talking.address_reg[15] ;
 wire \talking.address_reg[5] ;
 wire \talking.address_reg[6] ;
 wire \talking.address_reg[7] ;
 wire \talking.address_reg[8] ;
 wire \talking.address_reg[9] ;
 wire \talking.byte_count[0] ;
 wire \talking.byte_count[1] ;
 wire \talking.byte_count[2] ;
 wire \talking.byte_count[3] ;
 wire \talking.byte_count[4] ;
 wire \talking.byte_count[5] ;
 wire \talking.skip_address_bytes[0] ;
 wire \talking.skip_address_bytes[1] ;
 wire \talking.spi_bit_count[0] ;
 wire \talking.spi_bit_count[1] ;
 wire \talking.spi_bit_count[2] ;
 wire \talking.spi_bit_count[3] ;
 wire \talking.spi_shift_reg[0] ;
 wire \talking.spi_shift_reg[1] ;
 wire \talking.spi_shift_reg[2] ;
 wire \talking.spi_shift_reg[3] ;
 wire \talking.spi_shift_reg[4] ;
 wire \talking.spi_shift_reg[5] ;
 wire \talking.spi_shift_reg[6] ;
 wire \talking.state[0] ;
 wire \talking.state[1] ;
 wire \talking.state[2] ;
 wire \talking.uart_active ;
 wire \talking.uart_bit_count[0] ;
 wire \talking.uart_bit_count[1] ;
 wire \talking.uart_bit_count[2] ;
 wire \talking.uart_bit_count[3] ;
 wire \talking.uart_shift_reg[0] ;
 wire \talking.uart_shift_reg[1] ;
 wire \talking.uart_shift_reg[2] ;
 wire \talking.uart_shift_reg[3] ;
 wire \talking.uart_shift_reg[4] ;
 wire \talking.uart_shift_reg[5] ;
 wire \talking.uart_shift_reg[6] ;
 wire \talking.uart_shift_reg[7] ;
 wire \talking.uart_shift_reg[8] ;
 wire \talking.uart_shift_reg[9] ;
 wire \talking.uart_tx ;
 wire net13;
 wire net14;
 wire net15;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire clknet_0_clk;
 wire net16;
 wire net17;
 wire net18;
 wire \vital_energy_sys.vital_energy[0] ;
 wire \vital_energy_sys.vital_energy[1] ;
 wire \vital_energy_sys.vital_energy[2] ;
 wire \vital_energy_sys.vital_energy[3] ;
 wire \vital_energy_sys.vital_energy[4] ;
 wire \vital_energy_sys.vital_energy[5] ;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;

 sg13g2_inv_1 _1492_ (.Y(_0838_),
    .A(net27));
 sg13g2_inv_1 _1493_ (.Y(_0839_),
    .A(net29));
 sg13g2_inv_1 _1494_ (.Y(_0840_),
    .A(_0070_));
 sg13g2_inv_1 _1495_ (.Y(_0841_),
    .A(net481));
 sg13g2_inv_1 _1496_ (.Y(_0842_),
    .A(\emotions.NE[0] ));
 sg13g2_inv_1 _1497_ (.Y(_0843_),
    .A(\emotions.CORT[0] ));
 sg13g2_inv_2 _1498_ (.Y(_0844_),
    .A(net462));
 sg13g2_inv_1 _1499_ (.Y(_0845_),
    .A(\emotions.GABA[1] ));
 sg13g2_inv_1 _1500_ (.Y(_0846_),
    .A(\nourishment.glucose[6] ));
 sg13g2_inv_1 _1501_ (.Y(_0847_),
    .A(net465));
 sg13g2_inv_4 _1502_ (.A(net476),
    .Y(_0848_));
 sg13g2_inv_2 _1503_ (.Y(_0849_),
    .A(\emotions.DOP[1] ));
 sg13g2_inv_2 _1504_ (.Y(_0850_),
    .A(net473));
 sg13g2_inv_1 _1505_ (.Y(_0851_),
    .A(_0046_));
 sg13g2_inv_1 _1506_ (.Y(_0852_),
    .A(\development_stage_sys.development_stage_level[1] ));
 sg13g2_inv_1 _1507_ (.Y(_0853_),
    .A(\development_stage_sys.development_stage_level[0] ));
 sg13g2_inv_2 _1508_ (.Y(_0854_),
    .A(\development_stage_sys.development_stage_level[4] ));
 sg13g2_inv_1 _1509_ (.Y(_0855_),
    .A(net457));
 sg13g2_inv_1 _1510_ (.Y(_0856_),
    .A(\nourishment.glucose[0] ));
 sg13g2_inv_1 _1511_ (.Y(_0857_),
    .A(\neurotransmitter.cortisol_system.cortisol_regulator.GABA[1] ));
 sg13g2_inv_1 _1512_ (.Y(_0858_),
    .A(\neurotransmitter.cortisol_system.cortisol_regulator.play ));
 sg13g2_inv_1 _1513_ (.Y(_0859_),
    .A(\neurotransmitter.dopamine_system.dopamine[0] ));
 sg13g2_inv_1 _1514_ (.Y(_0860_),
    .A(\talking.uart_active ));
 sg13g2_inv_1 _1515_ (.Y(_0861_),
    .A(\counter_.count[3] ));
 sg13g2_inv_1 _1516_ (.Y(_0862_),
    .A(\neurotransmitter.gaba_system.gaba[0] ));
 sg13g2_inv_1 _1517_ (.Y(_0863_),
    .A(\neurotransmitter.gaba_system.gaba[3] ));
 sg13g2_inv_1 _1518_ (.Y(_0864_),
    .A(\neurotransmitter.gaba_system.gaba[4] ));
 sg13g2_inv_1 _1519_ (.Y(_0865_),
    .A(spi_sck));
 sg13g2_inv_1 _1520_ (.Y(_0866_),
    .A(\neurotransmitter.norepinephrine_system.norepinephrine[3] ));
 sg13g2_inv_1 _1521_ (.Y(_0867_),
    .A(\neurotransmitter.serotonin_system.serotonin[0] ));
 sg13g2_inv_1 _1522_ (.Y(_0868_),
    .A(net88));
 sg13g2_inv_1 _1523_ (.Y(_0869_),
    .A(\talking.byte_count[3] ));
 sg13g2_inv_1 _1524_ (.Y(_0870_),
    .A(\talking.byte_count[5] ));
 sg13g2_inv_1 _1525_ (.Y(_0871_),
    .A(\vital_energy_sys.vital_energy[2] ));
 sg13g2_inv_1 _1526_ (.Y(_0872_),
    .A(\neurotransmitter.cortisol_system.cortisol[3] ));
 sg13g2_inv_1 _1527_ (.Y(_0873_),
    .A(\neurotransmitter.cortisol_system.cortisol[2] ));
 sg13g2_inv_1 _1528_ (.Y(_0874_),
    .A(\neurotransmitter.cortisol_system.cortisol[4] ));
 sg13g2_inv_1 _1529_ (.Y(_0875_),
    .A(_0010_));
 sg13g2_inv_1 _1530_ (.Y(_0876_),
    .A(_0011_));
 sg13g2_inv_1 _1531_ (.Y(_0877_),
    .A(_0016_));
 sg13g2_inv_1 _1532_ (.Y(_0878_),
    .A(_0019_));
 sg13g2_inv_1 _1533_ (.Y(_0879_),
    .A(_0020_));
 sg13g2_inv_1 _1534_ (.Y(_0880_),
    .A(_0029_));
 sg13g2_inv_1 _1535_ (.Y(_0881_),
    .A(_0032_));
 sg13g2_inv_1 _1536_ (.Y(_0882_),
    .A(\talking.uart_shift_reg[3] ));
 sg13g2_inv_1 _1537_ (.Y(_0883_),
    .A(\talking.spi_shift_reg[1] ));
 sg13g2_inv_1 _1538_ (.Y(_0884_),
    .A(net82));
 sg13g2_inv_1 _1539_ (.Y(_0885_),
    .A(\talking.uart_shift_reg[5] ));
 sg13g2_inv_1 _1540_ (.Y(_0886_),
    .A(net105));
 sg13g2_inv_1 _1541_ (.Y(_0887_),
    .A(net100));
 sg13g2_inv_1 _1542_ (.Y(_0888_),
    .A(net84));
 sg13g2_inv_1 _1543_ (.Y(_0889_),
    .A(net90));
 sg13g2_inv_1 _1544_ (.Y(_0890_),
    .A(net57));
 sg13g2_inv_1 _1545_ (.Y(_0891_),
    .A(\heartbeat_divider.counter[3] ));
 sg13g2_inv_1 _1546_ (.Y(_0892_),
    .A(net35));
 sg13g2_inv_1 _1547_ (.Y(_0893_),
    .A(net47));
 sg13g2_nor2_1 _1548_ (.A(net468),
    .B(net467),
    .Y(_0894_));
 sg13g2_or2_2 _1549_ (.X(_0895_),
    .B(net467),
    .A(net468));
 sg13g2_and2_1 _1550_ (.A(\emotions.SER[1] ),
    .B(\emotions.GABA[1] ),
    .X(_0896_));
 sg13g2_nand2_2 _1551_ (.Y(_0897_),
    .A(net498),
    .B(net476));
 sg13g2_nor2_2 _1552_ (.A(net463),
    .B(net462),
    .Y(_0898_));
 sg13g2_nor4_2 _1553_ (.A(\emotions.NE[0] ),
    .B(_0896_),
    .C(_0897_),
    .Y(_0899_),
    .D(_0898_));
 sg13g2_a21oi_1 _1554_ (.A1(\emotions.SER[1] ),
    .A2(_0849_),
    .Y(_0900_),
    .B1(net454));
 sg13g2_nor2_1 _1555_ (.A(net498),
    .B(\emotions.CORT[1] ),
    .Y(_0901_));
 sg13g2_nand2_1 _1556_ (.Y(_0902_),
    .A(net455),
    .B(_0901_));
 sg13g2_nor2_2 _1557_ (.A(_0900_),
    .B(_0902_),
    .Y(_0903_));
 sg13g2_xnor2_1 _1558_ (.Y(_0904_),
    .A(net463),
    .B(net462));
 sg13g2_inv_1 _1559_ (.Y(_0905_),
    .A(_0904_));
 sg13g2_nor4_2 _1560_ (.A(\emotions.DOP[1] ),
    .B(_0896_),
    .C(_0897_),
    .Y(_0906_),
    .D(_0905_));
 sg13g2_nor2_1 _1561_ (.A(_0903_),
    .B(_0906_),
    .Y(_0907_));
 sg13g2_nor3_1 _1562_ (.A(_0899_),
    .B(_0903_),
    .C(_0906_),
    .Y(_0908_));
 sg13g2_nor2_1 _1563_ (.A(_0895_),
    .B(_0908_),
    .Y(_0909_));
 sg13g2_and2_2 _1564_ (.A(\emotions.NE[0] ),
    .B(net497),
    .X(_0910_));
 sg13g2_nand2_2 _1565_ (.Y(_0911_),
    .A(\emotions.NE[0] ),
    .B(net497));
 sg13g2_nor2_2 _1566_ (.A(\nourishment.glucose[6] ),
    .B(net465),
    .Y(_0912_));
 sg13g2_or2_2 _1567_ (.X(_0913_),
    .B(net465),
    .A(\nourishment.glucose[6] ));
 sg13g2_nor4_2 _1568_ (.A(\nourishment.glucose[6] ),
    .B(net465),
    .C(net468),
    .Y(_0914_),
    .D(net467));
 sg13g2_nand2_1 _1569_ (.Y(_0915_),
    .A(net455),
    .B(_0904_));
 sg13g2_or4_2 _1570_ (.A(_0896_),
    .B(_0911_),
    .C(_0914_),
    .D(_0915_),
    .X(_0916_));
 sg13g2_nor2_1 _1571_ (.A(net3),
    .B(net1),
    .Y(_0917_));
 sg13g2_nor3_2 _1572_ (.A(net2),
    .B(net3),
    .C(net1),
    .Y(_0918_));
 sg13g2_nand2b_1 _1573_ (.Y(_0919_),
    .B(net454),
    .A_N(_0918_));
 sg13g2_or3_1 _1574_ (.A(net466),
    .B(net468),
    .C(net467),
    .X(_0920_));
 sg13g2_nand4_1 _1575_ (.B(_0916_),
    .C(_0919_),
    .A(_0913_),
    .Y(_0921_),
    .D(_0920_));
 sg13g2_nor3_1 _1576_ (.A(_0848_),
    .B(\development_stage_sys.dev_stage_reg.cry ),
    .C(net474),
    .Y(_0922_));
 sg13g2_o21ai_1 _1577_ (.B1(_0922_),
    .Y(_0923_),
    .A1(_0909_),
    .A2(_0921_));
 sg13g2_nor3_1 _1578_ (.A(net482),
    .B(\emotions.GABA[1] ),
    .C(\emotions.DOP[1] ),
    .Y(_0924_));
 sg13g2_nor4_2 _1579_ (.A(net498),
    .B(net462),
    .C(_0848_),
    .Y(_0925_),
    .D(_0924_));
 sg13g2_nor4_2 _1580_ (.A(net462),
    .B(\emotions.GABA[1] ),
    .C(_0849_),
    .Y(_0926_),
    .D(_0897_));
 sg13g2_nor2_1 _1581_ (.A(_0925_),
    .B(_0926_),
    .Y(_0927_));
 sg13g2_or2_2 _1582_ (.X(_0928_),
    .B(_0926_),
    .A(_0925_));
 sg13g2_o21ai_1 _1583_ (.B1(_0895_),
    .Y(_0929_),
    .A1(_0903_),
    .A2(_0928_));
 sg13g2_nor4_2 _1584_ (.A(_0848_),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.babble ),
    .C(_0917_),
    .Y(_0930_),
    .D(_0929_));
 sg13g2_nand2_1 _1585_ (.Y(_0931_),
    .A(net477),
    .B(net2));
 sg13g2_nor3_1 _1586_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.play ),
    .B(_0929_),
    .C(_0931_),
    .Y(_0932_));
 sg13g2_nor2_1 _1587_ (.A(_0930_),
    .B(_0932_),
    .Y(_0933_));
 sg13g2_and2_1 _1588_ (.A(_0923_),
    .B(_0933_),
    .X(_0934_));
 sg13g2_nor2_1 _1589_ (.A(\development_stage_sys.dev_stage_reg.cry ),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.idle ),
    .Y(_0935_));
 sg13g2_or2_2 _1590_ (.X(_0936_),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.idle ),
    .A(\development_stage_sys.dev_stage_reg.cry ));
 sg13g2_nor2_1 _1591_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.play ),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.babble ),
    .Y(_0937_));
 sg13g2_nor3_2 _1592_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.play ),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.kick_legs ),
    .C(_0936_),
    .Y(_0938_));
 sg13g2_nor2b_1 _1593_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.babble ),
    .B_N(_0938_),
    .Y(_0939_));
 sg13g2_nor2_1 _1594_ (.A(net480),
    .B(net475),
    .Y(_0940_));
 sg13g2_nand3_1 _1595_ (.B(_0939_),
    .C(_0940_),
    .A(\neurotransmitter.cortisol_system.cortisol_regulator.smile ),
    .Y(_0941_));
 sg13g2_o21ai_1 _1596_ (.B1(net466),
    .Y(_0942_),
    .A1(net468),
    .A2(net467));
 sg13g2_nand2_2 _1597_ (.Y(_0943_),
    .A(\actions.vital_energy_level[0] ),
    .B(\actions.vital_energy_level[1] ));
 sg13g2_nor2b_1 _1598_ (.A(net481),
    .B_N(net474),
    .Y(_0944_));
 sg13g2_nand2_2 _1599_ (.Y(_0945_),
    .A(net455),
    .B(net475));
 sg13g2_nand2b_1 _1600_ (.Y(_0946_),
    .B(_0937_),
    .A_N(\neurotransmitter.cortisol_system.cortisol_regulator.smile ));
 sg13g2_nor4_2 _1601_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.kick_legs ),
    .B(_0936_),
    .C(_0945_),
    .Y(_0947_),
    .D(_0946_));
 sg13g2_nand2b_1 _1602_ (.Y(_0948_),
    .B(_0947_),
    .A_N(_0943_));
 sg13g2_o21ai_1 _1603_ (.B1(_0948_),
    .Y(_0949_),
    .A1(_0941_),
    .A2(_0942_));
 sg13g2_nand2_1 _1604_ (.Y(_0086_),
    .A(_0934_),
    .B(_0949_));
 sg13g2_nor2_1 _1605_ (.A(\counter_.count[2] ),
    .B(_0861_),
    .Y(_0950_));
 sg13g2_nand2b_1 _1606_ (.Y(_0951_),
    .B(\counter_.count[0] ),
    .A_N(\counter_.count[1] ));
 sg13g2_nor3_2 _1607_ (.A(\counter_.count[2] ),
    .B(_0861_),
    .C(_0951_),
    .Y(_0049_));
 sg13g2_nor2_1 _1608_ (.A(net500),
    .B(net501),
    .Y(_0952_));
 sg13g2_nor2b_1 _1609_ (.A(\talking.state[1] ),
    .B_N(_0048_),
    .Y(_0953_));
 sg13g2_nand2_1 _1610_ (.Y(_0954_),
    .A(_0048_),
    .B(_0952_));
 sg13g2_inv_1 _1611_ (.Y(spi_cs),
    .A(_0954_));
 sg13g2_nor2_1 _1612_ (.A(net7),
    .B(net9),
    .Y(_0955_));
 sg13g2_nor3_2 _1613_ (.A(net10),
    .B(net7),
    .C(net9),
    .Y(_0956_));
 sg13g2_nand4_1 _1614_ (.B(_0913_),
    .C(_0918_),
    .A(_0901_),
    .Y(_0957_),
    .D(_0956_));
 sg13g2_nor2_2 _1615_ (.A(\vital_energy_sys.vital_energy[1] ),
    .B(\vital_energy_sys.vital_energy[0] ),
    .Y(_0958_));
 sg13g2_nor2_2 _1616_ (.A(\vital_energy_sys.vital_energy[3] ),
    .B(\vital_energy_sys.vital_energy[2] ),
    .Y(_0959_));
 sg13g2_nor4_2 _1617_ (.A(\vital_energy_sys.vital_energy[3] ),
    .B(\vital_energy_sys.vital_energy[2] ),
    .C(\vital_energy_sys.vital_energy[5] ),
    .Y(_0960_),
    .D(\vital_energy_sys.vital_energy[4] ));
 sg13g2_nand2_2 _1618_ (.Y(_0961_),
    .A(_0958_),
    .B(_0960_));
 sg13g2_nand2_1 _1619_ (.Y(_0962_),
    .A(net456),
    .B(_0894_));
 sg13g2_a21oi_2 _1620_ (.B1(_0962_),
    .Y(_0963_),
    .A2(_0961_),
    .A1(_0957_));
 sg13g2_nand2b_1 _1621_ (.Y(_0964_),
    .B(_0908_),
    .A_N(_0925_));
 sg13g2_nor3_1 _1622_ (.A(net466),
    .B(_0848_),
    .C(net474),
    .Y(_0965_));
 sg13g2_nand3_1 _1623_ (.B(_0964_),
    .C(_0965_),
    .A(net5),
    .Y(_0966_));
 sg13g2_nand2b_1 _1624_ (.Y(_0967_),
    .B(_0943_),
    .A_N(_0957_));
 sg13g2_nand3_1 _1625_ (.B(_0895_),
    .C(_0967_),
    .A(net480),
    .Y(_0968_));
 sg13g2_nand2_1 _1626_ (.Y(_0969_),
    .A(net480),
    .B(_0939_));
 sg13g2_nor3_1 _1627_ (.A(net474),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.smile ),
    .C(_0969_),
    .Y(_0970_));
 sg13g2_nand4_1 _1628_ (.B(_0966_),
    .C(_0968_),
    .A(_0923_),
    .Y(_0971_),
    .D(_0970_));
 sg13g2_nand2b_1 _1629_ (.Y(\actions.next_action[0] ),
    .B(_0971_),
    .A_N(_0963_));
 sg13g2_nor2_2 _1630_ (.A(_0848_),
    .B(_0895_),
    .Y(_0972_));
 sg13g2_nand2_1 _1631_ (.Y(_0973_),
    .A(net477),
    .B(net454));
 sg13g2_nor3_2 _1632_ (.A(_0843_),
    .B(_0844_),
    .C(_0913_),
    .Y(_0974_));
 sg13g2_nor2_2 _1633_ (.A(net482),
    .B(\emotions.SER[0] ),
    .Y(_0975_));
 sg13g2_and4_1 _1634_ (.A(_0910_),
    .B(_0972_),
    .C(_0974_),
    .D(_0975_),
    .X(_0976_));
 sg13g2_nand4_1 _1635_ (.B(_0972_),
    .C(_0974_),
    .A(_0910_),
    .Y(_0977_),
    .D(_0975_));
 sg13g2_nand4_1 _1636_ (.B(_0943_),
    .C(_0947_),
    .A(_0933_),
    .Y(_0978_),
    .D(_0977_));
 sg13g2_nand2b_1 _1637_ (.Y(_0979_),
    .B(_0968_),
    .A_N(_0963_));
 sg13g2_a21oi_1 _1638_ (.A1(_0966_),
    .A2(_0978_),
    .Y(\actions.next_action[1] ),
    .B1(_0979_));
 sg13g2_nor3_1 _1639_ (.A(net481),
    .B(net474),
    .C(\neurotransmitter.cortisol_system.cortisol_regulator.smile ),
    .Y(_0980_));
 sg13g2_nand2b_1 _1640_ (.Y(_0981_),
    .B(_0940_),
    .A_N(\neurotransmitter.cortisol_system.cortisol_regulator.smile ));
 sg13g2_nor3_1 _1641_ (.A(_0858_),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.kick_legs ),
    .C(_0936_),
    .Y(_0982_));
 sg13g2_nand3b_1 _1642_ (.B(_0980_),
    .C(_0982_),
    .Y(_0983_),
    .A_N(\neurotransmitter.cortisol_system.cortisol_regulator.babble ));
 sg13g2_nor2_1 _1643_ (.A(net454),
    .B(_0983_),
    .Y(_0984_));
 sg13g2_a21oi_1 _1644_ (.A1(_0923_),
    .A2(_0984_),
    .Y(_0985_),
    .B1(_0932_));
 sg13g2_nand2b_1 _1645_ (.Y(_0986_),
    .B(_0966_),
    .A_N(_0979_));
 sg13g2_nor3_1 _1646_ (.A(_0930_),
    .B(_0985_),
    .C(_0986_),
    .Y(\actions.next_action[2] ));
 sg13g2_nand3_1 _1647_ (.B(_0938_),
    .C(_0980_),
    .A(\neurotransmitter.cortisol_system.cortisol_regulator.babble ),
    .Y(_0987_));
 sg13g2_nor3_1 _1648_ (.A(_0932_),
    .B(_0942_),
    .C(_0987_),
    .Y(_0988_));
 sg13g2_a21oi_1 _1649_ (.A1(_0923_),
    .A2(_0988_),
    .Y(_0989_),
    .B1(_0930_));
 sg13g2_nor2_1 _1650_ (.A(_0986_),
    .B(_0989_),
    .Y(\actions.next_action[4] ));
 sg13g2_nand2_1 _1651_ (.Y(_0990_),
    .A(_0934_),
    .B(_0966_));
 sg13g2_nand2_1 _1652_ (.Y(_0991_),
    .A(_0941_),
    .B(_0987_));
 sg13g2_nand2_1 _1653_ (.Y(_0992_),
    .A(_0942_),
    .B(_0991_));
 sg13g2_and2_1 _1654_ (.A(_0937_),
    .B(_0980_),
    .X(_0993_));
 sg13g2_nand3_1 _1655_ (.B(_0935_),
    .C(_0993_),
    .A(\neurotransmitter.cortisol_system.cortisol_regulator.kick_legs ),
    .Y(_0994_));
 sg13g2_and2_1 _1656_ (.A(_0992_),
    .B(_0994_),
    .X(_0995_));
 sg13g2_nor3_1 _1657_ (.A(_0963_),
    .B(_0990_),
    .C(_0995_),
    .Y(\actions.next_action[5] ));
 sg13g2_nor2_1 _1658_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.idle ),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.kick_legs ),
    .Y(_0996_));
 sg13g2_nand3_1 _1659_ (.B(_0993_),
    .C(_0996_),
    .A(\development_stage_sys.dev_stage_reg.cry ),
    .Y(_0997_));
 sg13g2_nand3_1 _1660_ (.B(_0994_),
    .C(_0997_),
    .A(_0983_),
    .Y(_0998_));
 sg13g2_nor4_1 _1661_ (.A(_0947_),
    .B(_0970_),
    .C(_0991_),
    .D(_0998_),
    .Y(_0999_));
 sg13g2_nor2_1 _1662_ (.A(_0895_),
    .B(_0983_),
    .Y(_1000_));
 sg13g2_nand3_1 _1663_ (.B(net4),
    .C(_0972_),
    .A(net466),
    .Y(_1001_));
 sg13g2_o21ai_1 _1664_ (.B1(_0977_),
    .Y(_1002_),
    .A1(_0997_),
    .A2(_1001_));
 sg13g2_or3_1 _1665_ (.A(_0999_),
    .B(_1000_),
    .C(_1002_),
    .X(_1003_));
 sg13g2_nand3_1 _1666_ (.B(_0966_),
    .C(_1003_),
    .A(_0934_),
    .Y(_1004_));
 sg13g2_a21oi_1 _1667_ (.A1(_0968_),
    .A2(_1004_),
    .Y(\actions.next_action[6] ),
    .B1(_0963_));
 sg13g2_nand3b_1 _1668_ (.B(_1001_),
    .C(_0977_),
    .Y(_1005_),
    .A_N(_0997_));
 sg13g2_a21oi_1 _1669_ (.A1(_0923_),
    .A2(_1005_),
    .Y(_1006_),
    .B1(_0986_));
 sg13g2_and2_1 _1670_ (.A(_0933_),
    .B(_1006_),
    .X(\actions.next_action[7] ));
 sg13g2_nor2b_1 _1671_ (.A(\counter_.count[0] ),
    .B_N(\counter_.count[1] ),
    .Y(_1007_));
 sg13g2_nand2b_1 _1672_ (.Y(_1008_),
    .B(\counter_.count[1] ),
    .A_N(\counter_.count[0] ));
 sg13g2_a21oi_1 _1673_ (.A1(\counter_.count[1] ),
    .A2(_0950_),
    .Y(_0000_),
    .B1(\counter_.count[0] ));
 sg13g2_o21ai_1 _1674_ (.B1(_0951_),
    .Y(_0001_),
    .A1(_0950_),
    .A2(_1008_));
 sg13g2_nand3_1 _1675_ (.B(\counter_.count[1] ),
    .C(\counter_.count[2] ),
    .A(\counter_.count[0] ),
    .Y(_1009_));
 sg13g2_a21o_1 _1676_ (.A2(\counter_.count[1] ),
    .A1(\counter_.count[0] ),
    .B1(\counter_.count[2] ),
    .X(_1010_));
 sg13g2_and2_1 _1677_ (.A(_1009_),
    .B(_1010_),
    .X(_0002_));
 sg13g2_xnor2_1 _1678_ (.Y(_1011_),
    .A(_0861_),
    .B(_1009_));
 sg13g2_a21oi_1 _1679_ (.A1(_0950_),
    .A2(_1007_),
    .Y(_0003_),
    .B1(_1011_));
 sg13g2_nand2b_1 _1680_ (.Y(\talking.uart_tx ),
    .B(\talking.uart_active ),
    .A_N(\talking.uart_shift_reg[0] ));
 sg13g2_xor2_1 _1681_ (.B(net61),
    .A(\heartbeat_divider.counter[1] ),
    .X(_0057_));
 sg13g2_nand3_1 _1682_ (.B(net61),
    .C(net123),
    .A(\heartbeat_divider.counter[1] ),
    .Y(_1012_));
 sg13g2_a21o_1 _1683_ (.A2(net61),
    .A1(\heartbeat_divider.counter[1] ),
    .B1(net123),
    .X(_1013_));
 sg13g2_and2_1 _1684_ (.A(_1012_),
    .B(net124),
    .X(_0058_));
 sg13g2_nor2_1 _1685_ (.A(_0891_),
    .B(_1012_),
    .Y(_1014_));
 sg13g2_xnor2_1 _1686_ (.Y(_0059_),
    .A(net52),
    .B(_1012_));
 sg13g2_and2_1 _1687_ (.A(net31),
    .B(_1014_),
    .X(_1015_));
 sg13g2_xor2_1 _1688_ (.B(_1014_),
    .A(net31),
    .X(_0060_));
 sg13g2_xor2_1 _1689_ (.B(_1015_),
    .A(net70),
    .X(_0061_));
 sg13g2_nand3_1 _1690_ (.B(net121),
    .C(_1015_),
    .A(net70),
    .Y(_1016_));
 sg13g2_a21o_1 _1691_ (.A2(_1015_),
    .A1(net70),
    .B1(net121),
    .X(_1017_));
 sg13g2_and2_1 _1692_ (.A(_1016_),
    .B(_1017_),
    .X(_0062_));
 sg13g2_nor2_1 _1693_ (.A(_0892_),
    .B(_1016_),
    .Y(_1018_));
 sg13g2_xnor2_1 _1694_ (.Y(_0063_),
    .A(net35),
    .B(_1016_));
 sg13g2_xor2_1 _1695_ (.B(_1018_),
    .A(net49),
    .X(_0064_));
 sg13g2_nand3_1 _1696_ (.B(net122),
    .C(_1018_),
    .A(net49),
    .Y(_1019_));
 sg13g2_a21o_1 _1697_ (.A2(_1018_),
    .A1(net49),
    .B1(net122),
    .X(_1020_));
 sg13g2_and2_1 _1698_ (.A(_1019_),
    .B(_1020_),
    .X(_0065_));
 sg13g2_nor2_1 _1699_ (.A(_0893_),
    .B(_1019_),
    .Y(_1021_));
 sg13g2_xnor2_1 _1700_ (.Y(_0053_),
    .A(net47),
    .B(_1019_));
 sg13g2_xor2_1 _1701_ (.B(_1021_),
    .A(net66),
    .X(_0054_));
 sg13g2_nand3_1 _1702_ (.B(net103),
    .C(_1021_),
    .A(net66),
    .Y(_1022_));
 sg13g2_a21o_1 _1703_ (.A2(_1021_),
    .A1(net66),
    .B1(net103),
    .X(_1023_));
 sg13g2_and2_1 _1704_ (.A(_1022_),
    .B(_1023_),
    .X(_0055_));
 sg13g2_xnor2_1 _1705_ (.Y(_0056_),
    .A(net504),
    .B(net104));
 sg13g2_nor2b_1 _1706_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.GABA[1] ),
    .B_N(net476),
    .Y(_1024_));
 sg13g2_nor3_1 _1707_ (.A(net474),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.SER[1] ),
    .C(\neurotransmitter.cortisol_system.cortisol_regulator.smile ),
    .Y(_1025_));
 sg13g2_nand3_1 _1708_ (.B(_1024_),
    .C(_1025_),
    .A(_0937_),
    .Y(_1026_));
 sg13g2_nor2_2 _1709_ (.A(net3),
    .B(net4),
    .Y(_1027_));
 sg13g2_nand2_2 _1710_ (.Y(_1028_),
    .A(net476),
    .B(_1027_));
 sg13g2_nor2_1 _1711_ (.A(_1026_),
    .B(_1028_),
    .Y(_1029_));
 sg13g2_nand3b_1 _1712_ (.B(_0918_),
    .C(_0956_),
    .Y(_1030_),
    .A_N(net4));
 sg13g2_and2_1 _1713_ (.A(net477),
    .B(_0942_),
    .X(_1031_));
 sg13g2_nor3_1 _1714_ (.A(net10),
    .B(net2),
    .C(net9),
    .Y(_1032_));
 sg13g2_nand2_1 _1715_ (.Y(_1033_),
    .A(_0917_),
    .B(_1032_));
 sg13g2_a221oi_1 _1716_ (.B2(_1033_),
    .C1(net7),
    .B1(_1031_),
    .A1(net481),
    .Y(_1034_),
    .A2(_1030_));
 sg13g2_nor2_1 _1717_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.kick_legs ),
    .B(_0942_),
    .Y(_1035_));
 sg13g2_and2_1 _1718_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.DOP[0] ),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.DOP[1] ),
    .X(_1036_));
 sg13g2_nor2_2 _1719_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.GABA[0] ),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.GABA[1] ),
    .Y(_1037_));
 sg13g2_nor4_1 _1720_ (.A(\development_stage_sys.dev_stage_reg.cry ),
    .B(net473),
    .C(_1036_),
    .D(_1037_),
    .Y(_1038_));
 sg13g2_a21o_1 _1721_ (.A2(_1038_),
    .A1(_1035_),
    .B1(_1026_),
    .X(_1039_));
 sg13g2_o21ai_1 _1722_ (.B1(_1039_),
    .Y(_1040_),
    .A1(_1028_),
    .A2(_1034_));
 sg13g2_nor2_1 _1723_ (.A(_1029_),
    .B(_1040_),
    .Y(_1041_));
 sg13g2_nand2b_1 _1724_ (.Y(_1042_),
    .B(_1040_),
    .A_N(_1029_));
 sg13g2_nor3_1 _1725_ (.A(_1028_),
    .B(_1034_),
    .C(_1039_),
    .Y(_1043_));
 sg13g2_a21oi_2 _1726_ (.B1(_1043_),
    .Y(_1044_),
    .A2(_1028_),
    .A1(_1026_));
 sg13g2_a21o_1 _1727_ (.A2(_1028_),
    .A1(_1026_),
    .B1(_1043_),
    .X(_1045_));
 sg13g2_nor2_1 _1728_ (.A(\emotions.NE[0] ),
    .B(net496),
    .Y(_1046_));
 sg13g2_nor2_2 _1729_ (.A(\neurotransmitter.norepinephrine_system.norepinephrine[1] ),
    .B(\neurotransmitter.norepinephrine_system.norepinephrine[0] ),
    .Y(_1047_));
 sg13g2_or2_2 _1730_ (.X(_1048_),
    .B(\neurotransmitter.norepinephrine_system.norepinephrine[0] ),
    .A(\neurotransmitter.norepinephrine_system.norepinephrine[1] ));
 sg13g2_nor2_1 _1731_ (.A(net499),
    .B(_1048_),
    .Y(_1049_));
 sg13g2_nand2_1 _1732_ (.Y(_1050_),
    .A(_0866_),
    .B(_1049_));
 sg13g2_nor4_2 _1733_ (.A(\emotions.NE[0] ),
    .B(net496),
    .C(\neurotransmitter.norepinephrine_system.norepinephrine[3] ),
    .Y(_1051_),
    .D(net499));
 sg13g2_and2_1 _1734_ (.A(_1047_),
    .B(_1051_),
    .X(_1052_));
 sg13g2_and2_1 _1735_ (.A(\neurotransmitter.norepinephrine_system.norepinephrine[1] ),
    .B(\neurotransmitter.norepinephrine_system.norepinephrine[0] ),
    .X(_1053_));
 sg13g2_nand2_1 _1736_ (.Y(_1054_),
    .A(\neurotransmitter.norepinephrine_system.norepinephrine[1] ),
    .B(\neurotransmitter.norepinephrine_system.norepinephrine[0] ));
 sg13g2_nand3_1 _1737_ (.B(\neurotransmitter.norepinephrine_system.norepinephrine[2] ),
    .C(_1053_),
    .A(\neurotransmitter.norepinephrine_system.norepinephrine[3] ),
    .Y(_1055_));
 sg13g2_nand3_1 _1738_ (.B(net499),
    .C(_0910_),
    .A(\neurotransmitter.norepinephrine_system.norepinephrine[3] ),
    .Y(_1056_));
 sg13g2_nor2_1 _1739_ (.A(_0911_),
    .B(_1055_),
    .Y(_1057_));
 sg13g2_a22oi_1 _1740_ (.Y(_1058_),
    .B1(_1057_),
    .B2(_1029_),
    .A2(_1052_),
    .A1(net434));
 sg13g2_o21ai_1 _1741_ (.B1(_1042_),
    .Y(_1059_),
    .A1(_1045_),
    .A2(_1058_));
 sg13g2_nand3_1 _1742_ (.B(\neurotransmitter.norepinephrine_system.norepinephrine[2] ),
    .C(_1048_),
    .A(\neurotransmitter.norepinephrine_system.norepinephrine[3] ),
    .Y(_1060_));
 sg13g2_nor2_1 _1743_ (.A(_0911_),
    .B(_1060_),
    .Y(_1061_));
 sg13g2_o21ai_1 _1744_ (.B1(net432),
    .Y(_1062_),
    .A1(net434),
    .A2(_1061_));
 sg13g2_o21ai_1 _1745_ (.B1(net433),
    .Y(_1063_),
    .A1(\neurotransmitter.norepinephrine_system.norepinephrine[0] ),
    .A2(_1051_));
 sg13g2_nor2_1 _1746_ (.A(_1044_),
    .B(_1063_),
    .Y(_1064_));
 sg13g2_a21oi_1 _1747_ (.A1(_0876_),
    .A2(_1062_),
    .Y(_1065_),
    .B1(_1064_));
 sg13g2_mux2_1 _1748_ (.A0(_1065_),
    .A1(\neurotransmitter.norepinephrine_system.norepinephrine[0] ),
    .S(net416),
    .X(_0087_));
 sg13g2_nor4_1 _1749_ (.A(_1044_),
    .B(_1047_),
    .C(_1051_),
    .D(_1053_),
    .Y(_1066_));
 sg13g2_o21ai_1 _1750_ (.B1(_1044_),
    .Y(_1067_),
    .A1(_1047_),
    .A2(_1053_));
 sg13g2_nor2b_1 _1751_ (.A(_1066_),
    .B_N(_1067_),
    .Y(_1068_));
 sg13g2_nand4_1 _1752_ (.B(_1048_),
    .C(_1054_),
    .A(net432),
    .Y(_1069_),
    .D(_1056_));
 sg13g2_a21oi_1 _1753_ (.A1(_1067_),
    .A2(_1069_),
    .Y(_1070_),
    .B1(net433));
 sg13g2_a21oi_1 _1754_ (.A1(net433),
    .A2(_1068_),
    .Y(_1071_),
    .B1(_1070_));
 sg13g2_mux2_1 _1755_ (.A0(_1071_),
    .A1(\neurotransmitter.norepinephrine_system.norepinephrine[1] ),
    .S(net416),
    .X(_0088_));
 sg13g2_xnor2_1 _1756_ (.Y(_1072_),
    .A(net499),
    .B(_1054_));
 sg13g2_nand2_1 _1757_ (.Y(_1073_),
    .A(_1044_),
    .B(_1072_));
 sg13g2_a21oi_1 _1758_ (.A1(_1048_),
    .A2(_1056_),
    .Y(_1074_),
    .B1(_0012_));
 sg13g2_a21o_1 _1759_ (.A2(_1048_),
    .A1(_0012_),
    .B1(_1074_),
    .X(_1075_));
 sg13g2_a21oi_1 _1760_ (.A1(net432),
    .A2(_1075_),
    .Y(_1076_),
    .B1(net433));
 sg13g2_nand2_1 _1761_ (.Y(_1077_),
    .A(_1073_),
    .B(_1076_));
 sg13g2_nor3_1 _1762_ (.A(_1044_),
    .B(_1051_),
    .C(_1072_),
    .Y(_1078_));
 sg13g2_xnor2_1 _1763_ (.Y(_1079_),
    .A(net499),
    .B(_1047_));
 sg13g2_o21ai_1 _1764_ (.B1(net433),
    .Y(_1080_),
    .A1(net432),
    .A2(_1079_));
 sg13g2_o21ai_1 _1765_ (.B1(_1077_),
    .Y(_1081_),
    .A1(_1078_),
    .A2(_1080_));
 sg13g2_nand2_1 _1766_ (.Y(_1082_),
    .A(net499),
    .B(net416));
 sg13g2_o21ai_1 _1767_ (.B1(_1082_),
    .Y(_0089_),
    .A1(net416),
    .A2(_1081_));
 sg13g2_nor2_1 _1768_ (.A(_0012_),
    .B(_1054_),
    .Y(_1083_));
 sg13g2_mux2_1 _1769_ (.A0(_1083_),
    .A1(_1049_),
    .S(net433),
    .X(_1084_));
 sg13g2_xnor2_1 _1770_ (.Y(_1085_),
    .A(_0866_),
    .B(_1084_));
 sg13g2_a21o_1 _1771_ (.A2(_1048_),
    .A1(net499),
    .B1(\neurotransmitter.norepinephrine_system.norepinephrine[3] ),
    .X(_1086_));
 sg13g2_nand3_1 _1772_ (.B(_1060_),
    .C(_1086_),
    .A(net432),
    .Y(_1087_));
 sg13g2_nand2_1 _1773_ (.Y(_1088_),
    .A(_1062_),
    .B(_1087_));
 sg13g2_o21ai_1 _1774_ (.B1(\neurotransmitter.norepinephrine_system.norepinephrine[3] ),
    .Y(_1089_),
    .A1(\neurotransmitter.norepinephrine_system.norepinephrine[2] ),
    .A2(_1053_));
 sg13g2_or3_1 _1775_ (.A(\neurotransmitter.norepinephrine_system.norepinephrine[3] ),
    .B(net499),
    .C(_1053_),
    .X(_1090_));
 sg13g2_or2_1 _1776_ (.X(_1091_),
    .B(_1090_),
    .A(_1046_));
 sg13g2_nand3_1 _1777_ (.B(_1089_),
    .C(_1091_),
    .A(net434),
    .Y(_1092_));
 sg13g2_a221oi_1 _1778_ (.B2(_1092_),
    .C1(_1059_),
    .B1(_1088_),
    .A1(_1044_),
    .Y(_1093_),
    .A2(_1085_));
 sg13g2_a21oi_1 _1779_ (.A1(_0866_),
    .A2(net416),
    .Y(_0090_),
    .B1(_1093_));
 sg13g2_mux2_1 _1780_ (.A0(_1055_),
    .A1(_1050_),
    .S(net433),
    .X(_1094_));
 sg13g2_a21oi_1 _1781_ (.A1(_0842_),
    .A2(_1094_),
    .Y(_1095_),
    .B1(net432));
 sg13g2_o21ai_1 _1782_ (.B1(_1095_),
    .Y(_1096_),
    .A1(_0842_),
    .A2(_1094_));
 sg13g2_nand2_1 _1783_ (.Y(_1097_),
    .A(_0013_),
    .B(_1091_));
 sg13g2_o21ai_1 _1784_ (.B1(_1097_),
    .Y(_1098_),
    .A1(_0013_),
    .A2(_1090_));
 sg13g2_nand2b_1 _1785_ (.Y(_1099_),
    .B(_0842_),
    .A_N(_1060_));
 sg13g2_o21ai_1 _1786_ (.B1(\emotions.NE[0] ),
    .Y(_1100_),
    .A1(net495),
    .A2(_1060_));
 sg13g2_nand2_1 _1787_ (.Y(_1101_),
    .A(_1099_),
    .B(_1100_));
 sg13g2_o21ai_1 _1788_ (.B1(net432),
    .Y(_1102_),
    .A1(net434),
    .A2(_1101_));
 sg13g2_a21oi_1 _1789_ (.A1(net434),
    .A2(_1098_),
    .Y(_1103_),
    .B1(_1102_));
 sg13g2_nor2_1 _1790_ (.A(_1059_),
    .B(_1103_),
    .Y(_1104_));
 sg13g2_a22oi_1 _1791_ (.Y(_0091_),
    .B1(_1096_),
    .B2(_1104_),
    .A2(net416),
    .A1(_0842_));
 sg13g2_a21oi_1 _1792_ (.A1(net495),
    .A2(_1050_),
    .Y(_1105_),
    .B1(_1052_));
 sg13g2_nand2b_1 _1793_ (.Y(_1106_),
    .B(net495),
    .A_N(_0013_));
 sg13g2_nand2b_1 _1794_ (.Y(_1107_),
    .B(_0013_),
    .A_N(net495));
 sg13g2_a21oi_1 _1795_ (.A1(_1106_),
    .A2(_1107_),
    .Y(_1108_),
    .B1(_1091_));
 sg13g2_a21oi_1 _1796_ (.A1(net495),
    .A2(_1090_),
    .Y(_1109_),
    .B1(_1108_));
 sg13g2_nand3_1 _1797_ (.B(_1044_),
    .C(_1105_),
    .A(_0911_),
    .Y(_1110_));
 sg13g2_nand2_1 _1798_ (.Y(_1111_),
    .A(_1045_),
    .B(_1109_));
 sg13g2_nand3_1 _1799_ (.B(_1110_),
    .C(_1111_),
    .A(net434),
    .Y(_1112_));
 sg13g2_mux2_1 _1800_ (.A0(_1106_),
    .A1(net495),
    .S(_1055_),
    .X(_1113_));
 sg13g2_o21ai_1 _1801_ (.B1(net496),
    .Y(_1114_),
    .A1(_0013_),
    .A2(_1099_));
 sg13g2_o21ai_1 _1802_ (.B1(_1114_),
    .Y(_1115_),
    .A1(net495),
    .A2(_1060_));
 sg13g2_nor2_1 _1803_ (.A(_1044_),
    .B(_1115_),
    .Y(_1116_));
 sg13g2_o21ai_1 _1804_ (.B1(_1107_),
    .Y(_1117_),
    .A1(net432),
    .A2(_1113_));
 sg13g2_or3_1 _1805_ (.A(net433),
    .B(_1116_),
    .C(_1117_),
    .X(_1118_));
 sg13g2_a21oi_1 _1806_ (.A1(_1112_),
    .A2(_1118_),
    .Y(_1119_),
    .B1(net416));
 sg13g2_a21o_1 _1807_ (.A2(net416),
    .A1(net495),
    .B1(_1119_),
    .X(_0092_));
 sg13g2_nand2_1 _1808_ (.Y(_1120_),
    .A(\neurotransmitter.cortisol_system.cortisol_regulator.SER[0] ),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.SER[1] ));
 sg13g2_or2_1 _1809_ (.X(_1121_),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.CORT[1] ),
    .A(\neurotransmitter.cortisol_system.cortisol_regulator.CORT[0] ));
 sg13g2_or2_1 _1810_ (.X(_1122_),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.NE[1] ),
    .A(\neurotransmitter.cortisol_system.cortisol_regulator.NE[0] ));
 sg13g2_nand4_1 _1811_ (.B(_1120_),
    .C(_1121_),
    .A(_0895_),
    .Y(_1123_),
    .D(_1122_));
 sg13g2_nor2b_1 _1812_ (.A(net1),
    .B_N(_0956_),
    .Y(_1124_));
 sg13g2_or4_2 _1813_ (.A(net10),
    .B(net7),
    .C(net9),
    .D(net1),
    .X(_1125_));
 sg13g2_nor2_1 _1814_ (.A(net8),
    .B(net4),
    .Y(_1126_));
 sg13g2_nor2_1 _1815_ (.A(_1125_),
    .B(_1126_),
    .Y(_1127_));
 sg13g2_or2_1 _1816_ (.X(_1128_),
    .B(_1126_),
    .A(_1125_));
 sg13g2_o21ai_1 _1817_ (.B1(_1127_),
    .Y(_1129_),
    .A1(_0981_),
    .A2(_1123_));
 sg13g2_and2_2 _1818_ (.A(\neurotransmitter.gaba_system.gaba[1] ),
    .B(\neurotransmitter.gaba_system.gaba[0] ),
    .X(_1130_));
 sg13g2_nand2_1 _1819_ (.Y(_1131_),
    .A(\neurotransmitter.gaba_system.gaba[1] ),
    .B(\neurotransmitter.gaba_system.gaba[0] ));
 sg13g2_nand3_1 _1820_ (.B(net494),
    .C(_1130_),
    .A(\neurotransmitter.gaba_system.gaba[3] ),
    .Y(_1132_));
 sg13g2_nand2_1 _1821_ (.Y(_1133_),
    .A(\emotions.GABA[0] ),
    .B(\neurotransmitter.gaba_system.gaba[4] ));
 sg13g2_nor2_1 _1822_ (.A(_1132_),
    .B(_1133_),
    .Y(_1134_));
 sg13g2_and3_1 _1823_ (.X(_1135_),
    .A(\emotions.GABA[1] ),
    .B(_1129_),
    .C(_1134_));
 sg13g2_or2_1 _1824_ (.X(_1136_),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.NE[1] ),
    .A(net473));
 sg13g2_nor2_1 _1825_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.SER[0] ),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.SER[1] ),
    .Y(_1137_));
 sg13g2_nor4_2 _1826_ (.A(_0847_),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.CORT[1] ),
    .C(_1136_),
    .Y(_1138_),
    .D(_1137_));
 sg13g2_a21oi_2 _1827_ (.B1(net480),
    .Y(_1139_),
    .A2(_1138_),
    .A1(_0938_));
 sg13g2_nor3_1 _1828_ (.A(_1125_),
    .B(_1135_),
    .C(_1139_),
    .Y(_1140_));
 sg13g2_nor3_1 _1829_ (.A(_0981_),
    .B(_1123_),
    .C(_1124_),
    .Y(_1141_));
 sg13g2_a21o_1 _1830_ (.A2(_1139_),
    .A1(_1128_),
    .B1(_1141_),
    .X(_1142_));
 sg13g2_a21oi_2 _1831_ (.B1(_1141_),
    .Y(_1143_),
    .A2(_1139_),
    .A1(_1128_));
 sg13g2_or2_1 _1832_ (.X(_1144_),
    .B(\emotions.GABA[1] ),
    .A(\emotions.GABA[0] ));
 sg13g2_o21ai_1 _1833_ (.B1(_1144_),
    .Y(_1145_),
    .A1(_1140_),
    .A2(net449));
 sg13g2_nand2_1 _1834_ (.Y(_1146_),
    .A(_1125_),
    .B(_1139_));
 sg13g2_mux2_1 _1835_ (.A0(_1129_),
    .A1(_1124_),
    .S(_1139_),
    .X(_1147_));
 sg13g2_o21ai_1 _1836_ (.B1(_1146_),
    .Y(_1148_),
    .A1(_1129_),
    .A2(_1139_));
 sg13g2_nor2_2 _1837_ (.A(net494),
    .B(_1130_),
    .Y(_1149_));
 sg13g2_nor3_1 _1838_ (.A(\emotions.GABA[0] ),
    .B(\neurotransmitter.gaba_system.gaba[3] ),
    .C(\neurotransmitter.gaba_system.gaba[4] ),
    .Y(_1150_));
 sg13g2_nand2_1 _1839_ (.Y(_1151_),
    .A(_1149_),
    .B(_1150_));
 sg13g2_nor2_2 _1840_ (.A(\neurotransmitter.gaba_system.gaba[1] ),
    .B(\neurotransmitter.gaba_system.gaba[0] ),
    .Y(_1152_));
 sg13g2_or2_1 _1841_ (.X(_1153_),
    .B(\neurotransmitter.gaba_system.gaba[0] ),
    .A(\neurotransmitter.gaba_system.gaba[1] ));
 sg13g2_nand2b_1 _1842_ (.Y(_1154_),
    .B(_1152_),
    .A_N(net494));
 sg13g2_nor4_1 _1843_ (.A(\emotions.GABA[0] ),
    .B(\neurotransmitter.gaba_system.gaba[3] ),
    .C(\neurotransmitter.gaba_system.gaba[4] ),
    .D(_1154_),
    .Y(_1155_));
 sg13g2_xnor2_1 _1844_ (.Y(_1156_),
    .A(_0845_),
    .B(_1155_));
 sg13g2_o21ai_1 _1845_ (.B1(_1156_),
    .Y(_1157_),
    .A1(net448),
    .A2(_1151_));
 sg13g2_nand2_1 _1846_ (.Y(_1158_),
    .A(net449),
    .B(_1157_));
 sg13g2_nand2_1 _1847_ (.Y(_1159_),
    .A(net494),
    .B(_1153_));
 sg13g2_nand3_1 _1848_ (.B(net494),
    .C(_1153_),
    .A(\neurotransmitter.gaba_system.gaba[3] ),
    .Y(_1160_));
 sg13g2_nor2_1 _1849_ (.A(_1133_),
    .B(_1160_),
    .Y(_1161_));
 sg13g2_inv_1 _1850_ (.Y(_1162_),
    .A(_1161_));
 sg13g2_xnor2_1 _1851_ (.Y(_1163_),
    .A(_0845_),
    .B(_1134_));
 sg13g2_o21ai_1 _1852_ (.B1(_1140_),
    .Y(_1164_),
    .A1(net448),
    .A2(_1162_));
 sg13g2_o21ai_1 _1853_ (.B1(_1158_),
    .Y(_1165_),
    .A1(_1163_),
    .A2(_1164_));
 sg13g2_nor2b_2 _1854_ (.A(_1165_),
    .B_N(_1145_),
    .Y(_1166_));
 sg13g2_a21oi_2 _1855_ (.B1(net449),
    .Y(_1167_),
    .A2(_1161_),
    .A1(\emotions.GABA[1] ));
 sg13g2_nor2_1 _1856_ (.A(net448),
    .B(_1167_),
    .Y(_1168_));
 sg13g2_nor2_1 _1857_ (.A(_0014_),
    .B(_1168_),
    .Y(_1169_));
 sg13g2_and2_1 _1858_ (.A(_0845_),
    .B(_1150_),
    .X(_1170_));
 sg13g2_nand2b_1 _1859_ (.Y(_1171_),
    .B(_1170_),
    .A_N(net494));
 sg13g2_a21oi_1 _1860_ (.A1(_0862_),
    .A2(_1171_),
    .Y(_1172_),
    .B1(net447));
 sg13g2_a21oi_1 _1861_ (.A1(_1142_),
    .A2(_1172_),
    .Y(_1173_),
    .B1(_1169_));
 sg13g2_mux2_1 _1862_ (.A0(_1173_),
    .A1(\neurotransmitter.gaba_system.gaba[0] ),
    .S(_1166_),
    .X(_0093_));
 sg13g2_a21oi_1 _1863_ (.A1(_1131_),
    .A2(_1153_),
    .Y(_1174_),
    .B1(_1148_));
 sg13g2_o21ai_1 _1864_ (.B1(net447),
    .Y(_1175_),
    .A1(_1130_),
    .A2(_1152_));
 sg13g2_nor3_1 _1865_ (.A(_1130_),
    .B(net447),
    .C(_1152_),
    .Y(_1176_));
 sg13g2_a21oi_1 _1866_ (.A1(_1171_),
    .A2(_1176_),
    .Y(_1177_),
    .B1(_1174_));
 sg13g2_o21ai_1 _1867_ (.B1(_1176_),
    .Y(_1178_),
    .A1(_0845_),
    .A2(_1162_));
 sg13g2_nand3_1 _1868_ (.B(_1175_),
    .C(_1178_),
    .A(_1143_),
    .Y(_1179_));
 sg13g2_o21ai_1 _1869_ (.B1(_1179_),
    .Y(_1180_),
    .A1(_1143_),
    .A2(_1177_));
 sg13g2_mux2_1 _1870_ (.A0(_1180_),
    .A1(\neurotransmitter.gaba_system.gaba[1] ),
    .S(_1166_),
    .X(_0094_));
 sg13g2_and2_1 _1871_ (.A(net449),
    .B(_1154_),
    .X(_1181_));
 sg13g2_xnor2_1 _1872_ (.Y(_1182_),
    .A(\neurotransmitter.gaba_system.gaba[2] ),
    .B(_1130_));
 sg13g2_a22oi_1 _1873_ (.Y(_1183_),
    .B1(_1182_),
    .B2(_1143_),
    .A2(_1181_),
    .A1(_1159_));
 sg13g2_xnor2_1 _1874_ (.Y(_1184_),
    .A(_0015_),
    .B(_1152_));
 sg13g2_nand2_2 _1875_ (.Y(_1185_),
    .A(_1149_),
    .B(_1170_));
 sg13g2_nand2_1 _1876_ (.Y(_1186_),
    .A(_1182_),
    .B(_1185_));
 sg13g2_a221oi_1 _1877_ (.B2(net449),
    .C1(net447),
    .B1(_1186_),
    .A1(_1167_),
    .Y(_1187_),
    .A2(_1184_));
 sg13g2_a21o_1 _1878_ (.A2(_1183_),
    .A1(net447),
    .B1(_1187_),
    .X(_1188_));
 sg13g2_mux2_1 _1879_ (.A0(_1188_),
    .A1(net494),
    .S(_1166_),
    .X(_0095_));
 sg13g2_o21ai_1 _1880_ (.B1(_1143_),
    .Y(_1189_),
    .A1(_0015_),
    .A2(_1131_));
 sg13g2_nor2b_1 _1881_ (.A(_1181_),
    .B_N(_1189_),
    .Y(_1190_));
 sg13g2_xnor2_1 _1882_ (.Y(_1191_),
    .A(_0863_),
    .B(_1190_));
 sg13g2_nor2_1 _1883_ (.A(_0863_),
    .B(_1149_),
    .Y(_1192_));
 sg13g2_nor3_2 _1884_ (.A(\neurotransmitter.gaba_system.gaba[3] ),
    .B(net494),
    .C(_1130_),
    .Y(_1193_));
 sg13g2_o21ai_1 _1885_ (.B1(_1185_),
    .Y(_1194_),
    .A1(_1192_),
    .A2(_1193_));
 sg13g2_xnor2_1 _1886_ (.Y(_1195_),
    .A(_0863_),
    .B(_1159_));
 sg13g2_a221oi_1 _1887_ (.B2(_1167_),
    .C1(net448),
    .B1(_1195_),
    .A1(net449),
    .Y(_1196_),
    .A2(_1194_));
 sg13g2_a21o_1 _1888_ (.A2(_1191_),
    .A1(net448),
    .B1(_1196_),
    .X(_1197_));
 sg13g2_mux2_1 _1889_ (.A0(_1197_),
    .A1(\neurotransmitter.gaba_system.gaba[3] ),
    .S(_1166_),
    .X(_0096_));
 sg13g2_nor2_1 _1890_ (.A(_1132_),
    .B(net449),
    .Y(_1198_));
 sg13g2_nor3_2 _1891_ (.A(\neurotransmitter.gaba_system.gaba[3] ),
    .B(_1143_),
    .C(_1154_),
    .Y(_1199_));
 sg13g2_o21ai_1 _1892_ (.B1(\neurotransmitter.gaba_system.gaba[4] ),
    .Y(_1200_),
    .A1(_1198_),
    .A2(_1199_));
 sg13g2_or3_1 _1893_ (.A(\neurotransmitter.gaba_system.gaba[4] ),
    .B(_1198_),
    .C(_1199_),
    .X(_1201_));
 sg13g2_nand3_1 _1894_ (.B(_1200_),
    .C(_1201_),
    .A(net447),
    .Y(_1202_));
 sg13g2_nand2_1 _1895_ (.Y(_1203_),
    .A(_0016_),
    .B(_1193_));
 sg13g2_xnor2_1 _1896_ (.Y(_1204_),
    .A(_0016_),
    .B(_1193_));
 sg13g2_a21oi_1 _1897_ (.A1(_1185_),
    .A2(_1204_),
    .Y(_1205_),
    .B1(_1143_));
 sg13g2_xnor2_1 _1898_ (.Y(_1206_),
    .A(\neurotransmitter.gaba_system.gaba[4] ),
    .B(_1160_));
 sg13g2_a21oi_1 _1899_ (.A1(_1148_),
    .A2(_1206_),
    .Y(_1207_),
    .B1(_1168_));
 sg13g2_o21ai_1 _1900_ (.B1(_1202_),
    .Y(_1208_),
    .A1(_1205_),
    .A2(_1207_));
 sg13g2_mux2_1 _1901_ (.A0(_1208_),
    .A1(\neurotransmitter.gaba_system.gaba[4] ),
    .S(_1166_),
    .X(_0097_));
 sg13g2_a22oi_1 _1902_ (.Y(_1209_),
    .B1(_1199_),
    .B2(_0864_),
    .A2(_1198_),
    .A1(_0877_));
 sg13g2_xnor2_1 _1903_ (.Y(_1210_),
    .A(\emotions.GABA[0] ),
    .B(_1209_));
 sg13g2_xnor2_1 _1904_ (.Y(_1211_),
    .A(\emotions.GABA[0] ),
    .B(_1203_));
 sg13g2_nand2_1 _1905_ (.Y(_1212_),
    .A(_1185_),
    .B(_1211_));
 sg13g2_nor2_1 _1906_ (.A(_0016_),
    .B(_1160_),
    .Y(_1213_));
 sg13g2_xnor2_1 _1907_ (.Y(_1214_),
    .A(\emotions.GABA[0] ),
    .B(_1213_));
 sg13g2_a221oi_1 _1908_ (.B2(_1167_),
    .C1(net447),
    .B1(_1214_),
    .A1(net449),
    .Y(_1215_),
    .A2(_1212_));
 sg13g2_a21oi_1 _1909_ (.A1(net447),
    .A2(_1210_),
    .Y(_1216_),
    .B1(_1215_));
 sg13g2_mux2_1 _1910_ (.A0(_1216_),
    .A1(_0066_),
    .S(_1166_),
    .X(_0098_));
 sg13g2_a21o_1 _1911_ (.A2(_1145_),
    .A1(_0067_),
    .B1(_1165_),
    .X(_0099_));
 sg13g2_nor3_1 _1912_ (.A(net10),
    .B(net2),
    .C(net3),
    .Y(_1217_));
 sg13g2_o21ai_1 _1913_ (.B1(_0955_),
    .Y(_1218_),
    .A1(net454),
    .A2(_1217_));
 sg13g2_and2_1 _1914_ (.A(net477),
    .B(_1218_),
    .X(_1219_));
 sg13g2_a21oi_1 _1915_ (.A1(_0857_),
    .A2(_1120_),
    .Y(_1220_),
    .B1(_1036_));
 sg13g2_nand2_1 _1916_ (.Y(_1221_),
    .A(\neurotransmitter.cortisol_system.cortisol_regulator.CORT[1] ),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.NE[1] ));
 sg13g2_or4_1 _1917_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.play ),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.kick_legs ),
    .C(_0942_),
    .D(_1221_),
    .X(_1222_));
 sg13g2_o21ai_1 _1918_ (.B1(net455),
    .Y(_1223_),
    .A1(_1220_),
    .A2(_1222_));
 sg13g2_nor2_1 _1919_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.DOP[0] ),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.DOP[1] ),
    .Y(_1224_));
 sg13g2_nor3_1 _1920_ (.A(_0936_),
    .B(_1037_),
    .C(_1137_),
    .Y(_1225_));
 sg13g2_and2_1 _1921_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.CORT[0] ),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.CORT[1] ),
    .X(_1226_));
 sg13g2_a22oi_1 _1922_ (.Y(_1227_),
    .B1(\neurotransmitter.cortisol_system.cortisol_regulator.NE[0] ),
    .B2(\neurotransmitter.cortisol_system.cortisol_regulator.NE[1] ),
    .A2(\neurotransmitter.cortisol_system.cortisol_regulator.CORT[1] ),
    .A1(\neurotransmitter.cortisol_system.cortisol_regulator.CORT[0] ));
 sg13g2_and4_1 _1923_ (.A(net476),
    .B(_0913_),
    .C(_0920_),
    .D(_1227_),
    .X(_1228_));
 sg13g2_o21ai_1 _1924_ (.B1(_1228_),
    .Y(_1229_),
    .A1(_1224_),
    .A2(_1225_));
 sg13g2_nand2_2 _1925_ (.Y(_1230_),
    .A(_1219_),
    .B(_1229_));
 sg13g2_nor2_1 _1926_ (.A(net6),
    .B(net10),
    .Y(_1231_));
 sg13g2_o21ai_1 _1927_ (.B1(_1231_),
    .Y(_1232_),
    .A1(net454),
    .A2(_1217_));
 sg13g2_nand2_1 _1928_ (.Y(_1233_),
    .A(net455),
    .B(_1232_));
 sg13g2_a221oi_1 _1929_ (.B2(_1233_),
    .C1(_1226_),
    .B1(_1229_),
    .A1(_1219_),
    .Y(_1234_),
    .A2(_1223_));
 sg13g2_and2_1 _1930_ (.A(_1230_),
    .B(_1234_),
    .X(_1235_));
 sg13g2_nand2_2 _1931_ (.Y(_1236_),
    .A(_1230_),
    .B(_1234_));
 sg13g2_nand2_2 _1932_ (.Y(_1237_),
    .A(\neurotransmitter.dopamine_system.dopamine[1] ),
    .B(\neurotransmitter.dopamine_system.dopamine[0] ));
 sg13g2_and4_1 _1933_ (.A(\neurotransmitter.dopamine_system.dopamine[1] ),
    .B(\neurotransmitter.dopamine_system.dopamine[0] ),
    .C(\neurotransmitter.dopamine_system.dopamine[3] ),
    .D(net493),
    .X(_1238_));
 sg13g2_nand3_1 _1934_ (.B(\neurotransmitter.dopamine_system.dopamine[4] ),
    .C(_1238_),
    .A(net490),
    .Y(_1239_));
 sg13g2_nor2_1 _1935_ (.A(_0849_),
    .B(_1239_),
    .Y(_1240_));
 sg13g2_xnor2_1 _1936_ (.Y(_1241_),
    .A(_0849_),
    .B(_1239_));
 sg13g2_or4_2 _1937_ (.A(_1218_),
    .B(_1223_),
    .C(_1229_),
    .D(_1231_),
    .X(_1242_));
 sg13g2_nand2_1 _1938_ (.Y(_1243_),
    .A(_1230_),
    .B(_1242_));
 sg13g2_nor2_2 _1939_ (.A(\neurotransmitter.dopamine_system.dopamine[1] ),
    .B(\neurotransmitter.dopamine_system.dopamine[0] ),
    .Y(_1244_));
 sg13g2_or2_2 _1940_ (.X(_1245_),
    .B(\neurotransmitter.dopamine_system.dopamine[0] ),
    .A(\neurotransmitter.dopamine_system.dopamine[1] ));
 sg13g2_nand3_1 _1941_ (.B(net493),
    .C(_1245_),
    .A(\neurotransmitter.dopamine_system.dopamine[3] ),
    .Y(_1246_));
 sg13g2_inv_1 _1942_ (.Y(_1247_),
    .A(_1246_));
 sg13g2_nand4_1 _1943_ (.B(net492),
    .C(net429),
    .A(net491),
    .Y(_1248_),
    .D(_1247_));
 sg13g2_a21oi_1 _1944_ (.A1(_1241_),
    .A2(_1248_),
    .Y(_1249_),
    .B1(_1236_));
 sg13g2_nand2b_1 _1945_ (.Y(_1250_),
    .B(_1237_),
    .A_N(net493));
 sg13g2_nor2_2 _1946_ (.A(\neurotransmitter.dopamine_system.dopamine[3] ),
    .B(net493),
    .Y(_1251_));
 sg13g2_nand2_2 _1947_ (.Y(_1252_),
    .A(_1237_),
    .B(_1251_));
 sg13g2_nor3_1 _1948_ (.A(net490),
    .B(net492),
    .C(_1252_),
    .Y(_1253_));
 sg13g2_or3_1 _1949_ (.A(_1218_),
    .B(_1229_),
    .C(_1240_),
    .X(_1254_));
 sg13g2_nand3_1 _1950_ (.B(_1242_),
    .C(_1254_),
    .A(net431),
    .Y(_1255_));
 sg13g2_nor2_1 _1951_ (.A(net493),
    .B(_1245_),
    .Y(_1256_));
 sg13g2_nand2_1 _1952_ (.Y(_1257_),
    .A(_1244_),
    .B(_1251_));
 sg13g2_nor3_1 _1953_ (.A(net490),
    .B(\neurotransmitter.dopamine_system.dopamine[4] ),
    .C(_1257_),
    .Y(_1258_));
 sg13g2_xnor2_1 _1954_ (.Y(_1259_),
    .A(_0849_),
    .B(_1258_));
 sg13g2_nand2_1 _1955_ (.Y(_1260_),
    .A(_1236_),
    .B(_1259_));
 sg13g2_a22oi_1 _1956_ (.Y(_1261_),
    .B1(_1255_),
    .B2(_1260_),
    .A2(_1253_),
    .A1(net430));
 sg13g2_nor3_1 _1957_ (.A(\emotions.DOP[1] ),
    .B(net490),
    .C(net492),
    .Y(_1262_));
 sg13g2_nand2_2 _1958_ (.Y(_1263_),
    .A(_1251_),
    .B(_1262_));
 sg13g2_nand2_1 _1959_ (.Y(_1264_),
    .A(_1255_),
    .B(_1263_));
 sg13g2_o21ai_1 _1960_ (.B1(_1264_),
    .Y(_1265_),
    .A1(_1249_),
    .A2(_1261_));
 sg13g2_nand4_1 _1961_ (.B(net490),
    .C(net492),
    .A(\emotions.DOP[1] ),
    .Y(_1266_),
    .D(_1247_));
 sg13g2_nand2_1 _1962_ (.Y(_1267_),
    .A(net431),
    .B(_1266_));
 sg13g2_a21oi_1 _1963_ (.A1(net430),
    .A2(_1267_),
    .Y(_1268_),
    .B1(_0017_));
 sg13g2_a21oi_1 _1964_ (.A1(_0859_),
    .A2(_1263_),
    .Y(_1269_),
    .B1(_1235_));
 sg13g2_a21oi_1 _1965_ (.A1(net429),
    .A2(_1269_),
    .Y(_1270_),
    .B1(_1268_));
 sg13g2_mux2_1 _1966_ (.A0(\neurotransmitter.dopamine_system.dopamine[0] ),
    .A1(_1270_),
    .S(_1265_),
    .X(_0100_));
 sg13g2_nand4_1 _1967_ (.B(net430),
    .C(_1245_),
    .A(_1237_),
    .Y(_1271_),
    .D(_1266_));
 sg13g2_a21o_1 _1968_ (.A2(_1245_),
    .A1(_1237_),
    .B1(net430),
    .X(_1272_));
 sg13g2_nand4_1 _1969_ (.B(net430),
    .C(_1245_),
    .A(_1237_),
    .Y(_1273_),
    .D(_1263_));
 sg13g2_nand2_1 _1970_ (.Y(_1274_),
    .A(_1271_),
    .B(_1272_));
 sg13g2_and2_1 _1971_ (.A(_1236_),
    .B(_1272_),
    .X(_1275_));
 sg13g2_a22oi_1 _1972_ (.Y(_1276_),
    .B1(_1275_),
    .B2(_1273_),
    .A2(_1274_),
    .A1(net431));
 sg13g2_mux2_1 _1973_ (.A0(\neurotransmitter.dopamine_system.dopamine[1] ),
    .A1(_1276_),
    .S(_1265_),
    .X(_0101_));
 sg13g2_xnor2_1 _1974_ (.Y(_1277_),
    .A(net493),
    .B(_1244_));
 sg13g2_xor2_1 _1975_ (.B(_1237_),
    .A(\neurotransmitter.dopamine_system.dopamine[2] ),
    .X(_1278_));
 sg13g2_nand2_1 _1976_ (.Y(_1279_),
    .A(_1263_),
    .B(_1278_));
 sg13g2_mux2_1 _1977_ (.A0(_1277_),
    .A1(_1279_),
    .S(net430),
    .X(_1280_));
 sg13g2_xnor2_1 _1978_ (.Y(_1281_),
    .A(_0018_),
    .B(_1244_));
 sg13g2_nand3_1 _1979_ (.B(_1266_),
    .C(_1281_),
    .A(net430),
    .Y(_1282_));
 sg13g2_nand3_1 _1980_ (.B(_1242_),
    .C(_1278_),
    .A(_1230_),
    .Y(_1283_));
 sg13g2_nand3_1 _1981_ (.B(_1282_),
    .C(_1283_),
    .A(_1235_),
    .Y(_1284_));
 sg13g2_o21ai_1 _1982_ (.B1(_1284_),
    .Y(_1285_),
    .A1(net431),
    .A2(_1280_));
 sg13g2_mux2_1 _1983_ (.A0(net493),
    .A1(_1285_),
    .S(_1265_),
    .X(_0102_));
 sg13g2_nor2_1 _1984_ (.A(_0018_),
    .B(_1237_),
    .Y(_1286_));
 sg13g2_mux2_1 _1985_ (.A0(_1256_),
    .A1(_1286_),
    .S(net431),
    .X(_1287_));
 sg13g2_nor2_1 _1986_ (.A(\neurotransmitter.dopamine_system.dopamine[3] ),
    .B(_1287_),
    .Y(_1288_));
 sg13g2_a21o_1 _1987_ (.A2(_1287_),
    .A1(\neurotransmitter.dopamine_system.dopamine[3] ),
    .B1(net429),
    .X(_1289_));
 sg13g2_nor2_1 _1988_ (.A(_1252_),
    .B(_1262_),
    .Y(_1290_));
 sg13g2_a21oi_1 _1989_ (.A1(\neurotransmitter.dopamine_system.dopamine[3] ),
    .A2(_1250_),
    .Y(_1291_),
    .B1(_1290_));
 sg13g2_nand2_1 _1990_ (.Y(_1292_),
    .A(_1236_),
    .B(_1291_));
 sg13g2_a21oi_1 _1991_ (.A1(net493),
    .A2(_1245_),
    .Y(_1293_),
    .B1(\neurotransmitter.dopamine_system.dopamine[3] ));
 sg13g2_or2_1 _1992_ (.X(_1294_),
    .B(_1293_),
    .A(_1247_));
 sg13g2_nand3_1 _1993_ (.B(_1266_),
    .C(_1294_),
    .A(net431),
    .Y(_1295_));
 sg13g2_nand3_1 _1994_ (.B(_1292_),
    .C(_1295_),
    .A(net429),
    .Y(_1296_));
 sg13g2_o21ai_1 _1995_ (.B1(_1296_),
    .Y(_1297_),
    .A1(_1288_),
    .A2(_1289_));
 sg13g2_mux2_1 _1996_ (.A0(\neurotransmitter.dopamine_system.dopamine[3] ),
    .A1(_1297_),
    .S(_1265_),
    .X(_0103_));
 sg13g2_a21o_1 _1997_ (.A2(_1234_),
    .A1(_1230_),
    .B1(_1257_),
    .X(_1298_));
 sg13g2_nand3_1 _1998_ (.B(_1234_),
    .C(_1238_),
    .A(_1230_),
    .Y(_1299_));
 sg13g2_nand2_1 _1999_ (.Y(_1300_),
    .A(_1298_),
    .B(_1299_));
 sg13g2_nor2_1 _2000_ (.A(net492),
    .B(_1300_),
    .Y(_1301_));
 sg13g2_a21o_1 _2001_ (.A2(_1300_),
    .A1(net492),
    .B1(net429),
    .X(_1302_));
 sg13g2_nand2_1 _2002_ (.Y(_1303_),
    .A(_0878_),
    .B(_1252_));
 sg13g2_nand2_1 _2003_ (.Y(_1304_),
    .A(_0019_),
    .B(_1290_));
 sg13g2_nand3_1 _2004_ (.B(_1303_),
    .C(_1304_),
    .A(_1236_),
    .Y(_1305_));
 sg13g2_xor2_1 _2005_ (.B(_1246_),
    .A(net492),
    .X(_1306_));
 sg13g2_nand3_1 _2006_ (.B(_1266_),
    .C(_1306_),
    .A(net431),
    .Y(_1307_));
 sg13g2_nand3_1 _2007_ (.B(_1305_),
    .C(_1307_),
    .A(net429),
    .Y(_1308_));
 sg13g2_o21ai_1 _2008_ (.B1(_1308_),
    .Y(_1309_),
    .A1(_1301_),
    .A2(_1302_));
 sg13g2_mux2_1 _2009_ (.A0(net492),
    .A1(_1309_),
    .S(_1265_),
    .X(_0104_));
 sg13g2_nand4_1 _2010_ (.B(_1230_),
    .C(_1234_),
    .A(_0878_),
    .Y(_1310_),
    .D(_1238_));
 sg13g2_o21ai_1 _2011_ (.B1(_1310_),
    .Y(_1311_),
    .A1(\neurotransmitter.dopamine_system.dopamine[4] ),
    .A2(_1298_));
 sg13g2_xnor2_1 _2012_ (.Y(_1312_),
    .A(net490),
    .B(_1311_));
 sg13g2_nor2_1 _2013_ (.A(_0019_),
    .B(_1246_),
    .Y(_1313_));
 sg13g2_xnor2_1 _2014_ (.Y(_1314_),
    .A(net490),
    .B(_1313_));
 sg13g2_nand3_1 _2015_ (.B(_1266_),
    .C(_1314_),
    .A(_1235_),
    .Y(_1315_));
 sg13g2_o21ai_1 _2016_ (.B1(net491),
    .Y(_1316_),
    .A1(_0878_),
    .A2(_1252_));
 sg13g2_o21ai_1 _2017_ (.B1(_1316_),
    .Y(_1317_),
    .A1(net491),
    .A2(_1304_));
 sg13g2_o21ai_1 _2018_ (.B1(net429),
    .Y(_1318_),
    .A1(net431),
    .A2(_1317_));
 sg13g2_nand2b_1 _2019_ (.Y(_1319_),
    .B(_1315_),
    .A_N(_1318_));
 sg13g2_o21ai_1 _2020_ (.B1(_1319_),
    .Y(_1320_),
    .A1(net429),
    .A2(_1312_));
 sg13g2_mux2_1 _2021_ (.A0(net490),
    .A1(_1320_),
    .S(_1265_),
    .X(_0105_));
 sg13g2_nand2_1 _2022_ (.Y(_1321_),
    .A(_0068_),
    .B(_1264_));
 sg13g2_o21ai_1 _2023_ (.B1(_1321_),
    .Y(_0106_),
    .A1(_1249_),
    .A2(_1261_));
 sg13g2_nand2_1 _2024_ (.Y(_1322_),
    .A(\nourishment.glucose[3] ),
    .B(\nourishment.glucose[2] ));
 sg13g2_and4_1 _2025_ (.A(\nourishment.glucose[3] ),
    .B(\nourishment.glucose[2] ),
    .C(\nourishment.glucose[5] ),
    .D(\nourishment.glucose[4] ),
    .X(_1323_));
 sg13g2_nand3_1 _2026_ (.B(net465),
    .C(_1323_),
    .A(\nourishment.glucose[6] ),
    .Y(_1324_));
 sg13g2_nand2_1 _2027_ (.Y(_1325_),
    .A(net453),
    .B(_1324_));
 sg13g2_inv_1 _2028_ (.Y(_1326_),
    .A(_1325_));
 sg13g2_nor2_1 _2029_ (.A(\nourishment.glucose[1] ),
    .B(\nourishment.glucose[0] ),
    .Y(_1327_));
 sg13g2_nor3_2 _2030_ (.A(\nourishment.glucose[1] ),
    .B(\nourishment.glucose[0] ),
    .C(\nourishment.glucose[2] ),
    .Y(_1328_));
 sg13g2_nand2b_2 _2031_ (.Y(_1329_),
    .B(_1328_),
    .A_N(\nourishment.glucose[3] ));
 sg13g2_nor3_2 _2032_ (.A(\nourishment.glucose[5] ),
    .B(\nourishment.glucose[4] ),
    .C(_1329_),
    .Y(_1330_));
 sg13g2_nand2_2 _2033_ (.Y(_1331_),
    .A(_0912_),
    .B(_1330_));
 sg13g2_nand2_2 _2034_ (.Y(_1332_),
    .A(_1325_),
    .B(_1331_));
 sg13g2_nor3_1 _2035_ (.A(_0028_),
    .B(net453),
    .C(_1332_),
    .Y(_1333_));
 sg13g2_a21oi_1 _2036_ (.A1(_0856_),
    .A2(_1332_),
    .Y(_0107_),
    .B1(_1333_));
 sg13g2_o21ai_1 _2037_ (.B1(\nourishment.glucose[1] ),
    .Y(_1334_),
    .A1(\nourishment.glucose[0] ),
    .A2(_1332_));
 sg13g2_nor2_1 _2038_ (.A(net453),
    .B(_1327_),
    .Y(_1335_));
 sg13g2_o21ai_1 _2039_ (.B1(_1334_),
    .Y(_0108_),
    .A1(_1332_),
    .A2(_1335_));
 sg13g2_nor3_1 _2040_ (.A(_0914_),
    .B(_1037_),
    .C(_1136_),
    .Y(_1336_));
 sg13g2_nand2b_1 _2041_ (.Y(_1337_),
    .B(net478),
    .A_N(_1336_));
 sg13g2_o21ai_1 _2042_ (.B1(_0955_),
    .Y(_1338_),
    .A1(_0895_),
    .A2(_0918_));
 sg13g2_a22oi_1 _2043_ (.Y(_1339_),
    .B1(_1338_),
    .B2(net478),
    .A2(\neurotransmitter.cortisol_system.cortisol_regulator.NE[1] ),
    .A1(\neurotransmitter.cortisol_system.cortisol_regulator.NE[0] ));
 sg13g2_nand3_1 _2044_ (.B(_1025_),
    .C(_1122_),
    .A(_1024_),
    .Y(_1340_));
 sg13g2_nor2_1 _2045_ (.A(net481),
    .B(_1027_),
    .Y(_1341_));
 sg13g2_or2_1 _2046_ (.X(_1342_),
    .B(_1341_),
    .A(_1340_));
 sg13g2_nand3_1 _2047_ (.B(_1339_),
    .C(_1342_),
    .A(_1337_),
    .Y(_1343_));
 sg13g2_or2_1 _2048_ (.X(_1344_),
    .B(_1339_),
    .A(_1337_));
 sg13g2_nand2b_1 _2049_ (.Y(_1345_),
    .B(_1338_),
    .A_N(_1340_));
 sg13g2_or2_1 _2050_ (.X(_1346_),
    .B(_1341_),
    .A(_1337_));
 sg13g2_nand3_1 _2051_ (.B(_1345_),
    .C(_1346_),
    .A(_1344_),
    .Y(_1347_));
 sg13g2_nand4_1 _2052_ (.B(_1344_),
    .C(_1345_),
    .A(net446),
    .Y(_1348_),
    .D(_1346_));
 sg13g2_nand4_1 _2053_ (.B(_1339_),
    .C(_1340_),
    .A(_1337_),
    .Y(_1349_),
    .D(_1341_));
 sg13g2_inv_1 _2054_ (.Y(_1350_),
    .A(_1349_));
 sg13g2_and2_1 _2055_ (.A(_1344_),
    .B(_1349_),
    .X(_1351_));
 sg13g2_nand2_1 _2056_ (.Y(_1352_),
    .A(_1344_),
    .B(_1349_));
 sg13g2_and2_2 _2057_ (.A(net464),
    .B(\neurotransmitter.cortisol_system.cortisol[2] ),
    .X(_1353_));
 sg13g2_and3_2 _2058_ (.X(_1354_),
    .A(\neurotransmitter.cortisol_system.cortisol[3] ),
    .B(\neurotransmitter.cortisol_system.cortisol[4] ),
    .C(_1353_));
 sg13g2_nand3b_1 _2059_ (.B(_1354_),
    .C(net463),
    .Y(_1355_),
    .A_N(_0052_));
 sg13g2_nand2_1 _2060_ (.Y(_1356_),
    .A(net488),
    .B(_1353_));
 sg13g2_nand3_1 _2061_ (.B(\neurotransmitter.cortisol_system.cortisol[3] ),
    .C(_1353_),
    .A(net488),
    .Y(_1357_));
 sg13g2_nand3_1 _2062_ (.B(net489),
    .C(_1354_),
    .A(net463),
    .Y(_1358_));
 sg13g2_nor2_1 _2063_ (.A(_0052_),
    .B(_1358_),
    .Y(_1359_));
 sg13g2_or2_2 _2064_ (.X(_1360_),
    .B(\neurotransmitter.cortisol_system.cortisol[2] ),
    .A(net464));
 sg13g2_nor2_2 _2065_ (.A(\neurotransmitter.cortisol_system.cortisol[3] ),
    .B(_1360_),
    .Y(_1361_));
 sg13g2_nand2b_2 _2066_ (.Y(_1362_),
    .B(_1361_),
    .A_N(net488));
 sg13g2_nand3_1 _2067_ (.B(_0874_),
    .C(_0052_),
    .A(_0843_),
    .Y(_1363_));
 sg13g2_nor3_1 _2068_ (.A(net445),
    .B(_1362_),
    .C(_1363_),
    .Y(_1364_));
 sg13g2_a21oi_1 _2069_ (.A1(_1347_),
    .A2(_1359_),
    .Y(_1365_),
    .B1(_1364_));
 sg13g2_o21ai_1 _2070_ (.B1(_1348_),
    .Y(_1366_),
    .A1(net426),
    .A2(_1365_));
 sg13g2_and2_2 _2071_ (.A(_1352_),
    .B(_1355_),
    .X(_1367_));
 sg13g2_a21oi_1 _2072_ (.A1(net464),
    .A2(net489),
    .Y(_1368_),
    .B1(\neurotransmitter.cortisol_system.cortisol[2] ));
 sg13g2_and4_1 _2073_ (.A(_0872_),
    .B(_0874_),
    .C(_0898_),
    .D(_1368_),
    .X(_1369_));
 sg13g2_nand2b_1 _2074_ (.Y(_1370_),
    .B(\neurotransmitter.cortisol_system.cortisol[1] ),
    .A_N(net488));
 sg13g2_o21ai_1 _2075_ (.B1(_1369_),
    .Y(_1371_),
    .A1(_1363_),
    .A2(_1370_));
 sg13g2_a221oi_1 _2076_ (.B2(_1350_),
    .C1(net415),
    .B1(_1371_),
    .A1(net446),
    .Y(_1372_),
    .A2(_1367_));
 sg13g2_a21oi_1 _2077_ (.A1(_0879_),
    .A2(net428),
    .Y(_1373_),
    .B1(_1367_));
 sg13g2_nor3_1 _2078_ (.A(net489),
    .B(net445),
    .C(net426),
    .Y(_1374_));
 sg13g2_a21o_1 _2079_ (.A2(_1373_),
    .A1(net445),
    .B1(_1374_),
    .X(_1375_));
 sg13g2_mux2_1 _2080_ (.A0(net489),
    .A1(_1375_),
    .S(_1372_),
    .X(_0109_));
 sg13g2_nor2b_1 _2081_ (.A(net500),
    .B_N(\talking.state[2] ),
    .Y(_1376_));
 sg13g2_and2_1 _2082_ (.A(net502),
    .B(_1376_),
    .X(_1377_));
 sg13g2_nand2_1 _2083_ (.Y(_1378_),
    .A(net502),
    .B(_1376_));
 sg13g2_nand2_2 _2084_ (.Y(_1379_),
    .A(net500),
    .B(net501));
 sg13g2_inv_1 _2085_ (.Y(_1380_),
    .A(_1379_));
 sg13g2_o21ai_1 _2086_ (.B1(_1378_),
    .Y(_1381_),
    .A1(\talking.state[2] ),
    .A2(_1379_));
 sg13g2_nor2b_2 _2087_ (.A(net502),
    .B_N(_1376_),
    .Y(_1382_));
 sg13g2_nand2_1 _2088_ (.Y(_1383_),
    .A(\talking.state[2] ),
    .B(_0952_));
 sg13g2_nor2_1 _2089_ (.A(\talking.byte_count[4] ),
    .B(\talking.byte_count[3] ),
    .Y(_1384_));
 sg13g2_nor2_1 _2090_ (.A(\talking.byte_count[2] ),
    .B(\talking.byte_count[1] ),
    .Y(_1385_));
 sg13g2_nand3_1 _2091_ (.B(_1384_),
    .C(_1385_),
    .A(_0051_),
    .Y(_1386_));
 sg13g2_and2_1 _2092_ (.A(_1382_),
    .B(_1386_),
    .X(_1387_));
 sg13g2_nand2_2 _2093_ (.Y(_1388_),
    .A(_1382_),
    .B(_1386_));
 sg13g2_or2_1 _2094_ (.X(_1389_),
    .B(_1386_),
    .A(_1383_));
 sg13g2_a21oi_1 _2095_ (.A1(_0870_),
    .A2(\talking.byte_count[0] ),
    .Y(_1390_),
    .B1(_1389_));
 sg13g2_nor2_2 _2096_ (.A(_1387_),
    .B(_1390_),
    .Y(_1391_));
 sg13g2_nand2_1 _2097_ (.Y(_1392_),
    .A(net500),
    .B(_0048_));
 sg13g2_nor2_2 _2098_ (.A(net501),
    .B(_1392_),
    .Y(_1393_));
 sg13g2_or2_1 _2099_ (.X(_1394_),
    .B(_1392_),
    .A(net501));
 sg13g2_nor3_1 _2100_ (.A(net451),
    .B(_1382_),
    .C(_1393_),
    .Y(_1395_));
 sg13g2_nor2_2 _2101_ (.A(\talking.spi_bit_count[3] ),
    .B(net452),
    .Y(_1396_));
 sg13g2_nor2_1 _2102_ (.A(_1395_),
    .B(_1396_),
    .Y(_1397_));
 sg13g2_o21ai_1 _2103_ (.B1(_1393_),
    .Y(_1398_),
    .A1(\talking.skip_address_bytes[0] ),
    .A2(\talking.skip_address_bytes[1] ));
 sg13g2_nand3_1 _2104_ (.B(_1397_),
    .C(_1398_),
    .A(_1391_),
    .Y(_1399_));
 sg13g2_nor2_1 _2105_ (.A(\talking.uart_bit_count[1] ),
    .B(\talking.uart_bit_count[2] ),
    .Y(_1400_));
 sg13g2_and3_1 _2106_ (.X(_1401_),
    .A(\talking.uart_bit_count[0] ),
    .B(\talking.uart_bit_count[3] ),
    .C(_1400_));
 sg13g2_nand3_1 _2107_ (.B(net108),
    .C(_1400_),
    .A(\talking.uart_bit_count[0] ),
    .Y(_1402_));
 sg13g2_o21ai_1 _2108_ (.B1(net115),
    .Y(_1403_),
    .A1(_1399_),
    .A2(_1402_));
 sg13g2_o21ai_1 _2109_ (.B1(net116),
    .Y(_0110_),
    .A1(net451),
    .A2(_1399_));
 sg13g2_nor2b_1 _2110_ (.A(_0956_),
    .B_N(_1031_),
    .Y(_0206_));
 sg13g2_nand3b_1 _2111_ (.B(net477),
    .C(_0942_),
    .Y(_0207_),
    .A_N(_0956_));
 sg13g2_nand2b_1 _2112_ (.Y(_0208_),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.DOP[1] ),
    .A_N(net473));
 sg13g2_nor4_1 _2113_ (.A(_0936_),
    .B(_0942_),
    .C(_1037_),
    .D(_0208_),
    .Y(_0209_));
 sg13g2_o21ai_1 _2114_ (.B1(_1227_),
    .Y(_0210_),
    .A1(_1137_),
    .A2(_0209_));
 sg13g2_nand2_1 _2115_ (.Y(_0211_),
    .A(net476),
    .B(_0210_));
 sg13g2_a21oi_2 _2116_ (.B1(_0206_),
    .Y(_0212_),
    .A2(_0210_),
    .A1(net476));
 sg13g2_and2_1 _2117_ (.A(_0206_),
    .B(_0210_),
    .X(_0213_));
 sg13g2_nand3_1 _2118_ (.B(net4),
    .C(_0207_),
    .A(net455),
    .Y(_0214_));
 sg13g2_and2_1 _2119_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.GABA[0] ),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.GABA[1] ),
    .X(_0215_));
 sg13g2_or3_1 _2120_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.DOP[1] ),
    .B(_1221_),
    .C(_0215_),
    .X(_0216_));
 sg13g2_a21oi_1 _2121_ (.A1(_1120_),
    .A2(_0216_),
    .Y(_0217_),
    .B1(_0946_));
 sg13g2_a21oi_1 _2122_ (.A1(net476),
    .A2(_0217_),
    .Y(_0218_),
    .B1(_0214_));
 sg13g2_a21oi_1 _2123_ (.A1(_0211_),
    .A2(_0218_),
    .Y(_0219_),
    .B1(_0213_));
 sg13g2_a21o_2 _2124_ (.A2(_0218_),
    .A1(_0211_),
    .B1(_0213_),
    .X(_0220_));
 sg13g2_o21ai_1 _2125_ (.B1(_0214_),
    .Y(_0221_),
    .A1(_0207_),
    .A2(_0217_));
 sg13g2_a21oi_2 _2126_ (.B1(_0212_),
    .Y(_0222_),
    .A2(_0221_),
    .A1(net425));
 sg13g2_a21o_2 _2127_ (.A2(_0221_),
    .A1(net425),
    .B1(_0212_),
    .X(_0223_));
 sg13g2_nand2_2 _2128_ (.Y(_0224_),
    .A(\neurotransmitter.serotonin_system.serotonin[1] ),
    .B(\neurotransmitter.serotonin_system.serotonin[0] ));
 sg13g2_and4_2 _2129_ (.A(\neurotransmitter.serotonin_system.serotonin[1] ),
    .B(\neurotransmitter.serotonin_system.serotonin[0] ),
    .C(\neurotransmitter.serotonin_system.serotonin[3] ),
    .D(net487),
    .X(_0225_));
 sg13g2_nand3_1 _2130_ (.B(net485),
    .C(_0225_),
    .A(net483),
    .Y(_0226_));
 sg13g2_nand4_1 _2131_ (.B(net483),
    .C(net485),
    .A(net482),
    .Y(_0227_),
    .D(_0225_));
 sg13g2_o21ai_1 _2132_ (.B1(_0212_),
    .Y(_0228_),
    .A1(_0220_),
    .A2(_0227_));
 sg13g2_a21oi_1 _2133_ (.A1(_0223_),
    .A2(_0228_),
    .Y(_0229_),
    .B1(_0975_));
 sg13g2_nand2b_1 _2134_ (.Y(_0230_),
    .B(_0224_),
    .A_N(net487));
 sg13g2_nor2_2 _2135_ (.A(\neurotransmitter.serotonin_system.serotonin[3] ),
    .B(net487),
    .Y(_0231_));
 sg13g2_nand2_2 _2136_ (.Y(_0232_),
    .A(_0224_),
    .B(_0231_));
 sg13g2_or4_1 _2137_ (.A(net483),
    .B(net485),
    .C(net425),
    .D(_0232_),
    .X(_0233_));
 sg13g2_nor2_2 _2138_ (.A(\neurotransmitter.serotonin_system.serotonin[1] ),
    .B(\neurotransmitter.serotonin_system.serotonin[0] ),
    .Y(_0234_));
 sg13g2_or2_1 _2139_ (.X(_0235_),
    .B(\neurotransmitter.serotonin_system.serotonin[0] ),
    .A(\neurotransmitter.serotonin_system.serotonin[1] ));
 sg13g2_nand2_2 _2140_ (.Y(_0236_),
    .A(_0231_),
    .B(_0234_));
 sg13g2_nor3_1 _2141_ (.A(net483),
    .B(net486),
    .C(_0236_),
    .Y(_0237_));
 sg13g2_xor2_1 _2142_ (.B(_0237_),
    .A(net482),
    .X(_0238_));
 sg13g2_nand3_1 _2143_ (.B(_0233_),
    .C(_0238_),
    .A(_0222_),
    .Y(_0239_));
 sg13g2_and3_2 _2144_ (.X(_0240_),
    .A(\neurotransmitter.serotonin_system.serotonin[3] ),
    .B(net487),
    .C(_0235_));
 sg13g2_nand3_1 _2145_ (.B(net485),
    .C(_0240_),
    .A(net483),
    .Y(_0241_));
 sg13g2_xor2_1 _2146_ (.B(_0226_),
    .A(net482),
    .X(_0242_));
 sg13g2_o21ai_1 _2147_ (.B1(_0242_),
    .Y(_0243_),
    .A1(net425),
    .A2(_0241_));
 sg13g2_o21ai_1 _2148_ (.B1(_0223_),
    .Y(_0244_),
    .A1(_0228_),
    .A2(_0243_));
 sg13g2_nand2_1 _2149_ (.Y(_0245_),
    .A(_0239_),
    .B(_0244_));
 sg13g2_a21oi_2 _2150_ (.B1(_0229_),
    .Y(_0246_),
    .A2(_0244_),
    .A1(_0239_));
 sg13g2_nand4_1 _2151_ (.B(net483),
    .C(net485),
    .A(net482),
    .Y(_0247_),
    .D(_0240_));
 sg13g2_nand2_1 _2152_ (.Y(_0248_),
    .A(_0212_),
    .B(_0247_));
 sg13g2_a21oi_1 _2153_ (.A1(_0220_),
    .A2(_0248_),
    .Y(_0249_),
    .B1(_0008_));
 sg13g2_nor3_1 _2154_ (.A(net482),
    .B(net484),
    .C(net485),
    .Y(_0250_));
 sg13g2_nand2_2 _2155_ (.Y(_0251_),
    .A(_0231_),
    .B(_0250_));
 sg13g2_a21oi_1 _2156_ (.A1(_0867_),
    .A2(_0251_),
    .Y(_0252_),
    .B1(_0212_));
 sg13g2_a21oi_1 _2157_ (.A1(_0220_),
    .A2(_0252_),
    .Y(_0253_),
    .B1(_0249_));
 sg13g2_mux2_1 _2158_ (.A0(_0253_),
    .A1(\neurotransmitter.serotonin_system.serotonin[0] ),
    .S(_0246_),
    .X(_0111_));
 sg13g2_and2_1 _2159_ (.A(_0224_),
    .B(_0235_),
    .X(_0254_));
 sg13g2_and2_2 _2160_ (.A(_0220_),
    .B(_0247_),
    .X(_0255_));
 sg13g2_nand2b_1 _2161_ (.Y(_0256_),
    .B(net425),
    .A_N(_0254_));
 sg13g2_a21oi_1 _2162_ (.A1(_0254_),
    .A2(_0255_),
    .Y(_0257_),
    .B1(_0222_));
 sg13g2_nand3_1 _2163_ (.B(_0251_),
    .C(_0254_),
    .A(_0220_),
    .Y(_0258_));
 sg13g2_a21oi_1 _2164_ (.A1(_0256_),
    .A2(_0258_),
    .Y(_0259_),
    .B1(_0223_));
 sg13g2_a21o_1 _2165_ (.A2(_0257_),
    .A1(_0256_),
    .B1(_0259_),
    .X(_0260_));
 sg13g2_mux2_1 _2166_ (.A0(_0260_),
    .A1(\neurotransmitter.serotonin_system.serotonin[1] ),
    .S(_0246_),
    .X(_0112_));
 sg13g2_xor2_1 _2167_ (.B(_0224_),
    .A(net487),
    .X(_0261_));
 sg13g2_nand3_1 _2168_ (.B(_0251_),
    .C(_0261_),
    .A(_0220_),
    .Y(_0262_));
 sg13g2_xnor2_1 _2169_ (.Y(_0263_),
    .A(net487),
    .B(_0234_));
 sg13g2_o21ai_1 _2170_ (.B1(_0262_),
    .Y(_0264_),
    .A1(_0220_),
    .A2(_0263_));
 sg13g2_xnor2_1 _2171_ (.Y(_0265_),
    .A(_0009_),
    .B(_0234_));
 sg13g2_a22oi_1 _2172_ (.Y(_0266_),
    .B1(_0265_),
    .B2(_0255_),
    .A2(_0261_),
    .A1(net424));
 sg13g2_mux2_1 _2173_ (.A0(_0264_),
    .A1(_0266_),
    .S(_0223_),
    .X(_0267_));
 sg13g2_mux2_1 _2174_ (.A0(_0267_),
    .A1(\neurotransmitter.serotonin_system.serotonin[2] ),
    .S(_0246_),
    .X(_0113_));
 sg13g2_nor2_1 _2175_ (.A(_0232_),
    .B(_0250_),
    .Y(_0268_));
 sg13g2_a21oi_1 _2176_ (.A1(\neurotransmitter.serotonin_system.serotonin[3] ),
    .A2(_0230_),
    .Y(_0269_),
    .B1(_0268_));
 sg13g2_o21ai_1 _2177_ (.B1(\neurotransmitter.serotonin_system.serotonin[3] ),
    .Y(_0270_),
    .A1(net487),
    .A2(_0235_));
 sg13g2_a21o_1 _2178_ (.A2(_0270_),
    .A1(_0236_),
    .B1(_0220_),
    .X(_0271_));
 sg13g2_o21ai_1 _2179_ (.B1(_0271_),
    .Y(_0272_),
    .A1(net425),
    .A2(_0269_));
 sg13g2_a21oi_1 _2180_ (.A1(net487),
    .A2(_0235_),
    .Y(_0273_),
    .B1(\neurotransmitter.serotonin_system.serotonin[3] ));
 sg13g2_or2_1 _2181_ (.X(_0274_),
    .B(_0273_),
    .A(_0240_));
 sg13g2_nor2_1 _2182_ (.A(_0009_),
    .B(_0224_),
    .Y(_0275_));
 sg13g2_xnor2_1 _2183_ (.Y(_0276_),
    .A(\neurotransmitter.serotonin_system.serotonin[3] ),
    .B(_0275_));
 sg13g2_a22oi_1 _2184_ (.Y(_0277_),
    .B1(_0276_),
    .B2(net424),
    .A2(_0274_),
    .A1(_0255_));
 sg13g2_mux2_1 _2185_ (.A0(_0272_),
    .A1(_0277_),
    .S(_0223_),
    .X(_0278_));
 sg13g2_mux2_1 _2186_ (.A0(_0278_),
    .A1(\neurotransmitter.serotonin_system.serotonin[3] ),
    .S(_0246_),
    .X(_0114_));
 sg13g2_xor2_1 _2187_ (.B(_0236_),
    .A(net485),
    .X(_0279_));
 sg13g2_nand2_1 _2188_ (.Y(_0280_),
    .A(_0010_),
    .B(_0268_));
 sg13g2_a21oi_1 _2189_ (.A1(_0875_),
    .A2(_0232_),
    .Y(_0281_),
    .B1(net424));
 sg13g2_a22oi_1 _2190_ (.Y(_0282_),
    .B1(_0280_),
    .B2(_0281_),
    .A2(_0279_),
    .A1(net424));
 sg13g2_xnor2_1 _2191_ (.Y(_0283_),
    .A(net486),
    .B(_0240_));
 sg13g2_xnor2_1 _2192_ (.Y(_0284_),
    .A(net486),
    .B(_0225_));
 sg13g2_a221oi_1 _2193_ (.B2(net424),
    .C1(_0222_),
    .B1(_0284_),
    .A1(_0255_),
    .Y(_0285_),
    .A2(_0283_));
 sg13g2_a21o_1 _2194_ (.A2(_0282_),
    .A1(_0222_),
    .B1(_0285_),
    .X(_0286_));
 sg13g2_mux2_1 _2195_ (.A0(_0286_),
    .A1(net486),
    .S(_0246_),
    .X(_0115_));
 sg13g2_nor2b_1 _2196_ (.A(_0010_),
    .B_N(_0240_),
    .Y(_0287_));
 sg13g2_xnor2_1 _2197_ (.Y(_0288_),
    .A(net484),
    .B(_0287_));
 sg13g2_nor2b_1 _2198_ (.A(_0010_),
    .B_N(_0225_),
    .Y(_0289_));
 sg13g2_xnor2_1 _2199_ (.Y(_0290_),
    .A(net484),
    .B(_0289_));
 sg13g2_a22oi_1 _2200_ (.Y(_0291_),
    .B1(_0290_),
    .B2(net424),
    .A2(_0288_),
    .A1(_0255_));
 sg13g2_xor2_1 _2201_ (.B(_0010_),
    .A(net484),
    .X(_0292_));
 sg13g2_a221oi_1 _2202_ (.B2(_0292_),
    .C1(net424),
    .B1(_0268_),
    .A1(net483),
    .Y(_0293_),
    .A2(_0232_));
 sg13g2_o21ai_1 _2203_ (.B1(net483),
    .Y(_0294_),
    .A1(net485),
    .A2(_0236_));
 sg13g2_nor2b_1 _2204_ (.A(_0237_),
    .B_N(_0294_),
    .Y(_0295_));
 sg13g2_and2_1 _2205_ (.A(net424),
    .B(_0295_),
    .X(_0296_));
 sg13g2_o21ai_1 _2206_ (.B1(_0222_),
    .Y(_0297_),
    .A1(_0293_),
    .A2(_0296_));
 sg13g2_o21ai_1 _2207_ (.B1(_0297_),
    .Y(_0298_),
    .A1(_0222_),
    .A2(_0291_));
 sg13g2_mux2_1 _2208_ (.A0(_0298_),
    .A1(_0069_),
    .S(_0246_),
    .X(_0116_));
 sg13g2_o21ai_1 _2209_ (.B1(_0245_),
    .Y(_0117_),
    .A1(_0840_),
    .A2(_0229_));
 sg13g2_nor2_1 _2210_ (.A(net471),
    .B(\illness_sys.illness[8] ),
    .Y(_0299_));
 sg13g2_a21oi_1 _2211_ (.A1(net470),
    .A2(\illness_sys.illness[8] ),
    .Y(_0300_),
    .B1(\illness_sys.illness[7] ));
 sg13g2_nor2_1 _2212_ (.A(_0299_),
    .B(_0300_),
    .Y(_0118_));
 sg13g2_nor4_2 _2213_ (.A(\emotions.CORT[1] ),
    .B(_0851_),
    .C(net454),
    .Y(_0301_),
    .D(_0912_));
 sg13g2_o21ai_1 _2214_ (.B1(net478),
    .Y(_0302_),
    .A1(_0047_),
    .A2(_0301_));
 sg13g2_nor2_1 _2215_ (.A(_0850_),
    .B(_0302_),
    .Y(_0303_));
 sg13g2_a21o_2 _2216_ (.A2(_0301_),
    .A1(_0850_),
    .B1(_0302_),
    .X(_0304_));
 sg13g2_a21oi_2 _2217_ (.B1(_0302_),
    .Y(_0305_),
    .A2(_0301_),
    .A1(_0850_));
 sg13g2_and2_1 _2218_ (.A(\illness_sys.illness[3] ),
    .B(net461),
    .X(_0306_));
 sg13g2_nand3_1 _2219_ (.B(\illness_sys.illness[5] ),
    .C(_0306_),
    .A(\illness_sys.illness[4] ),
    .Y(_0307_));
 sg13g2_nand2_1 _2220_ (.Y(_0308_),
    .A(\illness_sys.illness[7] ),
    .B(\illness_sys.illness[6] ));
 sg13g2_nor2_1 _2221_ (.A(_0307_),
    .B(_0308_),
    .Y(_0309_));
 sg13g2_and2_2 _2222_ (.A(\illness_sys.illness[1] ),
    .B(\illness_sys.illness[0] ),
    .X(_0310_));
 sg13g2_nand2_2 _2223_ (.Y(_0311_),
    .A(\illness_sys.illness[1] ),
    .B(\illness_sys.illness[0] ));
 sg13g2_nor2_1 _2224_ (.A(net471),
    .B(_0311_),
    .Y(_0312_));
 sg13g2_nand3_1 _2225_ (.B(_0309_),
    .C(_0312_),
    .A(\illness_sys.illness[8] ),
    .Y(_0313_));
 sg13g2_nor2_2 _2226_ (.A(\illness_sys.illness[1] ),
    .B(\illness_sys.illness[0] ),
    .Y(_0314_));
 sg13g2_inv_1 _2227_ (.Y(_0315_),
    .A(_0314_));
 sg13g2_nor2_1 _2228_ (.A(\illness_sys.illness[7] ),
    .B(\illness_sys.illness[6] ),
    .Y(_0316_));
 sg13g2_nor2_1 _2229_ (.A(\illness_sys.illness[4] ),
    .B(\illness_sys.illness[5] ),
    .Y(_0317_));
 sg13g2_nor2_1 _2230_ (.A(\illness_sys.illness[3] ),
    .B(net461),
    .Y(_0318_));
 sg13g2_nor4_2 _2231_ (.A(\illness_sys.illness[4] ),
    .B(\illness_sys.illness[5] ),
    .C(\illness_sys.illness[3] ),
    .Y(_0319_),
    .D(net461));
 sg13g2_nand2_1 _2232_ (.Y(_0320_),
    .A(_0316_),
    .B(_0319_));
 sg13g2_nor2_1 _2233_ (.A(net461),
    .B(_0315_),
    .Y(_0321_));
 sg13g2_nor2b_1 _2234_ (.A(\illness_sys.illness[3] ),
    .B_N(_0321_),
    .Y(_0322_));
 sg13g2_nand2_1 _2235_ (.Y(_0323_),
    .A(_0314_),
    .B(_0319_));
 sg13g2_nor2_1 _2236_ (.A(_0315_),
    .B(_0320_),
    .Y(_0324_));
 sg13g2_nand3b_1 _2237_ (.B(_0324_),
    .C(net471),
    .Y(_0325_),
    .A_N(\illness_sys.illness[8] ));
 sg13g2_a21oi_1 _2238_ (.A1(_0313_),
    .A2(_0325_),
    .Y(_0326_),
    .B1(net443));
 sg13g2_nor3_2 _2239_ (.A(_0006_),
    .B(_0307_),
    .C(_0308_),
    .Y(_0327_));
 sg13g2_or2_1 _2240_ (.X(_0328_),
    .B(_0327_),
    .A(net471));
 sg13g2_nor2_1 _2241_ (.A(\illness_sys.illness[3] ),
    .B(\illness_sys.illness[8] ),
    .Y(_0329_));
 sg13g2_nand2_1 _2242_ (.Y(_0330_),
    .A(net461),
    .B(_0006_));
 sg13g2_nand4_1 _2243_ (.B(_0317_),
    .C(_0329_),
    .A(_0316_),
    .Y(_0331_),
    .D(_0330_));
 sg13g2_a21oi_2 _2244_ (.B1(_0331_),
    .Y(_0332_),
    .A2(_0315_),
    .A1(\illness_sys.illness[2] ));
 sg13g2_o21ai_1 _2245_ (.B1(_0328_),
    .Y(_0333_),
    .A1(_0047_),
    .A2(_0332_));
 sg13g2_a21oi_2 _2246_ (.B1(_0326_),
    .Y(_0334_),
    .A2(_0333_),
    .A1(net442));
 sg13g2_nand3_1 _2247_ (.B(net442),
    .C(_0327_),
    .A(_0850_),
    .Y(_0335_));
 sg13g2_o21ai_1 _2248_ (.B1(_0335_),
    .Y(_0336_),
    .A1(_0881_),
    .A2(net442));
 sg13g2_mux2_1 _2249_ (.A0(\illness_sys.illness[0] ),
    .A1(_0336_),
    .S(_0334_),
    .X(_0119_));
 sg13g2_nor2_1 _2250_ (.A(_0310_),
    .B(_0314_),
    .Y(_0337_));
 sg13g2_xnor2_1 _2251_ (.Y(_0338_),
    .A(net470),
    .B(_0337_));
 sg13g2_o21ai_1 _2252_ (.B1(_0335_),
    .Y(_0339_),
    .A1(net442),
    .A2(_0338_));
 sg13g2_mux2_1 _2253_ (.A0(\illness_sys.illness[1] ),
    .A1(_0339_),
    .S(_0334_),
    .X(_0120_));
 sg13g2_a21o_2 _2254_ (.A2(_0977_),
    .A1(_0916_),
    .B1(_0848_),
    .X(_0340_));
 sg13g2_nor4_2 _2255_ (.A(net473),
    .B(_0851_),
    .C(_0912_),
    .Y(_0341_),
    .D(_0927_));
 sg13g2_nor2_2 _2256_ (.A(_0340_),
    .B(_0341_),
    .Y(_0342_));
 sg13g2_or2_2 _2257_ (.X(_0343_),
    .B(_0341_),
    .A(_0340_));
 sg13g2_nor4_2 _2258_ (.A(net481),
    .B(net473),
    .C(_0912_),
    .Y(_0344_),
    .D(_0927_));
 sg13g2_nand4_1 _2259_ (.B(_0850_),
    .C(_0913_),
    .A(net455),
    .Y(_0345_),
    .D(_0928_));
 sg13g2_nor2_2 _2260_ (.A(net460),
    .B(\development_stage_sys.development_stage_level[2] ),
    .Y(_0346_));
 sg13g2_nor3_1 _2261_ (.A(net460),
    .B(net459),
    .C(\development_stage_sys.development_stage_level[2] ),
    .Y(_0347_));
 sg13g2_nand2_1 _2262_ (.Y(_0348_),
    .A(_0854_),
    .B(_0347_));
 sg13g2_nor3_2 _2263_ (.A(net459),
    .B(\development_stage_sys.development_stage_level[5] ),
    .C(\development_stage_sys.development_stage_level[4] ),
    .Y(_0349_));
 sg13g2_nand2_2 _2264_ (.Y(_0350_),
    .A(_0346_),
    .B(_0349_));
 sg13g2_nor3_2 _2265_ (.A(net460),
    .B(net469),
    .C(\development_stage_sys.development_stage_level[2] ),
    .Y(_0351_));
 sg13g2_nand2_1 _2266_ (.Y(_0352_),
    .A(_0349_),
    .B(_0351_));
 sg13g2_nor2_1 _2267_ (.A(\development_stage_sys.development_stage_level[6] ),
    .B(_0350_),
    .Y(_0353_));
 sg13g2_nor3_1 _2268_ (.A(net457),
    .B(net458),
    .C(_0350_),
    .Y(_0354_));
 sg13g2_nand2_1 _2269_ (.Y(_0355_),
    .A(_0853_),
    .B(_0353_));
 sg13g2_nand3_1 _2270_ (.B(net440),
    .C(_0354_),
    .A(_0853_),
    .Y(_0356_));
 sg13g2_nor3_1 _2271_ (.A(net457),
    .B(net458),
    .C(\actions.development_stage[1] ),
    .Y(_0357_));
 sg13g2_o21ai_1 _2272_ (.B1(_0342_),
    .Y(_0358_),
    .A1(\actions.development_stage[1] ),
    .A2(_0356_));
 sg13g2_nand2_1 _2273_ (.Y(_0359_),
    .A(\development_stage_sys.development_stage_level[5] ),
    .B(\development_stage_sys.development_stage_level[4] ));
 sg13g2_and2_2 _2274_ (.A(net460),
    .B(\development_stage_sys.development_stage_level[2] ),
    .X(_0360_));
 sg13g2_and3_2 _2275_ (.X(_0361_),
    .A(net460),
    .B(\development_stage_sys.development_stage_level[3] ),
    .C(\development_stage_sys.development_stage_level[2] ));
 sg13g2_nand2_1 _2276_ (.Y(_0362_),
    .A(net459),
    .B(_0360_));
 sg13g2_nand2_1 _2277_ (.Y(_0363_),
    .A(net469),
    .B(_0361_));
 sg13g2_nand4_1 _2278_ (.B(\development_stage_sys.development_stage_level[5] ),
    .C(\development_stage_sys.development_stage_level[4] ),
    .A(\development_stage_sys.development_stage_level[0] ),
    .Y(_0364_),
    .D(_0361_));
 sg13g2_nand2_1 _2279_ (.Y(_0365_),
    .A(net457),
    .B(net458));
 sg13g2_nor2_1 _2280_ (.A(_0364_),
    .B(_0365_),
    .Y(_0366_));
 sg13g2_and2_1 _2281_ (.A(\actions.development_stage[1] ),
    .B(_0366_),
    .X(_0367_));
 sg13g2_nand2_1 _2282_ (.Y(_0368_),
    .A(net481),
    .B(_0367_));
 sg13g2_nand3_1 _2283_ (.B(_0341_),
    .C(_0368_),
    .A(_0340_),
    .Y(_0369_));
 sg13g2_nand2_1 _2284_ (.Y(_0370_),
    .A(_0358_),
    .B(_0369_));
 sg13g2_a21oi_1 _2285_ (.A1(net460),
    .A2(net469),
    .Y(_0371_),
    .B1(\development_stage_sys.development_stage_level[2] ));
 sg13g2_nand2_1 _2286_ (.Y(_0372_),
    .A(net460),
    .B(_0007_));
 sg13g2_nand4_1 _2287_ (.B(_0357_),
    .C(_0371_),
    .A(_0349_),
    .Y(_0373_),
    .D(_0372_));
 sg13g2_nand2_2 _2288_ (.Y(_0374_),
    .A(net441),
    .B(_0373_));
 sg13g2_nor2_1 _2289_ (.A(_0036_),
    .B(net441),
    .Y(_0375_));
 sg13g2_a21oi_1 _2290_ (.A1(net422),
    .A2(_0374_),
    .Y(_0376_),
    .B1(_0375_));
 sg13g2_a21oi_1 _2291_ (.A1(_0358_),
    .A2(_0369_),
    .Y(_0377_),
    .B1(_0376_));
 sg13g2_a21oi_1 _2292_ (.A1(_0343_),
    .A2(_0375_),
    .Y(_0378_),
    .B1(\development_stage_sys.development_stage_level[0] ));
 sg13g2_nand2_1 _2293_ (.Y(_0379_),
    .A(\development_stage_sys.development_stage_level[4] ),
    .B(_0361_));
 sg13g2_nor4_2 _2294_ (.A(_0007_),
    .B(_0359_),
    .C(_0362_),
    .Y(_0380_),
    .D(_0365_));
 sg13g2_nor2_2 _2295_ (.A(net439),
    .B(_0380_),
    .Y(_0381_));
 sg13g2_a21oi_1 _2296_ (.A1(_0343_),
    .A2(_0380_),
    .Y(_0382_),
    .B1(_0345_));
 sg13g2_nand3b_1 _2297_ (.B(net413),
    .C(_0378_),
    .Y(_0383_),
    .A_N(_0382_));
 sg13g2_o21ai_1 _2298_ (.B1(_0383_),
    .Y(_0121_),
    .A1(_0853_),
    .A2(_0377_));
 sg13g2_and2_2 _2299_ (.A(net501),
    .B(_0953_),
    .X(_0384_));
 sg13g2_nand2_2 _2300_ (.Y(_0385_),
    .A(net501),
    .B(_0953_));
 sg13g2_and2_2 _2301_ (.A(\talking.spi_bit_count[3] ),
    .B(_0384_),
    .X(_0386_));
 sg13g2_nand2_1 _2302_ (.Y(_0387_),
    .A(\talking.spi_bit_count[3] ),
    .B(_0384_));
 sg13g2_nor3_1 _2303_ (.A(\talking.address_reg[14] ),
    .B(\talking.address_reg[13] ),
    .C(\talking.address_reg[15] ),
    .Y(_0388_));
 sg13g2_nor4_1 _2304_ (.A(\talking.address_reg[10] ),
    .B(\talking.address_reg[9] ),
    .C(\talking.address_reg[12] ),
    .D(\talking.address_reg[11] ),
    .Y(_0389_));
 sg13g2_nor4_1 _2305_ (.A(\talking.address_reg[6] ),
    .B(\talking.address_reg[5] ),
    .C(\talking.address_reg[8] ),
    .D(\talking.address_reg[7] ),
    .Y(_0390_));
 sg13g2_nand3_1 _2306_ (.B(_0389_),
    .C(_0390_),
    .A(_0388_),
    .Y(_0391_));
 sg13g2_or2_1 _2307_ (.X(_0392_),
    .B(_0391_),
    .A(_0387_));
 sg13g2_nand2_1 _2308_ (.Y(_0393_),
    .A(_0954_),
    .B(_0387_));
 sg13g2_or2_1 _2309_ (.X(_0394_),
    .B(_0954_),
    .A(_0049_));
 sg13g2_nand3_1 _2310_ (.B(_0393_),
    .C(_0394_),
    .A(_0392_),
    .Y(_0395_));
 sg13g2_inv_1 _2311_ (.Y(_0396_),
    .A(net437));
 sg13g2_and3_1 _2312_ (.X(_0397_),
    .A(net529),
    .B(_0385_),
    .C(_0396_));
 sg13g2_nand3_1 _2313_ (.B(_0385_),
    .C(_0396_),
    .A(net529),
    .Y(_0398_));
 sg13g2_a22oi_1 _2314_ (.Y(_0399_),
    .B1(_0397_),
    .B2(\speech_planner_.variant_bit ),
    .A2(net437),
    .A1(net79));
 sg13g2_inv_1 _2315_ (.Y(_0122_),
    .A(_0399_));
 sg13g2_nand2_1 _2316_ (.Y(_0400_),
    .A(net51),
    .B(net438));
 sg13g2_or3_1 _2317_ (.A(_0899_),
    .B(_0906_),
    .C(_0976_),
    .X(_0401_));
 sg13g2_a21oi_1 _2318_ (.A1(_0916_),
    .A2(_0401_),
    .Y(_0402_),
    .B1(_0926_));
 sg13g2_o21ai_1 _2319_ (.B1(_0400_),
    .Y(_0123_),
    .A1(_0398_),
    .A2(_0402_));
 sg13g2_nand2b_1 _2320_ (.Y(_0403_),
    .B(_0916_),
    .A_N(_0899_));
 sg13g2_a21o_1 _2321_ (.A2(_0925_),
    .A1(_0849_),
    .B1(_0976_),
    .X(_0404_));
 sg13g2_a21oi_1 _2322_ (.A1(_0907_),
    .A2(_0404_),
    .Y(_0405_),
    .B1(_0403_));
 sg13g2_nor3_1 _2323_ (.A(_0928_),
    .B(_0398_),
    .C(_0405_),
    .Y(_0406_));
 sg13g2_a21o_1 _2324_ (.A2(net438),
    .A1(net76),
    .B1(_0406_),
    .X(_0124_));
 sg13g2_nor3_1 _2325_ (.A(_0903_),
    .B(_0906_),
    .C(_0404_),
    .Y(_0407_));
 sg13g2_nor4_1 _2326_ (.A(_0925_),
    .B(_0398_),
    .C(_0403_),
    .D(_0407_),
    .Y(_0408_));
 sg13g2_a21o_1 _2327_ (.A2(net438),
    .A1(net113),
    .B1(_0408_),
    .X(_0125_));
 sg13g2_nand2_1 _2328_ (.Y(_0409_),
    .A(net56),
    .B(net438));
 sg13g2_a21oi_1 _2329_ (.A1(\development_stage_sys.dev_stage_reg.cry ),
    .A2(_0858_),
    .Y(_0410_),
    .B1(net474));
 sg13g2_o21ai_1 _2330_ (.B1(_0409_),
    .Y(_0126_),
    .A1(_0398_),
    .A2(_0410_));
 sg13g2_nor2_1 _2331_ (.A(\development_stage_sys.dev_stage_reg.cry ),
    .B(\neurotransmitter.cortisol_system.cortisol_regulator.play ),
    .Y(_0411_));
 sg13g2_nor3_1 _2332_ (.A(net474),
    .B(_0398_),
    .C(_0411_),
    .Y(_0412_));
 sg13g2_a21o_1 _2333_ (.A2(net438),
    .A1(net102),
    .B1(_0412_),
    .X(_0127_));
 sg13g2_a22oi_1 _2334_ (.Y(_0413_),
    .B1(_0397_),
    .B2(\actions.development_stage[0] ),
    .A2(net437),
    .A1(net107));
 sg13g2_inv_1 _2335_ (.Y(_0128_),
    .A(_0413_));
 sg13g2_a22oi_1 _2336_ (.Y(_0414_),
    .B1(_0397_),
    .B2(\actions.development_stage[1] ),
    .A2(net437),
    .A1(net114));
 sg13g2_inv_1 _2337_ (.Y(_0129_),
    .A(_0414_));
 sg13g2_nand2_1 _2338_ (.Y(_0415_),
    .A(net79),
    .B(_0384_));
 sg13g2_nand2_1 _2339_ (.Y(_0416_),
    .A(\talking.address_reg[13] ),
    .B(net438));
 sg13g2_o21ai_1 _2340_ (.B1(_0416_),
    .Y(_0130_),
    .A1(net438),
    .A2(net80));
 sg13g2_nand2_1 _2341_ (.Y(_0417_),
    .A(net51),
    .B(_0384_));
 sg13g2_nand2_1 _2342_ (.Y(_0418_),
    .A(net74),
    .B(net437));
 sg13g2_o21ai_1 _2343_ (.B1(_0418_),
    .Y(_0131_),
    .A1(net437),
    .A2(_0417_));
 sg13g2_nand2_1 _2344_ (.Y(_0419_),
    .A(net76),
    .B(_0384_));
 sg13g2_nand2_1 _2345_ (.Y(_0420_),
    .A(\talking.address_reg[15] ),
    .B(net437));
 sg13g2_o21ai_1 _2346_ (.B1(_0420_),
    .Y(_0132_),
    .A1(net437),
    .A2(net77));
 sg13g2_nand2b_1 _2347_ (.Y(_0421_),
    .B(_1393_),
    .A_N(_0050_));
 sg13g2_or3_1 _2348_ (.A(\talking.skip_address_bytes[0] ),
    .B(\talking.skip_address_bytes[1] ),
    .C(net452),
    .X(_0422_));
 sg13g2_nor2b_1 _2349_ (.A(_1396_),
    .B_N(_0394_),
    .Y(_0423_));
 sg13g2_o21ai_1 _2350_ (.B1(_0423_),
    .Y(_0424_),
    .A1(_0050_),
    .A2(_0422_));
 sg13g2_nand2_1 _2351_ (.Y(_0425_),
    .A(_0954_),
    .B(_1394_));
 sg13g2_nor2_1 _2352_ (.A(_1382_),
    .B(_0425_),
    .Y(_0426_));
 sg13g2_or3_2 _2353_ (.A(_1390_),
    .B(_0424_),
    .C(_0426_),
    .X(_0427_));
 sg13g2_a21oi_2 _2354_ (.B1(_0427_),
    .Y(_0428_),
    .A2(net452),
    .A1(_1383_));
 sg13g2_mux2_1 _2355_ (.A0(_0428_),
    .A1(_0427_),
    .S(net127),
    .X(_0133_));
 sg13g2_nor2_2 _2356_ (.A(\talking.byte_count[1] ),
    .B(\talking.byte_count[0] ),
    .Y(_0429_));
 sg13g2_nand2_1 _2357_ (.Y(_0430_),
    .A(\talking.byte_count[1] ),
    .B(\talking.byte_count[0] ));
 sg13g2_nor2b_1 _2358_ (.A(_0429_),
    .B_N(_0430_),
    .Y(_0431_));
 sg13g2_nand2_1 _2359_ (.Y(_0432_),
    .A(_1393_),
    .B(_0431_));
 sg13g2_o21ai_1 _2360_ (.B1(_0432_),
    .Y(_0433_),
    .A1(_1388_),
    .A2(_0431_));
 sg13g2_mux2_1 _2361_ (.A0(_0433_),
    .A1(net126),
    .S(_0427_),
    .X(_0134_));
 sg13g2_o21ai_1 _2362_ (.B1(_1393_),
    .Y(_0434_),
    .A1(_0042_),
    .A2(_0430_));
 sg13g2_a21o_1 _2363_ (.A2(_0430_),
    .A1(_0042_),
    .B1(_0434_),
    .X(_0435_));
 sg13g2_xor2_1 _2364_ (.B(_0429_),
    .A(_0042_),
    .X(_0436_));
 sg13g2_o21ai_1 _2365_ (.B1(_0435_),
    .Y(_0437_),
    .A1(_1388_),
    .A2(_0436_));
 sg13g2_mux2_1 _2366_ (.A0(_0437_),
    .A1(net117),
    .S(_0427_),
    .X(_0135_));
 sg13g2_nand2b_2 _2367_ (.Y(_0438_),
    .B(_0429_),
    .A_N(\talking.byte_count[2] ));
 sg13g2_or3_1 _2368_ (.A(_0042_),
    .B(net452),
    .C(_0430_),
    .X(_0439_));
 sg13g2_nand2_1 _2369_ (.Y(_0440_),
    .A(_1387_),
    .B(_0438_));
 sg13g2_o21ai_1 _2370_ (.B1(_0439_),
    .Y(_0441_),
    .A1(_1388_),
    .A2(_0438_));
 sg13g2_a21oi_1 _2371_ (.A1(_0434_),
    .A2(_0440_),
    .Y(_0442_),
    .B1(net91));
 sg13g2_a21oi_1 _2372_ (.A1(net91),
    .A2(_0441_),
    .Y(_0443_),
    .B1(_0442_));
 sg13g2_a22oi_1 _2373_ (.Y(_0136_),
    .B1(_0428_),
    .B2(_0443_),
    .A2(_0427_),
    .A1(_0869_));
 sg13g2_nand4_1 _2374_ (.B(\talking.byte_count[2] ),
    .C(\talking.byte_count[1] ),
    .A(\talking.byte_count[3] ),
    .Y(_0444_),
    .D(\talking.byte_count[0] ));
 sg13g2_nand2_1 _2375_ (.Y(_0445_),
    .A(_0044_),
    .B(_0444_));
 sg13g2_nor2_1 _2376_ (.A(_0044_),
    .B(_0444_),
    .Y(_0446_));
 sg13g2_nor2_1 _2377_ (.A(net452),
    .B(_0446_),
    .Y(_0447_));
 sg13g2_nor3_1 _2378_ (.A(\talking.byte_count[3] ),
    .B(_0044_),
    .C(_0438_),
    .Y(_0448_));
 sg13g2_o21ai_1 _2379_ (.B1(_0044_),
    .Y(_0449_),
    .A1(\talking.byte_count[3] ),
    .A2(_0438_));
 sg13g2_nor2_1 _2380_ (.A(_1388_),
    .B(_0448_),
    .Y(_0450_));
 sg13g2_a22oi_1 _2381_ (.Y(_0451_),
    .B1(_0449_),
    .B2(_0450_),
    .A2(_0447_),
    .A1(_0445_));
 sg13g2_a22oi_1 _2382_ (.Y(_0137_),
    .B1(_0428_),
    .B2(_0451_),
    .A2(_0427_),
    .A1(_0868_));
 sg13g2_nand2_1 _2383_ (.Y(_0452_),
    .A(_1393_),
    .B(_0446_));
 sg13g2_nor2_1 _2384_ (.A(_1383_),
    .B(_1384_),
    .Y(_0453_));
 sg13g2_nor3_1 _2385_ (.A(_0051_),
    .B(_0447_),
    .C(_0453_),
    .Y(_0454_));
 sg13g2_a22oi_1 _2386_ (.Y(_0455_),
    .B1(_0454_),
    .B2(_0440_),
    .A2(_0452_),
    .A1(_0051_));
 sg13g2_mux2_1 _2387_ (.A0(_0455_),
    .A1(net93),
    .S(_0427_),
    .X(_0138_));
 sg13g2_nand2_1 _2388_ (.Y(_0456_),
    .A(net452),
    .B(_0385_));
 sg13g2_and2_2 _2389_ (.A(_0050_),
    .B(_0456_),
    .X(_0457_));
 sg13g2_nand2_1 _2390_ (.Y(_0458_),
    .A(net24),
    .B(_0457_));
 sg13g2_o21ai_1 _2391_ (.B1(net25),
    .Y(_0139_),
    .A1(_0865_),
    .A2(_0457_));
 sg13g2_and3_1 _2392_ (.X(_0459_),
    .A(_0048_),
    .B(_1379_),
    .C(_0394_));
 sg13g2_nand2_1 _2393_ (.Y(_0460_),
    .A(_0865_),
    .B(_0457_));
 sg13g2_and2_2 _2394_ (.A(_0459_),
    .B(_0460_),
    .X(_0461_));
 sg13g2_nor2_1 _2395_ (.A(\talking.spi_bit_count[3] ),
    .B(_0385_),
    .Y(_0462_));
 sg13g2_a21oi_2 _2396_ (.B1(\talking.spi_bit_count[3] ),
    .Y(_0463_),
    .A2(_0385_),
    .A1(net452));
 sg13g2_a21oi_1 _2397_ (.A1(_0461_),
    .A2(_0463_),
    .Y(_0464_),
    .B1(net86));
 sg13g2_a21oi_1 _2398_ (.A1(net86),
    .A2(_0461_),
    .Y(_0140_),
    .B1(net87));
 sg13g2_nand2_1 _2399_ (.Y(_0465_),
    .A(net86),
    .B(net63));
 sg13g2_nand2_1 _2400_ (.Y(_0466_),
    .A(_0457_),
    .B(_0465_));
 sg13g2_nand2_1 _2401_ (.Y(_0467_),
    .A(_0461_),
    .B(_0466_));
 sg13g2_a21oi_1 _2402_ (.A1(\talking.spi_bit_count[0] ),
    .A2(_0461_),
    .Y(_0468_),
    .B1(net63));
 sg13g2_a21oi_1 _2403_ (.A1(_0461_),
    .A2(_0466_),
    .Y(_0141_),
    .B1(net64));
 sg13g2_nand2_1 _2404_ (.Y(_0469_),
    .A(_0457_),
    .B(_0461_));
 sg13g2_nor3_1 _2405_ (.A(net97),
    .B(_0465_),
    .C(_0469_),
    .Y(_0470_));
 sg13g2_a21o_1 _2406_ (.A2(_0467_),
    .A1(net97),
    .B1(_0470_),
    .X(_0142_));
 sg13g2_nand2b_1 _2407_ (.Y(_0471_),
    .B(\talking.spi_bit_count[3] ),
    .A_N(_0461_));
 sg13g2_nand3_1 _2408_ (.B(net63),
    .C(net97),
    .A(net86),
    .Y(_0472_));
 sg13g2_o21ai_1 _2409_ (.B1(_0471_),
    .Y(_0143_),
    .A1(_0469_),
    .A2(_0472_));
 sg13g2_and2_1 _2410_ (.A(_0423_),
    .B(_0425_),
    .X(_0473_));
 sg13g2_o21ai_1 _2411_ (.B1(_0473_),
    .Y(_0474_),
    .A1(_0050_),
    .A2(_0422_));
 sg13g2_inv_1 _2412_ (.Y(_0475_),
    .A(_0474_));
 sg13g2_a21oi_1 _2413_ (.A1(net500),
    .A2(_0475_),
    .Y(_0476_),
    .B1(net95));
 sg13g2_a21oi_1 _2414_ (.A1(net95),
    .A2(_0473_),
    .Y(_0144_),
    .B1(net96));
 sg13g2_a21oi_1 _2415_ (.A1(\talking.skip_address_bytes[0] ),
    .A2(\talking.skip_address_bytes[1] ),
    .Y(_0477_),
    .B1(_1398_));
 sg13g2_a22oi_1 _2416_ (.Y(_0478_),
    .B1(_0477_),
    .B2(_0473_),
    .A2(_0474_),
    .A1(net33));
 sg13g2_inv_1 _2417_ (.Y(_0145_),
    .A(net34));
 sg13g2_a22oi_1 _2418_ (.Y(_0479_),
    .B1(_0462_),
    .B2(net24),
    .A2(_1396_),
    .A1(_0865_));
 sg13g2_nand4_1 _2419_ (.B(_0421_),
    .C(_0459_),
    .A(_0392_),
    .Y(_0480_),
    .D(_0479_));
 sg13g2_a22oi_1 _2420_ (.Y(_0481_),
    .B1(_0386_),
    .B2(\talking.address_reg[8] ),
    .A2(_1393_),
    .A1(net11));
 sg13g2_a21oi_1 _2421_ (.A1(_0456_),
    .A2(_0481_),
    .Y(_0482_),
    .B1(net420));
 sg13g2_a21o_1 _2422_ (.A2(net420),
    .A1(net111),
    .B1(_0482_),
    .X(_0146_));
 sg13g2_o21ai_1 _2423_ (.B1(net452),
    .Y(_0483_),
    .A1(\talking.spi_bit_count[3] ),
    .A2(_0385_));
 sg13g2_a22oi_1 _2424_ (.Y(_0484_),
    .B1(_0483_),
    .B2(\talking.spi_shift_reg[0] ),
    .A2(_0386_),
    .A1(net56));
 sg13g2_a21oi_1 _2425_ (.A1(_0456_),
    .A2(_0484_),
    .Y(_0485_),
    .B1(net420));
 sg13g2_a21o_1 _2426_ (.A2(net420),
    .A1(net109),
    .B1(_0485_),
    .X(_0147_));
 sg13g2_a221oi_1 _2427_ (.B2(\talking.spi_shift_reg[1] ),
    .C1(net421),
    .B1(_0483_),
    .A1(\talking.address_reg[10] ),
    .Y(_0486_),
    .A2(_0386_));
 sg13g2_a21oi_1 _2428_ (.A1(_0884_),
    .A2(net420),
    .Y(_0148_),
    .B1(_0486_));
 sg13g2_a221oi_1 _2429_ (.B2(net82),
    .C1(net420),
    .B1(_0483_),
    .A1(\talking.address_reg[11] ),
    .Y(_0487_),
    .A2(_0386_));
 sg13g2_a21oi_1 _2430_ (.A1(_0886_),
    .A2(net421),
    .Y(_0149_),
    .B1(_0487_));
 sg13g2_a221oi_1 _2431_ (.B2(\talking.spi_shift_reg[3] ),
    .C1(net420),
    .B1(_0483_),
    .A1(\talking.address_reg[12] ),
    .Y(_0488_),
    .A2(_0386_));
 sg13g2_a21oi_1 _2432_ (.A1(_0887_),
    .A2(net420),
    .Y(_0150_),
    .B1(_0488_));
 sg13g2_a221oi_1 _2433_ (.B2(\talking.spi_shift_reg[4] ),
    .C1(net421),
    .B1(_0483_),
    .A1(\talking.address_reg[13] ),
    .Y(_0489_),
    .A2(_0386_));
 sg13g2_a21oi_1 _2434_ (.A1(_0888_),
    .A2(net421),
    .Y(_0151_),
    .B1(_0489_));
 sg13g2_a221oi_1 _2435_ (.B2(net84),
    .C1(net421),
    .B1(_0483_),
    .A1(net74),
    .Y(_0490_),
    .A2(_0386_));
 sg13g2_a21oi_1 _2436_ (.A1(_0889_),
    .A2(net421),
    .Y(_0152_),
    .B1(_0490_));
 sg13g2_a221oi_1 _2437_ (.B2(\talking.spi_shift_reg[6] ),
    .C1(net421),
    .B1(_0483_),
    .A1(\talking.address_reg[15] ),
    .Y(_0491_),
    .A2(_0386_));
 sg13g2_a21oi_1 _2438_ (.A1(_0890_),
    .A2(net421),
    .Y(_0153_),
    .B1(_0491_));
 sg13g2_nor2_1 _2439_ (.A(_0050_),
    .B(_1398_),
    .Y(_0492_));
 sg13g2_a21oi_1 _2440_ (.A1(_0860_),
    .A2(net451),
    .Y(_0493_),
    .B1(_0492_));
 sg13g2_nand3_1 _2441_ (.B(_1397_),
    .C(_0493_),
    .A(_1391_),
    .Y(_0494_));
 sg13g2_nand2_1 _2442_ (.Y(_0495_),
    .A(\talking.uart_shift_reg[1] ),
    .B(net450));
 sg13g2_mux2_1 _2443_ (.A0(_0495_),
    .A1(net59),
    .S(net419),
    .X(_0154_));
 sg13g2_nor2_2 _2444_ (.A(net451),
    .B(_1382_),
    .Y(_0496_));
 sg13g2_a221oi_1 _2445_ (.B2(\talking.spi_shift_reg[0] ),
    .C1(net417),
    .B1(_0496_),
    .A1(\talking.uart_shift_reg[2] ),
    .Y(_0497_),
    .A2(net450));
 sg13g2_a21o_1 _2446_ (.A2(net417),
    .A1(net43),
    .B1(_0497_),
    .X(_0155_));
 sg13g2_a221oi_1 _2447_ (.B2(_0883_),
    .C1(net417),
    .B1(_0496_),
    .A1(_0882_),
    .Y(_0498_),
    .A2(net450));
 sg13g2_a21oi_1 _2448_ (.A1(_0839_),
    .A2(net417),
    .Y(_0156_),
    .B1(_0498_));
 sg13g2_a221oi_1 _2449_ (.B2(\talking.spi_shift_reg[2] ),
    .C1(net418),
    .B1(_0496_),
    .A1(\talking.uart_shift_reg[4] ),
    .Y(_0499_),
    .A2(net451));
 sg13g2_a21o_1 _2450_ (.A2(net417),
    .A1(net37),
    .B1(_0499_),
    .X(_0157_));
 sg13g2_a221oi_1 _2451_ (.B2(_0886_),
    .C1(net418),
    .B1(_0496_),
    .A1(_0885_),
    .Y(_0500_),
    .A2(net450));
 sg13g2_a21oi_1 _2452_ (.A1(_0838_),
    .A2(net418),
    .Y(_0158_),
    .B1(_0500_));
 sg13g2_a221oi_1 _2453_ (.B2(\talking.spi_shift_reg[4] ),
    .C1(net417),
    .B1(_0496_),
    .A1(\talking.uart_shift_reg[6] ),
    .Y(_0501_),
    .A2(net450));
 sg13g2_a21o_1 _2454_ (.A2(net417),
    .A1(net68),
    .B1(_0501_),
    .X(_0159_));
 sg13g2_a221oi_1 _2455_ (.B2(\talking.spi_shift_reg[5] ),
    .C1(net419),
    .B1(_0496_),
    .A1(\talking.uart_shift_reg[7] ),
    .Y(_0502_),
    .A2(net450));
 sg13g2_a21o_1 _2456_ (.A2(net417),
    .A1(net45),
    .B1(_0502_),
    .X(_0160_));
 sg13g2_a221oi_1 _2457_ (.B2(\talking.spi_shift_reg[6] ),
    .C1(net419),
    .B1(_0496_),
    .A1(\talking.uart_shift_reg[8] ),
    .Y(_0503_),
    .A2(net450));
 sg13g2_a21o_1 _2458_ (.A2(net419),
    .A1(net41),
    .B1(_0503_),
    .X(_0161_));
 sg13g2_a221oi_1 _2459_ (.B2(spi_mosi),
    .C1(net419),
    .B1(_0496_),
    .A1(\talking.uart_shift_reg[9] ),
    .Y(_0504_),
    .A2(net450));
 sg13g2_a21o_1 _2460_ (.A2(net419),
    .A1(net39),
    .B1(_0504_),
    .X(_0162_));
 sg13g2_mux2_1 _2461_ (.A0(net502),
    .A1(net54),
    .S(net419),
    .X(_0163_));
 sg13g2_a21oi_1 _2462_ (.A1(\talking.state[2] ),
    .A2(_1379_),
    .Y(_0505_),
    .B1(_0048_));
 sg13g2_o21ai_1 _2463_ (.B1(_1391_),
    .Y(_0506_),
    .A1(_0952_),
    .A2(_0505_));
 sg13g2_nand2b_1 _2464_ (.Y(_0507_),
    .B(_0394_),
    .A_N(_0463_));
 sg13g2_a21oi_2 _2465_ (.B1(_1377_),
    .Y(_0508_),
    .A2(_1380_),
    .A1(_0048_));
 sg13g2_a21oi_1 _2466_ (.A1(\talking.uart_active ),
    .A2(_1401_),
    .Y(_0509_),
    .B1(_0508_));
 sg13g2_nand2_1 _2467_ (.Y(_0510_),
    .A(_0384_),
    .B(_0391_));
 sg13g2_a21oi_1 _2468_ (.A1(\talking.state[2] ),
    .A2(_0049_),
    .Y(_0511_),
    .B1(net501));
 sg13g2_nor3_1 _2469_ (.A(\talking.state[2] ),
    .B(net500),
    .C(_0048_),
    .Y(_0512_));
 sg13g2_a21oi_1 _2470_ (.A1(\talking.state[2] ),
    .A2(net500),
    .Y(_0513_),
    .B1(_0512_));
 sg13g2_o21ai_1 _2471_ (.B1(_0510_),
    .Y(_0514_),
    .A1(_0511_),
    .A2(_0513_));
 sg13g2_or3_2 _2472_ (.A(_0507_),
    .B(_0509_),
    .C(_0514_),
    .X(_0515_));
 sg13g2_a21oi_1 _2473_ (.A1(_0422_),
    .A2(_0506_),
    .Y(_0516_),
    .B1(_0515_));
 sg13g2_a21o_1 _2474_ (.A2(_0515_),
    .A1(net501),
    .B1(_0516_),
    .X(_0164_));
 sg13g2_nand4_1 _2475_ (.B(_1391_),
    .C(_0385_),
    .A(_1378_),
    .Y(_0517_),
    .D(_0422_));
 sg13g2_mux2_1 _2476_ (.A0(_0517_),
    .A1(net500),
    .S(_0515_),
    .X(_0165_));
 sg13g2_nand3_1 _2477_ (.B(_1398_),
    .C(_0508_),
    .A(_1389_),
    .Y(_0518_));
 sg13g2_mux2_1 _2478_ (.A0(_0518_),
    .A1(net128),
    .S(_0515_),
    .X(_0166_));
 sg13g2_nor3_2 _2479_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.play ),
    .B(_0902_),
    .C(_0975_),
    .Y(_0519_));
 sg13g2_nand3_1 _2480_ (.B(net498),
    .C(net462),
    .A(net481),
    .Y(_0520_));
 sg13g2_or2_1 _2481_ (.X(_0521_),
    .B(_0520_),
    .A(_1144_));
 sg13g2_nor2b_2 _2482_ (.A(_0519_),
    .B_N(_0521_),
    .Y(_0522_));
 sg13g2_nand2b_1 _2483_ (.Y(_0523_),
    .B(_0521_),
    .A_N(_0519_));
 sg13g2_nand2_1 _2484_ (.Y(_0524_),
    .A(\vital_energy_sys.vital_energy[3] ),
    .B(\vital_energy_sys.vital_energy[2] ));
 sg13g2_nand2_1 _2485_ (.Y(_0525_),
    .A(\vital_energy_sys.vital_energy[5] ),
    .B(\vital_energy_sys.vital_energy[4] ));
 sg13g2_nor3_1 _2486_ (.A(_0943_),
    .B(_0524_),
    .C(_0525_),
    .Y(_0526_));
 sg13g2_and2_1 _2487_ (.A(_0848_),
    .B(_0526_),
    .X(_0527_));
 sg13g2_nand2_2 _2488_ (.Y(_0528_),
    .A(\vital_energy_sys.vital_energy[1] ),
    .B(\vital_energy_sys.vital_energy[0] ));
 sg13g2_nand3_1 _2489_ (.B(\vital_energy_sys.vital_energy[0] ),
    .C(_0527_),
    .A(\vital_energy_sys.vital_energy[1] ),
    .Y(_0529_));
 sg13g2_o21ai_1 _2490_ (.B1(_0529_),
    .Y(_0530_),
    .A1(_0961_),
    .A2(_0973_));
 sg13g2_and2_2 _2491_ (.A(net436),
    .B(_0530_),
    .X(_0531_));
 sg13g2_nand2_2 _2492_ (.Y(_0532_),
    .A(net436),
    .B(_0530_));
 sg13g2_a21oi_1 _2493_ (.A1(_0960_),
    .A2(_0972_),
    .Y(_0533_),
    .B1(_0527_));
 sg13g2_a21oi_2 _2494_ (.B1(_0531_),
    .Y(_0534_),
    .A2(_0533_),
    .A1(_0522_));
 sg13g2_nand2b_1 _2495_ (.Y(_0535_),
    .B(\vital_energy_sys.vital_energy[0] ),
    .A_N(_0534_));
 sg13g2_nand2_1 _2496_ (.Y(_0536_),
    .A(_0522_),
    .B(_0526_));
 sg13g2_nand2_2 _2497_ (.Y(_0537_),
    .A(net479),
    .B(_0536_));
 sg13g2_a21oi_1 _2498_ (.A1(_0024_),
    .A2(net436),
    .Y(_0538_),
    .B1(_0537_));
 sg13g2_o21ai_1 _2499_ (.B1(net456),
    .Y(_0539_),
    .A1(\vital_energy_sys.vital_energy[0] ),
    .A2(_0522_));
 sg13g2_nand2_1 _2500_ (.Y(_0540_),
    .A(_0534_),
    .B(_0539_));
 sg13g2_o21ai_1 _2501_ (.B1(_0535_),
    .Y(_0167_),
    .A1(_0538_),
    .A2(_0540_));
 sg13g2_nand2_1 _2502_ (.Y(_0541_),
    .A(net436),
    .B(_0528_));
 sg13g2_o21ai_1 _2503_ (.B1(_0536_),
    .Y(_0542_),
    .A1(_0958_),
    .A2(_0541_));
 sg13g2_nor2_1 _2504_ (.A(_0519_),
    .B(_0542_),
    .Y(_0543_));
 sg13g2_a21oi_1 _2505_ (.A1(net456),
    .A2(_0542_),
    .Y(_0544_),
    .B1(_0543_));
 sg13g2_mux2_1 _2506_ (.A0(\vital_energy_sys.vital_energy[1] ),
    .A1(_0544_),
    .S(_0534_),
    .X(_0168_));
 sg13g2_a21oi_1 _2507_ (.A1(_1394_),
    .A2(_0508_),
    .Y(_0545_),
    .B1(_1396_));
 sg13g2_nor2b_1 _2508_ (.A(_0492_),
    .B_N(_0545_),
    .Y(_0546_));
 sg13g2_o21ai_1 _2509_ (.B1(_0546_),
    .Y(_0547_),
    .A1(\talking.uart_active ),
    .A2(_0508_));
 sg13g2_nand2b_2 _2510_ (.Y(_0548_),
    .B(net451),
    .A_N(_0547_));
 sg13g2_nand2_1 _2511_ (.Y(_0549_),
    .A(net119),
    .B(_0547_));
 sg13g2_o21ai_1 _2512_ (.B1(_0549_),
    .Y(_0169_),
    .A1(net119),
    .A2(_0548_));
 sg13g2_nor2_1 _2513_ (.A(_1377_),
    .B(_1402_),
    .Y(_0550_));
 sg13g2_xnor2_1 _2514_ (.Y(_0551_),
    .A(net119),
    .B(net120));
 sg13g2_nor3_1 _2515_ (.A(_0548_),
    .B(_0550_),
    .C(_0551_),
    .Y(_0552_));
 sg13g2_a21o_1 _2516_ (.A2(_0547_),
    .A1(net120),
    .B1(_0552_),
    .X(_0170_));
 sg13g2_nand2_1 _2517_ (.Y(_0553_),
    .A(net72),
    .B(_0547_));
 sg13g2_a21oi_1 _2518_ (.A1(\talking.uart_bit_count[0] ),
    .A2(\talking.uart_bit_count[1] ),
    .Y(_0554_),
    .B1(net72));
 sg13g2_nand3_1 _2519_ (.B(\talking.uart_bit_count[1] ),
    .C(net72),
    .A(\talking.uart_bit_count[0] ),
    .Y(_0555_));
 sg13g2_nand2b_1 _2520_ (.Y(_0556_),
    .B(_0555_),
    .A_N(_0554_));
 sg13g2_o21ai_1 _2521_ (.B1(_0553_),
    .Y(_0171_),
    .A1(_0548_),
    .A2(_0556_));
 sg13g2_xor2_1 _2522_ (.B(_0555_),
    .A(net108),
    .X(_0557_));
 sg13g2_nor3_1 _2523_ (.A(_0548_),
    .B(_0550_),
    .C(_0557_),
    .Y(_0558_));
 sg13g2_a21o_1 _2524_ (.A2(_0547_),
    .A1(net108),
    .B1(_0558_),
    .X(_0172_));
 sg13g2_nand2_1 _2525_ (.Y(_0559_),
    .A(\vital_energy_sys.vital_energy[2] ),
    .B(_0531_));
 sg13g2_a21oi_2 _2526_ (.B1(net436),
    .Y(_0560_),
    .A2(_0960_),
    .A1(net454));
 sg13g2_nor3_1 _2527_ (.A(\vital_energy_sys.vital_energy[1] ),
    .B(\vital_energy_sys.vital_energy[0] ),
    .C(\vital_energy_sys.vital_energy[2] ),
    .Y(_0561_));
 sg13g2_xnor2_1 _2528_ (.Y(_0562_),
    .A(_0871_),
    .B(_0958_));
 sg13g2_a221oi_1 _2529_ (.B2(_0523_),
    .C1(net479),
    .B1(_0562_),
    .A1(_0871_),
    .Y(_0563_),
    .A2(_0560_));
 sg13g2_xnor2_1 _2530_ (.Y(_0564_),
    .A(_0871_),
    .B(_0528_));
 sg13g2_nor2_1 _2531_ (.A(_0025_),
    .B(net435),
    .Y(_0565_));
 sg13g2_a21oi_1 _2532_ (.A1(net435),
    .A2(_0564_),
    .Y(_0566_),
    .B1(_0565_));
 sg13g2_o21ai_1 _2533_ (.B1(_0532_),
    .Y(_0567_),
    .A1(_0537_),
    .A2(_0566_));
 sg13g2_o21ai_1 _2534_ (.B1(_0559_),
    .Y(_0173_),
    .A1(_0563_),
    .A2(_0567_));
 sg13g2_nand2b_1 _2535_ (.Y(_0568_),
    .B(_0524_),
    .A_N(_0959_));
 sg13g2_nand2_1 _2536_ (.Y(_0569_),
    .A(_0958_),
    .B(_0959_));
 sg13g2_xor2_1 _2537_ (.B(_0561_),
    .A(\vital_energy_sys.vital_energy[3] ),
    .X(_0570_));
 sg13g2_a221oi_1 _2538_ (.B2(net435),
    .C1(net480),
    .B1(_0570_),
    .A1(_0560_),
    .Y(_0571_),
    .A2(_0568_));
 sg13g2_nor2_1 _2539_ (.A(_0025_),
    .B(_0528_),
    .Y(_0572_));
 sg13g2_xor2_1 _2540_ (.B(_0572_),
    .A(\vital_energy_sys.vital_energy[3] ),
    .X(_0573_));
 sg13g2_nand2_1 _2541_ (.Y(_0574_),
    .A(net435),
    .B(_0573_));
 sg13g2_o21ai_1 _2542_ (.B1(_0574_),
    .Y(_0575_),
    .A1(net435),
    .A2(_0568_));
 sg13g2_o21ai_1 _2543_ (.B1(_0532_),
    .Y(_0576_),
    .A1(_0537_),
    .A2(_0575_));
 sg13g2_o21ai_1 _2544_ (.B1(_0559_),
    .Y(_0174_),
    .A1(_0571_),
    .A2(_0576_));
 sg13g2_nand2_1 _2545_ (.Y(_0577_),
    .A(_0026_),
    .B(_0959_));
 sg13g2_xnor2_1 _2546_ (.Y(_0578_),
    .A(_0026_),
    .B(_0959_));
 sg13g2_xnor2_1 _2547_ (.Y(_0579_),
    .A(\vital_energy_sys.vital_energy[4] ),
    .B(_0569_));
 sg13g2_a221oi_1 _2548_ (.B2(net435),
    .C1(net479),
    .B1(_0579_),
    .A1(_0560_),
    .Y(_0580_),
    .A2(_0578_));
 sg13g2_a21o_2 _2549_ (.A2(_0528_),
    .A1(net435),
    .B1(_0524_),
    .X(_0581_));
 sg13g2_nor2_1 _2550_ (.A(_0537_),
    .B(_0581_),
    .Y(_0582_));
 sg13g2_a21o_1 _2551_ (.A2(_0582_),
    .A1(\vital_energy_sys.vital_energy[4] ),
    .B1(_0580_),
    .X(_0583_));
 sg13g2_nand2_1 _2552_ (.Y(_0584_),
    .A(net479),
    .B(_0581_));
 sg13g2_a21oi_1 _2553_ (.A1(_0532_),
    .A2(_0584_),
    .Y(_0585_),
    .B1(\vital_energy_sys.vital_energy[4] ));
 sg13g2_a21oi_1 _2554_ (.A1(_0532_),
    .A2(_0583_),
    .Y(_0175_),
    .B1(_0585_));
 sg13g2_o21ai_1 _2555_ (.B1(net479),
    .Y(_0586_),
    .A1(_0026_),
    .A2(_0581_));
 sg13g2_nand2_1 _2556_ (.Y(_0587_),
    .A(_0532_),
    .B(_0586_));
 sg13g2_nor3_1 _2557_ (.A(\vital_energy_sys.vital_energy[5] ),
    .B(_0026_),
    .C(_0581_),
    .Y(_0588_));
 sg13g2_nor2_1 _2558_ (.A(_0537_),
    .B(_0588_),
    .Y(_0589_));
 sg13g2_xnor2_1 _2559_ (.Y(_0590_),
    .A(\vital_energy_sys.vital_energy[5] ),
    .B(_0577_));
 sg13g2_o21ai_1 _2560_ (.B1(\vital_energy_sys.vital_energy[5] ),
    .Y(_0591_),
    .A1(\vital_energy_sys.vital_energy[4] ),
    .A2(_0569_));
 sg13g2_nand2_1 _2561_ (.Y(_0592_),
    .A(_0961_),
    .B(_0591_));
 sg13g2_a221oi_1 _2562_ (.B2(net435),
    .C1(net479),
    .B1(_0592_),
    .A1(_0560_),
    .Y(_0593_),
    .A2(_0590_));
 sg13g2_nor3_1 _2563_ (.A(_0531_),
    .B(_0589_),
    .C(_0593_),
    .Y(_0594_));
 sg13g2_a21o_1 _2564_ (.A2(_0587_),
    .A1(\vital_energy_sys.vital_energy[5] ),
    .B1(_0594_),
    .X(_0176_));
 sg13g2_nor2_1 _2565_ (.A(_0525_),
    .B(_0581_),
    .Y(_0595_));
 sg13g2_xnor2_1 _2566_ (.Y(_0596_),
    .A(net468),
    .B(_0595_));
 sg13g2_nand2b_1 _2567_ (.Y(_0597_),
    .B(_0522_),
    .A_N(_0943_));
 sg13g2_and3_1 _2568_ (.X(_0598_),
    .A(net479),
    .B(_0596_),
    .C(_0597_));
 sg13g2_nor2_1 _2569_ (.A(net468),
    .B(_0961_),
    .Y(_0599_));
 sg13g2_nand2_1 _2570_ (.Y(_0600_),
    .A(_0027_),
    .B(_0960_));
 sg13g2_xnor2_1 _2571_ (.Y(_0601_),
    .A(_0027_),
    .B(_0960_));
 sg13g2_xnor2_1 _2572_ (.Y(_0602_),
    .A(net468),
    .B(_0961_));
 sg13g2_a22oi_1 _2573_ (.Y(_0603_),
    .B1(_0602_),
    .B2(net436),
    .A2(_0601_),
    .A1(_0560_));
 sg13g2_a21o_1 _2574_ (.A2(_0603_),
    .A1(net456),
    .B1(_0531_),
    .X(_0604_));
 sg13g2_o21ai_1 _2575_ (.B1(_0559_),
    .Y(_0177_),
    .A1(_0598_),
    .A2(_0604_));
 sg13g2_nand2_1 _2576_ (.Y(_0605_),
    .A(_0083_),
    .B(_0531_));
 sg13g2_nor3_1 _2577_ (.A(_0027_),
    .B(_0525_),
    .C(_0581_),
    .Y(_0606_));
 sg13g2_xnor2_1 _2578_ (.Y(_0607_),
    .A(net467),
    .B(_0606_));
 sg13g2_a21oi_1 _2579_ (.A1(_0597_),
    .A2(_0607_),
    .Y(_0608_),
    .B1(net455));
 sg13g2_xnor2_1 _2580_ (.Y(_0609_),
    .A(net467),
    .B(_0600_));
 sg13g2_xor2_1 _2581_ (.B(_0599_),
    .A(net467),
    .X(_0610_));
 sg13g2_a22oi_1 _2582_ (.Y(_0611_),
    .B1(_0610_),
    .B2(net436),
    .A2(_0609_),
    .A1(_0560_));
 sg13g2_o21ai_1 _2583_ (.B1(_0532_),
    .Y(_0612_),
    .A1(net479),
    .A2(_0611_));
 sg13g2_o21ai_1 _2584_ (.B1(_0605_),
    .Y(_0178_),
    .A1(_0608_),
    .A2(_0612_));
 sg13g2_nor2_2 _2585_ (.A(_0944_),
    .B(_1331_),
    .Y(_0613_));
 sg13g2_xnor2_1 _2586_ (.Y(_0614_),
    .A(\nourishment.glucose[2] ),
    .B(_1327_));
 sg13g2_a221oi_1 _2587_ (.B2(_0945_),
    .C1(_0613_),
    .B1(_0614_),
    .A1(_0880_),
    .Y(_0179_),
    .A2(_1326_));
 sg13g2_xnor2_1 _2588_ (.Y(_0615_),
    .A(\nourishment.glucose[3] ),
    .B(\nourishment.glucose[2] ));
 sg13g2_xnor2_1 _2589_ (.Y(_0616_),
    .A(\nourishment.glucose[3] ),
    .B(_1328_));
 sg13g2_a221oi_1 _2590_ (.B2(_0945_),
    .C1(_0613_),
    .B1(_0616_),
    .A1(_1326_),
    .Y(_0180_),
    .A2(_0615_));
 sg13g2_xor2_1 _2591_ (.B(_1322_),
    .A(\nourishment.glucose[4] ),
    .X(_0617_));
 sg13g2_xor2_1 _2592_ (.B(_1329_),
    .A(\nourishment.glucose[4] ),
    .X(_0618_));
 sg13g2_a221oi_1 _2593_ (.B2(_0945_),
    .C1(_0613_),
    .B1(_0618_),
    .A1(_1326_),
    .Y(_0181_),
    .A2(_0617_));
 sg13g2_nor2_1 _2594_ (.A(_0030_),
    .B(_1322_),
    .Y(_0619_));
 sg13g2_xnor2_1 _2595_ (.Y(_0620_),
    .A(\nourishment.glucose[5] ),
    .B(_0619_));
 sg13g2_o21ai_1 _2596_ (.B1(\nourishment.glucose[5] ),
    .Y(_0621_),
    .A1(\nourishment.glucose[4] ),
    .A2(_1329_));
 sg13g2_nor2_1 _2597_ (.A(net453),
    .B(_1330_),
    .Y(_0622_));
 sg13g2_a221oi_1 _2598_ (.B2(_0622_),
    .C1(_0613_),
    .B1(_0621_),
    .A1(_1326_),
    .Y(_0182_),
    .A2(_0620_));
 sg13g2_nand2b_1 _2599_ (.Y(_0623_),
    .B(\nourishment.glucose[6] ),
    .A_N(_1330_));
 sg13g2_a21oi_1 _2600_ (.A1(_0846_),
    .A2(_1330_),
    .Y(_0624_),
    .B1(net453));
 sg13g2_nand3_1 _2601_ (.B(_0847_),
    .C(_1323_),
    .A(\nourishment.glucose[6] ),
    .Y(_0625_));
 sg13g2_o21ai_1 _2602_ (.B1(_0625_),
    .Y(_0626_),
    .A1(\nourishment.glucose[6] ),
    .A2(_1323_));
 sg13g2_a221oi_1 _2603_ (.B2(net453),
    .C1(_0613_),
    .B1(_0626_),
    .A1(_0623_),
    .Y(_0183_),
    .A2(_0624_));
 sg13g2_nand2b_1 _2604_ (.Y(_0627_),
    .B(_1323_),
    .A_N(_0031_));
 sg13g2_a21oi_1 _2605_ (.A1(_0846_),
    .A2(net465),
    .Y(_0628_),
    .B1(_0627_));
 sg13g2_a21o_1 _2606_ (.A2(_0627_),
    .A1(net465),
    .B1(_0628_),
    .X(_0629_));
 sg13g2_nor3_1 _2607_ (.A(_0084_),
    .B(net453),
    .C(_1331_),
    .Y(_0630_));
 sg13g2_a221oi_1 _2608_ (.B2(net453),
    .C1(_0630_),
    .B1(_0629_),
    .A1(net465),
    .Y(_0184_),
    .A2(_0624_));
 sg13g2_xnor2_1 _2609_ (.Y(_0631_),
    .A(net464),
    .B(net488));
 sg13g2_nor2_1 _2610_ (.A(net464),
    .B(_1369_),
    .Y(_0632_));
 sg13g2_mux2_1 _2611_ (.A0(_0631_),
    .A1(_0632_),
    .S(net426),
    .X(_0633_));
 sg13g2_a22oi_1 _2612_ (.Y(_0634_),
    .B1(_0631_),
    .B2(net427),
    .A2(_1367_),
    .A1(net464));
 sg13g2_mux2_1 _2613_ (.A0(_0633_),
    .A1(_0634_),
    .S(net444),
    .X(_0635_));
 sg13g2_mux2_1 _2614_ (.A0(_0635_),
    .A1(net464),
    .S(net414),
    .X(_0185_));
 sg13g2_o21ai_1 _2615_ (.B1(\neurotransmitter.cortisol_system.cortisol[2] ),
    .Y(_0636_),
    .A1(net464),
    .A2(net488));
 sg13g2_o21ai_1 _2616_ (.B1(_0636_),
    .Y(_0637_),
    .A1(net489),
    .A2(_1360_));
 sg13g2_nand2b_1 _2617_ (.Y(_0638_),
    .B(_1360_),
    .A_N(_1353_));
 sg13g2_nand2_1 _2618_ (.Y(_0639_),
    .A(_1371_),
    .B(_0638_));
 sg13g2_a21oi_1 _2619_ (.A1(net426),
    .A2(_0639_),
    .Y(_0640_),
    .B1(net444));
 sg13g2_o21ai_1 _2620_ (.B1(_0640_),
    .Y(_0641_),
    .A1(net426),
    .A2(_0637_));
 sg13g2_a21o_1 _2621_ (.A2(_1353_),
    .A1(net488),
    .B1(_1368_),
    .X(_0642_));
 sg13g2_a22oi_1 _2622_ (.Y(_0643_),
    .B1(_0642_),
    .B2(net427),
    .A2(_0638_),
    .A1(_1367_));
 sg13g2_a21oi_1 _2623_ (.A1(net444),
    .A2(_0643_),
    .Y(_0644_),
    .B1(net414));
 sg13g2_a22oi_1 _2624_ (.Y(_0186_),
    .B1(_0641_),
    .B2(_0644_),
    .A2(net414),
    .A1(_0873_));
 sg13g2_o21ai_1 _2625_ (.B1(\neurotransmitter.cortisol_system.cortisol[3] ),
    .Y(_0645_),
    .A1(net488),
    .A2(_1360_));
 sg13g2_nand3_1 _2626_ (.B(_1362_),
    .C(_0645_),
    .A(net427),
    .Y(_0646_));
 sg13g2_o21ai_1 _2627_ (.B1(_1371_),
    .Y(_0647_),
    .A1(_0021_),
    .A2(_1360_));
 sg13g2_a21o_1 _2628_ (.A2(_1360_),
    .A1(_0021_),
    .B1(_0647_),
    .X(_0648_));
 sg13g2_a21oi_1 _2629_ (.A1(net426),
    .A2(_0648_),
    .Y(_0649_),
    .B1(net444));
 sg13g2_xnor2_1 _2630_ (.Y(_0650_),
    .A(\neurotransmitter.cortisol_system.cortisol[3] ),
    .B(_1353_));
 sg13g2_xnor2_1 _2631_ (.Y(_0651_),
    .A(_0872_),
    .B(_1356_));
 sg13g2_a22oi_1 _2632_ (.Y(_0652_),
    .B1(_0651_),
    .B2(net427),
    .A2(_0650_),
    .A1(_1367_));
 sg13g2_a221oi_1 _2633_ (.B2(net444),
    .C1(net414),
    .B1(_0652_),
    .A1(_0646_),
    .Y(_0653_),
    .A2(_0649_));
 sg13g2_a21oi_1 _2634_ (.A1(_0872_),
    .A2(net414),
    .Y(_0187_),
    .B1(_0653_));
 sg13g2_nor2b_1 _2635_ (.A(_0021_),
    .B_N(_1353_),
    .Y(_0654_));
 sg13g2_xnor2_1 _2636_ (.Y(_0655_),
    .A(\neurotransmitter.cortisol_system.cortisol[4] ),
    .B(_0654_));
 sg13g2_xnor2_1 _2637_ (.Y(_0656_),
    .A(\neurotransmitter.cortisol_system.cortisol[4] ),
    .B(_1357_));
 sg13g2_o21ai_1 _2638_ (.B1(net444),
    .Y(_0657_),
    .A1(net426),
    .A2(_0656_));
 sg13g2_a21oi_1 _2639_ (.A1(_1367_),
    .A2(_0655_),
    .Y(_0658_),
    .B1(_0657_));
 sg13g2_xnor2_1 _2640_ (.Y(_0659_),
    .A(_0022_),
    .B(_1361_));
 sg13g2_a21oi_1 _2641_ (.A1(_1371_),
    .A2(_0659_),
    .Y(_0660_),
    .B1(net427));
 sg13g2_nand2_2 _2642_ (.Y(_0661_),
    .A(_0874_),
    .B(_1361_));
 sg13g2_nor2_2 _2643_ (.A(net489),
    .B(_0661_),
    .Y(_0662_));
 sg13g2_a21oi_1 _2644_ (.A1(\neurotransmitter.cortisol_system.cortisol[4] ),
    .A2(_1362_),
    .Y(_0663_),
    .B1(_0662_));
 sg13g2_a21oi_1 _2645_ (.A1(net427),
    .A2(_0663_),
    .Y(_0664_),
    .B1(net444));
 sg13g2_nor2b_1 _2646_ (.A(_0660_),
    .B_N(_0664_),
    .Y(_0665_));
 sg13g2_nor3_1 _2647_ (.A(net414),
    .B(_0658_),
    .C(_0665_),
    .Y(_0666_));
 sg13g2_a21oi_1 _2648_ (.A1(_0874_),
    .A2(net414),
    .Y(_0188_),
    .B1(_0666_));
 sg13g2_xnor2_1 _2649_ (.Y(_0667_),
    .A(net463),
    .B(_1354_));
 sg13g2_nor2_1 _2650_ (.A(_0022_),
    .B(_1357_),
    .Y(_0668_));
 sg13g2_xnor2_1 _2651_ (.Y(_0669_),
    .A(net463),
    .B(_0668_));
 sg13g2_a22oi_1 _2652_ (.Y(_0670_),
    .B1(_0669_),
    .B2(net427),
    .A2(_0667_),
    .A1(_1367_));
 sg13g2_o21ai_1 _2653_ (.B1(_1371_),
    .Y(_0671_),
    .A1(_0023_),
    .A2(_0661_));
 sg13g2_a21oi_1 _2654_ (.A1(_0023_),
    .A2(_0661_),
    .Y(_0672_),
    .B1(_0671_));
 sg13g2_nor2_1 _2655_ (.A(net463),
    .B(_0661_),
    .Y(_0673_));
 sg13g2_xnor2_1 _2656_ (.Y(_0674_),
    .A(net463),
    .B(_0662_));
 sg13g2_a21oi_1 _2657_ (.A1(net428),
    .A2(_0674_),
    .Y(_0675_),
    .B1(net445));
 sg13g2_o21ai_1 _2658_ (.B1(_0675_),
    .Y(_0676_),
    .A1(net428),
    .A2(_0672_));
 sg13g2_a21oi_1 _2659_ (.A1(net444),
    .A2(_0670_),
    .Y(_0677_),
    .B1(net415));
 sg13g2_a22oi_1 _2660_ (.Y(_0189_),
    .B1(_0676_),
    .B2(_0677_),
    .A2(net415),
    .A1(_0843_));
 sg13g2_nand2_1 _2661_ (.Y(_0678_),
    .A(_0904_),
    .B(_0662_));
 sg13g2_o21ai_1 _2662_ (.B1(_0678_),
    .Y(_0679_),
    .A1(_0844_),
    .A2(_0662_));
 sg13g2_xnor2_1 _2663_ (.Y(_0680_),
    .A(_0052_),
    .B(_0673_));
 sg13g2_a21oi_1 _2664_ (.A1(_1371_),
    .A2(_0680_),
    .Y(_0681_),
    .B1(net428));
 sg13g2_nor2_1 _2665_ (.A(net446),
    .B(_0681_),
    .Y(_0682_));
 sg13g2_o21ai_1 _2666_ (.B1(_0682_),
    .Y(_0683_),
    .A1(net426),
    .A2(_0679_));
 sg13g2_nor2b_1 _2667_ (.A(_0023_),
    .B_N(_1354_),
    .Y(_0684_));
 sg13g2_xnor2_1 _2668_ (.Y(_0685_),
    .A(net462),
    .B(_0684_));
 sg13g2_xnor2_1 _2669_ (.Y(_0686_),
    .A(_0844_),
    .B(_1358_));
 sg13g2_a22oi_1 _2670_ (.Y(_0687_),
    .B1(_0686_),
    .B2(net427),
    .A2(_0685_),
    .A1(_1367_));
 sg13g2_a21oi_1 _2671_ (.A1(net446),
    .A2(_0687_),
    .Y(_0688_),
    .B1(net415));
 sg13g2_a22oi_1 _2672_ (.Y(_0190_),
    .B1(_0683_),
    .B2(_0688_),
    .A2(net414),
    .A1(_0844_));
 sg13g2_nand2_2 _2673_ (.Y(_0689_),
    .A(\illness_sys.illness[3] ),
    .B(net423));
 sg13g2_nor2_1 _2674_ (.A(_0304_),
    .B(_0327_),
    .Y(_0690_));
 sg13g2_xnor2_1 _2675_ (.Y(_0691_),
    .A(net461),
    .B(_0310_));
 sg13g2_nor2_1 _2676_ (.A(_0033_),
    .B(_0327_),
    .Y(_0692_));
 sg13g2_nand2b_1 _2677_ (.Y(_0693_),
    .B(_0331_),
    .A_N(net461));
 sg13g2_xnor2_1 _2678_ (.Y(_0694_),
    .A(net461),
    .B(_0314_));
 sg13g2_mux4_1 _2679_ (.S0(net442),
    .A0(_0691_),
    .A1(_0692_),
    .A2(_0694_),
    .A3(_0693_),
    .S1(net470),
    .X(_0695_));
 sg13g2_o21ai_1 _2680_ (.B1(_0689_),
    .Y(_0191_),
    .A1(net423),
    .A2(_0695_));
 sg13g2_a21oi_1 _2681_ (.A1(_0305_),
    .A2(_0327_),
    .Y(_0696_),
    .B1(net470));
 sg13g2_nor2_1 _2682_ (.A(_0306_),
    .B(_0318_),
    .Y(_0697_));
 sg13g2_nor2_1 _2683_ (.A(_0304_),
    .B(_0697_),
    .Y(_0698_));
 sg13g2_nor2_1 _2684_ (.A(_0033_),
    .B(_0311_),
    .Y(_0699_));
 sg13g2_xor2_1 _2685_ (.B(_0699_),
    .A(\illness_sys.illness[3] ),
    .X(_0700_));
 sg13g2_nor2_1 _2686_ (.A(net443),
    .B(_0700_),
    .Y(_0701_));
 sg13g2_o21ai_1 _2687_ (.B1(_0696_),
    .Y(_0702_),
    .A1(_0698_),
    .A2(_0701_));
 sg13g2_xnor2_1 _2688_ (.Y(_0703_),
    .A(\illness_sys.illness[3] ),
    .B(_0321_));
 sg13g2_nor3_1 _2689_ (.A(_0302_),
    .B(_0332_),
    .C(_0697_),
    .Y(_0704_));
 sg13g2_o21ai_1 _2690_ (.B1(net470),
    .Y(_0705_),
    .A1(net443),
    .A2(_0703_));
 sg13g2_o21ai_1 _2691_ (.B1(_0702_),
    .Y(_0706_),
    .A1(_0704_),
    .A2(_0705_));
 sg13g2_o21ai_1 _2692_ (.B1(_0689_),
    .Y(_0192_),
    .A1(net423),
    .A2(_0706_));
 sg13g2_o21ai_1 _2693_ (.B1(_0306_),
    .Y(_0707_),
    .A1(_0305_),
    .A2(_0310_));
 sg13g2_xor2_1 _2694_ (.B(_0707_),
    .A(\illness_sys.illness[4] ),
    .X(_0708_));
 sg13g2_nand2_1 _2695_ (.Y(_0709_),
    .A(_0696_),
    .B(_0708_));
 sg13g2_nand2_1 _2696_ (.Y(_0710_),
    .A(_0034_),
    .B(_0318_));
 sg13g2_xor2_1 _2697_ (.B(_0318_),
    .A(_0034_),
    .X(_0711_));
 sg13g2_o21ai_1 _2698_ (.B1(_0303_),
    .Y(_0712_),
    .A1(_0332_),
    .A2(_0711_));
 sg13g2_nor2b_1 _2699_ (.A(\illness_sys.illness[4] ),
    .B_N(_0322_),
    .Y(_0713_));
 sg13g2_xnor2_1 _2700_ (.Y(_0714_),
    .A(\illness_sys.illness[4] ),
    .B(_0322_));
 sg13g2_nand3_1 _2701_ (.B(_0302_),
    .C(_0714_),
    .A(net472),
    .Y(_0715_));
 sg13g2_nand3_1 _2702_ (.B(_0712_),
    .C(_0715_),
    .A(_0709_),
    .Y(_0716_));
 sg13g2_o21ai_1 _2703_ (.B1(_0689_),
    .Y(_0193_),
    .A1(net423),
    .A2(_0716_));
 sg13g2_nor2b_1 _2704_ (.A(_0034_),
    .B_N(_0306_),
    .Y(_0717_));
 sg13g2_a22oi_1 _2705_ (.Y(_0718_),
    .B1(_0717_),
    .B2(_0312_),
    .A2(_0713_),
    .A1(net470));
 sg13g2_a21oi_1 _2706_ (.A1(_0304_),
    .A2(_0718_),
    .Y(_0719_),
    .B1(net423));
 sg13g2_xor2_1 _2707_ (.B(_0717_),
    .A(\illness_sys.illness[5] ),
    .X(_0720_));
 sg13g2_xor2_1 _2708_ (.B(_0710_),
    .A(\illness_sys.illness[5] ),
    .X(_0721_));
 sg13g2_o21ai_1 _2709_ (.B1(net472),
    .Y(_0722_),
    .A1(_0332_),
    .A2(_0721_));
 sg13g2_o21ai_1 _2710_ (.B1(_0722_),
    .Y(_0723_),
    .A1(_0328_),
    .A2(_0720_));
 sg13g2_nand2b_1 _2711_ (.Y(_0724_),
    .B(net443),
    .A_N(_0723_));
 sg13g2_o21ai_1 _2712_ (.B1(_0724_),
    .Y(_0725_),
    .A1(\illness_sys.illness[5] ),
    .A2(net443));
 sg13g2_mux2_1 _2713_ (.A0(\illness_sys.illness[5] ),
    .A1(_0725_),
    .S(_0719_),
    .X(_0194_));
 sg13g2_xnor2_1 _2714_ (.Y(_0726_),
    .A(\illness_sys.illness[6] ),
    .B(_0323_));
 sg13g2_xor2_1 _2715_ (.B(_0319_),
    .A(_0035_),
    .X(_0727_));
 sg13g2_o21ai_1 _2716_ (.B1(net443),
    .Y(_0728_),
    .A1(_0332_),
    .A2(_0727_));
 sg13g2_o21ai_1 _2717_ (.B1(net470),
    .Y(_0729_),
    .A1(net442),
    .A2(_0726_));
 sg13g2_inv_1 _2718_ (.Y(_0730_),
    .A(_0729_));
 sg13g2_xor2_1 _2719_ (.B(_0307_),
    .A(\illness_sys.illness[6] ),
    .X(_0731_));
 sg13g2_nor2_1 _2720_ (.A(_0307_),
    .B(_0311_),
    .Y(_0732_));
 sg13g2_xnor2_1 _2721_ (.Y(_0733_),
    .A(\illness_sys.illness[6] ),
    .B(_0732_));
 sg13g2_a221oi_1 _2722_ (.B2(_0304_),
    .C1(net470),
    .B1(_0733_),
    .A1(_0690_),
    .Y(_0734_),
    .A2(_0731_));
 sg13g2_a21oi_1 _2723_ (.A1(_0728_),
    .A2(_0730_),
    .Y(_0735_),
    .B1(_0734_));
 sg13g2_o21ai_1 _2724_ (.B1(_0689_),
    .Y(_0195_),
    .A1(net423),
    .A2(_0735_));
 sg13g2_nand2_1 _2725_ (.Y(_0736_),
    .A(_0085_),
    .B(net423));
 sg13g2_nor2_1 _2726_ (.A(_0035_),
    .B(_0307_),
    .Y(_0737_));
 sg13g2_o21ai_1 _2727_ (.B1(_0737_),
    .Y(_0738_),
    .A1(net442),
    .A2(_0310_));
 sg13g2_xor2_1 _2728_ (.B(_0738_),
    .A(\illness_sys.illness[7] ),
    .X(_0739_));
 sg13g2_o21ai_1 _2729_ (.B1(\illness_sys.illness[7] ),
    .Y(_0740_),
    .A1(\illness_sys.illness[6] ),
    .A2(_0323_));
 sg13g2_nor2_1 _2730_ (.A(net442),
    .B(_0324_),
    .Y(_0741_));
 sg13g2_nand3_1 _2731_ (.B(_0035_),
    .C(_0319_),
    .A(\illness_sys.illness[7] ),
    .Y(_0742_));
 sg13g2_a21oi_1 _2732_ (.A1(_0035_),
    .A2(_0319_),
    .Y(_0743_),
    .B1(\illness_sys.illness[7] ));
 sg13g2_nor2_1 _2733_ (.A(_0332_),
    .B(_0743_),
    .Y(_0744_));
 sg13g2_a21oi_1 _2734_ (.A1(_0742_),
    .A2(_0744_),
    .Y(_0745_),
    .B1(_0302_));
 sg13g2_a21oi_1 _2735_ (.A1(_0740_),
    .A2(_0741_),
    .Y(_0746_),
    .B1(_0745_));
 sg13g2_nand2b_1 _2736_ (.Y(_0747_),
    .B(_0335_),
    .A_N(net423));
 sg13g2_a21oi_1 _2737_ (.A1(net471),
    .A2(_0746_),
    .Y(_0748_),
    .B1(_0747_));
 sg13g2_o21ai_1 _2738_ (.B1(_0748_),
    .Y(_0749_),
    .A1(net471),
    .A2(_0739_));
 sg13g2_nand2_1 _2739_ (.Y(_0196_),
    .A(_0736_),
    .B(_0749_));
 sg13g2_and2_1 _2740_ (.A(_0006_),
    .B(_0309_),
    .X(_0750_));
 sg13g2_a21oi_1 _2741_ (.A1(net443),
    .A2(_0750_),
    .Y(_0751_),
    .B1(net471));
 sg13g2_o21ai_1 _2742_ (.B1(\illness_sys.illness[8] ),
    .Y(_0752_),
    .A1(_0741_),
    .A2(_0751_));
 sg13g2_nor2_1 _2743_ (.A(_0006_),
    .B(_0320_),
    .Y(_0753_));
 sg13g2_a21oi_1 _2744_ (.A1(_0006_),
    .A2(_0320_),
    .Y(_0754_),
    .B1(_0332_));
 sg13g2_nand3b_1 _2745_ (.B(_0754_),
    .C(_0303_),
    .Y(_0755_),
    .A_N(_0753_));
 sg13g2_o21ai_1 _2746_ (.B1(_0311_),
    .Y(_0756_),
    .A1(_0301_),
    .A2(_0302_));
 sg13g2_nand3_1 _2747_ (.B(_0309_),
    .C(_0756_),
    .A(_0299_),
    .Y(_0757_));
 sg13g2_nand3_1 _2748_ (.B(_0755_),
    .C(_0757_),
    .A(_0752_),
    .Y(_0197_));
 sg13g2_o21ai_1 _2749_ (.B1(_0852_),
    .Y(_0758_),
    .A1(_0343_),
    .A2(_0373_));
 sg13g2_xor2_1 _2750_ (.B(net469),
    .A(\development_stage_sys.development_stage_level[1] ),
    .X(_0759_));
 sg13g2_xnor2_1 _2751_ (.Y(_0760_),
    .A(net422),
    .B(_0759_));
 sg13g2_a22oi_1 _2752_ (.Y(_0761_),
    .B1(_0760_),
    .B2(net440),
    .A2(_0758_),
    .A1(_0382_));
 sg13g2_nand2_1 _2753_ (.Y(_0762_),
    .A(net412),
    .B(_0761_));
 sg13g2_o21ai_1 _2754_ (.B1(_0762_),
    .Y(_0198_),
    .A1(_0852_),
    .A2(net412));
 sg13g2_a21oi_1 _2755_ (.A1(net469),
    .A2(_0360_),
    .Y(_0763_),
    .B1(_0371_));
 sg13g2_nor2_1 _2756_ (.A(_0346_),
    .B(_0360_),
    .Y(_0764_));
 sg13g2_nand2b_1 _2757_ (.Y(_0765_),
    .B(_0381_),
    .A_N(_0764_));
 sg13g2_o21ai_1 _2758_ (.B1(_0765_),
    .Y(_0766_),
    .A1(net441),
    .A2(_0763_));
 sg13g2_o21ai_1 _2759_ (.B1(\development_stage_sys.development_stage_level[2] ),
    .Y(_0767_),
    .A1(net460),
    .A2(net469));
 sg13g2_nand2b_1 _2760_ (.Y(_0768_),
    .B(_0767_),
    .A_N(_0351_));
 sg13g2_o21ai_1 _2761_ (.B1(net422),
    .Y(_0769_),
    .A1(_0374_),
    .A2(_0764_));
 sg13g2_a21oi_1 _2762_ (.A1(net440),
    .A2(_0768_),
    .Y(_0770_),
    .B1(_0769_));
 sg13g2_a21oi_1 _2763_ (.A1(_0343_),
    .A2(_0766_),
    .Y(_0771_),
    .B1(_0770_));
 sg13g2_mux2_1 _2764_ (.A0(\development_stage_sys.development_stage_level[2] ),
    .A1(_0771_),
    .S(net412),
    .X(_0199_));
 sg13g2_a21o_1 _2765_ (.A2(_0360_),
    .A1(net469),
    .B1(net459),
    .X(_0772_));
 sg13g2_nand3_1 _2766_ (.B(_0363_),
    .C(_0772_),
    .A(net439),
    .Y(_0773_));
 sg13g2_nor2_1 _2767_ (.A(net459),
    .B(_0360_),
    .Y(_0774_));
 sg13g2_nor3_1 _2768_ (.A(_0007_),
    .B(_0359_),
    .C(_0365_),
    .Y(_0775_));
 sg13g2_nor2_1 _2769_ (.A(_0362_),
    .B(_0775_),
    .Y(_0776_));
 sg13g2_nor3_1 _2770_ (.A(net439),
    .B(_0774_),
    .C(_0776_),
    .Y(_0777_));
 sg13g2_nor2_1 _2771_ (.A(net422),
    .B(_0777_),
    .Y(_0778_));
 sg13g2_xnor2_1 _2772_ (.Y(_0779_),
    .A(_0037_),
    .B(_0346_));
 sg13g2_nand3_1 _2773_ (.B(_0373_),
    .C(_0779_),
    .A(net441),
    .Y(_0780_));
 sg13g2_nor2b_1 _2774_ (.A(net459),
    .B_N(_0351_),
    .Y(_0781_));
 sg13g2_xor2_1 _2775_ (.B(_0351_),
    .A(net459),
    .X(_0782_));
 sg13g2_a21oi_1 _2776_ (.A1(net440),
    .A2(_0782_),
    .Y(_0783_),
    .B1(_0343_));
 sg13g2_a22oi_1 _2777_ (.Y(_0784_),
    .B1(_0780_),
    .B2(_0783_),
    .A2(_0778_),
    .A1(_0773_));
 sg13g2_mux2_1 _2778_ (.A0(net459),
    .A1(_0784_),
    .S(net412),
    .X(_0200_));
 sg13g2_nand2b_1 _2779_ (.Y(_0785_),
    .B(_0360_),
    .A_N(_0037_));
 sg13g2_xnor2_1 _2780_ (.Y(_0786_),
    .A(_0854_),
    .B(_0785_));
 sg13g2_xnor2_1 _2781_ (.Y(_0787_),
    .A(_0854_),
    .B(_0363_));
 sg13g2_a22oi_1 _2782_ (.Y(_0788_),
    .B1(_0787_),
    .B2(net439),
    .A2(_0786_),
    .A1(_0381_));
 sg13g2_or2_1 _2783_ (.X(_0789_),
    .B(_0788_),
    .A(net422));
 sg13g2_xor2_1 _2784_ (.B(_0347_),
    .A(_0038_),
    .X(_0790_));
 sg13g2_xnor2_1 _2785_ (.Y(_0791_),
    .A(_0854_),
    .B(_0781_));
 sg13g2_a21oi_1 _2786_ (.A1(net439),
    .A2(_0791_),
    .Y(_0792_),
    .B1(_0343_));
 sg13g2_o21ai_1 _2787_ (.B1(_0792_),
    .Y(_0793_),
    .A1(_0374_),
    .A2(_0790_));
 sg13g2_nand3_1 _2788_ (.B(_0789_),
    .C(_0793_),
    .A(net412),
    .Y(_0794_));
 sg13g2_o21ai_1 _2789_ (.B1(_0794_),
    .Y(_0201_),
    .A1(_0854_),
    .A2(net412));
 sg13g2_xor2_1 _2790_ (.B(_0379_),
    .A(\development_stage_sys.development_stage_level[5] ),
    .X(_0795_));
 sg13g2_nor2_1 _2791_ (.A(_0038_),
    .B(_0363_),
    .Y(_0796_));
 sg13g2_xnor2_1 _2792_ (.Y(_0797_),
    .A(\development_stage_sys.development_stage_level[5] ),
    .B(_0796_));
 sg13g2_a22oi_1 _2793_ (.Y(_0798_),
    .B1(_0797_),
    .B2(net439),
    .A2(_0795_),
    .A1(_0381_));
 sg13g2_xnor2_1 _2794_ (.Y(_0799_),
    .A(_0039_),
    .B(_0348_));
 sg13g2_o21ai_1 _2795_ (.B1(\development_stage_sys.development_stage_level[5] ),
    .Y(_0800_),
    .A1(net469),
    .A2(_0348_));
 sg13g2_a21o_1 _2796_ (.A2(_0800_),
    .A1(_0352_),
    .B1(net441),
    .X(_0801_));
 sg13g2_o21ai_1 _2797_ (.B1(_0801_),
    .Y(_0802_),
    .A1(_0374_),
    .A2(_0799_));
 sg13g2_mux2_1 _2798_ (.A0(_0798_),
    .A1(_0802_),
    .S(net422),
    .X(_0803_));
 sg13g2_mux2_1 _2799_ (.A0(\development_stage_sys.development_stage_level[5] ),
    .A1(_0803_),
    .S(net412),
    .X(_0202_));
 sg13g2_xnor2_1 _2800_ (.Y(_0804_),
    .A(_0040_),
    .B(_0350_));
 sg13g2_xnor2_1 _2801_ (.Y(_0805_),
    .A(net458),
    .B(_0352_));
 sg13g2_a21oi_1 _2802_ (.A1(net439),
    .A2(_0805_),
    .Y(_0806_),
    .B1(_0343_));
 sg13g2_o21ai_1 _2803_ (.B1(_0806_),
    .Y(_0807_),
    .A1(_0374_),
    .A2(_0804_));
 sg13g2_nor2_1 _2804_ (.A(_0039_),
    .B(_0379_),
    .Y(_0808_));
 sg13g2_xnor2_1 _2805_ (.Y(_0809_),
    .A(net458),
    .B(_0808_));
 sg13g2_xor2_1 _2806_ (.B(_0364_),
    .A(net458),
    .X(_0810_));
 sg13g2_a22oi_1 _2807_ (.Y(_0811_),
    .B1(_0810_),
    .B2(net439),
    .A2(_0809_),
    .A1(_0381_));
 sg13g2_o21ai_1 _2808_ (.B1(_0807_),
    .Y(_0812_),
    .A1(_0342_),
    .A2(_0811_));
 sg13g2_nor2_1 _2809_ (.A(net458),
    .B(net413),
    .Y(_0813_));
 sg13g2_a21oi_1 _2810_ (.A1(net412),
    .A2(_0812_),
    .Y(_0203_),
    .B1(_0813_));
 sg13g2_xnor2_1 _2811_ (.Y(_0814_),
    .A(_0041_),
    .B(_0353_));
 sg13g2_nand3_1 _2812_ (.B(_0373_),
    .C(_0814_),
    .A(_0344_),
    .Y(_0815_));
 sg13g2_nand3_1 _2813_ (.B(net440),
    .C(_0355_),
    .A(net457),
    .Y(_0816_));
 sg13g2_nand4_1 _2814_ (.B(_0356_),
    .C(_0815_),
    .A(net422),
    .Y(_0817_),
    .D(_0816_));
 sg13g2_nor2_1 _2815_ (.A(_0040_),
    .B(_0364_),
    .Y(_0818_));
 sg13g2_xnor2_1 _2816_ (.Y(_0819_),
    .A(_0855_),
    .B(_0818_));
 sg13g2_nand4_1 _2817_ (.B(\development_stage_sys.development_stage_level[4] ),
    .C(net458),
    .A(\development_stage_sys.development_stage_level[5] ),
    .Y(_0820_),
    .D(_0361_));
 sg13g2_a21oi_1 _2818_ (.A1(net457),
    .A2(_0007_),
    .Y(_0821_),
    .B1(_0820_));
 sg13g2_a21oi_1 _2819_ (.A1(net457),
    .A2(_0820_),
    .Y(_0822_),
    .B1(_0821_));
 sg13g2_a21oi_1 _2820_ (.A1(_0345_),
    .A2(_0819_),
    .Y(_0823_),
    .B1(net422));
 sg13g2_o21ai_1 _2821_ (.B1(_0823_),
    .Y(_0824_),
    .A1(net440),
    .A2(_0822_));
 sg13g2_nand3_1 _2822_ (.B(_0817_),
    .C(_0824_),
    .A(net413),
    .Y(_0825_));
 sg13g2_o21ai_1 _2823_ (.B1(_0825_),
    .Y(_0204_),
    .A1(_0855_),
    .A2(net413));
 sg13g2_xnor2_1 _2824_ (.Y(_0826_),
    .A(_0007_),
    .B(_0354_));
 sg13g2_nand3_1 _2825_ (.B(_0373_),
    .C(_0826_),
    .A(net441),
    .Y(_0827_));
 sg13g2_o21ai_1 _2826_ (.B1(\actions.development_stage[1] ),
    .Y(_0828_),
    .A1(net457),
    .A2(_0355_));
 sg13g2_o21ai_1 _2827_ (.B1(_0827_),
    .Y(_0829_),
    .A1(net441),
    .A2(_0828_));
 sg13g2_nor2_1 _2828_ (.A(_0041_),
    .B(_0820_),
    .Y(_0830_));
 sg13g2_xor2_1 _2829_ (.B(_0830_),
    .A(\actions.development_stage[1] ),
    .X(_0831_));
 sg13g2_o21ai_1 _2830_ (.B1(net441),
    .Y(_0832_),
    .A1(_0380_),
    .A2(_0831_));
 sg13g2_o21ai_1 _2831_ (.B1(net440),
    .Y(_0833_),
    .A1(\actions.development_stage[1] ),
    .A2(_0366_));
 sg13g2_o21ai_1 _2832_ (.B1(_0343_),
    .Y(_0834_),
    .A1(_0367_),
    .A2(_0833_));
 sg13g2_nand2b_1 _2833_ (.Y(_0835_),
    .B(_0832_),
    .A_N(_0834_));
 sg13g2_o21ai_1 _2834_ (.B1(_0835_),
    .Y(_0836_),
    .A1(_0358_),
    .A2(_0829_));
 sg13g2_nor2_1 _2835_ (.A(\actions.development_stage[1] ),
    .B(net413),
    .Y(_0837_));
 sg13g2_a21oi_1 _2836_ (.A1(net413),
    .A2(_0836_),
    .Y(_0205_),
    .B1(_0837_));
 sg13g2_dfrbp_1 _2837_ (.CLK(net508),
    .RESET_B(net524),
    .D(\emotions.CORT[0] ),
    .Q_N(_1462_),
    .Q(\neurotransmitter.cortisol_system.cortisol_regulator.CORT[0] ));
 sg13g2_dfrbp_1 _2838_ (.CLK(net508),
    .RESET_B(net539),
    .D(net462),
    .Q_N(_1463_),
    .Q(\neurotransmitter.cortisol_system.cortisol_regulator.CORT[1] ));
 sg13g2_dfrbp_1 _2839_ (.CLK(net513),
    .RESET_B(net538),
    .D(net491),
    .Q_N(_1464_),
    .Q(\neurotransmitter.cortisol_system.cortisol_regulator.DOP[0] ));
 sg13g2_dfrbp_1 _2840_ (.CLK(net514),
    .RESET_B(net538),
    .D(\emotions.DOP[1] ),
    .Q_N(_1465_),
    .Q(\neurotransmitter.cortisol_system.cortisol_regulator.DOP[1] ));
 sg13g2_dfrbp_1 _2841_ (.CLK(net514),
    .RESET_B(net538),
    .D(\emotions.GABA[0] ),
    .Q_N(_1466_),
    .Q(\neurotransmitter.cortisol_system.cortisol_regulator.GABA[0] ));
 sg13g2_dfrbp_1 _2842_ (.CLK(net514),
    .RESET_B(net538),
    .D(\emotions.GABA[1] ),
    .Q_N(_1467_),
    .Q(\neurotransmitter.cortisol_system.cortisol_regulator.GABA[1] ));
 sg13g2_dfrbp_1 _2843_ (.CLK(net508),
    .RESET_B(net524),
    .D(\emotions.NE[0] ),
    .Q_N(_1468_),
    .Q(\neurotransmitter.cortisol_system.cortisol_regulator.NE[0] ));
 sg13g2_dfrbp_1 _2844_ (.CLK(net508),
    .RESET_B(net524),
    .D(net497),
    .Q_N(_1469_),
    .Q(\neurotransmitter.cortisol_system.cortisol_regulator.NE[1] ));
 sg13g2_dfrbp_1 _2845_ (.CLK(net509),
    .RESET_B(net525),
    .D(\emotions.SER[0] ),
    .Q_N(_1470_),
    .Q(\neurotransmitter.cortisol_system.cortisol_regulator.SER[0] ));
 sg13g2_dfrbp_1 _2846_ (.CLK(net514),
    .RESET_B(net539),
    .D(net482),
    .Q_N(_1471_),
    .Q(\neurotransmitter.cortisol_system.cortisol_regulator.SER[1] ));
 sg13g2_dfrbp_1 _2847_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net519),
    .D(net23),
    .Q_N(_1404_),
    .Q(\heartbeat_divider.counter[0] ));
 sg13g2_dfrbp_1 _2848_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net519),
    .D(net62),
    .Q_N(_1472_),
    .Q(\heartbeat_divider.counter[1] ));
 sg13g2_dfrbp_1 _2849_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net519),
    .D(net125),
    .Q_N(_1473_),
    .Q(\heartbeat_divider.counter[2] ));
 sg13g2_dfrbp_1 _2850_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net519),
    .D(net53),
    .Q_N(_1474_),
    .Q(\heartbeat_divider.counter[3] ));
 sg13g2_dfrbp_1 _2851_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net520),
    .D(net32),
    .Q_N(_1475_),
    .Q(\heartbeat_divider.counter[4] ));
 sg13g2_dfrbp_1 _2852_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net518),
    .D(net71),
    .Q_N(_1476_),
    .Q(\heartbeat_divider.counter[5] ));
 sg13g2_dfrbp_1 _2853_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net518),
    .D(_0062_),
    .Q_N(_1477_),
    .Q(\heartbeat_divider.counter[6] ));
 sg13g2_dfrbp_1 _2854_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net518),
    .D(net36),
    .Q_N(_1478_),
    .Q(\heartbeat_divider.counter[7] ));
 sg13g2_dfrbp_1 _2855_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net518),
    .D(net50),
    .Q_N(_1479_),
    .Q(\heartbeat_divider.counter[8] ));
 sg13g2_dfrbp_1 _2856_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net518),
    .D(_0065_),
    .Q_N(_1480_),
    .Q(\heartbeat_divider.counter[9] ));
 sg13g2_dfrbp_1 _2857_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net519),
    .D(net48),
    .Q_N(_1481_),
    .Q(\heartbeat_divider.counter[10] ));
 sg13g2_dfrbp_1 _2858_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net518),
    .D(net67),
    .Q_N(_1482_),
    .Q(\heartbeat_divider.counter[11] ));
 sg13g2_dfrbp_1 _2859_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net518),
    .D(_0055_),
    .Q_N(_1483_),
    .Q(\heartbeat_divider.counter[12] ));
 sg13g2_dfrbp_1 _2860_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net518),
    .D(_0056_),
    .Q_N(_1461_),
    .Q(\actions.clk ));
 sg13g2_dfrbp_1 _2861_ (.CLK(net507),
    .RESET_B(net522),
    .D(_0087_),
    .Q_N(_0011_),
    .Q(\neurotransmitter.norepinephrine_system.norepinephrine[0] ));
 sg13g2_dfrbp_1 _2862_ (.CLK(net507),
    .RESET_B(net522),
    .D(_0088_),
    .Q_N(_1460_),
    .Q(\neurotransmitter.norepinephrine_system.norepinephrine[1] ));
 sg13g2_dfrbp_1 _2863_ (.CLK(net505),
    .RESET_B(net524),
    .D(_0089_),
    .Q_N(_0012_),
    .Q(\neurotransmitter.norepinephrine_system.norepinephrine[2] ));
 sg13g2_dfrbp_1 _2864_ (.CLK(net508),
    .RESET_B(net524),
    .D(_0090_),
    .Q_N(_1459_),
    .Q(\neurotransmitter.norepinephrine_system.norepinephrine[3] ));
 sg13g2_dfrbp_1 _2865_ (.CLK(net505),
    .RESET_B(net524),
    .D(_0091_),
    .Q_N(_0013_),
    .Q(\emotions.NE[0] ));
 sg13g2_dfrbp_1 _2866_ (.CLK(net505),
    .RESET_B(net524),
    .D(_0092_),
    .Q_N(_1458_),
    .Q(\emotions.NE[1] ));
 sg13g2_dfrbp_1 _2867_ (.CLK(net516),
    .RESET_B(net543),
    .D(_0093_),
    .Q_N(_0014_),
    .Q(\neurotransmitter.gaba_system.gaba[0] ));
 sg13g2_dfrbp_1 _2868_ (.CLK(net516),
    .RESET_B(net542),
    .D(_0094_),
    .Q_N(_1457_),
    .Q(\neurotransmitter.gaba_system.gaba[1] ));
 sg13g2_dfrbp_1 _2869_ (.CLK(net516),
    .RESET_B(net542),
    .D(_0095_),
    .Q_N(_0015_),
    .Q(\neurotransmitter.gaba_system.gaba[2] ));
 sg13g2_dfrbp_1 _2870_ (.CLK(net516),
    .RESET_B(net542),
    .D(_0096_),
    .Q_N(_1456_),
    .Q(\neurotransmitter.gaba_system.gaba[3] ));
 sg13g2_dfrbp_1 _2871_ (.CLK(net515),
    .RESET_B(net542),
    .D(_0097_),
    .Q_N(_0016_),
    .Q(\neurotransmitter.gaba_system.gaba[4] ));
 sg13g2_dfrbp_1 _2872_ (.CLK(net515),
    .RESET_B(net542),
    .D(_0098_),
    .Q_N(\emotions.GABA[0] ),
    .Q(_0066_));
 sg13g2_dfrbp_1 _2873_ (.CLK(net516),
    .RESET_B(net542),
    .D(_0099_),
    .Q_N(\emotions.GABA[1] ),
    .Q(_0067_));
 sg13g2_dfrbp_1 _2874_ (.CLK(net513),
    .RESET_B(net539),
    .D(_0100_),
    .Q_N(_0017_),
    .Q(\neurotransmitter.dopamine_system.dopamine[0] ));
 sg13g2_dfrbp_1 _2875_ (.CLK(net513),
    .RESET_B(net542),
    .D(_0101_),
    .Q_N(_1455_),
    .Q(\neurotransmitter.dopamine_system.dopamine[1] ));
 sg13g2_dfrbp_1 _2876_ (.CLK(net513),
    .RESET_B(net538),
    .D(_0102_),
    .Q_N(_0018_),
    .Q(\neurotransmitter.dopamine_system.dopamine[2] ));
 sg13g2_dfrbp_1 _2877_ (.CLK(net513),
    .RESET_B(net538),
    .D(_0103_),
    .Q_N(_1454_),
    .Q(\neurotransmitter.dopamine_system.dopamine[3] ));
 sg13g2_dfrbp_1 _2878_ (.CLK(net513),
    .RESET_B(net538),
    .D(_0104_),
    .Q_N(_0019_),
    .Q(\neurotransmitter.dopamine_system.dopamine[4] ));
 sg13g2_dfrbp_1 _2879_ (.CLK(net513),
    .RESET_B(net538),
    .D(_0105_),
    .Q_N(_1453_),
    .Q(\emotions.DOP[0] ));
 sg13g2_dfrbp_1 _2880_ (.CLK(net513),
    .RESET_B(net539),
    .D(_0106_),
    .Q_N(\emotions.DOP[1] ),
    .Q(_0068_));
 sg13g2_dfrbp_1 _2881_ (.CLK(net512),
    .RESET_B(net530),
    .D(_0107_),
    .Q_N(_0028_),
    .Q(\nourishment.glucose[0] ));
 sg13g2_dfrbp_1 _2882_ (.CLK(net512),
    .RESET_B(net530),
    .D(_0108_),
    .Q_N(_1452_),
    .Q(\nourishment.glucose[1] ));
 sg13g2_dfrbp_1 _2883_ (.CLK(net510),
    .RESET_B(net523),
    .D(_0109_),
    .Q_N(_0020_),
    .Q(\neurotransmitter.cortisol_system.cortisol[0] ));
 sg13g2_dfrbp_1 _2884_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net532),
    .D(_0110_),
    .Q_N(_1451_),
    .Q(\talking.uart_active ));
 sg13g2_dfrbp_1 _2885_ (.CLK(net509),
    .RESET_B(net525),
    .D(_0111_),
    .Q_N(_0008_),
    .Q(\neurotransmitter.serotonin_system.serotonin[0] ));
 sg13g2_dfrbp_1 _2886_ (.CLK(net509),
    .RESET_B(net525),
    .D(_0112_),
    .Q_N(_1450_),
    .Q(\neurotransmitter.serotonin_system.serotonin[1] ));
 sg13g2_dfrbp_1 _2887_ (.CLK(net509),
    .RESET_B(net525),
    .D(_0113_),
    .Q_N(_0009_),
    .Q(\neurotransmitter.serotonin_system.serotonin[2] ));
 sg13g2_dfrbp_1 _2888_ (.CLK(net509),
    .RESET_B(net525),
    .D(_0114_),
    .Q_N(_1449_),
    .Q(\neurotransmitter.serotonin_system.serotonin[3] ));
 sg13g2_dfrbp_1 _2889_ (.CLK(net508),
    .RESET_B(net525),
    .D(_0115_),
    .Q_N(_0010_),
    .Q(\neurotransmitter.serotonin_system.serotonin[4] ));
 sg13g2_dfrbp_1 _2890_ (.CLK(net509),
    .RESET_B(net525),
    .D(_0116_),
    .Q_N(\emotions.SER[0] ),
    .Q(_0069_));
 sg13g2_dfrbp_1 _2891_ (.CLK(net508),
    .RESET_B(net525),
    .D(_0117_),
    .Q_N(\emotions.SER[1] ),
    .Q(_0070_));
 sg13g2_dfrbp_1 _2892_ (.CLK(net515),
    .RESET_B(net541),
    .D(\actions.next_action[0] ),
    .Q_N(_0045_),
    .Q(\actions.is_asleep ));
 sg13g2_dfrbp_1 _2893_ (.CLK(net511),
    .RESET_B(net541),
    .D(\actions.next_action[1] ),
    .Q_N(_1484_),
    .Q(\neurotransmitter.cortisol_system.cortisol_regulator.eat ));
 sg13g2_dfrbp_1 _2894_ (.CLK(net511),
    .RESET_B(net541),
    .D(\actions.next_action[2] ),
    .Q_N(_1448_),
    .Q(\neurotransmitter.cortisol_system.cortisol_regulator.play ));
 sg13g2_dfrbp_1 _2895_ (.CLK(net517),
    .RESET_B(net540),
    .D(_0086_),
    .Q_N(\neurotransmitter.cortisol_system.cortisol_regulator.smile ),
    .Q(_0071_));
 sg13g2_dfrbp_1 _2896_ (.CLK(net511),
    .RESET_B(net541),
    .D(\actions.next_action[4] ),
    .Q_N(_1485_),
    .Q(\neurotransmitter.cortisol_system.cortisol_regulator.babble ));
 sg13g2_dfrbp_1 _2897_ (.CLK(net511),
    .RESET_B(net540),
    .D(\actions.next_action[5] ),
    .Q_N(_1486_),
    .Q(\neurotransmitter.cortisol_system.cortisol_regulator.kick_legs ));
 sg13g2_dfrbp_1 _2898_ (.CLK(net511),
    .RESET_B(net536),
    .D(\actions.next_action[6] ),
    .Q_N(_1487_),
    .Q(\neurotransmitter.cortisol_system.cortisol_regulator.idle ));
 sg13g2_dfrbp_1 _2899_ (.CLK(net512),
    .RESET_B(net539),
    .D(\actions.next_action[7] ),
    .Q_N(_0046_),
    .Q(\development_stage_sys.dev_stage_reg.cry ));
 sg13g2_dfrbp_1 _2900_ (.CLK(net503),
    .RESET_B(net523),
    .D(_0118_),
    .Q_N(_0047_),
    .Q(\development_stage_sys.dev_stage_reg.is_ill ));
 sg13g2_dfrbp_1 _2901_ (.CLK(net503),
    .RESET_B(net521),
    .D(_0119_),
    .Q_N(_0032_),
    .Q(\illness_sys.illness[0] ));
 sg13g2_dfrbp_1 _2902_ (.CLK(net503),
    .RESET_B(net521),
    .D(_0120_),
    .Q_N(_1447_),
    .Q(\illness_sys.illness[1] ));
 sg13g2_dfrbp_1 _2903_ (.CLK(net506),
    .RESET_B(net520),
    .D(_0121_),
    .Q_N(_0036_),
    .Q(\development_stage_sys.development_stage_level[0] ));
 sg13g2_dfrbp_1 _2904_ (.CLK(net504),
    .RESET_B(net519),
    .D(_0000_),
    .Q_N(_1488_),
    .Q(\counter_.count[0] ));
 sg13g2_dfrbp_1 _2905_ (.CLK(net504),
    .RESET_B(net527),
    .D(_0001_),
    .Q_N(_1489_),
    .Q(\counter_.count[1] ));
 sg13g2_dfrbp_1 _2906_ (.CLK(net512),
    .RESET_B(net527),
    .D(_0002_),
    .Q_N(_1490_),
    .Q(\counter_.count[2] ));
 sg13g2_dfrbp_1 _2907_ (.CLK(net504),
    .RESET_B(net527),
    .D(_0003_),
    .Q_N(_1491_),
    .Q(\counter_.count[3] ));
 sg13g2_dfrbp_1 _2908_ (.CLK(_0049_),
    .RESET_B(net527),
    .D(_0004_),
    .Q_N(_0004_),
    .Q(\speech_planner_.variant_bit ));
 sg13g2_dfrbp_1 _2909_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net529),
    .D(_0122_),
    .Q_N(_1446_),
    .Q(\talking.address_reg[5] ));
 sg13g2_dfrbp_1 _2910_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net530),
    .D(_0123_),
    .Q_N(_1445_),
    .Q(\talking.address_reg[6] ));
 sg13g2_dfrbp_1 _2911_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net530),
    .D(_0124_),
    .Q_N(_1444_),
    .Q(\talking.address_reg[7] ));
 sg13g2_dfrbp_1 _2912_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net531),
    .D(_0125_),
    .Q_N(_1443_),
    .Q(\talking.address_reg[8] ));
 sg13g2_dfrbp_1 _2913_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net536),
    .D(_0126_),
    .Q_N(_1442_),
    .Q(\talking.address_reg[9] ));
 sg13g2_dfrbp_1 _2914_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net536),
    .D(_0127_),
    .Q_N(_1441_),
    .Q(\talking.address_reg[10] ));
 sg13g2_dfrbp_1 _2915_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net529),
    .D(_0128_),
    .Q_N(_1440_),
    .Q(\talking.address_reg[11] ));
 sg13g2_dfrbp_1 _2916_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net529),
    .D(_0129_),
    .Q_N(_1439_),
    .Q(\talking.address_reg[12] ));
 sg13g2_dfrbp_1 _2917_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net529),
    .D(net81),
    .Q_N(_1438_),
    .Q(\talking.address_reg[13] ));
 sg13g2_dfrbp_1 _2918_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net529),
    .D(net75),
    .Q_N(_1437_),
    .Q(\talking.address_reg[14] ));
 sg13g2_dfrbp_1 _2919_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net529),
    .D(net78),
    .Q_N(_1436_),
    .Q(\talking.address_reg[15] ));
 sg13g2_dfrbp_1 _2920_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net527),
    .D(_0133_),
    .Q_N(_1435_),
    .Q(\talking.byte_count[0] ));
 sg13g2_dfrbp_1 _2921_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net527),
    .D(_0134_),
    .Q_N(_1434_),
    .Q(\talking.byte_count[1] ));
 sg13g2_dfrbp_1 _2922_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net527),
    .D(net118),
    .Q_N(_0042_),
    .Q(\talking.byte_count[2] ));
 sg13g2_dfrbp_1 _2923_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net528),
    .D(net92),
    .Q_N(_0043_),
    .Q(\talking.byte_count[3] ));
 sg13g2_dfrbp_1 _2924_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net528),
    .D(net89),
    .Q_N(_0044_),
    .Q(\talking.byte_count[4] ));
 sg13g2_dfrbp_1 _2925_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net528),
    .D(net94),
    .Q_N(_0051_),
    .Q(\talking.byte_count[5] ));
 sg13g2_dfrbp_1 _2926_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net533),
    .D(net26),
    .Q_N(_0005_),
    .Q(spi_sck));
 sg13g2_dfrbp_1 _2927_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net532),
    .D(_0140_),
    .Q_N(_1433_),
    .Q(\talking.spi_bit_count[0] ));
 sg13g2_dfrbp_1 _2928_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net532),
    .D(net65),
    .Q_N(_1432_),
    .Q(\talking.spi_bit_count[1] ));
 sg13g2_dfrbp_1 _2929_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net532),
    .D(_0142_),
    .Q_N(_1431_),
    .Q(\talking.spi_bit_count[2] ));
 sg13g2_dfrbp_1 _2930_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net532),
    .D(net98),
    .Q_N(_0050_),
    .Q(\talking.spi_bit_count[3] ));
 sg13g2_dfrbp_1 _2931_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net528),
    .D(_0144_),
    .Q_N(_1430_),
    .Q(\talking.skip_address_bytes[0] ));
 sg13g2_dfrbp_1 _2932_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net528),
    .D(_0145_),
    .Q_N(\talking.skip_address_bytes[1] ),
    .Q(_0072_));
 sg13g2_dfrbp_1 _2933_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net535),
    .D(net112),
    .Q_N(_1429_),
    .Q(\talking.spi_shift_reg[0] ));
 sg13g2_dfrbp_1 _2934_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net536),
    .D(net110),
    .Q_N(_1428_),
    .Q(\talking.spi_shift_reg[1] ));
 sg13g2_dfrbp_1 _2935_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net537),
    .D(net83),
    .Q_N(_1427_),
    .Q(\talking.spi_shift_reg[2] ));
 sg13g2_dfrbp_1 _2936_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net536),
    .D(net106),
    .Q_N(_1426_),
    .Q(\talking.spi_shift_reg[3] ));
 sg13g2_dfrbp_1 _2937_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net536),
    .D(net101),
    .Q_N(_1425_),
    .Q(\talking.spi_shift_reg[4] ));
 sg13g2_dfrbp_1 _2938_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net536),
    .D(net85),
    .Q_N(_1424_),
    .Q(\talking.spi_shift_reg[5] ));
 sg13g2_dfrbp_1 _2939_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net536),
    .D(_0152_),
    .Q_N(_1423_),
    .Q(\talking.spi_shift_reg[6] ));
 sg13g2_dfrbp_1 _2940_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net533),
    .D(net58),
    .Q_N(_1422_),
    .Q(spi_mosi));
 sg13g2_dfrbp_1 _2941_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net532),
    .D(net60),
    .Q_N(\talking.uart_shift_reg[0] ),
    .Q(_0073_));
 sg13g2_dfrbp_1 _2942_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net535),
    .D(net44),
    .Q_N(\talking.uart_shift_reg[1] ),
    .Q(_0074_));
 sg13g2_dfrbp_1 _2943_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net535),
    .D(net30),
    .Q_N(\talking.uart_shift_reg[2] ),
    .Q(_0075_));
 sg13g2_dfrbp_1 _2944_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net535),
    .D(net38),
    .Q_N(\talking.uart_shift_reg[3] ),
    .Q(_0076_));
 sg13g2_dfrbp_1 _2945_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net535),
    .D(net28),
    .Q_N(\talking.uart_shift_reg[4] ),
    .Q(_0077_));
 sg13g2_dfrbp_1 _2946_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net535),
    .D(net69),
    .Q_N(\talking.uart_shift_reg[5] ),
    .Q(_0078_));
 sg13g2_dfrbp_1 _2947_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net535),
    .D(net46),
    .Q_N(\talking.uart_shift_reg[6] ),
    .Q(_0079_));
 sg13g2_dfrbp_1 _2948_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net535),
    .D(net42),
    .Q_N(\talking.uart_shift_reg[7] ),
    .Q(_0080_));
 sg13g2_dfrbp_1 _2949_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net533),
    .D(net40),
    .Q_N(\talking.uart_shift_reg[8] ),
    .Q(_0081_));
 sg13g2_dfrbp_1 _2950_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net533),
    .D(net55),
    .Q_N(\talking.uart_shift_reg[9] ),
    .Q(_0082_));
 sg13g2_dfrbp_1 _2951_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net527),
    .D(_0164_),
    .Q_N(_1421_),
    .Q(\talking.state[0] ));
 sg13g2_dfrbp_1 _2952_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net528),
    .D(_0165_),
    .Q_N(_1420_),
    .Q(\talking.state[1] ));
 sg13g2_dfrbp_1 _2953_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net534),
    .D(_0166_),
    .Q_N(_0048_),
    .Q(\talking.state[2] ));
 sg13g2_dfrbp_1 _2954_ (.CLK(net515),
    .RESET_B(net541),
    .D(_0167_),
    .Q_N(_0024_),
    .Q(\vital_energy_sys.vital_energy[0] ));
 sg13g2_dfrbp_1 _2955_ (.CLK(net515),
    .RESET_B(net542),
    .D(_0168_),
    .Q_N(_1419_),
    .Q(\vital_energy_sys.vital_energy[1] ));
 sg13g2_dfrbp_1 _2956_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net534),
    .D(_0169_),
    .Q_N(_1418_),
    .Q(\talking.uart_bit_count[0] ));
 sg13g2_dfrbp_1 _2957_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net532),
    .D(_0170_),
    .Q_N(_1417_),
    .Q(\talking.uart_bit_count[1] ));
 sg13g2_dfrbp_1 _2958_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net532),
    .D(net73),
    .Q_N(_1416_),
    .Q(\talking.uart_bit_count[2] ));
 sg13g2_dfrbp_1 _2959_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net534),
    .D(_0172_),
    .Q_N(_1415_),
    .Q(\talking.uart_bit_count[3] ));
 sg13g2_dfrbp_1 _2960_ (.CLK(net515),
    .RESET_B(net540),
    .D(_0173_),
    .Q_N(_0025_),
    .Q(\vital_energy_sys.vital_energy[2] ));
 sg13g2_dfrbp_1 _2961_ (.CLK(net515),
    .RESET_B(net540),
    .D(_0174_),
    .Q_N(_1414_),
    .Q(\vital_energy_sys.vital_energy[3] ));
 sg13g2_dfrbp_1 _2962_ (.CLK(net515),
    .RESET_B(net540),
    .D(_0175_),
    .Q_N(_0026_),
    .Q(\vital_energy_sys.vital_energy[4] ));
 sg13g2_dfrbp_1 _2963_ (.CLK(net511),
    .RESET_B(net540),
    .D(_0176_),
    .Q_N(_1413_),
    .Q(\vital_energy_sys.vital_energy[5] ));
 sg13g2_dfrbp_1 _2964_ (.CLK(net511),
    .RESET_B(net540),
    .D(_0177_),
    .Q_N(_0027_),
    .Q(\actions.vital_energy_level[0] ));
 sg13g2_dfrbp_1 _2965_ (.CLK(net511),
    .RESET_B(net540),
    .D(_0178_),
    .Q_N(\actions.vital_energy_level[1] ),
    .Q(_0083_));
 sg13g2_dfrbp_1 _2966_ (.CLK(net512),
    .RESET_B(net530),
    .D(_0179_),
    .Q_N(_0029_),
    .Q(\nourishment.glucose[2] ));
 sg13g2_dfrbp_1 _2967_ (.CLK(net512),
    .RESET_B(net530),
    .D(_0180_),
    .Q_N(_1412_),
    .Q(\nourishment.glucose[3] ));
 sg13g2_dfrbp_1 _2968_ (.CLK(net505),
    .RESET_B(net520),
    .D(_0181_),
    .Q_N(_0030_),
    .Q(\nourishment.glucose[4] ));
 sg13g2_dfrbp_1 _2969_ (.CLK(net505),
    .RESET_B(net520),
    .D(_0182_),
    .Q_N(_1411_),
    .Q(\nourishment.glucose[5] ));
 sg13g2_dfrbp_1 _2970_ (.CLK(net512),
    .RESET_B(net539),
    .D(_0183_),
    .Q_N(_0031_),
    .Q(\nourishment.glucose[6] ));
 sg13g2_dfrbp_1 _2971_ (.CLK(net512),
    .RESET_B(net530),
    .D(_0184_),
    .Q_N(\nourishment.glucose[7] ),
    .Q(_0084_));
 sg13g2_dfrbp_1 _2972_ (.CLK(net510),
    .RESET_B(net523),
    .D(_0185_),
    .Q_N(_1410_),
    .Q(\neurotransmitter.cortisol_system.cortisol[1] ));
 sg13g2_dfrbp_1 _2973_ (.CLK(net510),
    .RESET_B(net523),
    .D(_0186_),
    .Q_N(_1409_),
    .Q(\neurotransmitter.cortisol_system.cortisol[2] ));
 sg13g2_dfrbp_1 _2974_ (.CLK(net507),
    .RESET_B(net522),
    .D(_0187_),
    .Q_N(_0021_),
    .Q(\neurotransmitter.cortisol_system.cortisol[3] ));
 sg13g2_dfrbp_1 _2975_ (.CLK(net507),
    .RESET_B(net522),
    .D(_0188_),
    .Q_N(_0022_),
    .Q(\neurotransmitter.cortisol_system.cortisol[4] ));
 sg13g2_dfrbp_1 _2976_ (.CLK(net507),
    .RESET_B(net522),
    .D(_0189_),
    .Q_N(_0023_),
    .Q(\emotions.CORT[0] ));
 sg13g2_dfrbp_1 _2977_ (.CLK(net508),
    .RESET_B(net524),
    .D(_0190_),
    .Q_N(_0052_),
    .Q(\emotions.CORT[1] ));
 sg13g2_dfrbp_1 _2978_ (.CLK(net506),
    .RESET_B(net521),
    .D(_0191_),
    .Q_N(_0033_),
    .Q(\illness_sys.illness[2] ));
 sg13g2_dfrbp_1 _2979_ (.CLK(net507),
    .RESET_B(net522),
    .D(_0192_),
    .Q_N(_1408_),
    .Q(\illness_sys.illness[3] ));
 sg13g2_dfrbp_1 _2980_ (.CLK(net507),
    .RESET_B(net522),
    .D(_0193_),
    .Q_N(_0034_),
    .Q(\illness_sys.illness[4] ));
 sg13g2_dfrbp_1 _2981_ (.CLK(net507),
    .RESET_B(net522),
    .D(_0194_),
    .Q_N(_1407_),
    .Q(\illness_sys.illness[5] ));
 sg13g2_dfrbp_1 _2982_ (.CLK(net503),
    .RESET_B(net521),
    .D(_0195_),
    .Q_N(_0035_),
    .Q(\illness_sys.illness[6] ));
 sg13g2_dfrbp_1 _2983_ (.CLK(net503),
    .RESET_B(net521),
    .D(_0196_),
    .Q_N(\illness_sys.illness[7] ),
    .Q(_0085_));
 sg13g2_dfrbp_1 _2984_ (.CLK(net503),
    .RESET_B(net521),
    .D(_0197_),
    .Q_N(_0006_),
    .Q(\illness_sys.illness[8] ));
 sg13g2_dfrbp_1 _2985_ (.CLK(net505),
    .RESET_B(net526),
    .D(_0198_),
    .Q_N(_1406_),
    .Q(\development_stage_sys.development_stage_level[1] ));
 sg13g2_dfrbp_1 _2986_ (.CLK(net503),
    .RESET_B(net526),
    .D(_0199_),
    .Q_N(_1405_),
    .Q(\development_stage_sys.development_stage_level[2] ));
 sg13g2_dfrbp_1 _2987_ (.CLK(net503),
    .RESET_B(net521),
    .D(_0200_),
    .Q_N(_0037_),
    .Q(\development_stage_sys.development_stage_level[3] ));
 sg13g2_dfrbp_1 _2988_ (.CLK(net504),
    .RESET_B(net526),
    .D(_0201_),
    .Q_N(_0038_),
    .Q(\development_stage_sys.development_stage_level[4] ));
 sg13g2_dfrbp_1 _2989_ (.CLK(net504),
    .RESET_B(net519),
    .D(_0202_),
    .Q_N(_0039_),
    .Q(\development_stage_sys.development_stage_level[5] ));
 sg13g2_dfrbp_1 _2990_ (.CLK(net505),
    .RESET_B(net520),
    .D(_0203_),
    .Q_N(_0040_),
    .Q(\development_stage_sys.development_stage_level[6] ));
 sg13g2_dfrbp_1 _2991_ (.CLK(net504),
    .RESET_B(net520),
    .D(_0204_),
    .Q_N(_0041_),
    .Q(\actions.development_stage[0] ));
 sg13g2_dfrbp_1 _2992_ (.CLK(net504),
    .RESET_B(net520),
    .D(_0205_),
    .Q_N(_0007_),
    .Q(\actions.development_stage[1] ));
 sg13g2_tiehi tt_um_moody_mimosa_19 (.L_HI(net19));
 sg13g2_tiehi tt_um_moody_mimosa_20 (.L_HI(net20));
 sg13g2_tiehi tt_um_moody_mimosa_21 (.L_HI(net21));
 sg13g2_tiehi tt_um_moody_mimosa_22 (.L_HI(net22));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_moody_mimosa_13 (.L_LO(net13));
 sg13g2_tielo tt_um_moody_mimosa_14 (.L_LO(net14));
 sg13g2_tielo tt_um_moody_mimosa_15 (.L_LO(net15));
 sg13g2_tielo tt_um_moody_mimosa_16 (.L_LO(net16));
 sg13g2_tielo tt_um_moody_mimosa_17 (.L_LO(net17));
 sg13g2_tiehi tt_um_moody_mimosa_18 (.L_HI(net18));
 sg13g2_buf_1 _3004_ (.A(spi_sck),
    .X(uio_out[3]));
 sg13g2_buf_1 _3005_ (.A(spi_cs),
    .X(uio_out[4]));
 sg13g2_buf_1 _3006_ (.A(spi_mosi),
    .X(uio_out[5]));
 sg13g2_buf_1 _3007_ (.A(\talking.uart_tx ),
    .X(uio_out[6]));
 sg13g2_buf_2 _3008_ (.A(net517),
    .X(uio_out[7]));
 sg13g2_buf_1 _3009_ (.A(net480),
    .X(uo_out[0]));
 sg13g2_buf_2 _3010_ (.A(net475),
    .X(uo_out[1]));
 sg13g2_buf_2 _3011_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.play ),
    .X(uo_out[2]));
 sg13g2_buf_2 _3012_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.smile ),
    .X(uo_out[3]));
 sg13g2_buf_2 _3013_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.babble ),
    .X(uo_out[4]));
 sg13g2_buf_2 _3014_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.kick_legs ),
    .X(uo_out[5]));
 sg13g2_buf_2 _3015_ (.A(\neurotransmitter.cortisol_system.cortisol_regulator.idle ),
    .X(uo_out[6]));
 sg13g2_buf_2 _3016_ (.A(\development_stage_sys.dev_stage_reg.cry ),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout412 (.X(net412),
    .A(_0370_));
 sg13g2_buf_2 fanout413 (.A(_0370_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_1366_),
    .X(net414));
 sg13g2_buf_1 fanout415 (.A(_1366_),
    .X(net415));
 sg13g2_buf_4 fanout416 (.X(net416),
    .A(_1059_));
 sg13g2_buf_2 fanout417 (.A(net418),
    .X(net417));
 sg13g2_buf_1 fanout418 (.A(net419),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(_0494_),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(_0480_),
    .X(net420));
 sg13g2_buf_2 fanout421 (.A(_0480_),
    .X(net421));
 sg13g2_buf_4 fanout422 (.X(net422),
    .A(_0342_));
 sg13g2_buf_4 fanout423 (.X(net423),
    .A(_0326_));
 sg13g2_buf_2 fanout424 (.A(net425),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(_0219_),
    .X(net425));
 sg13g2_buf_4 fanout426 (.X(net426),
    .A(_1352_));
 sg13g2_buf_4 fanout427 (.X(net427),
    .A(_1351_));
 sg13g2_buf_1 fanout428 (.A(_1351_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(_1243_),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(_1243_),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(_1235_),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(_1045_),
    .X(net432));
 sg13g2_buf_4 fanout433 (.X(net433),
    .A(_1041_));
 sg13g2_buf_2 fanout434 (.A(_1041_),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(net436),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(_0523_),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(net438),
    .X(net437));
 sg13g2_buf_2 fanout438 (.A(_0395_),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(net440),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(_0345_),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(_0344_),
    .X(net441));
 sg13g2_buf_4 fanout442 (.X(net442),
    .A(net443));
 sg13g2_buf_2 fanout443 (.A(_0305_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(net446),
    .X(net444));
 sg13g2_buf_1 fanout445 (.A(net446),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(_1343_),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(net448),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_1147_),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(_1142_),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(net451),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(_1381_),
    .X(net451));
 sg13g2_buf_4 fanout452 (.X(net452),
    .A(_1394_));
 sg13g2_buf_2 fanout453 (.A(_0944_),
    .X(net453));
 sg13g2_buf_4 fanout454 (.X(net454),
    .A(_0894_));
 sg13g2_buf_4 fanout455 (.X(net455),
    .A(_0841_));
 sg13g2_buf_1 fanout456 (.A(_0841_),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(\actions.development_stage[0] ),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(\development_stage_sys.development_stage_level[6] ),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(\development_stage_sys.development_stage_level[3] ),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(\development_stage_sys.development_stage_level[1] ),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(\illness_sys.illness[2] ),
    .X(net461));
 sg13g2_buf_4 fanout462 (.X(net462),
    .A(\emotions.CORT[1] ));
 sg13g2_buf_4 fanout463 (.X(net463),
    .A(\emotions.CORT[0] ));
 sg13g2_buf_2 fanout464 (.A(\neurotransmitter.cortisol_system.cortisol[1] ),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(\nourishment.glucose[7] ),
    .X(net465));
 sg13g2_buf_1 fanout466 (.A(\nourishment.glucose[7] ),
    .X(net466));
 sg13g2_buf_4 fanout467 (.X(net467),
    .A(\actions.vital_energy_level[1] ));
 sg13g2_buf_4 fanout468 (.X(net468),
    .A(\actions.vital_energy_level[0] ));
 sg13g2_buf_2 fanout469 (.A(\development_stage_sys.development_stage_level[0] ),
    .X(net469));
 sg13g2_buf_4 fanout470 (.X(net470),
    .A(net472));
 sg13g2_buf_2 fanout471 (.A(net472),
    .X(net471));
 sg13g2_buf_1 fanout472 (.A(net473),
    .X(net472));
 sg13g2_buf_4 fanout473 (.X(net473),
    .A(\development_stage_sys.dev_stage_reg.is_ill ));
 sg13g2_buf_2 fanout474 (.A(net475),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(\neurotransmitter.cortisol_system.cortisol_regulator.eat ),
    .X(net475));
 sg13g2_buf_4 fanout476 (.X(net476),
    .A(net478));
 sg13g2_buf_2 fanout477 (.A(net478),
    .X(net477));
 sg13g2_buf_4 fanout478 (.X(net478),
    .A(_0045_));
 sg13g2_buf_2 fanout479 (.A(net480),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(\actions.is_asleep ),
    .X(net480));
 sg13g2_buf_4 fanout481 (.X(net481),
    .A(\actions.is_asleep ));
 sg13g2_buf_4 fanout482 (.X(net482),
    .A(\emotions.SER[1] ));
 sg13g2_buf_2 fanout483 (.A(net484),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(\emotions.SER[0] ),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(net486),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(\neurotransmitter.serotonin_system.serotonin[4] ),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(\neurotransmitter.serotonin_system.serotonin[2] ),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(net489),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(\neurotransmitter.cortisol_system.cortisol[0] ),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(net491),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(\emotions.DOP[0] ),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(\neurotransmitter.dopamine_system.dopamine[4] ),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(\neurotransmitter.dopamine_system.dopamine[2] ),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(\neurotransmitter.gaba_system.gaba[2] ),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(net496),
    .X(net495));
 sg13g2_buf_1 fanout496 (.A(net497),
    .X(net496));
 sg13g2_buf_1 fanout497 (.A(net498),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(\emotions.NE[1] ),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(\neurotransmitter.norepinephrine_system.norepinephrine[2] ),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(net99),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(net502),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(\talking.state[0] ),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(net506),
    .X(net503));
 sg13g2_buf_4 fanout504 (.X(net504),
    .A(net505));
 sg13g2_buf_4 fanout505 (.X(net505),
    .A(net506));
 sg13g2_buf_2 fanout506 (.A(\actions.clk ),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(net510),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(net510),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(net510),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(\actions.clk ),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(net517),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(net517),
    .X(net512));
 sg13g2_buf_4 fanout513 (.X(net513),
    .A(net514));
 sg13g2_buf_2 fanout514 (.A(net517),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(net517),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(net517),
    .X(net516));
 sg13g2_buf_4 fanout517 (.X(net517),
    .A(\actions.clk ));
 sg13g2_buf_4 fanout518 (.X(net518),
    .A(net519));
 sg13g2_buf_4 fanout519 (.X(net519),
    .A(net520));
 sg13g2_buf_4 fanout520 (.X(net520),
    .A(net521));
 sg13g2_buf_4 fanout521 (.X(net521),
    .A(net526));
 sg13g2_buf_4 fanout522 (.X(net522),
    .A(net523));
 sg13g2_buf_4 fanout523 (.X(net523),
    .A(net526));
 sg13g2_buf_4 fanout524 (.X(net524),
    .A(net526));
 sg13g2_buf_4 fanout525 (.X(net525),
    .A(net526));
 sg13g2_buf_4 fanout526 (.X(net526),
    .A(net544));
 sg13g2_buf_4 fanout527 (.X(net527),
    .A(net531));
 sg13g2_buf_4 fanout528 (.X(net528),
    .A(net531));
 sg13g2_buf_4 fanout529 (.X(net529),
    .A(net530));
 sg13g2_buf_4 fanout530 (.X(net530),
    .A(net531));
 sg13g2_buf_2 fanout531 (.A(net544),
    .X(net531));
 sg13g2_buf_4 fanout532 (.X(net532),
    .A(net534));
 sg13g2_buf_2 fanout533 (.A(net534),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(net537),
    .X(net534));
 sg13g2_buf_4 fanout535 (.X(net535),
    .A(net537));
 sg13g2_buf_4 fanout536 (.X(net536),
    .A(net537));
 sg13g2_buf_2 fanout537 (.A(net544),
    .X(net537));
 sg13g2_buf_4 fanout538 (.X(net538),
    .A(net539));
 sg13g2_buf_4 fanout539 (.X(net539),
    .A(net543));
 sg13g2_buf_4 fanout540 (.X(net540),
    .A(net541));
 sg13g2_buf_4 fanout541 (.X(net541),
    .A(net543));
 sg13g2_buf_4 fanout542 (.X(net542),
    .A(net543));
 sg13g2_buf_2 fanout543 (.A(net544),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(rst_n),
    .X(net544));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_tielo tt_um_moody_mimosa_12 (.L_LO(net12));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_1404_),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0005_),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0458_),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0139_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0077_),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0158_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0075_),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0156_),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold9 (.A(\heartbeat_divider.counter[4] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0060_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0072_),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0478_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold13 (.A(\heartbeat_divider.counter[7] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0063_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0076_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0157_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0081_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0162_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0080_),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0161_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0074_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0155_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0079_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0160_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold25 (.A(\heartbeat_divider.counter[10] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0053_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold27 (.A(\heartbeat_divider.counter[8] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0064_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold29 (.A(\talking.address_reg[6] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold30 (.A(\heartbeat_divider.counter[3] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0059_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0082_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0163_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold34 (.A(\talking.address_reg[9] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold35 (.A(spi_mosi),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0153_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0073_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0154_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold39 (.A(\heartbeat_divider.counter[0] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0057_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold41 (.A(\talking.spi_bit_count[1] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0468_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0141_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold44 (.A(\heartbeat_divider.counter[11] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0054_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0078_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0159_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold48 (.A(\heartbeat_divider.counter[5] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0061_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold50 (.A(\talking.uart_bit_count[2] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0171_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold52 (.A(\talking.address_reg[14] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0131_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold54 (.A(\talking.address_reg[7] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0419_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0132_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold57 (.A(\talking.address_reg[5] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0415_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0130_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold60 (.A(\talking.spi_shift_reg[2] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0148_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold62 (.A(\talking.spi_shift_reg[5] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0151_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold64 (.A(\talking.spi_bit_count[0] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0464_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold66 (.A(\talking.byte_count[4] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0137_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold68 (.A(\talking.spi_shift_reg[6] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0043_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0136_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold71 (.A(\talking.byte_count[5] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0138_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold73 (.A(\talking.skip_address_bytes[0] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0476_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold75 (.A(\talking.spi_bit_count[2] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0143_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold77 (.A(\talking.state[1] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold78 (.A(\talking.spi_shift_reg[4] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0150_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold80 (.A(\talking.address_reg[10] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold81 (.A(\heartbeat_divider.counter[12] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold82 (.A(_1022_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold83 (.A(\talking.spi_shift_reg[3] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0149_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold85 (.A(\talking.address_reg[11] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold86 (.A(\talking.uart_bit_count[3] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold87 (.A(\talking.spi_shift_reg[1] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0147_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold89 (.A(\talking.spi_shift_reg[0] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0146_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold91 (.A(\talking.address_reg[8] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold92 (.A(\talking.address_reg[12] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold93 (.A(\talking.uart_active ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold94 (.A(_1403_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold95 (.A(\talking.byte_count[2] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0135_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold97 (.A(\talking.uart_bit_count[0] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold98 (.A(\talking.uart_bit_count[1] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold99 (.A(\heartbeat_divider.counter[6] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold100 (.A(\heartbeat_divider.counter[9] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold101 (.A(\heartbeat_divider.counter[2] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold102 (.A(_1013_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0058_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold104 (.A(\talking.byte_count[1] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold105 (.A(\talking.byte_count[0] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold106 (.A(\talking.state[2] ),
    .X(net128));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_4 FILLER_10_189 ();
 sg13g2_fill_2 FILLER_10_193 ();
 sg13g2_decap_4 FILLER_10_212 ();
 sg13g2_fill_2 FILLER_10_216 ();
 sg13g2_fill_2 FILLER_10_222 ();
 sg13g2_decap_8 FILLER_10_228 ();
 sg13g2_decap_8 FILLER_10_235 ();
 sg13g2_decap_8 FILLER_10_242 ();
 sg13g2_decap_8 FILLER_10_249 ();
 sg13g2_decap_8 FILLER_10_256 ();
 sg13g2_decap_8 FILLER_10_263 ();
 sg13g2_decap_8 FILLER_10_270 ();
 sg13g2_decap_8 FILLER_10_277 ();
 sg13g2_decap_8 FILLER_10_284 ();
 sg13g2_decap_8 FILLER_10_291 ();
 sg13g2_decap_8 FILLER_10_298 ();
 sg13g2_decap_8 FILLER_10_305 ();
 sg13g2_decap_8 FILLER_10_312 ();
 sg13g2_decap_8 FILLER_10_319 ();
 sg13g2_decap_8 FILLER_10_326 ();
 sg13g2_decap_8 FILLER_10_333 ();
 sg13g2_decap_8 FILLER_10_340 ();
 sg13g2_decap_8 FILLER_10_347 ();
 sg13g2_decap_8 FILLER_10_354 ();
 sg13g2_decap_8 FILLER_10_361 ();
 sg13g2_decap_8 FILLER_10_368 ();
 sg13g2_decap_8 FILLER_10_375 ();
 sg13g2_decap_8 FILLER_10_382 ();
 sg13g2_decap_8 FILLER_10_389 ();
 sg13g2_decap_8 FILLER_10_396 ();
 sg13g2_decap_4 FILLER_10_403 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_fill_1 FILLER_11_182 ();
 sg13g2_fill_1 FILLER_11_219 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_4 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_246 ();
 sg13g2_decap_8 FILLER_12_253 ();
 sg13g2_decap_8 FILLER_12_260 ();
 sg13g2_decap_8 FILLER_12_267 ();
 sg13g2_decap_8 FILLER_12_274 ();
 sg13g2_decap_8 FILLER_12_281 ();
 sg13g2_decap_8 FILLER_12_288 ();
 sg13g2_decap_8 FILLER_12_295 ();
 sg13g2_decap_8 FILLER_12_302 ();
 sg13g2_decap_8 FILLER_12_309 ();
 sg13g2_decap_8 FILLER_12_316 ();
 sg13g2_decap_8 FILLER_12_323 ();
 sg13g2_decap_8 FILLER_12_330 ();
 sg13g2_decap_8 FILLER_12_337 ();
 sg13g2_decap_8 FILLER_12_344 ();
 sg13g2_decap_8 FILLER_12_351 ();
 sg13g2_decap_8 FILLER_12_358 ();
 sg13g2_decap_8 FILLER_12_365 ();
 sg13g2_decap_8 FILLER_12_372 ();
 sg13g2_decap_8 FILLER_12_379 ();
 sg13g2_decap_8 FILLER_12_386 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_4 FILLER_13_168 ();
 sg13g2_decap_4 FILLER_13_196 ();
 sg13g2_fill_1 FILLER_13_213 ();
 sg13g2_fill_2 FILLER_13_223 ();
 sg13g2_fill_1 FILLER_13_225 ();
 sg13g2_fill_1 FILLER_13_236 ();
 sg13g2_decap_8 FILLER_13_246 ();
 sg13g2_decap_8 FILLER_13_253 ();
 sg13g2_decap_8 FILLER_13_260 ();
 sg13g2_decap_8 FILLER_13_267 ();
 sg13g2_decap_8 FILLER_13_274 ();
 sg13g2_decap_8 FILLER_13_281 ();
 sg13g2_decap_8 FILLER_13_288 ();
 sg13g2_decap_8 FILLER_13_295 ();
 sg13g2_decap_8 FILLER_13_302 ();
 sg13g2_decap_8 FILLER_13_309 ();
 sg13g2_decap_8 FILLER_13_316 ();
 sg13g2_decap_8 FILLER_13_323 ();
 sg13g2_decap_8 FILLER_13_330 ();
 sg13g2_decap_8 FILLER_13_337 ();
 sg13g2_decap_8 FILLER_13_344 ();
 sg13g2_decap_8 FILLER_13_351 ();
 sg13g2_decap_8 FILLER_13_358 ();
 sg13g2_decap_8 FILLER_13_365 ();
 sg13g2_decap_8 FILLER_13_372 ();
 sg13g2_decap_8 FILLER_13_379 ();
 sg13g2_decap_8 FILLER_13_386 ();
 sg13g2_decap_8 FILLER_13_393 ();
 sg13g2_decap_8 FILLER_13_400 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_4 FILLER_14_189 ();
 sg13g2_fill_1 FILLER_14_198 ();
 sg13g2_fill_2 FILLER_14_204 ();
 sg13g2_fill_1 FILLER_14_206 ();
 sg13g2_decap_4 FILLER_14_211 ();
 sg13g2_decap_4 FILLER_14_219 ();
 sg13g2_fill_1 FILLER_14_228 ();
 sg13g2_decap_8 FILLER_14_237 ();
 sg13g2_decap_8 FILLER_14_244 ();
 sg13g2_decap_8 FILLER_14_251 ();
 sg13g2_decap_8 FILLER_14_258 ();
 sg13g2_decap_8 FILLER_14_265 ();
 sg13g2_decap_8 FILLER_14_272 ();
 sg13g2_decap_8 FILLER_14_279 ();
 sg13g2_decap_8 FILLER_14_286 ();
 sg13g2_decap_8 FILLER_14_293 ();
 sg13g2_decap_8 FILLER_14_300 ();
 sg13g2_decap_8 FILLER_14_307 ();
 sg13g2_decap_8 FILLER_14_314 ();
 sg13g2_decap_8 FILLER_14_321 ();
 sg13g2_decap_8 FILLER_14_328 ();
 sg13g2_decap_8 FILLER_14_335 ();
 sg13g2_decap_8 FILLER_14_342 ();
 sg13g2_decap_8 FILLER_14_349 ();
 sg13g2_decap_8 FILLER_14_356 ();
 sg13g2_decap_8 FILLER_14_363 ();
 sg13g2_decap_8 FILLER_14_370 ();
 sg13g2_decap_8 FILLER_14_377 ();
 sg13g2_decap_8 FILLER_14_384 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_4 FILLER_15_161 ();
 sg13g2_fill_2 FILLER_15_165 ();
 sg13g2_fill_1 FILLER_15_193 ();
 sg13g2_decap_4 FILLER_15_213 ();
 sg13g2_fill_2 FILLER_15_217 ();
 sg13g2_fill_2 FILLER_15_229 ();
 sg13g2_decap_8 FILLER_15_241 ();
 sg13g2_decap_8 FILLER_15_248 ();
 sg13g2_decap_8 FILLER_15_255 ();
 sg13g2_decap_8 FILLER_15_262 ();
 sg13g2_decap_8 FILLER_15_269 ();
 sg13g2_decap_8 FILLER_15_276 ();
 sg13g2_decap_8 FILLER_15_283 ();
 sg13g2_decap_8 FILLER_15_290 ();
 sg13g2_decap_8 FILLER_15_297 ();
 sg13g2_decap_8 FILLER_15_304 ();
 sg13g2_decap_8 FILLER_15_311 ();
 sg13g2_decap_8 FILLER_15_318 ();
 sg13g2_decap_8 FILLER_15_325 ();
 sg13g2_decap_8 FILLER_15_332 ();
 sg13g2_decap_8 FILLER_15_339 ();
 sg13g2_decap_8 FILLER_15_346 ();
 sg13g2_decap_8 FILLER_15_353 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_decap_8 FILLER_15_367 ();
 sg13g2_decap_8 FILLER_15_374 ();
 sg13g2_decap_8 FILLER_15_381 ();
 sg13g2_decap_8 FILLER_15_388 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_fill_2 FILLER_16_194 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_fill_1 FILLER_17_175 ();
 sg13g2_fill_2 FILLER_17_236 ();
 sg13g2_decap_8 FILLER_17_264 ();
 sg13g2_decap_8 FILLER_17_271 ();
 sg13g2_fill_2 FILLER_17_278 ();
 sg13g2_fill_1 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_291 ();
 sg13g2_decap_8 FILLER_17_298 ();
 sg13g2_decap_8 FILLER_17_305 ();
 sg13g2_decap_8 FILLER_17_312 ();
 sg13g2_decap_8 FILLER_17_319 ();
 sg13g2_decap_8 FILLER_17_326 ();
 sg13g2_decap_8 FILLER_17_333 ();
 sg13g2_decap_8 FILLER_17_340 ();
 sg13g2_decap_8 FILLER_17_347 ();
 sg13g2_decap_8 FILLER_17_354 ();
 sg13g2_decap_8 FILLER_17_361 ();
 sg13g2_decap_8 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_fill_2 FILLER_18_154 ();
 sg13g2_fill_1 FILLER_18_156 ();
 sg13g2_decap_4 FILLER_18_191 ();
 sg13g2_fill_2 FILLER_18_199 ();
 sg13g2_fill_1 FILLER_18_201 ();
 sg13g2_decap_4 FILLER_18_218 ();
 sg13g2_fill_2 FILLER_18_222 ();
 sg13g2_fill_2 FILLER_18_234 ();
 sg13g2_decap_8 FILLER_18_253 ();
 sg13g2_decap_8 FILLER_18_260 ();
 sg13g2_decap_4 FILLER_18_267 ();
 sg13g2_fill_2 FILLER_18_296 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_4 FILLER_19_154 ();
 sg13g2_fill_2 FILLER_19_158 ();
 sg13g2_fill_2 FILLER_19_191 ();
 sg13g2_decap_4 FILLER_19_198 ();
 sg13g2_decap_8 FILLER_19_211 ();
 sg13g2_decap_8 FILLER_19_218 ();
 sg13g2_decap_4 FILLER_19_225 ();
 sg13g2_fill_2 FILLER_19_229 ();
 sg13g2_decap_4 FILLER_19_236 ();
 sg13g2_decap_4 FILLER_19_248 ();
 sg13g2_fill_1 FILLER_19_252 ();
 sg13g2_fill_1 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_324 ();
 sg13g2_decap_8 FILLER_19_331 ();
 sg13g2_decap_8 FILLER_19_338 ();
 sg13g2_decap_8 FILLER_19_345 ();
 sg13g2_decap_8 FILLER_19_352 ();
 sg13g2_decap_8 FILLER_19_359 ();
 sg13g2_decap_8 FILLER_19_366 ();
 sg13g2_decap_8 FILLER_19_373 ();
 sg13g2_decap_8 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_fill_2 FILLER_20_154 ();
 sg13g2_fill_2 FILLER_20_200 ();
 sg13g2_fill_2 FILLER_20_214 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_fill_2 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_262 ();
 sg13g2_fill_2 FILLER_20_269 ();
 sg13g2_decap_8 FILLER_20_327 ();
 sg13g2_decap_8 FILLER_20_334 ();
 sg13g2_decap_8 FILLER_20_341 ();
 sg13g2_decap_8 FILLER_20_348 ();
 sg13g2_decap_8 FILLER_20_355 ();
 sg13g2_decap_8 FILLER_20_362 ();
 sg13g2_decap_8 FILLER_20_369 ();
 sg13g2_decap_8 FILLER_20_376 ();
 sg13g2_decap_8 FILLER_20_383 ();
 sg13g2_decap_8 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_397 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_4 FILLER_21_168 ();
 sg13g2_fill_2 FILLER_21_172 ();
 sg13g2_fill_2 FILLER_21_177 ();
 sg13g2_fill_2 FILLER_21_200 ();
 sg13g2_fill_1 FILLER_21_202 ();
 sg13g2_fill_2 FILLER_21_220 ();
 sg13g2_fill_1 FILLER_21_222 ();
 sg13g2_fill_1 FILLER_21_228 ();
 sg13g2_decap_8 FILLER_21_265 ();
 sg13g2_decap_8 FILLER_21_272 ();
 sg13g2_fill_2 FILLER_21_279 ();
 sg13g2_decap_8 FILLER_21_316 ();
 sg13g2_decap_8 FILLER_21_323 ();
 sg13g2_decap_8 FILLER_21_330 ();
 sg13g2_decap_8 FILLER_21_337 ();
 sg13g2_decap_8 FILLER_21_344 ();
 sg13g2_decap_8 FILLER_21_351 ();
 sg13g2_decap_8 FILLER_21_358 ();
 sg13g2_decap_8 FILLER_21_365 ();
 sg13g2_decap_8 FILLER_21_372 ();
 sg13g2_decap_8 FILLER_21_379 ();
 sg13g2_decap_8 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_393 ();
 sg13g2_decap_8 FILLER_21_400 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_4 FILLER_22_182 ();
 sg13g2_fill_1 FILLER_22_186 ();
 sg13g2_fill_2 FILLER_22_195 ();
 sg13g2_decap_4 FILLER_22_202 ();
 sg13g2_fill_1 FILLER_22_219 ();
 sg13g2_decap_8 FILLER_22_244 ();
 sg13g2_fill_1 FILLER_22_251 ();
 sg13g2_decap_8 FILLER_22_257 ();
 sg13g2_decap_8 FILLER_22_264 ();
 sg13g2_fill_1 FILLER_22_271 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_fill_1 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_307 ();
 sg13g2_decap_8 FILLER_22_314 ();
 sg13g2_decap_8 FILLER_22_321 ();
 sg13g2_decap_8 FILLER_22_328 ();
 sg13g2_decap_8 FILLER_22_335 ();
 sg13g2_decap_8 FILLER_22_342 ();
 sg13g2_decap_8 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_decap_8 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_370 ();
 sg13g2_decap_8 FILLER_22_377 ();
 sg13g2_decap_8 FILLER_22_384 ();
 sg13g2_decap_8 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_fill_2 FILLER_23_194 ();
 sg13g2_fill_1 FILLER_23_196 ();
 sg13g2_fill_1 FILLER_23_212 ();
 sg13g2_fill_2 FILLER_23_223 ();
 sg13g2_decap_8 FILLER_23_241 ();
 sg13g2_fill_2 FILLER_23_248 ();
 sg13g2_fill_2 FILLER_23_292 ();
 sg13g2_decap_8 FILLER_23_317 ();
 sg13g2_decap_8 FILLER_23_324 ();
 sg13g2_decap_8 FILLER_23_331 ();
 sg13g2_decap_8 FILLER_23_338 ();
 sg13g2_decap_8 FILLER_23_345 ();
 sg13g2_decap_8 FILLER_23_352 ();
 sg13g2_decap_8 FILLER_23_359 ();
 sg13g2_decap_8 FILLER_23_366 ();
 sg13g2_decap_8 FILLER_23_373 ();
 sg13g2_decap_8 FILLER_23_380 ();
 sg13g2_decap_8 FILLER_23_387 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_fill_2 FILLER_24_189 ();
 sg13g2_fill_1 FILLER_24_221 ();
 sg13g2_fill_2 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_237 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_fill_2 FILLER_25_154 ();
 sg13g2_fill_1 FILLER_25_156 ();
 sg13g2_decap_8 FILLER_25_188 ();
 sg13g2_decap_8 FILLER_25_195 ();
 sg13g2_fill_2 FILLER_25_202 ();
 sg13g2_decap_8 FILLER_25_213 ();
 sg13g2_decap_4 FILLER_25_220 ();
 sg13g2_fill_1 FILLER_25_224 ();
 sg13g2_decap_4 FILLER_25_268 ();
 sg13g2_decap_8 FILLER_25_317 ();
 sg13g2_decap_8 FILLER_25_324 ();
 sg13g2_decap_8 FILLER_25_331 ();
 sg13g2_decap_8 FILLER_25_338 ();
 sg13g2_decap_8 FILLER_25_345 ();
 sg13g2_decap_8 FILLER_25_352 ();
 sg13g2_decap_8 FILLER_25_359 ();
 sg13g2_decap_8 FILLER_25_366 ();
 sg13g2_decap_8 FILLER_25_373 ();
 sg13g2_decap_8 FILLER_25_380 ();
 sg13g2_decap_8 FILLER_25_387 ();
 sg13g2_decap_8 FILLER_25_394 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_4 FILLER_26_154 ();
 sg13g2_decap_4 FILLER_26_168 ();
 sg13g2_fill_1 FILLER_26_172 ();
 sg13g2_decap_4 FILLER_26_194 ();
 sg13g2_fill_2 FILLER_26_198 ();
 sg13g2_fill_2 FILLER_26_205 ();
 sg13g2_fill_1 FILLER_26_233 ();
 sg13g2_fill_1 FILLER_26_244 ();
 sg13g2_decap_8 FILLER_26_255 ();
 sg13g2_fill_1 FILLER_26_262 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_fill_1 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_4 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_307 ();
 sg13g2_decap_8 FILLER_26_314 ();
 sg13g2_decap_8 FILLER_26_321 ();
 sg13g2_decap_8 FILLER_26_328 ();
 sg13g2_decap_8 FILLER_26_335 ();
 sg13g2_decap_8 FILLER_26_342 ();
 sg13g2_decap_8 FILLER_26_349 ();
 sg13g2_decap_8 FILLER_26_356 ();
 sg13g2_decap_8 FILLER_26_363 ();
 sg13g2_decap_8 FILLER_26_370 ();
 sg13g2_decap_8 FILLER_26_377 ();
 sg13g2_decap_8 FILLER_26_384 ();
 sg13g2_decap_8 FILLER_26_391 ();
 sg13g2_decap_8 FILLER_26_398 ();
 sg13g2_decap_4 FILLER_26_405 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_4 FILLER_27_175 ();
 sg13g2_fill_1 FILLER_27_179 ();
 sg13g2_decap_8 FILLER_27_200 ();
 sg13g2_decap_8 FILLER_27_207 ();
 sg13g2_decap_8 FILLER_27_214 ();
 sg13g2_decap_8 FILLER_27_221 ();
 sg13g2_decap_8 FILLER_27_228 ();
 sg13g2_decap_4 FILLER_27_235 ();
 sg13g2_fill_1 FILLER_27_239 ();
 sg13g2_fill_2 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_257 ();
 sg13g2_decap_8 FILLER_27_264 ();
 sg13g2_decap_8 FILLER_27_271 ();
 sg13g2_fill_1 FILLER_27_278 ();
 sg13g2_decap_8 FILLER_27_305 ();
 sg13g2_decap_8 FILLER_27_312 ();
 sg13g2_decap_8 FILLER_27_319 ();
 sg13g2_decap_8 FILLER_27_326 ();
 sg13g2_decap_8 FILLER_27_333 ();
 sg13g2_decap_8 FILLER_27_340 ();
 sg13g2_decap_8 FILLER_27_347 ();
 sg13g2_decap_8 FILLER_27_354 ();
 sg13g2_decap_8 FILLER_27_361 ();
 sg13g2_decap_8 FILLER_27_368 ();
 sg13g2_decap_8 FILLER_27_375 ();
 sg13g2_decap_8 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_27_396 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_fill_2 FILLER_28_147 ();
 sg13g2_fill_2 FILLER_28_180 ();
 sg13g2_fill_1 FILLER_28_182 ();
 sg13g2_fill_2 FILLER_28_232 ();
 sg13g2_fill_1 FILLER_28_234 ();
 sg13g2_fill_1 FILLER_28_245 ();
 sg13g2_decap_4 FILLER_28_266 ();
 sg13g2_fill_2 FILLER_28_284 ();
 sg13g2_fill_1 FILLER_28_299 ();
 sg13g2_decap_8 FILLER_28_320 ();
 sg13g2_decap_8 FILLER_28_327 ();
 sg13g2_decap_8 FILLER_28_334 ();
 sg13g2_decap_8 FILLER_28_341 ();
 sg13g2_decap_8 FILLER_28_348 ();
 sg13g2_decap_8 FILLER_28_355 ();
 sg13g2_decap_8 FILLER_28_362 ();
 sg13g2_decap_8 FILLER_28_369 ();
 sg13g2_decap_8 FILLER_28_376 ();
 sg13g2_decap_8 FILLER_28_383 ();
 sg13g2_decap_8 FILLER_28_390 ();
 sg13g2_decap_8 FILLER_28_397 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_4 FILLER_29_133 ();
 sg13g2_fill_1 FILLER_29_137 ();
 sg13g2_decap_4 FILLER_29_202 ();
 sg13g2_fill_2 FILLER_29_206 ();
 sg13g2_decap_8 FILLER_29_216 ();
 sg13g2_fill_2 FILLER_29_223 ();
 sg13g2_fill_1 FILLER_29_239 ();
 sg13g2_fill_1 FILLER_29_246 ();
 sg13g2_fill_1 FILLER_29_300 ();
 sg13g2_decap_8 FILLER_29_327 ();
 sg13g2_decap_8 FILLER_29_334 ();
 sg13g2_decap_8 FILLER_29_341 ();
 sg13g2_decap_8 FILLER_29_348 ();
 sg13g2_decap_8 FILLER_29_355 ();
 sg13g2_decap_8 FILLER_29_362 ();
 sg13g2_decap_8 FILLER_29_369 ();
 sg13g2_decap_8 FILLER_29_376 ();
 sg13g2_decap_8 FILLER_29_383 ();
 sg13g2_decap_8 FILLER_29_390 ();
 sg13g2_decap_8 FILLER_29_397 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_fill_2 FILLER_30_133 ();
 sg13g2_fill_1 FILLER_30_135 ();
 sg13g2_fill_1 FILLER_30_158 ();
 sg13g2_fill_1 FILLER_30_169 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_fill_2 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_213 ();
 sg13g2_fill_1 FILLER_30_220 ();
 sg13g2_decap_4 FILLER_30_242 ();
 sg13g2_decap_8 FILLER_30_261 ();
 sg13g2_decap_8 FILLER_30_268 ();
 sg13g2_fill_2 FILLER_30_296 ();
 sg13g2_decap_8 FILLER_30_321 ();
 sg13g2_decap_8 FILLER_30_328 ();
 sg13g2_decap_8 FILLER_30_335 ();
 sg13g2_decap_8 FILLER_30_342 ();
 sg13g2_decap_8 FILLER_30_349 ();
 sg13g2_decap_8 FILLER_30_356 ();
 sg13g2_decap_8 FILLER_30_363 ();
 sg13g2_decap_8 FILLER_30_370 ();
 sg13g2_decap_8 FILLER_30_377 ();
 sg13g2_decap_8 FILLER_30_384 ();
 sg13g2_decap_8 FILLER_30_391 ();
 sg13g2_decap_8 FILLER_30_398 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_fill_2 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_186 ();
 sg13g2_fill_2 FILLER_31_193 ();
 sg13g2_decap_8 FILLER_31_204 ();
 sg13g2_decap_8 FILLER_31_211 ();
 sg13g2_fill_2 FILLER_31_218 ();
 sg13g2_fill_1 FILLER_31_229 ();
 sg13g2_fill_2 FILLER_31_235 ();
 sg13g2_fill_1 FILLER_31_237 ();
 sg13g2_decap_8 FILLER_31_254 ();
 sg13g2_decap_8 FILLER_31_261 ();
 sg13g2_decap_4 FILLER_31_268 ();
 sg13g2_fill_2 FILLER_31_285 ();
 sg13g2_fill_1 FILLER_31_287 ();
 sg13g2_decap_4 FILLER_31_296 ();
 sg13g2_fill_2 FILLER_31_304 ();
 sg13g2_decap_8 FILLER_31_310 ();
 sg13g2_decap_8 FILLER_31_317 ();
 sg13g2_decap_8 FILLER_31_324 ();
 sg13g2_decap_8 FILLER_31_331 ();
 sg13g2_decap_8 FILLER_31_338 ();
 sg13g2_decap_8 FILLER_31_345 ();
 sg13g2_decap_8 FILLER_31_352 ();
 sg13g2_decap_8 FILLER_31_359 ();
 sg13g2_decap_8 FILLER_31_366 ();
 sg13g2_decap_8 FILLER_31_373 ();
 sg13g2_decap_8 FILLER_31_380 ();
 sg13g2_decap_8 FILLER_31_387 ();
 sg13g2_decap_8 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_4 FILLER_32_161 ();
 sg13g2_fill_2 FILLER_32_174 ();
 sg13g2_decap_4 FILLER_32_186 ();
 sg13g2_fill_1 FILLER_32_190 ();
 sg13g2_fill_1 FILLER_32_202 ();
 sg13g2_fill_2 FILLER_32_211 ();
 sg13g2_decap_8 FILLER_32_243 ();
 sg13g2_decap_8 FILLER_32_263 ();
 sg13g2_decap_8 FILLER_32_270 ();
 sg13g2_fill_2 FILLER_32_301 ();
 sg13g2_decap_8 FILLER_32_315 ();
 sg13g2_decap_8 FILLER_32_322 ();
 sg13g2_decap_8 FILLER_32_329 ();
 sg13g2_decap_8 FILLER_32_336 ();
 sg13g2_decap_8 FILLER_32_343 ();
 sg13g2_decap_8 FILLER_32_350 ();
 sg13g2_decap_8 FILLER_32_357 ();
 sg13g2_decap_8 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_decap_8 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_fill_2 FILLER_33_140 ();
 sg13g2_fill_1 FILLER_33_163 ();
 sg13g2_fill_2 FILLER_33_169 ();
 sg13g2_fill_1 FILLER_33_171 ();
 sg13g2_fill_2 FILLER_33_187 ();
 sg13g2_decap_8 FILLER_33_223 ();
 sg13g2_decap_4 FILLER_33_230 ();
 sg13g2_decap_4 FILLER_33_239 ();
 sg13g2_fill_2 FILLER_33_248 ();
 sg13g2_fill_1 FILLER_33_271 ();
 sg13g2_fill_1 FILLER_33_299 ();
 sg13g2_decap_8 FILLER_33_319 ();
 sg13g2_decap_8 FILLER_33_326 ();
 sg13g2_decap_8 FILLER_33_333 ();
 sg13g2_decap_8 FILLER_33_340 ();
 sg13g2_decap_8 FILLER_33_347 ();
 sg13g2_decap_8 FILLER_33_354 ();
 sg13g2_decap_8 FILLER_33_361 ();
 sg13g2_decap_8 FILLER_33_368 ();
 sg13g2_decap_8 FILLER_33_375 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_33_389 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_4 FILLER_34_140 ();
 sg13g2_fill_2 FILLER_34_144 ();
 sg13g2_fill_1 FILLER_34_164 ();
 sg13g2_fill_2 FILLER_34_172 ();
 sg13g2_decap_8 FILLER_34_183 ();
 sg13g2_fill_2 FILLER_34_190 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_fill_2 FILLER_34_231 ();
 sg13g2_fill_2 FILLER_34_269 ();
 sg13g2_fill_2 FILLER_34_291 ();
 sg13g2_fill_2 FILLER_34_298 ();
 sg13g2_fill_1 FILLER_34_300 ();
 sg13g2_decap_8 FILLER_34_311 ();
 sg13g2_decap_8 FILLER_34_318 ();
 sg13g2_decap_8 FILLER_34_325 ();
 sg13g2_decap_8 FILLER_34_332 ();
 sg13g2_decap_8 FILLER_34_339 ();
 sg13g2_decap_8 FILLER_34_346 ();
 sg13g2_decap_8 FILLER_34_353 ();
 sg13g2_decap_8 FILLER_34_360 ();
 sg13g2_decap_8 FILLER_34_367 ();
 sg13g2_decap_8 FILLER_34_374 ();
 sg13g2_decap_8 FILLER_34_381 ();
 sg13g2_decap_8 FILLER_34_388 ();
 sg13g2_decap_8 FILLER_34_395 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_4 FILLER_35_133 ();
 sg13g2_fill_2 FILLER_35_137 ();
 sg13g2_fill_2 FILLER_35_163 ();
 sg13g2_fill_1 FILLER_35_165 ();
 sg13g2_fill_2 FILLER_35_176 ();
 sg13g2_decap_8 FILLER_35_190 ();
 sg13g2_fill_2 FILLER_35_197 ();
 sg13g2_fill_1 FILLER_35_199 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_fill_2 FILLER_35_217 ();
 sg13g2_decap_4 FILLER_35_237 ();
 sg13g2_fill_2 FILLER_35_241 ();
 sg13g2_fill_2 FILLER_35_295 ();
 sg13g2_fill_1 FILLER_35_297 ();
 sg13g2_decap_8 FILLER_35_309 ();
 sg13g2_decap_8 FILLER_35_316 ();
 sg13g2_decap_4 FILLER_35_323 ();
 sg13g2_fill_1 FILLER_35_327 ();
 sg13g2_decap_4 FILLER_35_333 ();
 sg13g2_decap_8 FILLER_35_353 ();
 sg13g2_decap_8 FILLER_35_360 ();
 sg13g2_decap_8 FILLER_35_367 ();
 sg13g2_decap_8 FILLER_35_374 ();
 sg13g2_decap_8 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_35_388 ();
 sg13g2_decap_8 FILLER_35_395 ();
 sg13g2_decap_8 FILLER_35_402 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_4 FILLER_36_126 ();
 sg13g2_fill_2 FILLER_36_164 ();
 sg13g2_fill_1 FILLER_36_166 ();
 sg13g2_fill_2 FILLER_36_175 ();
 sg13g2_fill_1 FILLER_36_177 ();
 sg13g2_fill_2 FILLER_36_184 ();
 sg13g2_decap_4 FILLER_36_189 ();
 sg13g2_fill_1 FILLER_36_193 ();
 sg13g2_fill_2 FILLER_36_208 ();
 sg13g2_fill_1 FILLER_36_241 ();
 sg13g2_fill_2 FILLER_36_246 ();
 sg13g2_fill_2 FILLER_36_253 ();
 sg13g2_fill_1 FILLER_36_255 ();
 sg13g2_decap_8 FILLER_36_265 ();
 sg13g2_decap_8 FILLER_36_272 ();
 sg13g2_decap_8 FILLER_36_279 ();
 sg13g2_decap_8 FILLER_36_286 ();
 sg13g2_decap_8 FILLER_36_293 ();
 sg13g2_decap_4 FILLER_36_300 ();
 sg13g2_decap_8 FILLER_36_362 ();
 sg13g2_decap_8 FILLER_36_369 ();
 sg13g2_decap_8 FILLER_36_376 ();
 sg13g2_decap_8 FILLER_36_383 ();
 sg13g2_decap_8 FILLER_36_390 ();
 sg13g2_decap_8 FILLER_36_397 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_4 FILLER_37_133 ();
 sg13g2_fill_1 FILLER_37_137 ();
 sg13g2_decap_4 FILLER_37_146 ();
 sg13g2_fill_2 FILLER_37_150 ();
 sg13g2_fill_2 FILLER_37_171 ();
 sg13g2_fill_2 FILLER_37_179 ();
 sg13g2_fill_2 FILLER_37_219 ();
 sg13g2_fill_1 FILLER_37_227 ();
 sg13g2_fill_2 FILLER_37_238 ();
 sg13g2_decap_4 FILLER_37_263 ();
 sg13g2_fill_2 FILLER_37_267 ();
 sg13g2_decap_4 FILLER_37_316 ();
 sg13g2_fill_1 FILLER_37_320 ();
 sg13g2_decap_8 FILLER_37_354 ();
 sg13g2_decap_8 FILLER_37_361 ();
 sg13g2_decap_8 FILLER_37_368 ();
 sg13g2_decap_8 FILLER_37_375 ();
 sg13g2_decap_8 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_396 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_fill_2 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_122 ();
 sg13g2_decap_8 FILLER_38_129 ();
 sg13g2_decap_8 FILLER_38_136 ();
 sg13g2_decap_8 FILLER_38_143 ();
 sg13g2_decap_4 FILLER_38_150 ();
 sg13g2_decap_4 FILLER_38_169 ();
 sg13g2_fill_1 FILLER_38_183 ();
 sg13g2_decap_8 FILLER_38_207 ();
 sg13g2_decap_4 FILLER_38_214 ();
 sg13g2_fill_2 FILLER_38_218 ();
 sg13g2_fill_2 FILLER_38_248 ();
 sg13g2_fill_1 FILLER_38_265 ();
 sg13g2_decap_4 FILLER_38_304 ();
 sg13g2_decap_8 FILLER_38_321 ();
 sg13g2_fill_1 FILLER_38_328 ();
 sg13g2_fill_1 FILLER_38_342 ();
 sg13g2_fill_2 FILLER_38_358 ();
 sg13g2_fill_1 FILLER_38_360 ();
 sg13g2_decap_8 FILLER_38_376 ();
 sg13g2_decap_8 FILLER_38_383 ();
 sg13g2_decap_8 FILLER_38_390 ();
 sg13g2_decap_8 FILLER_38_397 ();
 sg13g2_decap_4 FILLER_38_404 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_fill_2 FILLER_39_105 ();
 sg13g2_fill_2 FILLER_39_142 ();
 sg13g2_fill_2 FILLER_39_178 ();
 sg13g2_fill_1 FILLER_39_180 ();
 sg13g2_decap_4 FILLER_39_194 ();
 sg13g2_decap_8 FILLER_39_210 ();
 sg13g2_fill_2 FILLER_39_217 ();
 sg13g2_fill_1 FILLER_39_219 ();
 sg13g2_fill_2 FILLER_39_249 ();
 sg13g2_fill_1 FILLER_39_251 ();
 sg13g2_fill_2 FILLER_39_275 ();
 sg13g2_decap_8 FILLER_39_289 ();
 sg13g2_fill_2 FILLER_39_296 ();
 sg13g2_fill_1 FILLER_39_339 ();
 sg13g2_fill_2 FILLER_39_358 ();
 sg13g2_fill_1 FILLER_39_360 ();
 sg13g2_decap_8 FILLER_39_387 ();
 sg13g2_decap_8 FILLER_39_394 ();
 sg13g2_decap_8 FILLER_39_401 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_4 FILLER_40_84 ();
 sg13g2_fill_1 FILLER_40_123 ();
 sg13g2_decap_4 FILLER_40_150 ();
 sg13g2_fill_1 FILLER_40_163 ();
 sg13g2_fill_2 FILLER_40_168 ();
 sg13g2_fill_1 FILLER_40_170 ();
 sg13g2_fill_2 FILLER_40_183 ();
 sg13g2_fill_2 FILLER_40_200 ();
 sg13g2_decap_4 FILLER_40_224 ();
 sg13g2_fill_2 FILLER_40_245 ();
 sg13g2_decap_4 FILLER_40_278 ();
 sg13g2_fill_1 FILLER_40_282 ();
 sg13g2_decap_8 FILLER_40_291 ();
 sg13g2_fill_2 FILLER_40_298 ();
 sg13g2_fill_2 FILLER_40_305 ();
 sg13g2_decap_8 FILLER_40_312 ();
 sg13g2_fill_2 FILLER_40_319 ();
 sg13g2_fill_1 FILLER_40_321 ();
 sg13g2_decap_4 FILLER_40_327 ();
 sg13g2_fill_2 FILLER_40_349 ();
 sg13g2_fill_1 FILLER_40_351 ();
 sg13g2_fill_1 FILLER_40_362 ();
 sg13g2_decap_8 FILLER_40_376 ();
 sg13g2_decap_8 FILLER_40_383 ();
 sg13g2_decap_8 FILLER_40_390 ();
 sg13g2_decap_8 FILLER_40_397 ();
 sg13g2_decap_4 FILLER_40_404 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_4 FILLER_41_77 ();
 sg13g2_fill_2 FILLER_41_81 ();
 sg13g2_decap_8 FILLER_41_163 ();
 sg13g2_fill_2 FILLER_41_170 ();
 sg13g2_fill_2 FILLER_41_191 ();
 sg13g2_fill_1 FILLER_41_193 ();
 sg13g2_fill_2 FILLER_41_199 ();
 sg13g2_fill_2 FILLER_41_210 ();
 sg13g2_decap_8 FILLER_41_232 ();
 sg13g2_decap_8 FILLER_41_244 ();
 sg13g2_decap_4 FILLER_41_251 ();
 sg13g2_fill_1 FILLER_41_255 ();
 sg13g2_decap_4 FILLER_41_285 ();
 sg13g2_fill_2 FILLER_41_295 ();
 sg13g2_fill_1 FILLER_41_301 ();
 sg13g2_fill_2 FILLER_41_307 ();
 sg13g2_decap_8 FILLER_41_317 ();
 sg13g2_decap_4 FILLER_41_324 ();
 sg13g2_fill_2 FILLER_41_328 ();
 sg13g2_decap_8 FILLER_41_391 ();
 sg13g2_decap_8 FILLER_41_398 ();
 sg13g2_decap_4 FILLER_41_405 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_fill_2 FILLER_42_102 ();
 sg13g2_fill_1 FILLER_42_122 ();
 sg13g2_decap_4 FILLER_42_163 ();
 sg13g2_fill_2 FILLER_42_177 ();
 sg13g2_decap_4 FILLER_42_184 ();
 sg13g2_decap_8 FILLER_42_203 ();
 sg13g2_decap_8 FILLER_42_210 ();
 sg13g2_decap_8 FILLER_42_217 ();
 sg13g2_decap_8 FILLER_42_224 ();
 sg13g2_decap_8 FILLER_42_231 ();
 sg13g2_decap_8 FILLER_42_238 ();
 sg13g2_decap_8 FILLER_42_245 ();
 sg13g2_decap_8 FILLER_42_256 ();
 sg13g2_decap_4 FILLER_42_263 ();
 sg13g2_decap_8 FILLER_42_312 ();
 sg13g2_fill_2 FILLER_42_319 ();
 sg13g2_fill_1 FILLER_42_321 ();
 sg13g2_decap_8 FILLER_42_327 ();
 sg13g2_decap_4 FILLER_42_334 ();
 sg13g2_fill_1 FILLER_42_338 ();
 sg13g2_decap_8 FILLER_42_344 ();
 sg13g2_fill_2 FILLER_42_351 ();
 sg13g2_fill_1 FILLER_42_353 ();
 sg13g2_fill_2 FILLER_42_360 ();
 sg13g2_decap_8 FILLER_42_373 ();
 sg13g2_decap_8 FILLER_42_380 ();
 sg13g2_decap_8 FILLER_42_387 ();
 sg13g2_decap_8 FILLER_42_394 ();
 sg13g2_decap_8 FILLER_42_401 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_fill_2 FILLER_43_77 ();
 sg13g2_fill_2 FILLER_43_112 ();
 sg13g2_fill_2 FILLER_43_155 ();
 sg13g2_fill_2 FILLER_43_170 ();
 sg13g2_fill_1 FILLER_43_180 ();
 sg13g2_fill_2 FILLER_43_192 ();
 sg13g2_decap_8 FILLER_43_199 ();
 sg13g2_decap_8 FILLER_43_206 ();
 sg13g2_decap_8 FILLER_43_213 ();
 sg13g2_decap_4 FILLER_43_220 ();
 sg13g2_decap_8 FILLER_43_250 ();
 sg13g2_decap_4 FILLER_43_257 ();
 sg13g2_fill_1 FILLER_43_261 ();
 sg13g2_fill_2 FILLER_43_267 ();
 sg13g2_fill_1 FILLER_43_269 ();
 sg13g2_decap_4 FILLER_43_296 ();
 sg13g2_fill_2 FILLER_43_300 ();
 sg13g2_fill_2 FILLER_43_328 ();
 sg13g2_fill_2 FILLER_43_348 ();
 sg13g2_fill_1 FILLER_43_350 ();
 sg13g2_decap_8 FILLER_43_380 ();
 sg13g2_decap_8 FILLER_43_387 ();
 sg13g2_decap_8 FILLER_43_394 ();
 sg13g2_decap_8 FILLER_43_401 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_fill_2 FILLER_44_84 ();
 sg13g2_fill_1 FILLER_44_112 ();
 sg13g2_fill_2 FILLER_44_139 ();
 sg13g2_fill_1 FILLER_44_141 ();
 sg13g2_fill_1 FILLER_44_184 ();
 sg13g2_fill_2 FILLER_44_190 ();
 sg13g2_decap_4 FILLER_44_227 ();
 sg13g2_fill_2 FILLER_44_231 ();
 sg13g2_decap_4 FILLER_44_249 ();
 sg13g2_fill_2 FILLER_44_253 ();
 sg13g2_decap_8 FILLER_44_276 ();
 sg13g2_decap_8 FILLER_44_283 ();
 sg13g2_decap_8 FILLER_44_290 ();
 sg13g2_fill_1 FILLER_44_297 ();
 sg13g2_decap_4 FILLER_44_324 ();
 sg13g2_fill_2 FILLER_44_349 ();
 sg13g2_fill_1 FILLER_44_351 ();
 sg13g2_decap_4 FILLER_44_369 ();
 sg13g2_decap_8 FILLER_44_394 ();
 sg13g2_decap_8 FILLER_44_401 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_fill_2 FILLER_45_91 ();
 sg13g2_fill_1 FILLER_45_117 ();
 sg13g2_fill_2 FILLER_45_179 ();
 sg13g2_fill_1 FILLER_45_181 ();
 sg13g2_decap_8 FILLER_45_232 ();
 sg13g2_decap_4 FILLER_45_239 ();
 sg13g2_decap_8 FILLER_45_267 ();
 sg13g2_fill_1 FILLER_45_274 ();
 sg13g2_decap_4 FILLER_45_278 ();
 sg13g2_fill_2 FILLER_45_282 ();
 sg13g2_decap_8 FILLER_45_288 ();
 sg13g2_decap_8 FILLER_45_295 ();
 sg13g2_decap_4 FILLER_45_302 ();
 sg13g2_fill_2 FILLER_45_306 ();
 sg13g2_fill_1 FILLER_45_333 ();
 sg13g2_fill_1 FILLER_45_350 ();
 sg13g2_decap_8 FILLER_45_385 ();
 sg13g2_decap_8 FILLER_45_392 ();
 sg13g2_decap_8 FILLER_45_399 ();
 sg13g2_fill_2 FILLER_45_406 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_fill_2 FILLER_46_84 ();
 sg13g2_fill_1 FILLER_46_112 ();
 sg13g2_fill_1 FILLER_46_118 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_decap_4 FILLER_46_168 ();
 sg13g2_fill_1 FILLER_46_172 ();
 sg13g2_decap_8 FILLER_46_188 ();
 sg13g2_decap_8 FILLER_46_195 ();
 sg13g2_fill_2 FILLER_46_202 ();
 sg13g2_decap_8 FILLER_46_236 ();
 sg13g2_decap_4 FILLER_46_243 ();
 sg13g2_decap_8 FILLER_46_260 ();
 sg13g2_decap_8 FILLER_46_289 ();
 sg13g2_decap_8 FILLER_46_296 ();
 sg13g2_decap_8 FILLER_46_303 ();
 sg13g2_decap_8 FILLER_46_310 ();
 sg13g2_decap_8 FILLER_46_317 ();
 sg13g2_decap_8 FILLER_46_338 ();
 sg13g2_decap_4 FILLER_46_345 ();
 sg13g2_decap_4 FILLER_46_354 ();
 sg13g2_decap_4 FILLER_46_371 ();
 sg13g2_fill_1 FILLER_46_375 ();
 sg13g2_decap_8 FILLER_46_388 ();
 sg13g2_decap_8 FILLER_46_395 ();
 sg13g2_decap_8 FILLER_46_402 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_4 FILLER_47_84 ();
 sg13g2_fill_1 FILLER_47_88 ();
 sg13g2_fill_1 FILLER_47_149 ();
 sg13g2_decap_8 FILLER_47_155 ();
 sg13g2_fill_2 FILLER_47_162 ();
 sg13g2_decap_8 FILLER_47_167 ();
 sg13g2_decap_8 FILLER_47_174 ();
 sg13g2_decap_8 FILLER_47_181 ();
 sg13g2_fill_1 FILLER_47_188 ();
 sg13g2_decap_8 FILLER_47_198 ();
 sg13g2_fill_2 FILLER_47_245 ();
 sg13g2_fill_2 FILLER_47_253 ();
 sg13g2_fill_1 FILLER_47_255 ();
 sg13g2_fill_2 FILLER_47_262 ();
 sg13g2_fill_1 FILLER_47_273 ();
 sg13g2_decap_8 FILLER_47_316 ();
 sg13g2_decap_4 FILLER_47_323 ();
 sg13g2_decap_8 FILLER_47_331 ();
 sg13g2_decap_4 FILLER_47_338 ();
 sg13g2_decap_4 FILLER_47_347 ();
 sg13g2_decap_8 FILLER_47_391 ();
 sg13g2_decap_8 FILLER_47_398 ();
 sg13g2_decap_4 FILLER_47_405 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_4 FILLER_48_91 ();
 sg13g2_decap_4 FILLER_48_142 ();
 sg13g2_decap_4 FILLER_48_207 ();
 sg13g2_fill_1 FILLER_48_211 ();
 sg13g2_fill_2 FILLER_48_220 ();
 sg13g2_fill_1 FILLER_48_222 ();
 sg13g2_fill_1 FILLER_48_260 ();
 sg13g2_fill_1 FILLER_48_274 ();
 sg13g2_fill_1 FILLER_48_366 ();
 sg13g2_decap_8 FILLER_48_393 ();
 sg13g2_decap_8 FILLER_48_400 ();
 sg13g2_fill_2 FILLER_48_407 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_fill_2 FILLER_49_91 ();
 sg13g2_fill_1 FILLER_49_93 ();
 sg13g2_fill_2 FILLER_49_172 ();
 sg13g2_fill_1 FILLER_49_214 ();
 sg13g2_fill_2 FILLER_49_249 ();
 sg13g2_fill_1 FILLER_49_260 ();
 sg13g2_fill_1 FILLER_49_276 ();
 sg13g2_fill_2 FILLER_49_315 ();
 sg13g2_fill_1 FILLER_49_317 ();
 sg13g2_fill_1 FILLER_49_354 ();
 sg13g2_decap_8 FILLER_49_385 ();
 sg13g2_decap_8 FILLER_49_392 ();
 sg13g2_decap_8 FILLER_49_399 ();
 sg13g2_fill_2 FILLER_49_406 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_fill_2 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_177 ();
 sg13g2_fill_1 FILLER_50_184 ();
 sg13g2_decap_8 FILLER_50_217 ();
 sg13g2_fill_2 FILLER_50_224 ();
 sg13g2_fill_1 FILLER_50_226 ();
 sg13g2_decap_4 FILLER_50_233 ();
 sg13g2_fill_2 FILLER_50_254 ();
 sg13g2_decap_8 FILLER_50_286 ();
 sg13g2_decap_8 FILLER_50_293 ();
 sg13g2_decap_4 FILLER_50_305 ();
 sg13g2_fill_1 FILLER_50_309 ();
 sg13g2_decap_8 FILLER_50_342 ();
 sg13g2_decap_8 FILLER_50_369 ();
 sg13g2_decap_8 FILLER_50_376 ();
 sg13g2_decap_8 FILLER_50_383 ();
 sg13g2_decap_8 FILLER_50_390 ();
 sg13g2_decap_8 FILLER_50_397 ();
 sg13g2_decap_4 FILLER_50_404 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_4 FILLER_51_98 ();
 sg13g2_decap_4 FILLER_51_145 ();
 sg13g2_decap_8 FILLER_51_170 ();
 sg13g2_decap_8 FILLER_51_177 ();
 sg13g2_fill_2 FILLER_51_184 ();
 sg13g2_fill_2 FILLER_51_228 ();
 sg13g2_fill_1 FILLER_51_230 ();
 sg13g2_decap_8 FILLER_51_244 ();
 sg13g2_decap_8 FILLER_51_251 ();
 sg13g2_decap_4 FILLER_51_258 ();
 sg13g2_fill_1 FILLER_51_262 ();
 sg13g2_decap_8 FILLER_51_269 ();
 sg13g2_decap_8 FILLER_51_276 ();
 sg13g2_decap_4 FILLER_51_290 ();
 sg13g2_fill_1 FILLER_51_294 ();
 sg13g2_fill_1 FILLER_51_315 ();
 sg13g2_decap_8 FILLER_51_333 ();
 sg13g2_decap_8 FILLER_51_340 ();
 sg13g2_decap_8 FILLER_51_347 ();
 sg13g2_decap_8 FILLER_51_354 ();
 sg13g2_decap_8 FILLER_51_361 ();
 sg13g2_decap_8 FILLER_51_368 ();
 sg13g2_decap_8 FILLER_51_375 ();
 sg13g2_decap_8 FILLER_51_382 ();
 sg13g2_decap_8 FILLER_51_389 ();
 sg13g2_decap_8 FILLER_51_396 ();
 sg13g2_decap_4 FILLER_51_403 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_fill_2 FILLER_52_105 ();
 sg13g2_fill_1 FILLER_52_107 ();
 sg13g2_fill_2 FILLER_52_122 ();
 sg13g2_decap_4 FILLER_52_138 ();
 sg13g2_fill_2 FILLER_52_142 ();
 sg13g2_fill_2 FILLER_52_180 ();
 sg13g2_fill_1 FILLER_52_182 ();
 sg13g2_decap_8 FILLER_52_191 ();
 sg13g2_fill_2 FILLER_52_198 ();
 sg13g2_fill_1 FILLER_52_200 ();
 sg13g2_decap_4 FILLER_52_261 ();
 sg13g2_decap_8 FILLER_52_274 ();
 sg13g2_fill_1 FILLER_52_281 ();
 sg13g2_decap_8 FILLER_52_354 ();
 sg13g2_decap_8 FILLER_52_361 ();
 sg13g2_fill_2 FILLER_52_368 ();
 sg13g2_fill_1 FILLER_52_370 ();
 sg13g2_decap_8 FILLER_52_397 ();
 sg13g2_decap_4 FILLER_52_404 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_fill_2 FILLER_53_105 ();
 sg13g2_fill_1 FILLER_53_107 ();
 sg13g2_decap_8 FILLER_53_134 ();
 sg13g2_decap_8 FILLER_53_141 ();
 sg13g2_decap_8 FILLER_53_148 ();
 sg13g2_decap_8 FILLER_53_155 ();
 sg13g2_decap_8 FILLER_53_162 ();
 sg13g2_fill_2 FILLER_53_169 ();
 sg13g2_decap_8 FILLER_53_206 ();
 sg13g2_decap_4 FILLER_53_213 ();
 sg13g2_decap_4 FILLER_53_222 ();
 sg13g2_fill_1 FILLER_53_226 ();
 sg13g2_decap_8 FILLER_53_237 ();
 sg13g2_decap_8 FILLER_53_244 ();
 sg13g2_decap_4 FILLER_53_251 ();
 sg13g2_fill_1 FILLER_53_259 ();
 sg13g2_fill_1 FILLER_53_265 ();
 sg13g2_fill_2 FILLER_53_326 ();
 sg13g2_fill_1 FILLER_53_354 ();
 sg13g2_decap_8 FILLER_53_391 ();
 sg13g2_decap_8 FILLER_53_398 ();
 sg13g2_decap_4 FILLER_53_405 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_4 FILLER_54_105 ();
 sg13g2_fill_2 FILLER_54_109 ();
 sg13g2_decap_4 FILLER_54_163 ();
 sg13g2_fill_2 FILLER_54_167 ();
 sg13g2_fill_1 FILLER_54_172 ();
 sg13g2_fill_2 FILLER_54_176 ();
 sg13g2_decap_8 FILLER_54_210 ();
 sg13g2_decap_8 FILLER_54_217 ();
 sg13g2_decap_8 FILLER_54_224 ();
 sg13g2_fill_2 FILLER_54_231 ();
 sg13g2_fill_2 FILLER_54_283 ();
 sg13g2_fill_1 FILLER_54_285 ();
 sg13g2_decap_8 FILLER_54_301 ();
 sg13g2_decap_8 FILLER_54_308 ();
 sg13g2_fill_1 FILLER_54_315 ();
 sg13g2_fill_1 FILLER_54_366 ();
 sg13g2_decap_8 FILLER_54_377 ();
 sg13g2_decap_8 FILLER_54_384 ();
 sg13g2_decap_8 FILLER_54_391 ();
 sg13g2_decap_8 FILLER_54_398 ();
 sg13g2_decap_4 FILLER_54_405 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_fill_2 FILLER_55_98 ();
 sg13g2_fill_1 FILLER_55_100 ();
 sg13g2_decap_8 FILLER_55_121 ();
 sg13g2_fill_1 FILLER_55_180 ();
 sg13g2_fill_1 FILLER_55_213 ();
 sg13g2_decap_4 FILLER_55_222 ();
 sg13g2_fill_2 FILLER_55_226 ();
 sg13g2_fill_2 FILLER_55_240 ();
 sg13g2_decap_4 FILLER_55_287 ();
 sg13g2_decap_8 FILLER_55_301 ();
 sg13g2_fill_1 FILLER_55_308 ();
 sg13g2_fill_2 FILLER_55_313 ();
 sg13g2_fill_1 FILLER_55_322 ();
 sg13g2_decap_8 FILLER_55_328 ();
 sg13g2_decap_8 FILLER_55_335 ();
 sg13g2_decap_8 FILLER_55_342 ();
 sg13g2_decap_8 FILLER_55_349 ();
 sg13g2_decap_8 FILLER_55_371 ();
 sg13g2_decap_8 FILLER_55_378 ();
 sg13g2_decap_8 FILLER_55_385 ();
 sg13g2_decap_8 FILLER_55_392 ();
 sg13g2_decap_8 FILLER_55_399 ();
 sg13g2_fill_2 FILLER_55_406 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_4 FILLER_56_98 ();
 sg13g2_decap_4 FILLER_56_137 ();
 sg13g2_decap_4 FILLER_56_151 ();
 sg13g2_fill_2 FILLER_56_171 ();
 sg13g2_decap_4 FILLER_56_258 ();
 sg13g2_decap_8 FILLER_56_272 ();
 sg13g2_fill_2 FILLER_56_279 ();
 sg13g2_fill_1 FILLER_56_281 ();
 sg13g2_decap_8 FILLER_56_286 ();
 sg13g2_decap_8 FILLER_56_293 ();
 sg13g2_fill_1 FILLER_56_300 ();
 sg13g2_fill_2 FILLER_56_307 ();
 sg13g2_fill_2 FILLER_56_314 ();
 sg13g2_fill_2 FILLER_56_325 ();
 sg13g2_fill_1 FILLER_56_327 ();
 sg13g2_decap_8 FILLER_56_337 ();
 sg13g2_decap_4 FILLER_56_344 ();
 sg13g2_fill_2 FILLER_56_348 ();
 sg13g2_decap_8 FILLER_56_389 ();
 sg13g2_decap_8 FILLER_56_396 ();
 sg13g2_decap_4 FILLER_56_403 ();
 sg13g2_fill_2 FILLER_56_407 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_4 FILLER_57_91 ();
 sg13g2_fill_1 FILLER_57_95 ();
 sg13g2_fill_2 FILLER_57_128 ();
 sg13g2_fill_1 FILLER_57_130 ();
 sg13g2_fill_1 FILLER_57_134 ();
 sg13g2_fill_1 FILLER_57_144 ();
 sg13g2_fill_1 FILLER_57_157 ();
 sg13g2_fill_2 FILLER_57_175 ();
 sg13g2_fill_2 FILLER_57_202 ();
 sg13g2_fill_1 FILLER_57_204 ();
 sg13g2_fill_2 FILLER_57_219 ();
 sg13g2_decap_8 FILLER_57_247 ();
 sg13g2_fill_1 FILLER_57_254 ();
 sg13g2_decap_8 FILLER_57_258 ();
 sg13g2_fill_2 FILLER_57_265 ();
 sg13g2_decap_4 FILLER_57_272 ();
 sg13g2_fill_1 FILLER_57_276 ();
 sg13g2_fill_1 FILLER_57_291 ();
 sg13g2_fill_2 FILLER_57_326 ();
 sg13g2_fill_1 FILLER_57_336 ();
 sg13g2_fill_2 FILLER_57_350 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_fill_2 FILLER_58_186 ();
 sg13g2_decap_4 FILLER_58_237 ();
 sg13g2_fill_2 FILLER_58_241 ();
 sg13g2_fill_2 FILLER_58_252 ();
 sg13g2_fill_1 FILLER_58_264 ();
 sg13g2_fill_1 FILLER_58_307 ();
 sg13g2_fill_2 FILLER_58_384 ();
 sg13g2_fill_1 FILLER_58_386 ();
 sg13g2_fill_2 FILLER_58_406 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_fill_2 FILLER_59_131 ();
 sg13g2_fill_1 FILLER_59_146 ();
 sg13g2_fill_2 FILLER_59_220 ();
 sg13g2_fill_1 FILLER_59_222 ();
 sg13g2_fill_2 FILLER_59_237 ();
 sg13g2_fill_1 FILLER_59_239 ();
 sg13g2_fill_1 FILLER_59_281 ();
 sg13g2_fill_2 FILLER_59_297 ();
 sg13g2_fill_2 FILLER_59_308 ();
 sg13g2_fill_1 FILLER_59_310 ();
 sg13g2_fill_1 FILLER_59_316 ();
 sg13g2_decap_4 FILLER_59_335 ();
 sg13g2_fill_2 FILLER_59_339 ();
 sg13g2_decap_4 FILLER_59_345 ();
 sg13g2_fill_2 FILLER_59_365 ();
 sg13g2_fill_1 FILLER_59_367 ();
 sg13g2_fill_2 FILLER_59_407 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_4 FILLER_60_91 ();
 sg13g2_fill_2 FILLER_60_95 ();
 sg13g2_fill_2 FILLER_60_112 ();
 sg13g2_fill_1 FILLER_60_114 ();
 sg13g2_fill_1 FILLER_60_206 ();
 sg13g2_fill_2 FILLER_60_268 ();
 sg13g2_fill_1 FILLER_60_270 ();
 sg13g2_decap_8 FILLER_60_284 ();
 sg13g2_decap_8 FILLER_60_291 ();
 sg13g2_decap_8 FILLER_60_298 ();
 sg13g2_fill_2 FILLER_60_323 ();
 sg13g2_fill_1 FILLER_60_325 ();
 sg13g2_fill_1 FILLER_60_352 ();
 sg13g2_fill_1 FILLER_60_358 ();
 sg13g2_decap_8 FILLER_60_365 ();
 sg13g2_fill_2 FILLER_60_372 ();
 sg13g2_fill_1 FILLER_60_374 ();
 sg13g2_fill_1 FILLER_60_385 ();
 sg13g2_fill_1 FILLER_60_395 ();
 sg13g2_decap_8 FILLER_60_401 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_4 FILLER_61_84 ();
 sg13g2_fill_2 FILLER_61_119 ();
 sg13g2_fill_1 FILLER_61_121 ();
 sg13g2_fill_1 FILLER_61_144 ();
 sg13g2_fill_2 FILLER_61_216 ();
 sg13g2_fill_1 FILLER_61_218 ();
 sg13g2_decap_8 FILLER_61_245 ();
 sg13g2_decap_4 FILLER_61_252 ();
 sg13g2_decap_4 FILLER_61_260 ();
 sg13g2_decap_8 FILLER_61_268 ();
 sg13g2_fill_2 FILLER_61_275 ();
 sg13g2_fill_2 FILLER_61_294 ();
 sg13g2_decap_8 FILLER_61_306 ();
 sg13g2_decap_8 FILLER_61_313 ();
 sg13g2_decap_4 FILLER_61_320 ();
 sg13g2_fill_2 FILLER_61_324 ();
 sg13g2_decap_8 FILLER_61_331 ();
 sg13g2_decap_8 FILLER_61_338 ();
 sg13g2_decap_8 FILLER_61_345 ();
 sg13g2_fill_2 FILLER_61_352 ();
 sg13g2_decap_4 FILLER_61_381 ();
 sg13g2_fill_2 FILLER_61_395 ();
 sg13g2_decap_8 FILLER_61_401 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_4 FILLER_62_98 ();
 sg13g2_fill_2 FILLER_62_102 ();
 sg13g2_fill_2 FILLER_62_107 ();
 sg13g2_fill_1 FILLER_62_159 ();
 sg13g2_fill_2 FILLER_62_195 ();
 sg13g2_fill_1 FILLER_62_197 ();
 sg13g2_decap_8 FILLER_62_203 ();
 sg13g2_decap_4 FILLER_62_210 ();
 sg13g2_decap_4 FILLER_62_219 ();
 sg13g2_fill_1 FILLER_62_223 ();
 sg13g2_decap_8 FILLER_62_240 ();
 sg13g2_decap_8 FILLER_62_247 ();
 sg13g2_decap_4 FILLER_62_254 ();
 sg13g2_fill_2 FILLER_62_258 ();
 sg13g2_fill_1 FILLER_62_265 ();
 sg13g2_fill_2 FILLER_62_281 ();
 sg13g2_fill_1 FILLER_62_283 ();
 sg13g2_fill_2 FILLER_62_320 ();
 sg13g2_fill_1 FILLER_62_322 ();
 sg13g2_fill_2 FILLER_62_373 ();
 sg13g2_fill_1 FILLER_62_379 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_fill_2 FILLER_63_98 ();
 sg13g2_fill_1 FILLER_63_118 ();
 sg13g2_fill_1 FILLER_63_155 ();
 sg13g2_fill_2 FILLER_63_172 ();
 sg13g2_decap_8 FILLER_63_188 ();
 sg13g2_fill_2 FILLER_63_235 ();
 sg13g2_fill_1 FILLER_63_242 ();
 sg13g2_fill_2 FILLER_63_295 ();
 sg13g2_fill_2 FILLER_63_328 ();
 sg13g2_fill_1 FILLER_63_330 ();
 sg13g2_decap_8 FILLER_63_343 ();
 sg13g2_fill_2 FILLER_63_350 ();
 sg13g2_fill_2 FILLER_63_370 ();
 sg13g2_fill_1 FILLER_63_372 ();
 sg13g2_fill_1 FILLER_63_379 ();
 sg13g2_fill_1 FILLER_63_394 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_fill_2 FILLER_64_91 ();
 sg13g2_fill_1 FILLER_64_118 ();
 sg13g2_fill_2 FILLER_64_146 ();
 sg13g2_fill_1 FILLER_64_157 ();
 sg13g2_decap_4 FILLER_64_163 ();
 sg13g2_fill_1 FILLER_64_167 ();
 sg13g2_fill_1 FILLER_64_181 ();
 sg13g2_decap_8 FILLER_64_193 ();
 sg13g2_fill_2 FILLER_64_211 ();
 sg13g2_decap_4 FILLER_64_265 ();
 sg13g2_fill_2 FILLER_64_295 ();
 sg13g2_fill_1 FILLER_64_297 ();
 sg13g2_decap_4 FILLER_64_307 ();
 sg13g2_decap_4 FILLER_64_316 ();
 sg13g2_fill_2 FILLER_64_320 ();
 sg13g2_decap_8 FILLER_64_351 ();
 sg13g2_fill_1 FILLER_64_358 ();
 sg13g2_fill_2 FILLER_64_364 ();
 sg13g2_decap_4 FILLER_64_370 ();
 sg13g2_fill_1 FILLER_64_374 ();
 sg13g2_fill_1 FILLER_64_379 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_fill_2 FILLER_65_84 ();
 sg13g2_fill_1 FILLER_65_86 ();
 sg13g2_fill_2 FILLER_65_150 ();
 sg13g2_fill_1 FILLER_65_152 ();
 sg13g2_decap_4 FILLER_65_165 ();
 sg13g2_decap_4 FILLER_65_206 ();
 sg13g2_fill_1 FILLER_65_233 ();
 sg13g2_decap_4 FILLER_65_269 ();
 sg13g2_fill_2 FILLER_65_273 ();
 sg13g2_fill_2 FILLER_65_280 ();
 sg13g2_decap_8 FILLER_65_299 ();
 sg13g2_decap_4 FILLER_65_306 ();
 sg13g2_fill_1 FILLER_65_310 ();
 sg13g2_decap_8 FILLER_65_319 ();
 sg13g2_decap_8 FILLER_65_326 ();
 sg13g2_fill_2 FILLER_65_333 ();
 sg13g2_fill_2 FILLER_65_350 ();
 sg13g2_fill_2 FILLER_65_386 ();
 sg13g2_fill_1 FILLER_65_388 ();
 sg13g2_fill_2 FILLER_65_395 ();
 sg13g2_fill_1 FILLER_65_397 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_fill_1 FILLER_66_173 ();
 sg13g2_fill_1 FILLER_66_216 ();
 sg13g2_decap_8 FILLER_66_260 ();
 sg13g2_decap_8 FILLER_66_267 ();
 sg13g2_decap_4 FILLER_66_274 ();
 sg13g2_fill_1 FILLER_66_286 ();
 sg13g2_decap_4 FILLER_66_329 ();
 sg13g2_fill_1 FILLER_66_395 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_fill_2 FILLER_67_98 ();
 sg13g2_fill_1 FILLER_67_100 ();
 sg13g2_fill_1 FILLER_67_127 ();
 sg13g2_fill_1 FILLER_67_186 ();
 sg13g2_decap_8 FILLER_67_247 ();
 sg13g2_decap_4 FILLER_67_254 ();
 sg13g2_fill_2 FILLER_67_258 ();
 sg13g2_fill_2 FILLER_67_272 ();
 sg13g2_decap_8 FILLER_67_278 ();
 sg13g2_decap_4 FILLER_67_285 ();
 sg13g2_fill_1 FILLER_67_289 ();
 sg13g2_decap_4 FILLER_67_303 ();
 sg13g2_fill_1 FILLER_67_307 ();
 sg13g2_decap_4 FILLER_67_318 ();
 sg13g2_decap_8 FILLER_67_340 ();
 sg13g2_decap_8 FILLER_67_347 ();
 sg13g2_decap_8 FILLER_67_354 ();
 sg13g2_fill_2 FILLER_67_371 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_fill_2 FILLER_68_105 ();
 sg13g2_fill_1 FILLER_68_116 ();
 sg13g2_decap_8 FILLER_68_121 ();
 sg13g2_decap_4 FILLER_68_128 ();
 sg13g2_fill_2 FILLER_68_135 ();
 sg13g2_fill_2 FILLER_68_142 ();
 sg13g2_fill_2 FILLER_68_157 ();
 sg13g2_fill_2 FILLER_68_171 ();
 sg13g2_fill_2 FILLER_68_195 ();
 sg13g2_fill_2 FILLER_68_215 ();
 sg13g2_fill_1 FILLER_68_240 ();
 sg13g2_decap_4 FILLER_68_246 ();
 sg13g2_fill_2 FILLER_68_262 ();
 sg13g2_fill_2 FILLER_68_281 ();
 sg13g2_fill_1 FILLER_68_283 ();
 sg13g2_decap_8 FILLER_68_300 ();
 sg13g2_decap_8 FILLER_68_307 ();
 sg13g2_fill_2 FILLER_68_314 ();
 sg13g2_fill_2 FILLER_68_334 ();
 sg13g2_decap_8 FILLER_68_353 ();
 sg13g2_decap_4 FILLER_68_360 ();
 sg13g2_fill_2 FILLER_68_364 ();
 sg13g2_decap_4 FILLER_68_369 ();
 sg13g2_fill_2 FILLER_68_373 ();
 sg13g2_decap_4 FILLER_68_393 ();
 sg13g2_fill_1 FILLER_68_397 ();
 sg13g2_decap_4 FILLER_68_403 ();
 sg13g2_fill_2 FILLER_68_407 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_8 FILLER_69_119 ();
 sg13g2_decap_4 FILLER_69_126 ();
 sg13g2_fill_1 FILLER_69_130 ();
 sg13g2_fill_2 FILLER_69_173 ();
 sg13g2_fill_1 FILLER_69_217 ();
 sg13g2_fill_2 FILLER_69_308 ();
 sg13g2_fill_2 FILLER_69_318 ();
 sg13g2_fill_1 FILLER_69_320 ();
 sg13g2_decap_8 FILLER_69_360 ();
 sg13g2_decap_8 FILLER_69_367 ();
 sg13g2_decap_8 FILLER_69_374 ();
 sg13g2_fill_2 FILLER_69_381 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_fill_2 FILLER_70_119 ();
 sg13g2_fill_1 FILLER_70_130 ();
 sg13g2_decap_8 FILLER_70_236 ();
 sg13g2_decap_8 FILLER_70_243 ();
 sg13g2_fill_2 FILLER_70_283 ();
 sg13g2_decap_8 FILLER_70_312 ();
 sg13g2_decap_8 FILLER_70_319 ();
 sg13g2_decap_8 FILLER_70_326 ();
 sg13g2_decap_8 FILLER_70_333 ();
 sg13g2_fill_1 FILLER_70_340 ();
 sg13g2_fill_1 FILLER_70_348 ();
 sg13g2_decap_4 FILLER_70_361 ();
 sg13g2_fill_2 FILLER_70_370 ();
 sg13g2_decap_8 FILLER_70_377 ();
 sg13g2_decap_8 FILLER_70_384 ();
 sg13g2_decap_8 FILLER_70_391 ();
 sg13g2_decap_8 FILLER_70_398 ();
 sg13g2_decap_4 FILLER_70_405 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_4 FILLER_71_105 ();
 sg13g2_fill_2 FILLER_71_135 ();
 sg13g2_fill_2 FILLER_71_182 ();
 sg13g2_fill_1 FILLER_71_193 ();
 sg13g2_decap_4 FILLER_71_231 ();
 sg13g2_fill_2 FILLER_71_238 ();
 sg13g2_fill_2 FILLER_71_249 ();
 sg13g2_fill_1 FILLER_71_251 ();
 sg13g2_fill_1 FILLER_71_271 ();
 sg13g2_fill_2 FILLER_71_298 ();
 sg13g2_decap_8 FILLER_71_326 ();
 sg13g2_decap_8 FILLER_71_333 ();
 sg13g2_decap_4 FILLER_71_340 ();
 sg13g2_fill_1 FILLER_71_344 ();
 sg13g2_fill_2 FILLER_71_355 ();
 sg13g2_fill_2 FILLER_71_385 ();
 sg13g2_fill_2 FILLER_71_392 ();
 sg13g2_decap_8 FILLER_71_400 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_4 FILLER_72_98 ();
 sg13g2_fill_2 FILLER_72_167 ();
 sg13g2_fill_1 FILLER_72_169 ();
 sg13g2_fill_1 FILLER_72_201 ();
 sg13g2_fill_2 FILLER_72_216 ();
 sg13g2_fill_1 FILLER_72_286 ();
 sg13g2_fill_1 FILLER_72_293 ();
 sg13g2_fill_1 FILLER_72_344 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_4 FILLER_73_105 ();
 sg13g2_fill_1 FILLER_73_109 ();
 sg13g2_fill_1 FILLER_73_154 ();
 sg13g2_fill_2 FILLER_73_181 ();
 sg13g2_fill_2 FILLER_73_206 ();
 sg13g2_decap_8 FILLER_73_246 ();
 sg13g2_fill_2 FILLER_73_253 ();
 sg13g2_decap_4 FILLER_73_270 ();
 sg13g2_fill_2 FILLER_73_280 ();
 sg13g2_fill_1 FILLER_73_296 ();
 sg13g2_decap_8 FILLER_73_308 ();
 sg13g2_fill_2 FILLER_73_315 ();
 sg13g2_fill_1 FILLER_73_317 ();
 sg13g2_fill_1 FILLER_73_344 ();
 sg13g2_fill_2 FILLER_73_363 ();
 sg13g2_fill_1 FILLER_73_365 ();
 sg13g2_fill_2 FILLER_73_392 ();
 sg13g2_fill_1 FILLER_73_394 ();
 sg13g2_decap_4 FILLER_73_405 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_4 FILLER_74_112 ();
 sg13g2_decap_4 FILLER_74_254 ();
 sg13g2_fill_1 FILLER_74_258 ();
 sg13g2_decap_4 FILLER_74_263 ();
 sg13g2_fill_2 FILLER_74_267 ();
 sg13g2_fill_2 FILLER_74_274 ();
 sg13g2_fill_2 FILLER_74_287 ();
 sg13g2_decap_8 FILLER_74_298 ();
 sg13g2_decap_4 FILLER_74_305 ();
 sg13g2_fill_1 FILLER_74_309 ();
 sg13g2_decap_8 FILLER_74_316 ();
 sg13g2_fill_1 FILLER_74_331 ();
 sg13g2_decap_8 FILLER_74_354 ();
 sg13g2_fill_2 FILLER_74_361 ();
 sg13g2_fill_1 FILLER_74_363 ();
 sg13g2_fill_1 FILLER_74_389 ();
 sg13g2_fill_1 FILLER_74_395 ();
 sg13g2_decap_8 FILLER_74_401 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_4 FILLER_75_105 ();
 sg13g2_fill_1 FILLER_75_109 ();
 sg13g2_fill_1 FILLER_75_172 ();
 sg13g2_fill_2 FILLER_75_182 ();
 sg13g2_fill_2 FILLER_75_193 ();
 sg13g2_fill_1 FILLER_75_195 ();
 sg13g2_fill_2 FILLER_75_269 ();
 sg13g2_fill_1 FILLER_75_271 ();
 sg13g2_fill_1 FILLER_75_289 ();
 sg13g2_fill_2 FILLER_75_310 ();
 sg13g2_fill_1 FILLER_75_312 ();
 sg13g2_decap_8 FILLER_75_322 ();
 sg13g2_decap_8 FILLER_75_329 ();
 sg13g2_decap_8 FILLER_75_336 ();
 sg13g2_fill_2 FILLER_75_343 ();
 sg13g2_fill_1 FILLER_75_345 ();
 sg13g2_fill_1 FILLER_75_355 ();
 sg13g2_fill_2 FILLER_75_365 ();
 sg13g2_fill_1 FILLER_75_376 ();
 sg13g2_fill_1 FILLER_75_391 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_fill_1 FILLER_76_143 ();
 sg13g2_fill_2 FILLER_76_174 ();
 sg13g2_fill_1 FILLER_76_293 ();
 sg13g2_decap_8 FILLER_76_322 ();
 sg13g2_decap_8 FILLER_76_329 ();
 sg13g2_fill_1 FILLER_76_336 ();
 sg13g2_fill_2 FILLER_76_356 ();
 sg13g2_fill_1 FILLER_76_367 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_4 FILLER_77_105 ();
 sg13g2_fill_2 FILLER_77_255 ();
 sg13g2_fill_1 FILLER_77_301 ();
 sg13g2_fill_2 FILLER_77_332 ();
 sg13g2_fill_1 FILLER_77_344 ();
 sg13g2_fill_2 FILLER_77_368 ();
 sg13g2_fill_1 FILLER_77_370 ();
 sg13g2_fill_2 FILLER_77_385 ();
 sg13g2_decap_8 FILLER_77_396 ();
 sg13g2_decap_4 FILLER_77_403 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_fill_2 FILLER_78_119 ();
 sg13g2_fill_2 FILLER_78_132 ();
 sg13g2_fill_2 FILLER_78_266 ();
 sg13g2_fill_1 FILLER_78_268 ();
 sg13g2_fill_1 FILLER_78_370 ();
 sg13g2_decap_8 FILLER_78_398 ();
 sg13g2_decap_4 FILLER_78_405 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_4 FILLER_79_112 ();
 sg13g2_fill_1 FILLER_79_158 ();
 sg13g2_fill_1 FILLER_79_185 ();
 sg13g2_fill_1 FILLER_79_219 ();
 sg13g2_fill_1 FILLER_79_268 ();
 sg13g2_decap_4 FILLER_79_287 ();
 sg13g2_fill_1 FILLER_79_291 ();
 sg13g2_fill_2 FILLER_79_313 ();
 sg13g2_fill_1 FILLER_79_366 ();
 sg13g2_fill_1 FILLER_79_382 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_8 FILLER_80_116 ();
 sg13g2_decap_8 FILLER_80_123 ();
 sg13g2_fill_2 FILLER_80_151 ();
 sg13g2_fill_1 FILLER_80_153 ();
 sg13g2_fill_2 FILLER_80_208 ();
 sg13g2_decap_8 FILLER_80_255 ();
 sg13g2_decap_8 FILLER_80_262 ();
 sg13g2_decap_8 FILLER_80_269 ();
 sg13g2_decap_8 FILLER_80_276 ();
 sg13g2_decap_4 FILLER_80_283 ();
 sg13g2_fill_1 FILLER_80_287 ();
 sg13g2_decap_4 FILLER_80_292 ();
 sg13g2_fill_2 FILLER_80_301 ();
 sg13g2_fill_1 FILLER_80_303 ();
 sg13g2_fill_2 FILLER_80_317 ();
 sg13g2_fill_1 FILLER_80_319 ();
 sg13g2_fill_2 FILLER_80_325 ();
 sg13g2_fill_1 FILLER_80_327 ();
 sg13g2_decap_4 FILLER_80_332 ();
 sg13g2_fill_2 FILLER_80_341 ();
 sg13g2_fill_1 FILLER_80_343 ();
 sg13g2_fill_2 FILLER_80_349 ();
 sg13g2_fill_1 FILLER_80_351 ();
 sg13g2_fill_2 FILLER_80_357 ();
 sg13g2_fill_1 FILLER_80_359 ();
 sg13g2_fill_2 FILLER_80_365 ();
 sg13g2_fill_1 FILLER_80_367 ();
 sg13g2_decap_8 FILLER_80_381 ();
 sg13g2_decap_8 FILLER_80_388 ();
 sg13g2_decap_8 FILLER_80_395 ();
 sg13g2_decap_8 FILLER_80_402 ();
 assign uio_oe[0] = net12;
 assign uio_oe[1] = net13;
 assign uio_oe[2] = net14;
 assign uio_oe[3] = net18;
 assign uio_oe[4] = net19;
 assign uio_oe[5] = net20;
 assign uio_oe[6] = net21;
 assign uio_oe[7] = net22;
 assign uio_out[0] = net15;
 assign uio_out[1] = net16;
 assign uio_out[2] = net17;
endmodule

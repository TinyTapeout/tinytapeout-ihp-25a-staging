module tt_um_wokwi_group_4 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire \proj_10.net10 ;
 wire \proj_10.net11 ;
 wire \proj_10.net14 ;
 wire \proj_10.net4 ;
 wire \proj_10.net5 ;
 wire \proj_11.net15 ;
 wire \proj_11.net16 ;
 wire \proj_11.net17 ;
 wire \proj_11.net18 ;
 wire \proj_11.net6 ;
 wire \proj_11.net7 ;
 wire \proj_11.net8 ;
 wire \proj_11.net9 ;
 wire \proj_12.net3 ;
 wire \proj_12.net4 ;
 wire \proj_13.net10 ;
 wire \proj_13.net11 ;
 wire \proj_13.net8 ;
 wire \proj_13.net9 ;
 wire \proj_14.net14 ;
 wire \proj_14.net15 ;
 wire \proj_14.net16 ;
 wire \proj_14.net17 ;
 wire \proj_14.net18 ;
 wire \proj_14.net19 ;
 wire \proj_14.net20 ;
 wire \proj_14.net6 ;
 wire \proj_14.net7 ;
 wire \proj_14.net8 ;
 wire \proj_15.net3 ;
 wire \proj_15.net4 ;
 wire \proj_15.net6 ;
 wire \proj_15.net7 ;
 wire \proj__0.net10 ;
 wire \proj__0.net11 ;
 wire \proj__0.net12 ;
 wire \proj__0.net13 ;
 wire \proj__1.net4 ;
 wire \proj__1.net5 ;
 wire \proj__1.net6 ;
 wire \proj__1.net7 ;
 wire \proj__1.net8 ;
 wire \proj__1.net9 ;
 wire \proj__2.net10 ;
 wire \proj__2.net11 ;
 wire \proj__2.net12 ;
 wire \proj__2.net9 ;
 wire \proj__3.net10 ;
 wire \proj__3.net11 ;
 wire \proj__3.net12 ;
 wire \proj__3.net13 ;
 wire \proj__3.net14 ;
 wire \proj__3.net20 ;
 wire \proj__3.net9 ;
 wire \proj__4.net10 ;
 wire \proj__4.net11 ;
 wire \proj__4.net12 ;
 wire \proj__4.net13 ;
 wire \proj__5.net10 ;
 wire \proj__5.net9 ;
 wire \proj__6.net10 ;
 wire \proj__6.net100 ;
 wire \proj__6.net101 ;
 wire \proj__6.net102 ;
 wire \proj__6.net103 ;
 wire \proj__6.net104 ;
 wire \proj__6.net105 ;
 wire \proj__6.net106 ;
 wire \proj__6.net107 ;
 wire \proj__6.net108 ;
 wire \proj__6.net109 ;
 wire \proj__6.net11 ;
 wire \proj__6.net110 ;
 wire \proj__6.net111 ;
 wire \proj__6.net112 ;
 wire \proj__6.net113 ;
 wire \proj__6.net114 ;
 wire \proj__6.net115 ;
 wire \proj__6.net116 ;
 wire \proj__6.net117 ;
 wire \proj__6.net118 ;
 wire \proj__6.net119 ;
 wire \proj__6.net12 ;
 wire \proj__6.net120 ;
 wire \proj__6.net121 ;
 wire \proj__6.net122 ;
 wire \proj__6.net123 ;
 wire \proj__6.net124 ;
 wire \proj__6.net125 ;
 wire \proj__6.net126 ;
 wire \proj__6.net127 ;
 wire \proj__6.net128 ;
 wire \proj__6.net129 ;
 wire \proj__6.net13 ;
 wire \proj__6.net130 ;
 wire \proj__6.net131 ;
 wire \proj__6.net132 ;
 wire \proj__6.net133 ;
 wire \proj__6.net134 ;
 wire \proj__6.net135 ;
 wire \proj__6.net136 ;
 wire \proj__6.net137 ;
 wire \proj__6.net138 ;
 wire \proj__6.net139 ;
 wire \proj__6.net14 ;
 wire \proj__6.net140 ;
 wire \proj__6.net141 ;
 wire \proj__6.net142 ;
 wire \proj__6.net143 ;
 wire \proj__6.net144 ;
 wire \proj__6.net145 ;
 wire \proj__6.net146 ;
 wire \proj__6.net147 ;
 wire \proj__6.net148 ;
 wire \proj__6.net149 ;
 wire \proj__6.net15 ;
 wire \proj__6.net150 ;
 wire \proj__6.net151 ;
 wire \proj__6.net152 ;
 wire \proj__6.net153 ;
 wire \proj__6.net154 ;
 wire \proj__6.net155 ;
 wire \proj__6.net156 ;
 wire \proj__6.net157 ;
 wire \proj__6.net158 ;
 wire \proj__6.net159 ;
 wire \proj__6.net16 ;
 wire \proj__6.net160 ;
 wire \proj__6.net161 ;
 wire \proj__6.net162 ;
 wire \proj__6.net163 ;
 wire \proj__6.net164 ;
 wire \proj__6.net165 ;
 wire \proj__6.net166 ;
 wire \proj__6.net167 ;
 wire \proj__6.net168 ;
 wire \proj__6.net169 ;
 wire \proj__6.net170 ;
 wire \proj__6.net171 ;
 wire \proj__6.net172 ;
 wire \proj__6.net173 ;
 wire \proj__6.net174 ;
 wire \proj__6.net175 ;
 wire \proj__6.net176 ;
 wire \proj__6.net177 ;
 wire \proj__6.net178 ;
 wire \proj__6.net179 ;
 wire \proj__6.net180 ;
 wire \proj__6.net181 ;
 wire \proj__6.net182 ;
 wire \proj__6.net183 ;
 wire \proj__6.net184 ;
 wire \proj__6.net185 ;
 wire \proj__6.net186 ;
 wire \proj__6.net187 ;
 wire \proj__6.net188 ;
 wire \proj__6.net189 ;
 wire \proj__6.net190 ;
 wire \proj__6.net191 ;
 wire \proj__6.net192 ;
 wire \proj__6.net193 ;
 wire \proj__6.net194 ;
 wire \proj__6.net195 ;
 wire \proj__6.net22 ;
 wire \proj__6.net23 ;
 wire \proj__6.net24 ;
 wire \proj__6.net25 ;
 wire \proj__6.net26 ;
 wire \proj__6.net27 ;
 wire \proj__6.net28 ;
 wire \proj__6.net29 ;
 wire \proj__6.net30 ;
 wire \proj__6.net31 ;
 wire \proj__6.net32 ;
 wire \proj__6.net33 ;
 wire \proj__6.net34 ;
 wire \proj__6.net35 ;
 wire \proj__6.net36 ;
 wire \proj__6.net37 ;
 wire \proj__6.net38 ;
 wire \proj__6.net39 ;
 wire \proj__6.net40 ;
 wire \proj__6.net41 ;
 wire \proj__6.net42 ;
 wire \proj__6.net43 ;
 wire \proj__6.net44 ;
 wire \proj__6.net45 ;
 wire \proj__6.net46 ;
 wire \proj__6.net47 ;
 wire \proj__6.net48 ;
 wire \proj__6.net49 ;
 wire \proj__6.net50 ;
 wire \proj__6.net51 ;
 wire \proj__6.net52 ;
 wire \proj__6.net53 ;
 wire \proj__6.net54 ;
 wire \proj__6.net55 ;
 wire \proj__6.net56 ;
 wire \proj__6.net57 ;
 wire \proj__6.net58 ;
 wire \proj__6.net59 ;
 wire \proj__6.net60 ;
 wire \proj__6.net61 ;
 wire \proj__6.net62 ;
 wire \proj__6.net63 ;
 wire \proj__6.net64 ;
 wire \proj__6.net65 ;
 wire \proj__6.net66 ;
 wire \proj__6.net67 ;
 wire \proj__6.net68 ;
 wire \proj__6.net69 ;
 wire \proj__6.net70 ;
 wire \proj__6.net71 ;
 wire \proj__6.net72 ;
 wire \proj__6.net73 ;
 wire \proj__6.net74 ;
 wire \proj__6.net75 ;
 wire \proj__6.net76 ;
 wire \proj__6.net77 ;
 wire \proj__6.net78 ;
 wire \proj__6.net79 ;
 wire \proj__6.net80 ;
 wire \proj__6.net81 ;
 wire \proj__6.net82 ;
 wire \proj__6.net83 ;
 wire \proj__6.net84 ;
 wire \proj__6.net85 ;
 wire \proj__6.net86 ;
 wire \proj__6.net87 ;
 wire \proj__6.net88 ;
 wire \proj__6.net89 ;
 wire \proj__6.net9 ;
 wire \proj__6.net90 ;
 wire \proj__6.net91 ;
 wire \proj__6.net92 ;
 wire \proj__6.net93 ;
 wire \proj__6.net94 ;
 wire \proj__6.net95 ;
 wire \proj__6.net96 ;
 wire \proj__6.net97 ;
 wire \proj__6.net98 ;
 wire \proj__6.net99 ;
 wire \proj__7.net7 ;
 wire \proj__8.net10 ;
 wire \proj__8.net11 ;
 wire \proj__8.net12 ;
 wire \proj__8.net13 ;
 wire \proj__8.net14 ;
 wire \proj__8.net15 ;
 wire \proj__8.net18 ;
 wire \proj__8.net19 ;
 wire \proj__8.net20 ;
 wire \proj__8.net21 ;
 wire \proj__8.net22 ;
 wire \proj__8.net23 ;
 wire \proj__8.net24 ;
 wire \proj__8.net25 ;
 wire \proj__8.net26 ;
 wire \proj__8.net27 ;
 wire \proj__8.net28 ;
 wire \proj__8.net29 ;
 wire \proj__8.net30 ;
 wire \proj__8.net31 ;
 wire \proj__8.net32 ;
 wire \proj__8.net33 ;
 wire \proj__8.net34 ;
 wire \proj__8.net35 ;
 wire \proj__8.net36 ;
 wire \proj__8.net37 ;
 wire \proj__8.net38 ;
 wire \proj__8.net39 ;
 wire \proj__8.net40 ;
 wire \proj__8.net9 ;
 wire \proj__9.net10 ;
 wire \proj__9.net11 ;
 wire \proj__9.net12 ;
 wire \proj__9.net13 ;
 wire \proj__9.net19 ;
 wire \proj__9.net20 ;
 wire \proj__9.net21 ;
 wire \proj__9.net22 ;
 wire \proj__9.net23 ;
 wire \proj__9.net24 ;
 wire \proj__9.net25 ;
 wire \proj__9.net26 ;
 wire \proj__9.net27 ;
 wire \proj__9.net28 ;
 wire \proj__9.net29 ;
 wire \proj__9.net30 ;
 wire \proj__9.net9 ;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire \proj__1.flop1/notq ;
 wire net35;
 wire \proj__1.flop2/notq ;
 wire net36;
 wire \proj__1.flop3/notq ;
 wire net37;
 wire \proj__1.flop4/notq ;
 wire net38;
 wire \proj__1.flop5/notq ;
 wire net39;
 wire \proj__1.flop6/notq ;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;

 sg13g2_inv_1 _094_ (.Y(_066_),
    .A(net3));
 sg13g2_inv_2 _095_ (.Y(_067_),
    .A(net6));
 sg13g2_inv_1 _096_ (.Y(_068_),
    .A(net5));
 sg13g2_inv_1 _097_ (.Y(_069_),
    .A(\proj__0.net10 ));
 sg13g2_inv_1 _098_ (.Y(_070_),
    .A(\proj__0.net11 ));
 sg13g2_inv_1 _099_ (.Y(_071_),
    .A(\proj__0.net12 ));
 sg13g2_inv_1 _100_ (.Y(_072_),
    .A(\proj__0.net13 ));
 sg13g2_nor2_2 _101_ (.A(net6),
    .B(net5),
    .Y(_073_));
 sg13g2_nor2b_1 _102_ (.A(net107),
    .B_N(net3),
    .Y(_074_));
 sg13g2_and2_2 _103_ (.A(_073_),
    .B(_074_),
    .X(_075_));
 sg13g2_nor2b_2 _104_ (.A(net6),
    .B_N(net5),
    .Y(_076_));
 sg13g2_inv_1 _105_ (.Y(_077_),
    .A(_076_));
 sg13g2_and2_2 _106_ (.A(_074_),
    .B(_076_),
    .X(_078_));
 sg13g2_nor2_1 _107_ (.A(net3),
    .B(net107),
    .Y(_079_));
 sg13g2_and2_2 _108_ (.A(_076_),
    .B(_079_),
    .X(_080_));
 sg13g2_and2_1 _109_ (.A(net3),
    .B(net107),
    .X(_081_));
 sg13g2_and2_1 _110_ (.A(_076_),
    .B(_081_),
    .X(_082_));
 sg13g2_a22oi_1 _111_ (.Y(_083_),
    .B1(_076_),
    .B2(_081_),
    .A2(_073_),
    .A1(_066_));
 sg13g2_inv_1 _112_ (.Y(_000_),
    .A(_083_));
 sg13g2_o21ai_1 _113_ (.B1(_083_),
    .Y(_001_),
    .A1(net107),
    .A2(_077_));
 sg13g2_o21ai_1 _114_ (.B1(net109),
    .Y(_002_),
    .A1(_075_),
    .A2(_001_));
 sg13g2_nor4_2 _115_ (.A(_066_),
    .B(net4),
    .C(_067_),
    .Y(_003_),
    .D(_068_));
 sg13g2_nand2_1 _116_ (.Y(_004_),
    .A(\proj_13.net11 ),
    .B(_003_));
 sg13g2_nand3_1 _117_ (.B(net107),
    .C(net6),
    .A(net3),
    .Y(_005_));
 sg13g2_nor2_1 _118_ (.A(_068_),
    .B(_005_),
    .Y(_006_));
 sg13g2_nand2_1 _119_ (.Y(_007_),
    .A(\proj_15.net4 ),
    .B(_006_));
 sg13g2_and2_2 _120_ (.A(_073_),
    .B(_081_),
    .X(_008_));
 sg13g2_nor2b_2 _121_ (.A(net3),
    .B_N(net107),
    .Y(_009_));
 sg13g2_and2_2 _122_ (.A(_076_),
    .B(_009_),
    .X(_010_));
 sg13g2_a22oi_1 _123_ (.Y(_011_),
    .B1(_010_),
    .B2(\proj__6.net16 ),
    .A2(_008_),
    .A1(\proj__3.net14 ));
 sg13g2_nand4_1 _124_ (.B(_004_),
    .C(_007_),
    .A(_002_),
    .Y(uo_out[7]),
    .D(_011_));
 sg13g2_and2_2 _125_ (.A(_073_),
    .B(_079_),
    .X(_012_));
 sg13g2_nor2_2 _126_ (.A(net5),
    .B(_005_),
    .Y(_013_));
 sg13g2_nor4_2 _127_ (.A(_066_),
    .B(net107),
    .C(_067_),
    .Y(_014_),
    .D(net5));
 sg13g2_nand2_1 _128_ (.Y(_015_),
    .A(\proj__9.net9 ),
    .B(_014_));
 sg13g2_nor4_2 _129_ (.A(net3),
    .B(net107),
    .C(_067_),
    .Y(_016_),
    .D(net5));
 sg13g2_and3_1 _130_ (.X(_017_),
    .A(net6),
    .B(net5),
    .C(_009_));
 sg13g2_nor4_2 _131_ (.A(net3),
    .B(net4),
    .C(_067_),
    .Y(_018_),
    .D(_068_));
 sg13g2_a22oi_1 _132_ (.Y(_019_),
    .B1(_018_),
    .B2(\proj_12.net3 ),
    .A2(_003_),
    .A1(\proj_13.net8 ));
 sg13g2_and3_1 _133_ (.X(_020_),
    .A(net6),
    .B(_068_),
    .C(_009_));
 sg13g2_a22oi_1 _134_ (.Y(_021_),
    .B1(_008_),
    .B2(\proj__3.net9 ),
    .A2(_082_),
    .A1(\proj__7.net7 ));
 sg13g2_and2_2 _135_ (.A(_073_),
    .B(_009_),
    .X(_022_));
 sg13g2_a22oi_1 _136_ (.Y(_023_),
    .B1(_022_),
    .B2(\proj__2.net9 ),
    .A2(_075_),
    .A1(\proj__1.net4 ));
 sg13g2_a22oi_1 _137_ (.Y(_024_),
    .B1(_017_),
    .B2(\proj_14.net6 ),
    .A2(_080_),
    .A1(\proj__4.net10 ));
 sg13g2_and4_1 _138_ (.A(_015_),
    .B(_021_),
    .C(_023_),
    .D(_024_),
    .X(_025_));
 sg13g2_a22oi_1 _139_ (.Y(_026_),
    .B1(_020_),
    .B2(\proj_10.net4 ),
    .A2(_013_),
    .A1(\proj_11.net6 ));
 sg13g2_a221oi_1 _140_ (.B2(\proj__6.net9 ),
    .C1(_012_),
    .B1(_010_),
    .A1(\proj__5.net9 ),
    .Y(_027_),
    .A2(_078_));
 sg13g2_a22oi_1 _141_ (.Y(_028_),
    .B1(_016_),
    .B2(\proj__8.net9 ),
    .A2(_006_),
    .A1(\proj_15.net3 ));
 sg13g2_and4_1 _142_ (.A(_019_),
    .B(_026_),
    .C(_027_),
    .D(_028_),
    .X(_029_));
 sg13g2_a22oi_1 _143_ (.Y(uo_out[0]),
    .B1(_025_),
    .B2(_029_),
    .A2(_012_),
    .A1(_069_));
 sg13g2_nand2_1 _144_ (.Y(_030_),
    .A(\proj_12.net4 ),
    .B(_018_));
 sg13g2_nand2_1 _145_ (.Y(_031_),
    .A(\proj_13.net9 ),
    .B(_003_));
 sg13g2_a22oi_1 _146_ (.Y(_032_),
    .B1(_020_),
    .B2(\proj_10.net5 ),
    .A2(_013_),
    .A1(\proj_11.net7 ));
 sg13g2_a22oi_1 _147_ (.Y(_033_),
    .B1(_022_),
    .B2(\proj__2.net10 ),
    .A2(_008_),
    .A1(\proj__3.net10 ));
 sg13g2_a21oi_1 _148_ (.A1(\proj__6.net10 ),
    .A2(_010_),
    .Y(_034_),
    .B1(_012_));
 sg13g2_and4_1 _149_ (.A(_030_),
    .B(_031_),
    .C(_033_),
    .D(_034_),
    .X(_035_));
 sg13g2_a22oi_1 _150_ (.Y(_036_),
    .B1(_017_),
    .B2(\proj_14.net7 ),
    .A2(_014_),
    .A1(\proj__9.net10 ));
 sg13g2_a22oi_1 _151_ (.Y(_037_),
    .B1(_080_),
    .B2(net125),
    .A2(_078_),
    .A1(\proj__5.net10 ));
 sg13g2_a22oi_1 _152_ (.Y(_038_),
    .B1(_016_),
    .B2(\proj__8.net10 ),
    .A2(_075_),
    .A1(\proj__1.net5 ));
 sg13g2_and4_1 _153_ (.A(_032_),
    .B(_036_),
    .C(_037_),
    .D(_038_),
    .X(_039_));
 sg13g2_a22oi_1 _154_ (.Y(uo_out[1]),
    .B1(_035_),
    .B2(_039_),
    .A2(_012_),
    .A1(_070_));
 sg13g2_nand2_1 _155_ (.Y(_040_),
    .A(\proj__8.net11 ),
    .B(_016_));
 sg13g2_a22oi_1 _156_ (.Y(_041_),
    .B1(_017_),
    .B2(\proj_14.net8 ),
    .A2(_014_),
    .A1(\proj__9.net11 ));
 sg13g2_and2_1 _157_ (.A(_040_),
    .B(_041_),
    .X(_042_));
 sg13g2_a22oi_1 _158_ (.Y(_043_),
    .B1(_008_),
    .B2(\proj__3.net11 ),
    .A2(_003_),
    .A1(\proj_13.net10 ));
 sg13g2_a22oi_1 _159_ (.Y(_044_),
    .B1(_022_),
    .B2(\proj__2.net11 ),
    .A2(_080_),
    .A1(\proj__4.net11 ));
 sg13g2_a22oi_1 _160_ (.Y(_045_),
    .B1(_010_),
    .B2(\proj__6.net11 ),
    .A2(_075_),
    .A1(\proj__1.net6 ));
 sg13g2_a221oi_1 _161_ (.B2(\proj_11.net8 ),
    .C1(_012_),
    .B1(_013_),
    .A1(\proj__5.net10 ),
    .Y(_046_),
    .A2(_078_));
 sg13g2_and4_1 _162_ (.A(_043_),
    .B(_044_),
    .C(_045_),
    .D(_046_),
    .X(_047_));
 sg13g2_a22oi_1 _163_ (.Y(uo_out[2]),
    .B1(_042_),
    .B2(_047_),
    .A2(_012_),
    .A1(_071_));
 sg13g2_a221oi_1 _164_ (.B2(\proj__9.net12 ),
    .C1(_012_),
    .B1(_014_),
    .A1(\proj__5.net9 ),
    .Y(_048_),
    .A2(_078_));
 sg13g2_a22oi_1 _165_ (.Y(_049_),
    .B1(_016_),
    .B2(\proj__8.net12 ),
    .A2(_013_),
    .A1(\proj_11.net9 ));
 sg13g2_and2_1 _166_ (.A(_048_),
    .B(_049_),
    .X(_050_));
 sg13g2_nand2_1 _167_ (.Y(_051_),
    .A(\proj__6.net12 ),
    .B(_010_));
 sg13g2_a22oi_1 _168_ (.Y(_052_),
    .B1(_080_),
    .B2(\proj__4.net12 ),
    .A2(_075_),
    .A1(\proj__1.net7 ));
 sg13g2_a22oi_1 _169_ (.Y(_053_),
    .B1(_022_),
    .B2(\proj__2.net12 ),
    .A2(_008_),
    .A1(\proj__3.net12 ));
 sg13g2_and4_1 _170_ (.A(_004_),
    .B(_051_),
    .C(_052_),
    .D(_053_),
    .X(_054_));
 sg13g2_a22oi_1 _171_ (.Y(uo_out[3]),
    .B1(_050_),
    .B2(_054_),
    .A2(_012_),
    .A1(_072_));
 sg13g2_a22oi_1 _172_ (.Y(_055_),
    .B1(_016_),
    .B2(\proj__8.net13 ),
    .A2(_014_),
    .A1(\proj__9.net13 ));
 sg13g2_a22oi_1 _173_ (.Y(_056_),
    .B1(_078_),
    .B2(net113),
    .A2(_075_),
    .A1(\proj__1.net8 ));
 sg13g2_a22oi_1 _174_ (.Y(_057_),
    .B1(_010_),
    .B2(\proj__6.net13 ),
    .A2(_080_),
    .A1(\proj__4.net13 ));
 sg13g2_nand4_1 _175_ (.B(_055_),
    .C(_056_),
    .A(_043_),
    .Y(_058_),
    .D(_057_));
 sg13g2_a21o_1 _176_ (.A2(_000_),
    .A1(net115),
    .B1(_058_),
    .X(uo_out[4]));
 sg13g2_o21ai_1 _177_ (.B1(net113),
    .Y(_059_),
    .A1(_080_),
    .A2(_000_));
 sg13g2_a22oi_1 _178_ (.Y(_060_),
    .B1(_016_),
    .B2(\proj__8.net14 ),
    .A2(_003_),
    .A1(\proj_13.net8 ));
 sg13g2_a22oi_1 _179_ (.Y(_061_),
    .B1(_008_),
    .B2(\proj__3.net10 ),
    .A2(_075_),
    .A1(\proj__1.net9 ));
 sg13g2_a22oi_1 _180_ (.Y(_062_),
    .B1(_010_),
    .B2(\proj__6.net14 ),
    .A2(_078_),
    .A1(net114));
 sg13g2_nand4_1 _181_ (.B(_060_),
    .C(_061_),
    .A(_059_),
    .Y(uo_out[5]),
    .D(_062_));
 sg13g2_nand2_1 _182_ (.Y(_063_),
    .A(net110),
    .B(_001_));
 sg13g2_a22oi_1 _183_ (.Y(_064_),
    .B1(_008_),
    .B2(\proj__3.net13 ),
    .A2(_003_),
    .A1(\proj_13.net9 ));
 sg13g2_a22oi_1 _184_ (.Y(_065_),
    .B1(_016_),
    .B2(\proj__8.net15 ),
    .A2(_010_),
    .A1(\proj__6.net15 ));
 sg13g2_nand3_1 _185_ (.B(_064_),
    .C(_065_),
    .A(_063_),
    .Y(uo_out[6]));
 sg13g2_tielo \proj_15.gate8/_0__8  (.L_LO(net8));
 sg13g2_tielo \proj__0.and2/_0__9  (.L_LO(net9));
 sg13g2_tielo \proj__1.flop1/_1__10  (.L_LO(net10));
 sg13g2_tielo \proj__1.flop2/_1__11  (.L_LO(net11));
 sg13g2_tielo \proj__1.flop3/_1__12  (.L_LO(net12));
 sg13g2_tielo \proj__1.flop4/_1__13  (.L_LO(net13));
 sg13g2_tielo \proj__1.flop5/_1__14  (.L_LO(net14));
 sg13g2_tielo \proj__1.flop6/_1__15  (.L_LO(net15));
 sg13g2_tielo \proj__4.nand1/_0__16  (.L_LO(net16));
 sg13g2_tielo tt_um_wokwi_group_4_17 (.L_LO(net17));
 sg13g2_tielo tt_um_wokwi_group_4_18 (.L_LO(net18));
 sg13g2_tielo tt_um_wokwi_group_4_19 (.L_LO(net19));
 sg13g2_tielo tt_um_wokwi_group_4_20 (.L_LO(net20));
 sg13g2_tielo tt_um_wokwi_group_4_21 (.L_LO(net21));
 sg13g2_tielo tt_um_wokwi_group_4_22 (.L_LO(net22));
 sg13g2_tielo tt_um_wokwi_group_4_23 (.L_LO(net23));
 sg13g2_tielo tt_um_wokwi_group_4_24 (.L_LO(net24));
 sg13g2_tielo tt_um_wokwi_group_4_25 (.L_LO(net25));
 sg13g2_tielo tt_um_wokwi_group_4_26 (.L_LO(net26));
 sg13g2_tielo tt_um_wokwi_group_4_27 (.L_LO(net27));
 sg13g2_tielo tt_um_wokwi_group_4_28 (.L_LO(net28));
 sg13g2_tielo tt_um_wokwi_group_4_29 (.L_LO(net29));
 sg13g2_tielo tt_um_wokwi_group_4_30 (.L_LO(net30));
 sg13g2_tielo tt_um_wokwi_group_4_31 (.L_LO(net31));
 sg13g2_tielo tt_um_wokwi_group_4_32 (.L_LO(net32));
 sg13g2_tiehi \proj__1.flop1/_1__33  (.L_HI(net33));
 sg13g2_and2_1 \proj_10.and1/_0_  (.A(net124),
    .B(net129),
    .X(\proj_10.net11 ));
 sg13g2_and2_1 \proj_10.and2/_0_  (.A(net120),
    .B(\proj_10.net10 ),
    .X(\proj_10.net14 ));
 sg13g2_or2_1 \proj_10.or1/_0_  (.X(\proj_10.net5 ),
    .B(\proj_10.net14 ),
    .A(\proj_10.net11 ));
 sg13g2_xor2_1 \proj_10.xor1/_0_  (.B(net129),
    .A(net124),
    .X(\proj_10.net10 ));
 sg13g2_xor2_1 \proj_10.xor2/_0_  (.B(\proj_10.net10 ),
    .A(net120),
    .X(\proj_10.net4 ));
 sg13g2_and2_1 \proj_11.and1/_0_  (.A(net121),
    .B(net125),
    .X(\proj_11.net15 ));
 sg13g2_and2_1 \proj_11.and2/_0_  (.A(net1),
    .B(net117),
    .X(\proj_11.net17 ));
 sg13g2_and2_1 \proj_11.and3/_0_  (.A(\proj_11.net15 ),
    .B(\proj_11.net16 ),
    .X(\proj_11.net18 ));
 sg13g2_inv_1 \proj_11.not5/_0_  (.Y(\proj_11.net6 ),
    .A(net129));
 sg13g2_or2_1 \proj_11.or1/_0_  (.X(\proj_11.net9 ),
    .B(\proj_11.net18 ),
    .A(\proj_11.net17 ));
 sg13g2_xor2_1 \proj_11.xor1/_0_  (.B(net124),
    .A(net120),
    .X(\proj_11.net7 ));
 sg13g2_xor2_1 \proj_11.xor2/_0_  (.B(net116),
    .A(net115),
    .X(\proj_11.net16 ));
 sg13g2_xor2_1 \proj_11.xor3/_0_  (.B(\proj_11.net16 ),
    .A(\proj_11.net15 ),
    .X(\proj_11.net8 ));
 sg13g2_and2_1 \proj_12.and1/_0_  (.A(net122),
    .B(net127),
    .X(\proj_12.net4 ));
 sg13g2_xor2_1 \proj_12.xor1/_0_  (.B(net127),
    .A(net122),
    .X(\proj_12.net3 ));
 sg13g2_and2_1 \proj_13.and1/_0_  (.A(net122),
    .B(net127),
    .X(\proj_13.net8 ));
 sg13g2_and2_1 \proj_13.and2/_0_  (.A(net114),
    .B(net116),
    .X(\proj_13.net10 ));
 sg13g2_or2_1 \proj_13.or1/_0_  (.X(\proj_13.net9 ),
    .B(net121),
    .A(net122));
 sg13g2_xor2_1 \proj_13.xor1/_0_  (.B(net113),
    .A(net110),
    .X(\proj_13.net11 ));
 sg13g2_and2_1 \proj_14.and1/_0_  (.A(net120),
    .B(net129),
    .X(\proj_14.net15 ));
 sg13g2_and2_1 \proj_14.and2/_0_  (.A(net108),
    .B(\proj_14.net14 ),
    .X(\proj_14.net16 ));
 sg13g2_and2_1 \proj_14.and3/_0_  (.A(net117),
    .B(net123),
    .X(\proj_14.net19 ));
 sg13g2_and2_1 \proj_14.and4/_0_  (.A(\proj_14.net17 ),
    .B(\proj_14.net18 ),
    .X(\proj_14.net20 ));
 sg13g2_or2_1 \proj_14.or1/_0_  (.X(\proj_14.net17 ),
    .B(\proj_14.net16 ),
    .A(\proj_14.net15 ));
 sg13g2_or2_1 \proj_14.or2/_0_  (.X(\proj_14.net8 ),
    .B(\proj_14.net20 ),
    .A(\proj_14.net19 ));
 sg13g2_xor2_1 \proj_14.xor1/_0_  (.B(\proj_14.net14 ),
    .A(net108),
    .X(\proj_14.net6 ));
 sg13g2_xor2_1 \proj_14.xor2/_0_  (.B(net129),
    .A(net120),
    .X(\proj_14.net14 ));
 sg13g2_xor2_1 \proj_14.xor4/_0_  (.B(\proj_14.net18 ),
    .A(\proj_14.net17 ),
    .X(\proj_14.net7 ));
 sg13g2_xor2_1 \proj_14.xor5/_0_  (.B(net123),
    .A(net117),
    .X(\proj_14.net18 ));
 sg13g2_nand2_1 \proj_15.gate10/_0_  (.Y(\proj_15.net4 ),
    .A(\proj_15.net7 ),
    .B(\proj_15.net3 ));
 sg13g2_nand2_1 \proj_15.gate7/_0_  (.Y(\proj_15.net6 ),
    .A(net7),
    .B(net127));
 sg13g2_nand2_1 \proj_15.gate8/_0_  (.Y(\proj_15.net7 ),
    .A(net8),
    .B(\proj_15.net6 ));
 sg13g2_nand2_1 \proj_15.gate9/_0_  (.Y(\proj_15.net3 ),
    .A(\proj_15.net4 ),
    .B(\proj_15.net6 ));
 sg13g2_and2_1 \proj__0.and1/_0_  (.A(net122),
    .B(net127),
    .X(\proj__0.net11 ));
 sg13g2_and2_1 \proj__0.and2/_0_  (.A(net9),
    .B(net127),
    .X(\proj__0.net10 ));
 sg13g2_inv_1 \proj__0.not3/_0_  (.Y(\proj__0.net12 ),
    .A(net121));
 sg13g2_inv_1 \proj__0.not4/_0_  (.Y(\proj__0.net13 ),
    .A(net118));
 sg13g2_dfrbp_1 \proj__1.flop1/_1_  (.CLK(net10),
    .RESET_B(net33),
    .D(net122),
    .Q_N(\proj__1.flop1/notq ),
    .Q(\proj__1.net4 ));
 sg13g2_tiehi \proj__1.flop2/_1__34  (.L_HI(net34));
 sg13g2_dfrbp_1 \proj__1.flop2/_1_  (.CLK(net11),
    .RESET_B(net34),
    .D(\proj__1.net4 ),
    .Q_N(\proj__1.flop2/notq ),
    .Q(\proj__1.net5 ));
 sg13g2_tiehi \proj__1.flop3/_1__35  (.L_HI(net35));
 sg13g2_dfrbp_1 \proj__1.flop3/_1_  (.CLK(net12),
    .RESET_B(net35),
    .D(\proj__1.net5 ),
    .Q_N(\proj__1.flop3/notq ),
    .Q(\proj__1.net6 ));
 sg13g2_tiehi \proj__1.flop4/_1__36  (.L_HI(net36));
 sg13g2_dfrbp_1 \proj__1.flop4/_1_  (.CLK(net13),
    .RESET_B(net36),
    .D(\proj__1.net6 ),
    .Q_N(\proj__1.flop4/notq ),
    .Q(\proj__1.net7 ));
 sg13g2_tiehi \proj__1.flop5/_1__37  (.L_HI(net37));
 sg13g2_dfrbp_1 \proj__1.flop5/_1_  (.CLK(net14),
    .RESET_B(net37),
    .D(\proj__1.net7 ),
    .Q_N(\proj__1.flop5/notq ),
    .Q(\proj__1.net8 ));
 sg13g2_tiehi \proj__1.flop6/_1__38  (.L_HI(net38));
 sg13g2_dfrbp_1 \proj__1.flop6/_1_  (.CLK(net15),
    .RESET_B(net38),
    .D(\proj__1.net8 ),
    .Q_N(\proj__1.flop6/notq ),
    .Q(\proj__1.net9 ));
 sg13g2_tiehi \proj__4.flop1/_1__39  (.L_HI(net39));
 sg13g2_inv_1 \proj__2.not1/_0_  (.Y(\proj__2.net9 ),
    .A(net127));
 sg13g2_inv_1 \proj__2.not2/_0_  (.Y(\proj__2.net10 ),
    .A(net122));
 sg13g2_inv_1 \proj__2.not3/_0_  (.Y(\proj__2.net11 ),
    .A(net121));
 sg13g2_inv_1 \proj__2.not4/_0_  (.Y(\proj__2.net12 ),
    .A(net116));
 sg13g2_and2_1 \proj__3.and1/_0_  (.A(net109),
    .B(net110),
    .X(\proj__3.net13 ));
 sg13g2_nand2_1 \proj__3.nand1/_0_  (.Y(\proj__3.net12 ),
    .A(net109),
    .B(net110));
 sg13g2_inv_1 \proj__3.not1/_0_  (.Y(\proj__3.net9 ),
    .A(net128));
 sg13g2_inv_1 \proj__3.not2/_0_  (.Y(\proj__3.net14 ),
    .A(\proj__3.net10 ));
 sg13g2_or2_1 \proj__3.or1/_0_  (.X(\proj__3.net10 ),
    .B(net122),
    .A(net113));
 sg13g2_xor2_1 \proj__3.xor1/_0_  (.B(\proj__3.net20 ),
    .A(net114),
    .X(\proj__3.net11 ));
 sg13g2_xor2_1 \proj__3.xor2/_0_  (.B(net121),
    .A(net116),
    .X(\proj__3.net20 ));
 sg13g2_dfrbp_1 \proj__4.flop1/_1_  (.CLK(net116),
    .RESET_B(net39),
    .D(net121),
    .Q_N(\proj__4.net12 ),
    .Q(\proj__4.net11 ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_nand2_1 \proj__4.nand1/_0_  (.Y(\proj__4.net10 ),
    .A(net129),
    .B(net16));
 sg13g2_inv_1 \proj__4.not1/_0_  (.Y(\proj__4.net13 ),
    .A(net114));
 sg13g2_and2_1 \proj__5.and1/_0_  (.A(net125),
    .B(net128),
    .X(\proj__5.net9 ));
 sg13g2_or2_1 \proj__5.or1/_0_  (.X(\proj__5.net10 ),
    .B(net121),
    .A(net116));
 sg13g2_and2_1 \proj__6.and1/_0_  (.A(\proj__6.net23 ),
    .B(\proj__6.net22 ),
    .X(\proj__6.net25 ));
 sg13g2_and2_1 \proj__6.and10/_0_  (.A(net108),
    .B(\proj__6.net29 ),
    .X(\proj__6.net31 ));
 sg13g2_and2_1 \proj__6.and11/_0_  (.A(net110),
    .B(\proj__6.net28 ),
    .X(\proj__6.net34 ));
 sg13g2_and2_1 \proj__6.and12/_0_  (.A(\proj__6.net31 ),
    .B(\proj__6.net28 ),
    .X(\proj__6.net35 ));
 sg13g2_and2_1 \proj__6.and13/_0_  (.A(\proj__6.net31 ),
    .B(net110),
    .X(\proj__6.net36 ));
 sg13g2_and2_1 \proj__6.and14/_0_  (.A(net112),
    .B(\proj__6.net24 ),
    .X(\proj__6.net41 ));
 sg13g2_and2_1 \proj__6.and15/_0_  (.A(\proj__6.net38 ),
    .B(\proj__6.net24 ),
    .X(\proj__6.net42 ));
 sg13g2_and2_1 \proj__6.and16/_0_  (.A(\proj__6.net38 ),
    .B(net112),
    .X(\proj__6.net43 ));
 sg13g2_and2_1 \proj__6.and17/_0_  (.A(net1),
    .B(\proj__6.net25 ),
    .X(\proj__6.net48 ));
 sg13g2_and2_1 \proj__6.and18/_0_  (.A(\proj__6.net45 ),
    .B(\proj__6.net25 ),
    .X(\proj__6.net49 ));
 sg13g2_and2_1 \proj__6.and19/_0_  (.A(\proj__6.net45 ),
    .B(net115),
    .X(\proj__6.net50 ));
 sg13g2_and2_1 \proj__6.and2/_0_  (.A(\proj__6.net27 ),
    .B(\proj__6.net26 ),
    .X(\proj__6.net22 ));
 sg13g2_and2_1 \proj__6.and20/_0_  (.A(\proj__6.net53 ),
    .B(\proj__6.net52 ),
    .X(\proj__6.net54 ));
 sg13g2_and2_1 \proj__6.and21/_0_  (.A(\proj__6.net56 ),
    .B(\proj__6.net55 ),
    .X(\proj__6.net57 ));
 sg13g2_and2_1 \proj__6.and22/_0_  (.A(\proj__6.net57 ),
    .B(\proj__6.net54 ),
    .X(\proj__6.net58 ));
 sg13g2_and2_1 \proj__6.and23/_0_  (.A(\proj__6.net59 ),
    .B(net106),
    .X(\proj__6.net60 ));
 sg13g2_and2_1 \proj__6.and24/_0_  (.A(\proj__6.net62 ),
    .B(\proj__6.net61 ),
    .X(\proj__6.net63 ));
 sg13g2_and2_1 \proj__6.and25/_0_  (.A(\proj__6.net63 ),
    .B(\proj__6.net60 ),
    .X(\proj__6.net64 ));
 sg13g2_and2_1 \proj__6.and26/_0_  (.A(net104),
    .B(net106),
    .X(\proj__6.net71 ));
 sg13g2_and2_1 \proj__6.and27/_0_  (.A(\proj__6.net73 ),
    .B(\proj__6.net72 ),
    .X(\proj__6.net74 ));
 sg13g2_and2_1 \proj__6.and28/_0_  (.A(\proj__6.net74 ),
    .B(\proj__6.net71 ),
    .X(\proj__6.net75 ));
 sg13g2_and2_1 \proj__6.and29/_0_  (.A(\proj__6.net77 ),
    .B(\proj__6.net76 ),
    .X(\proj__6.net78 ));
 sg13g2_and2_1 \proj__6.and3/_0_  (.A(net117),
    .B(net130),
    .X(\proj__6.net26 ));
 sg13g2_and2_1 \proj__6.and30/_0_  (.A(\proj__6.net79 ),
    .B(\proj__6.net40 ),
    .X(\proj__6.net80 ));
 sg13g2_and2_1 \proj__6.and31/_0_  (.A(\proj__6.net80 ),
    .B(\proj__6.net78 ),
    .X(\proj__6.net81 ));
 sg13g2_and2_1 \proj__6.and32/_0_  (.A(\proj__6.net82 ),
    .B(\proj__6.net30 ),
    .X(\proj__6.net83 ));
 sg13g2_and2_1 \proj__6.and33/_0_  (.A(\proj__6.net84 ),
    .B(net102),
    .X(\proj__6.net85 ));
 sg13g2_and2_1 \proj__6.and34/_0_  (.A(\proj__6.net85 ),
    .B(\proj__6.net83 ),
    .X(\proj__6.net86 ));
 sg13g2_and2_1 \proj__6.and35/_0_  (.A(net104),
    .B(\proj__6.net87 ),
    .X(\proj__6.net88 ));
 sg13g2_and2_1 \proj__6.and36/_0_  (.A(\proj__6.net89 ),
    .B(net102),
    .X(\proj__6.net90 ));
 sg13g2_and2_1 \proj__6.and37/_0_  (.A(\proj__6.net90 ),
    .B(\proj__6.net88 ),
    .X(\proj__6.net91 ));
 sg13g2_and2_1 \proj__6.and38/_0_  (.A(net104),
    .B(net106),
    .X(\proj__6.net92 ));
 sg13g2_and2_1 \proj__6.and39/_0_  (.A(\proj__6.net93 ),
    .B(net102),
    .X(\proj__6.net94 ));
 sg13g2_and2_1 \proj__6.and4/_0_  (.A(net117),
    .B(net125),
    .X(\proj__6.net29 ));
 sg13g2_and2_1 \proj__6.and40/_0_  (.A(\proj__6.net94 ),
    .B(\proj__6.net92 ),
    .X(\proj__6.net95 ));
 sg13g2_and2_1 \proj__6.and41/_0_  (.A(\proj__6.net97 ),
    .B(\proj__6.net96 ),
    .X(\proj__6.net98 ));
 sg13g2_and2_1 \proj__6.and42/_0_  (.A(net99),
    .B(\proj__6.net99 ),
    .X(\proj__6.net100 ));
 sg13g2_and2_2 \proj__6.and43/_0_  (.A(\proj__6.net100 ),
    .B(\proj__6.net98 ),
    .X(\proj__6.net101 ));
 sg13g2_and2_1 \proj__6.and44/_0_  (.A(\proj__6.net102 ),
    .B(net105),
    .X(\proj__6.net103 ));
 sg13g2_and2_1 \proj__6.and45/_0_  (.A(net99),
    .B(\proj__6.net104 ),
    .X(\proj__6.net105 ));
 sg13g2_and2_1 \proj__6.and46/_0_  (.A(\proj__6.net105 ),
    .B(\proj__6.net103 ),
    .X(\proj__6.net106 ));
 sg13g2_and2_1 \proj__6.and47/_0_  (.A(net104),
    .B(\proj__6.net65 ),
    .X(\proj__6.net66 ));
 sg13g2_and2_1 \proj__6.and48/_0_  (.A(\proj__6.net68 ),
    .B(\proj__6.net67 ),
    .X(\proj__6.net69 ));
 sg13g2_and2_1 \proj__6.and49/_0_  (.A(\proj__6.net69 ),
    .B(\proj__6.net66 ),
    .X(\proj__6.net70 ));
 sg13g2_and2_1 \proj__6.and5/_0_  (.A(net119),
    .B(net129),
    .X(\proj__6.net23 ));
 sg13g2_and2_1 \proj__6.and50/_0_  (.A(net103),
    .B(\proj__6.net107 ),
    .X(\proj__6.net108 ));
 sg13g2_and2_1 \proj__6.and51/_0_  (.A(net99),
    .B(\proj__6.net109 ),
    .X(\proj__6.net110 ));
 sg13g2_and2_1 \proj__6.and52/_0_  (.A(\proj__6.net110 ),
    .B(\proj__6.net108 ),
    .X(\proj__6.net111 ));
 sg13g2_and2_1 \proj__6.and53/_0_  (.A(net103),
    .B(net105),
    .X(\proj__6.net112 ));
 sg13g2_and2_1 \proj__6.and54/_0_  (.A(net99),
    .B(\proj__6.net113 ),
    .X(\proj__6.net114 ));
 sg13g2_and2_1 \proj__6.and55/_0_  (.A(\proj__6.net114 ),
    .B(\proj__6.net112 ),
    .X(\proj__6.net115 ));
 sg13g2_and2_1 \proj__6.and56/_0_  (.A(\proj__6.net117 ),
    .B(\proj__6.net116 ),
    .X(\proj__6.net118 ));
 sg13g2_and2_1 \proj__6.and57/_0_  (.A(net99),
    .B(net101),
    .X(\proj__6.net119 ));
 sg13g2_and2_1 \proj__6.and58/_0_  (.A(\proj__6.net119 ),
    .B(\proj__6.net118 ),
    .X(\proj__6.net120 ));
 sg13g2_and2_1 \proj__6.and59/_0_  (.A(\proj__6.net121 ),
    .B(net105),
    .X(\proj__6.net122 ));
 sg13g2_and2_1 \proj__6.and6/_0_  (.A(net119),
    .B(net123),
    .X(\proj__6.net27 ));
 sg13g2_and2_1 \proj__6.and60/_0_  (.A(net99),
    .B(net101),
    .X(\proj__6.net123 ));
 sg13g2_and2_1 \proj__6.and61/_0_  (.A(\proj__6.net123 ),
    .B(\proj__6.net122 ),
    .X(\proj__6.net124 ));
 sg13g2_and2_1 \proj__6.and62/_0_  (.A(net103),
    .B(\proj__6.net125 ),
    .X(\proj__6.net126 ));
 sg13g2_and2_1 \proj__6.and63/_0_  (.A(net99),
    .B(net101),
    .X(\proj__6.net127 ));
 sg13g2_and2_1 \proj__6.and64/_0_  (.A(\proj__6.net127 ),
    .B(\proj__6.net126 ),
    .X(\proj__6.net128 ));
 sg13g2_and2_1 \proj__6.and65/_0_  (.A(net103),
    .B(net105),
    .X(\proj__6.net129 ));
 sg13g2_and2_1 \proj__6.and66/_0_  (.A(net99),
    .B(net101),
    .X(\proj__6.net130 ));
 sg13g2_and2_1 \proj__6.and67/_0_  (.A(\proj__6.net130 ),
    .B(\proj__6.net129 ),
    .X(\proj__6.net131 ));
 sg13g2_inv_1 \proj__6.not10/_0_  (.Y(\proj__6.net62 ),
    .A(\proj__6.net47 ));
 sg13g2_inv_1 \proj__6.not11/_0_  (.Y(\proj__6.net61 ),
    .A(net102));
 sg13g2_inv_1 \proj__6.not12/_0_  (.Y(\proj__6.net59 ),
    .A(net104));
 sg13g2_inv_1 \proj__6.not14/_0_  (.Y(\proj__6.net73 ),
    .A(net100));
 sg13g2_inv_1 \proj__6.not15/_0_  (.Y(\proj__6.net72 ),
    .A(net102));
 sg13g2_inv_1 \proj__6.not17/_0_  (.Y(\proj__6.net76 ),
    .A(net106));
 sg13g2_inv_1 \proj__6.not18/_0_  (.Y(\proj__6.net79 ),
    .A(net100));
 sg13g2_inv_1 \proj__6.not20/_0_  (.Y(\proj__6.net77 ),
    .A(net104));
 sg13g2_inv_1 \proj__6.not22/_0_  (.Y(\proj__6.net84 ),
    .A(net100));
 sg13g2_inv_1 \proj__6.not24/_0_  (.Y(\proj__6.net82 ),
    .A(\proj__6.net33 ));
 sg13g2_inv_1 \proj__6.not25/_0_  (.Y(\proj__6.net87 ),
    .A(net106));
 sg13g2_inv_1 \proj__6.not26/_0_  (.Y(\proj__6.net89 ),
    .A(net100));
 sg13g2_inv_1 \proj__6.not30/_0_  (.Y(\proj__6.net93 ),
    .A(net100));
 sg13g2_inv_1 \proj__6.not33/_0_  (.Y(\proj__6.net96 ),
    .A(net105));
 sg13g2_inv_1 \proj__6.not35/_0_  (.Y(\proj__6.net99 ),
    .A(net101));
 sg13g2_inv_1 \proj__6.not36/_0_  (.Y(\proj__6.net97 ),
    .A(net103));
 sg13g2_inv_1 \proj__6.not39/_0_  (.Y(\proj__6.net104 ),
    .A(net101));
 sg13g2_inv_1 \proj__6.not40/_0_  (.Y(\proj__6.net102 ),
    .A(net103));
 sg13g2_inv_1 \proj__6.not41/_0_  (.Y(\proj__6.net65 ),
    .A(net106));
 sg13g2_inv_1 \proj__6.not42/_0_  (.Y(\proj__6.net68 ),
    .A(net100));
 sg13g2_inv_1 \proj__6.not43/_0_  (.Y(\proj__6.net67 ),
    .A(net102));
 sg13g2_inv_1 \proj__6.not45/_0_  (.Y(\proj__6.net107 ),
    .A(net105));
 sg13g2_inv_1 \proj__6.not47/_0_  (.Y(\proj__6.net109 ),
    .A(net101));
 sg13g2_inv_1 \proj__6.not5/_0_  (.Y(\proj__6.net52 ),
    .A(net106));
 sg13g2_inv_1 \proj__6.not51/_0_  (.Y(\proj__6.net113 ),
    .A(net101));
 sg13g2_inv_1 \proj__6.not53/_0_  (.Y(\proj__6.net116 ),
    .A(net105));
 sg13g2_inv_1 \proj__6.not56/_0_  (.Y(\proj__6.net117 ),
    .A(net103));
 sg13g2_inv_1 \proj__6.not6/_0_  (.Y(\proj__6.net56 ),
    .A(net100));
 sg13g2_inv_1 \proj__6.not60/_0_  (.Y(\proj__6.net121 ),
    .A(net103));
 sg13g2_inv_1 \proj__6.not61/_0_  (.Y(\proj__6.net125 ),
    .A(net105));
 sg13g2_inv_1 \proj__6.not7/_0_  (.Y(\proj__6.net55 ),
    .A(net102));
 sg13g2_inv_1 \proj__6.not8/_0_  (.Y(\proj__6.net53 ),
    .A(net104));
 sg13g2_or2_1 \proj__6.or1/_0_  (.X(\proj__6.net132 ),
    .B(\proj__6.net58 ),
    .A(\proj__6.net70 ));
 sg13g2_or2_1 \proj__6.or10/_0_  (.X(\proj__6.net135 ),
    .B(\proj__6.net101 ),
    .A(\proj__6.net106 ));
 sg13g2_or2_1 \proj__6.or11/_0_  (.X(\proj__6.net136 ),
    .B(\proj__6.net111 ),
    .A(\proj__6.net120 ));
 sg13g2_or2_1 \proj__6.or12/_0_  (.X(\proj__6.net137 ),
    .B(\proj__6.net128 ),
    .A(\proj__6.net131 ));
 sg13g2_or2_1 \proj__6.or13/_0_  (.X(\proj__6.net138 ),
    .B(\proj__6.net132 ),
    .A(\proj__6.net133 ));
 sg13g2_or2_1 \proj__6.or14/_0_  (.X(\proj__6.net139 ),
    .B(\proj__6.net134 ),
    .A(\proj__6.net135 ));
 sg13g2_or2_1 \proj__6.or15/_0_  (.X(\proj__6.net140 ),
    .B(\proj__6.net136 ),
    .A(\proj__6.net137 ));
 sg13g2_or2_1 \proj__6.or16/_0_  (.X(\proj__6.net142 ),
    .B(\proj__6.net58 ),
    .A(\proj__6.net64 ));
 sg13g2_or2_1 \proj__6.or17/_0_  (.X(\proj__6.net143 ),
    .B(\proj__6.net70 ),
    .A(\proj__6.net75 ));
 sg13g2_or2_1 \proj__6.or18/_0_  (.X(\proj__6.net144 ),
    .B(\proj__6.net81 ),
    .A(\proj__6.net95 ));
 sg13g2_or2_1 \proj__6.or19/_0_  (.X(\proj__6.net141 ),
    .B(\proj__6.net138 ),
    .A(\proj__6.net139 ));
 sg13g2_or2_1 \proj__6.or2/_0_  (.X(\proj__6.net133 ),
    .B(\proj__6.net75 ),
    .A(\proj__6.net86 ));
 sg13g2_or2_1 \proj__6.or20/_0_  (.X(\proj__6.net145 ),
    .B(\proj__6.net101 ),
    .A(\proj__6.net106 ));
 sg13g2_or2_1 \proj__6.or21/_0_  (.X(\proj__6.net9 ),
    .B(\proj__6.net141 ),
    .A(\proj__6.net140 ));
 sg13g2_or2_1 \proj__6.or3/_0_  (.X(\proj__6.net37 ),
    .B(\proj__6.net34 ),
    .A(\proj__6.net36 ));
 sg13g2_or2_1 \proj__6.or37/_0_  (.X(\proj__6.net146 ),
    .B(\proj__6.net120 ),
    .A(\proj__6.net124 ));
 sg13g2_or2_1 \proj__6.or38/_0_  (.X(\proj__6.net150 ),
    .B(\proj__6.net58 ),
    .A(\proj__6.net64 ));
 sg13g2_or2_1 \proj__6.or39/_0_  (.X(\proj__6.net147 ),
    .B(\proj__6.net142 ),
    .A(\proj__6.net143 ));
 sg13g2_or2_1 \proj__6.or4/_0_  (.X(\proj__6.net38 ),
    .B(\proj__6.net37 ),
    .A(\proj__6.net35 ));
 sg13g2_or2_1 \proj__6.or40/_0_  (.X(\proj__6.net148 ),
    .B(\proj__6.net144 ),
    .A(\proj__6.net145 ));
 sg13g2_or2_1 \proj__6.or41/_0_  (.X(\proj__6.net151 ),
    .B(\proj__6.net75 ),
    .A(\proj__6.net81 ));
 sg13g2_or2_1 \proj__6.or42/_0_  (.X(\proj__6.net152 ),
    .B(\proj__6.net86 ),
    .A(\proj__6.net91 ));
 sg13g2_or2_1 \proj__6.or43/_0_  (.X(\proj__6.net153 ),
    .B(\proj__6.net95 ),
    .A(\proj__6.net101 ));
 sg13g2_or2_1 \proj__6.or44/_0_  (.X(\proj__6.net154 ),
    .B(\proj__6.net106 ),
    .A(\proj__6.net111 ));
 sg13g2_or2_1 \proj__6.or45/_0_  (.X(\proj__6.net149 ),
    .B(\proj__6.net147 ),
    .A(\proj__6.net148 ));
 sg13g2_or2_1 \proj__6.or46/_0_  (.X(\proj__6.net155 ),
    .B(\proj__6.net115 ),
    .A(\proj__6.net124 ));
 sg13g2_or2_1 \proj__6.or47/_0_  (.X(\proj__6.net10 ),
    .B(\proj__6.net149 ),
    .A(\proj__6.net146 ));
 sg13g2_or2_1 \proj__6.or48/_0_  (.X(\proj__6.net156 ),
    .B(\proj__6.net150 ),
    .A(\proj__6.net151 ));
 sg13g2_or2_1 \proj__6.or49/_0_  (.X(\proj__6.net157 ),
    .B(\proj__6.net152 ),
    .A(\proj__6.net153 ));
 sg13g2_or2_1 \proj__6.or5/_0_  (.X(\proj__6.net44 ),
    .B(\proj__6.net41 ),
    .A(\proj__6.net43 ));
 sg13g2_or2_1 \proj__6.or50/_0_  (.X(\proj__6.net158 ),
    .B(\proj__6.net154 ),
    .A(\proj__6.net155 ));
 sg13g2_or2_1 \proj__6.or51/_0_  (.X(\proj__6.net159 ),
    .B(\proj__6.net156 ),
    .A(\proj__6.net157 ));
 sg13g2_or2_1 \proj__6.or52/_0_  (.X(\proj__6.net11 ),
    .B(\proj__6.net159 ),
    .A(\proj__6.net158 ));
 sg13g2_or2_1 \proj__6.or53/_0_  (.X(\proj__6.net160 ),
    .B(\proj__6.net58 ),
    .A(\proj__6.net70 ));
 sg13g2_or2_1 \proj__6.or54/_0_  (.X(\proj__6.net161 ),
    .B(\proj__6.net75 ),
    .A(\proj__6.net86 ));
 sg13g2_or2_1 \proj__6.or55/_0_  (.X(\proj__6.net162 ),
    .B(\proj__6.net91 ),
    .A(\proj__6.net101 ));
 sg13g2_or2_1 \proj__6.or56/_0_  (.X(\proj__6.net163 ),
    .B(\proj__6.net106 ),
    .A(\proj__6.net115 ));
 sg13g2_or2_1 \proj__6.or57/_0_  (.X(\proj__6.net164 ),
    .B(\proj__6.net120 ),
    .A(\proj__6.net124 ));
 sg13g2_or2_1 \proj__6.or58/_0_  (.X(\proj__6.net169 ),
    .B(\proj__6.net58 ),
    .A(\proj__6.net70 ));
 sg13g2_or2_1 \proj__6.or59/_0_  (.X(\proj__6.net165 ),
    .B(\proj__6.net160 ),
    .A(\proj__6.net161 ));
 sg13g2_or2_1 \proj__6.or6/_0_  (.X(\proj__6.net45 ),
    .B(\proj__6.net44 ),
    .A(\proj__6.net42 ));
 sg13g2_or2_1 \proj__6.or60/_0_  (.X(\proj__6.net166 ),
    .B(\proj__6.net162 ),
    .A(\proj__6.net163 ));
 sg13g2_or2_1 \proj__6.or61/_0_  (.X(\proj__6.net167 ),
    .B(\proj__6.net164 ),
    .A(\proj__6.net128 ));
 sg13g2_or2_1 \proj__6.or62/_0_  (.X(\proj__6.net168 ),
    .B(\proj__6.net165 ),
    .A(\proj__6.net166 ));
 sg13g2_or2_1 \proj__6.or63/_0_  (.X(\proj__6.net12 ),
    .B(\proj__6.net168 ),
    .A(\proj__6.net167 ));
 sg13g2_or2_1 \proj__6.or64/_0_  (.X(\proj__6.net170 ),
    .B(\proj__6.net91 ),
    .A(\proj__6.net101 ));
 sg13g2_or2_1 \proj__6.or65/_0_  (.X(\proj__6.net171 ),
    .B(\proj__6.net111 ),
    .A(\proj__6.net115 ));
 sg13g2_or2_1 \proj__6.or66/_0_  (.X(\proj__6.net172 ),
    .B(\proj__6.net120 ),
    .A(\proj__6.net124 ));
 sg13g2_or2_1 \proj__6.or67/_0_  (.X(\proj__6.net173 ),
    .B(\proj__6.net128 ),
    .A(\proj__6.net131 ));
 sg13g2_or2_1 \proj__6.or68/_0_  (.X(\proj__6.net174 ),
    .B(\proj__6.net169 ),
    .A(\proj__6.net170 ));
 sg13g2_or2_1 \proj__6.or69/_0_  (.X(\proj__6.net175 ),
    .B(\proj__6.net171 ),
    .A(\proj__6.net172 ));
 sg13g2_or2_1 \proj__6.or7/_0_  (.X(\proj__6.net51 ),
    .B(\proj__6.net48 ),
    .A(\proj__6.net50 ));
 sg13g2_or2_1 \proj__6.or70/_0_  (.X(\proj__6.net176 ),
    .B(\proj__6.net174 ),
    .A(\proj__6.net175 ));
 sg13g2_or2_1 \proj__6.or71/_0_  (.X(\proj__6.net13 ),
    .B(\proj__6.net176 ),
    .A(\proj__6.net173 ));
 sg13g2_or2_1 \proj__6.or72/_0_  (.X(\proj__6.net177 ),
    .B(\proj__6.net58 ),
    .A(\proj__6.net81 ));
 sg13g2_or2_1 \proj__6.or73/_0_  (.X(\proj__6.net178 ),
    .B(\proj__6.net86 ),
    .A(\proj__6.net91 ));
 sg13g2_or2_1 \proj__6.or74/_0_  (.X(\proj__6.net179 ),
    .B(\proj__6.net101 ),
    .A(\proj__6.net106 ));
 sg13g2_or2_1 \proj__6.or75/_0_  (.X(\proj__6.net180 ),
    .B(\proj__6.net111 ),
    .A(\proj__6.net115 ));
 sg13g2_or2_1 \proj__6.or76/_0_  (.X(\proj__6.net181 ),
    .B(\proj__6.net120 ),
    .A(\proj__6.net128 ));
 sg13g2_or2_1 \proj__6.or77/_0_  (.X(\proj__6.net182 ),
    .B(\proj__6.net177 ),
    .A(\proj__6.net178 ));
 sg13g2_or2_1 \proj__6.or78/_0_  (.X(\proj__6.net183 ),
    .B(\proj__6.net179 ),
    .A(\proj__6.net180 ));
 sg13g2_or2_1 \proj__6.or79/_0_  (.X(\proj__6.net184 ),
    .B(\proj__6.net181 ),
    .A(\proj__6.net131 ));
 sg13g2_or2_1 \proj__6.or8/_0_  (.X(\proj__6.net16 ),
    .B(\proj__6.net51 ),
    .A(\proj__6.net49 ));
 sg13g2_or2_1 \proj__6.or80/_0_  (.X(\proj__6.net185 ),
    .B(\proj__6.net182 ),
    .A(\proj__6.net183 ));
 sg13g2_or2_1 \proj__6.or81/_0_  (.X(\proj__6.net14 ),
    .B(\proj__6.net185 ),
    .A(\proj__6.net184 ));
 sg13g2_or2_1 \proj__6.or82/_0_  (.X(\proj__6.net186 ),
    .B(\proj__6.net70 ),
    .A(\proj__6.net75 ));
 sg13g2_or2_1 \proj__6.or83/_0_  (.X(\proj__6.net187 ),
    .B(\proj__6.net81 ),
    .A(\proj__6.net86 ));
 sg13g2_or2_1 \proj__6.or84/_0_  (.X(\proj__6.net188 ),
    .B(\proj__6.net91 ),
    .A(\proj__6.net101 ));
 sg13g2_or2_1 \proj__6.or85/_0_  (.X(\proj__6.net189 ),
    .B(\proj__6.net106 ),
    .A(\proj__6.net111 ));
 sg13g2_or2_1 \proj__6.or86/_0_  (.X(\proj__6.net190 ),
    .B(\proj__6.net115 ),
    .A(\proj__6.net124 ));
 sg13g2_or2_1 \proj__6.or87/_0_  (.X(\proj__6.net191 ),
    .B(\proj__6.net128 ),
    .A(\proj__6.net131 ));
 sg13g2_or2_1 \proj__6.or88/_0_  (.X(\proj__6.net192 ),
    .B(\proj__6.net186 ),
    .A(\proj__6.net187 ));
 sg13g2_or2_1 \proj__6.or89/_0_  (.X(\proj__6.net193 ),
    .B(\proj__6.net188 ),
    .A(\proj__6.net189 ));
 sg13g2_or2_1 \proj__6.or9/_0_  (.X(\proj__6.net134 ),
    .B(\proj__6.net91 ),
    .A(\proj__6.net95 ));
 sg13g2_or2_1 \proj__6.or90/_0_  (.X(\proj__6.net194 ),
    .B(\proj__6.net190 ),
    .A(\proj__6.net191 ));
 sg13g2_or2_1 \proj__6.or91/_0_  (.X(\proj__6.net195 ),
    .B(\proj__6.net192 ),
    .A(\proj__6.net193 ));
 sg13g2_or2_1 \proj__6.or92/_0_  (.X(\proj__6.net15 ),
    .B(\proj__6.net195 ),
    .A(\proj__6.net194 ));
 sg13g2_xor2_1 \proj__6.xor1/_0_  (.B(\proj__6.net22 ),
    .A(\proj__6.net23 ),
    .X(\proj__6.net24 ));
 sg13g2_xor2_1 \proj__6.xor10/_0_  (.B(\proj__6.net25 ),
    .A(net114),
    .X(\proj__6.net46 ));
 sg13g2_xor2_1 \proj__6.xor11/_0_  (.B(\proj__6.net46 ),
    .A(\proj__6.net45 ),
    .X(\proj__6.net47 ));
 sg13g2_xor2_1 \proj__6.xor2/_0_  (.B(\proj__6.net26 ),
    .A(\proj__6.net27 ),
    .X(\proj__6.net28 ));
 sg13g2_xor2_1 \proj__6.xor5/_0_  (.B(\proj__6.net29 ),
    .A(net108),
    .X(\proj__6.net30 ));
 sg13g2_xor2_1 \proj__6.xor6/_0_  (.B(\proj__6.net28 ),
    .A(net110),
    .X(\proj__6.net32 ));
 sg13g2_xor2_1 \proj__6.xor7/_0_  (.B(\proj__6.net32 ),
    .A(\proj__6.net31 ),
    .X(\proj__6.net33 ));
 sg13g2_xor2_1 \proj__6.xor8/_0_  (.B(\proj__6.net24 ),
    .A(net112),
    .X(\proj__6.net39 ));
 sg13g2_xor2_1 \proj__6.xor9/_0_  (.B(\proj__6.net39 ),
    .A(\proj__6.net38 ),
    .X(\proj__6.net40 ));
 sg13g2_and2_1 \proj__7.and1/_0_  (.A(net126),
    .B(net127),
    .X(\proj__7.net7 ));
 sg13g2_or2_1 \proj__8.gate1/_0_  (.X(\proj__8.net18 ),
    .B(net124),
    .A(net119));
 sg13g2_or2_1 \proj__8.gate10/_0_  (.X(\proj__8.net22 ),
    .B(net130),
    .A(net123));
 sg13g2_or2_1 \proj__8.gate11/_0_  (.X(\proj__8.net27 ),
    .B(\proj__8.net26 ),
    .A(net117));
 sg13g2_or2_1 \proj__8.gate12/_0_  (.X(\proj__8.net28 ),
    .B(\proj__8.net27 ),
    .A(net115));
 sg13g2_or2_1 \proj__8.gate13/_0_  (.X(\proj__8.net30 ),
    .B(\proj__8.net29 ),
    .A(net111));
 sg13g2_or2_1 \proj__8.gate14/_0_  (.X(\proj__8.net29 ),
    .B(\proj__8.net28 ),
    .A(net112));
 sg13g2_or2_1 \proj__8.gate15/_0_  (.X(\proj__8.net26 ),
    .B(net130),
    .A(net119));
 sg13g2_or2_1 \proj__8.gate16/_0_  (.X(\proj__8.net11 ),
    .B(\proj__8.net30 ),
    .A(net108));
 sg13g2_or2_1 \proj__8.gate17/_0_  (.X(\proj__8.net32 ),
    .B(\proj__8.net31 ),
    .A(net115));
 sg13g2_or2_1 \proj__8.gate18/_0_  (.X(\proj__8.net33 ),
    .B(\proj__8.net32 ),
    .A(net112));
 sg13g2_or2_1 \proj__8.gate19/_0_  (.X(\proj__8.net12 ),
    .B(\proj__8.net33 ),
    .A(net108));
 sg13g2_or2_1 \proj__8.gate2/_0_  (.X(\proj__8.net19 ),
    .B(\proj__8.net18 ),
    .A(net115));
 sg13g2_or2_1 \proj__8.gate20/_0_  (.X(\proj__8.net31 ),
    .B(net123),
    .A(net119));
 sg13g2_or2_1 \proj__8.gate21/_0_  (.X(\proj__8.net13 ),
    .B(\proj__8.net34 ),
    .A(net2));
 sg13g2_or2_1 \proj__8.gate22/_0_  (.X(\proj__8.net34 ),
    .B(net123),
    .A(net113));
 sg13g2_or2_1 \proj__8.gate23/_0_  (.X(\proj__8.net36 ),
    .B(\proj__8.net35 ),
    .A(net113));
 sg13g2_or2_1 \proj__8.gate24/_0_  (.X(\proj__8.net14 ),
    .B(\proj__8.net36 ),
    .A(net109));
 sg13g2_or2_1 \proj__8.gate25/_0_  (.X(\proj__8.net35 ),
    .B(net116),
    .A(net114));
 sg13g2_or2_1 \proj__8.gate26/_0_  (.X(\proj__8.net38 ),
    .B(\proj__8.net37 ),
    .A(net116));
 sg13g2_or2_1 \proj__8.gate27/_0_  (.X(\proj__8.net39 ),
    .B(\proj__8.net38 ),
    .A(net114));
 sg13g2_or2_1 \proj__8.gate28/_0_  (.X(\proj__8.net15 ),
    .B(\proj__8.net40 ),
    .A(net109));
 sg13g2_or2_1 \proj__8.gate29/_0_  (.X(\proj__8.net40 ),
    .B(\proj__8.net39 ),
    .A(net113));
 sg13g2_or2_1 \proj__8.gate3/_0_  (.X(\proj__8.net21 ),
    .B(\proj__8.net20 ),
    .A(net111));
 sg13g2_or2_1 \proj__8.gate30/_0_  (.X(\proj__8.net37 ),
    .B(net126),
    .A(net121));
 sg13g2_or2_1 \proj__8.gate4/_0_  (.X(\proj__8.net20 ),
    .B(\proj__8.net19 ),
    .A(net112));
 sg13g2_or2_1 \proj__8.gate5/_0_  (.X(\proj__8.net9 ),
    .B(\proj__8.net21 ),
    .A(net109));
 sg13g2_or2_1 \proj__8.gate6/_0_  (.X(\proj__8.net23 ),
    .B(\proj__8.net22 ),
    .A(net119));
 sg13g2_or2_1 \proj__8.gate7/_0_  (.X(\proj__8.net24 ),
    .B(\proj__8.net23 ),
    .A(net118));
 sg13g2_or2_1 \proj__8.gate8/_0_  (.X(\proj__8.net10 ),
    .B(\proj__8.net25 ),
    .A(net109));
 sg13g2_or2_1 \proj__8.gate9/_0_  (.X(\proj__8.net25 ),
    .B(\proj__8.net24 ),
    .A(net111));
 sg13g2_and2_1 \proj__9.and1/_0_  (.A(net112),
    .B(net123),
    .X(\proj__9.net20 ));
 sg13g2_and2_1 \proj__9.and2/_0_  (.A(\proj__9.net19 ),
    .B(\proj__9.net21 ),
    .X(\proj__9.net22 ));
 sg13g2_and2_1 \proj__9.and3/_0_  (.A(net111),
    .B(net119),
    .X(\proj__9.net25 ));
 sg13g2_and2_1 \proj__9.and4/_0_  (.A(\proj__9.net24 ),
    .B(\proj__9.net23 ),
    .X(\proj__9.net26 ));
 sg13g2_and2_1 \proj__9.and5/_0_  (.A(net108),
    .B(net117),
    .X(\proj__9.net29 ));
 sg13g2_and2_1 \proj__9.and6/_0_  (.A(\proj__9.net28 ),
    .B(\proj__9.net27 ),
    .X(\proj__9.net30 ));
 sg13g2_and2_1 \proj__9.and7/_0_  (.A(net115),
    .B(net129),
    .X(\proj__9.net21 ));
 sg13g2_or2_1 \proj__9.or1/_0_  (.X(\proj__9.net23 ),
    .B(\proj__9.net22 ),
    .A(\proj__9.net20 ));
 sg13g2_or2_1 \proj__9.or2/_0_  (.X(\proj__9.net27 ),
    .B(\proj__9.net26 ),
    .A(\proj__9.net25 ));
 sg13g2_or2_1 \proj__9.or3/_0_  (.X(\proj__9.net13 ),
    .B(\proj__9.net30 ),
    .A(\proj__9.net29 ));
 sg13g2_xor2_1 \proj__9.xor1/_0_  (.B(net123),
    .A(net112),
    .X(\proj__9.net19 ));
 sg13g2_xor2_1 \proj__9.xor2/_0_  (.B(\proj__9.net21 ),
    .A(\proj__9.net19 ),
    .X(\proj__9.net10 ));
 sg13g2_xor2_1 \proj__9.xor3/_0_  (.B(net119),
    .A(net110),
    .X(\proj__9.net24 ));
 sg13g2_xor2_1 \proj__9.xor4/_0_  (.B(\proj__9.net23 ),
    .A(\proj__9.net24 ),
    .X(\proj__9.net11 ));
 sg13g2_xor2_1 \proj__9.xor5/_0_  (.B(net117),
    .A(net108),
    .X(\proj__9.net28 ));
 sg13g2_xor2_1 \proj__9.xor6/_0_  (.B(\proj__9.net27 ),
    .A(\proj__9.net28 ),
    .X(\proj__9.net12 ));
 sg13g2_xor2_1 \proj__9.xor7/_0_  (.B(net128),
    .A(net114),
    .X(\proj__9.net9 ));
 sg13g2_buf_2 fanout99 (.A(net100),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(\proj__6.net47 ),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(net102),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(\proj__6.net40 ),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(net104),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(\proj__6.net33 ),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(net106),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(\proj__6.net30 ),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(net4),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(net109),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(net2),
    .X(net109));
 sg13g2_buf_4 fanout110 (.X(net110),
    .A(ui_in[6]));
 sg13g2_buf_1 fanout111 (.A(ui_in[6]),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(net113),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(ui_in[5]),
    .X(net113));
 sg13g2_buf_4 fanout114 (.X(net114),
    .A(net115));
 sg13g2_buf_2 fanout115 (.A(net1),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(net118),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(net118),
    .X(net117));
 sg13g2_buf_1 fanout118 (.A(ui_in[3]),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(ui_in[2]),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(ui_in[2]),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(ui_in[2]),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(net126),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(net125),
    .X(net123));
 sg13g2_buf_1 fanout124 (.A(net125),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(net126),
    .X(net125));
 sg13g2_buf_1 fanout126 (.A(ui_in[1]),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(net128),
    .X(net127));
 sg13g2_buf_1 fanout128 (.A(net130),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(net130),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(ui_in[0]),
    .X(net130));
 sg13g2_buf_1 input1 (.A(ui_in[4]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[7]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(uio_in[0]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[1]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(uio_in[2]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(uio_in[3]),
    .X(net6));
 sg13g2_tielo \proj_15.gate7/_0__7  (.L_LO(net7));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_fill_2 FILLER_19_245 ();
 sg13g2_fill_1 FILLER_19_247 ();
 sg13g2_decap_8 FILLER_19_253 ();
 sg13g2_fill_2 FILLER_19_260 ();
 sg13g2_fill_1 FILLER_19_268 ();
 sg13g2_decap_8 FILLER_19_277 ();
 sg13g2_decap_4 FILLER_19_284 ();
 sg13g2_fill_2 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_293 ();
 sg13g2_decap_8 FILLER_19_300 ();
 sg13g2_decap_8 FILLER_19_307 ();
 sg13g2_decap_8 FILLER_19_314 ();
 sg13g2_decap_8 FILLER_19_321 ();
 sg13g2_decap_8 FILLER_19_328 ();
 sg13g2_decap_8 FILLER_19_335 ();
 sg13g2_decap_8 FILLER_19_342 ();
 sg13g2_decap_8 FILLER_19_349 ();
 sg13g2_decap_8 FILLER_19_356 ();
 sg13g2_decap_8 FILLER_19_363 ();
 sg13g2_decap_8 FILLER_19_370 ();
 sg13g2_decap_8 FILLER_19_377 ();
 sg13g2_decap_8 FILLER_19_384 ();
 sg13g2_decap_8 FILLER_19_391 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_fill_1 FILLER_20_210 ();
 sg13g2_fill_2 FILLER_20_219 ();
 sg13g2_fill_2 FILLER_20_224 ();
 sg13g2_fill_2 FILLER_20_247 ();
 sg13g2_decap_4 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_fill_2 FILLER_20_315 ();
 sg13g2_fill_1 FILLER_20_317 ();
 sg13g2_decap_8 FILLER_20_321 ();
 sg13g2_decap_8 FILLER_20_328 ();
 sg13g2_decap_8 FILLER_20_335 ();
 sg13g2_decap_8 FILLER_20_342 ();
 sg13g2_decap_8 FILLER_20_349 ();
 sg13g2_decap_8 FILLER_20_356 ();
 sg13g2_decap_8 FILLER_20_363 ();
 sg13g2_decap_8 FILLER_20_370 ();
 sg13g2_decap_8 FILLER_20_377 ();
 sg13g2_decap_8 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_fill_2 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_fill_2 FILLER_21_203 ();
 sg13g2_fill_2 FILLER_21_208 ();
 sg13g2_decap_8 FILLER_21_239 ();
 sg13g2_fill_2 FILLER_21_249 ();
 sg13g2_fill_1 FILLER_21_251 ();
 sg13g2_decap_8 FILLER_21_257 ();
 sg13g2_decap_4 FILLER_21_264 ();
 sg13g2_fill_1 FILLER_21_268 ();
 sg13g2_fill_1 FILLER_21_272 ();
 sg13g2_decap_8 FILLER_21_283 ();
 sg13g2_fill_1 FILLER_21_290 ();
 sg13g2_fill_1 FILLER_21_296 ();
 sg13g2_decap_4 FILLER_21_302 ();
 sg13g2_fill_1 FILLER_21_306 ();
 sg13g2_decap_4 FILLER_21_310 ();
 sg13g2_fill_2 FILLER_21_314 ();
 sg13g2_fill_1 FILLER_21_324 ();
 sg13g2_decap_8 FILLER_21_335 ();
 sg13g2_decap_8 FILLER_21_342 ();
 sg13g2_decap_8 FILLER_21_349 ();
 sg13g2_decap_8 FILLER_21_356 ();
 sg13g2_decap_8 FILLER_21_363 ();
 sg13g2_decap_8 FILLER_21_370 ();
 sg13g2_decap_8 FILLER_21_377 ();
 sg13g2_decap_8 FILLER_21_384 ();
 sg13g2_decap_8 FILLER_21_391 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_4 FILLER_22_182 ();
 sg13g2_fill_2 FILLER_22_209 ();
 sg13g2_decap_8 FILLER_22_236 ();
 sg13g2_fill_1 FILLER_22_243 ();
 sg13g2_fill_2 FILLER_22_269 ();
 sg13g2_fill_2 FILLER_22_291 ();
 sg13g2_fill_2 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_339 ();
 sg13g2_decap_8 FILLER_22_346 ();
 sg13g2_decap_8 FILLER_22_353 ();
 sg13g2_decap_8 FILLER_22_360 ();
 sg13g2_decap_8 FILLER_22_367 ();
 sg13g2_decap_8 FILLER_22_374 ();
 sg13g2_decap_8 FILLER_22_381 ();
 sg13g2_decap_8 FILLER_22_388 ();
 sg13g2_decap_8 FILLER_22_395 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_4 FILLER_23_175 ();
 sg13g2_fill_1 FILLER_23_179 ();
 sg13g2_fill_1 FILLER_23_183 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_4 FILLER_23_211 ();
 sg13g2_decap_4 FILLER_23_250 ();
 sg13g2_fill_1 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_270 ();
 sg13g2_decap_4 FILLER_23_297 ();
 sg13g2_fill_2 FILLER_23_301 ();
 sg13g2_fill_1 FILLER_23_316 ();
 sg13g2_fill_2 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_332 ();
 sg13g2_decap_8 FILLER_23_339 ();
 sg13g2_fill_2 FILLER_23_346 ();
 sg13g2_decap_8 FILLER_23_353 ();
 sg13g2_decap_8 FILLER_23_360 ();
 sg13g2_decap_8 FILLER_23_367 ();
 sg13g2_decap_8 FILLER_23_374 ();
 sg13g2_decap_8 FILLER_23_381 ();
 sg13g2_decap_8 FILLER_23_388 ();
 sg13g2_decap_8 FILLER_23_395 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_4 FILLER_24_168 ();
 sg13g2_fill_1 FILLER_24_172 ();
 sg13g2_decap_4 FILLER_24_201 ();
 sg13g2_fill_1 FILLER_24_205 ();
 sg13g2_decap_8 FILLER_24_216 ();
 sg13g2_decap_4 FILLER_24_223 ();
 sg13g2_fill_2 FILLER_24_237 ();
 sg13g2_fill_1 FILLER_24_239 ();
 sg13g2_fill_1 FILLER_24_255 ();
 sg13g2_decap_4 FILLER_24_271 ();
 sg13g2_fill_2 FILLER_24_275 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_4 FILLER_24_294 ();
 sg13g2_fill_2 FILLER_24_298 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_fill_2 FILLER_24_315 ();
 sg13g2_fill_1 FILLER_24_317 ();
 sg13g2_fill_1 FILLER_24_341 ();
 sg13g2_decap_8 FILLER_24_363 ();
 sg13g2_decap_8 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_377 ();
 sg13g2_decap_8 FILLER_24_384 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_4 FILLER_25_175 ();
 sg13g2_fill_2 FILLER_25_179 ();
 sg13g2_decap_8 FILLER_25_199 ();
 sg13g2_fill_2 FILLER_25_206 ();
 sg13g2_fill_1 FILLER_25_208 ();
 sg13g2_fill_2 FILLER_25_239 ();
 sg13g2_fill_1 FILLER_25_241 ();
 sg13g2_fill_2 FILLER_25_247 ();
 sg13g2_decap_4 FILLER_25_264 ();
 sg13g2_fill_2 FILLER_25_268 ();
 sg13g2_fill_2 FILLER_25_295 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_fill_2 FILLER_25_322 ();
 sg13g2_fill_2 FILLER_25_329 ();
 sg13g2_fill_1 FILLER_25_339 ();
 sg13g2_fill_2 FILLER_25_345 ();
 sg13g2_fill_1 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_25_363 ();
 sg13g2_decap_8 FILLER_25_370 ();
 sg13g2_decap_8 FILLER_25_377 ();
 sg13g2_decap_8 FILLER_25_384 ();
 sg13g2_decap_8 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_fill_2 FILLER_26_182 ();
 sg13g2_fill_2 FILLER_26_199 ();
 sg13g2_fill_1 FILLER_26_201 ();
 sg13g2_decap_4 FILLER_26_207 ();
 sg13g2_fill_1 FILLER_26_211 ();
 sg13g2_decap_8 FILLER_26_227 ();
 sg13g2_decap_4 FILLER_26_234 ();
 sg13g2_decap_8 FILLER_26_243 ();
 sg13g2_fill_2 FILLER_26_250 ();
 sg13g2_fill_1 FILLER_26_252 ();
 sg13g2_fill_1 FILLER_26_258 ();
 sg13g2_decap_8 FILLER_26_264 ();
 sg13g2_decap_8 FILLER_26_271 ();
 sg13g2_fill_2 FILLER_26_278 ();
 sg13g2_decap_4 FILLER_26_288 ();
 sg13g2_fill_2 FILLER_26_297 ();
 sg13g2_fill_1 FILLER_26_304 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_fill_1 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_361 ();
 sg13g2_decap_8 FILLER_26_368 ();
 sg13g2_decap_8 FILLER_26_375 ();
 sg13g2_decap_8 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_fill_1 FILLER_27_224 ();
 sg13g2_fill_1 FILLER_27_230 ();
 sg13g2_fill_1 FILLER_27_236 ();
 sg13g2_decap_8 FILLER_27_241 ();
 sg13g2_fill_1 FILLER_27_248 ();
 sg13g2_decap_8 FILLER_27_254 ();
 sg13g2_decap_4 FILLER_27_261 ();
 sg13g2_fill_2 FILLER_27_281 ();
 sg13g2_fill_1 FILLER_27_283 ();
 sg13g2_decap_4 FILLER_27_300 ();
 sg13g2_decap_8 FILLER_27_314 ();
 sg13g2_fill_2 FILLER_27_321 ();
 sg13g2_decap_8 FILLER_27_338 ();
 sg13g2_fill_2 FILLER_27_345 ();
 sg13g2_fill_1 FILLER_27_347 ();
 sg13g2_decap_8 FILLER_27_363 ();
 sg13g2_decap_8 FILLER_27_370 ();
 sg13g2_decap_8 FILLER_27_377 ();
 sg13g2_decap_8 FILLER_27_384 ();
 sg13g2_decap_8 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_fill_2 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_167 ();
 sg13g2_decap_8 FILLER_28_174 ();
 sg13g2_fill_2 FILLER_28_181 ();
 sg13g2_fill_1 FILLER_28_183 ();
 sg13g2_fill_2 FILLER_28_188 ();
 sg13g2_decap_8 FILLER_28_194 ();
 sg13g2_decap_8 FILLER_28_201 ();
 sg13g2_decap_8 FILLER_28_208 ();
 sg13g2_decap_8 FILLER_28_215 ();
 sg13g2_decap_4 FILLER_28_222 ();
 sg13g2_fill_1 FILLER_28_259 ();
 sg13g2_fill_2 FILLER_28_269 ();
 sg13g2_decap_4 FILLER_28_280 ();
 sg13g2_fill_1 FILLER_28_284 ();
 sg13g2_decap_4 FILLER_28_290 ();
 sg13g2_fill_1 FILLER_28_302 ();
 sg13g2_fill_1 FILLER_28_308 ();
 sg13g2_fill_2 FILLER_28_314 ();
 sg13g2_fill_1 FILLER_28_316 ();
 sg13g2_decap_4 FILLER_28_342 ();
 sg13g2_decap_8 FILLER_28_366 ();
 sg13g2_decap_8 FILLER_28_373 ();
 sg13g2_decap_8 FILLER_28_380 ();
 sg13g2_decap_8 FILLER_28_387 ();
 sg13g2_decap_8 FILLER_28_394 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_206 ();
 sg13g2_decap_4 FILLER_29_213 ();
 sg13g2_fill_1 FILLER_29_222 ();
 sg13g2_decap_4 FILLER_29_240 ();
 sg13g2_fill_2 FILLER_29_244 ();
 sg13g2_decap_4 FILLER_29_272 ();
 sg13g2_fill_1 FILLER_29_284 ();
 sg13g2_fill_2 FILLER_29_291 ();
 sg13g2_decap_4 FILLER_29_326 ();
 sg13g2_fill_2 FILLER_29_340 ();
 sg13g2_fill_1 FILLER_29_342 ();
 sg13g2_fill_1 FILLER_29_347 ();
 sg13g2_decap_8 FILLER_29_358 ();
 sg13g2_decap_4 FILLER_29_365 ();
 sg13g2_fill_1 FILLER_29_369 ();
 sg13g2_decap_8 FILLER_29_382 ();
 sg13g2_decap_8 FILLER_29_389 ();
 sg13g2_decap_8 FILLER_29_396 ();
 sg13g2_decap_4 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_fill_1 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_173 ();
 sg13g2_decap_8 FILLER_30_180 ();
 sg13g2_fill_2 FILLER_30_187 ();
 sg13g2_fill_1 FILLER_30_189 ();
 sg13g2_fill_2 FILLER_30_216 ();
 sg13g2_fill_1 FILLER_30_218 ();
 sg13g2_decap_4 FILLER_30_224 ();
 sg13g2_decap_4 FILLER_30_260 ();
 sg13g2_fill_2 FILLER_30_264 ();
 sg13g2_decap_4 FILLER_30_283 ();
 sg13g2_decap_8 FILLER_30_309 ();
 sg13g2_fill_2 FILLER_30_316 ();
 sg13g2_decap_4 FILLER_30_323 ();
 sg13g2_fill_1 FILLER_30_337 ();
 sg13g2_fill_1 FILLER_30_354 ();
 sg13g2_fill_1 FILLER_30_368 ();
 sg13g2_decap_8 FILLER_30_387 ();
 sg13g2_decap_8 FILLER_30_394 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_fill_1 FILLER_31_182 ();
 sg13g2_fill_2 FILLER_31_187 ();
 sg13g2_fill_1 FILLER_31_193 ();
 sg13g2_fill_2 FILLER_31_198 ();
 sg13g2_decap_8 FILLER_31_204 ();
 sg13g2_fill_2 FILLER_31_211 ();
 sg13g2_fill_1 FILLER_31_218 ();
 sg13g2_decap_4 FILLER_31_234 ();
 sg13g2_decap_4 FILLER_31_241 ();
 sg13g2_fill_1 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_268 ();
 sg13g2_decap_8 FILLER_31_287 ();
 sg13g2_decap_4 FILLER_31_304 ();
 sg13g2_fill_2 FILLER_31_318 ();
 sg13g2_fill_2 FILLER_31_340 ();
 sg13g2_fill_1 FILLER_31_342 ();
 sg13g2_decap_8 FILLER_31_348 ();
 sg13g2_decap_4 FILLER_31_355 ();
 sg13g2_fill_2 FILLER_31_364 ();
 sg13g2_fill_1 FILLER_31_371 ();
 sg13g2_decap_8 FILLER_31_382 ();
 sg13g2_decap_8 FILLER_31_389 ();
 sg13g2_decap_8 FILLER_31_396 ();
 sg13g2_decap_4 FILLER_31_403 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_fill_2 FILLER_32_175 ();
 sg13g2_fill_1 FILLER_32_177 ();
 sg13g2_decap_8 FILLER_32_204 ();
 sg13g2_fill_1 FILLER_32_211 ();
 sg13g2_decap_4 FILLER_32_227 ();
 sg13g2_decap_4 FILLER_32_251 ();
 sg13g2_decap_8 FILLER_32_266 ();
 sg13g2_fill_1 FILLER_32_273 ();
 sg13g2_decap_8 FILLER_32_280 ();
 sg13g2_decap_4 FILLER_32_292 ();
 sg13g2_fill_2 FILLER_32_296 ();
 sg13g2_decap_8 FILLER_32_310 ();
 sg13g2_decap_4 FILLER_32_317 ();
 sg13g2_fill_2 FILLER_32_321 ();
 sg13g2_fill_2 FILLER_32_333 ();
 sg13g2_fill_1 FILLER_32_354 ();
 sg13g2_fill_1 FILLER_32_368 ();
 sg13g2_decap_8 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_4 FILLER_33_201 ();
 sg13g2_fill_1 FILLER_33_205 ();
 sg13g2_decap_4 FILLER_33_220 ();
 sg13g2_fill_1 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_243 ();
 sg13g2_fill_1 FILLER_33_255 ();
 sg13g2_fill_2 FILLER_33_268 ();
 sg13g2_fill_2 FILLER_33_287 ();
 sg13g2_decap_8 FILLER_33_309 ();
 sg13g2_fill_1 FILLER_33_316 ();
 sg13g2_decap_8 FILLER_33_331 ();
 sg13g2_decap_4 FILLER_33_357 ();
 sg13g2_decap_8 FILLER_33_379 ();
 sg13g2_decap_8 FILLER_33_386 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_4 FILLER_34_175 ();
 sg13g2_fill_1 FILLER_34_179 ();
 sg13g2_fill_2 FILLER_34_184 ();
 sg13g2_decap_4 FILLER_34_190 ();
 sg13g2_fill_2 FILLER_34_194 ();
 sg13g2_fill_2 FILLER_34_200 ();
 sg13g2_decap_8 FILLER_34_206 ();
 sg13g2_decap_4 FILLER_34_213 ();
 sg13g2_fill_2 FILLER_34_217 ();
 sg13g2_fill_1 FILLER_34_250 ();
 sg13g2_decap_4 FILLER_34_268 ();
 sg13g2_fill_2 FILLER_34_284 ();
 sg13g2_fill_1 FILLER_34_286 ();
 sg13g2_decap_8 FILLER_34_303 ();
 sg13g2_fill_2 FILLER_34_310 ();
 sg13g2_fill_1 FILLER_34_312 ();
 sg13g2_decap_8 FILLER_34_328 ();
 sg13g2_decap_4 FILLER_34_335 ();
 sg13g2_fill_2 FILLER_34_339 ();
 sg13g2_decap_8 FILLER_34_359 ();
 sg13g2_decap_8 FILLER_34_366 ();
 sg13g2_decap_8 FILLER_34_373 ();
 sg13g2_decap_8 FILLER_34_380 ();
 sg13g2_decap_8 FILLER_34_387 ();
 sg13g2_decap_8 FILLER_34_394 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_fill_2 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_fill_1 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_235 ();
 sg13g2_decap_8 FILLER_35_242 ();
 sg13g2_fill_1 FILLER_35_249 ();
 sg13g2_fill_2 FILLER_35_253 ();
 sg13g2_fill_1 FILLER_35_269 ();
 sg13g2_fill_2 FILLER_35_275 ();
 sg13g2_fill_1 FILLER_35_297 ();
 sg13g2_decap_4 FILLER_35_305 ();
 sg13g2_fill_1 FILLER_35_309 ();
 sg13g2_fill_2 FILLER_35_316 ();
 sg13g2_fill_2 FILLER_35_343 ();
 sg13g2_fill_1 FILLER_35_345 ();
 sg13g2_decap_8 FILLER_35_359 ();
 sg13g2_decap_8 FILLER_35_366 ();
 sg13g2_decap_8 FILLER_35_373 ();
 sg13g2_decap_8 FILLER_35_380 ();
 sg13g2_decap_8 FILLER_35_387 ();
 sg13g2_decap_8 FILLER_35_394 ();
 sg13g2_decap_8 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_fill_2 FILLER_36_217 ();
 sg13g2_fill_2 FILLER_36_242 ();
 sg13g2_fill_1 FILLER_36_244 ();
 sg13g2_decap_4 FILLER_36_254 ();
 sg13g2_fill_2 FILLER_36_285 ();
 sg13g2_fill_1 FILLER_36_287 ();
 sg13g2_fill_1 FILLER_36_310 ();
 sg13g2_decap_4 FILLER_36_320 ();
 sg13g2_fill_2 FILLER_36_324 ();
 sg13g2_decap_8 FILLER_36_344 ();
 sg13g2_decap_8 FILLER_36_351 ();
 sg13g2_decap_8 FILLER_36_358 ();
 sg13g2_decap_8 FILLER_36_365 ();
 sg13g2_decap_8 FILLER_36_372 ();
 sg13g2_decap_8 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_36_386 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_fill_2 FILLER_37_245 ();
 sg13g2_fill_2 FILLER_37_267 ();
 sg13g2_fill_1 FILLER_37_269 ();
 sg13g2_decap_8 FILLER_37_309 ();
 sg13g2_decap_8 FILLER_37_316 ();
 sg13g2_decap_8 FILLER_37_323 ();
 sg13g2_decap_8 FILLER_37_330 ();
 sg13g2_decap_8 FILLER_37_337 ();
 sg13g2_decap_8 FILLER_37_344 ();
 sg13g2_decap_8 FILLER_37_351 ();
 sg13g2_decap_8 FILLER_37_358 ();
 sg13g2_decap_8 FILLER_37_365 ();
 sg13g2_decap_8 FILLER_37_372 ();
 sg13g2_decap_8 FILLER_37_379 ();
 sg13g2_decap_8 FILLER_37_386 ();
 sg13g2_decap_8 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_250 ();
 sg13g2_fill_2 FILLER_38_257 ();
 sg13g2_decap_8 FILLER_38_263 ();
 sg13g2_fill_2 FILLER_38_270 ();
 sg13g2_fill_2 FILLER_38_277 ();
 sg13g2_fill_1 FILLER_38_279 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_fill_1 FILLER_38_287 ();
 sg13g2_fill_2 FILLER_38_309 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_decap_8 FILLER_38_316 ();
 sg13g2_decap_8 FILLER_38_323 ();
 sg13g2_decap_4 FILLER_38_330 ();
 sg13g2_fill_2 FILLER_38_334 ();
 sg13g2_decap_8 FILLER_38_340 ();
 sg13g2_decap_8 FILLER_38_347 ();
 sg13g2_decap_8 FILLER_38_354 ();
 sg13g2_decap_8 FILLER_38_361 ();
 sg13g2_decap_8 FILLER_38_368 ();
 sg13g2_decap_8 FILLER_38_375 ();
 sg13g2_decap_8 FILLER_38_382 ();
 sg13g2_decap_8 FILLER_38_389 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net17;
 assign uio_oe[1] = net18;
 assign uio_oe[2] = net19;
 assign uio_oe[3] = net20;
 assign uio_oe[4] = net21;
 assign uio_oe[5] = net22;
 assign uio_oe[6] = net23;
 assign uio_oe[7] = net24;
 assign uio_out[0] = net25;
 assign uio_out[1] = net26;
 assign uio_out[2] = net27;
 assign uio_out[3] = net28;
 assign uio_out[4] = net29;
 assign uio_out[5] = net30;
 assign uio_out[6] = net31;
 assign uio_out[7] = net32;
endmodule

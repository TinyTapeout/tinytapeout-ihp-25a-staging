module tt_um_tmkong_rgb_mixer (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire \enc0[0] ;
 wire \enc0[1] ;
 wire \enc0[2] ;
 wire \enc0[3] ;
 wire \enc0[4] ;
 wire \enc0[5] ;
 wire \enc0[6] ;
 wire \enc0[7] ;
 wire \enc1[0] ;
 wire \enc1[1] ;
 wire \enc1[2] ;
 wire \enc1[3] ;
 wire \enc1[4] ;
 wire \enc1[5] ;
 wire \enc1[6] ;
 wire \enc1[7] ;
 wire \enc2[0] ;
 wire \enc2[1] ;
 wire \enc2[2] ;
 wire \enc2[3] ;
 wire \enc2[4] ;
 wire \enc2[5] ;
 wire \enc2[6] ;
 wire \enc2[7] ;
 wire \rgb_mixer.debounce0_a.button_hist[0] ;
 wire \rgb_mixer.debounce0_a.button_hist[1] ;
 wire \rgb_mixer.debounce0_a.button_hist[2] ;
 wire \rgb_mixer.debounce0_a.button_hist[3] ;
 wire \rgb_mixer.debounce0_a.button_hist[4] ;
 wire \rgb_mixer.debounce0_a.button_hist[5] ;
 wire \rgb_mixer.debounce0_a.button_hist[6] ;
 wire \rgb_mixer.debounce0_a.button_hist[7] ;
 wire \rgb_mixer.debounce0_a.debounced ;
 wire \rgb_mixer.debounce0_b.button_hist[0] ;
 wire \rgb_mixer.debounce0_b.button_hist[1] ;
 wire \rgb_mixer.debounce0_b.button_hist[2] ;
 wire \rgb_mixer.debounce0_b.button_hist[3] ;
 wire \rgb_mixer.debounce0_b.button_hist[4] ;
 wire \rgb_mixer.debounce0_b.button_hist[5] ;
 wire \rgb_mixer.debounce0_b.button_hist[6] ;
 wire \rgb_mixer.debounce0_b.button_hist[7] ;
 wire \rgb_mixer.debounce0_b.debounced ;
 wire \rgb_mixer.debounce1_a.button_hist[0] ;
 wire \rgb_mixer.debounce1_a.button_hist[1] ;
 wire \rgb_mixer.debounce1_a.button_hist[2] ;
 wire \rgb_mixer.debounce1_a.button_hist[3] ;
 wire \rgb_mixer.debounce1_a.button_hist[4] ;
 wire \rgb_mixer.debounce1_a.button_hist[5] ;
 wire \rgb_mixer.debounce1_a.button_hist[6] ;
 wire \rgb_mixer.debounce1_a.button_hist[7] ;
 wire \rgb_mixer.debounce1_a.debounced ;
 wire \rgb_mixer.debounce1_b.button_hist[0] ;
 wire \rgb_mixer.debounce1_b.button_hist[1] ;
 wire \rgb_mixer.debounce1_b.button_hist[2] ;
 wire \rgb_mixer.debounce1_b.button_hist[3] ;
 wire \rgb_mixer.debounce1_b.button_hist[4] ;
 wire \rgb_mixer.debounce1_b.button_hist[5] ;
 wire \rgb_mixer.debounce1_b.button_hist[6] ;
 wire \rgb_mixer.debounce1_b.button_hist[7] ;
 wire \rgb_mixer.debounce1_b.debounced ;
 wire \rgb_mixer.debounce2_a.button_hist[0] ;
 wire \rgb_mixer.debounce2_a.button_hist[1] ;
 wire \rgb_mixer.debounce2_a.button_hist[2] ;
 wire \rgb_mixer.debounce2_a.button_hist[3] ;
 wire \rgb_mixer.debounce2_a.button_hist[4] ;
 wire \rgb_mixer.debounce2_a.button_hist[5] ;
 wire \rgb_mixer.debounce2_a.button_hist[6] ;
 wire \rgb_mixer.debounce2_a.button_hist[7] ;
 wire \rgb_mixer.debounce2_a.debounced ;
 wire \rgb_mixer.debounce2_b.button_hist[0] ;
 wire \rgb_mixer.debounce2_b.button_hist[1] ;
 wire \rgb_mixer.debounce2_b.button_hist[2] ;
 wire \rgb_mixer.debounce2_b.button_hist[3] ;
 wire \rgb_mixer.debounce2_b.button_hist[4] ;
 wire \rgb_mixer.debounce2_b.button_hist[5] ;
 wire \rgb_mixer.debounce2_b.button_hist[6] ;
 wire \rgb_mixer.debounce2_b.button_hist[7] ;
 wire \rgb_mixer.debounce2_b.debounced ;
 wire \rgb_mixer.encoder0.old_a ;
 wire \rgb_mixer.encoder0.old_b ;
 wire \rgb_mixer.encoder1.old_a ;
 wire \rgb_mixer.encoder1.old_b ;
 wire \rgb_mixer.encoder2.old_a ;
 wire \rgb_mixer.encoder2.old_b ;
 wire \rgb_mixer.pwm0.count[0] ;
 wire \rgb_mixer.pwm0.count[1] ;
 wire \rgb_mixer.pwm0.count[2] ;
 wire \rgb_mixer.pwm0.count[3] ;
 wire \rgb_mixer.pwm0.count[4] ;
 wire \rgb_mixer.pwm0.count[5] ;
 wire \rgb_mixer.pwm0.count[6] ;
 wire \rgb_mixer.pwm0.count[7] ;
 wire \rgb_mixer.pwm0.out ;
 wire \rgb_mixer.pwm1.count[0] ;
 wire \rgb_mixer.pwm1.count[1] ;
 wire \rgb_mixer.pwm1.count[2] ;
 wire \rgb_mixer.pwm1.count[3] ;
 wire \rgb_mixer.pwm1.count[4] ;
 wire \rgb_mixer.pwm1.count[5] ;
 wire \rgb_mixer.pwm1.count[6] ;
 wire \rgb_mixer.pwm1.count[7] ;
 wire \rgb_mixer.pwm1.out ;
 wire \rgb_mixer.pwm2.count[0] ;
 wire \rgb_mixer.pwm2.count[1] ;
 wire \rgb_mixer.pwm2.count[2] ;
 wire \rgb_mixer.pwm2.count[3] ;
 wire \rgb_mixer.pwm2.count[4] ;
 wire \rgb_mixer.pwm2.count[5] ;
 wire \rgb_mixer.pwm2.count[6] ;
 wire \rgb_mixer.pwm2.count[7] ;
 wire \rgb_mixer.pwm2.out ;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire clknet_0_clk;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;

 sg13g2_inv_1 _0692_ (.Y(_0117_),
    .A(\enc0[2] ));
 sg13g2_inv_1 _0693_ (.Y(_0118_),
    .A(\enc0[1] ));
 sg13g2_inv_1 _0694_ (.Y(_0119_),
    .A(\enc0[0] ));
 sg13g2_inv_1 _0695_ (.Y(_0120_),
    .A(net285));
 sg13g2_inv_1 _0696_ (.Y(_0121_),
    .A(net291));
 sg13g2_inv_1 _0697_ (.Y(_0122_),
    .A(\enc1[4] ));
 sg13g2_inv_1 _0698_ (.Y(_0123_),
    .A(\enc1[1] ));
 sg13g2_inv_1 _0699_ (.Y(_0124_),
    .A(\enc1[0] ));
 sg13g2_inv_1 _0700_ (.Y(_0125_),
    .A(net287));
 sg13g2_inv_1 _0701_ (.Y(_0126_),
    .A(\enc2[4] ));
 sg13g2_inv_1 _0702_ (.Y(_0127_),
    .A(\enc2[2] ));
 sg13g2_inv_1 _0703_ (.Y(_0128_),
    .A(\enc2[1] ));
 sg13g2_inv_1 _0704_ (.Y(_0129_),
    .A(\enc2[0] ));
 sg13g2_inv_1 _0705_ (.Y(_0130_),
    .A(net201));
 sg13g2_inv_1 _0706_ (.Y(_0131_),
    .A(net193));
 sg13g2_inv_1 _0707_ (.Y(_0132_),
    .A(net236));
 sg13g2_inv_1 _0708_ (.Y(_0133_),
    .A(\rgb_mixer.pwm1.count[6] ));
 sg13g2_inv_1 _0709_ (.Y(_0134_),
    .A(net282));
 sg13g2_inv_1 _0710_ (.Y(_0135_),
    .A(\rgb_mixer.pwm1.count[2] ));
 sg13g2_inv_1 _0711_ (.Y(_0136_),
    .A(net263));
 sg13g2_inv_1 _0712_ (.Y(_0137_),
    .A(\rgb_mixer.pwm2.count[4] ));
 sg13g2_inv_1 _0713_ (.Y(_0138_),
    .A(net299));
 sg13g2_inv_1 _0714_ (.Y(_0139_),
    .A(net239));
 sg13g2_inv_1 _0715_ (.Y(_0140_),
    .A(\rgb_mixer.pwm0.count[6] ));
 sg13g2_inv_1 _0716_ (.Y(_0141_),
    .A(\rgb_mixer.pwm0.count[5] ));
 sg13g2_inv_1 _0717_ (.Y(_0142_),
    .A(net279));
 sg13g2_inv_1 _0718_ (.Y(_0143_),
    .A(net91));
 sg13g2_nor2b_2 _0719_ (.A(net8),
    .B_N(net7),
    .Y(_0144_));
 sg13g2_nand2_1 _0720_ (.Y(_0145_),
    .A(\enc1[0] ),
    .B(_0144_));
 sg13g2_nor2_2 _0721_ (.A(net7),
    .B(net8),
    .Y(_0146_));
 sg13g2_nor2b_2 _0722_ (.A(net7),
    .B_N(net8),
    .Y(_0147_));
 sg13g2_a22oi_1 _0723_ (.Y(_0148_),
    .B1(_0147_),
    .B2(\enc2[0] ),
    .A2(_0146_),
    .A1(\enc0[0] ));
 sg13g2_nand2_2 _0724_ (.Y(uio_out[0]),
    .A(_0145_),
    .B(_0148_));
 sg13g2_nand2_1 _0725_ (.Y(_0149_),
    .A(\enc1[1] ),
    .B(_0144_));
 sg13g2_a22oi_1 _0726_ (.Y(_0150_),
    .B1(_0147_),
    .B2(\enc2[1] ),
    .A2(_0146_),
    .A1(\enc0[1] ));
 sg13g2_nand2_2 _0727_ (.Y(uio_out[1]),
    .A(_0149_),
    .B(_0150_));
 sg13g2_nand2_1 _0728_ (.Y(_0151_),
    .A(\enc1[2] ),
    .B(_0144_));
 sg13g2_a22oi_1 _0729_ (.Y(_0152_),
    .B1(_0147_),
    .B2(\enc2[2] ),
    .A2(_0146_),
    .A1(\enc0[2] ));
 sg13g2_nand2_2 _0730_ (.Y(uio_out[2]),
    .A(_0151_),
    .B(_0152_));
 sg13g2_nand2_1 _0731_ (.Y(_0153_),
    .A(\enc1[3] ),
    .B(_0144_));
 sg13g2_a22oi_1 _0732_ (.Y(_0154_),
    .B1(_0147_),
    .B2(\enc2[3] ),
    .A2(_0146_),
    .A1(\enc0[3] ));
 sg13g2_nand2_2 _0733_ (.Y(uio_out[3]),
    .A(_0153_),
    .B(_0154_));
 sg13g2_nand2_1 _0734_ (.Y(_0155_),
    .A(\enc1[4] ),
    .B(_0144_));
 sg13g2_a22oi_1 _0735_ (.Y(_0156_),
    .B1(_0147_),
    .B2(\enc2[4] ),
    .A2(_0146_),
    .A1(\enc0[4] ));
 sg13g2_nand2_2 _0736_ (.Y(uio_out[4]),
    .A(_0155_),
    .B(_0156_));
 sg13g2_nand2_1 _0737_ (.Y(_0157_),
    .A(\enc1[5] ),
    .B(_0144_));
 sg13g2_a22oi_1 _0738_ (.Y(_0158_),
    .B1(_0147_),
    .B2(\enc2[5] ),
    .A2(_0146_),
    .A1(\enc0[5] ));
 sg13g2_nand2_2 _0739_ (.Y(uio_out[5]),
    .A(_0157_),
    .B(_0158_));
 sg13g2_nand2_1 _0740_ (.Y(_0159_),
    .A(\enc1[6] ),
    .B(_0144_));
 sg13g2_a22oi_1 _0741_ (.Y(_0160_),
    .B1(_0147_),
    .B2(\enc2[6] ),
    .A2(_0146_),
    .A1(\enc0[6] ));
 sg13g2_nand2_2 _0742_ (.Y(uio_out[6]),
    .A(_0159_),
    .B(_0160_));
 sg13g2_nand2_1 _0743_ (.Y(_0161_),
    .A(\enc1[7] ),
    .B(_0144_));
 sg13g2_a22oi_1 _0744_ (.Y(_0162_),
    .B1(_0147_),
    .B2(\enc2[7] ),
    .A2(_0146_),
    .A1(\enc0[7] ));
 sg13g2_nand2_2 _0745_ (.Y(uio_out[7]),
    .A(_0161_),
    .B(_0162_));
 sg13g2_and2_1 _0746_ (.A(net158),
    .B(net88),
    .X(_0006_));
 sg13g2_xnor2_1 _0747_ (.Y(_0163_),
    .A(\rgb_mixer.pwm2.count[0] ),
    .B(net270));
 sg13g2_nor2_1 _0748_ (.A(net84),
    .B(net271),
    .Y(_0007_));
 sg13g2_a21oi_1 _0749_ (.A1(\rgb_mixer.pwm2.count[0] ),
    .A2(\rgb_mixer.pwm2.count[1] ),
    .Y(_0164_),
    .B1(net243));
 sg13g2_nand3_1 _0750_ (.B(\rgb_mixer.pwm2.count[2] ),
    .C(\rgb_mixer.pwm2.count[1] ),
    .A(\rgb_mixer.pwm2.count[0] ),
    .Y(_0165_));
 sg13g2_nand2_1 _0751_ (.Y(_0166_),
    .A(net91),
    .B(_0165_));
 sg13g2_nor2_1 _0752_ (.A(net244),
    .B(_0166_),
    .Y(_0008_));
 sg13g2_nor2_1 _0753_ (.A(_0138_),
    .B(_0165_),
    .Y(_0167_));
 sg13g2_a21oi_1 _0754_ (.A1(_0138_),
    .A2(_0165_),
    .Y(_0168_),
    .B1(net84));
 sg13g2_nor2b_1 _0755_ (.A(_0167_),
    .B_N(_0168_),
    .Y(_0009_));
 sg13g2_nor2_1 _0756_ (.A(net259),
    .B(_0167_),
    .Y(_0169_));
 sg13g2_nor3_2 _0757_ (.A(_0137_),
    .B(_0138_),
    .C(_0165_),
    .Y(_0170_));
 sg13g2_nor3_1 _0758_ (.A(net84),
    .B(net260),
    .C(_0170_),
    .Y(_0010_));
 sg13g2_o21ai_1 _0759_ (.B1(net91),
    .Y(_0171_),
    .A1(net251),
    .A2(_0170_));
 sg13g2_a21oi_1 _0760_ (.A1(net251),
    .A2(_0170_),
    .Y(_0011_),
    .B1(_0171_));
 sg13g2_a21oi_1 _0761_ (.A1(\rgb_mixer.pwm2.count[5] ),
    .A2(_0170_),
    .Y(_0172_),
    .B1(net208));
 sg13g2_nand3_1 _0762_ (.B(net251),
    .C(_0170_),
    .A(net208),
    .Y(_0173_));
 sg13g2_nand2_1 _0763_ (.Y(_0174_),
    .A(net91),
    .B(_0173_));
 sg13g2_nor2_1 _0764_ (.A(net209),
    .B(_0174_),
    .Y(_0012_));
 sg13g2_o21ai_1 _0765_ (.B1(net92),
    .Y(_0175_),
    .A1(_0136_),
    .A2(_0173_));
 sg13g2_a21oi_1 _0766_ (.A1(_0136_),
    .A2(_0173_),
    .Y(_0013_),
    .B1(_0175_));
 sg13g2_and2_1 _0767_ (.A(net85),
    .B(net159),
    .X(_0014_));
 sg13g2_xnor2_1 _0768_ (.Y(_0176_),
    .A(\rgb_mixer.pwm1.count[0] ),
    .B(net267));
 sg13g2_nor2_1 _0769_ (.A(net83),
    .B(net268),
    .Y(_0015_));
 sg13g2_a21oi_1 _0770_ (.A1(\rgb_mixer.pwm1.count[0] ),
    .A2(\rgb_mixer.pwm1.count[1] ),
    .Y(_0177_),
    .B1(net217));
 sg13g2_nand3_1 _0771_ (.B(net217),
    .C(net267),
    .A(\rgb_mixer.pwm1.count[0] ),
    .Y(_0178_));
 sg13g2_nand2_1 _0772_ (.Y(_0179_),
    .A(net85),
    .B(_0178_));
 sg13g2_nor2_1 _0773_ (.A(net218),
    .B(_0179_),
    .Y(_0016_));
 sg13g2_nor2_1 _0774_ (.A(_0134_),
    .B(_0178_),
    .Y(_0180_));
 sg13g2_a21oi_1 _0775_ (.A1(_0134_),
    .A2(_0178_),
    .Y(_0181_),
    .B1(net83));
 sg13g2_nor2b_1 _0776_ (.A(_0180_),
    .B_N(net283),
    .Y(_0017_));
 sg13g2_nor2_1 _0777_ (.A(net265),
    .B(_0180_),
    .Y(_0182_));
 sg13g2_and2_1 _0778_ (.A(net265),
    .B(_0180_),
    .X(_0183_));
 sg13g2_nor3_1 _0779_ (.A(net83),
    .B(net266),
    .C(_0183_),
    .Y(_0018_));
 sg13g2_o21ai_1 _0780_ (.B1(net85),
    .Y(_0184_),
    .A1(net253),
    .A2(_0183_));
 sg13g2_a21oi_1 _0781_ (.A1(net253),
    .A2(_0183_),
    .Y(_0019_),
    .B1(_0184_));
 sg13g2_a21oi_1 _0782_ (.A1(\rgb_mixer.pwm1.count[5] ),
    .A2(_0183_),
    .Y(_0185_),
    .B1(net223));
 sg13g2_nand3_1 _0783_ (.B(\rgb_mixer.pwm1.count[5] ),
    .C(_0183_),
    .A(net223),
    .Y(_0186_));
 sg13g2_nand2_1 _0784_ (.Y(_0187_),
    .A(net85),
    .B(_0186_));
 sg13g2_nor2_1 _0785_ (.A(net224),
    .B(_0187_),
    .Y(_0020_));
 sg13g2_o21ai_1 _0786_ (.B1(net85),
    .Y(_0188_),
    .A1(_0132_),
    .A2(_0186_));
 sg13g2_a21oi_1 _0787_ (.A1(_0132_),
    .A2(_0186_),
    .Y(_0021_),
    .B1(_0188_));
 sg13g2_nand2_1 _0788_ (.Y(_0189_),
    .A(net275),
    .B(_0136_));
 sg13g2_nand2b_1 _0789_ (.Y(_0190_),
    .B(net208),
    .A_N(\enc2[6] ));
 sg13g2_nand2b_1 _0790_ (.Y(_0191_),
    .B(\enc2[6] ),
    .A_N(\rgb_mixer.pwm2.count[6] ));
 sg13g2_o21ai_1 _0791_ (.B1(_0191_),
    .Y(_0192_),
    .A1(_0125_),
    .A2(\rgb_mixer.pwm2.count[5] ));
 sg13g2_nand2_1 _0792_ (.Y(_0193_),
    .A(_0125_),
    .B(\rgb_mixer.pwm2.count[5] ));
 sg13g2_o21ai_1 _0793_ (.B1(_0193_),
    .Y(_0194_),
    .A1(\enc2[4] ),
    .A2(_0137_));
 sg13g2_nand2b_1 _0794_ (.Y(_0195_),
    .B(\rgb_mixer.pwm2.count[3] ),
    .A_N(\enc2[3] ));
 sg13g2_nor2_1 _0795_ (.A(_0127_),
    .B(\rgb_mixer.pwm2.count[2] ),
    .Y(_0196_));
 sg13g2_nand2b_1 _0796_ (.Y(_0197_),
    .B(\enc2[2] ),
    .A_N(\rgb_mixer.pwm2.count[2] ));
 sg13g2_nor2b_1 _0797_ (.A(\rgb_mixer.pwm2.count[3] ),
    .B_N(\enc2[3] ),
    .Y(_0198_));
 sg13g2_a21o_1 _0798_ (.A2(\rgb_mixer.pwm2.count[2] ),
    .A1(_0127_),
    .B1(_0198_),
    .X(_0199_));
 sg13g2_nand2b_1 _0799_ (.Y(_0200_),
    .B(\enc2[1] ),
    .A_N(\rgb_mixer.pwm2.count[1] ));
 sg13g2_nor2b_1 _0800_ (.A(\enc2[0] ),
    .B_N(\rgb_mixer.pwm2.count[0] ),
    .Y(_0201_));
 sg13g2_a21o_1 _0801_ (.A2(\rgb_mixer.pwm2.count[1] ),
    .A1(_0128_),
    .B1(_0201_),
    .X(_0202_));
 sg13g2_a21oi_1 _0802_ (.A1(_0200_),
    .A2(_0202_),
    .Y(_0203_),
    .B1(_0199_));
 sg13g2_o21ai_1 _0803_ (.B1(_0195_),
    .Y(_0204_),
    .A1(_0196_),
    .A2(_0203_));
 sg13g2_a21oi_1 _0804_ (.A1(\enc2[4] ),
    .A2(_0137_),
    .Y(_0205_),
    .B1(_0198_));
 sg13g2_a21oi_1 _0805_ (.A1(_0204_),
    .A2(_0205_),
    .Y(_0206_),
    .B1(_0194_));
 sg13g2_o21ai_1 _0806_ (.B1(_0190_),
    .Y(_0207_),
    .A1(_0192_),
    .A2(_0206_));
 sg13g2_nor4_1 _0807_ (.A(_0192_),
    .B(_0194_),
    .C(_0199_),
    .D(_0202_),
    .Y(_0208_));
 sg13g2_nor2_1 _0808_ (.A(_0129_),
    .B(\rgb_mixer.pwm2.count[0] ),
    .Y(_0209_));
 sg13g2_o21ai_1 _0809_ (.B1(_0200_),
    .Y(_0210_),
    .A1(_0126_),
    .A2(\rgb_mixer.pwm2.count[4] ));
 sg13g2_nand4_1 _0810_ (.B(_0190_),
    .C(_0195_),
    .A(_0189_),
    .Y(_0211_),
    .D(_0197_));
 sg13g2_nor3_1 _0811_ (.A(_0209_),
    .B(_0210_),
    .C(_0211_),
    .Y(_0212_));
 sg13g2_o21ai_1 _0812_ (.B1(net93),
    .Y(_0213_),
    .A1(net275),
    .A2(_0136_));
 sg13g2_a221oi_1 _0813_ (.B2(_0212_),
    .C1(_0213_),
    .B1(_0208_),
    .A1(_0189_),
    .Y(_0022_),
    .A2(_0207_));
 sg13g2_and2_1 _0814_ (.A(net86),
    .B(net160),
    .X(_0023_));
 sg13g2_o21ai_1 _0815_ (.B1(net86),
    .Y(_0214_),
    .A1(\rgb_mixer.pwm0.count[0] ),
    .A2(net241));
 sg13g2_a21oi_1 _0816_ (.A1(\rgb_mixer.pwm0.count[0] ),
    .A2(net241),
    .Y(_0024_),
    .B1(_0214_));
 sg13g2_a21oi_1 _0817_ (.A1(\rgb_mixer.pwm0.count[0] ),
    .A2(\rgb_mixer.pwm0.count[1] ),
    .Y(_0215_),
    .B1(net204));
 sg13g2_nand3_1 _0818_ (.B(net204),
    .C(net241),
    .A(\rgb_mixer.pwm0.count[0] ),
    .Y(_0216_));
 sg13g2_nand2_1 _0819_ (.Y(_0217_),
    .A(net86),
    .B(_0216_));
 sg13g2_nor2_1 _0820_ (.A(net205),
    .B(_0217_),
    .Y(_0025_));
 sg13g2_nor2_1 _0821_ (.A(_0142_),
    .B(_0216_),
    .Y(_0218_));
 sg13g2_a21oi_1 _0822_ (.A1(_0142_),
    .A2(_0216_),
    .Y(_0219_),
    .B1(net83));
 sg13g2_nor2b_1 _0823_ (.A(_0218_),
    .B_N(net280),
    .Y(_0026_));
 sg13g2_nor2_1 _0824_ (.A(net257),
    .B(_0218_),
    .Y(_0220_));
 sg13g2_and2_1 _0825_ (.A(net257),
    .B(_0218_),
    .X(_0221_));
 sg13g2_nor3_1 _0826_ (.A(net83),
    .B(net258),
    .C(_0221_),
    .Y(_0027_));
 sg13g2_o21ai_1 _0827_ (.B1(net86),
    .Y(_0222_),
    .A1(net249),
    .A2(_0221_));
 sg13g2_a21oi_1 _0828_ (.A1(net249),
    .A2(_0221_),
    .Y(_0028_),
    .B1(_0222_));
 sg13g2_a21oi_1 _0829_ (.A1(\rgb_mixer.pwm0.count[5] ),
    .A2(_0221_),
    .Y(_0223_),
    .B1(net220));
 sg13g2_nand3_1 _0830_ (.B(\rgb_mixer.pwm0.count[5] ),
    .C(_0221_),
    .A(net220),
    .Y(_0224_));
 sg13g2_nand2_1 _0831_ (.Y(_0225_),
    .A(net86),
    .B(_0224_));
 sg13g2_nor2_1 _0832_ (.A(net221),
    .B(_0225_),
    .Y(_0029_));
 sg13g2_o21ai_1 _0833_ (.B1(net86),
    .Y(_0226_),
    .A1(_0139_),
    .A2(_0224_));
 sg13g2_a21oi_1 _0834_ (.A1(_0139_),
    .A2(_0224_),
    .Y(_0030_),
    .B1(_0226_));
 sg13g2_nand2_1 _0835_ (.Y(_0227_),
    .A(net273),
    .B(_0132_));
 sg13g2_nor2_1 _0836_ (.A(\enc1[6] ),
    .B(_0133_),
    .Y(_0228_));
 sg13g2_nand2_1 _0837_ (.Y(_0229_),
    .A(_0120_),
    .B(\rgb_mixer.pwm1.count[6] ));
 sg13g2_nor2_1 _0838_ (.A(_0121_),
    .B(\rgb_mixer.pwm1.count[5] ),
    .Y(_0230_));
 sg13g2_a21oi_1 _0839_ (.A1(\enc1[6] ),
    .A2(_0133_),
    .Y(_0231_),
    .B1(_0230_));
 sg13g2_a22oi_1 _0840_ (.Y(_0232_),
    .B1(\rgb_mixer.pwm1.count[4] ),
    .B2(_0122_),
    .A2(\rgb_mixer.pwm1.count[5] ),
    .A1(_0121_));
 sg13g2_nand2b_1 _0841_ (.Y(_0233_),
    .B(\rgb_mixer.pwm1.count[3] ),
    .A_N(\enc1[3] ));
 sg13g2_nor2b_1 _0842_ (.A(\rgb_mixer.pwm1.count[2] ),
    .B_N(\enc1[2] ),
    .Y(_0234_));
 sg13g2_nand2_1 _0843_ (.Y(_0235_),
    .A(\enc1[3] ),
    .B(_0134_));
 sg13g2_o21ai_1 _0844_ (.B1(_0235_),
    .Y(_0236_),
    .A1(\enc1[2] ),
    .A2(_0135_));
 sg13g2_nand2b_1 _0845_ (.Y(_0237_),
    .B(\enc1[1] ),
    .A_N(\rgb_mixer.pwm1.count[1] ));
 sg13g2_nor2b_1 _0846_ (.A(\enc1[0] ),
    .B_N(\rgb_mixer.pwm1.count[0] ),
    .Y(_0238_));
 sg13g2_a21o_1 _0847_ (.A2(\rgb_mixer.pwm1.count[1] ),
    .A1(_0123_),
    .B1(_0238_),
    .X(_0239_));
 sg13g2_a21oi_1 _0848_ (.A1(_0237_),
    .A2(_0239_),
    .Y(_0240_),
    .B1(_0236_));
 sg13g2_o21ai_1 _0849_ (.B1(_0233_),
    .Y(_0241_),
    .A1(_0234_),
    .A2(_0240_));
 sg13g2_nand2b_1 _0850_ (.Y(_0242_),
    .B(\enc1[4] ),
    .A_N(\rgb_mixer.pwm1.count[4] ));
 sg13g2_nand3_1 _0851_ (.B(_0241_),
    .C(_0242_),
    .A(_0235_),
    .Y(_0243_));
 sg13g2_a221oi_1 _0852_ (.B2(_0243_),
    .C1(_0230_),
    .B1(_0232_),
    .A1(\enc1[6] ),
    .Y(_0244_),
    .A2(_0133_));
 sg13g2_o21ai_1 _0853_ (.B1(_0227_),
    .Y(_0245_),
    .A1(_0228_),
    .A2(_0244_));
 sg13g2_nor2_1 _0854_ (.A(_0124_),
    .B(\rgb_mixer.pwm1.count[0] ),
    .Y(_0246_));
 sg13g2_and4_1 _0855_ (.A(_0227_),
    .B(_0229_),
    .C(_0233_),
    .D(_0237_),
    .X(_0247_));
 sg13g2_nand2b_1 _0856_ (.Y(_0248_),
    .B(_0242_),
    .A_N(_0234_));
 sg13g2_nor4_1 _0857_ (.A(_0236_),
    .B(_0239_),
    .C(_0246_),
    .D(_0248_),
    .Y(_0249_));
 sg13g2_nand4_1 _0858_ (.B(_0232_),
    .C(_0247_),
    .A(_0231_),
    .Y(_0250_),
    .D(_0249_));
 sg13g2_nand2b_1 _0859_ (.Y(_0251_),
    .B(net236),
    .A_N(net273));
 sg13g2_and4_1 _0860_ (.A(net85),
    .B(_0245_),
    .C(_0250_),
    .D(_0251_),
    .X(_0031_));
 sg13g2_nand2_1 _0861_ (.Y(_0252_),
    .A(net229),
    .B(net96));
 sg13g2_inv_1 _0862_ (.Y(_0032_),
    .A(_0252_));
 sg13g2_nor2b_1 _0863_ (.A(net239),
    .B_N(net255),
    .Y(_0253_));
 sg13g2_nand2b_1 _0864_ (.Y(_0254_),
    .B(net220),
    .A_N(\enc0[6] ));
 sg13g2_a22oi_1 _0865_ (.Y(_0255_),
    .B1(_0141_),
    .B2(\enc0[5] ),
    .A2(_0140_),
    .A1(\enc0[6] ));
 sg13g2_nand2b_1 _0866_ (.Y(_0256_),
    .B(\rgb_mixer.pwm0.count[5] ),
    .A_N(\enc0[5] ));
 sg13g2_nand2b_1 _0867_ (.Y(_0257_),
    .B(\rgb_mixer.pwm0.count[4] ),
    .A_N(\enc0[4] ));
 sg13g2_nand2_1 _0868_ (.Y(_0258_),
    .A(_0256_),
    .B(_0257_));
 sg13g2_nor2b_1 _0869_ (.A(\enc0[1] ),
    .B_N(\rgb_mixer.pwm0.count[1] ),
    .Y(_0259_));
 sg13g2_a21o_1 _0870_ (.A2(\rgb_mixer.pwm0.count[0] ),
    .A1(_0119_),
    .B1(_0259_),
    .X(_0260_));
 sg13g2_nand2b_1 _0871_ (.Y(_0261_),
    .B(\enc0[2] ),
    .A_N(\rgb_mixer.pwm0.count[2] ));
 sg13g2_nand2b_1 _0872_ (.Y(_0262_),
    .B(\enc0[1] ),
    .A_N(\rgb_mixer.pwm0.count[1] ));
 sg13g2_and2_1 _0873_ (.A(_0261_),
    .B(_0262_),
    .X(_0263_));
 sg13g2_nor2_1 _0874_ (.A(\enc0[3] ),
    .B(_0142_),
    .Y(_0264_));
 sg13g2_nor2b_1 _0875_ (.A(\rgb_mixer.pwm0.count[3] ),
    .B_N(\enc0[3] ),
    .Y(_0265_));
 sg13g2_a21o_1 _0876_ (.A2(\rgb_mixer.pwm0.count[2] ),
    .A1(_0117_),
    .B1(_0265_),
    .X(_0266_));
 sg13g2_a221oi_1 _0877_ (.B2(_0261_),
    .C1(_0264_),
    .B1(_0266_),
    .A1(_0260_),
    .Y(_0267_),
    .A2(_0263_));
 sg13g2_nor2b_1 _0878_ (.A(\rgb_mixer.pwm0.count[4] ),
    .B_N(\enc0[4] ),
    .Y(_0268_));
 sg13g2_nor3_1 _0879_ (.A(_0265_),
    .B(_0267_),
    .C(_0268_),
    .Y(_0269_));
 sg13g2_o21ai_1 _0880_ (.B1(_0255_),
    .Y(_0270_),
    .A1(_0258_),
    .A2(_0269_));
 sg13g2_a21oi_1 _0881_ (.A1(_0254_),
    .A2(_0270_),
    .Y(_0271_),
    .B1(_0253_));
 sg13g2_nor2b_1 _0882_ (.A(_0253_),
    .B_N(_0254_),
    .Y(_0272_));
 sg13g2_nand4_1 _0883_ (.B(_0256_),
    .C(_0257_),
    .A(_0255_),
    .Y(_0273_),
    .D(_0272_));
 sg13g2_o21ai_1 _0884_ (.B1(_0263_),
    .Y(_0274_),
    .A1(_0119_),
    .A2(\rgb_mixer.pwm0.count[0] ));
 sg13g2_or4_1 _0885_ (.A(_0264_),
    .B(_0268_),
    .C(_0273_),
    .D(_0274_),
    .X(_0275_));
 sg13g2_nor3_1 _0886_ (.A(_0260_),
    .B(_0266_),
    .C(_0275_),
    .Y(_0276_));
 sg13g2_o21ai_1 _0887_ (.B1(net86),
    .Y(_0277_),
    .A1(net255),
    .A2(_0139_));
 sg13g2_nor3_1 _0888_ (.A(_0271_),
    .B(_0276_),
    .C(_0277_),
    .Y(_0033_));
 sg13g2_nor2_1 _0889_ (.A(\rgb_mixer.encoder2.old_b ),
    .B(\rgb_mixer.encoder2.old_a ),
    .Y(_0278_));
 sg13g2_inv_1 _0890_ (.Y(_0279_),
    .A(_0278_));
 sg13g2_and2_1 _0891_ (.A(\rgb_mixer.encoder2.old_b ),
    .B(\rgb_mixer.encoder2.old_a ),
    .X(_0280_));
 sg13g2_or2_1 _0892_ (.X(_0281_),
    .B(_0280_),
    .A(_0278_));
 sg13g2_nor2b_1 _0893_ (.A(\rgb_mixer.debounce2_a.debounced ),
    .B_N(\rgb_mixer.debounce2_b.debounced ),
    .Y(_0282_));
 sg13g2_nor2b_1 _0894_ (.A(\rgb_mixer.debounce2_b.debounced ),
    .B_N(\rgb_mixer.debounce2_a.debounced ),
    .Y(_0283_));
 sg13g2_nand2b_1 _0895_ (.Y(_0284_),
    .B(\rgb_mixer.debounce2_a.debounced ),
    .A_N(\rgb_mixer.debounce2_b.debounced ));
 sg13g2_nand2b_1 _0896_ (.Y(_0285_),
    .B(_0284_),
    .A_N(_0282_));
 sg13g2_and2_1 _0897_ (.A(_0281_),
    .B(_0285_),
    .X(_0286_));
 sg13g2_nand2_2 _0898_ (.Y(_0287_),
    .A(_0281_),
    .B(_0285_));
 sg13g2_o21ai_1 _0899_ (.B1(net89),
    .Y(_0288_),
    .A1(net247),
    .A2(_0287_));
 sg13g2_a21oi_1 _0900_ (.A1(_0129_),
    .A2(_0287_),
    .Y(_0034_),
    .B1(_0288_));
 sg13g2_nor2_1 _0901_ (.A(_0280_),
    .B(_0282_),
    .Y(_0289_));
 sg13g2_a21oi_2 _0902_ (.B1(_0289_),
    .Y(_0290_),
    .A2(_0284_),
    .A1(_0279_));
 sg13g2_a22oi_1 _0903_ (.Y(_0291_),
    .B1(_0283_),
    .B2(_0280_),
    .A2(_0282_),
    .A1(_0278_));
 sg13g2_nand2_1 _0904_ (.Y(_0292_),
    .A(_0128_),
    .B(_0291_));
 sg13g2_xnor2_1 _0905_ (.Y(_0293_),
    .A(_0128_),
    .B(net82));
 sg13g2_nor3_1 _0906_ (.A(net247),
    .B(_0287_),
    .C(_0293_),
    .Y(_0294_));
 sg13g2_and3_1 _0907_ (.X(_0295_),
    .A(net247),
    .B(net79),
    .C(_0293_));
 sg13g2_o21ai_1 _0908_ (.B1(net89),
    .Y(_0296_),
    .A1(net272),
    .A2(net79));
 sg13g2_nor3_1 _0909_ (.A(_0294_),
    .B(_0295_),
    .C(_0296_),
    .Y(_0035_));
 sg13g2_xnor2_1 _0910_ (.Y(_0297_),
    .A(\enc2[2] ),
    .B(_0291_));
 sg13g2_o21ai_1 _0911_ (.B1(_0129_),
    .Y(_0298_),
    .A1(_0128_),
    .A2(net82));
 sg13g2_nand3_1 _0912_ (.B(_0297_),
    .C(_0298_),
    .A(_0292_),
    .Y(_0299_));
 sg13g2_a21o_1 _0913_ (.A2(_0298_),
    .A1(_0292_),
    .B1(_0297_),
    .X(_0300_));
 sg13g2_a21oi_1 _0914_ (.A1(_0299_),
    .A2(_0300_),
    .Y(_0301_),
    .B1(_0287_));
 sg13g2_o21ai_1 _0915_ (.B1(net92),
    .Y(_0302_),
    .A1(net289),
    .A2(_0286_));
 sg13g2_nor2_1 _0916_ (.A(_0301_),
    .B(_0302_),
    .Y(_0036_));
 sg13g2_xnor2_1 _0917_ (.Y(_0303_),
    .A(\enc2[3] ),
    .B(net82));
 sg13g2_o21ai_1 _0918_ (.B1(_0299_),
    .Y(_0304_),
    .A1(_0127_),
    .A2(net82));
 sg13g2_xnor2_1 _0919_ (.Y(_0305_),
    .A(_0303_),
    .B(_0304_));
 sg13g2_o21ai_1 _0920_ (.B1(net92),
    .Y(_0306_),
    .A1(net290),
    .A2(_0286_));
 sg13g2_a21oi_1 _0921_ (.A1(_0286_),
    .A2(_0305_),
    .Y(_0037_),
    .B1(_0306_));
 sg13g2_nand4_1 _0922_ (.B(_0297_),
    .C(_0298_),
    .A(_0292_),
    .Y(_0307_),
    .D(_0303_));
 sg13g2_o21ai_1 _0923_ (.B1(_0290_),
    .Y(_0308_),
    .A1(\enc2[3] ),
    .A2(\enc2[2] ));
 sg13g2_nand2_1 _0924_ (.Y(_0309_),
    .A(_0307_),
    .B(_0308_));
 sg13g2_nor2_1 _0925_ (.A(_0126_),
    .B(net82),
    .Y(_0310_));
 sg13g2_xnor2_1 _0926_ (.Y(_0311_),
    .A(\enc2[4] ),
    .B(net82));
 sg13g2_xnor2_1 _0927_ (.Y(_0312_),
    .A(_0309_),
    .B(_0311_));
 sg13g2_o21ai_1 _0928_ (.B1(net89),
    .Y(_0313_),
    .A1(net298),
    .A2(net79));
 sg13g2_a21oi_1 _0929_ (.A1(net79),
    .A2(_0312_),
    .Y(_0038_),
    .B1(_0313_));
 sg13g2_xnor2_1 _0930_ (.Y(_0314_),
    .A(\enc2[5] ),
    .B(net82));
 sg13g2_a21oi_1 _0931_ (.A1(_0309_),
    .A2(_0311_),
    .Y(_0315_),
    .B1(_0310_));
 sg13g2_or2_1 _0932_ (.X(_0316_),
    .B(_0315_),
    .A(_0314_));
 sg13g2_a21oi_1 _0933_ (.A1(_0314_),
    .A2(_0315_),
    .Y(_0317_),
    .B1(_0287_));
 sg13g2_a221oi_1 _0934_ (.B2(_0317_),
    .C1(net84),
    .B1(_0316_),
    .A1(_0125_),
    .Y(_0039_),
    .A2(_0287_));
 sg13g2_nor2_1 _0935_ (.A(\enc2[6] ),
    .B(_0290_),
    .Y(_0318_));
 sg13g2_nand2_1 _0936_ (.Y(_0319_),
    .A(\enc2[6] ),
    .B(_0290_));
 sg13g2_nor2b_1 _0937_ (.A(_0318_),
    .B_N(_0319_),
    .Y(_0320_));
 sg13g2_and2_1 _0938_ (.A(_0311_),
    .B(_0314_),
    .X(_0321_));
 sg13g2_a221oi_1 _0939_ (.B2(_0321_),
    .C1(_0310_),
    .B1(_0309_),
    .A1(\enc2[5] ),
    .Y(_0322_),
    .A2(_0290_));
 sg13g2_xor2_1 _0940_ (.B(_0322_),
    .A(_0320_),
    .X(_0323_));
 sg13g2_o21ai_1 _0941_ (.B1(net93),
    .Y(_0324_),
    .A1(net295),
    .A2(net79));
 sg13g2_a21oi_1 _0942_ (.A1(net79),
    .A2(_0323_),
    .Y(_0040_),
    .B1(_0324_));
 sg13g2_o21ai_1 _0943_ (.B1(_0319_),
    .Y(_0325_),
    .A1(_0318_),
    .A2(_0322_));
 sg13g2_xnor2_1 _0944_ (.Y(_0326_),
    .A(\enc2[7] ),
    .B(net82));
 sg13g2_xnor2_1 _0945_ (.Y(_0327_),
    .A(_0325_),
    .B(_0326_));
 sg13g2_o21ai_1 _0946_ (.B1(net89),
    .Y(_0328_),
    .A1(net275),
    .A2(net79));
 sg13g2_a21oi_1 _0947_ (.A1(net79),
    .A2(_0327_),
    .Y(_0041_),
    .B1(_0328_));
 sg13g2_nand2_1 _0948_ (.Y(_0329_),
    .A(net211),
    .B(net92));
 sg13g2_inv_1 _0949_ (.Y(_0042_),
    .A(_0329_));
 sg13g2_nand2_1 _0950_ (.Y(_0330_),
    .A(net226),
    .B(net96));
 sg13g2_inv_1 _0951_ (.Y(_0043_),
    .A(_0330_));
 sg13g2_nor2_1 _0952_ (.A(\rgb_mixer.encoder1.old_b ),
    .B(\rgb_mixer.encoder1.old_a ),
    .Y(_0331_));
 sg13g2_inv_1 _0953_ (.Y(_0332_),
    .A(_0331_));
 sg13g2_and2_1 _0954_ (.A(\rgb_mixer.encoder1.old_b ),
    .B(\rgb_mixer.encoder1.old_a ),
    .X(_0333_));
 sg13g2_or2_1 _0955_ (.X(_0334_),
    .B(_0333_),
    .A(_0331_));
 sg13g2_nor2b_1 _0956_ (.A(\rgb_mixer.debounce1_a.debounced ),
    .B_N(\rgb_mixer.debounce1_b.debounced ),
    .Y(_0335_));
 sg13g2_nor2b_1 _0957_ (.A(\rgb_mixer.debounce1_b.debounced ),
    .B_N(\rgb_mixer.debounce1_a.debounced ),
    .Y(_0336_));
 sg13g2_nand2b_1 _0958_ (.Y(_0337_),
    .B(\rgb_mixer.debounce1_a.debounced ),
    .A_N(\rgb_mixer.debounce1_b.debounced ));
 sg13g2_nand2b_1 _0959_ (.Y(_0338_),
    .B(_0337_),
    .A_N(_0335_));
 sg13g2_and2_1 _0960_ (.A(_0334_),
    .B(_0338_),
    .X(_0339_));
 sg13g2_nand2_2 _0961_ (.Y(_0340_),
    .A(_0334_),
    .B(_0338_));
 sg13g2_o21ai_1 _0962_ (.B1(net89),
    .Y(_0341_),
    .A1(net234),
    .A2(_0340_));
 sg13g2_a21oi_1 _0963_ (.A1(_0124_),
    .A2(_0340_),
    .Y(_0044_),
    .B1(_0341_));
 sg13g2_nor2_1 _0964_ (.A(_0333_),
    .B(_0335_),
    .Y(_0342_));
 sg13g2_a21oi_2 _0965_ (.B1(_0342_),
    .Y(_0343_),
    .A2(_0337_),
    .A1(_0332_));
 sg13g2_a22oi_1 _0966_ (.Y(_0344_),
    .B1(_0336_),
    .B2(_0333_),
    .A2(_0335_),
    .A1(_0331_));
 sg13g2_nand2_1 _0967_ (.Y(_0345_),
    .A(_0123_),
    .B(net81));
 sg13g2_xnor2_1 _0968_ (.Y(_0346_),
    .A(_0123_),
    .B(net81));
 sg13g2_nor3_1 _0969_ (.A(net234),
    .B(_0340_),
    .C(_0346_),
    .Y(_0347_));
 sg13g2_and3_1 _0970_ (.X(_0348_),
    .A(net234),
    .B(net78),
    .C(_0346_));
 sg13g2_o21ai_1 _0971_ (.B1(net89),
    .Y(_0349_),
    .A1(net262),
    .A2(net78));
 sg13g2_nor3_1 _0972_ (.A(_0347_),
    .B(_0348_),
    .C(_0349_),
    .Y(_0045_));
 sg13g2_xnor2_1 _0973_ (.Y(_0350_),
    .A(\enc1[2] ),
    .B(net81));
 sg13g2_o21ai_1 _0974_ (.B1(_0124_),
    .Y(_0351_),
    .A1(_0123_),
    .A2(net81));
 sg13g2_and3_1 _0975_ (.X(_0352_),
    .A(_0345_),
    .B(_0350_),
    .C(_0351_));
 sg13g2_a21oi_1 _0976_ (.A1(_0345_),
    .A2(_0351_),
    .Y(_0353_),
    .B1(_0350_));
 sg13g2_o21ai_1 _0977_ (.B1(net78),
    .Y(_0354_),
    .A1(_0352_),
    .A2(_0353_));
 sg13g2_o21ai_1 _0978_ (.B1(_0354_),
    .Y(_0355_),
    .A1(net300),
    .A2(net78));
 sg13g2_nor2_1 _0979_ (.A(net83),
    .B(_0355_),
    .Y(_0046_));
 sg13g2_xnor2_1 _0980_ (.Y(_0356_),
    .A(\enc1[3] ),
    .B(net81));
 sg13g2_a21oi_1 _0981_ (.A1(\enc1[2] ),
    .A2(_0343_),
    .Y(_0357_),
    .B1(_0352_));
 sg13g2_o21ai_1 _0982_ (.B1(net78),
    .Y(_0358_),
    .A1(_0356_),
    .A2(_0357_));
 sg13g2_a21oi_1 _0983_ (.A1(_0356_),
    .A2(_0357_),
    .Y(_0359_),
    .B1(_0358_));
 sg13g2_o21ai_1 _0984_ (.B1(net90),
    .Y(_0360_),
    .A1(net294),
    .A2(net78));
 sg13g2_nor2_1 _0985_ (.A(_0359_),
    .B(_0360_),
    .Y(_0047_));
 sg13g2_nand4_1 _0986_ (.B(_0350_),
    .C(_0351_),
    .A(_0345_),
    .Y(_0361_),
    .D(_0356_));
 sg13g2_o21ai_1 _0987_ (.B1(_0343_),
    .Y(_0362_),
    .A1(\enc1[3] ),
    .A2(\enc1[2] ));
 sg13g2_nand2_1 _0988_ (.Y(_0363_),
    .A(_0361_),
    .B(_0362_));
 sg13g2_nor2_1 _0989_ (.A(_0122_),
    .B(net81),
    .Y(_0364_));
 sg13g2_xnor2_1 _0990_ (.Y(_0365_),
    .A(\enc1[4] ),
    .B(net81));
 sg13g2_xnor2_1 _0991_ (.Y(_0366_),
    .A(_0363_),
    .B(_0365_));
 sg13g2_o21ai_1 _0992_ (.B1(net90),
    .Y(_0367_),
    .A1(net288),
    .A2(_0339_));
 sg13g2_a21oi_1 _0993_ (.A1(net78),
    .A2(_0366_),
    .Y(_0048_),
    .B1(_0367_));
 sg13g2_xnor2_1 _0994_ (.Y(_0368_),
    .A(\enc1[5] ),
    .B(net81));
 sg13g2_a21oi_1 _0995_ (.A1(_0363_),
    .A2(_0365_),
    .Y(_0369_),
    .B1(_0364_));
 sg13g2_or2_1 _0996_ (.X(_0370_),
    .B(_0369_),
    .A(_0368_));
 sg13g2_a21oi_1 _0997_ (.A1(_0368_),
    .A2(_0369_),
    .Y(_0371_),
    .B1(_0340_));
 sg13g2_a221oi_1 _0998_ (.B2(_0371_),
    .C1(net83),
    .B1(_0370_),
    .A1(_0121_),
    .Y(_0049_),
    .A2(_0340_));
 sg13g2_nand2_1 _0999_ (.Y(_0372_),
    .A(\enc1[6] ),
    .B(_0343_));
 sg13g2_xnor2_1 _1000_ (.Y(_0373_),
    .A(\enc1[6] ),
    .B(_0344_));
 sg13g2_nand2_1 _1001_ (.Y(_0374_),
    .A(_0365_),
    .B(_0368_));
 sg13g2_a21oi_1 _1002_ (.A1(_0361_),
    .A2(_0362_),
    .Y(_0375_),
    .B1(_0374_));
 sg13g2_a21oi_1 _1003_ (.A1(_0121_),
    .A2(_0122_),
    .Y(_0376_),
    .B1(_0344_));
 sg13g2_nor3_1 _1004_ (.A(_0373_),
    .B(_0375_),
    .C(_0376_),
    .Y(_0377_));
 sg13g2_o21ai_1 _1005_ (.B1(_0373_),
    .Y(_0378_),
    .A1(_0375_),
    .A2(_0376_));
 sg13g2_nor2b_1 _1006_ (.A(_0377_),
    .B_N(_0378_),
    .Y(_0379_));
 sg13g2_o21ai_1 _1007_ (.B1(net85),
    .Y(_0380_),
    .A1(_0340_),
    .A2(_0379_));
 sg13g2_a21oi_1 _1008_ (.A1(_0120_),
    .A2(_0340_),
    .Y(_0050_),
    .B1(_0380_));
 sg13g2_xnor2_1 _1009_ (.Y(_0381_),
    .A(net296),
    .B(_0344_));
 sg13g2_a21oi_1 _1010_ (.A1(_0372_),
    .A2(_0378_),
    .Y(_0382_),
    .B1(_0381_));
 sg13g2_nand3_1 _1011_ (.B(_0378_),
    .C(_0381_),
    .A(_0372_),
    .Y(_0383_));
 sg13g2_nor2_1 _1012_ (.A(_0340_),
    .B(_0382_),
    .Y(_0384_));
 sg13g2_o21ai_1 _1013_ (.B1(net85),
    .Y(_0385_),
    .A1(net273),
    .A2(net78));
 sg13g2_a21oi_1 _1014_ (.A1(net297),
    .A2(_0384_),
    .Y(_0051_),
    .B1(_0385_));
 sg13g2_and2_1 _1015_ (.A(net203),
    .B(net88),
    .X(_0052_));
 sg13g2_nand2_2 _1016_ (.Y(_0386_),
    .A(net214),
    .B(net92));
 sg13g2_inv_1 _1017_ (.Y(_0053_),
    .A(_0386_));
 sg13g2_nor2_1 _1018_ (.A(\rgb_mixer.encoder0.old_b ),
    .B(\rgb_mixer.encoder0.old_a ),
    .Y(_0387_));
 sg13g2_inv_1 _1019_ (.Y(_0388_),
    .A(_0387_));
 sg13g2_and2_1 _1020_ (.A(\rgb_mixer.encoder0.old_b ),
    .B(\rgb_mixer.encoder0.old_a ),
    .X(_0389_));
 sg13g2_or2_1 _1021_ (.X(_0390_),
    .B(_0389_),
    .A(_0387_));
 sg13g2_nor2b_1 _1022_ (.A(\rgb_mixer.debounce0_a.debounced ),
    .B_N(\rgb_mixer.debounce0_b.debounced ),
    .Y(_0391_));
 sg13g2_nor2b_1 _1023_ (.A(\rgb_mixer.debounce0_b.debounced ),
    .B_N(\rgb_mixer.debounce0_a.debounced ),
    .Y(_0392_));
 sg13g2_nand2b_1 _1024_ (.Y(_0393_),
    .B(\rgb_mixer.debounce0_a.debounced ),
    .A_N(\rgb_mixer.debounce0_b.debounced ));
 sg13g2_nand2b_1 _1025_ (.Y(_0394_),
    .B(_0393_),
    .A_N(_0391_));
 sg13g2_and2_1 _1026_ (.A(_0390_),
    .B(_0394_),
    .X(_0395_));
 sg13g2_nand2_2 _1027_ (.Y(_0396_),
    .A(_0390_),
    .B(_0394_));
 sg13g2_o21ai_1 _1028_ (.B1(net87),
    .Y(_0397_),
    .A1(net245),
    .A2(_0396_));
 sg13g2_a21oi_1 _1029_ (.A1(_0119_),
    .A2(_0396_),
    .Y(_0054_),
    .B1(_0397_));
 sg13g2_nor2_1 _1030_ (.A(_0389_),
    .B(_0391_),
    .Y(_0398_));
 sg13g2_a21oi_2 _1031_ (.B1(_0398_),
    .Y(_0399_),
    .A2(_0393_),
    .A1(_0388_));
 sg13g2_a22oi_1 _1032_ (.Y(_0400_),
    .B1(_0392_),
    .B2(_0389_),
    .A2(_0391_),
    .A1(_0387_));
 sg13g2_nand2_1 _1033_ (.Y(_0401_),
    .A(_0118_),
    .B(net80));
 sg13g2_xnor2_1 _1034_ (.Y(_0402_),
    .A(_0118_),
    .B(net80));
 sg13g2_nor3_1 _1035_ (.A(net245),
    .B(_0396_),
    .C(_0402_),
    .Y(_0403_));
 sg13g2_and3_1 _1036_ (.X(_0404_),
    .A(net245),
    .B(net76),
    .C(_0402_));
 sg13g2_o21ai_1 _1037_ (.B1(net88),
    .Y(_0405_),
    .A1(net269),
    .A2(net76));
 sg13g2_nor3_1 _1038_ (.A(_0403_),
    .B(_0404_),
    .C(_0405_),
    .Y(_0055_));
 sg13g2_xnor2_1 _1039_ (.Y(_0406_),
    .A(\enc0[2] ),
    .B(net80));
 sg13g2_o21ai_1 _1040_ (.B1(_0119_),
    .Y(_0407_),
    .A1(_0118_),
    .A2(net80));
 sg13g2_nand3_1 _1041_ (.B(_0406_),
    .C(_0407_),
    .A(_0401_),
    .Y(_0408_));
 sg13g2_a21o_1 _1042_ (.A2(_0407_),
    .A1(_0401_),
    .B1(_0406_),
    .X(_0409_));
 sg13g2_a21oi_1 _1043_ (.A1(_0408_),
    .A2(_0409_),
    .Y(_0410_),
    .B1(_0396_));
 sg13g2_o21ai_1 _1044_ (.B1(net87),
    .Y(_0411_),
    .A1(net293),
    .A2(net76));
 sg13g2_nor2_1 _1045_ (.A(_0410_),
    .B(_0411_),
    .Y(_0056_));
 sg13g2_xnor2_1 _1046_ (.Y(_0412_),
    .A(\enc0[3] ),
    .B(net80));
 sg13g2_inv_1 _1047_ (.Y(_0413_),
    .A(_0412_));
 sg13g2_o21ai_1 _1048_ (.B1(_0408_),
    .Y(_0414_),
    .A1(_0117_),
    .A2(net80));
 sg13g2_xnor2_1 _1049_ (.Y(_0415_),
    .A(_0412_),
    .B(_0414_));
 sg13g2_o21ai_1 _1050_ (.B1(net87),
    .Y(_0416_),
    .A1(net292),
    .A2(net76));
 sg13g2_a21oi_1 _1051_ (.A1(net76),
    .A2(_0415_),
    .Y(_0057_),
    .B1(_0416_));
 sg13g2_o21ai_1 _1052_ (.B1(_0399_),
    .Y(_0417_),
    .A1(\enc0[3] ),
    .A2(\enc0[2] ));
 sg13g2_o21ai_1 _1053_ (.B1(_0417_),
    .Y(_0418_),
    .A1(_0408_),
    .A2(_0413_));
 sg13g2_and2_1 _1054_ (.A(\enc0[4] ),
    .B(_0399_),
    .X(_0419_));
 sg13g2_xnor2_1 _1055_ (.Y(_0420_),
    .A(\enc0[4] ),
    .B(_0400_));
 sg13g2_xnor2_1 _1056_ (.Y(_0421_),
    .A(_0418_),
    .B(_0420_));
 sg13g2_o21ai_1 _1057_ (.B1(net87),
    .Y(_0422_),
    .A1(net278),
    .A2(net77));
 sg13g2_a21oi_1 _1058_ (.A1(net77),
    .A2(_0421_),
    .Y(_0058_),
    .B1(_0422_));
 sg13g2_xnor2_1 _1059_ (.Y(_0423_),
    .A(\enc0[5] ),
    .B(net80));
 sg13g2_a21oi_1 _1060_ (.A1(_0418_),
    .A2(_0420_),
    .Y(_0424_),
    .B1(_0419_));
 sg13g2_nand2_1 _1061_ (.Y(_0425_),
    .A(_0423_),
    .B(_0424_));
 sg13g2_nor2_1 _1062_ (.A(_0423_),
    .B(_0424_),
    .Y(_0426_));
 sg13g2_nor2_1 _1063_ (.A(_0396_),
    .B(_0426_),
    .Y(_0427_));
 sg13g2_o21ai_1 _1064_ (.B1(net87),
    .Y(_0428_),
    .A1(net286),
    .A2(net77));
 sg13g2_a21oi_1 _1065_ (.A1(_0425_),
    .A2(_0427_),
    .Y(_0059_),
    .B1(_0428_));
 sg13g2_nor2_1 _1066_ (.A(\enc0[6] ),
    .B(_0399_),
    .Y(_0429_));
 sg13g2_nand2_1 _1067_ (.Y(_0430_),
    .A(\enc0[6] ),
    .B(_0399_));
 sg13g2_nand2b_1 _1068_ (.Y(_0431_),
    .B(_0430_),
    .A_N(_0429_));
 sg13g2_and2_1 _1069_ (.A(_0420_),
    .B(_0423_),
    .X(_0432_));
 sg13g2_a221oi_1 _1070_ (.B2(_0432_),
    .C1(_0419_),
    .B1(_0418_),
    .A1(\enc0[5] ),
    .Y(_0433_),
    .A2(_0399_));
 sg13g2_xnor2_1 _1071_ (.Y(_0434_),
    .A(_0431_),
    .B(_0433_));
 sg13g2_o21ai_1 _1072_ (.B1(net87),
    .Y(_0435_),
    .A1(net274),
    .A2(net77));
 sg13g2_a21oi_1 _1073_ (.A1(net76),
    .A2(_0434_),
    .Y(_0060_),
    .B1(_0435_));
 sg13g2_o21ai_1 _1074_ (.B1(_0430_),
    .Y(_0436_),
    .A1(_0429_),
    .A2(_0433_));
 sg13g2_xnor2_1 _1075_ (.Y(_0437_),
    .A(net277),
    .B(net80));
 sg13g2_xnor2_1 _1076_ (.Y(_0438_),
    .A(_0436_),
    .B(_0437_));
 sg13g2_o21ai_1 _1077_ (.B1(net87),
    .Y(_0439_),
    .A1(net255),
    .A2(net76));
 sg13g2_a21oi_1 _1078_ (.A1(net76),
    .A2(_0438_),
    .Y(_0061_),
    .B1(_0439_));
 sg13g2_and2_1 _1079_ (.A(net99),
    .B(net6),
    .X(_0062_));
 sg13g2_and2_1 _1080_ (.A(net185),
    .B(net95),
    .X(_0063_));
 sg13g2_and2_1 _1081_ (.A(net178),
    .B(net95),
    .X(_0064_));
 sg13g2_and2_1 _1082_ (.A(net173),
    .B(net95),
    .X(_0065_));
 sg13g2_and2_1 _1083_ (.A(net163),
    .B(net95),
    .X(_0066_));
 sg13g2_and2_1 _1084_ (.A(net172),
    .B(net95),
    .X(_0067_));
 sg13g2_and2_1 _1085_ (.A(net187),
    .B(net95),
    .X(_0068_));
 sg13g2_and2_1 _1086_ (.A(net194),
    .B(net95),
    .X(_0069_));
 sg13g2_and2_1 _1087_ (.A(net238),
    .B(net94),
    .X(_0070_));
 sg13g2_nand3_1 _1088_ (.B(net173),
    .C(_0064_),
    .A(net185),
    .Y(_0440_));
 sg13g2_nand4_1 _1089_ (.B(net187),
    .C(\rgb_mixer.debounce2_b.button_hist[7] ),
    .A(net172),
    .Y(_0441_),
    .D(net194));
 sg13g2_o21ai_1 _1090_ (.B1(_0252_),
    .Y(_0442_),
    .A1(_0440_),
    .A2(_0441_));
 sg13g2_nor3_1 _1091_ (.A(net187),
    .B(\rgb_mixer.debounce2_b.button_hist[7] ),
    .C(net194),
    .Y(_0443_));
 sg13g2_nor4_1 _1092_ (.A(net185),
    .B(net178),
    .C(net173),
    .D(net172),
    .Y(_0444_));
 sg13g2_a21oi_1 _1093_ (.A1(_0443_),
    .A2(_0444_),
    .Y(_0445_),
    .B1(_0252_));
 sg13g2_a21o_1 _1094_ (.A2(_0442_),
    .A1(net163),
    .B1(net230),
    .X(_0071_));
 sg13g2_and2_1 _1095_ (.A(net99),
    .B(net5),
    .X(_0072_));
 sg13g2_and2_1 _1096_ (.A(net175),
    .B(net97),
    .X(_0073_));
 sg13g2_and2_1 _1097_ (.A(net174),
    .B(net97),
    .X(_0074_));
 sg13g2_and2_1 _1098_ (.A(net177),
    .B(net97),
    .X(_0075_));
 sg13g2_and2_1 _1099_ (.A(net198),
    .B(net97),
    .X(_0076_));
 sg13g2_and2_1 _1100_ (.A(net171),
    .B(net95),
    .X(_0077_));
 sg13g2_and2_1 _1101_ (.A(net197),
    .B(net96),
    .X(_0078_));
 sg13g2_and2_1 _1102_ (.A(net182),
    .B(net100),
    .X(_0079_));
 sg13g2_nor4_1 _1103_ (.A(net174),
    .B(net175),
    .C(net198),
    .D(net177),
    .Y(_0446_));
 sg13g2_nand4_1 _1104_ (.B(net177),
    .C(\rgb_mixer.debounce2_a.button_hist[7] ),
    .A(net198),
    .Y(_0447_),
    .D(net182));
 sg13g2_nand3_1 _1105_ (.B(net175),
    .C(_0078_),
    .A(net174),
    .Y(_0448_));
 sg13g2_o21ai_1 _1106_ (.B1(_0330_),
    .Y(_0449_),
    .A1(_0447_),
    .A2(_0448_));
 sg13g2_nor3_1 _1107_ (.A(net197),
    .B(\rgb_mixer.debounce2_a.button_hist[7] ),
    .C(net182),
    .Y(_0450_));
 sg13g2_a21oi_1 _1108_ (.A1(_0446_),
    .A2(_0450_),
    .Y(_0451_),
    .B1(_0330_));
 sg13g2_a21o_1 _1109_ (.A2(_0449_),
    .A1(net171),
    .B1(net227),
    .X(_0080_));
 sg13g2_and2_1 _1110_ (.A(net99),
    .B(net4),
    .X(_0081_));
 sg13g2_and2_1 _1111_ (.A(net191),
    .B(net92),
    .X(_0082_));
 sg13g2_and2_1 _1112_ (.A(net176),
    .B(net99),
    .X(_0083_));
 sg13g2_and2_1 _1113_ (.A(net192),
    .B(net99),
    .X(_0084_));
 sg13g2_and2_1 _1114_ (.A(net166),
    .B(net93),
    .X(_0085_));
 sg13g2_and2_1 _1115_ (.A(net164),
    .B(net92),
    .X(_0086_));
 sg13g2_and2_1 _1116_ (.A(net199),
    .B(net99),
    .X(_0087_));
 sg13g2_and2_1 _1117_ (.A(net195),
    .B(net99),
    .X(_0088_));
 sg13g2_nor4_1 _1118_ (.A(net176),
    .B(net191),
    .C(net166),
    .D(net192),
    .Y(_0452_));
 sg13g2_nand4_1 _1119_ (.B(net192),
    .C(\rgb_mixer.debounce1_b.button_hist[7] ),
    .A(net166),
    .Y(_0453_),
    .D(net195));
 sg13g2_nand3_1 _1120_ (.B(net191),
    .C(_0087_),
    .A(net176),
    .Y(_0454_));
 sg13g2_o21ai_1 _1121_ (.B1(_0329_),
    .Y(_0455_),
    .A1(_0453_),
    .A2(_0454_));
 sg13g2_nor3_1 _1122_ (.A(net199),
    .B(\rgb_mixer.debounce1_b.button_hist[7] ),
    .C(net195),
    .Y(_0456_));
 sg13g2_a21oi_1 _1123_ (.A1(_0452_),
    .A2(_0456_),
    .Y(_0457_),
    .B1(_0329_));
 sg13g2_a21o_1 _1124_ (.A2(_0455_),
    .A1(net164),
    .B1(net212),
    .X(_0089_));
 sg13g2_and2_1 _1125_ (.A(net98),
    .B(net3),
    .X(_0090_));
 sg13g2_and2_1 _1126_ (.A(net167),
    .B(net97),
    .X(_0091_));
 sg13g2_and2_1 _1127_ (.A(net179),
    .B(net97),
    .X(_0092_));
 sg13g2_and2_1 _1128_ (.A(net190),
    .B(net97),
    .X(_0093_));
 sg13g2_and2_1 _1129_ (.A(net202),
    .B(net98),
    .X(_0094_));
 sg13g2_and2_1 _1130_ (.A(net161),
    .B(net98),
    .X(_0095_));
 sg13g2_and2_1 _1131_ (.A(net168),
    .B(net98),
    .X(_0096_));
 sg13g2_and2_1 _1132_ (.A(net200),
    .B(net97),
    .X(_0097_));
 sg13g2_nor4_1 _1133_ (.A(net179),
    .B(net167),
    .C(net202),
    .D(net190),
    .Y(_0458_));
 sg13g2_nand4_1 _1134_ (.B(net190),
    .C(\rgb_mixer.debounce1_a.button_hist[7] ),
    .A(net202),
    .Y(_0459_),
    .D(net200));
 sg13g2_nand3_1 _1135_ (.B(net167),
    .C(_0096_),
    .A(net179),
    .Y(_0460_));
 sg13g2_o21ai_1 _1136_ (.B1(_0386_),
    .Y(_0461_),
    .A1(_0459_),
    .A2(_0460_));
 sg13g2_nor3_1 _1137_ (.A(net168),
    .B(\rgb_mixer.debounce1_a.button_hist[7] ),
    .C(net200),
    .Y(_0462_));
 sg13g2_a21oi_1 _1138_ (.A1(_0458_),
    .A2(_0462_),
    .Y(_0463_),
    .B1(_0386_));
 sg13g2_a21o_1 _1139_ (.A2(_0461_),
    .A1(net161),
    .B1(net215),
    .X(_0098_));
 sg13g2_and2_1 _1140_ (.A(net92),
    .B(net2),
    .X(_0099_));
 sg13g2_and2_1 _1141_ (.A(net183),
    .B(net91),
    .X(_0100_));
 sg13g2_and2_1 _1142_ (.A(net184),
    .B(net91),
    .X(_0101_));
 sg13g2_and2_1 _1143_ (.A(net165),
    .B(net91),
    .X(_0102_));
 sg13g2_and2_1 _1144_ (.A(net170),
    .B(net91),
    .X(_0103_));
 sg13g2_and2_1 _1145_ (.A(net180),
    .B(net88),
    .X(_0104_));
 sg13g2_nor2_1 _1146_ (.A(_0131_),
    .B(net83),
    .Y(_0105_));
 sg13g2_and2_1 _1147_ (.A(net186),
    .B(net87),
    .X(_0106_));
 sg13g2_or4_1 _1148_ (.A(net184),
    .B(net183),
    .C(net170),
    .D(net165),
    .X(_0464_));
 sg13g2_nand4_1 _1149_ (.B(net183),
    .C(net165),
    .A(net184),
    .Y(_0465_),
    .D(net186));
 sg13g2_nand3_1 _1150_ (.B(net207),
    .C(_0103_),
    .A(net180),
    .Y(_0466_));
 sg13g2_nor3_1 _1151_ (.A(_0131_),
    .B(_0465_),
    .C(_0466_),
    .Y(_0467_));
 sg13g2_nor2_1 _1152_ (.A(_0052_),
    .B(_0467_),
    .Y(_0468_));
 sg13g2_nor4_1 _1153_ (.A(net180),
    .B(net207),
    .C(net186),
    .D(_0464_),
    .Y(_0469_));
 sg13g2_a21oi_1 _1154_ (.A1(_0131_),
    .A2(_0469_),
    .Y(_0107_),
    .B1(_0468_));
 sg13g2_and2_1 _1155_ (.A(net99),
    .B(net1),
    .X(_0108_));
 sg13g2_and2_1 _1156_ (.A(net181),
    .B(net96),
    .X(_0109_));
 sg13g2_and2_1 _1157_ (.A(net162),
    .B(net96),
    .X(_0110_));
 sg13g2_and2_1 _1158_ (.A(net189),
    .B(net96),
    .X(_0111_));
 sg13g2_and2_1 _1159_ (.A(net169),
    .B(net96),
    .X(_0112_));
 sg13g2_and2_1 _1160_ (.A(net196),
    .B(net94),
    .X(_0113_));
 sg13g2_nor2_1 _1161_ (.A(_0130_),
    .B(net84),
    .Y(_0114_));
 sg13g2_and2_1 _1162_ (.A(net188),
    .B(net94),
    .X(_0115_));
 sg13g2_or4_1 _1163_ (.A(net162),
    .B(net181),
    .C(net169),
    .D(net189),
    .X(_0470_));
 sg13g2_nand4_1 _1164_ (.B(net196),
    .C(net232),
    .A(net189),
    .Y(_0471_),
    .D(net188));
 sg13g2_nand3_1 _1165_ (.B(net169),
    .C(_0109_),
    .A(net162),
    .Y(_0472_));
 sg13g2_nor3_1 _1166_ (.A(_0130_),
    .B(_0471_),
    .C(_0472_),
    .Y(_0473_));
 sg13g2_nor2_1 _1167_ (.A(_0070_),
    .B(_0473_),
    .Y(_0474_));
 sg13g2_nor4_1 _1168_ (.A(net196),
    .B(net232),
    .C(net188),
    .D(_0470_),
    .Y(_0475_));
 sg13g2_a21oi_1 _1169_ (.A1(_0130_),
    .A2(_0475_),
    .Y(_0116_),
    .B1(_0474_));
 sg13g2_dfrbp_1 _1170_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net59),
    .D(_0006_),
    .Q_N(_0005_),
    .Q(\rgb_mixer.pwm2.count[0] ));
 sg13g2_dfrbp_1 _1171_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net16),
    .D(_0007_),
    .Q_N(_0580_),
    .Q(\rgb_mixer.pwm2.count[1] ));
 sg13g2_dfrbp_1 _1172_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net15),
    .D(_0008_),
    .Q_N(_0579_),
    .Q(\rgb_mixer.pwm2.count[2] ));
 sg13g2_dfrbp_1 _1173_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net14),
    .D(_0009_),
    .Q_N(_0578_),
    .Q(\rgb_mixer.pwm2.count[3] ));
 sg13g2_dfrbp_1 _1174_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net149),
    .D(net261),
    .Q_N(_0577_),
    .Q(\rgb_mixer.pwm2.count[4] ));
 sg13g2_dfrbp_1 _1175_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net148),
    .D(net252),
    .Q_N(_0576_),
    .Q(\rgb_mixer.pwm2.count[5] ));
 sg13g2_dfrbp_1 _1176_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net147),
    .D(net210),
    .Q_N(_0575_),
    .Q(\rgb_mixer.pwm2.count[6] ));
 sg13g2_dfrbp_1 _1177_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net146),
    .D(net264),
    .Q_N(_0574_),
    .Q(\rgb_mixer.pwm2.count[7] ));
 sg13g2_dfrbp_1 _1178_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net145),
    .D(_0014_),
    .Q_N(_0004_),
    .Q(\rgb_mixer.pwm1.count[0] ));
 sg13g2_dfrbp_1 _1179_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net144),
    .D(_0015_),
    .Q_N(_0573_),
    .Q(\rgb_mixer.pwm1.count[1] ));
 sg13g2_dfrbp_1 _1180_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net143),
    .D(net219),
    .Q_N(_0572_),
    .Q(\rgb_mixer.pwm1.count[2] ));
 sg13g2_dfrbp_1 _1181_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net142),
    .D(net284),
    .Q_N(_0571_),
    .Q(\rgb_mixer.pwm1.count[3] ));
 sg13g2_dfrbp_1 _1182_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net141),
    .D(_0018_),
    .Q_N(_0570_),
    .Q(\rgb_mixer.pwm1.count[4] ));
 sg13g2_dfrbp_1 _1183_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net140),
    .D(net254),
    .Q_N(_0569_),
    .Q(\rgb_mixer.pwm1.count[5] ));
 sg13g2_dfrbp_1 _1184_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net139),
    .D(net225),
    .Q_N(_0568_),
    .Q(\rgb_mixer.pwm1.count[6] ));
 sg13g2_dfrbp_1 _1185_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net138),
    .D(net237),
    .Q_N(_0567_),
    .Q(\rgb_mixer.pwm1.count[7] ));
 sg13g2_dfrbp_1 _1186_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net137),
    .D(_0022_),
    .Q_N(_0566_),
    .Q(\rgb_mixer.pwm2.out ));
 sg13g2_dfrbp_1 _1187_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net136),
    .D(_0023_),
    .Q_N(_0003_),
    .Q(\rgb_mixer.pwm0.count[0] ));
 sg13g2_dfrbp_1 _1188_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net135),
    .D(net242),
    .Q_N(_0565_),
    .Q(\rgb_mixer.pwm0.count[1] ));
 sg13g2_dfrbp_1 _1189_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net134),
    .D(net206),
    .Q_N(_0564_),
    .Q(\rgb_mixer.pwm0.count[2] ));
 sg13g2_dfrbp_1 _1190_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net133),
    .D(net281),
    .Q_N(_0563_),
    .Q(\rgb_mixer.pwm0.count[3] ));
 sg13g2_dfrbp_1 _1191_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net132),
    .D(_0027_),
    .Q_N(_0562_),
    .Q(\rgb_mixer.pwm0.count[4] ));
 sg13g2_dfrbp_1 _1192_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net131),
    .D(net250),
    .Q_N(_0561_),
    .Q(\rgb_mixer.pwm0.count[5] ));
 sg13g2_dfrbp_1 _1193_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net130),
    .D(net222),
    .Q_N(_0560_),
    .Q(\rgb_mixer.pwm0.count[6] ));
 sg13g2_dfrbp_1 _1194_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net129),
    .D(net240),
    .Q_N(_0559_),
    .Q(\rgb_mixer.pwm0.count[7] ));
 sg13g2_dfrbp_1 _1195_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net128),
    .D(_0031_),
    .Q_N(_0558_),
    .Q(\rgb_mixer.pwm1.out ));
 sg13g2_dfrbp_1 _1196_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net127),
    .D(_0032_),
    .Q_N(_0557_),
    .Q(\rgb_mixer.encoder2.old_b ));
 sg13g2_dfrbp_1 _1197_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net126),
    .D(net256),
    .Q_N(_0556_),
    .Q(\rgb_mixer.pwm0.out ));
 sg13g2_dfrbp_1 _1198_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net125),
    .D(net248),
    .Q_N(_0002_),
    .Q(\enc2[0] ));
 sg13g2_dfrbp_1 _1199_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net123),
    .D(_0035_),
    .Q_N(_0555_),
    .Q(\enc2[1] ));
 sg13g2_dfrbp_1 _1200_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net121),
    .D(_0036_),
    .Q_N(_0554_),
    .Q(\enc2[2] ));
 sg13g2_dfrbp_1 _1201_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net119),
    .D(_0037_),
    .Q_N(_0553_),
    .Q(\enc2[3] ));
 sg13g2_dfrbp_1 _1202_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net117),
    .D(_0038_),
    .Q_N(_0552_),
    .Q(\enc2[4] ));
 sg13g2_dfrbp_1 _1203_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net115),
    .D(_0039_),
    .Q_N(_0551_),
    .Q(\enc2[5] ));
 sg13g2_dfrbp_1 _1204_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net113),
    .D(_0040_),
    .Q_N(_0550_),
    .Q(\enc2[6] ));
 sg13g2_dfrbp_1 _1205_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net111),
    .D(net276),
    .Q_N(_0549_),
    .Q(\enc2[7] ));
 sg13g2_dfrbp_1 _1206_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net109),
    .D(_0042_),
    .Q_N(_0548_),
    .Q(\rgb_mixer.encoder1.old_b ));
 sg13g2_dfrbp_1 _1207_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net108),
    .D(_0043_),
    .Q_N(_0547_),
    .Q(\rgb_mixer.encoder2.old_a ));
 sg13g2_dfrbp_1 _1208_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net107),
    .D(net235),
    .Q_N(_0001_),
    .Q(\enc1[0] ));
 sg13g2_dfrbp_1 _1209_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net105),
    .D(_0045_),
    .Q_N(_0546_),
    .Q(\enc1[1] ));
 sg13g2_dfrbp_1 _1210_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net103),
    .D(_0046_),
    .Q_N(_0545_),
    .Q(\enc1[2] ));
 sg13g2_dfrbp_1 _1211_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net101),
    .D(_0047_),
    .Q_N(_0544_),
    .Q(\enc1[3] ));
 sg13g2_dfrbp_1 _1212_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net74),
    .D(_0048_),
    .Q_N(_0543_),
    .Q(\enc1[4] ));
 sg13g2_dfrbp_1 _1213_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net72),
    .D(_0049_),
    .Q_N(_0542_),
    .Q(\enc1[5] ));
 sg13g2_dfrbp_1 _1214_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net70),
    .D(_0050_),
    .Q_N(_0541_),
    .Q(\enc1[6] ));
 sg13g2_dfrbp_1 _1215_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net68),
    .D(_0051_),
    .Q_N(_0540_),
    .Q(\enc1[7] ));
 sg13g2_dfrbp_1 _1216_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net66),
    .D(_0052_),
    .Q_N(_0539_),
    .Q(\rgb_mixer.encoder0.old_b ));
 sg13g2_dfrbp_1 _1217_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net65),
    .D(_0053_),
    .Q_N(_0538_),
    .Q(\rgb_mixer.encoder1.old_a ));
 sg13g2_dfrbp_1 _1218_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net64),
    .D(net246),
    .Q_N(_0000_),
    .Q(\enc0[0] ));
 sg13g2_dfrbp_1 _1219_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net62),
    .D(_0055_),
    .Q_N(_0537_),
    .Q(\enc0[1] ));
 sg13g2_dfrbp_1 _1220_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net60),
    .D(_0056_),
    .Q_N(_0536_),
    .Q(\enc0[2] ));
 sg13g2_dfrbp_1 _1221_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net58),
    .D(_0057_),
    .Q_N(_0535_),
    .Q(\enc0[3] ));
 sg13g2_dfrbp_1 _1222_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net56),
    .D(_0058_),
    .Q_N(_0534_),
    .Q(\enc0[4] ));
 sg13g2_dfrbp_1 _1223_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net54),
    .D(_0059_),
    .Q_N(_0533_),
    .Q(\enc0[5] ));
 sg13g2_dfrbp_1 _1224_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net52),
    .D(_0060_),
    .Q_N(_0532_),
    .Q(\enc0[6] ));
 sg13g2_dfrbp_1 _1225_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net50),
    .D(_0061_),
    .Q_N(_0531_),
    .Q(\enc0[7] ));
 sg13g2_dfrbp_1 _1226_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net48),
    .D(_0062_),
    .Q_N(_0530_),
    .Q(\rgb_mixer.debounce2_b.button_hist[0] ));
 sg13g2_dfrbp_1 _1227_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net47),
    .D(_0063_),
    .Q_N(_0529_),
    .Q(\rgb_mixer.debounce2_b.button_hist[1] ));
 sg13g2_dfrbp_1 _1228_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net46),
    .D(_0064_),
    .Q_N(_0528_),
    .Q(\rgb_mixer.debounce2_b.button_hist[2] ));
 sg13g2_dfrbp_1 _1229_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net45),
    .D(_0065_),
    .Q_N(_0527_),
    .Q(\rgb_mixer.debounce2_b.button_hist[3] ));
 sg13g2_dfrbp_1 _1230_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net44),
    .D(_0066_),
    .Q_N(_0526_),
    .Q(\rgb_mixer.debounce2_b.button_hist[4] ));
 sg13g2_dfrbp_1 _1231_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net43),
    .D(_0067_),
    .Q_N(_0525_),
    .Q(\rgb_mixer.debounce2_b.button_hist[5] ));
 sg13g2_dfrbp_1 _1232_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net42),
    .D(_0068_),
    .Q_N(_0524_),
    .Q(\rgb_mixer.debounce2_b.button_hist[6] ));
 sg13g2_dfrbp_1 _1233_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net41),
    .D(_0069_),
    .Q_N(_0523_),
    .Q(\rgb_mixer.debounce2_b.button_hist[7] ));
 sg13g2_dfrbp_1 _1234_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net40),
    .D(_0070_),
    .Q_N(_0522_),
    .Q(\rgb_mixer.encoder0.old_a ));
 sg13g2_dfrbp_1 _1235_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net39),
    .D(net231),
    .Q_N(_0521_),
    .Q(\rgb_mixer.debounce2_b.debounced ));
 sg13g2_dfrbp_1 _1236_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net37),
    .D(_0072_),
    .Q_N(_0520_),
    .Q(\rgb_mixer.debounce2_a.button_hist[0] ));
 sg13g2_dfrbp_1 _1237_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net36),
    .D(_0073_),
    .Q_N(_0519_),
    .Q(\rgb_mixer.debounce2_a.button_hist[1] ));
 sg13g2_dfrbp_1 _1238_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net35),
    .D(_0074_),
    .Q_N(_0518_),
    .Q(\rgb_mixer.debounce2_a.button_hist[2] ));
 sg13g2_dfrbp_1 _1239_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net34),
    .D(_0075_),
    .Q_N(_0517_),
    .Q(\rgb_mixer.debounce2_a.button_hist[3] ));
 sg13g2_dfrbp_1 _1240_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net33),
    .D(_0076_),
    .Q_N(_0516_),
    .Q(\rgb_mixer.debounce2_a.button_hist[4] ));
 sg13g2_dfrbp_1 _1241_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net32),
    .D(_0077_),
    .Q_N(_0515_),
    .Q(\rgb_mixer.debounce2_a.button_hist[5] ));
 sg13g2_dfrbp_1 _1242_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net31),
    .D(_0078_),
    .Q_N(_0514_),
    .Q(\rgb_mixer.debounce2_a.button_hist[6] ));
 sg13g2_dfrbp_1 _1243_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net30),
    .D(_0079_),
    .Q_N(_0513_),
    .Q(\rgb_mixer.debounce2_a.button_hist[7] ));
 sg13g2_dfrbp_1 _1244_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net29),
    .D(net228),
    .Q_N(_0512_),
    .Q(\rgb_mixer.debounce2_a.debounced ));
 sg13g2_dfrbp_1 _1245_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net27),
    .D(_0081_),
    .Q_N(_0511_),
    .Q(\rgb_mixer.debounce1_b.button_hist[0] ));
 sg13g2_dfrbp_1 _1246_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net26),
    .D(_0082_),
    .Q_N(_0510_),
    .Q(\rgb_mixer.debounce1_b.button_hist[1] ));
 sg13g2_dfrbp_1 _1247_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net25),
    .D(_0083_),
    .Q_N(_0509_),
    .Q(\rgb_mixer.debounce1_b.button_hist[2] ));
 sg13g2_dfrbp_1 _1248_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net24),
    .D(_0084_),
    .Q_N(_0508_),
    .Q(\rgb_mixer.debounce1_b.button_hist[3] ));
 sg13g2_dfrbp_1 _1249_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net23),
    .D(_0085_),
    .Q_N(_0507_),
    .Q(\rgb_mixer.debounce1_b.button_hist[4] ));
 sg13g2_dfrbp_1 _1250_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net22),
    .D(_0086_),
    .Q_N(_0506_),
    .Q(\rgb_mixer.debounce1_b.button_hist[5] ));
 sg13g2_dfrbp_1 _1251_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net21),
    .D(_0087_),
    .Q_N(_0505_),
    .Q(\rgb_mixer.debounce1_b.button_hist[6] ));
 sg13g2_dfrbp_1 _1252_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net20),
    .D(_0088_),
    .Q_N(_0504_),
    .Q(\rgb_mixer.debounce1_b.button_hist[7] ));
 sg13g2_dfrbp_1 _1253_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net19),
    .D(net213),
    .Q_N(_0503_),
    .Q(\rgb_mixer.debounce1_b.debounced ));
 sg13g2_dfrbp_1 _1254_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net17),
    .D(_0090_),
    .Q_N(_0502_),
    .Q(\rgb_mixer.debounce1_a.button_hist[0] ));
 sg13g2_dfrbp_1 _1255_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net124),
    .D(_0091_),
    .Q_N(_0501_),
    .Q(\rgb_mixer.debounce1_a.button_hist[1] ));
 sg13g2_dfrbp_1 _1256_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net122),
    .D(_0092_),
    .Q_N(_0500_),
    .Q(\rgb_mixer.debounce1_a.button_hist[2] ));
 sg13g2_dfrbp_1 _1257_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net120),
    .D(_0093_),
    .Q_N(_0499_),
    .Q(\rgb_mixer.debounce1_a.button_hist[3] ));
 sg13g2_dfrbp_1 _1258_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net118),
    .D(_0094_),
    .Q_N(_0498_),
    .Q(\rgb_mixer.debounce1_a.button_hist[4] ));
 sg13g2_dfrbp_1 _1259_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net116),
    .D(_0095_),
    .Q_N(_0497_),
    .Q(\rgb_mixer.debounce1_a.button_hist[5] ));
 sg13g2_dfrbp_1 _1260_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net114),
    .D(_0096_),
    .Q_N(_0496_),
    .Q(\rgb_mixer.debounce1_a.button_hist[6] ));
 sg13g2_dfrbp_1 _1261_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net112),
    .D(_0097_),
    .Q_N(_0495_),
    .Q(\rgb_mixer.debounce1_a.button_hist[7] ));
 sg13g2_dfrbp_1 _1262_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net110),
    .D(net216),
    .Q_N(_0494_),
    .Q(\rgb_mixer.debounce1_a.debounced ));
 sg13g2_dfrbp_1 _1263_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net104),
    .D(_0099_),
    .Q_N(_0493_),
    .Q(\rgb_mixer.debounce0_b.button_hist[0] ));
 sg13g2_dfrbp_1 _1264_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net102),
    .D(_0100_),
    .Q_N(_0492_),
    .Q(\rgb_mixer.debounce0_b.button_hist[1] ));
 sg13g2_dfrbp_1 _1265_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net75),
    .D(_0101_),
    .Q_N(_0491_),
    .Q(\rgb_mixer.debounce0_b.button_hist[2] ));
 sg13g2_dfrbp_1 _1266_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net73),
    .D(_0102_),
    .Q_N(_0490_),
    .Q(\rgb_mixer.debounce0_b.button_hist[3] ));
 sg13g2_dfrbp_1 _1267_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net71),
    .D(_0103_),
    .Q_N(_0489_),
    .Q(\rgb_mixer.debounce0_b.button_hist[4] ));
 sg13g2_dfrbp_1 _1268_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net69),
    .D(_0104_),
    .Q_N(_0488_),
    .Q(\rgb_mixer.debounce0_b.button_hist[5] ));
 sg13g2_dfrbp_1 _1269_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net67),
    .D(_0105_),
    .Q_N(_0487_),
    .Q(\rgb_mixer.debounce0_b.button_hist[6] ));
 sg13g2_dfrbp_1 _1270_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net63),
    .D(_0106_),
    .Q_N(_0486_),
    .Q(\rgb_mixer.debounce0_b.button_hist[7] ));
 sg13g2_dfrbp_1 _1271_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net61),
    .D(_0107_),
    .Q_N(_0485_),
    .Q(\rgb_mixer.debounce0_b.debounced ));
 sg13g2_dfrbp_1 _1272_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net57),
    .D(_0108_),
    .Q_N(_0484_),
    .Q(\rgb_mixer.debounce0_a.button_hist[0] ));
 sg13g2_dfrbp_1 _1273_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net55),
    .D(_0109_),
    .Q_N(_0483_),
    .Q(\rgb_mixer.debounce0_a.button_hist[1] ));
 sg13g2_dfrbp_1 _1274_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net53),
    .D(_0110_),
    .Q_N(_0482_),
    .Q(\rgb_mixer.debounce0_a.button_hist[2] ));
 sg13g2_dfrbp_1 _1275_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net51),
    .D(_0111_),
    .Q_N(_0481_),
    .Q(\rgb_mixer.debounce0_a.button_hist[3] ));
 sg13g2_dfrbp_1 _1276_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net49),
    .D(_0112_),
    .Q_N(_0480_),
    .Q(\rgb_mixer.debounce0_a.button_hist[4] ));
 sg13g2_dfrbp_1 _1277_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net38),
    .D(_0113_),
    .Q_N(_0479_),
    .Q(\rgb_mixer.debounce0_a.button_hist[5] ));
 sg13g2_dfrbp_1 _1278_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net28),
    .D(_0114_),
    .Q_N(_0478_),
    .Q(\rgb_mixer.debounce0_a.button_hist[6] ));
 sg13g2_dfrbp_1 _1279_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net18),
    .D(_0115_),
    .Q_N(_0477_),
    .Q(\rgb_mixer.debounce0_a.button_hist[7] ));
 sg13g2_dfrbp_1 _1280_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net106),
    .D(net233),
    .Q_N(_0476_),
    .Q(\rgb_mixer.debounce0_a.debounced ));
 sg13g2_tiehi _1172__15 (.L_HI(net15));
 sg13g2_tiehi _1171__16 (.L_HI(net16));
 sg13g2_tiehi _1254__17 (.L_HI(net17));
 sg13g2_tiehi _1279__18 (.L_HI(net18));
 sg13g2_tiehi _1253__19 (.L_HI(net19));
 sg13g2_tiehi _1252__20 (.L_HI(net20));
 sg13g2_tiehi _1251__21 (.L_HI(net21));
 sg13g2_tiehi _1250__22 (.L_HI(net22));
 sg13g2_tiehi _1249__23 (.L_HI(net23));
 sg13g2_tiehi _1248__24 (.L_HI(net24));
 sg13g2_tiehi _1247__25 (.L_HI(net25));
 sg13g2_tiehi _1246__26 (.L_HI(net26));
 sg13g2_tiehi _1245__27 (.L_HI(net27));
 sg13g2_tiehi _1278__28 (.L_HI(net28));
 sg13g2_tiehi _1244__29 (.L_HI(net29));
 sg13g2_tiehi _1243__30 (.L_HI(net30));
 sg13g2_tiehi _1242__31 (.L_HI(net31));
 sg13g2_tiehi _1241__32 (.L_HI(net32));
 sg13g2_tiehi _1240__33 (.L_HI(net33));
 sg13g2_tiehi _1239__34 (.L_HI(net34));
 sg13g2_tiehi _1238__35 (.L_HI(net35));
 sg13g2_tiehi _1237__36 (.L_HI(net36));
 sg13g2_tiehi _1236__37 (.L_HI(net37));
 sg13g2_tiehi _1277__38 (.L_HI(net38));
 sg13g2_tiehi _1235__39 (.L_HI(net39));
 sg13g2_tiehi _1234__40 (.L_HI(net40));
 sg13g2_tiehi _1233__41 (.L_HI(net41));
 sg13g2_tiehi _1232__42 (.L_HI(net42));
 sg13g2_tiehi _1231__43 (.L_HI(net43));
 sg13g2_tiehi _1230__44 (.L_HI(net44));
 sg13g2_tiehi _1229__45 (.L_HI(net45));
 sg13g2_tiehi _1228__46 (.L_HI(net46));
 sg13g2_tiehi _1227__47 (.L_HI(net47));
 sg13g2_tiehi _1226__48 (.L_HI(net48));
 sg13g2_tiehi _1276__49 (.L_HI(net49));
 sg13g2_tiehi _1225__50 (.L_HI(net50));
 sg13g2_tiehi _1275__51 (.L_HI(net51));
 sg13g2_tiehi _1224__52 (.L_HI(net52));
 sg13g2_tiehi _1274__53 (.L_HI(net53));
 sg13g2_tiehi _1223__54 (.L_HI(net54));
 sg13g2_tiehi _1273__55 (.L_HI(net55));
 sg13g2_tiehi _1222__56 (.L_HI(net56));
 sg13g2_tiehi _1272__57 (.L_HI(net57));
 sg13g2_tiehi _1221__58 (.L_HI(net58));
 sg13g2_tiehi _1170__59 (.L_HI(net59));
 sg13g2_tiehi _1220__60 (.L_HI(net60));
 sg13g2_tiehi _1271__61 (.L_HI(net61));
 sg13g2_tiehi _1219__62 (.L_HI(net62));
 sg13g2_tiehi _1270__63 (.L_HI(net63));
 sg13g2_tiehi _1218__64 (.L_HI(net64));
 sg13g2_tiehi _1217__65 (.L_HI(net65));
 sg13g2_tiehi _1216__66 (.L_HI(net66));
 sg13g2_tiehi _1269__67 (.L_HI(net67));
 sg13g2_tiehi _1215__68 (.L_HI(net68));
 sg13g2_tiehi _1268__69 (.L_HI(net69));
 sg13g2_tiehi _1214__70 (.L_HI(net70));
 sg13g2_tiehi _1267__71 (.L_HI(net71));
 sg13g2_tiehi _1213__72 (.L_HI(net72));
 sg13g2_tiehi _1266__73 (.L_HI(net73));
 sg13g2_tiehi _1212__74 (.L_HI(net74));
 sg13g2_tiehi _1265__75 (.L_HI(net75));
 sg13g2_tiehi _1211__76 (.L_HI(net101));
 sg13g2_tiehi _1264__77 (.L_HI(net102));
 sg13g2_tiehi _1210__78 (.L_HI(net103));
 sg13g2_tiehi _1263__79 (.L_HI(net104));
 sg13g2_tiehi _1209__80 (.L_HI(net105));
 sg13g2_tiehi _1280__81 (.L_HI(net106));
 sg13g2_tiehi _1208__82 (.L_HI(net107));
 sg13g2_tiehi _1207__83 (.L_HI(net108));
 sg13g2_tiehi _1206__84 (.L_HI(net109));
 sg13g2_tiehi _1262__85 (.L_HI(net110));
 sg13g2_tiehi _1205__86 (.L_HI(net111));
 sg13g2_tiehi _1261__87 (.L_HI(net112));
 sg13g2_tiehi _1204__88 (.L_HI(net113));
 sg13g2_tiehi _1260__89 (.L_HI(net114));
 sg13g2_tiehi _1203__90 (.L_HI(net115));
 sg13g2_tiehi _1259__91 (.L_HI(net116));
 sg13g2_tiehi _1202__92 (.L_HI(net117));
 sg13g2_tiehi _1258__93 (.L_HI(net118));
 sg13g2_tiehi _1201__94 (.L_HI(net119));
 sg13g2_tiehi _1257__95 (.L_HI(net120));
 sg13g2_tiehi _1200__96 (.L_HI(net121));
 sg13g2_tiehi _1256__97 (.L_HI(net122));
 sg13g2_tiehi _1199__98 (.L_HI(net123));
 sg13g2_tiehi _1255__99 (.L_HI(net124));
 sg13g2_tiehi _1198__100 (.L_HI(net125));
 sg13g2_tiehi _1197__101 (.L_HI(net126));
 sg13g2_tiehi _1196__102 (.L_HI(net127));
 sg13g2_tiehi _1195__103 (.L_HI(net128));
 sg13g2_tiehi _1194__104 (.L_HI(net129));
 sg13g2_tiehi _1193__105 (.L_HI(net130));
 sg13g2_tiehi _1192__106 (.L_HI(net131));
 sg13g2_tiehi _1191__107 (.L_HI(net132));
 sg13g2_tiehi _1190__108 (.L_HI(net133));
 sg13g2_tiehi _1189__109 (.L_HI(net134));
 sg13g2_tiehi _1188__110 (.L_HI(net135));
 sg13g2_tiehi _1187__111 (.L_HI(net136));
 sg13g2_tiehi _1186__112 (.L_HI(net137));
 sg13g2_tiehi _1185__113 (.L_HI(net138));
 sg13g2_tiehi _1184__114 (.L_HI(net139));
 sg13g2_tiehi _1183__115 (.L_HI(net140));
 sg13g2_tiehi _1182__116 (.L_HI(net141));
 sg13g2_tiehi _1181__117 (.L_HI(net142));
 sg13g2_tiehi _1180__118 (.L_HI(net143));
 sg13g2_tiehi _1179__119 (.L_HI(net144));
 sg13g2_tiehi _1178__120 (.L_HI(net145));
 sg13g2_tiehi _1177__121 (.L_HI(net146));
 sg13g2_tiehi _1176__122 (.L_HI(net147));
 sg13g2_tiehi _1175__123 (.L_HI(net148));
 sg13g2_tiehi _1174__124 (.L_HI(net149));
 sg13g2_tiehi tt_um_tmkong_rgb_mixer_125 (.L_HI(net150));
 sg13g2_tiehi tt_um_tmkong_rgb_mixer_126 (.L_HI(net151));
 sg13g2_tiehi tt_um_tmkong_rgb_mixer_127 (.L_HI(net152));
 sg13g2_tiehi tt_um_tmkong_rgb_mixer_128 (.L_HI(net153));
 sg13g2_tiehi tt_um_tmkong_rgb_mixer_129 (.L_HI(net154));
 sg13g2_tiehi tt_um_tmkong_rgb_mixer_130 (.L_HI(net155));
 sg13g2_tiehi tt_um_tmkong_rgb_mixer_131 (.L_HI(net156));
 sg13g2_tiehi tt_um_tmkong_rgb_mixer_132 (.L_HI(net157));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_tmkong_rgb_mixer_10 (.L_LO(net10));
 sg13g2_tielo tt_um_tmkong_rgb_mixer_11 (.L_LO(net11));
 sg13g2_tielo tt_um_tmkong_rgb_mixer_12 (.L_LO(net12));
 sg13g2_tielo tt_um_tmkong_rgb_mixer_13 (.L_LO(net13));
 sg13g2_tiehi _1173__14 (.L_HI(net14));
 sg13g2_buf_2 _1405_ (.A(\rgb_mixer.pwm0.out ),
    .X(uo_out[0]));
 sg13g2_buf_1 _1406_ (.A(\rgb_mixer.pwm1.out ),
    .X(uo_out[1]));
 sg13g2_buf_1 _1407_ (.A(\rgb_mixer.pwm2.out ),
    .X(uo_out[2]));
 sg13g2_buf_2 fanout76 (.A(_0395_),
    .X(net76));
 sg13g2_buf_1 fanout77 (.A(_0395_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0339_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_0286_),
    .X(net79));
 sg13g2_buf_4 fanout80 (.X(net80),
    .A(_0400_));
 sg13g2_buf_4 fanout81 (.X(net81),
    .A(_0344_));
 sg13g2_buf_4 fanout82 (.X(net82),
    .A(_0291_));
 sg13g2_buf_4 fanout83 (.X(net83),
    .A(_0143_));
 sg13g2_buf_2 fanout84 (.A(_0143_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(net86),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(net90),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(net89),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(net89),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(net90),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(rst_n),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(net94),
    .X(net91));
 sg13g2_buf_4 fanout92 (.X(net92),
    .A(net93));
 sg13g2_buf_1 fanout93 (.A(net94),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(rst_n),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(net96),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(net100),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(net100),
    .X(net97));
 sg13g2_buf_1 fanout98 (.A(net100),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(net100),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(rst_n),
    .X(net100));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_tmkong_rgb_mixer_9 (.L_LO(net9));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0005_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0004_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0003_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold4 (.A(\rgb_mixer.debounce1_a.button_hist[4] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold5 (.A(\rgb_mixer.debounce0_a.button_hist[1] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold6 (.A(\rgb_mixer.debounce2_b.button_hist[3] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold7 (.A(\rgb_mixer.debounce1_b.button_hist[4] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold8 (.A(\rgb_mixer.debounce0_b.button_hist[2] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold9 (.A(\rgb_mixer.debounce1_b.button_hist[3] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold10 (.A(\rgb_mixer.debounce1_a.button_hist[0] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold11 (.A(\rgb_mixer.debounce1_a.button_hist[5] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold12 (.A(\rgb_mixer.debounce0_a.button_hist[3] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold13 (.A(\rgb_mixer.debounce0_b.button_hist[3] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold14 (.A(\rgb_mixer.debounce2_a.button_hist[4] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold15 (.A(\rgb_mixer.debounce2_b.button_hist[4] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold16 (.A(\rgb_mixer.debounce2_b.button_hist[2] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold17 (.A(\rgb_mixer.debounce2_a.button_hist[1] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold18 (.A(\rgb_mixer.debounce2_a.button_hist[0] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold19 (.A(\rgb_mixer.debounce1_b.button_hist[1] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold20 (.A(\rgb_mixer.debounce2_a.button_hist[2] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold21 (.A(\rgb_mixer.debounce2_b.button_hist[1] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold22 (.A(\rgb_mixer.debounce1_a.button_hist[1] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold23 (.A(\rgb_mixer.debounce0_b.button_hist[4] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold24 (.A(\rgb_mixer.debounce0_a.button_hist[0] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold25 (.A(\rgb_mixer.debounce2_a.button_hist[6] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold26 (.A(\rgb_mixer.debounce0_b.button_hist[0] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold27 (.A(\rgb_mixer.debounce0_b.button_hist[1] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold28 (.A(\rgb_mixer.debounce2_b.button_hist[0] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold29 (.A(\rgb_mixer.debounce0_b.button_hist[6] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold30 (.A(\rgb_mixer.debounce2_b.button_hist[5] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold31 (.A(\rgb_mixer.debounce0_a.button_hist[6] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold32 (.A(\rgb_mixer.debounce0_a.button_hist[2] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold33 (.A(\rgb_mixer.debounce1_a.button_hist[2] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold34 (.A(\rgb_mixer.debounce1_b.button_hist[0] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold35 (.A(\rgb_mixer.debounce1_b.button_hist[2] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold36 (.A(\rgb_mixer.debounce0_b.button_hist[5] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold37 (.A(\rgb_mixer.debounce2_b.button_hist[6] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold38 (.A(\rgb_mixer.debounce1_b.button_hist[6] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold39 (.A(\rgb_mixer.debounce0_a.button_hist[4] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold40 (.A(\rgb_mixer.debounce2_a.button_hist[5] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold41 (.A(\rgb_mixer.debounce2_a.button_hist[3] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold42 (.A(\rgb_mixer.debounce1_b.button_hist[5] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold43 (.A(\rgb_mixer.debounce1_a.button_hist[6] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold44 (.A(\rgb_mixer.debounce0_a.button_hist[5] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold45 (.A(\rgb_mixer.debounce1_a.button_hist[3] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold46 (.A(\rgb_mixer.debounce0_b.debounced ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold47 (.A(\rgb_mixer.pwm0.count[2] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0215_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0025_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold50 (.A(\rgb_mixer.debounce0_b.button_hist[7] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold51 (.A(\rgb_mixer.pwm2.count[6] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0172_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0012_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold54 (.A(\rgb_mixer.debounce1_b.debounced ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0457_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0089_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold57 (.A(\rgb_mixer.debounce1_a.debounced ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0463_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0098_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold60 (.A(\rgb_mixer.pwm1.count[2] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0177_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0016_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold63 (.A(\rgb_mixer.pwm0.count[6] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0223_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0029_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold66 (.A(\rgb_mixer.pwm1.count[6] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0185_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0020_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold69 (.A(\rgb_mixer.debounce2_a.debounced ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0451_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0080_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold72 (.A(\rgb_mixer.debounce2_b.debounced ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0445_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0071_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold75 (.A(\rgb_mixer.debounce0_a.button_hist[7] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0116_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0001_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0044_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold79 (.A(\rgb_mixer.pwm1.count[7] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0021_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold81 (.A(\rgb_mixer.debounce0_a.debounced ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold82 (.A(\rgb_mixer.pwm0.count[7] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0030_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold84 (.A(\rgb_mixer.pwm0.count[1] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0024_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold86 (.A(\rgb_mixer.pwm2.count[2] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0164_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0000_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0054_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0002_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0034_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold92 (.A(\rgb_mixer.pwm0.count[5] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0028_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold94 (.A(\rgb_mixer.pwm2.count[5] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0011_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold96 (.A(\rgb_mixer.pwm1.count[5] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0019_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold98 (.A(\enc0[7] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0033_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold100 (.A(\rgb_mixer.pwm0.count[4] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0220_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold102 (.A(\rgb_mixer.pwm2.count[4] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0169_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0010_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold105 (.A(\enc1[1] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold106 (.A(\rgb_mixer.pwm2.count[7] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0013_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold108 (.A(\rgb_mixer.pwm1.count[4] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0182_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold110 (.A(\rgb_mixer.pwm1.count[1] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0176_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold112 (.A(\enc0[1] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold113 (.A(\rgb_mixer.pwm2.count[1] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0163_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold115 (.A(\enc2[1] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold116 (.A(\enc1[7] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold117 (.A(\enc0[6] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold118 (.A(\enc2[7] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0041_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold120 (.A(\enc0[7] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold121 (.A(\enc0[4] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold122 (.A(\rgb_mixer.pwm0.count[3] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0219_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0026_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold125 (.A(\rgb_mixer.pwm1.count[3] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0181_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0017_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold128 (.A(\enc1[6] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold129 (.A(\enc0[5] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold130 (.A(\enc2[5] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold131 (.A(\enc1[4] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold132 (.A(\enc2[2] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold133 (.A(\enc2[3] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold134 (.A(\enc1[5] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold135 (.A(\enc0[3] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold136 (.A(\enc0[2] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold137 (.A(\enc1[3] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold138 (.A(\enc2[6] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold139 (.A(\enc1[7] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0383_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold141 (.A(\enc2[4] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold142 (.A(\rgb_mixer.pwm2.count[3] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold143 (.A(\enc1[2] ),
    .X(net300));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_4 FILLER_14_154 ();
 sg13g2_fill_2 FILLER_14_158 ();
 sg13g2_decap_8 FILLER_14_164 ();
 sg13g2_decap_4 FILLER_14_183 ();
 sg13g2_fill_1 FILLER_14_187 ();
 sg13g2_decap_8 FILLER_14_192 ();
 sg13g2_decap_8 FILLER_14_199 ();
 sg13g2_decap_8 FILLER_14_206 ();
 sg13g2_decap_4 FILLER_14_213 ();
 sg13g2_fill_1 FILLER_14_217 ();
 sg13g2_decap_4 FILLER_14_228 ();
 sg13g2_decap_8 FILLER_14_237 ();
 sg13g2_decap_8 FILLER_14_244 ();
 sg13g2_decap_8 FILLER_14_251 ();
 sg13g2_decap_8 FILLER_14_258 ();
 sg13g2_decap_8 FILLER_14_265 ();
 sg13g2_decap_8 FILLER_14_272 ();
 sg13g2_decap_8 FILLER_14_279 ();
 sg13g2_decap_8 FILLER_14_286 ();
 sg13g2_decap_8 FILLER_14_293 ();
 sg13g2_decap_8 FILLER_14_300 ();
 sg13g2_decap_8 FILLER_14_307 ();
 sg13g2_decap_8 FILLER_14_314 ();
 sg13g2_decap_8 FILLER_14_321 ();
 sg13g2_decap_8 FILLER_14_328 ();
 sg13g2_decap_8 FILLER_14_335 ();
 sg13g2_decap_8 FILLER_14_342 ();
 sg13g2_decap_8 FILLER_14_349 ();
 sg13g2_decap_8 FILLER_14_356 ();
 sg13g2_decap_8 FILLER_14_363 ();
 sg13g2_decap_8 FILLER_14_370 ();
 sg13g2_decap_8 FILLER_14_377 ();
 sg13g2_decap_8 FILLER_14_384 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_fill_2 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_43 ();
 sg13g2_decap_8 FILLER_15_50 ();
 sg13g2_decap_8 FILLER_15_57 ();
 sg13g2_decap_8 FILLER_15_64 ();
 sg13g2_decap_8 FILLER_15_71 ();
 sg13g2_decap_8 FILLER_15_78 ();
 sg13g2_decap_8 FILLER_15_85 ();
 sg13g2_decap_8 FILLER_15_92 ();
 sg13g2_decap_8 FILLER_15_99 ();
 sg13g2_decap_8 FILLER_15_106 ();
 sg13g2_decap_8 FILLER_15_113 ();
 sg13g2_decap_8 FILLER_15_120 ();
 sg13g2_decap_8 FILLER_15_127 ();
 sg13g2_decap_4 FILLER_15_134 ();
 sg13g2_fill_2 FILLER_15_142 ();
 sg13g2_fill_2 FILLER_15_175 ();
 sg13g2_fill_2 FILLER_15_203 ();
 sg13g2_fill_1 FILLER_15_205 ();
 sg13g2_fill_1 FILLER_15_232 ();
 sg13g2_decap_8 FILLER_15_246 ();
 sg13g2_decap_8 FILLER_15_253 ();
 sg13g2_decap_8 FILLER_15_260 ();
 sg13g2_decap_8 FILLER_15_267 ();
 sg13g2_decap_8 FILLER_15_274 ();
 sg13g2_decap_8 FILLER_15_281 ();
 sg13g2_decap_8 FILLER_15_288 ();
 sg13g2_decap_8 FILLER_15_295 ();
 sg13g2_decap_8 FILLER_15_302 ();
 sg13g2_decap_8 FILLER_15_309 ();
 sg13g2_decap_8 FILLER_15_316 ();
 sg13g2_decap_8 FILLER_15_323 ();
 sg13g2_decap_8 FILLER_15_330 ();
 sg13g2_decap_8 FILLER_15_337 ();
 sg13g2_decap_8 FILLER_15_344 ();
 sg13g2_decap_8 FILLER_15_351 ();
 sg13g2_decap_8 FILLER_15_358 ();
 sg13g2_decap_8 FILLER_15_365 ();
 sg13g2_decap_8 FILLER_15_372 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_60 ();
 sg13g2_decap_8 FILLER_16_67 ();
 sg13g2_decap_8 FILLER_16_74 ();
 sg13g2_decap_8 FILLER_16_81 ();
 sg13g2_decap_8 FILLER_16_88 ();
 sg13g2_fill_2 FILLER_16_95 ();
 sg13g2_fill_1 FILLER_16_97 ();
 sg13g2_fill_1 FILLER_16_107 ();
 sg13g2_fill_1 FILLER_16_121 ();
 sg13g2_fill_2 FILLER_16_153 ();
 sg13g2_fill_2 FILLER_16_189 ();
 sg13g2_fill_1 FILLER_16_191 ();
 sg13g2_fill_1 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_251 ();
 sg13g2_decap_8 FILLER_16_258 ();
 sg13g2_decap_8 FILLER_16_265 ();
 sg13g2_decap_8 FILLER_16_272 ();
 sg13g2_decap_8 FILLER_16_279 ();
 sg13g2_decap_8 FILLER_16_286 ();
 sg13g2_decap_8 FILLER_16_293 ();
 sg13g2_decap_8 FILLER_16_300 ();
 sg13g2_decap_8 FILLER_16_307 ();
 sg13g2_decap_8 FILLER_16_314 ();
 sg13g2_decap_8 FILLER_16_321 ();
 sg13g2_decap_8 FILLER_16_328 ();
 sg13g2_decap_8 FILLER_16_335 ();
 sg13g2_decap_8 FILLER_16_342 ();
 sg13g2_decap_8 FILLER_16_349 ();
 sg13g2_decap_8 FILLER_16_356 ();
 sg13g2_decap_8 FILLER_16_363 ();
 sg13g2_decap_8 FILLER_16_370 ();
 sg13g2_decap_8 FILLER_16_377 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_fill_1 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_27 ();
 sg13g2_fill_1 FILLER_17_29 ();
 sg13g2_fill_1 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_fill_1 FILLER_17_70 ();
 sg13g2_fill_2 FILLER_17_97 ();
 sg13g2_fill_1 FILLER_17_99 ();
 sg13g2_fill_2 FILLER_17_126 ();
 sg13g2_decap_4 FILLER_17_133 ();
 sg13g2_fill_1 FILLER_17_142 ();
 sg13g2_fill_2 FILLER_17_182 ();
 sg13g2_fill_2 FILLER_17_218 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_4 FILLER_18_7 ();
 sg13g2_fill_1 FILLER_18_11 ();
 sg13g2_fill_2 FILLER_18_16 ();
 sg13g2_decap_8 FILLER_18_66 ();
 sg13g2_fill_2 FILLER_18_73 ();
 sg13g2_fill_1 FILLER_18_89 ();
 sg13g2_fill_2 FILLER_18_119 ();
 sg13g2_fill_2 FILLER_18_154 ();
 sg13g2_fill_1 FILLER_18_156 ();
 sg13g2_fill_2 FILLER_18_171 ();
 sg13g2_fill_2 FILLER_18_182 ();
 sg13g2_fill_1 FILLER_18_184 ();
 sg13g2_fill_2 FILLER_18_193 ();
 sg13g2_decap_4 FILLER_18_200 ();
 sg13g2_fill_2 FILLER_18_207 ();
 sg13g2_fill_2 FILLER_18_240 ();
 sg13g2_fill_1 FILLER_18_242 ();
 sg13g2_decap_8 FILLER_18_269 ();
 sg13g2_decap_8 FILLER_18_276 ();
 sg13g2_decap_8 FILLER_18_283 ();
 sg13g2_fill_2 FILLER_18_290 ();
 sg13g2_fill_1 FILLER_18_292 ();
 sg13g2_decap_4 FILLER_18_297 ();
 sg13g2_decap_8 FILLER_18_306 ();
 sg13g2_fill_2 FILLER_18_313 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_fill_2 FILLER_19_37 ();
 sg13g2_fill_1 FILLER_19_61 ();
 sg13g2_fill_2 FILLER_19_67 ();
 sg13g2_decap_4 FILLER_19_90 ();
 sg13g2_fill_2 FILLER_19_114 ();
 sg13g2_fill_2 FILLER_19_156 ();
 sg13g2_fill_1 FILLER_19_158 ();
 sg13g2_fill_2 FILLER_19_208 ();
 sg13g2_decap_4 FILLER_19_215 ();
 sg13g2_fill_1 FILLER_19_219 ();
 sg13g2_fill_1 FILLER_19_237 ();
 sg13g2_decap_8 FILLER_19_263 ();
 sg13g2_fill_2 FILLER_19_270 ();
 sg13g2_decap_4 FILLER_19_277 ();
 sg13g2_fill_1 FILLER_19_281 ();
 sg13g2_decap_8 FILLER_19_337 ();
 sg13g2_decap_8 FILLER_19_344 ();
 sg13g2_decap_8 FILLER_19_351 ();
 sg13g2_decap_8 FILLER_19_358 ();
 sg13g2_decap_8 FILLER_19_365 ();
 sg13g2_decap_8 FILLER_19_372 ();
 sg13g2_decap_8 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_44 ();
 sg13g2_decap_4 FILLER_20_65 ();
 sg13g2_decap_8 FILLER_20_72 ();
 sg13g2_fill_2 FILLER_20_79 ();
 sg13g2_fill_1 FILLER_20_81 ();
 sg13g2_decap_4 FILLER_20_85 ();
 sg13g2_fill_1 FILLER_20_89 ();
 sg13g2_fill_2 FILLER_20_100 ();
 sg13g2_fill_2 FILLER_20_115 ();
 sg13g2_fill_1 FILLER_20_117 ();
 sg13g2_fill_2 FILLER_20_144 ();
 sg13g2_fill_1 FILLER_20_146 ();
 sg13g2_fill_2 FILLER_20_153 ();
 sg13g2_decap_8 FILLER_20_177 ();
 sg13g2_fill_2 FILLER_20_184 ();
 sg13g2_fill_1 FILLER_20_191 ();
 sg13g2_fill_2 FILLER_20_197 ();
 sg13g2_fill_1 FILLER_20_199 ();
 sg13g2_fill_2 FILLER_20_209 ();
 sg13g2_fill_2 FILLER_20_242 ();
 sg13g2_fill_2 FILLER_20_332 ();
 sg13g2_fill_1 FILLER_20_334 ();
 sg13g2_fill_2 FILLER_20_344 ();
 sg13g2_fill_1 FILLER_20_346 ();
 sg13g2_decap_8 FILLER_20_356 ();
 sg13g2_decap_8 FILLER_20_363 ();
 sg13g2_decap_8 FILLER_20_370 ();
 sg13g2_decap_8 FILLER_20_377 ();
 sg13g2_decap_8 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_25 ();
 sg13g2_decap_8 FILLER_21_62 ();
 sg13g2_decap_4 FILLER_21_69 ();
 sg13g2_fill_2 FILLER_21_77 ();
 sg13g2_fill_1 FILLER_21_79 ();
 sg13g2_fill_1 FILLER_21_95 ();
 sg13g2_fill_2 FILLER_21_101 ();
 sg13g2_fill_1 FILLER_21_103 ();
 sg13g2_fill_2 FILLER_21_112 ();
 sg13g2_fill_2 FILLER_21_118 ();
 sg13g2_fill_1 FILLER_21_120 ();
 sg13g2_fill_2 FILLER_21_126 ();
 sg13g2_decap_4 FILLER_21_150 ();
 sg13g2_fill_2 FILLER_21_176 ();
 sg13g2_decap_4 FILLER_21_221 ();
 sg13g2_fill_1 FILLER_21_337 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_2 ();
 sg13g2_decap_8 FILLER_22_52 ();
 sg13g2_fill_2 FILLER_22_59 ();
 sg13g2_fill_1 FILLER_22_61 ();
 sg13g2_fill_1 FILLER_22_88 ();
 sg13g2_fill_1 FILLER_22_97 ();
 sg13g2_fill_1 FILLER_22_111 ();
 sg13g2_fill_1 FILLER_22_125 ();
 sg13g2_fill_1 FILLER_22_152 ();
 sg13g2_fill_2 FILLER_22_184 ();
 sg13g2_fill_1 FILLER_22_186 ();
 sg13g2_fill_1 FILLER_22_214 ();
 sg13g2_decap_8 FILLER_22_244 ();
 sg13g2_decap_4 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_300 ();
 sg13g2_fill_2 FILLER_22_316 ();
 sg13g2_fill_2 FILLER_22_341 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_7 ();
 sg13g2_fill_2 FILLER_23_11 ();
 sg13g2_decap_8 FILLER_23_17 ();
 sg13g2_decap_4 FILLER_23_24 ();
 sg13g2_fill_1 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_34 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_4 FILLER_23_89 ();
 sg13g2_fill_1 FILLER_23_93 ();
 sg13g2_fill_2 FILLER_23_98 ();
 sg13g2_fill_1 FILLER_23_105 ();
 sg13g2_decap_4 FILLER_23_114 ();
 sg13g2_fill_1 FILLER_23_118 ();
 sg13g2_decap_4 FILLER_23_129 ();
 sg13g2_fill_2 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_148 ();
 sg13g2_fill_1 FILLER_23_155 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_fill_2 FILLER_23_168 ();
 sg13g2_fill_2 FILLER_23_174 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_fill_2 FILLER_23_238 ();
 sg13g2_fill_1 FILLER_23_240 ();
 sg13g2_fill_2 FILLER_23_245 ();
 sg13g2_fill_1 FILLER_23_247 ();
 sg13g2_fill_2 FILLER_23_266 ();
 sg13g2_fill_1 FILLER_23_268 ();
 sg13g2_fill_2 FILLER_23_278 ();
 sg13g2_fill_2 FILLER_23_306 ();
 sg13g2_fill_1 FILLER_23_308 ();
 sg13g2_fill_1 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_4 ();
 sg13g2_fill_2 FILLER_24_31 ();
 sg13g2_fill_1 FILLER_24_82 ();
 sg13g2_decap_8 FILLER_24_110 ();
 sg13g2_decap_4 FILLER_24_117 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_4 FILLER_24_140 ();
 sg13g2_fill_2 FILLER_24_144 ();
 sg13g2_fill_1 FILLER_24_152 ();
 sg13g2_fill_1 FILLER_24_203 ();
 sg13g2_fill_2 FILLER_24_221 ();
 sg13g2_fill_2 FILLER_24_262 ();
 sg13g2_fill_1 FILLER_24_264 ();
 sg13g2_fill_1 FILLER_24_293 ();
 sg13g2_fill_1 FILLER_24_303 ();
 sg13g2_fill_2 FILLER_24_330 ();
 sg13g2_fill_2 FILLER_24_355 ();
 sg13g2_decap_8 FILLER_24_375 ();
 sg13g2_decap_8 FILLER_24_382 ();
 sg13g2_decap_4 FILLER_24_389 ();
 sg13g2_fill_1 FILLER_24_393 ();
 sg13g2_fill_2 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_4 ();
 sg13g2_fill_2 FILLER_25_41 ();
 sg13g2_fill_1 FILLER_25_66 ();
 sg13g2_decap_4 FILLER_25_81 ();
 sg13g2_decap_8 FILLER_25_90 ();
 sg13g2_fill_1 FILLER_25_97 ();
 sg13g2_decap_4 FILLER_25_111 ();
 sg13g2_fill_2 FILLER_25_115 ();
 sg13g2_fill_1 FILLER_25_125 ();
 sg13g2_decap_8 FILLER_25_162 ();
 sg13g2_fill_2 FILLER_25_169 ();
 sg13g2_fill_1 FILLER_25_192 ();
 sg13g2_fill_2 FILLER_25_200 ();
 sg13g2_decap_4 FILLER_25_254 ();
 sg13g2_fill_1 FILLER_25_298 ();
 sg13g2_decap_8 FILLER_25_304 ();
 sg13g2_decap_4 FILLER_25_311 ();
 sg13g2_decap_8 FILLER_25_323 ();
 sg13g2_fill_1 FILLER_25_340 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_27 ();
 sg13g2_fill_1 FILLER_26_55 ();
 sg13g2_fill_2 FILLER_26_61 ();
 sg13g2_decap_4 FILLER_26_115 ();
 sg13g2_fill_1 FILLER_26_119 ();
 sg13g2_decap_4 FILLER_26_144 ();
 sg13g2_fill_1 FILLER_26_148 ();
 sg13g2_fill_2 FILLER_26_203 ();
 sg13g2_fill_1 FILLER_26_205 ();
 sg13g2_fill_2 FILLER_26_211 ();
 sg13g2_fill_1 FILLER_26_213 ();
 sg13g2_decap_4 FILLER_26_217 ();
 sg13g2_fill_1 FILLER_26_221 ();
 sg13g2_fill_2 FILLER_26_248 ();
 sg13g2_fill_1 FILLER_26_250 ();
 sg13g2_fill_1 FILLER_26_256 ();
 sg13g2_decap_8 FILLER_26_262 ();
 sg13g2_fill_2 FILLER_26_304 ();
 sg13g2_fill_2 FILLER_26_358 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_40 ();
 sg13g2_decap_8 FILLER_27_94 ();
 sg13g2_decap_8 FILLER_27_101 ();
 sg13g2_decap_4 FILLER_27_112 ();
 sg13g2_fill_2 FILLER_27_126 ();
 sg13g2_decap_4 FILLER_27_132 ();
 sg13g2_fill_1 FILLER_27_136 ();
 sg13g2_decap_8 FILLER_27_163 ();
 sg13g2_fill_1 FILLER_27_170 ();
 sg13g2_fill_2 FILLER_27_184 ();
 sg13g2_decap_4 FILLER_27_196 ();
 sg13g2_fill_1 FILLER_27_200 ();
 sg13g2_decap_8 FILLER_27_223 ();
 sg13g2_decap_4 FILLER_27_235 ();
 sg13g2_fill_2 FILLER_27_273 ();
 sg13g2_fill_1 FILLER_27_330 ();
 sg13g2_decap_4 FILLER_27_354 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_4 FILLER_28_14 ();
 sg13g2_fill_2 FILLER_28_53 ();
 sg13g2_fill_1 FILLER_28_60 ();
 sg13g2_fill_2 FILLER_28_123 ();
 sg13g2_fill_1 FILLER_28_125 ();
 sg13g2_decap_4 FILLER_28_135 ();
 sg13g2_fill_2 FILLER_28_139 ();
 sg13g2_decap_4 FILLER_28_146 ();
 sg13g2_decap_8 FILLER_28_163 ();
 sg13g2_decap_4 FILLER_28_170 ();
 sg13g2_fill_2 FILLER_28_174 ();
 sg13g2_decap_4 FILLER_28_186 ();
 sg13g2_decap_8 FILLER_28_236 ();
 sg13g2_fill_2 FILLER_28_267 ();
 sg13g2_fill_2 FILLER_28_287 ();
 sg13g2_fill_1 FILLER_28_289 ();
 sg13g2_decap_4 FILLER_28_307 ();
 sg13g2_fill_1 FILLER_28_311 ();
 sg13g2_fill_2 FILLER_28_316 ();
 sg13g2_fill_2 FILLER_28_341 ();
 sg13g2_fill_2 FILLER_28_352 ();
 sg13g2_fill_1 FILLER_28_377 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_fill_2 FILLER_29_28 ();
 sg13g2_fill_2 FILLER_29_70 ();
 sg13g2_fill_1 FILLER_29_72 ();
 sg13g2_fill_1 FILLER_29_108 ();
 sg13g2_fill_1 FILLER_29_118 ();
 sg13g2_fill_2 FILLER_29_128 ();
 sg13g2_fill_1 FILLER_29_130 ();
 sg13g2_decap_4 FILLER_29_199 ();
 sg13g2_fill_2 FILLER_29_211 ();
 sg13g2_fill_2 FILLER_29_223 ();
 sg13g2_fill_2 FILLER_29_230 ();
 sg13g2_fill_1 FILLER_29_232 ();
 sg13g2_fill_2 FILLER_29_238 ();
 sg13g2_fill_1 FILLER_29_240 ();
 sg13g2_fill_1 FILLER_29_251 ();
 sg13g2_fill_2 FILLER_29_260 ();
 sg13g2_fill_1 FILLER_29_262 ();
 sg13g2_fill_2 FILLER_29_272 ();
 sg13g2_fill_1 FILLER_29_274 ();
 sg13g2_fill_2 FILLER_29_290 ();
 sg13g2_decap_4 FILLER_29_315 ();
 sg13g2_fill_1 FILLER_29_371 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_fill_1 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_fill_2 FILLER_30_154 ();
 sg13g2_fill_2 FILLER_30_165 ();
 sg13g2_fill_1 FILLER_30_167 ();
 sg13g2_fill_2 FILLER_30_173 ();
 sg13g2_fill_1 FILLER_30_179 ();
 sg13g2_fill_1 FILLER_30_224 ();
 sg13g2_fill_2 FILLER_30_281 ();
 sg13g2_fill_1 FILLER_30_283 ();
 sg13g2_decap_4 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_292 ();
 sg13g2_decap_8 FILLER_30_303 ();
 sg13g2_decap_8 FILLER_30_310 ();
 sg13g2_decap_4 FILLER_30_321 ();
 sg13g2_fill_1 FILLER_30_325 ();
 sg13g2_decap_4 FILLER_30_338 ();
 sg13g2_fill_2 FILLER_30_351 ();
 sg13g2_fill_1 FILLER_30_353 ();
 sg13g2_fill_1 FILLER_30_359 ();
 sg13g2_fill_1 FILLER_30_377 ();
 sg13g2_fill_2 FILLER_30_388 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_fill_2 FILLER_31_28 ();
 sg13g2_fill_2 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_58 ();
 sg13g2_fill_2 FILLER_31_86 ();
 sg13g2_fill_1 FILLER_31_100 ();
 sg13g2_fill_1 FILLER_31_137 ();
 sg13g2_fill_1 FILLER_31_164 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_fill_2 FILLER_31_224 ();
 sg13g2_fill_1 FILLER_31_226 ();
 sg13g2_fill_2 FILLER_31_255 ();
 sg13g2_decap_4 FILLER_31_261 ();
 sg13g2_fill_1 FILLER_31_282 ();
 sg13g2_fill_1 FILLER_31_288 ();
 sg13g2_decap_4 FILLER_31_299 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_fill_1 FILLER_32_86 ();
 sg13g2_fill_2 FILLER_32_108 ();
 sg13g2_fill_2 FILLER_32_125 ();
 sg13g2_decap_4 FILLER_32_149 ();
 sg13g2_fill_2 FILLER_32_153 ();
 sg13g2_fill_1 FILLER_32_167 ();
 sg13g2_fill_1 FILLER_32_177 ();
 sg13g2_decap_8 FILLER_32_187 ();
 sg13g2_decap_8 FILLER_32_194 ();
 sg13g2_fill_1 FILLER_32_201 ();
 sg13g2_decap_8 FILLER_32_206 ();
 sg13g2_fill_2 FILLER_32_213 ();
 sg13g2_fill_1 FILLER_32_215 ();
 sg13g2_fill_2 FILLER_32_272 ();
 sg13g2_fill_2 FILLER_32_305 ();
 sg13g2_fill_1 FILLER_32_307 ();
 sg13g2_fill_1 FILLER_32_359 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_fill_1 FILLER_33_28 ();
 sg13g2_fill_2 FILLER_33_55 ();
 sg13g2_fill_1 FILLER_33_57 ();
 sg13g2_fill_1 FILLER_33_104 ();
 sg13g2_fill_1 FILLER_33_131 ();
 sg13g2_fill_2 FILLER_33_137 ();
 sg13g2_fill_2 FILLER_33_144 ();
 sg13g2_fill_1 FILLER_33_151 ();
 sg13g2_fill_2 FILLER_33_229 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_fill_1 FILLER_33_242 ();
 sg13g2_fill_1 FILLER_33_258 ();
 sg13g2_fill_2 FILLER_33_273 ();
 sg13g2_fill_1 FILLER_33_350 ();
 sg13g2_fill_1 FILLER_33_371 ();
 sg13g2_fill_2 FILLER_33_381 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_4 FILLER_34_21 ();
 sg13g2_fill_1 FILLER_34_25 ();
 sg13g2_fill_2 FILLER_34_48 ();
 sg13g2_fill_1 FILLER_34_50 ();
 sg13g2_fill_2 FILLER_34_78 ();
 sg13g2_fill_2 FILLER_34_128 ();
 sg13g2_fill_2 FILLER_34_153 ();
 sg13g2_fill_1 FILLER_34_155 ();
 sg13g2_fill_1 FILLER_34_169 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_4 FILLER_34_203 ();
 sg13g2_fill_2 FILLER_34_207 ();
 sg13g2_fill_1 FILLER_34_213 ();
 sg13g2_fill_2 FILLER_34_223 ();
 sg13g2_fill_1 FILLER_34_225 ();
 sg13g2_fill_2 FILLER_34_242 ();
 sg13g2_decap_4 FILLER_34_250 ();
 sg13g2_fill_2 FILLER_34_311 ();
 sg13g2_fill_1 FILLER_34_317 ();
 sg13g2_fill_2 FILLER_34_352 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_fill_2 FILLER_35_92 ();
 sg13g2_fill_2 FILLER_35_145 ();
 sg13g2_decap_4 FILLER_35_164 ();
 sg13g2_fill_2 FILLER_35_201 ();
 sg13g2_fill_2 FILLER_35_238 ();
 sg13g2_fill_2 FILLER_35_249 ();
 sg13g2_fill_1 FILLER_35_265 ();
 sg13g2_decap_4 FILLER_35_292 ();
 sg13g2_fill_1 FILLER_35_308 ();
 sg13g2_fill_1 FILLER_35_318 ();
 sg13g2_fill_2 FILLER_35_343 ();
 sg13g2_fill_1 FILLER_35_345 ();
 sg13g2_fill_1 FILLER_35_360 ();
 sg13g2_fill_2 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_fill_2 FILLER_36_35 ();
 sg13g2_fill_1 FILLER_36_123 ();
 sg13g2_decap_8 FILLER_36_155 ();
 sg13g2_decap_8 FILLER_36_162 ();
 sg13g2_decap_4 FILLER_36_169 ();
 sg13g2_fill_1 FILLER_36_173 ();
 sg13g2_decap_4 FILLER_36_179 ();
 sg13g2_fill_2 FILLER_36_183 ();
 sg13g2_decap_8 FILLER_36_201 ();
 sg13g2_fill_1 FILLER_36_208 ();
 sg13g2_fill_2 FILLER_36_224 ();
 sg13g2_fill_1 FILLER_36_226 ();
 sg13g2_fill_2 FILLER_36_279 ();
 sg13g2_fill_2 FILLER_36_329 ();
 sg13g2_fill_2 FILLER_36_357 ();
 sg13g2_fill_2 FILLER_36_390 ();
 sg13g2_fill_1 FILLER_36_392 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_4 FILLER_37_49 ();
 sg13g2_fill_1 FILLER_37_53 ();
 sg13g2_fill_2 FILLER_37_69 ();
 sg13g2_fill_1 FILLER_37_71 ();
 sg13g2_fill_1 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_129 ();
 sg13g2_fill_2 FILLER_37_136 ();
 sg13g2_fill_2 FILLER_37_164 ();
 sg13g2_decap_4 FILLER_37_200 ();
 sg13g2_fill_2 FILLER_37_215 ();
 sg13g2_fill_1 FILLER_37_217 ();
 sg13g2_fill_1 FILLER_37_244 ();
 sg13g2_fill_1 FILLER_37_255 ();
 sg13g2_decap_8 FILLER_37_270 ();
 sg13g2_fill_1 FILLER_37_281 ();
 sg13g2_fill_2 FILLER_37_291 ();
 sg13g2_fill_1 FILLER_37_293 ();
 sg13g2_fill_2 FILLER_37_310 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_fill_2 FILLER_38_49 ();
 sg13g2_fill_1 FILLER_38_72 ();
 sg13g2_fill_2 FILLER_38_86 ();
 sg13g2_fill_1 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_131 ();
 sg13g2_decap_8 FILLER_38_139 ();
 sg13g2_fill_2 FILLER_38_146 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_fill_2 FILLER_38_175 ();
 sg13g2_fill_1 FILLER_38_177 ();
 sg13g2_fill_2 FILLER_38_194 ();
 sg13g2_fill_2 FILLER_38_230 ();
 sg13g2_fill_1 FILLER_38_232 ();
 sg13g2_fill_1 FILLER_38_259 ();
 sg13g2_fill_2 FILLER_38_268 ();
 sg13g2_fill_2 FILLER_38_296 ();
 sg13g2_fill_1 FILLER_38_298 ();
 assign uio_oe[0] = net150;
 assign uio_oe[1] = net151;
 assign uio_oe[2] = net152;
 assign uio_oe[3] = net153;
 assign uio_oe[4] = net154;
 assign uio_oe[5] = net155;
 assign uio_oe[6] = net156;
 assign uio_oe[7] = net157;
 assign uo_out[3] = net9;
 assign uo_out[4] = net10;
 assign uo_out[5] = net11;
 assign uo_out[6] = net12;
 assign uo_out[7] = net13;
endmodule

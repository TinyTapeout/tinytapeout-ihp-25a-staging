module tt_um_wokwi_413386991502909441 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire clk_regs;
 wire \bi_en[0] ;
 wire \bi_en[1] ;
 wire \bi_en[2] ;
 wire \bi_en[3] ;
 wire \bi_en[4] ;
 wire \bi_en[5] ;
 wire \bi_en[6] ;
 wire \bi_en[7] ;
 wire \bi_frame_index[0] ;
 wire \bi_frame_index[1] ;
 wire \bi_out[0] ;
 wire \bi_out[1] ;
 wire \bi_out[2] ;
 wire \bi_out[3] ;
 wire \bi_out[4] ;
 wire \bi_out[5] ;
 wire \bi_out[6] ;
 wire \bi_out[7] ;
 wire \charlie_0.charlie_index[0] ;
 wire \charlie_0.charlie_index[1] ;
 wire \charlie_0.charlie_index[2] ;
 wire \charlie_0.charlie_index[3] ;
 wire \charlie_0.charlie_index[4] ;
 wire \charlie_0.charlie_index[5] ;
 wire \charlie_0.is_mirror ;
 wire \charlie_0.memory[0][0] ;
 wire \charlie_0.memory[0][1] ;
 wire \charlie_0.memory[0][2] ;
 wire \charlie_0.memory[0][3] ;
 wire \charlie_0.memory[0][4] ;
 wire \charlie_0.memory[0][5] ;
 wire \charlie_0.memory[0][6] ;
 wire \charlie_0.memory[0][7] ;
 wire \charlie_0.memory[10][0] ;
 wire \charlie_0.memory[10][1] ;
 wire \charlie_0.memory[10][2] ;
 wire \charlie_0.memory[10][3] ;
 wire \charlie_0.memory[10][4] ;
 wire \charlie_0.memory[10][5] ;
 wire \charlie_0.memory[10][6] ;
 wire \charlie_0.memory[10][7] ;
 wire \charlie_0.memory[11][0] ;
 wire \charlie_0.memory[11][1] ;
 wire \charlie_0.memory[11][2] ;
 wire \charlie_0.memory[11][3] ;
 wire \charlie_0.memory[11][4] ;
 wire \charlie_0.memory[11][5] ;
 wire \charlie_0.memory[11][6] ;
 wire \charlie_0.memory[11][7] ;
 wire \charlie_0.memory[12][0] ;
 wire \charlie_0.memory[12][1] ;
 wire \charlie_0.memory[12][2] ;
 wire \charlie_0.memory[12][3] ;
 wire \charlie_0.memory[12][4] ;
 wire \charlie_0.memory[12][5] ;
 wire \charlie_0.memory[12][6] ;
 wire \charlie_0.memory[12][7] ;
 wire \charlie_0.memory[13][0] ;
 wire \charlie_0.memory[13][1] ;
 wire \charlie_0.memory[13][2] ;
 wire \charlie_0.memory[13][3] ;
 wire \charlie_0.memory[13][4] ;
 wire \charlie_0.memory[13][5] ;
 wire \charlie_0.memory[13][6] ;
 wire \charlie_0.memory[13][7] ;
 wire \charlie_0.memory[14][0] ;
 wire \charlie_0.memory[14][1] ;
 wire \charlie_0.memory[14][2] ;
 wire \charlie_0.memory[14][3] ;
 wire \charlie_0.memory[14][4] ;
 wire \charlie_0.memory[14][5] ;
 wire \charlie_0.memory[14][6] ;
 wire \charlie_0.memory[14][7] ;
 wire \charlie_0.memory[15][0] ;
 wire \charlie_0.memory[15][1] ;
 wire \charlie_0.memory[15][2] ;
 wire \charlie_0.memory[15][3] ;
 wire \charlie_0.memory[15][4] ;
 wire \charlie_0.memory[15][5] ;
 wire \charlie_0.memory[15][6] ;
 wire \charlie_0.memory[15][7] ;
 wire \charlie_0.memory[16][0] ;
 wire \charlie_0.memory[16][1] ;
 wire \charlie_0.memory[16][2] ;
 wire \charlie_0.memory[16][3] ;
 wire \charlie_0.memory[16][4] ;
 wire \charlie_0.memory[16][5] ;
 wire \charlie_0.memory[16][6] ;
 wire \charlie_0.memory[16][7] ;
 wire \charlie_0.memory[17][0] ;
 wire \charlie_0.memory[17][1] ;
 wire \charlie_0.memory[17][2] ;
 wire \charlie_0.memory[17][3] ;
 wire \charlie_0.memory[17][4] ;
 wire \charlie_0.memory[17][5] ;
 wire \charlie_0.memory[17][6] ;
 wire \charlie_0.memory[17][7] ;
 wire \charlie_0.memory[18][0] ;
 wire \charlie_0.memory[18][1] ;
 wire \charlie_0.memory[18][2] ;
 wire \charlie_0.memory[18][3] ;
 wire \charlie_0.memory[18][4] ;
 wire \charlie_0.memory[18][5] ;
 wire \charlie_0.memory[18][6] ;
 wire \charlie_0.memory[18][7] ;
 wire \charlie_0.memory[19][3] ;
 wire \charlie_0.memory[19][4] ;
 wire \charlie_0.memory[19][5] ;
 wire \charlie_0.memory[19][6] ;
 wire \charlie_0.memory[19][7] ;
 wire \charlie_0.memory[1][0] ;
 wire \charlie_0.memory[1][1] ;
 wire \charlie_0.memory[1][2] ;
 wire \charlie_0.memory[1][3] ;
 wire \charlie_0.memory[1][4] ;
 wire \charlie_0.memory[1][5] ;
 wire \charlie_0.memory[1][6] ;
 wire \charlie_0.memory[1][7] ;
 wire \charlie_0.memory[20][0] ;
 wire \charlie_0.memory[20][1] ;
 wire \charlie_0.memory[20][2] ;
 wire \charlie_0.memory[20][3] ;
 wire \charlie_0.memory[20][4] ;
 wire \charlie_0.memory[20][5] ;
 wire \charlie_0.memory[20][6] ;
 wire \charlie_0.memory[20][7] ;
 wire \charlie_0.memory[21][0] ;
 wire \charlie_0.memory[21][1] ;
 wire \charlie_0.memory[21][2] ;
 wire \charlie_0.memory[21][3] ;
 wire \charlie_0.memory[21][4] ;
 wire \charlie_0.memory[21][5] ;
 wire \charlie_0.memory[21][6] ;
 wire \charlie_0.memory[21][7] ;
 wire \charlie_0.memory[22][0] ;
 wire \charlie_0.memory[22][1] ;
 wire \charlie_0.memory[22][2] ;
 wire \charlie_0.memory[22][3] ;
 wire \charlie_0.memory[22][4] ;
 wire \charlie_0.memory[22][5] ;
 wire \charlie_0.memory[22][6] ;
 wire \charlie_0.memory[22][7] ;
 wire \charlie_0.memory[2][0] ;
 wire \charlie_0.memory[2][1] ;
 wire \charlie_0.memory[2][2] ;
 wire \charlie_0.memory[2][3] ;
 wire \charlie_0.memory[2][4] ;
 wire \charlie_0.memory[2][5] ;
 wire \charlie_0.memory[2][6] ;
 wire \charlie_0.memory[2][7] ;
 wire \charlie_0.memory[3][0] ;
 wire \charlie_0.memory[3][1] ;
 wire \charlie_0.memory[3][2] ;
 wire \charlie_0.memory[3][3] ;
 wire \charlie_0.memory[3][4] ;
 wire \charlie_0.memory[3][5] ;
 wire \charlie_0.memory[3][6] ;
 wire \charlie_0.memory[3][7] ;
 wire \charlie_0.memory[4][0] ;
 wire \charlie_0.memory[4][1] ;
 wire \charlie_0.memory[4][2] ;
 wire \charlie_0.memory[4][3] ;
 wire \charlie_0.memory[4][4] ;
 wire \charlie_0.memory[4][5] ;
 wire \charlie_0.memory[4][6] ;
 wire \charlie_0.memory[4][7] ;
 wire \charlie_0.memory[5][0] ;
 wire \charlie_0.memory[5][1] ;
 wire \charlie_0.memory[5][2] ;
 wire \charlie_0.memory[5][3] ;
 wire \charlie_0.memory[5][4] ;
 wire \charlie_0.memory[5][5] ;
 wire \charlie_0.memory[5][6] ;
 wire \charlie_0.memory[5][7] ;
 wire \charlie_0.memory[6][0] ;
 wire \charlie_0.memory[6][1] ;
 wire \charlie_0.memory[6][2] ;
 wire \charlie_0.memory[6][3] ;
 wire \charlie_0.memory[6][4] ;
 wire \charlie_0.memory[6][5] ;
 wire \charlie_0.memory[6][6] ;
 wire \charlie_0.memory[6][7] ;
 wire \charlie_0.memory[7][0] ;
 wire \charlie_0.memory[7][1] ;
 wire \charlie_0.memory[7][2] ;
 wire \charlie_0.memory[7][3] ;
 wire \charlie_0.memory[7][4] ;
 wire \charlie_0.memory[7][5] ;
 wire \charlie_0.memory[7][6] ;
 wire \charlie_0.memory[7][7] ;
 wire \charlie_0.memory[8][0] ;
 wire \charlie_0.memory[8][1] ;
 wire \charlie_0.memory[8][2] ;
 wire \charlie_0.memory[8][3] ;
 wire \charlie_0.memory[8][4] ;
 wire \charlie_0.memory[8][5] ;
 wire \charlie_0.memory[8][6] ;
 wire \charlie_0.memory[8][7] ;
 wire \charlie_0.memory[9][0] ;
 wire \charlie_0.memory[9][1] ;
 wire \charlie_0.memory[9][2] ;
 wire \charlie_0.memory[9][3] ;
 wire \charlie_0.memory[9][4] ;
 wire \charlie_0.memory[9][5] ;
 wire \charlie_0.memory[9][6] ;
 wire \charlie_0.memory[9][7] ;
 wire \counter[10] ;
 wire \counter[11] ;
 wire \counter[12] ;
 wire \counter[13] ;
 wire \counter[14] ;
 wire \counter[15] ;
 wire \counter[16] ;
 wire \counter[17] ;
 wire \counter[18] ;
 wire \counter[19] ;
 wire \counter[20] ;
 wire \counter[21] ;
 wire \counter[22] ;
 wire \counter[23] ;
 wire \counter[24] ;
 wire \counter[25] ;
 wire \counter[26] ;
 wire \counter[27] ;
 wire \counter[28] ;
 wire \counter[29] ;
 wire \counter[30] ;
 wire \counter[31] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire \gen_priority_write_blocks[0].this_priority_write.data_bits[10] ;
 wire \gen_priority_write_blocks[0].this_priority_write.data_bits[11] ;
 wire \gen_priority_write_blocks[0].this_priority_write.data_bits[12] ;
 wire \gen_priority_write_blocks[0].this_priority_write.data_bits[13] ;
 wire \gen_priority_write_blocks[0].this_priority_write.data_bits[14] ;
 wire \gen_priority_write_blocks[0].this_priority_write.data_bits[15] ;
 wire \gen_priority_write_blocks[0].this_priority_write.data_bits[9] ;
 wire miso;
 wire sig_gen_out;
 wire \signal_generator_0.index_reg[0] ;
 wire \signal_generator_0.index_reg[1] ;
 wire \signal_generator_0.index_reg[2] ;
 wire \signal_generator_0.index_reg[3] ;
 wire \signal_generator_0.index_reg[4] ;
 wire \signal_generator_0.index_reg[5] ;
 wire \signal_generator_0.index_reg[6] ;
 wire \signal_generator_0.index_reg[7] ;
 wire \signal_generator_0.prev_clk_div ;
 wire \signal_generator_0.prev_trigger ;
 wire \signal_generator_0.state_machine[0] ;
 wire \signal_generator_0.state_machine[1] ;
 wire \spi_address[0] ;
 wire \spi_address[1] ;
 wire \spi_address[2] ;
 wire \spi_address[3] ;
 wire \spi_address[4] ;
 wire \spi_slave_0.bit_cnt[0] ;
 wire \spi_slave_0.bit_cnt[1] ;
 wire \spi_slave_0.bit_cnt[2] ;
 wire \spi_slave_0.is_data_phase ;
 wire \spi_slave_0.is_mosi ;
 wire \spi_slave_0.reg_data[7] ;
 wire \spi_slave_0.spi_clk_prev ;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_leaf_0_clk_regs;
 wire clknet_leaf_1_clk_regs;
 wire clknet_leaf_2_clk_regs;
 wire clknet_leaf_3_clk_regs;
 wire clknet_leaf_4_clk_regs;
 wire clknet_leaf_5_clk_regs;
 wire clknet_leaf_6_clk_regs;
 wire clknet_leaf_7_clk_regs;
 wire clknet_leaf_8_clk_regs;
 wire clknet_leaf_9_clk_regs;
 wire clknet_leaf_10_clk_regs;
 wire clknet_leaf_11_clk_regs;
 wire clknet_leaf_12_clk_regs;
 wire clknet_leaf_13_clk_regs;
 wire clknet_leaf_14_clk_regs;
 wire clknet_leaf_15_clk_regs;
 wire clknet_leaf_16_clk_regs;
 wire clknet_leaf_17_clk_regs;
 wire clknet_leaf_18_clk_regs;
 wire clknet_leaf_19_clk_regs;
 wire clknet_leaf_20_clk_regs;
 wire clknet_leaf_21_clk_regs;
 wire clknet_leaf_22_clk_regs;
 wire clknet_leaf_24_clk_regs;
 wire clknet_leaf_25_clk_regs;
 wire clknet_leaf_26_clk_regs;
 wire clknet_leaf_27_clk_regs;
 wire clknet_leaf_28_clk_regs;
 wire clknet_leaf_29_clk_regs;
 wire clknet_leaf_30_clk_regs;
 wire clknet_leaf_31_clk_regs;
 wire clknet_leaf_32_clk_regs;
 wire clknet_leaf_33_clk_regs;
 wire clknet_leaf_34_clk_regs;
 wire clknet_leaf_35_clk_regs;
 wire clknet_0_clk_regs;
 wire clknet_3_0__leaf_clk_regs;
 wire clknet_3_1__leaf_clk_regs;
 wire clknet_3_2__leaf_clk_regs;
 wire clknet_3_3__leaf_clk_regs;
 wire clknet_3_4__leaf_clk_regs;
 wire clknet_3_5__leaf_clk_regs;
 wire clknet_3_6__leaf_clk_regs;
 wire clknet_3_7__leaf_clk_regs;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;

 sg13g2_inv_1 _2630_ (.Y(_1768_),
    .A(net1213));
 sg13g2_inv_1 _2631_ (.Y(_1769_),
    .A(net1184));
 sg13g2_inv_1 _2632_ (.Y(_1770_),
    .A(net1187));
 sg13g2_inv_1 _2633_ (.Y(_1771_),
    .A(net1189));
 sg13g2_inv_1 _2634_ (.Y(_1772_),
    .A(net1191));
 sg13g2_inv_2 _2635_ (.Y(_1773_),
    .A(net1194));
 sg13g2_inv_1 _2636_ (.Y(_1774_),
    .A(\charlie_0.memory[22][1] ));
 sg13g2_inv_4 _2637_ (.A(net1197),
    .Y(_1775_));
 sg13g2_inv_1 _2638_ (.Y(_1776_),
    .A(net1232));
 sg13g2_inv_1 _2639_ (.Y(_1777_),
    .A(\charlie_0.memory[20][3] ));
 sg13g2_inv_2 _2640_ (.Y(_1778_),
    .A(\charlie_0.memory[17][6] ));
 sg13g2_inv_4 _2641_ (.A(\charlie_0.memory[17][5] ),
    .Y(_1779_));
 sg13g2_inv_4 _2642_ (.A(\charlie_0.memory[17][4] ),
    .Y(_1780_));
 sg13g2_inv_4 _2643_ (.A(net1157),
    .Y(_1781_));
 sg13g2_inv_1 _2644_ (.Y(_1782_),
    .A(net1160));
 sg13g2_inv_1 _2645_ (.Y(_1783_),
    .A(net1161));
 sg13g2_inv_1 _2646_ (.Y(_1784_),
    .A(net1163));
 sg13g2_inv_1 _2647_ (.Y(_1785_),
    .A(net1165));
 sg13g2_inv_2 _2648_ (.Y(_1786_),
    .A(\charlie_0.memory[16][5] ));
 sg13g2_inv_1 _2649_ (.Y(_1787_),
    .A(\charlie_0.memory[16][4] ));
 sg13g2_inv_1 _2650_ (.Y(_1788_),
    .A(\charlie_0.memory[16][3] ));
 sg13g2_inv_2 _2651_ (.Y(_1789_),
    .A(\charlie_0.memory[16][2] ));
 sg13g2_inv_2 _2652_ (.Y(_1790_),
    .A(net1170));
 sg13g2_inv_1 _2653_ (.Y(_1791_),
    .A(net1173));
 sg13g2_inv_1 _2654_ (.Y(_1792_),
    .A(\charlie_0.memory[14][7] ));
 sg13g2_inv_1 _2655_ (.Y(_1793_),
    .A(\charlie_0.memory[14][6] ));
 sg13g2_inv_2 _2656_ (.Y(_1794_),
    .A(\charlie_0.memory[14][5] ));
 sg13g2_inv_1 _2657_ (.Y(_1795_),
    .A(\charlie_0.memory[14][4] ));
 sg13g2_inv_1 _2658_ (.Y(_1796_),
    .A(\charlie_0.memory[10][7] ));
 sg13g2_inv_1 _2659_ (.Y(_1797_),
    .A(\charlie_0.memory[10][6] ));
 sg13g2_inv_1 _2660_ (.Y(_1798_),
    .A(\charlie_0.memory[10][5] ));
 sg13g2_inv_1 _2661_ (.Y(_1799_),
    .A(\charlie_0.memory[10][3] ));
 sg13g2_inv_1 _2662_ (.Y(_1800_),
    .A(\charlie_0.memory[10][2] ));
 sg13g2_inv_1 _2663_ (.Y(_1801_),
    .A(\charlie_0.memory[10][1] ));
 sg13g2_inv_1 _2664_ (.Y(_1802_),
    .A(\charlie_0.memory[10][0] ));
 sg13g2_inv_1 _2665_ (.Y(_1803_),
    .A(\charlie_0.memory[7][7] ));
 sg13g2_inv_1 _2666_ (.Y(_1804_),
    .A(\charlie_0.memory[7][6] ));
 sg13g2_inv_1 _2667_ (.Y(_1805_),
    .A(\charlie_0.memory[7][5] ));
 sg13g2_inv_1 _2668_ (.Y(_1806_),
    .A(\charlie_0.memory[6][6] ));
 sg13g2_inv_1 _2669_ (.Y(_1807_),
    .A(\charlie_0.memory[5][7] ));
 sg13g2_inv_1 _2670_ (.Y(_1808_),
    .A(\charlie_0.memory[4][6] ));
 sg13g2_inv_1 _2671_ (.Y(_1809_),
    .A(\charlie_0.memory[4][5] ));
 sg13g2_inv_1 _2672_ (.Y(_1810_),
    .A(\charlie_0.memory[3][7] ));
 sg13g2_inv_1 _2673_ (.Y(_1811_),
    .A(\charlie_0.memory[2][7] ));
 sg13g2_inv_1 _2674_ (.Y(_1812_),
    .A(\charlie_0.memory[2][6] ));
 sg13g2_inv_1 _2675_ (.Y(_1813_),
    .A(\charlie_0.memory[2][5] ));
 sg13g2_inv_1 _2676_ (.Y(_1814_),
    .A(\charlie_0.memory[2][4] ));
 sg13g2_inv_1 _2677_ (.Y(_1815_),
    .A(\charlie_0.memory[1][7] ));
 sg13g2_inv_1 _2678_ (.Y(_1816_),
    .A(\charlie_0.memory[1][6] ));
 sg13g2_inv_1 _2679_ (.Y(_1817_),
    .A(\charlie_0.memory[0][4] ));
 sg13g2_inv_1 _2680_ (.Y(_1818_),
    .A(\signal_generator_0.index_reg[6] ));
 sg13g2_inv_2 _2681_ (.Y(_1819_),
    .A(\signal_generator_0.index_reg[5] ));
 sg13g2_inv_2 _2682_ (.Y(_1820_),
    .A(net1176));
 sg13g2_inv_2 _2683_ (.Y(_1821_),
    .A(\signal_generator_0.index_reg[3] ));
 sg13g2_inv_1 _2684_ (.Y(_1822_),
    .A(net1179));
 sg13g2_inv_1 _2685_ (.Y(_1823_),
    .A(net284));
 sg13g2_inv_1 _2686_ (.Y(_1824_),
    .A(net286));
 sg13g2_inv_1 _2687_ (.Y(_1825_),
    .A(\spi_slave_0.spi_clk_prev ));
 sg13g2_inv_1 _2688_ (.Y(_1826_),
    .A(net1211));
 sg13g2_inv_1 _2689_ (.Y(_1827_),
    .A(net1210));
 sg13g2_inv_2 _2690_ (.Y(_1828_),
    .A(net1208));
 sg13g2_inv_1 _2691_ (.Y(_1829_),
    .A(net493));
 sg13g2_inv_1 _2692_ (.Y(_1830_),
    .A(net360));
 sg13g2_inv_1 _2693_ (.Y(_1831_),
    .A(net465));
 sg13g2_inv_1 _2694_ (.Y(_1832_),
    .A(\counter[28] ));
 sg13g2_inv_1 _2695_ (.Y(_1833_),
    .A(\counter[29] ));
 sg13g2_inv_1 _2696_ (.Y(_1834_),
    .A(\signal_generator_0.state_machine[0] ));
 sg13g2_inv_1 _2697_ (.Y(_1835_),
    .A(net1237));
 sg13g2_inv_1 _2698_ (.Y(_1836_),
    .A(_0050_));
 sg13g2_inv_1 _2699_ (.Y(_1837_),
    .A(_0053_));
 sg13g2_nor2_1 _2700_ (.A(\charlie_0.memory[16][7] ),
    .B(net1222),
    .Y(_1838_));
 sg13g2_nand2b_1 _2701_ (.Y(_1839_),
    .B(net1234),
    .A_N(\charlie_0.memory[16][7] ));
 sg13g2_nand2_1 _2702_ (.Y(_1840_),
    .A(net1167),
    .B(net1112));
 sg13g2_xnor2_1 _2703_ (.Y(_1841_),
    .A(net1209),
    .B(\counter[21] ));
 sg13g2_o21ai_1 _2704_ (.B1(net1167),
    .Y(_1842_),
    .A1(\counter[31] ),
    .A2(_1841_));
 sg13g2_a21oi_1 _2705_ (.A1(\counter[31] ),
    .A2(_1841_),
    .Y(_1843_),
    .B1(_1842_));
 sg13g2_and2_1 _2706_ (.A(net295),
    .B(_1843_),
    .X(_1844_));
 sg13g2_a21oi_1 _2707_ (.A1(net295),
    .A2(_1838_),
    .Y(_1845_),
    .B1(_1843_));
 sg13g2_o21ai_1 _2708_ (.B1(_1840_),
    .Y(_0016_),
    .A1(_1844_),
    .A2(_1845_));
 sg13g2_nor2_2 _2709_ (.A(net1211),
    .B(net1210),
    .Y(_1846_));
 sg13g2_nand2_2 _2710_ (.Y(_1847_),
    .A(net1211),
    .B(net1209));
 sg13g2_nand2b_1 _2711_ (.Y(_1848_),
    .B(_1847_),
    .A_N(_1846_));
 sg13g2_nor2_2 _2712_ (.A(net1165),
    .B(net1106),
    .Y(_1849_));
 sg13g2_nand2b_1 _2713_ (.Y(_1850_),
    .B(net1119),
    .A_N(net1106));
 sg13g2_o21ai_1 _2714_ (.B1(net1167),
    .Y(_1851_),
    .A1(net1211),
    .A2(net1112));
 sg13g2_o21ai_1 _2715_ (.B1(_1851_),
    .Y(_0027_),
    .A1(_1848_),
    .A2(net1028));
 sg13g2_and3_1 _2716_ (.X(_1852_),
    .A(net1211),
    .B(net1209),
    .C(net1208));
 sg13g2_xnor2_1 _2717_ (.Y(_1853_),
    .A(net1208),
    .B(_1847_));
 sg13g2_a22oi_1 _2718_ (.Y(_1854_),
    .B1(_1849_),
    .B2(_1853_),
    .A2(net1209),
    .A1(net1167));
 sg13g2_nand2_1 _2719_ (.Y(_0038_),
    .A(_1840_),
    .B(_1854_));
 sg13g2_nor2_1 _2720_ (.A(net307),
    .B(_1847_),
    .Y(_1855_));
 sg13g2_xnor2_1 _2721_ (.Y(_1856_),
    .A(net1205),
    .B(_1855_));
 sg13g2_o21ai_1 _2722_ (.B1(net1167),
    .Y(_1857_),
    .A1(net1207),
    .A2(net1112));
 sg13g2_o21ai_1 _2723_ (.B1(_1857_),
    .Y(_0041_),
    .A1(net1028),
    .A2(_1856_));
 sg13g2_nor2_2 _2724_ (.A(net1205),
    .B(net1203),
    .Y(_1858_));
 sg13g2_a21oi_1 _2725_ (.A1(net1205),
    .A2(_1852_),
    .Y(_1859_),
    .B1(net1203));
 sg13g2_and2_2 _2726_ (.A(net1205),
    .B(net1203),
    .X(_1860_));
 sg13g2_nand2_2 _2727_ (.Y(_1861_),
    .A(net1206),
    .B(net1204));
 sg13g2_and2_1 _2728_ (.A(_1852_),
    .B(_1860_),
    .X(_1862_));
 sg13g2_nor3_1 _2729_ (.A(net1028),
    .B(_1859_),
    .C(_1862_),
    .Y(_1863_));
 sg13g2_o21ai_1 _2730_ (.B1(net1167),
    .Y(_1864_),
    .A1(net1205),
    .A2(net1112));
 sg13g2_nand2b_1 _2731_ (.Y(_0042_),
    .B(_1864_),
    .A_N(_1863_));
 sg13g2_and2_1 _2732_ (.A(net1201),
    .B(_1862_),
    .X(_1865_));
 sg13g2_o21ai_1 _2733_ (.B1(_1849_),
    .Y(_1866_),
    .A1(net1201),
    .A2(_1862_));
 sg13g2_o21ai_1 _2734_ (.B1(net1167),
    .Y(_1867_),
    .A1(net1203),
    .A2(net1112));
 sg13g2_o21ai_1 _2735_ (.B1(_1867_),
    .Y(_0043_),
    .A1(_1865_),
    .A2(_1866_));
 sg13g2_nand4_1 _2736_ (.B(\counter[6] ),
    .C(_1852_),
    .A(net1201),
    .Y(_1868_),
    .D(_1860_));
 sg13g2_nor2_1 _2737_ (.A(net355),
    .B(_1865_),
    .Y(_1869_));
 sg13g2_nor2_1 _2738_ (.A(net1028),
    .B(_1869_),
    .Y(_1870_));
 sg13g2_a22oi_1 _2739_ (.Y(_1871_),
    .B1(_1868_),
    .B2(_1870_),
    .A2(net1201),
    .A1(net1167));
 sg13g2_nand2_1 _2740_ (.Y(_0044_),
    .A(_1840_),
    .B(_1871_));
 sg13g2_or2_1 _2741_ (.X(_1872_),
    .B(_1868_),
    .A(_1829_));
 sg13g2_xnor2_1 _2742_ (.Y(_1873_),
    .A(_1829_),
    .B(_1868_));
 sg13g2_o21ai_1 _2743_ (.B1(net1166),
    .Y(_1874_),
    .A1(net355),
    .A2(net1107));
 sg13g2_o21ai_1 _2744_ (.B1(_1874_),
    .Y(_0045_),
    .A1(net1028),
    .A2(_1873_));
 sg13g2_nor2_1 _2745_ (.A(net333),
    .B(net1109),
    .Y(_1875_));
 sg13g2_a21oi_2 _2746_ (.B1(_1875_),
    .Y(_1876_),
    .A2(_1872_),
    .A1(_1849_));
 sg13g2_nor2_1 _2747_ (.A(net1166),
    .B(_1872_),
    .Y(_1877_));
 sg13g2_nor2_1 _2748_ (.A(net333),
    .B(_1877_),
    .Y(_1878_));
 sg13g2_o21ai_1 _2749_ (.B1(net1166),
    .Y(_1879_),
    .A1(\counter[7] ),
    .A2(net1111));
 sg13g2_o21ai_1 _2750_ (.B1(_1879_),
    .Y(_0046_),
    .A1(_1876_),
    .A2(_1878_));
 sg13g2_o21ai_1 _2751_ (.B1(net1120),
    .Y(_1880_),
    .A1(net472),
    .A2(net1109));
 sg13g2_xnor2_1 _2752_ (.Y(_0047_),
    .A(_1876_),
    .B(_1880_));
 sg13g2_o21ai_1 _2753_ (.B1(net1166),
    .Y(_1881_),
    .A1(\counter[9] ),
    .A2(net1109));
 sg13g2_nand2_1 _2754_ (.Y(_1882_),
    .A(\counter[8] ),
    .B(\counter[9] ));
 sg13g2_nor2_1 _2755_ (.A(_1872_),
    .B(_1882_),
    .Y(_1883_));
 sg13g2_nor2_1 _2756_ (.A(net376),
    .B(_1883_),
    .Y(_1884_));
 sg13g2_a21o_1 _2757_ (.A2(_1883_),
    .A1(\counter[10] ),
    .B1(net1027),
    .X(_1885_));
 sg13g2_o21ai_1 _2758_ (.B1(_1881_),
    .Y(_0017_),
    .A1(net377),
    .A2(_1885_));
 sg13g2_o21ai_1 _2759_ (.B1(net1120),
    .Y(_1886_),
    .A1(net486),
    .A2(net1110));
 sg13g2_o21ai_1 _2760_ (.B1(_1885_),
    .Y(_1887_),
    .A1(net376),
    .A2(net1109));
 sg13g2_xor2_1 _2761_ (.B(_1887_),
    .A(_1886_),
    .X(_0018_));
 sg13g2_nand2_1 _2762_ (.Y(_1888_),
    .A(\counter[10] ),
    .B(\counter[11] ));
 sg13g2_nor4_2 _2763_ (.A(_1829_),
    .B(_1868_),
    .C(_1882_),
    .Y(_1889_),
    .D(_1888_));
 sg13g2_nor2_1 _2764_ (.A(\counter[12] ),
    .B(_1889_),
    .Y(_1890_));
 sg13g2_a21o_1 _2765_ (.A2(_1889_),
    .A1(\counter[12] ),
    .B1(net1027),
    .X(_1891_));
 sg13g2_o21ai_1 _2766_ (.B1(net1169),
    .Y(_1892_),
    .A1(\counter[11] ),
    .A2(net1109));
 sg13g2_o21ai_1 _2767_ (.B1(net344),
    .Y(_0019_),
    .A1(_1890_),
    .A2(_1891_));
 sg13g2_o21ai_1 _2768_ (.B1(net1120),
    .Y(_1893_),
    .A1(net347),
    .A2(net1109));
 sg13g2_o21ai_1 _2769_ (.B1(_1891_),
    .Y(_1894_),
    .A1(net476),
    .A2(net1110));
 sg13g2_xor2_1 _2770_ (.B(_1894_),
    .A(_1893_),
    .X(_0020_));
 sg13g2_nand3_1 _2771_ (.B(\counter[13] ),
    .C(_1889_),
    .A(\counter[12] ),
    .Y(_1895_));
 sg13g2_and2_1 _2772_ (.A(_1830_),
    .B(_1895_),
    .X(_1896_));
 sg13g2_o21ai_1 _2773_ (.B1(_1849_),
    .Y(_1897_),
    .A1(_1830_),
    .A2(_1895_));
 sg13g2_o21ai_1 _2774_ (.B1(net1169),
    .Y(_1898_),
    .A1(net347),
    .A2(net1110));
 sg13g2_o21ai_1 _2775_ (.B1(_1898_),
    .Y(_0021_),
    .A1(_1896_),
    .A2(_1897_));
 sg13g2_nor2_1 _2776_ (.A(net419),
    .B(net1109),
    .Y(_1899_));
 sg13g2_nor2_1 _2777_ (.A(net1169),
    .B(_1899_),
    .Y(_1900_));
 sg13g2_o21ai_1 _2778_ (.B1(_1897_),
    .Y(_1901_),
    .A1(net360),
    .A2(net1109));
 sg13g2_xnor2_1 _2779_ (.Y(_0022_),
    .A(_1900_),
    .B(_1901_));
 sg13g2_nor2_1 _2780_ (.A(net1120),
    .B(_1899_),
    .Y(_1902_));
 sg13g2_and2_1 _2781_ (.A(\counter[14] ),
    .B(\counter[15] ),
    .X(_1903_));
 sg13g2_nand4_1 _2782_ (.B(\counter[13] ),
    .C(_1889_),
    .A(\counter[12] ),
    .Y(_1904_),
    .D(_1903_));
 sg13g2_nand2_1 _2783_ (.Y(_1905_),
    .A(_1831_),
    .B(_1904_));
 sg13g2_nor2_1 _2784_ (.A(_1831_),
    .B(_1904_),
    .Y(_1906_));
 sg13g2_nor2_1 _2785_ (.A(net1027),
    .B(_1906_),
    .Y(_1907_));
 sg13g2_a21o_1 _2786_ (.A2(_1907_),
    .A1(_1905_),
    .B1(_1902_),
    .X(_0023_));
 sg13g2_o21ai_1 _2787_ (.B1(net1120),
    .Y(_1908_),
    .A1(\counter[17] ),
    .A2(net1107));
 sg13g2_nor2_1 _2788_ (.A(net465),
    .B(net1111),
    .Y(_1909_));
 sg13g2_nor2_1 _2789_ (.A(_1907_),
    .B(_1909_),
    .Y(_1910_));
 sg13g2_xnor2_1 _2790_ (.Y(_0024_),
    .A(_1908_),
    .B(_1910_));
 sg13g2_a21oi_1 _2791_ (.A1(\counter[17] ),
    .A2(_1906_),
    .Y(_1911_),
    .B1(net403));
 sg13g2_nand3_1 _2792_ (.B(\counter[18] ),
    .C(_1906_),
    .A(\counter[17] ),
    .Y(_1912_));
 sg13g2_nand2_1 _2793_ (.Y(_1913_),
    .A(_1849_),
    .B(_1912_));
 sg13g2_o21ai_1 _2794_ (.B1(net1166),
    .Y(_1914_),
    .A1(\counter[17] ),
    .A2(net1107));
 sg13g2_o21ai_1 _2795_ (.B1(_1914_),
    .Y(_0025_),
    .A1(net404),
    .A2(_1913_));
 sg13g2_nor2_1 _2796_ (.A(\counter[19] ),
    .B(net1107),
    .Y(_1915_));
 sg13g2_nor2_1 _2797_ (.A(net1165),
    .B(_1915_),
    .Y(_1916_));
 sg13g2_o21ai_1 _2798_ (.B1(_1913_),
    .Y(_1917_),
    .A1(net482),
    .A2(net1107));
 sg13g2_xnor2_1 _2799_ (.Y(_0026_),
    .A(_1916_),
    .B(_1917_));
 sg13g2_nand4_1 _2800_ (.B(\counter[17] ),
    .C(\counter[18] ),
    .A(\counter[16] ),
    .Y(_1918_),
    .D(\counter[19] ));
 sg13g2_nor2_1 _2801_ (.A(_1904_),
    .B(_1918_),
    .Y(_1919_));
 sg13g2_a21oi_1 _2802_ (.A1(net488),
    .A2(_1919_),
    .Y(_1920_),
    .B1(net1027));
 sg13g2_o21ai_1 _2803_ (.B1(_1920_),
    .Y(_1921_),
    .A1(net408),
    .A2(_1919_));
 sg13g2_o21ai_1 _2804_ (.B1(net409),
    .Y(_0028_),
    .A1(net1119),
    .A2(_1915_));
 sg13g2_nor2_1 _2805_ (.A(\counter[21] ),
    .B(net1106),
    .Y(_1922_));
 sg13g2_nor2_1 _2806_ (.A(net1165),
    .B(_1922_),
    .Y(_1923_));
 sg13g2_nor2_1 _2807_ (.A(net408),
    .B(net1108),
    .Y(_1924_));
 sg13g2_nor2_1 _2808_ (.A(_1920_),
    .B(_1924_),
    .Y(_1925_));
 sg13g2_xor2_1 _2809_ (.B(_1925_),
    .A(_1923_),
    .X(_0029_));
 sg13g2_nand2_1 _2810_ (.Y(_1926_),
    .A(net488),
    .B(\counter[21] ));
 sg13g2_nor3_1 _2811_ (.A(_1904_),
    .B(_1918_),
    .C(_1926_),
    .Y(_1927_));
 sg13g2_a21oi_1 _2812_ (.A1(\counter[22] ),
    .A2(_1927_),
    .Y(_1928_),
    .B1(net1027));
 sg13g2_o21ai_1 _2813_ (.B1(_1928_),
    .Y(_1929_),
    .A1(net421),
    .A2(_1927_));
 sg13g2_o21ai_1 _2814_ (.B1(_1929_),
    .Y(_0030_),
    .A1(net1119),
    .A2(_1922_));
 sg13g2_nor2_1 _2815_ (.A(net379),
    .B(net1106),
    .Y(_1930_));
 sg13g2_nor2_1 _2816_ (.A(net1165),
    .B(_1930_),
    .Y(_1931_));
 sg13g2_nor2_1 _2817_ (.A(\counter[22] ),
    .B(net1106),
    .Y(_1932_));
 sg13g2_or2_1 _2818_ (.X(_1933_),
    .B(_1932_),
    .A(_1928_));
 sg13g2_xnor2_1 _2819_ (.Y(_0031_),
    .A(_1931_),
    .B(_1933_));
 sg13g2_nand2_1 _2820_ (.Y(_1934_),
    .A(\counter[22] ),
    .B(\counter[23] ));
 sg13g2_nor4_2 _2821_ (.A(_1904_),
    .B(_1918_),
    .C(_1926_),
    .Y(_1935_),
    .D(_1934_));
 sg13g2_a21oi_1 _2822_ (.A1(net496),
    .A2(_1935_),
    .Y(_1936_),
    .B1(net1027));
 sg13g2_o21ai_1 _2823_ (.B1(_1936_),
    .Y(_1937_),
    .A1(\counter[24] ),
    .A2(_1935_));
 sg13g2_o21ai_1 _2824_ (.B1(_1937_),
    .Y(_0032_),
    .A1(net1119),
    .A2(_1930_));
 sg13g2_nor2_1 _2825_ (.A(net353),
    .B(net1106),
    .Y(_1938_));
 sg13g2_nor2_1 _2826_ (.A(net1165),
    .B(_1938_),
    .Y(_1939_));
 sg13g2_nor2_1 _2827_ (.A(net487),
    .B(net1106),
    .Y(_1940_));
 sg13g2_nor2_1 _2828_ (.A(_1936_),
    .B(_1940_),
    .Y(_1941_));
 sg13g2_xor2_1 _2829_ (.B(_1941_),
    .A(_1939_),
    .X(_0033_));
 sg13g2_and3_1 _2830_ (.X(_1942_),
    .A(\counter[24] ),
    .B(\counter[25] ),
    .C(_1935_));
 sg13g2_a21oi_1 _2831_ (.A1(\counter[26] ),
    .A2(_1942_),
    .Y(_1943_),
    .B1(net1027));
 sg13g2_o21ai_1 _2832_ (.B1(_1943_),
    .Y(_1944_),
    .A1(\counter[26] ),
    .A2(_1942_));
 sg13g2_o21ai_1 _2833_ (.B1(_1944_),
    .Y(_0034_),
    .A1(net1119),
    .A2(_1938_));
 sg13g2_o21ai_1 _2834_ (.B1(net1119),
    .Y(_1945_),
    .A1(net396),
    .A2(net1107));
 sg13g2_nor2_1 _2835_ (.A(\counter[26] ),
    .B(net1106),
    .Y(_1946_));
 sg13g2_nor2_1 _2836_ (.A(_1943_),
    .B(_1946_),
    .Y(_1947_));
 sg13g2_xnor2_1 _2837_ (.Y(_0035_),
    .A(_1945_),
    .B(_1947_));
 sg13g2_nand3_1 _2838_ (.B(\counter[27] ),
    .C(_1942_),
    .A(\counter[26] ),
    .Y(_1948_));
 sg13g2_and2_1 _2839_ (.A(_1832_),
    .B(_1948_),
    .X(_1949_));
 sg13g2_o21ai_1 _2840_ (.B1(_1849_),
    .Y(_1950_),
    .A1(_1832_),
    .A2(_1948_));
 sg13g2_o21ai_1 _2841_ (.B1(net1165),
    .Y(_1951_),
    .A1(net396),
    .A2(net1107));
 sg13g2_o21ai_1 _2842_ (.B1(_1951_),
    .Y(_0036_),
    .A1(_1949_),
    .A2(_1950_));
 sg13g2_o21ai_1 _2843_ (.B1(net1119),
    .Y(_1952_),
    .A1(net369),
    .A2(net1108));
 sg13g2_o21ai_1 _2844_ (.B1(_1950_),
    .Y(_1953_),
    .A1(net406),
    .A2(net1108));
 sg13g2_xor2_1 _2845_ (.B(_1953_),
    .A(_1952_),
    .X(_0037_));
 sg13g2_o21ai_1 _2846_ (.B1(net1165),
    .Y(_1954_),
    .A1(net369),
    .A2(net1108));
 sg13g2_nor3_2 _2847_ (.A(_1832_),
    .B(_1833_),
    .C(_1948_),
    .Y(_1955_));
 sg13g2_and2_1 _2848_ (.A(\counter[30] ),
    .B(_1955_),
    .X(_1956_));
 sg13g2_o21ai_1 _2849_ (.B1(_1849_),
    .Y(_1957_),
    .A1(\counter[30] ),
    .A2(_1955_));
 sg13g2_o21ai_1 _2850_ (.B1(_1954_),
    .Y(_0039_),
    .A1(_1956_),
    .A2(_1957_));
 sg13g2_o21ai_1 _2851_ (.B1(net1119),
    .Y(_1958_),
    .A1(\counter[31] ),
    .A2(net1108));
 sg13g2_or2_1 _2852_ (.X(_1959_),
    .B(net1108),
    .A(\counter[30] ));
 sg13g2_o21ai_1 _2853_ (.B1(_1959_),
    .Y(_1960_),
    .A1(net1027),
    .A2(_1955_));
 sg13g2_xor2_1 _2854_ (.B(_1960_),
    .A(_1958_),
    .X(_0040_));
 sg13g2_xnor2_1 _2855_ (.Y(_1961_),
    .A(\charlie_0.memory[22][5] ),
    .B(net5));
 sg13g2_xor2_1 _2856_ (.B(net5),
    .A(\charlie_0.memory[22][5] ),
    .X(_1962_));
 sg13g2_xnor2_1 _2857_ (.Y(_1963_),
    .A(\charlie_0.memory[22][4] ),
    .B(net4));
 sg13g2_xor2_1 _2858_ (.B(net4),
    .A(\charlie_0.memory[22][4] ),
    .X(_1964_));
 sg13g2_nand2_2 _2859_ (.Y(_1965_),
    .A(_1962_),
    .B(_1963_));
 sg13g2_xnor2_1 _2860_ (.Y(_1966_),
    .A(\charlie_0.memory[22][7] ),
    .B(net7));
 sg13g2_xor2_1 _2861_ (.B(net7),
    .A(\charlie_0.memory[22][7] ),
    .X(_1967_));
 sg13g2_xnor2_1 _2862_ (.Y(_1968_),
    .A(\charlie_0.memory[22][6] ),
    .B(net6));
 sg13g2_xor2_1 _2863_ (.B(net6),
    .A(\charlie_0.memory[22][6] ),
    .X(_1969_));
 sg13g2_nand2_2 _2864_ (.Y(_1970_),
    .A(_1967_),
    .B(_1969_));
 sg13g2_nor2_2 _2865_ (.A(_1965_),
    .B(_1970_),
    .Y(_1971_));
 sg13g2_nand2_2 _2866_ (.Y(_1972_),
    .A(_1967_),
    .B(_1968_));
 sg13g2_nor2_2 _2867_ (.A(_1965_),
    .B(_1972_),
    .Y(_1973_));
 sg13g2_nand2_2 _2868_ (.Y(_1974_),
    .A(_1961_),
    .B(_1963_));
 sg13g2_nor2_2 _2869_ (.A(_1972_),
    .B(_1974_),
    .Y(_1975_));
 sg13g2_nand2_2 _2870_ (.Y(_1976_),
    .A(_1961_),
    .B(_1964_));
 sg13g2_nor2_2 _2871_ (.A(_1970_),
    .B(_1976_),
    .Y(_1977_));
 sg13g2_nand2_2 _2872_ (.Y(_1978_),
    .A(_1966_),
    .B(_1968_));
 sg13g2_nor2_1 _2873_ (.A(_1974_),
    .B(_1978_),
    .Y(_1979_));
 sg13g2_nand2_2 _2874_ (.Y(_1980_),
    .A(_1962_),
    .B(_1964_));
 sg13g2_nor2_2 _2875_ (.A(_1970_),
    .B(_1980_),
    .Y(_1981_));
 sg13g2_nand2_2 _2876_ (.Y(_1982_),
    .A(_1966_),
    .B(_1969_));
 sg13g2_nor2_2 _2877_ (.A(_1965_),
    .B(_1982_),
    .Y(_1983_));
 sg13g2_nor2_2 _2878_ (.A(_1976_),
    .B(_1982_),
    .Y(_1984_));
 sg13g2_nor2_2 _2879_ (.A(_1974_),
    .B(_1982_),
    .Y(_1985_));
 sg13g2_nor2_2 _2880_ (.A(_1970_),
    .B(_1974_),
    .Y(_1986_));
 sg13g2_nor2_2 _2881_ (.A(_1965_),
    .B(_1978_),
    .Y(_1987_));
 sg13g2_nor2_2 _2882_ (.A(_1972_),
    .B(_1976_),
    .Y(_1988_));
 sg13g2_nor2_2 _2883_ (.A(_1976_),
    .B(_1978_),
    .Y(_1989_));
 sg13g2_nor2_2 _2884_ (.A(_1978_),
    .B(_1980_),
    .Y(_1990_));
 sg13g2_nor2_2 _2885_ (.A(_1980_),
    .B(_1982_),
    .Y(_1991_));
 sg13g2_nor2_2 _2886_ (.A(_1972_),
    .B(_1980_),
    .Y(_1992_));
 sg13g2_a22oi_1 _2887_ (.Y(_1993_),
    .B1(_1981_),
    .B2(\charlie_0.memory[15][0] ),
    .A2(_1977_),
    .A1(\charlie_0.memory[13][0] ));
 sg13g2_a22oi_1 _2888_ (.Y(_1994_),
    .B1(_1987_),
    .B2(\charlie_0.memory[2][0] ),
    .A2(_1971_),
    .A1(\charlie_0.memory[14][0] ));
 sg13g2_a22oi_1 _2889_ (.Y(_1995_),
    .B1(_1990_),
    .B2(\charlie_0.memory[3][0] ),
    .A2(_1988_),
    .A1(\charlie_0.memory[9][0] ));
 sg13g2_a21oi_1 _2890_ (.A1(\charlie_0.memory[6][0] ),
    .A2(_1983_),
    .Y(_1996_),
    .B1(net1022));
 sg13g2_nand3_1 _2891_ (.B(_1995_),
    .C(_1996_),
    .A(_1994_),
    .Y(_1997_));
 sg13g2_a221oi_1 _2892_ (.B2(\charlie_0.memory[1][0] ),
    .C1(_1997_),
    .B1(_1989_),
    .A1(\charlie_0.memory[8][0] ),
    .Y(_1998_),
    .A2(_1975_));
 sg13g2_a22oi_1 _2893_ (.Y(_1999_),
    .B1(_1986_),
    .B2(\charlie_0.memory[12][0] ),
    .A2(_1984_),
    .A1(\charlie_0.memory[5][0] ));
 sg13g2_a22oi_1 _2894_ (.Y(_2000_),
    .B1(_1992_),
    .B2(\charlie_0.memory[11][0] ),
    .A2(_1973_),
    .A1(\charlie_0.memory[10][0] ));
 sg13g2_nand3_1 _2895_ (.B(_1999_),
    .C(_2000_),
    .A(_1993_),
    .Y(_2001_));
 sg13g2_a221oi_1 _2896_ (.B2(\charlie_0.memory[7][0] ),
    .C1(_2001_),
    .B1(_1991_),
    .A1(\charlie_0.memory[4][0] ),
    .Y(_2002_),
    .A2(_1985_));
 sg13g2_and2_1 _2897_ (.A(\charlie_0.memory[22][1] ),
    .B(_0056_),
    .X(_2003_));
 sg13g2_nand2b_1 _2898_ (.Y(_2004_),
    .B(\charlie_0.memory[22][0] ),
    .A_N(_2003_));
 sg13g2_a221oi_1 _2899_ (.B2(_2002_),
    .C1(_2004_),
    .B1(_1998_),
    .A1(_0055_),
    .Y(_2005_),
    .A2(net1022));
 sg13g2_nor2_1 _2900_ (.A(\charlie_0.memory[22][1] ),
    .B(net1146),
    .Y(_2006_));
 sg13g2_nor2_1 _2901_ (.A(\signal_generator_0.state_machine[0] ),
    .B(\signal_generator_0.state_machine[1] ),
    .Y(_2007_));
 sg13g2_or2_1 _2902_ (.X(_2008_),
    .B(\signal_generator_0.state_machine[1] ),
    .A(\signal_generator_0.state_machine[0] ));
 sg13g2_nor2_1 _2903_ (.A(_1774_),
    .B(net1146),
    .Y(_2009_));
 sg13g2_a221oi_1 _2904_ (.B2(_2009_),
    .C1(_2005_),
    .B1(_2008_),
    .A1(net2),
    .Y(_2010_),
    .A2(_2006_));
 sg13g2_xor2_1 _2905_ (.B(_2010_),
    .A(_0052_),
    .X(uo_out[0]));
 sg13g2_nand2_1 _2906_ (.Y(_2011_),
    .A(_0057_),
    .B(net1022));
 sg13g2_a22oi_1 _2907_ (.Y(_2012_),
    .B1(_1988_),
    .B2(\charlie_0.memory[9][1] ),
    .A2(_1971_),
    .A1(\charlie_0.memory[14][1] ));
 sg13g2_a22oi_1 _2908_ (.Y(_2013_),
    .B1(_1989_),
    .B2(\charlie_0.memory[1][1] ),
    .A2(_1981_),
    .A1(\charlie_0.memory[15][1] ));
 sg13g2_a22oi_1 _2909_ (.Y(_2014_),
    .B1(_1987_),
    .B2(\charlie_0.memory[2][1] ),
    .A2(_1984_),
    .A1(\charlie_0.memory[5][1] ));
 sg13g2_a21oi_1 _2910_ (.A1(\charlie_0.memory[11][1] ),
    .A2(_1992_),
    .Y(_2015_),
    .B1(net1022));
 sg13g2_nand4_1 _2911_ (.B(_2013_),
    .C(_2014_),
    .A(_2012_),
    .Y(_2016_),
    .D(_2015_));
 sg13g2_a22oi_1 _2912_ (.Y(_2017_),
    .B1(_1991_),
    .B2(\charlie_0.memory[7][1] ),
    .A2(_1977_),
    .A1(\charlie_0.memory[13][1] ));
 sg13g2_a22oi_1 _2913_ (.Y(_2018_),
    .B1(_1986_),
    .B2(\charlie_0.memory[12][1] ),
    .A2(_1985_),
    .A1(\charlie_0.memory[4][1] ));
 sg13g2_a22oi_1 _2914_ (.Y(_2019_),
    .B1(_1983_),
    .B2(\charlie_0.memory[6][1] ),
    .A2(_1975_),
    .A1(\charlie_0.memory[8][1] ));
 sg13g2_a22oi_1 _2915_ (.Y(_2020_),
    .B1(_1990_),
    .B2(\charlie_0.memory[3][1] ),
    .A2(_1973_),
    .A1(\charlie_0.memory[10][1] ));
 sg13g2_nand4_1 _2916_ (.B(_2018_),
    .C(_2019_),
    .A(_2017_),
    .Y(_2021_),
    .D(_2020_));
 sg13g2_o21ai_1 _2917_ (.B1(_2011_),
    .Y(_2022_),
    .A1(_2016_),
    .A2(_2021_));
 sg13g2_a221oi_1 _2918_ (.B2(net1146),
    .C1(_2003_),
    .B1(_2022_),
    .A1(net1228),
    .Y(_2023_),
    .A2(net1105));
 sg13g2_xnor2_1 _2919_ (.Y(uo_out[1]),
    .A(_0052_),
    .B(_2023_));
 sg13g2_o21ai_1 _2920_ (.B1(\charlie_0.memory[22][1] ),
    .Y(_2024_),
    .A1(_0056_),
    .A2(_0054_));
 sg13g2_a22oi_1 _2921_ (.Y(_2025_),
    .B1(_1990_),
    .B2(\charlie_0.memory[3][2] ),
    .A2(_1985_),
    .A1(\charlie_0.memory[4][2] ));
 sg13g2_a22oi_1 _2922_ (.Y(_2026_),
    .B1(_1989_),
    .B2(\charlie_0.memory[1][2] ),
    .A2(_1986_),
    .A1(\charlie_0.memory[12][2] ));
 sg13g2_a22oi_1 _2923_ (.Y(_2027_),
    .B1(_1992_),
    .B2(\charlie_0.memory[11][2] ),
    .A2(_1977_),
    .A1(\charlie_0.memory[13][2] ));
 sg13g2_a22oi_1 _2924_ (.Y(_2028_),
    .B1(_1987_),
    .B2(\charlie_0.memory[2][2] ),
    .A2(_1983_),
    .A1(\charlie_0.memory[6][2] ));
 sg13g2_a22oi_1 _2925_ (.Y(_2029_),
    .B1(_1981_),
    .B2(\charlie_0.memory[15][2] ),
    .A2(_1971_),
    .A1(\charlie_0.memory[14][2] ));
 sg13g2_a21oi_1 _2926_ (.A1(\charlie_0.memory[8][2] ),
    .A2(_1975_),
    .Y(_2030_),
    .B1(net1022));
 sg13g2_nand4_1 _2927_ (.B(_2028_),
    .C(_2029_),
    .A(_2025_),
    .Y(_2031_),
    .D(_2030_));
 sg13g2_a22oi_1 _2928_ (.Y(_2032_),
    .B1(_1991_),
    .B2(\charlie_0.memory[7][2] ),
    .A2(_1984_),
    .A1(\charlie_0.memory[5][2] ));
 sg13g2_a22oi_1 _2929_ (.Y(_2033_),
    .B1(_1988_),
    .B2(\charlie_0.memory[9][2] ),
    .A2(_1973_),
    .A1(\charlie_0.memory[10][2] ));
 sg13g2_nand4_1 _2930_ (.B(_2027_),
    .C(_2032_),
    .A(_2026_),
    .Y(_2034_),
    .D(_2033_));
 sg13g2_or2_1 _2931_ (.X(_2035_),
    .B(_2034_),
    .A(_2031_));
 sg13g2_a21oi_1 _2932_ (.A1(_0058_),
    .A2(net1023),
    .Y(_2036_),
    .B1(net1105));
 sg13g2_xor2_1 _2933_ (.B(net3),
    .A(\charlie_0.memory[22][3] ),
    .X(_2037_));
 sg13g2_a22oi_1 _2934_ (.Y(_2038_),
    .B1(_2037_),
    .B2(net1105),
    .A2(_2036_),
    .A1(_2035_));
 sg13g2_nor2b_1 _2935_ (.A(_2038_),
    .B_N(_2024_),
    .Y(_2039_));
 sg13g2_xnor2_1 _2936_ (.Y(uo_out[2]),
    .A(_0052_),
    .B(_2039_));
 sg13g2_a22oi_1 _2937_ (.Y(_2040_),
    .B1(_1991_),
    .B2(\charlie_0.memory[7][3] ),
    .A2(_1977_),
    .A1(\charlie_0.memory[13][3] ));
 sg13g2_a22oi_1 _2938_ (.Y(_2041_),
    .B1(_1984_),
    .B2(\charlie_0.memory[5][3] ),
    .A2(_1983_),
    .A1(\charlie_0.memory[6][3] ));
 sg13g2_a22oi_1 _2939_ (.Y(_2042_),
    .B1(_1989_),
    .B2(\charlie_0.memory[1][3] ),
    .A2(_1987_),
    .A1(\charlie_0.memory[2][3] ));
 sg13g2_a22oi_1 _2940_ (.Y(_2043_),
    .B1(_1973_),
    .B2(\charlie_0.memory[10][3] ),
    .A2(_1971_),
    .A1(\charlie_0.memory[14][3] ));
 sg13g2_a22oi_1 _2941_ (.Y(_2044_),
    .B1(_1988_),
    .B2(\charlie_0.memory[9][3] ),
    .A2(_1981_),
    .A1(\charlie_0.memory[15][3] ));
 sg13g2_a21oi_1 _2942_ (.A1(\charlie_0.memory[11][3] ),
    .A2(_1992_),
    .Y(_2045_),
    .B1(net1022));
 sg13g2_nand4_1 _2943_ (.B(_2043_),
    .C(_2044_),
    .A(_2040_),
    .Y(_2046_),
    .D(_2045_));
 sg13g2_a22oi_1 _2944_ (.Y(_2047_),
    .B1(_1985_),
    .B2(\charlie_0.memory[4][3] ),
    .A2(_1975_),
    .A1(\charlie_0.memory[8][3] ));
 sg13g2_a22oi_1 _2945_ (.Y(_2048_),
    .B1(_1990_),
    .B2(\charlie_0.memory[3][3] ),
    .A2(_1986_),
    .A1(\charlie_0.memory[12][3] ));
 sg13g2_nand4_1 _2946_ (.B(_2042_),
    .C(_2047_),
    .A(_2041_),
    .Y(_2049_),
    .D(_2048_));
 sg13g2_nor2_1 _2947_ (.A(_2046_),
    .B(_2049_),
    .Y(_2050_));
 sg13g2_a21oi_1 _2948_ (.A1(_0059_),
    .A2(net1023),
    .Y(_2051_),
    .B1(_2050_));
 sg13g2_o21ai_1 _2949_ (.B1(_2024_),
    .Y(_2052_),
    .A1(net1105),
    .A2(_2051_));
 sg13g2_a21oi_1 _2950_ (.A1(_1963_),
    .A2(net1105),
    .Y(_2053_),
    .B1(_2052_));
 sg13g2_xnor2_1 _2951_ (.Y(uo_out[3]),
    .A(_0052_),
    .B(_2053_));
 sg13g2_a22oi_1 _2952_ (.Y(_2054_),
    .B1(_1990_),
    .B2(\charlie_0.memory[3][4] ),
    .A2(_1987_),
    .A1(\charlie_0.memory[2][4] ));
 sg13g2_a22oi_1 _2953_ (.Y(_2055_),
    .B1(_1986_),
    .B2(\charlie_0.memory[12][4] ),
    .A2(_1984_),
    .A1(\charlie_0.memory[5][4] ));
 sg13g2_a22oi_1 _2954_ (.Y(_2056_),
    .B1(_1981_),
    .B2(\charlie_0.memory[15][4] ),
    .A2(_1977_),
    .A1(\charlie_0.memory[13][4] ));
 sg13g2_a22oi_1 _2955_ (.Y(_2057_),
    .B1(_1992_),
    .B2(\charlie_0.memory[11][4] ),
    .A2(_1985_),
    .A1(\charlie_0.memory[4][4] ));
 sg13g2_a22oi_1 _2956_ (.Y(_2058_),
    .B1(_1991_),
    .B2(\charlie_0.memory[7][4] ),
    .A2(_1989_),
    .A1(\charlie_0.memory[1][4] ));
 sg13g2_a21oi_1 _2957_ (.A1(\charlie_0.memory[14][4] ),
    .A2(_1971_),
    .Y(_2059_),
    .B1(net1022));
 sg13g2_nand4_1 _2958_ (.B(_2057_),
    .C(_2058_),
    .A(_2056_),
    .Y(_2060_),
    .D(_2059_));
 sg13g2_a22oi_1 _2959_ (.Y(_2061_),
    .B1(_1983_),
    .B2(\charlie_0.memory[6][4] ),
    .A2(_1975_),
    .A1(\charlie_0.memory[8][4] ));
 sg13g2_a22oi_1 _2960_ (.Y(_2062_),
    .B1(_1988_),
    .B2(\charlie_0.memory[9][4] ),
    .A2(_1973_),
    .A1(\charlie_0.memory[10][4] ));
 sg13g2_nand4_1 _2961_ (.B(_2055_),
    .C(_2061_),
    .A(_2054_),
    .Y(_2063_),
    .D(_2062_));
 sg13g2_nor2_1 _2962_ (.A(_2060_),
    .B(_2063_),
    .Y(_2064_));
 sg13g2_a21oi_1 _2963_ (.A1(_0060_),
    .A2(net1023),
    .Y(_2065_),
    .B1(_2064_));
 sg13g2_o21ai_1 _2964_ (.B1(_2024_),
    .Y(_2066_),
    .A1(net1105),
    .A2(_2065_));
 sg13g2_a21oi_1 _2965_ (.A1(_1961_),
    .A2(net1105),
    .Y(_2067_),
    .B1(_2066_));
 sg13g2_xnor2_1 _2966_ (.Y(uo_out[4]),
    .A(_0052_),
    .B(_2067_));
 sg13g2_a22oi_1 _2967_ (.Y(_2068_),
    .B1(_1991_),
    .B2(\charlie_0.memory[7][5] ),
    .A2(_1981_),
    .A1(\charlie_0.memory[15][5] ));
 sg13g2_a22oi_1 _2968_ (.Y(_2069_),
    .B1(_1992_),
    .B2(\charlie_0.memory[11][5] ),
    .A2(_1989_),
    .A1(\charlie_0.memory[1][5] ));
 sg13g2_a22oi_1 _2969_ (.Y(_2070_),
    .B1(_1986_),
    .B2(\charlie_0.memory[12][5] ),
    .A2(_1973_),
    .A1(\charlie_0.memory[10][5] ));
 sg13g2_a22oi_1 _2970_ (.Y(_2071_),
    .B1(_1987_),
    .B2(\charlie_0.memory[2][5] ),
    .A2(_1975_),
    .A1(\charlie_0.memory[8][5] ));
 sg13g2_a22oi_1 _2971_ (.Y(_2072_),
    .B1(_1988_),
    .B2(\charlie_0.memory[9][5] ),
    .A2(_1977_),
    .A1(\charlie_0.memory[13][5] ));
 sg13g2_a21oi_1 _2972_ (.A1(\charlie_0.memory[6][5] ),
    .A2(_1983_),
    .Y(_2073_),
    .B1(net1022));
 sg13g2_nand4_1 _2973_ (.B(_2071_),
    .C(_2072_),
    .A(_2070_),
    .Y(_2074_),
    .D(_2073_));
 sg13g2_a22oi_1 _2974_ (.Y(_2075_),
    .B1(_1990_),
    .B2(\charlie_0.memory[3][5] ),
    .A2(_1985_),
    .A1(\charlie_0.memory[4][5] ));
 sg13g2_a22oi_1 _2975_ (.Y(_2076_),
    .B1(_1984_),
    .B2(\charlie_0.memory[5][5] ),
    .A2(_1971_),
    .A1(\charlie_0.memory[14][5] ));
 sg13g2_nand4_1 _2976_ (.B(_2069_),
    .C(_2075_),
    .A(_2068_),
    .Y(_2077_),
    .D(_2076_));
 sg13g2_or2_1 _2977_ (.X(_2078_),
    .B(_2077_),
    .A(_2074_));
 sg13g2_a21oi_1 _2978_ (.A1(_0061_),
    .A2(net1023),
    .Y(_2079_),
    .B1(_2004_));
 sg13g2_mux4_1 _2979_ (.S0(net1172),
    .A0(\counter[8] ),
    .A1(\counter[9] ),
    .A2(\counter[10] ),
    .A3(\counter[11] ),
    .S1(net1170),
    .X(_2080_));
 sg13g2_inv_1 _2980_ (.Y(_2081_),
    .A(_2080_));
 sg13g2_mux2_1 _2981_ (.A0(\counter[12] ),
    .A1(\counter[13] ),
    .S(net1172),
    .X(_2082_));
 sg13g2_nand2_1 _2982_ (.Y(_2083_),
    .A(_1790_),
    .B(_2082_));
 sg13g2_mux2_1 _2983_ (.A0(\counter[14] ),
    .A1(\counter[15] ),
    .S(net1173),
    .X(_2084_));
 sg13g2_a21oi_1 _2984_ (.A1(net1170),
    .A2(_2084_),
    .Y(_2085_),
    .B1(_1789_));
 sg13g2_a221oi_1 _2985_ (.B2(_2085_),
    .C1(\charlie_0.memory[16][4] ),
    .B1(_2083_),
    .A1(_1789_),
    .Y(_2086_),
    .A2(_2081_));
 sg13g2_mux2_1 _2986_ (.A0(\counter[20] ),
    .A1(\counter[21] ),
    .S(net1173),
    .X(_2087_));
 sg13g2_nor2_1 _2987_ (.A(net1173),
    .B(\counter[22] ),
    .Y(_2088_));
 sg13g2_o21ai_1 _2988_ (.B1(net1171),
    .Y(_2089_),
    .A1(_1791_),
    .A2(\counter[23] ));
 sg13g2_a21oi_1 _2989_ (.A1(_1790_),
    .A2(_2087_),
    .Y(_2090_),
    .B1(_1789_));
 sg13g2_o21ai_1 _2990_ (.B1(_2090_),
    .Y(_2091_),
    .A1(_2088_),
    .A2(_2089_));
 sg13g2_mux2_1 _2991_ (.A0(\counter[16] ),
    .A1(\counter[17] ),
    .S(net1174),
    .X(_2092_));
 sg13g2_nand2b_1 _2992_ (.Y(_2093_),
    .B(net1173),
    .A_N(\counter[19] ));
 sg13g2_o21ai_1 _2993_ (.B1(_2093_),
    .Y(_2094_),
    .A1(net1173),
    .A2(\counter[18] ));
 sg13g2_a21oi_1 _2994_ (.A1(_1790_),
    .A2(_2092_),
    .Y(_2095_),
    .B1(\charlie_0.memory[16][2] ));
 sg13g2_o21ai_1 _2995_ (.B1(_2095_),
    .Y(_2096_),
    .A1(_1790_),
    .A2(_2094_));
 sg13g2_nand4_1 _2996_ (.B(\charlie_0.memory[16][3] ),
    .C(_2091_),
    .A(_1787_),
    .Y(_2097_),
    .D(_2096_));
 sg13g2_mux4_1 _2997_ (.S0(net1172),
    .A0(\counter[24] ),
    .A1(\counter[25] ),
    .A2(\counter[26] ),
    .A3(\counter[27] ),
    .S1(net1170),
    .X(_2098_));
 sg13g2_nor2_1 _2998_ (.A(\charlie_0.memory[16][2] ),
    .B(_2098_),
    .Y(_2099_));
 sg13g2_nor2b_1 _2999_ (.A(\counter[29] ),
    .B_N(net1172),
    .Y(_2100_));
 sg13g2_nor2_1 _3000_ (.A(net1172),
    .B(\counter[28] ),
    .Y(_2101_));
 sg13g2_nor3_1 _3001_ (.A(net1170),
    .B(_2100_),
    .C(_2101_),
    .Y(_2102_));
 sg13g2_nor2b_1 _3002_ (.A(\counter[31] ),
    .B_N(net1172),
    .Y(_2103_));
 sg13g2_o21ai_1 _3003_ (.B1(net1170),
    .Y(_2104_),
    .A1(net1173),
    .A2(\counter[30] ));
 sg13g2_o21ai_1 _3004_ (.B1(\charlie_0.memory[16][2] ),
    .Y(_2105_),
    .A1(_2103_),
    .A2(_2104_));
 sg13g2_o21ai_1 _3005_ (.B1(\charlie_0.memory[16][4] ),
    .Y(_2106_),
    .A1(_2102_),
    .A2(_2105_));
 sg13g2_nor2_1 _3006_ (.A(_2099_),
    .B(_2106_),
    .Y(_2107_));
 sg13g2_or2_1 _3007_ (.X(_2108_),
    .B(_2106_),
    .A(_2099_));
 sg13g2_a22oi_1 _3008_ (.Y(_2109_),
    .B1(_2107_),
    .B2(_0067_),
    .A2(_2086_),
    .A1(_1788_));
 sg13g2_nand3_1 _3009_ (.B(_2097_),
    .C(_2109_),
    .A(\charlie_0.memory[22][1] ),
    .Y(_2110_));
 sg13g2_a21oi_1 _3010_ (.A1(_1774_),
    .A2(_1968_),
    .Y(_2111_),
    .B1(net1146));
 sg13g2_a22oi_1 _3011_ (.Y(_2112_),
    .B1(_2110_),
    .B2(_2111_),
    .A2(_2079_),
    .A1(_2078_));
 sg13g2_xor2_1 _3012_ (.B(_2112_),
    .A(_0052_),
    .X(uo_out[5]));
 sg13g2_mux2_1 _3013_ (.A0(net1204),
    .A1(net1201),
    .S(net1174),
    .X(_2113_));
 sg13g2_nand2_1 _3014_ (.Y(_2114_),
    .A(_1790_),
    .B(_2113_));
 sg13g2_mux2_1 _3015_ (.A0(\counter[6] ),
    .A1(\counter[7] ),
    .S(net1172),
    .X(_2115_));
 sg13g2_a21oi_1 _3016_ (.A1(net1170),
    .A2(_2115_),
    .Y(_2116_),
    .B1(_1789_));
 sg13g2_mux4_1 _3017_ (.S0(net1174),
    .A0(_1826_),
    .A1(_1827_),
    .A2(_0069_),
    .A3(_0068_),
    .S1(net1171),
    .X(_2117_));
 sg13g2_a22oi_1 _3018_ (.Y(_2118_),
    .B1(_2117_),
    .B2(_1789_),
    .A2(_2116_),
    .A1(_2114_));
 sg13g2_nand3_1 _3019_ (.B(_2091_),
    .C(_2096_),
    .A(\charlie_0.memory[16][4] ),
    .Y(_2119_));
 sg13g2_a21oi_1 _3020_ (.A1(_1787_),
    .A2(_2118_),
    .Y(_2120_),
    .B1(\charlie_0.memory[16][3] ));
 sg13g2_nor2b_1 _3021_ (.A(_2086_),
    .B_N(\charlie_0.memory[16][3] ),
    .Y(_2121_));
 sg13g2_a22oi_1 _3022_ (.Y(_2122_),
    .B1(_2121_),
    .B2(_2108_),
    .A2(_2120_),
    .A1(_2119_));
 sg13g2_nor2_1 _3023_ (.A(\charlie_0.memory[16][5] ),
    .B(_2122_),
    .Y(_2123_));
 sg13g2_o21ai_1 _3024_ (.B1(_2009_),
    .Y(_2124_),
    .A1(_1786_),
    .A2(clknet_1_0__leaf_clk));
 sg13g2_a22oi_1 _3025_ (.Y(_2125_),
    .B1(_1985_),
    .B2(\charlie_0.memory[4][6] ),
    .A2(_1984_),
    .A1(\charlie_0.memory[5][6] ));
 sg13g2_a22oi_1 _3026_ (.Y(_2126_),
    .B1(_1986_),
    .B2(\charlie_0.memory[12][6] ),
    .A2(_1975_),
    .A1(\charlie_0.memory[8][6] ));
 sg13g2_a22oi_1 _3027_ (.Y(_2127_),
    .B1(_1987_),
    .B2(\charlie_0.memory[2][6] ),
    .A2(_1977_),
    .A1(\charlie_0.memory[13][6] ));
 sg13g2_a22oi_1 _3028_ (.Y(_2128_),
    .B1(_1983_),
    .B2(\charlie_0.memory[6][6] ),
    .A2(_1981_),
    .A1(\charlie_0.memory[15][6] ));
 sg13g2_a21oi_1 _3029_ (.A1(\charlie_0.memory[3][6] ),
    .A2(_1990_),
    .Y(_2129_),
    .B1(net1023));
 sg13g2_nand4_1 _3030_ (.B(_2127_),
    .C(_2128_),
    .A(_2126_),
    .Y(_2130_),
    .D(_2129_));
 sg13g2_a22oi_1 _3031_ (.Y(_2131_),
    .B1(_1991_),
    .B2(\charlie_0.memory[7][6] ),
    .A2(_1973_),
    .A1(\charlie_0.memory[10][6] ));
 sg13g2_a22oi_1 _3032_ (.Y(_2132_),
    .B1(_1989_),
    .B2(\charlie_0.memory[1][6] ),
    .A2(_1971_),
    .A1(\charlie_0.memory[14][6] ));
 sg13g2_a22oi_1 _3033_ (.Y(_0298_),
    .B1(_1992_),
    .B2(\charlie_0.memory[11][6] ),
    .A2(_1988_),
    .A1(\charlie_0.memory[9][6] ));
 sg13g2_nand4_1 _3034_ (.B(_2131_),
    .C(_2132_),
    .A(_2125_),
    .Y(_0299_),
    .D(_0298_));
 sg13g2_a21oi_1 _3035_ (.A1(_0062_),
    .A2(net1023),
    .Y(_0300_),
    .B1(_2004_));
 sg13g2_o21ai_1 _3036_ (.B1(_0300_),
    .Y(_0301_),
    .A1(_2130_),
    .A2(_0299_));
 sg13g2_o21ai_1 _3037_ (.B1(_0301_),
    .Y(_0302_),
    .A1(_2123_),
    .A2(_2124_));
 sg13g2_a21oi_1 _3038_ (.A1(_1967_),
    .A2(net1105),
    .Y(_0303_),
    .B1(_0302_));
 sg13g2_xor2_1 _3039_ (.B(_0303_),
    .A(_0052_),
    .X(uo_out[6]));
 sg13g2_xor2_1 _3040_ (.B(\bi_out[0] ),
    .A(net1148),
    .X(uio_out[0]));
 sg13g2_xor2_1 _3041_ (.B(\bi_out[1] ),
    .A(net1147),
    .X(uio_out[1]));
 sg13g2_xor2_1 _3042_ (.B(\bi_out[2] ),
    .A(net1147),
    .X(uio_out[2]));
 sg13g2_xor2_1 _3043_ (.B(\bi_out[3] ),
    .A(net1147),
    .X(uio_out[3]));
 sg13g2_xor2_1 _3044_ (.B(\bi_out[4] ),
    .A(net1147),
    .X(uio_out[4]));
 sg13g2_xor2_1 _3045_ (.B(\bi_out[5] ),
    .A(net1147),
    .X(uio_out[5]));
 sg13g2_xor2_1 _3046_ (.B(\bi_out[6] ),
    .A(net1147),
    .X(uio_out[6]));
 sg13g2_xor2_1 _3047_ (.B(\bi_out[7] ),
    .A(net1147),
    .X(uio_out[7]));
 sg13g2_xor2_1 _3048_ (.B(\bi_en[0] ),
    .A(net1149),
    .X(uio_oe[0]));
 sg13g2_xor2_1 _3049_ (.B(\bi_en[1] ),
    .A(net1149),
    .X(uio_oe[1]));
 sg13g2_xor2_1 _3050_ (.B(\bi_en[2] ),
    .A(net1149),
    .X(uio_oe[2]));
 sg13g2_xor2_1 _3051_ (.B(\bi_en[3] ),
    .A(net1149),
    .X(uio_oe[3]));
 sg13g2_xor2_1 _3052_ (.B(\bi_en[4] ),
    .A(net1149),
    .X(uio_oe[4]));
 sg13g2_xor2_1 _3053_ (.B(\bi_en[5] ),
    .A(net1149),
    .X(uio_oe[5]));
 sg13g2_xor2_1 _3054_ (.B(\bi_en[6] ),
    .A(net1149),
    .X(uio_oe[6]));
 sg13g2_xor2_1 _3055_ (.B(\bi_en[7] ),
    .A(net1149),
    .X(uio_oe[7]));
 sg13g2_nand2_1 _3056_ (.Y(_0304_),
    .A(net1200),
    .B(_1858_));
 sg13g2_nor3_2 _3057_ (.A(net1211),
    .B(net1209),
    .C(net1207),
    .Y(_0305_));
 sg13g2_a21oi_1 _3058_ (.A1(net295),
    .A2(_0305_),
    .Y(_0008_),
    .B1(_0304_));
 sg13g2_nand3_1 _3059_ (.B(_1827_),
    .C(_1828_),
    .A(net1212),
    .Y(_0306_));
 sg13g2_nor3_1 _3060_ (.A(_0068_),
    .B(_1858_),
    .C(_1860_),
    .Y(_0307_));
 sg13g2_or3_1 _3061_ (.A(net304),
    .B(_1858_),
    .C(_1860_),
    .X(_0308_));
 sg13g2_nand3_1 _3062_ (.B(_0306_),
    .C(_0307_),
    .A(net280),
    .Y(_0309_));
 sg13g2_inv_1 _3063_ (.Y(_0009_),
    .A(net281));
 sg13g2_nor2_1 _3064_ (.A(net1211),
    .B(_1827_),
    .Y(_0310_));
 sg13g2_nor2b_2 _3065_ (.A(net1205),
    .B_N(net1203),
    .Y(_0311_));
 sg13g2_nand2b_2 _3066_ (.Y(_0312_),
    .B(net1203),
    .A_N(net1205));
 sg13g2_nand2_1 _3067_ (.Y(_0313_),
    .A(net1200),
    .B(_0311_));
 sg13g2_a21oi_1 _3068_ (.A1(_1828_),
    .A2(_0310_),
    .Y(_0010_),
    .B1(_0313_));
 sg13g2_xor2_1 _3069_ (.B(_1858_),
    .A(net1200),
    .X(_0314_));
 sg13g2_o21ai_1 _3070_ (.B1(_0314_),
    .Y(_0315_),
    .A1(net1207),
    .A2(_1847_));
 sg13g2_nand2b_1 _3071_ (.Y(_0316_),
    .B(_1858_),
    .A_N(net1200));
 sg13g2_a21o_1 _3072_ (.A2(_0316_),
    .A1(_1861_),
    .B1(net304),
    .X(_0317_));
 sg13g2_nor2_1 _3073_ (.A(_0315_),
    .B(_0317_),
    .Y(_0011_));
 sg13g2_nand2_1 _3074_ (.Y(_0318_),
    .A(net1207),
    .B(_1846_));
 sg13g2_nor2b_1 _3075_ (.A(_0316_),
    .B_N(_0318_),
    .Y(_0012_));
 sg13g2_nor3_1 _3076_ (.A(_1826_),
    .B(net1209),
    .C(_1828_),
    .Y(_0319_));
 sg13g2_nor3_1 _3077_ (.A(net1200),
    .B(_0308_),
    .C(_0319_),
    .Y(_0013_));
 sg13g2_nor3_1 _3078_ (.A(net1211),
    .B(_1827_),
    .C(_1828_),
    .Y(_0320_));
 sg13g2_nor3_1 _3079_ (.A(net1200),
    .B(_0312_),
    .C(_0320_),
    .Y(_0014_));
 sg13g2_or2_1 _3080_ (.X(_0321_),
    .B(_0314_),
    .A(_1852_));
 sg13g2_nor2_1 _3081_ (.A(_0317_),
    .B(_0321_),
    .Y(_0015_));
 sg13g2_nand2_1 _3082_ (.Y(_0322_),
    .A(net1153),
    .B(net1155));
 sg13g2_nand2b_2 _3083_ (.Y(_0323_),
    .B(net1155),
    .A_N(net1202));
 sg13g2_nand2b_2 _3084_ (.Y(_0324_),
    .B(net1206),
    .A_N(net1204));
 sg13g2_nor3_2 _3085_ (.A(net1152),
    .B(_0323_),
    .C(_0324_),
    .Y(_0325_));
 sg13g2_or3_2 _3086_ (.A(net1154),
    .B(net1206),
    .C(net1204),
    .X(_0326_));
 sg13g2_nor2_2 _3087_ (.A(_0323_),
    .B(_0326_),
    .Y(_0327_));
 sg13g2_nand2b_2 _3088_ (.Y(_0328_),
    .B(net1202),
    .A_N(net1155));
 sg13g2_nor3_2 _3089_ (.A(net1152),
    .B(_0324_),
    .C(_0328_),
    .Y(_0329_));
 sg13g2_nor3_2 _3090_ (.A(net1152),
    .B(_0312_),
    .C(_0323_),
    .Y(_0330_));
 sg13g2_or2_2 _3091_ (.X(_0331_),
    .B(net1202),
    .A(net1155));
 sg13g2_nor2_1 _3092_ (.A(_0326_),
    .B(_0331_),
    .Y(_0332_));
 sg13g2_a21oi_2 _3093_ (.B1(_0332_),
    .Y(_0333_),
    .A2(net1155),
    .A1(net1153));
 sg13g2_o21ai_1 _3094_ (.B1(_0322_),
    .Y(_0334_),
    .A1(_0326_),
    .A2(_0331_));
 sg13g2_nor3_1 _3095_ (.A(_0064_),
    .B(_1861_),
    .C(_0328_),
    .Y(_0335_));
 sg13g2_nor2_2 _3096_ (.A(net1026),
    .B(_0335_),
    .Y(_0336_));
 sg13g2_nor3_2 _3097_ (.A(net1155),
    .B(net1202),
    .C(_0064_),
    .Y(_0337_));
 sg13g2_nor2_1 _3098_ (.A(_1861_),
    .B(_0331_),
    .Y(_0338_));
 sg13g2_and2_2 _3099_ (.A(_1860_),
    .B(_0337_),
    .X(_0339_));
 sg13g2_nand3b_1 _3100_ (.B(net1206),
    .C(net1204),
    .Y(_0340_),
    .A_N(net1154));
 sg13g2_nand2_2 _3101_ (.Y(_0341_),
    .A(net1155),
    .B(net1201));
 sg13g2_nor2_2 _3102_ (.A(_0340_),
    .B(_0341_),
    .Y(_0342_));
 sg13g2_nor2_2 _3103_ (.A(_0326_),
    .B(_0341_),
    .Y(_0343_));
 sg13g2_nor3_2 _3104_ (.A(net1152),
    .B(_0312_),
    .C(_0341_),
    .Y(_0344_));
 sg13g2_nor3_2 _3105_ (.A(net1153),
    .B(_0324_),
    .C(_0331_),
    .Y(_0345_));
 sg13g2_nor2_2 _3106_ (.A(_0328_),
    .B(_0340_),
    .Y(_0346_));
 sg13g2_nor4_2 _3107_ (.A(net1206),
    .B(net1204),
    .C(_0064_),
    .Y(_0347_),
    .D(_0328_));
 sg13g2_nor3_2 _3108_ (.A(_0064_),
    .B(_0312_),
    .C(_0328_),
    .Y(_0348_));
 sg13g2_nor2b_2 _3109_ (.A(_0324_),
    .B_N(_0337_),
    .Y(_0349_));
 sg13g2_nor3_2 _3110_ (.A(_0064_),
    .B(_0324_),
    .C(_0328_),
    .Y(_0350_));
 sg13g2_nor2_2 _3111_ (.A(_0323_),
    .B(_0340_),
    .Y(_0351_));
 sg13g2_nor3_2 _3112_ (.A(net1152),
    .B(_0312_),
    .C(_0328_),
    .Y(_0352_));
 sg13g2_and2_2 _3113_ (.A(_0311_),
    .B(_0337_),
    .X(_0353_));
 sg13g2_nor3_2 _3114_ (.A(net1152),
    .B(_0312_),
    .C(_0331_),
    .Y(_0354_));
 sg13g2_and2_2 _3115_ (.A(_1858_),
    .B(_0337_),
    .X(_0355_));
 sg13g2_nor3_2 _3116_ (.A(net1152),
    .B(_0324_),
    .C(_0341_),
    .Y(_0356_));
 sg13g2_nor2_2 _3117_ (.A(_0326_),
    .B(_0328_),
    .Y(_0357_));
 sg13g2_nor2_2 _3118_ (.A(_0331_),
    .B(_0340_),
    .Y(_0358_));
 sg13g2_a22oi_1 _3119_ (.Y(_0359_),
    .B1(_0357_),
    .B2(\charlie_0.memory[4][2] ),
    .A2(_0345_),
    .A1(\charlie_0.memory[1][2] ));
 sg13g2_a22oi_1 _3120_ (.Y(_0360_),
    .B1(_0358_),
    .B2(\charlie_0.memory[3][2] ),
    .A2(_0347_),
    .A1(\charlie_0.memory[20][2] ));
 sg13g2_a22oi_1 _3121_ (.Y(_0361_),
    .B1(_0349_),
    .B2(net1158),
    .A2(_0330_),
    .A1(\charlie_0.memory[10][2] ));
 sg13g2_a22oi_1 _3122_ (.Y(_0362_),
    .B1(_0356_),
    .B2(\charlie_0.memory[13][2] ),
    .A2(_0351_),
    .A1(\charlie_0.memory[11][2] ));
 sg13g2_a22oi_1 _3123_ (.Y(_0363_),
    .B1(_0354_),
    .B2(\charlie_0.memory[2][2] ),
    .A2(_0325_),
    .A1(\charlie_0.memory[9][2] ));
 sg13g2_a22oi_1 _3124_ (.Y(_0364_),
    .B1(_0339_),
    .B2(net1151),
    .A2(_0329_),
    .A1(\charlie_0.memory[5][2] ));
 sg13g2_nand4_1 _3125_ (.B(_0359_),
    .C(_0360_),
    .A(_0336_),
    .Y(_0365_),
    .D(_0364_));
 sg13g2_a22oi_1 _3126_ (.Y(_0366_),
    .B1(_0350_),
    .B2(\charlie_0.memory[21][2] ),
    .A2(_0343_),
    .A1(\charlie_0.memory[12][2] ));
 sg13g2_a22oi_1 _3127_ (.Y(_0367_),
    .B1(_0355_),
    .B2(\charlie_0.memory[16][2] ),
    .A2(_0344_),
    .A1(\charlie_0.memory[14][2] ));
 sg13g2_a22oi_1 _3128_ (.Y(_0368_),
    .B1(_0353_),
    .B2(\charlie_0.memory[18][2] ),
    .A2(_0348_),
    .A1(\charlie_0.memory[22][2] ));
 sg13g2_nand4_1 _3129_ (.B(_0366_),
    .C(_0367_),
    .A(_0361_),
    .Y(_0369_),
    .D(_0368_));
 sg13g2_a22oi_1 _3130_ (.Y(_0370_),
    .B1(_0346_),
    .B2(\charlie_0.memory[7][2] ),
    .A2(_0342_),
    .A1(\charlie_0.memory[15][2] ));
 sg13g2_a22oi_1 _3131_ (.Y(_0371_),
    .B1(_0352_),
    .B2(\charlie_0.memory[6][2] ),
    .A2(_0327_),
    .A1(\charlie_0.memory[8][2] ));
 sg13g2_nand4_1 _3132_ (.B(_0363_),
    .C(_0370_),
    .A(_0362_),
    .Y(_0372_),
    .D(_0371_));
 sg13g2_or3_1 _3133_ (.A(_0365_),
    .B(_0369_),
    .C(_0372_),
    .X(_0373_));
 sg13g2_xor2_1 _3134_ (.B(net1210),
    .A(net1151),
    .X(_0374_));
 sg13g2_xnor2_1 _3135_ (.Y(_0375_),
    .A(net1151),
    .B(net1210));
 sg13g2_a21oi_1 _3136_ (.A1(_0058_),
    .A2(_0334_),
    .Y(_0376_),
    .B1(_0375_));
 sg13g2_xor2_1 _3137_ (.B(\charlie_0.charlie_index[0] ),
    .A(net1151),
    .X(_0377_));
 sg13g2_xnor2_1 _3138_ (.Y(_0378_),
    .A(net1151),
    .B(\charlie_0.charlie_index[0] ));
 sg13g2_a22oi_1 _3139_ (.Y(_0379_),
    .B1(_0345_),
    .B2(\charlie_0.memory[1][0] ),
    .A2(_0329_),
    .A1(\charlie_0.memory[5][0] ));
 sg13g2_nand2_1 _3140_ (.Y(_0380_),
    .A(net1174),
    .B(_0355_));
 sg13g2_a22oi_1 _3141_ (.Y(_0381_),
    .B1(_0344_),
    .B2(\charlie_0.memory[14][0] ),
    .A2(_0342_),
    .A1(\charlie_0.memory[15][0] ));
 sg13g2_a22oi_1 _3142_ (.Y(_0382_),
    .B1(_0343_),
    .B2(\charlie_0.memory[12][0] ),
    .A2(_0327_),
    .A1(\charlie_0.memory[8][0] ));
 sg13g2_a22oi_1 _3143_ (.Y(_0383_),
    .B1(_0353_),
    .B2(\charlie_0.memory[18][0] ),
    .A2(_0351_),
    .A1(\charlie_0.memory[11][0] ));
 sg13g2_a22oi_1 _3144_ (.Y(_0384_),
    .B1(_0358_),
    .B2(\charlie_0.memory[3][0] ),
    .A2(_0357_),
    .A1(\charlie_0.memory[4][0] ));
 sg13g2_a22oi_1 _3145_ (.Y(_0385_),
    .B1(_0354_),
    .B2(\charlie_0.memory[2][0] ),
    .A2(_0325_),
    .A1(\charlie_0.memory[9][0] ));
 sg13g2_a22oi_1 _3146_ (.Y(_0386_),
    .B1(_0349_),
    .B2(net1164),
    .A2(_0348_),
    .A1(net1146));
 sg13g2_nand4_1 _3147_ (.B(_0383_),
    .C(_0384_),
    .A(_0336_),
    .Y(_0387_),
    .D(_0386_));
 sg13g2_a22oi_1 _3148_ (.Y(_0388_),
    .B1(_0350_),
    .B2(\charlie_0.memory[21][0] ),
    .A2(_0346_),
    .A1(\charlie_0.memory[7][0] ));
 sg13g2_a22oi_1 _3149_ (.Y(_0389_),
    .B1(_0356_),
    .B2(\charlie_0.memory[13][0] ),
    .A2(_0352_),
    .A1(\charlie_0.memory[6][0] ));
 sg13g2_nand4_1 _3150_ (.B(_0385_),
    .C(_0388_),
    .A(_0379_),
    .Y(_0390_),
    .D(_0389_));
 sg13g2_a22oi_1 _3151_ (.Y(_0391_),
    .B1(_0347_),
    .B2(\charlie_0.memory[20][0] ),
    .A2(_0330_),
    .A1(\charlie_0.memory[10][0] ));
 sg13g2_nand4_1 _3152_ (.B(_0381_),
    .C(_0382_),
    .A(_0380_),
    .Y(_0392_),
    .D(_0391_));
 sg13g2_or3_1 _3153_ (.A(_0387_),
    .B(_0390_),
    .C(_0392_),
    .X(_0393_));
 sg13g2_a21oi_1 _3154_ (.A1(_0055_),
    .A2(net1026),
    .Y(_0394_),
    .B1(_0374_));
 sg13g2_a221oi_1 _3155_ (.B2(_0394_),
    .C1(_0377_),
    .B1(_0393_),
    .A1(_0373_),
    .Y(_0395_),
    .A2(_0376_));
 sg13g2_xor2_1 _3156_ (.B(\charlie_0.charlie_index[2] ),
    .A(\charlie_0.is_mirror ),
    .X(_0396_));
 sg13g2_xnor2_1 _3157_ (.Y(_0397_),
    .A(net1151),
    .B(\charlie_0.charlie_index[2] ));
 sg13g2_a22oi_1 _3158_ (.Y(_0398_),
    .B1(_0351_),
    .B2(\charlie_0.memory[11][1] ),
    .A2(_0327_),
    .A1(\charlie_0.memory[8][1] ));
 sg13g2_a22oi_1 _3159_ (.Y(_0399_),
    .B1(_0354_),
    .B2(\charlie_0.memory[2][1] ),
    .A2(_0338_),
    .A1(net1152));
 sg13g2_a22oi_1 _3160_ (.Y(_0400_),
    .B1(_0355_),
    .B2(net1171),
    .A2(_0353_),
    .A1(\charlie_0.memory[18][1] ));
 sg13g2_a22oi_1 _3161_ (.Y(_0401_),
    .B1(_0348_),
    .B2(_1837_),
    .A2(_0346_),
    .A1(\charlie_0.memory[7][1] ));
 sg13g2_nand4_1 _3162_ (.B(_0399_),
    .C(_0400_),
    .A(_0333_),
    .Y(_0402_),
    .D(_0401_));
 sg13g2_a22oi_1 _3163_ (.Y(_0403_),
    .B1(_0358_),
    .B2(\charlie_0.memory[3][1] ),
    .A2(_0344_),
    .A1(\charlie_0.memory[14][1] ));
 sg13g2_a22oi_1 _3164_ (.Y(_0404_),
    .B1(_0357_),
    .B2(\charlie_0.memory[4][1] ),
    .A2(_0356_),
    .A1(\charlie_0.memory[13][1] ));
 sg13g2_a22oi_1 _3165_ (.Y(_0405_),
    .B1(_0347_),
    .B2(\charlie_0.memory[20][1] ),
    .A2(_0343_),
    .A1(\charlie_0.memory[12][1] ));
 sg13g2_a22oi_1 _3166_ (.Y(_0406_),
    .B1(_0352_),
    .B2(\charlie_0.memory[6][1] ),
    .A2(_0329_),
    .A1(\charlie_0.memory[5][1] ));
 sg13g2_nand4_1 _3167_ (.B(_0404_),
    .C(_0405_),
    .A(_0403_),
    .Y(_0407_),
    .D(_0406_));
 sg13g2_a22oi_1 _3168_ (.Y(_0408_),
    .B1(_0349_),
    .B2(net1162),
    .A2(_0345_),
    .A1(\charlie_0.memory[1][1] ));
 sg13g2_a22oi_1 _3169_ (.Y(_0409_),
    .B1(_0342_),
    .B2(\charlie_0.memory[15][1] ),
    .A2(_0325_),
    .A1(\charlie_0.memory[9][1] ));
 sg13g2_a22oi_1 _3170_ (.Y(_0410_),
    .B1(_0350_),
    .B2(\charlie_0.memory[21][1] ),
    .A2(_0330_),
    .A1(\charlie_0.memory[10][1] ));
 sg13g2_nand4_1 _3171_ (.B(_0408_),
    .C(_0409_),
    .A(_0398_),
    .Y(_0411_),
    .D(_0410_));
 sg13g2_or3_1 _3172_ (.A(_0402_),
    .B(_0407_),
    .C(_0411_),
    .X(_0412_));
 sg13g2_a21oi_1 _3173_ (.A1(_0057_),
    .A2(net1026),
    .Y(_0413_),
    .B1(_0374_));
 sg13g2_a22oi_1 _3174_ (.Y(_0414_),
    .B1(_0330_),
    .B2(\charlie_0.memory[10][3] ),
    .A2(_0325_),
    .A1(\charlie_0.memory[9][3] ));
 sg13g2_a22oi_1 _3175_ (.Y(_0415_),
    .B1(_0355_),
    .B2(\charlie_0.memory[16][3] ),
    .A2(_0345_),
    .A1(\charlie_0.memory[1][3] ));
 sg13g2_a22oi_1 _3176_ (.Y(_0416_),
    .B1(_0351_),
    .B2(\charlie_0.memory[11][3] ),
    .A2(_0342_),
    .A1(\charlie_0.memory[15][3] ));
 sg13g2_a22oi_1 _3177_ (.Y(_0417_),
    .B1(_0346_),
    .B2(\charlie_0.memory[7][3] ),
    .A2(_0327_),
    .A1(\charlie_0.memory[8][3] ));
 sg13g2_nand4_1 _3178_ (.B(_0415_),
    .C(_0416_),
    .A(_0333_),
    .Y(_0418_),
    .D(_0417_));
 sg13g2_a22oi_1 _3179_ (.Y(_0419_),
    .B1(_0350_),
    .B2(\charlie_0.memory[21][3] ),
    .A2(_0349_),
    .A1(net1156));
 sg13g2_a22oi_1 _3180_ (.Y(_0420_),
    .B1(_0354_),
    .B2(\charlie_0.memory[2][3] ),
    .A2(_0343_),
    .A1(\charlie_0.memory[12][3] ));
 sg13g2_a22oi_1 _3181_ (.Y(_0421_),
    .B1(_0358_),
    .B2(\charlie_0.memory[3][3] ),
    .A2(_0348_),
    .A1(\charlie_0.memory[22][3] ));
 sg13g2_nand4_1 _3182_ (.B(_0419_),
    .C(_0420_),
    .A(_0414_),
    .Y(_0422_),
    .D(_0421_));
 sg13g2_a22oi_1 _3183_ (.Y(_0423_),
    .B1(_0357_),
    .B2(\charlie_0.memory[4][3] ),
    .A2(_0356_),
    .A1(\charlie_0.memory[13][3] ));
 sg13g2_a22oi_1 _3184_ (.Y(_0424_),
    .B1(_0344_),
    .B2(\charlie_0.memory[14][3] ),
    .A2(_0329_),
    .A1(\charlie_0.memory[5][3] ));
 sg13g2_a22oi_1 _3185_ (.Y(_0425_),
    .B1(_0347_),
    .B2(\charlie_0.memory[20][3] ),
    .A2(_0339_),
    .A1(net1150));
 sg13g2_a22oi_1 _3186_ (.Y(_0426_),
    .B1(_0353_),
    .B2(\charlie_0.memory[18][3] ),
    .A2(_0352_),
    .A1(\charlie_0.memory[6][3] ));
 sg13g2_nand4_1 _3187_ (.B(_0424_),
    .C(_0425_),
    .A(_0423_),
    .Y(_0427_),
    .D(_0426_));
 sg13g2_or3_1 _3188_ (.A(_0418_),
    .B(_0422_),
    .C(_0427_),
    .X(_0428_));
 sg13g2_a21oi_1 _3189_ (.A1(_0059_),
    .A2(net1026),
    .Y(_0429_),
    .B1(_0375_));
 sg13g2_a221oi_1 _3190_ (.B2(_0429_),
    .C1(_0378_),
    .B1(_0428_),
    .A1(_0412_),
    .Y(_0430_),
    .A2(_0413_));
 sg13g2_nor3_1 _3191_ (.A(_0395_),
    .B(_0396_),
    .C(_0430_),
    .Y(_0431_));
 sg13g2_a22oi_1 _3192_ (.Y(_0432_),
    .B1(_0356_),
    .B2(\charlie_0.memory[13][7] ),
    .A2(_0344_),
    .A1(\charlie_0.memory[14][7] ));
 sg13g2_a22oi_1 _3193_ (.Y(_0433_),
    .B1(_0351_),
    .B2(\charlie_0.memory[11][7] ),
    .A2(_0348_),
    .A1(\charlie_0.memory[22][7] ));
 sg13g2_a22oi_1 _3194_ (.Y(_0434_),
    .B1(_0330_),
    .B2(\charlie_0.memory[10][7] ),
    .A2(_0325_),
    .A1(\charlie_0.memory[9][7] ));
 sg13g2_a22oi_1 _3195_ (.Y(_0435_),
    .B1(_0358_),
    .B2(\charlie_0.memory[3][7] ),
    .A2(_0349_),
    .A1(\charlie_0.memory[17][7] ));
 sg13g2_nand4_1 _3196_ (.B(_0433_),
    .C(_0434_),
    .A(_0432_),
    .Y(_0436_),
    .D(_0435_));
 sg13g2_a22oi_1 _3197_ (.Y(_0437_),
    .B1(_0346_),
    .B2(\charlie_0.memory[7][7] ),
    .A2(_0342_),
    .A1(\charlie_0.memory[15][7] ));
 sg13g2_a22oi_1 _3198_ (.Y(_0438_),
    .B1(_0357_),
    .B2(\charlie_0.memory[4][7] ),
    .A2(_0339_),
    .A1(\charlie_0.memory[19][7] ));
 sg13g2_a22oi_1 _3199_ (.Y(_0439_),
    .B1(_0355_),
    .B2(\charlie_0.memory[16][7] ),
    .A2(_0353_),
    .A1(\charlie_0.memory[18][7] ));
 sg13g2_a22oi_1 _3200_ (.Y(_0440_),
    .B1(_0354_),
    .B2(\charlie_0.memory[2][7] ),
    .A2(_0352_),
    .A1(\charlie_0.memory[6][7] ));
 sg13g2_a22oi_1 _3201_ (.Y(_0441_),
    .B1(_0347_),
    .B2(\charlie_0.memory[20][7] ),
    .A2(_0327_),
    .A1(\charlie_0.memory[8][7] ));
 sg13g2_a22oi_1 _3202_ (.Y(_0442_),
    .B1(_0350_),
    .B2(\charlie_0.memory[21][7] ),
    .A2(_0329_),
    .A1(\charlie_0.memory[5][7] ));
 sg13g2_nand4_1 _3203_ (.B(_0439_),
    .C(_0441_),
    .A(_0336_),
    .Y(_0443_),
    .D(_0442_));
 sg13g2_a22oi_1 _3204_ (.Y(_0444_),
    .B1(_0345_),
    .B2(\charlie_0.memory[1][7] ),
    .A2(_0343_),
    .A1(\charlie_0.memory[12][7] ));
 sg13g2_nand4_1 _3205_ (.B(_0438_),
    .C(_0440_),
    .A(_0437_),
    .Y(_0445_),
    .D(_0444_));
 sg13g2_or3_1 _3206_ (.A(_0436_),
    .B(_0443_),
    .C(_0445_),
    .X(_0446_));
 sg13g2_a21oi_1 _3207_ (.A1(_0065_),
    .A2(net1026),
    .Y(_0447_),
    .B1(_0378_));
 sg13g2_a22oi_1 _3208_ (.Y(_0448_),
    .B1(_0357_),
    .B2(\charlie_0.memory[4][6] ),
    .A2(_0329_),
    .A1(\charlie_0.memory[5][6] ));
 sg13g2_a22oi_1 _3209_ (.Y(_0449_),
    .B1(_0350_),
    .B2(\charlie_0.memory[21][6] ),
    .A2(_0344_),
    .A1(\charlie_0.memory[14][6] ));
 sg13g2_a22oi_1 _3210_ (.Y(_0450_),
    .B1(_0355_),
    .B2(net1169),
    .A2(_0351_),
    .A1(\charlie_0.memory[11][6] ));
 sg13g2_a22oi_1 _3211_ (.Y(_0451_),
    .B1(_0345_),
    .B2(\charlie_0.memory[1][6] ),
    .A2(_0342_),
    .A1(\charlie_0.memory[15][6] ));
 sg13g2_a22oi_1 _3212_ (.Y(_0452_),
    .B1(_0354_),
    .B2(\charlie_0.memory[2][6] ),
    .A2(_0352_),
    .A1(\charlie_0.memory[6][6] ));
 sg13g2_a22oi_1 _3213_ (.Y(_0453_),
    .B1(_0356_),
    .B2(\charlie_0.memory[13][6] ),
    .A2(_0353_),
    .A1(\charlie_0.memory[18][6] ));
 sg13g2_a22oi_1 _3214_ (.Y(_0454_),
    .B1(_0358_),
    .B2(\charlie_0.memory[3][6] ),
    .A2(_0348_),
    .A1(\charlie_0.memory[22][6] ));
 sg13g2_a22oi_1 _3215_ (.Y(_0455_),
    .B1(_0347_),
    .B2(\charlie_0.memory[20][6] ),
    .A2(_0330_),
    .A1(\charlie_0.memory[10][6] ));
 sg13g2_a22oi_1 _3216_ (.Y(_0456_),
    .B1(_0343_),
    .B2(\charlie_0.memory[12][6] ),
    .A2(_0339_),
    .A1(\charlie_0.memory[19][6] ));
 sg13g2_a22oi_1 _3217_ (.Y(_0457_),
    .B1(_0349_),
    .B2(\charlie_0.memory[17][6] ),
    .A2(_0327_),
    .A1(\charlie_0.memory[8][6] ));
 sg13g2_nand4_1 _3218_ (.B(_0449_),
    .C(_0456_),
    .A(_0336_),
    .Y(_0458_),
    .D(_0457_));
 sg13g2_a22oi_1 _3219_ (.Y(_0459_),
    .B1(_0346_),
    .B2(\charlie_0.memory[7][6] ),
    .A2(_0325_),
    .A1(\charlie_0.memory[9][6] ));
 sg13g2_nand4_1 _3220_ (.B(_0451_),
    .C(_0455_),
    .A(_0450_),
    .Y(_0460_),
    .D(_0459_));
 sg13g2_nand4_1 _3221_ (.B(_0452_),
    .C(_0453_),
    .A(_0448_),
    .Y(_0461_),
    .D(_0454_));
 sg13g2_or3_1 _3222_ (.A(_0458_),
    .B(_0460_),
    .C(_0461_),
    .X(_0462_));
 sg13g2_a21oi_1 _3223_ (.A1(_0062_),
    .A2(net1026),
    .Y(_0463_),
    .B1(_0377_));
 sg13g2_a22oi_1 _3224_ (.Y(_0464_),
    .B1(_0356_),
    .B2(\charlie_0.memory[13][5] ),
    .A2(_0330_),
    .A1(\charlie_0.memory[10][5] ));
 sg13g2_a22oi_1 _3225_ (.Y(_0465_),
    .B1(_0345_),
    .B2(\charlie_0.memory[1][5] ),
    .A2(_0344_),
    .A1(\charlie_0.memory[14][5] ));
 sg13g2_a22oi_1 _3226_ (.Y(_0466_),
    .B1(_0358_),
    .B2(\charlie_0.memory[3][5] ),
    .A2(_0357_),
    .A1(\charlie_0.memory[4][5] ));
 sg13g2_a22oi_1 _3227_ (.Y(_0467_),
    .B1(_0350_),
    .B2(\charlie_0.memory[21][5] ),
    .A2(_0339_),
    .A1(\charlie_0.memory[19][5] ));
 sg13g2_a22oi_1 _3228_ (.Y(_0468_),
    .B1(_0354_),
    .B2(\charlie_0.memory[2][5] ),
    .A2(_0348_),
    .A1(\charlie_0.memory[22][5] ));
 sg13g2_a22oi_1 _3229_ (.Y(_0469_),
    .B1(_0347_),
    .B2(\charlie_0.memory[20][5] ),
    .A2(_0325_),
    .A1(\charlie_0.memory[9][5] ));
 sg13g2_a22oi_1 _3230_ (.Y(_0470_),
    .B1(_0355_),
    .B2(\charlie_0.memory[16][5] ),
    .A2(_0342_),
    .A1(\charlie_0.memory[15][5] ));
 sg13g2_nand4_1 _3231_ (.B(_0465_),
    .C(_0466_),
    .A(_0336_),
    .Y(_0471_),
    .D(_0470_));
 sg13g2_a22oi_1 _3232_ (.Y(_0472_),
    .B1(_0343_),
    .B2(\charlie_0.memory[12][5] ),
    .A2(_0329_),
    .A1(\charlie_0.memory[5][5] ));
 sg13g2_a22oi_1 _3233_ (.Y(_0473_),
    .B1(_0352_),
    .B2(\charlie_0.memory[6][5] ),
    .A2(_0346_),
    .A1(\charlie_0.memory[7][5] ));
 sg13g2_nand4_1 _3234_ (.B(_0467_),
    .C(_0472_),
    .A(_0464_),
    .Y(_0474_),
    .D(_0473_));
 sg13g2_a22oi_1 _3235_ (.Y(_0475_),
    .B1(_0353_),
    .B2(\charlie_0.memory[18][5] ),
    .A2(_0351_),
    .A1(\charlie_0.memory[11][5] ));
 sg13g2_a22oi_1 _3236_ (.Y(_0476_),
    .B1(_0349_),
    .B2(\charlie_0.memory[17][5] ),
    .A2(_0327_),
    .A1(\charlie_0.memory[8][5] ));
 sg13g2_nand4_1 _3237_ (.B(_0469_),
    .C(_0475_),
    .A(_0468_),
    .Y(_0477_),
    .D(_0476_));
 sg13g2_or3_1 _3238_ (.A(_0471_),
    .B(_0474_),
    .C(_0477_),
    .X(_0478_));
 sg13g2_a22oi_1 _3239_ (.Y(_0479_),
    .B1(_0339_),
    .B2(net1148),
    .A2(_0329_),
    .A1(\charlie_0.memory[5][4] ));
 sg13g2_a22oi_1 _3240_ (.Y(_0480_),
    .B1(_0344_),
    .B2(\charlie_0.memory[14][4] ),
    .A2(_0330_),
    .A1(\charlie_0.memory[10][4] ));
 sg13g2_a22oi_1 _3241_ (.Y(_0481_),
    .B1(_0351_),
    .B2(\charlie_0.memory[11][4] ),
    .A2(_0343_),
    .A1(\charlie_0.memory[12][4] ));
 sg13g2_nand4_1 _3242_ (.B(_0479_),
    .C(_0480_),
    .A(_0333_),
    .Y(_0482_),
    .D(_0481_));
 sg13g2_a22oi_1 _3243_ (.Y(_0483_),
    .B1(_0358_),
    .B2(\charlie_0.memory[3][4] ),
    .A2(_0327_),
    .A1(\charlie_0.memory[8][4] ));
 sg13g2_a22oi_1 _3244_ (.Y(_0484_),
    .B1(_0353_),
    .B2(\charlie_0.memory[18][4] ),
    .A2(_0345_),
    .A1(\charlie_0.memory[1][4] ));
 sg13g2_a22oi_1 _3245_ (.Y(_0485_),
    .B1(_0350_),
    .B2(\charlie_0.memory[21][4] ),
    .A2(_0347_),
    .A1(\charlie_0.memory[20][4] ));
 sg13g2_a22oi_1 _3246_ (.Y(_0486_),
    .B1(_0349_),
    .B2(\charlie_0.memory[17][4] ),
    .A2(_0348_),
    .A1(\charlie_0.memory[22][4] ));
 sg13g2_nand4_1 _3247_ (.B(_0484_),
    .C(_0485_),
    .A(_0483_),
    .Y(_0487_),
    .D(_0486_));
 sg13g2_a22oi_1 _3248_ (.Y(_0488_),
    .B1(_0354_),
    .B2(\charlie_0.memory[2][4] ),
    .A2(_0352_),
    .A1(\charlie_0.memory[6][4] ));
 sg13g2_a22oi_1 _3249_ (.Y(_0489_),
    .B1(_0356_),
    .B2(\charlie_0.memory[13][4] ),
    .A2(_0325_),
    .A1(\charlie_0.memory[9][4] ));
 sg13g2_a22oi_1 _3250_ (.Y(_0490_),
    .B1(_0357_),
    .B2(\charlie_0.memory[4][4] ),
    .A2(_0346_),
    .A1(\charlie_0.memory[7][4] ));
 sg13g2_a22oi_1 _3251_ (.Y(_0491_),
    .B1(_0355_),
    .B2(\charlie_0.memory[16][4] ),
    .A2(_0342_),
    .A1(\charlie_0.memory[15][4] ));
 sg13g2_nand4_1 _3252_ (.B(_0489_),
    .C(_0490_),
    .A(_0488_),
    .Y(_0492_),
    .D(_0491_));
 sg13g2_or3_1 _3253_ (.A(_0482_),
    .B(_0487_),
    .C(_0492_),
    .X(_0493_));
 sg13g2_a221oi_1 _3254_ (.B2(_0463_),
    .C1(_0375_),
    .B1(_0462_),
    .A1(_0446_),
    .Y(_0494_),
    .A2(_0447_));
 sg13g2_a21oi_1 _3255_ (.A1(_0061_),
    .A2(net1026),
    .Y(_0495_),
    .B1(_0378_));
 sg13g2_a21oi_1 _3256_ (.A1(_0060_),
    .A2(net1026),
    .Y(_0496_),
    .B1(_0377_));
 sg13g2_a221oi_1 _3257_ (.B2(_0493_),
    .C1(_0374_),
    .B1(_0496_),
    .A1(_0478_),
    .Y(_0497_),
    .A2(_0495_));
 sg13g2_nor3_1 _3258_ (.A(_0397_),
    .B(_0494_),
    .C(_0497_),
    .Y(_0498_));
 sg13g2_o21ai_1 _3259_ (.B1(_0322_),
    .Y(_0499_),
    .A1(_0431_),
    .A2(_0498_));
 sg13g2_a21oi_1 _3260_ (.A1(net1200),
    .A2(_1858_),
    .Y(_0500_),
    .B1(_0305_));
 sg13g2_nor2_1 _3261_ (.A(_0499_),
    .B(_0500_),
    .Y(_0000_));
 sg13g2_nor2_1 _3262_ (.A(net295),
    .B(_0305_),
    .Y(_0501_));
 sg13g2_nor4_1 _3263_ (.A(net295),
    .B(_1848_),
    .C(_0305_),
    .D(net952),
    .Y(_0502_));
 sg13g2_nor2_1 _3264_ (.A(net281),
    .B(net952),
    .Y(_0503_));
 sg13g2_a21o_1 _3265_ (.A2(_0502_),
    .A1(_1828_),
    .B1(_0503_),
    .X(_0001_));
 sg13g2_a21oi_1 _3266_ (.A1(_1828_),
    .A2(_0310_),
    .Y(_0504_),
    .B1(_0010_));
 sg13g2_nor2_1 _3267_ (.A(_0499_),
    .B(_0504_),
    .Y(_0002_));
 sg13g2_xnor2_1 _3268_ (.Y(_0505_),
    .A(net1207),
    .B(_1846_));
 sg13g2_xnor2_1 _3269_ (.Y(_0506_),
    .A(_1828_),
    .B(_1846_));
 sg13g2_nand3b_1 _3270_ (.B(_0501_),
    .C(_1848_),
    .Y(_0507_),
    .A_N(net952));
 sg13g2_or3_1 _3271_ (.A(_0315_),
    .B(_0317_),
    .C(net952),
    .X(_0508_));
 sg13g2_o21ai_1 _3272_ (.B1(_0508_),
    .Y(_0003_),
    .A1(_0506_),
    .A2(_0507_));
 sg13g2_a21oi_1 _3273_ (.A1(_0316_),
    .A2(_0318_),
    .Y(_0004_),
    .B1(net952));
 sg13g2_nor4_1 _3274_ (.A(net1200),
    .B(_0308_),
    .C(_0319_),
    .D(net952),
    .Y(_0509_));
 sg13g2_a21o_1 _3275_ (.A2(_0502_),
    .A1(net1207),
    .B1(_0509_),
    .X(_0005_));
 sg13g2_nor2_1 _3276_ (.A(_0320_),
    .B(_0014_),
    .Y(_0510_));
 sg13g2_nor2_1 _3277_ (.A(net952),
    .B(_0510_),
    .Y(_0006_));
 sg13g2_or3_1 _3278_ (.A(_0317_),
    .B(_0321_),
    .C(net952),
    .X(_0511_));
 sg13g2_o21ai_1 _3279_ (.B1(_0511_),
    .Y(_0007_),
    .A1(_0505_),
    .A2(_0507_));
 sg13g2_and2_1 _3280_ (.A(net1197),
    .B(net1232),
    .X(_0512_));
 sg13g2_nand2_1 _3281_ (.Y(_0513_),
    .A(net1199),
    .B(net1233));
 sg13g2_o21ai_1 _3282_ (.B1(net1196),
    .Y(_0514_),
    .A1(\charlie_0.memory[7][6] ),
    .A2(net1098));
 sg13g2_nor2b_1 _3283_ (.A(net1197),
    .B_N(net1231),
    .Y(_0515_));
 sg13g2_nand2_1 _3284_ (.Y(_0516_),
    .A(net1125),
    .B(net1233));
 sg13g2_nor2_1 _3285_ (.A(net1197),
    .B(net1231),
    .Y(_0517_));
 sg13g2_or2_1 _3286_ (.X(_0518_),
    .B(net1233),
    .A(net1199));
 sg13g2_nor2b_1 _3287_ (.A(net1231),
    .B_N(net1197),
    .Y(_0519_));
 sg13g2_nand2_2 _3288_ (.Y(_0520_),
    .A(net1199),
    .B(net1228));
 sg13g2_a22oi_1 _3289_ (.Y(_0521_),
    .B1(net1084),
    .B2(_1806_),
    .A2(net1091),
    .A1(_1808_));
 sg13g2_o21ai_1 _3290_ (.B1(_0521_),
    .Y(_0522_),
    .A1(\charlie_0.memory[5][6] ),
    .A2(net1024));
 sg13g2_nand2_2 _3291_ (.Y(_0523_),
    .A(net1138),
    .B(net1135));
 sg13g2_o21ai_1 _3292_ (.B1(net1132),
    .Y(_0524_),
    .A1(\charlie_0.memory[0][6] ),
    .A2(net1086));
 sg13g2_a221oi_1 _3293_ (.B2(_1812_),
    .C1(_0524_),
    .B1(net1084),
    .A1(_1816_),
    .Y(_0525_),
    .A2(net1097));
 sg13g2_o21ai_1 _3294_ (.B1(_0525_),
    .Y(_0526_),
    .A1(\charlie_0.memory[3][6] ),
    .A2(net1099));
 sg13g2_o21ai_1 _3295_ (.B1(_0526_),
    .Y(_0527_),
    .A1(_0514_),
    .A2(_0522_));
 sg13g2_nand2_1 _3296_ (.Y(_0528_),
    .A(net1191),
    .B(net1194));
 sg13g2_nand2_1 _3297_ (.Y(_0529_),
    .A(\charlie_0.memory[12][6] ),
    .B(net1088));
 sg13g2_nand2_1 _3298_ (.Y(_0530_),
    .A(net1191),
    .B(net1128));
 sg13g2_a22oi_1 _3299_ (.Y(_0531_),
    .B1(net1092),
    .B2(\charlie_0.memory[9][6] ),
    .A2(net1101),
    .A1(\charlie_0.memory[11][6] ));
 sg13g2_a221oi_1 _3300_ (.B2(\charlie_0.memory[10][6] ),
    .C1(net1192),
    .B1(net1080),
    .A1(\charlie_0.memory[8][6] ),
    .Y(_0532_),
    .A2(net1088));
 sg13g2_nand2_1 _3301_ (.Y(_0533_),
    .A(_0531_),
    .B(_0532_));
 sg13g2_a21oi_1 _3302_ (.A1(\charlie_0.memory[15][6] ),
    .A2(net1101),
    .Y(_0534_),
    .B1(net1128));
 sg13g2_a22oi_1 _3303_ (.Y(_0535_),
    .B1(net1081),
    .B2(\charlie_0.memory[14][6] ),
    .A2(net1092),
    .A1(\charlie_0.memory[13][6] ));
 sg13g2_nand3_1 _3304_ (.B(_0534_),
    .C(_0535_),
    .A(_0529_),
    .Y(_0536_));
 sg13g2_nand2_1 _3305_ (.Y(_0537_),
    .A(_0533_),
    .B(_0536_));
 sg13g2_mux4_1 _3306_ (.S0(net1232),
    .A0(net1169),
    .A1(\charlie_0.memory[17][6] ),
    .A2(\charlie_0.memory[18][6] ),
    .A3(\charlie_0.memory[19][6] ),
    .S1(net1199),
    .X(_0538_));
 sg13g2_a21oi_1 _3307_ (.A1(\charlie_0.memory[22][6] ),
    .A2(net1083),
    .Y(_0539_),
    .B1(net1129));
 sg13g2_a22oi_1 _3308_ (.Y(_0540_),
    .B1(net1091),
    .B2(\charlie_0.memory[20][6] ),
    .A2(net1094),
    .A1(\charlie_0.memory[21][6] ));
 sg13g2_a21oi_1 _3309_ (.A1(_0539_),
    .A2(_0540_),
    .Y(_0541_),
    .B1(\gen_priority_write_blocks[0].this_priority_write.data_bits[11] ));
 sg13g2_o21ai_1 _3310_ (.B1(_0541_),
    .Y(_0542_),
    .A1(net1193),
    .A2(_0538_));
 sg13g2_a22oi_1 _3311_ (.Y(_0543_),
    .B1(_0542_),
    .B2(net1188),
    .A2(_0537_),
    .A1(\gen_priority_write_blocks[0].this_priority_write.data_bits[11] ));
 sg13g2_nor2_1 _3312_ (.A(net1137),
    .B(net1135),
    .Y(_0544_));
 sg13g2_o21ai_1 _3313_ (.B1(_0543_),
    .Y(_0545_),
    .A1(_0523_),
    .A2(_0527_));
 sg13g2_nand3_1 _3314_ (.B(net1193),
    .C(net1102),
    .A(net1189),
    .Y(_0546_));
 sg13g2_nor3_1 _3315_ (.A(net1185),
    .B(net1187),
    .C(_0546_),
    .Y(_0547_));
 sg13g2_nor4_2 _3316_ (.A(net1185),
    .B(net1186),
    .C(_0544_),
    .Y(_0548_),
    .D(_0547_));
 sg13g2_nand2_1 _3317_ (.Y(_0549_),
    .A(\spi_slave_0.is_data_phase ),
    .B(_1824_));
 sg13g2_nor4_2 _3318_ (.A(net2),
    .B(_1825_),
    .C(net1),
    .Y(_0550_),
    .D(_0549_));
 sg13g2_nand2_1 _3319_ (.Y(_0551_),
    .A(\spi_slave_0.is_data_phase ),
    .B(net439));
 sg13g2_nor2b_1 _3320_ (.A(\spi_slave_0.spi_clk_prev ),
    .B_N(net2),
    .Y(_0552_));
 sg13g2_nor2b_2 _3321_ (.A(net1),
    .B_N(_0552_),
    .Y(_0553_));
 sg13g2_a21oi_2 _3322_ (.B1(_0550_),
    .Y(_0554_),
    .A2(_0553_),
    .A1(_0551_));
 sg13g2_nand3_1 _3323_ (.B(net292),
    .C(\spi_slave_0.bit_cnt[0] ),
    .A(net296),
    .Y(_0555_));
 sg13g2_inv_1 _3324_ (.Y(_0556_),
    .A(_0555_));
 sg13g2_nor2_2 _3325_ (.A(\spi_slave_0.is_data_phase ),
    .B(_0555_),
    .Y(_0557_));
 sg13g2_or2_2 _3326_ (.X(_0558_),
    .B(_0555_),
    .A(\spi_slave_0.is_data_phase ));
 sg13g2_nand3_1 _3327_ (.B(_0545_),
    .C(_0548_),
    .A(net301),
    .Y(_0559_));
 sg13g2_o21ai_1 _3328_ (.B1(_0559_),
    .Y(_0560_),
    .A1(net1184),
    .A2(_0557_));
 sg13g2_mux2_1 _3329_ (.A0(_0560_),
    .A1(net1145),
    .S(_0554_),
    .X(_0561_));
 sg13g2_nor2_1 _3330_ (.A(net1223),
    .B(_0561_),
    .Y(_0081_));
 sg13g2_and4_2 _3331_ (.A(\charlie_0.memory[20][2] ),
    .B(_0070_),
    .C(_2007_),
    .D(_2037_),
    .X(_0562_));
 sg13g2_nor4_2 _3332_ (.A(_1777_),
    .B(_0070_),
    .C(_2008_),
    .Y(_0563_),
    .D(_2037_));
 sg13g2_nor2_2 _3333_ (.A(_0562_),
    .B(_0563_),
    .Y(_0564_));
 sg13g2_or2_2 _3334_ (.X(_0565_),
    .B(_0563_),
    .A(_0562_));
 sg13g2_nor2b_1 _3335_ (.A(\charlie_0.memory[20][1] ),
    .B_N(\charlie_0.memory[20][0] ),
    .Y(_0566_));
 sg13g2_nand2_1 _3336_ (.Y(_0567_),
    .A(_0565_),
    .B(_0566_));
 sg13g2_nand2_1 _3337_ (.Y(_0568_),
    .A(_0562_),
    .B(_0566_));
 sg13g2_nor3_2 _3338_ (.A(\spi_address[1] ),
    .B(\spi_address[0] ),
    .C(_0074_),
    .Y(_0569_));
 sg13g2_nor2_1 _3339_ (.A(_0073_),
    .B(_0555_),
    .Y(_0570_));
 sg13g2_nand3_1 _3340_ (.B(_0553_),
    .C(_0570_),
    .A(\spi_slave_0.is_data_phase ),
    .Y(_0571_));
 sg13g2_nor3_2 _3341_ (.A(\spi_address[3] ),
    .B(net411),
    .C(_0571_),
    .Y(_0572_));
 sg13g2_and2_1 _3342_ (.A(_0569_),
    .B(_0572_),
    .X(_0573_));
 sg13g2_nor3_2 _3343_ (.A(\spi_address[3] ),
    .B(_0071_),
    .C(_0571_),
    .Y(_0574_));
 sg13g2_and2_1 _3344_ (.A(_0569_),
    .B(_0574_),
    .X(_0575_));
 sg13g2_a21oi_1 _3345_ (.A1(\charlie_0.memory[20][2] ),
    .A2(_0568_),
    .Y(_0576_),
    .B1(net998));
 sg13g2_a21oi_1 _3346_ (.A1(net288),
    .A2(net999),
    .Y(_0577_),
    .B1(net1223));
 sg13g2_nor2b_1 _3347_ (.A(_0576_),
    .B_N(_0577_),
    .Y(_0082_));
 sg13g2_and2_1 _3348_ (.A(net2),
    .B(net1237),
    .X(_0083_));
 sg13g2_a21oi_1 _3349_ (.A1(\charlie_0.memory[20][3] ),
    .A2(\charlie_0.memory[20][2] ),
    .Y(_0578_),
    .B1(_0567_));
 sg13g2_nor2b_1 _3350_ (.A(_0578_),
    .B_N(\charlie_0.memory[20][0] ),
    .Y(_0579_));
 sg13g2_o21ai_1 _3351_ (.B1(net1238),
    .Y(_0580_),
    .A1(net998),
    .A2(_0579_));
 sg13g2_a21oi_1 _3352_ (.A1(net1230),
    .A2(net998),
    .Y(_0084_),
    .B1(_0580_));
 sg13g2_and2_1 _3353_ (.A(net301),
    .B(_0557_),
    .X(_0581_));
 sg13g2_nand2_1 _3354_ (.Y(_0582_),
    .A(net301),
    .B(_0557_));
 sg13g2_o21ai_1 _3355_ (.B1(net1196),
    .Y(_0583_),
    .A1(\charlie_0.memory[7][0] ),
    .A2(net1098));
 sg13g2_nor2_1 _3356_ (.A(\charlie_0.memory[5][0] ),
    .B(net1024),
    .Y(_0584_));
 sg13g2_nor2_1 _3357_ (.A(\charlie_0.memory[4][0] ),
    .B(net1085),
    .Y(_0585_));
 sg13g2_nor2_1 _3358_ (.A(\charlie_0.memory[6][0] ),
    .B(net1079),
    .Y(_0586_));
 sg13g2_nor4_1 _3359_ (.A(_0583_),
    .B(_0584_),
    .C(_0585_),
    .D(_0586_),
    .Y(_0587_));
 sg13g2_o21ai_1 _3360_ (.B1(net1130),
    .Y(_0588_),
    .A1(\charlie_0.memory[1][0] ),
    .A2(net1025));
 sg13g2_nor2_1 _3361_ (.A(\charlie_0.memory[2][0] ),
    .B(net1079),
    .Y(_0589_));
 sg13g2_nor2_1 _3362_ (.A(\charlie_0.memory[0][0] ),
    .B(net1086),
    .Y(_0590_));
 sg13g2_nor2_1 _3363_ (.A(\charlie_0.memory[3][0] ),
    .B(net1099),
    .Y(_0591_));
 sg13g2_nor4_1 _3364_ (.A(_0588_),
    .B(_0589_),
    .C(_0590_),
    .D(_0591_),
    .Y(_0592_));
 sg13g2_nor3_2 _3365_ (.A(_0523_),
    .B(_0587_),
    .C(_0592_),
    .Y(_0593_));
 sg13g2_a22oi_1 _3366_ (.Y(_0594_),
    .B1(net1089),
    .B2(\charlie_0.memory[20][0] ),
    .A2(net1094),
    .A1(\charlie_0.memory[21][0] ));
 sg13g2_nand2_1 _3367_ (.Y(_0595_),
    .A(net1146),
    .B(net1083));
 sg13g2_a21oi_1 _3368_ (.A1(_0594_),
    .A2(_0595_),
    .Y(_0596_),
    .B1(net1127));
 sg13g2_a22oi_1 _3369_ (.Y(_0597_),
    .B1(net1084),
    .B2(\charlie_0.memory[18][0] ),
    .A2(net1097),
    .A1(net1164));
 sg13g2_a22oi_1 _3370_ (.Y(_0598_),
    .B1(net1090),
    .B2(net1174),
    .A2(net1102),
    .A1(net1155));
 sg13g2_a21oi_1 _3371_ (.A1(_0597_),
    .A2(_0598_),
    .Y(_0599_),
    .B1(net1192));
 sg13g2_nor2_1 _3372_ (.A(_0596_),
    .B(_0599_),
    .Y(_0600_));
 sg13g2_a22oi_1 _3373_ (.Y(_0601_),
    .B1(net1092),
    .B2(\charlie_0.memory[9][0] ),
    .A2(net1101),
    .A1(\charlie_0.memory[11][0] ));
 sg13g2_a22oi_1 _3374_ (.Y(_0602_),
    .B1(net1081),
    .B2(\charlie_0.memory[10][0] ),
    .A2(net1088),
    .A1(\charlie_0.memory[8][0] ));
 sg13g2_a21oi_1 _3375_ (.A1(_0601_),
    .A2(_0602_),
    .Y(_0603_),
    .B1(net1192));
 sg13g2_a22oi_1 _3376_ (.Y(_0604_),
    .B1(net1093),
    .B2(\charlie_0.memory[13][0] ),
    .A2(net1100),
    .A1(\charlie_0.memory[15][0] ));
 sg13g2_a22oi_1 _3377_ (.Y(_0605_),
    .B1(net1080),
    .B2(\charlie_0.memory[14][0] ),
    .A2(net1087),
    .A1(\charlie_0.memory[12][0] ));
 sg13g2_a21oi_1 _3378_ (.A1(_0604_),
    .A2(_0605_),
    .Y(_0606_),
    .B1(net1128));
 sg13g2_nor2_1 _3379_ (.A(_0603_),
    .B(_0606_),
    .Y(_0607_));
 sg13g2_a221oi_1 _3380_ (.B2(net1190),
    .C1(_0593_),
    .B1(_0607_),
    .A1(net1188),
    .Y(_0608_),
    .A2(_0600_));
 sg13g2_nand2b_1 _3381_ (.Y(_0609_),
    .B(_0548_),
    .A_N(_0608_));
 sg13g2_a21o_2 _3382_ (.A2(_0557_),
    .A1(net1214),
    .B1(_0554_),
    .X(_0610_));
 sg13g2_a21oi_2 _3383_ (.B1(_0554_),
    .Y(_0611_),
    .A2(_0557_),
    .A1(net1214));
 sg13g2_a221oi_1 _3384_ (.B2(_0609_),
    .C1(_0610_),
    .B1(_0581_),
    .A1(net1232),
    .Y(_0612_),
    .A2(_0558_));
 sg13g2_o21ai_1 _3385_ (.B1(net1235),
    .Y(_0613_),
    .A1(net1198),
    .A2(_0611_));
 sg13g2_nor2_1 _3386_ (.A(_0612_),
    .B(_0613_),
    .Y(_0085_));
 sg13g2_a21oi_1 _3387_ (.A1(net1133),
    .A2(_0547_),
    .Y(_0614_),
    .B1(_0582_));
 sg13g2_o21ai_1 _3388_ (.B1(net1195),
    .Y(_0615_),
    .A1(\charlie_0.memory[4][1] ),
    .A2(net1085));
 sg13g2_nor2_1 _3389_ (.A(\charlie_0.memory[7][1] ),
    .B(net1098),
    .Y(_0616_));
 sg13g2_nor2_1 _3390_ (.A(\charlie_0.memory[6][1] ),
    .B(net1079),
    .Y(_0617_));
 sg13g2_nor2_1 _3391_ (.A(\charlie_0.memory[5][1] ),
    .B(net1024),
    .Y(_0618_));
 sg13g2_nor4_2 _3392_ (.A(_0615_),
    .B(_0616_),
    .C(_0617_),
    .Y(_0619_),
    .D(_0618_));
 sg13g2_o21ai_1 _3393_ (.B1(net1130),
    .Y(_0620_),
    .A1(\charlie_0.memory[1][1] ),
    .A2(net1025));
 sg13g2_nor2_1 _3394_ (.A(\charlie_0.memory[3][1] ),
    .B(net1099),
    .Y(_0621_));
 sg13g2_nor2_1 _3395_ (.A(\charlie_0.memory[2][1] ),
    .B(net1078),
    .Y(_0622_));
 sg13g2_nor2_1 _3396_ (.A(\charlie_0.memory[0][1] ),
    .B(net1086),
    .Y(_0623_));
 sg13g2_nor4_1 _3397_ (.A(_0620_),
    .B(_0621_),
    .C(_0622_),
    .D(_0623_),
    .Y(_0624_));
 sg13g2_nor3_2 _3398_ (.A(_0523_),
    .B(_0619_),
    .C(_0624_),
    .Y(_0625_));
 sg13g2_nand2_1 _3399_ (.Y(_0626_),
    .A(\charlie_0.memory[21][1] ),
    .B(net1096));
 sg13g2_a22oi_1 _3400_ (.Y(_0627_),
    .B1(net1083),
    .B2(\charlie_0.memory[22][1] ),
    .A2(net1089),
    .A1(\charlie_0.memory[20][1] ));
 sg13g2_a21oi_1 _3401_ (.A1(_0626_),
    .A2(_0627_),
    .Y(_0628_),
    .B1(net1127));
 sg13g2_a22oi_1 _3402_ (.Y(_0629_),
    .B1(net1089),
    .B2(net1171),
    .A2(net1102),
    .A1(net1154));
 sg13g2_a22oi_1 _3403_ (.Y(_0630_),
    .B1(net1082),
    .B2(\charlie_0.memory[18][1] ),
    .A2(net1095),
    .A1(net1162));
 sg13g2_a21oi_1 _3404_ (.A1(_0629_),
    .A2(_0630_),
    .Y(_0631_),
    .B1(net1192));
 sg13g2_nor2_1 _3405_ (.A(_0628_),
    .B(_0631_),
    .Y(_0632_));
 sg13g2_a22oi_1 _3406_ (.Y(_0633_),
    .B1(net1092),
    .B2(\charlie_0.memory[9][1] ),
    .A2(net1100),
    .A1(\charlie_0.memory[11][1] ));
 sg13g2_a22oi_1 _3407_ (.Y(_0634_),
    .B1(net1080),
    .B2(\charlie_0.memory[10][1] ),
    .A2(net1087),
    .A1(\charlie_0.memory[8][1] ));
 sg13g2_a21oi_1 _3408_ (.A1(_0633_),
    .A2(_0634_),
    .Y(_0635_),
    .B1(net1192));
 sg13g2_a22oi_1 _3409_ (.Y(_0636_),
    .B1(net1088),
    .B2(\charlie_0.memory[12][1] ),
    .A2(net1093),
    .A1(\charlie_0.memory[13][1] ));
 sg13g2_a22oi_1 _3410_ (.Y(_0637_),
    .B1(net1080),
    .B2(\charlie_0.memory[14][1] ),
    .A2(net1100),
    .A1(\charlie_0.memory[15][1] ));
 sg13g2_a21oi_1 _3411_ (.A1(_0636_),
    .A2(_0637_),
    .Y(_0638_),
    .B1(net1128));
 sg13g2_nor2_1 _3412_ (.A(_0635_),
    .B(_0638_),
    .Y(_0639_));
 sg13g2_a22oi_1 _3413_ (.Y(_0640_),
    .B1(_0639_),
    .B2(net1190),
    .A2(_0632_),
    .A1(net1188));
 sg13g2_inv_1 _3414_ (.Y(_0641_),
    .A(_0640_));
 sg13g2_o21ai_1 _3415_ (.B1(_0548_),
    .Y(_0642_),
    .A1(_0625_),
    .A2(_0641_));
 sg13g2_a221oi_1 _3416_ (.B2(_0642_),
    .C1(_0610_),
    .B1(_0614_),
    .A1(net1198),
    .Y(_0643_),
    .A2(_0558_));
 sg13g2_o21ai_1 _3417_ (.B1(net1235),
    .Y(_0644_),
    .A1(net1193),
    .A2(_0611_));
 sg13g2_nor2_1 _3418_ (.A(_0643_),
    .B(_0644_),
    .Y(_0086_));
 sg13g2_a21oi_1 _3419_ (.A1(\charlie_0.memory[22][2] ),
    .A2(net1082),
    .Y(_0645_),
    .B1(net1129));
 sg13g2_a22oi_1 _3420_ (.Y(_0646_),
    .B1(net1089),
    .B2(\charlie_0.memory[20][2] ),
    .A2(net1094),
    .A1(\charlie_0.memory[21][2] ));
 sg13g2_a22oi_1 _3421_ (.Y(_0647_),
    .B1(net1094),
    .B2(net1158),
    .A2(net1103),
    .A1(net1151));
 sg13g2_a221oi_1 _3422_ (.B2(\charlie_0.memory[18][2] ),
    .C1(net1192),
    .B1(net1083),
    .A1(\charlie_0.memory[16][2] ),
    .Y(_0648_),
    .A2(net1089));
 sg13g2_a22oi_1 _3423_ (.Y(_0649_),
    .B1(_0647_),
    .B2(_0648_),
    .A2(_0646_),
    .A1(_0645_));
 sg13g2_o21ai_1 _3424_ (.B1(net1195),
    .Y(_0650_),
    .A1(\charlie_0.memory[5][2] ),
    .A2(net1024));
 sg13g2_nor2_1 _3425_ (.A(\charlie_0.memory[7][2] ),
    .B(net1098),
    .Y(_0651_));
 sg13g2_nor2_1 _3426_ (.A(\charlie_0.memory[6][2] ),
    .B(net1078),
    .Y(_0652_));
 sg13g2_nor2_1 _3427_ (.A(\charlie_0.memory[4][2] ),
    .B(net1085),
    .Y(_0653_));
 sg13g2_nor4_2 _3428_ (.A(_0650_),
    .B(_0651_),
    .C(_0652_),
    .Y(_0654_),
    .D(_0653_));
 sg13g2_o21ai_1 _3429_ (.B1(net1131),
    .Y(_0655_),
    .A1(\charlie_0.memory[3][2] ),
    .A2(net1099));
 sg13g2_nor2_1 _3430_ (.A(\charlie_0.memory[0][2] ),
    .B(net1086),
    .Y(_0656_));
 sg13g2_nor2_1 _3431_ (.A(\charlie_0.memory[2][2] ),
    .B(net1078),
    .Y(_0657_));
 sg13g2_nor2_1 _3432_ (.A(\charlie_0.memory[1][2] ),
    .B(net1025),
    .Y(_0658_));
 sg13g2_nor4_1 _3433_ (.A(_0655_),
    .B(_0656_),
    .C(_0657_),
    .D(_0658_),
    .Y(_0659_));
 sg13g2_nor3_2 _3434_ (.A(_0523_),
    .B(_0654_),
    .C(_0659_),
    .Y(_0660_));
 sg13g2_a22oi_1 _3435_ (.Y(_0661_),
    .B1(net1088),
    .B2(\charlie_0.memory[12][2] ),
    .A2(net1096),
    .A1(\charlie_0.memory[13][2] ));
 sg13g2_a22oi_1 _3436_ (.Y(_0662_),
    .B1(net1081),
    .B2(\charlie_0.memory[14][2] ),
    .A2(net1103),
    .A1(\charlie_0.memory[15][2] ));
 sg13g2_a21oi_1 _3437_ (.A1(_0661_),
    .A2(_0662_),
    .Y(_0663_),
    .B1(net1128));
 sg13g2_a22oi_1 _3438_ (.Y(_0664_),
    .B1(net1081),
    .B2(\charlie_0.memory[10][2] ),
    .A2(net1103),
    .A1(\charlie_0.memory[11][2] ));
 sg13g2_a22oi_1 _3439_ (.Y(_0665_),
    .B1(net1088),
    .B2(\charlie_0.memory[8][2] ),
    .A2(net1093),
    .A1(\charlie_0.memory[9][2] ));
 sg13g2_a21oi_1 _3440_ (.A1(_0664_),
    .A2(_0665_),
    .Y(_0666_),
    .B1(net1192));
 sg13g2_or3_1 _3441_ (.A(net1133),
    .B(_0663_),
    .C(_0666_),
    .X(_0667_));
 sg13g2_o21ai_1 _3442_ (.B1(_0667_),
    .Y(_0668_),
    .A1(net1136),
    .A2(_0649_));
 sg13g2_o21ai_1 _3443_ (.B1(_0548_),
    .Y(_0669_),
    .A1(_0660_),
    .A2(_0668_));
 sg13g2_a221oi_1 _3444_ (.B2(_0669_),
    .C1(_0610_),
    .B1(_0581_),
    .A1(net1193),
    .Y(_0670_),
    .A2(_0558_));
 sg13g2_o21ai_1 _3445_ (.B1(net1237),
    .Y(_0671_),
    .A1(net1190),
    .A2(_0611_));
 sg13g2_nor2_1 _3446_ (.A(_0670_),
    .B(_0671_),
    .Y(_0087_));
 sg13g2_a22oi_1 _3447_ (.Y(_0672_),
    .B1(net1087),
    .B2(\charlie_0.memory[12][3] ),
    .A2(net1100),
    .A1(\charlie_0.memory[15][3] ));
 sg13g2_a221oi_1 _3448_ (.B2(\charlie_0.memory[14][3] ),
    .C1(_0528_),
    .B1(net1081),
    .A1(\charlie_0.memory[13][3] ),
    .Y(_0673_),
    .A2(net1093));
 sg13g2_a21oi_1 _3449_ (.A1(\charlie_0.memory[9][3] ),
    .A2(net1093),
    .Y(_0674_),
    .B1(_0530_));
 sg13g2_nor2_1 _3450_ (.A(_1799_),
    .B(_0520_),
    .Y(_0675_));
 sg13g2_a221oi_1 _3451_ (.B2(\charlie_0.memory[8][3] ),
    .C1(_0675_),
    .B1(net1088),
    .A1(\charlie_0.memory[11][3] ),
    .Y(_0676_),
    .A2(net1100));
 sg13g2_a22oi_1 _3452_ (.Y(_0677_),
    .B1(_0674_),
    .B2(_0676_),
    .A2(_0673_),
    .A1(_0672_));
 sg13g2_o21ai_1 _3453_ (.B1(net1195),
    .Y(_0678_),
    .A1(\charlie_0.memory[5][3] ),
    .A2(net1024));
 sg13g2_nor2_1 _3454_ (.A(\charlie_0.memory[4][3] ),
    .B(net1085),
    .Y(_0679_));
 sg13g2_nor2_1 _3455_ (.A(\charlie_0.memory[6][3] ),
    .B(net1078),
    .Y(_0680_));
 sg13g2_nor3_1 _3456_ (.A(_0678_),
    .B(_0679_),
    .C(_0680_),
    .Y(_0681_));
 sg13g2_o21ai_1 _3457_ (.B1(_0681_),
    .Y(_0682_),
    .A1(\charlie_0.memory[7][3] ),
    .A2(net1098));
 sg13g2_o21ai_1 _3458_ (.B1(net1131),
    .Y(_0683_),
    .A1(\charlie_0.memory[3][3] ),
    .A2(net1098));
 sg13g2_nor2_1 _3459_ (.A(\charlie_0.memory[1][3] ),
    .B(net1025),
    .Y(_0684_));
 sg13g2_nor2_1 _3460_ (.A(\charlie_0.memory[2][3] ),
    .B(net1078),
    .Y(_0685_));
 sg13g2_nor2_1 _3461_ (.A(\charlie_0.memory[0][3] ),
    .B(net1086),
    .Y(_0686_));
 sg13g2_nor4_2 _3462_ (.A(_0683_),
    .B(_0684_),
    .C(_0685_),
    .Y(_0687_),
    .D(_0686_));
 sg13g2_nor2_1 _3463_ (.A(net1190),
    .B(_0687_),
    .Y(_0688_));
 sg13g2_a21oi_1 _3464_ (.A1(_0682_),
    .A2(_0688_),
    .Y(_0689_),
    .B1(net1188));
 sg13g2_a22oi_1 _3465_ (.Y(_0690_),
    .B1(net1091),
    .B2(\charlie_0.memory[16][3] ),
    .A2(net1103),
    .A1(net1150));
 sg13g2_a221oi_1 _3466_ (.B2(\charlie_0.memory[18][3] ),
    .C1(net1196),
    .B1(net1084),
    .A1(net1156),
    .Y(_0691_),
    .A2(net1097));
 sg13g2_a21oi_1 _3467_ (.A1(\charlie_0.memory[22][3] ),
    .A2(net1082),
    .Y(_0692_),
    .B1(net1129));
 sg13g2_a22oi_1 _3468_ (.Y(_0693_),
    .B1(net1090),
    .B2(\charlie_0.memory[20][3] ),
    .A2(net1095),
    .A1(\charlie_0.memory[21][3] ));
 sg13g2_a221oi_1 _3469_ (.B2(_0693_),
    .C1(net1137),
    .B1(_0692_),
    .A1(_0690_),
    .Y(_0694_),
    .A2(_0691_));
 sg13g2_o21ai_1 _3470_ (.B1(_0677_),
    .Y(_0695_),
    .A1(_0689_),
    .A2(_0694_));
 sg13g2_nand2_1 _3471_ (.Y(_0696_),
    .A(_0548_),
    .B(_0695_));
 sg13g2_a221oi_1 _3472_ (.B2(_0696_),
    .C1(_0610_),
    .B1(_0614_),
    .A1(net1190),
    .Y(_0697_),
    .A2(_0558_));
 sg13g2_o21ai_1 _3473_ (.B1(net1235),
    .Y(_0698_),
    .A1(net303),
    .A2(_0611_));
 sg13g2_nor2_1 _3474_ (.A(_0697_),
    .B(_0698_),
    .Y(_0088_));
 sg13g2_nand2_1 _3475_ (.Y(_0699_),
    .A(\charlie_0.memory[20][4] ),
    .B(net1090));
 sg13g2_a22oi_1 _3476_ (.Y(_0700_),
    .B1(net1084),
    .B2(\charlie_0.memory[18][4] ),
    .A2(net1097),
    .A1(\charlie_0.memory[17][4] ));
 sg13g2_a22oi_1 _3477_ (.Y(_0701_),
    .B1(net1082),
    .B2(\charlie_0.memory[22][4] ),
    .A2(net1094),
    .A1(\charlie_0.memory[21][4] ));
 sg13g2_a21oi_1 _3478_ (.A1(_0699_),
    .A2(_0701_),
    .Y(_0702_),
    .B1(net1127));
 sg13g2_a22oi_1 _3479_ (.Y(_0703_),
    .B1(net1087),
    .B2(\charlie_0.memory[16][4] ),
    .A2(net1100),
    .A1(net1148));
 sg13g2_a21oi_1 _3480_ (.A1(_0700_),
    .A2(_0703_),
    .Y(_0704_),
    .B1(net1192));
 sg13g2_or3_1 _3481_ (.A(net1136),
    .B(_0702_),
    .C(_0704_),
    .X(_0705_));
 sg13g2_o21ai_1 _3482_ (.B1(net1195),
    .Y(_0706_),
    .A1(\charlie_0.memory[7][4] ),
    .A2(net1098));
 sg13g2_nor2_1 _3483_ (.A(\charlie_0.memory[4][4] ),
    .B(net1085),
    .Y(_0707_));
 sg13g2_nor2_1 _3484_ (.A(\charlie_0.memory[6][4] ),
    .B(net1078),
    .Y(_0708_));
 sg13g2_nor2_1 _3485_ (.A(\charlie_0.memory[5][4] ),
    .B(net1024),
    .Y(_0709_));
 sg13g2_nor4_1 _3486_ (.A(_0706_),
    .B(_0707_),
    .C(_0708_),
    .D(_0709_),
    .Y(_0710_));
 sg13g2_o21ai_1 _3487_ (.B1(net1130),
    .Y(_0711_),
    .A1(\charlie_0.memory[3][4] ),
    .A2(net1098));
 sg13g2_a22oi_1 _3488_ (.Y(_0712_),
    .B1(net1084),
    .B2(_1814_),
    .A2(net1091),
    .A1(_1817_));
 sg13g2_o21ai_1 _3489_ (.B1(_0712_),
    .Y(_0713_),
    .A1(\charlie_0.memory[1][4] ),
    .A2(net1025));
 sg13g2_nor2_1 _3490_ (.A(_0711_),
    .B(_0713_),
    .Y(_0714_));
 sg13g2_or3_1 _3491_ (.A(_0523_),
    .B(_0710_),
    .C(_0714_),
    .X(_0715_));
 sg13g2_a21oi_1 _3492_ (.A1(\charlie_0.memory[13][4] ),
    .A2(net1092),
    .Y(_0716_),
    .B1(_0528_));
 sg13g2_nand2_1 _3493_ (.Y(_0717_),
    .A(\charlie_0.memory[14][4] ),
    .B(net1080));
 sg13g2_a22oi_1 _3494_ (.Y(_0718_),
    .B1(net1087),
    .B2(\charlie_0.memory[12][4] ),
    .A2(net1101),
    .A1(\charlie_0.memory[15][4] ));
 sg13g2_nand3_1 _3495_ (.B(_0717_),
    .C(_0718_),
    .A(_0716_),
    .Y(_0719_));
 sg13g2_a21oi_1 _3496_ (.A1(\charlie_0.memory[11][4] ),
    .A2(net1100),
    .Y(_0720_),
    .B1(_0530_));
 sg13g2_nand2_1 _3497_ (.Y(_0721_),
    .A(\charlie_0.memory[8][4] ),
    .B(net1087));
 sg13g2_a22oi_1 _3498_ (.Y(_0722_),
    .B1(net1080),
    .B2(\charlie_0.memory[10][4] ),
    .A2(net1092),
    .A1(\charlie_0.memory[9][4] ));
 sg13g2_nand3_1 _3499_ (.B(_0721_),
    .C(_0722_),
    .A(_0720_),
    .Y(_0723_));
 sg13g2_nand4_1 _3500_ (.B(_0715_),
    .C(_0719_),
    .A(_0705_),
    .Y(_0724_),
    .D(_0723_));
 sg13g2_nand2_1 _3501_ (.Y(_0725_),
    .A(_0548_),
    .B(_0724_));
 sg13g2_a221oi_1 _3502_ (.B2(_0725_),
    .C1(_0610_),
    .B1(_0614_),
    .A1(net1188),
    .Y(_0726_),
    .A2(_0558_));
 sg13g2_o21ai_1 _3503_ (.B1(net1235),
    .Y(_0727_),
    .A1(net1186),
    .A2(_0611_));
 sg13g2_nor2_1 _3504_ (.A(_0726_),
    .B(_0727_),
    .Y(_0089_));
 sg13g2_a22oi_1 _3505_ (.Y(_0728_),
    .B1(net1090),
    .B2(\charlie_0.memory[16][5] ),
    .A2(net1095),
    .A1(\charlie_0.memory[17][5] ));
 sg13g2_a221oi_1 _3506_ (.B2(\charlie_0.memory[18][5] ),
    .C1(net1196),
    .B1(net1082),
    .A1(\charlie_0.memory[19][5] ),
    .Y(_0729_),
    .A2(net1103));
 sg13g2_a21oi_1 _3507_ (.A1(\charlie_0.memory[21][5] ),
    .A2(net1094),
    .Y(_0730_),
    .B1(net1127));
 sg13g2_a22oi_1 _3508_ (.Y(_0731_),
    .B1(net1082),
    .B2(\charlie_0.memory[22][5] ),
    .A2(net1090),
    .A1(\charlie_0.memory[20][5] ));
 sg13g2_a22oi_1 _3509_ (.Y(_0732_),
    .B1(_0730_),
    .B2(_0731_),
    .A2(_0729_),
    .A1(_0728_));
 sg13g2_nor2_1 _3510_ (.A(net1136),
    .B(_0732_),
    .Y(_0733_));
 sg13g2_nand2b_1 _3511_ (.Y(_0734_),
    .B(net1104),
    .A_N(\charlie_0.memory[3][5] ));
 sg13g2_o21ai_1 _3512_ (.B1(_0734_),
    .Y(_0735_),
    .A1(\charlie_0.memory[1][5] ),
    .A2(net1024));
 sg13g2_a21oi_1 _3513_ (.A1(_1813_),
    .A2(net1084),
    .Y(_0736_),
    .B1(net1196));
 sg13g2_o21ai_1 _3514_ (.B1(_0736_),
    .Y(_0737_),
    .A1(\charlie_0.memory[0][5] ),
    .A2(net1085));
 sg13g2_o21ai_1 _3515_ (.B1(net1195),
    .Y(_0738_),
    .A1(\charlie_0.memory[6][5] ),
    .A2(net1078));
 sg13g2_a221oi_1 _3516_ (.B2(_1809_),
    .C1(_0738_),
    .B1(net1091),
    .A1(_1805_),
    .Y(_0739_),
    .A2(net1104));
 sg13g2_o21ai_1 _3517_ (.B1(_0739_),
    .Y(_0740_),
    .A1(\charlie_0.memory[5][5] ),
    .A2(net1024));
 sg13g2_o21ai_1 _3518_ (.B1(_0740_),
    .Y(_0741_),
    .A1(_0735_),
    .A2(_0737_));
 sg13g2_a22oi_1 _3519_ (.Y(_0742_),
    .B1(net1081),
    .B2(\charlie_0.memory[10][5] ),
    .A2(net1089),
    .A1(\charlie_0.memory[8][5] ));
 sg13g2_a221oi_1 _3520_ (.B2(\charlie_0.memory[9][5] ),
    .C1(_0530_),
    .B1(net1093),
    .A1(\charlie_0.memory[11][5] ),
    .Y(_0743_),
    .A2(net1100));
 sg13g2_a21oi_1 _3521_ (.A1(\charlie_0.memory[12][5] ),
    .A2(net1089),
    .Y(_0744_),
    .B1(_0528_));
 sg13g2_nor2_1 _3522_ (.A(_1794_),
    .B(_0520_),
    .Y(_0745_));
 sg13g2_a221oi_1 _3523_ (.B2(\charlie_0.memory[13][5] ),
    .C1(_0745_),
    .B1(net1093),
    .A1(\charlie_0.memory[15][5] ),
    .Y(_0746_),
    .A2(net1103));
 sg13g2_a22oi_1 _3524_ (.Y(_0747_),
    .B1(_0744_),
    .B2(_0746_),
    .A2(_0743_),
    .A1(_0742_));
 sg13g2_o21ai_1 _3525_ (.B1(_0747_),
    .Y(_0748_),
    .A1(_0523_),
    .A2(_0741_));
 sg13g2_o21ai_1 _3526_ (.B1(_0548_),
    .Y(_0749_),
    .A1(_0733_),
    .A2(_0748_));
 sg13g2_a221oi_1 _3527_ (.B2(_0749_),
    .C1(_0610_),
    .B1(_0581_),
    .A1(net1186),
    .Y(_0750_),
    .A2(_0558_));
 sg13g2_o21ai_1 _3528_ (.B1(net1235),
    .Y(_0751_),
    .A1(net1184),
    .A2(_0611_));
 sg13g2_nor2_1 _3529_ (.A(_0750_),
    .B(_0751_),
    .Y(_0090_));
 sg13g2_o21ai_1 _3530_ (.B1(net1131),
    .Y(_0752_),
    .A1(\charlie_0.memory[0][7] ),
    .A2(net1085));
 sg13g2_a22oi_1 _3531_ (.Y(_0753_),
    .B1(net1097),
    .B2(_1815_),
    .A2(net1104),
    .A1(_1810_));
 sg13g2_o21ai_1 _3532_ (.B1(_0753_),
    .Y(_0754_),
    .A1(\charlie_0.memory[2][7] ),
    .A2(net1079));
 sg13g2_o21ai_1 _3533_ (.B1(net1195),
    .Y(_0755_),
    .A1(\charlie_0.memory[4][7] ),
    .A2(net1085));
 sg13g2_a221oi_1 _3534_ (.B2(_1807_),
    .C1(_0755_),
    .B1(net1097),
    .A1(_1803_),
    .Y(_0756_),
    .A2(net1104));
 sg13g2_o21ai_1 _3535_ (.B1(_0756_),
    .Y(_0757_),
    .A1(\charlie_0.memory[6][7] ),
    .A2(net1078));
 sg13g2_o21ai_1 _3536_ (.B1(_0757_),
    .Y(_0758_),
    .A1(_0752_),
    .A2(_0754_));
 sg13g2_a22oi_1 _3537_ (.Y(_0759_),
    .B1(net1080),
    .B2(\charlie_0.memory[14][7] ),
    .A2(net1087),
    .A1(\charlie_0.memory[12][7] ));
 sg13g2_a22oi_1 _3538_ (.Y(_0760_),
    .B1(net1080),
    .B2(\charlie_0.memory[10][7] ),
    .A2(net1087),
    .A1(\charlie_0.memory[8][7] ));
 sg13g2_a22oi_1 _3539_ (.Y(_0761_),
    .B1(net1092),
    .B2(\charlie_0.memory[9][7] ),
    .A2(net1101),
    .A1(\charlie_0.memory[11][7] ));
 sg13g2_a21oi_1 _3540_ (.A1(_0760_),
    .A2(_0761_),
    .Y(_0762_),
    .B1(net1194));
 sg13g2_a22oi_1 _3541_ (.Y(_0763_),
    .B1(net1092),
    .B2(\charlie_0.memory[13][7] ),
    .A2(net1101),
    .A1(\charlie_0.memory[15][7] ));
 sg13g2_a21oi_1 _3542_ (.A1(_0759_),
    .A2(_0763_),
    .Y(_0764_),
    .B1(net1128));
 sg13g2_nor2_1 _3543_ (.A(_0762_),
    .B(_0764_),
    .Y(_0765_));
 sg13g2_a22oi_1 _3544_ (.Y(_0766_),
    .B1(net1094),
    .B2(\charlie_0.memory[17][7] ),
    .A2(net1103),
    .A1(\charlie_0.memory[19][7] ));
 sg13g2_a221oi_1 _3545_ (.B2(\charlie_0.memory[18][7] ),
    .C1(net1196),
    .B1(net1082),
    .A1(\charlie_0.memory[16][7] ),
    .Y(_0767_),
    .A2(net1090));
 sg13g2_a22oi_1 _3546_ (.Y(_0768_),
    .B1(net1090),
    .B2(\charlie_0.memory[20][7] ),
    .A2(net1094),
    .A1(\charlie_0.memory[21][7] ));
 sg13g2_a21oi_1 _3547_ (.A1(\charlie_0.memory[22][7] ),
    .A2(net1082),
    .Y(_0769_),
    .B1(net1127));
 sg13g2_a22oi_1 _3548_ (.Y(_0770_),
    .B1(_0768_),
    .B2(_0769_),
    .A2(_0767_),
    .A1(_0766_));
 sg13g2_nor2_1 _3549_ (.A(net1136),
    .B(_0770_),
    .Y(_0771_));
 sg13g2_a21oi_1 _3550_ (.A1(net1190),
    .A2(_0765_),
    .Y(_0772_),
    .B1(_0771_));
 sg13g2_o21ai_1 _3551_ (.B1(_0772_),
    .Y(_0773_),
    .A1(_0523_),
    .A2(_0758_));
 sg13g2_a21oi_1 _3552_ (.A1(_0548_),
    .A2(_0773_),
    .Y(_0774_),
    .B1(_0582_));
 sg13g2_nor3_1 _3553_ (.A(net1213),
    .B(_0554_),
    .C(_0774_),
    .Y(_0775_));
 sg13g2_o21ai_1 _3554_ (.B1(net1237),
    .Y(_0776_),
    .A1(net284),
    .A2(_0611_));
 sg13g2_nor2_1 _3555_ (.A(net302),
    .B(_0776_),
    .Y(_0091_));
 sg13g2_nand2_2 _3556_ (.Y(_0777_),
    .A(_0553_),
    .B(_0557_));
 sg13g2_nor2_2 _3557_ (.A(net299),
    .B(_0777_),
    .Y(_0778_));
 sg13g2_o21ai_1 _3558_ (.B1(net1234),
    .Y(_0779_),
    .A1(net335),
    .A2(net1002));
 sg13g2_a21oi_1 _3559_ (.A1(net1230),
    .A2(net1002),
    .Y(_0092_),
    .B1(_0779_));
 sg13g2_o21ai_1 _3560_ (.B1(net1234),
    .Y(_0780_),
    .A1(net342),
    .A2(net1002));
 sg13g2_a21oi_1 _3561_ (.A1(net1126),
    .A2(net1002),
    .Y(_0093_),
    .B1(_0780_));
 sg13g2_o21ai_1 _3562_ (.B1(net1234),
    .Y(_0781_),
    .A1(net346),
    .A2(_0778_));
 sg13g2_a21oi_1 _3563_ (.A1(net1127),
    .A2(net1002),
    .Y(_0094_),
    .B1(_0781_));
 sg13g2_o21ai_1 _3564_ (.B1(net1234),
    .Y(_0782_),
    .A1(net331),
    .A2(_0778_));
 sg13g2_a21oi_1 _3565_ (.A1(net1133),
    .A2(net1002),
    .Y(_0095_),
    .B1(_0782_));
 sg13g2_o21ai_1 _3566_ (.B1(net1234),
    .Y(_0783_),
    .A1(net313),
    .A2(net1002));
 sg13g2_a21oi_1 _3567_ (.A1(net1136),
    .A2(net1002),
    .Y(_0096_),
    .B1(_0783_));
 sg13g2_o21ai_1 _3568_ (.B1(net1238),
    .Y(_0784_),
    .A1(net1213),
    .A2(_0777_));
 sg13g2_a21oi_1 _3569_ (.A1(_1824_),
    .A2(_0777_),
    .Y(_0097_),
    .B1(_0784_));
 sg13g2_and2_1 _3570_ (.A(_0549_),
    .B(_0552_),
    .X(_0785_));
 sg13g2_nand2_1 _3571_ (.Y(_0786_),
    .A(_0549_),
    .B(_0552_));
 sg13g2_nor2_1 _3572_ (.A(net274),
    .B(_0786_),
    .Y(_0787_));
 sg13g2_nor2_1 _3573_ (.A(\spi_slave_0.bit_cnt[0] ),
    .B(_0785_),
    .Y(_0788_));
 sg13g2_nand2b_2 _3574_ (.Y(_0789_),
    .B(net1238),
    .A_N(net1));
 sg13g2_nor3_1 _3575_ (.A(_0787_),
    .B(_0788_),
    .C(_0789_),
    .Y(_0098_));
 sg13g2_a21oi_1 _3576_ (.A1(\spi_slave_0.bit_cnt[0] ),
    .A2(_0785_),
    .Y(_0790_),
    .B1(net292));
 sg13g2_and3_1 _3577_ (.X(_0791_),
    .A(net292),
    .B(\spi_slave_0.bit_cnt[0] ),
    .C(_0785_));
 sg13g2_nor3_1 _3578_ (.A(_0789_),
    .B(net293),
    .C(_0791_),
    .Y(_0099_));
 sg13g2_nor2_1 _3579_ (.A(net296),
    .B(_0791_),
    .Y(_0792_));
 sg13g2_nor2_1 _3580_ (.A(_0555_),
    .B(_0786_),
    .Y(_0793_));
 sg13g2_nor3_1 _3581_ (.A(_0789_),
    .B(net297),
    .C(_0793_),
    .Y(_0100_));
 sg13g2_o21ai_1 _3582_ (.B1(net1238),
    .Y(_0794_),
    .A1(miso),
    .A2(_0550_));
 sg13g2_a21oi_1 _3583_ (.A1(_1823_),
    .A2(_0550_),
    .Y(_0101_),
    .B1(_0794_));
 sg13g2_and2_2 _3584_ (.A(\charlie_0.memory[20][1] ),
    .B(\charlie_0.memory[20][0] ),
    .X(_0795_));
 sg13g2_and3_1 _3585_ (.X(_0796_),
    .A(_1834_),
    .B(\signal_generator_0.state_machine[1] ),
    .C(_0795_));
 sg13g2_a21oi_1 _3586_ (.A1(_1786_),
    .A2(\signal_generator_0.prev_clk_div ),
    .Y(_0797_),
    .B1(_2007_));
 sg13g2_o21ai_1 _3587_ (.B1(_0797_),
    .Y(_0798_),
    .A1(\charlie_0.memory[16][5] ),
    .A2(_2122_));
 sg13g2_nor2_1 _3588_ (.A(net1182),
    .B(net1183),
    .Y(_0799_));
 sg13g2_or2_1 _3589_ (.X(_0800_),
    .B(\signal_generator_0.index_reg[0] ),
    .A(\signal_generator_0.index_reg[1] ));
 sg13g2_nor3_2 _3590_ (.A(\signal_generator_0.index_reg[3] ),
    .B(net1180),
    .C(net1074),
    .Y(_0801_));
 sg13g2_and2_1 _3591_ (.A(_1820_),
    .B(_0801_),
    .X(_0802_));
 sg13g2_nand2_2 _3592_ (.Y(_0803_),
    .A(_1819_),
    .B(_0802_));
 sg13g2_nor2_1 _3593_ (.A(\signal_generator_0.index_reg[6] ),
    .B(_0803_),
    .Y(_0804_));
 sg13g2_nand2b_1 _3594_ (.Y(_0805_),
    .B(_0804_),
    .A_N(net953));
 sg13g2_nor2_1 _3595_ (.A(\signal_generator_0.index_reg[7] ),
    .B(\signal_generator_0.index_reg[6] ),
    .Y(_0806_));
 sg13g2_nor2b_2 _3596_ (.A(_0803_),
    .B_N(_0806_),
    .Y(_0807_));
 sg13g2_nor2b_2 _3597_ (.A(net953),
    .B_N(_0807_),
    .Y(_0808_));
 sg13g2_and2_2 _3598_ (.A(_0796_),
    .B(_0807_),
    .X(_0809_));
 sg13g2_nor2b_1 _3599_ (.A(net953),
    .B_N(_0809_),
    .Y(_0810_));
 sg13g2_nor2_2 _3600_ (.A(_1834_),
    .B(\signal_generator_0.state_machine[1] ),
    .Y(_0811_));
 sg13g2_nand2b_2 _3601_ (.Y(_0812_),
    .B(\signal_generator_0.state_machine[0] ),
    .A_N(\signal_generator_0.state_machine[1] ));
 sg13g2_xor2_1 _3602_ (.B(\signal_generator_0.state_machine[1] ),
    .A(\signal_generator_0.state_machine[0] ),
    .X(_0813_));
 sg13g2_a22oi_1 _3603_ (.Y(_0814_),
    .B1(_0808_),
    .B2(_0813_),
    .A2(_0564_),
    .A1(_1834_));
 sg13g2_nor2_1 _3604_ (.A(_0810_),
    .B(_0814_),
    .Y(_0815_));
 sg13g2_nor2_1 _3605_ (.A(net1226),
    .B(_0815_),
    .Y(_0102_));
 sg13g2_o21ai_1 _3606_ (.B1(net1257),
    .Y(_0816_),
    .A1(net338),
    .A2(_0808_));
 sg13g2_a21oi_1 _3607_ (.A1(_1834_),
    .A2(_0808_),
    .Y(_0103_),
    .B1(_0816_));
 sg13g2_a21oi_1 _3608_ (.A1(_0552_),
    .A2(_0556_),
    .Y(_0817_),
    .B1(net305));
 sg13g2_nor2_1 _3609_ (.A(_0789_),
    .B(net306),
    .Y(_0104_));
 sg13g2_nor2b_2 _3610_ (.A(net1163),
    .B_N(net1161),
    .Y(_0818_));
 sg13g2_nand2b_1 _3611_ (.Y(_0819_),
    .B(net1162),
    .A_N(net1164));
 sg13g2_nor2_1 _3612_ (.A(\charlie_0.memory[2][2] ),
    .B(net1068),
    .Y(_0820_));
 sg13g2_nor2b_2 _3613_ (.A(net1161),
    .B_N(net1163),
    .Y(_0821_));
 sg13g2_nand2b_2 _3614_ (.Y(_0822_),
    .B(net1163),
    .A_N(net1161));
 sg13g2_nor2_1 _3615_ (.A(\charlie_0.memory[2][1] ),
    .B(net1064),
    .Y(_0823_));
 sg13g2_nor2_2 _3616_ (.A(net1162),
    .B(net1163),
    .Y(_0824_));
 sg13g2_or2_1 _3617_ (.X(_0825_),
    .B(net1163),
    .A(net1161));
 sg13g2_and2_2 _3618_ (.A(net1162),
    .B(net1163),
    .X(_0826_));
 sg13g2_nand2_1 _3619_ (.Y(_0827_),
    .A(net1161),
    .B(net1163));
 sg13g2_nor2_1 _3620_ (.A(\charlie_0.memory[2][3] ),
    .B(net1054),
    .Y(_0828_));
 sg13g2_a22oi_1 _3621_ (.Y(_0829_),
    .B1(_0824_),
    .B2(_1814_),
    .A2(_0821_),
    .A1(_1813_));
 sg13g2_nor2_1 _3622_ (.A(\charlie_0.memory[3][1] ),
    .B(net1064),
    .Y(_0830_));
 sg13g2_nor2_1 _3623_ (.A(\charlie_0.memory[3][0] ),
    .B(net1059),
    .Y(_0831_));
 sg13g2_nor2_1 _3624_ (.A(\charlie_0.memory[3][3] ),
    .B(net1054),
    .Y(_0832_));
 sg13g2_nor2_1 _3625_ (.A(\charlie_0.memory[3][6] ),
    .B(net1068),
    .Y(_0833_));
 sg13g2_nor2_1 _3626_ (.A(\charlie_0.memory[3][5] ),
    .B(net1064),
    .Y(_0834_));
 sg13g2_nor2_1 _3627_ (.A(\charlie_0.memory[3][7] ),
    .B(net1054),
    .Y(_0835_));
 sg13g2_nor2_1 _3628_ (.A(\charlie_0.memory[0][4] ),
    .B(net1060),
    .Y(_0836_));
 sg13g2_nor2_1 _3629_ (.A(\charlie_0.memory[0][6] ),
    .B(net1068),
    .Y(_0837_));
 sg13g2_nor2_1 _3630_ (.A(\charlie_0.memory[0][5] ),
    .B(net1064),
    .Y(_0838_));
 sg13g2_o21ai_1 _3631_ (.B1(net1159),
    .Y(_0839_),
    .A1(\charlie_0.memory[0][7] ),
    .A2(net1054));
 sg13g2_nor4_1 _3632_ (.A(_0836_),
    .B(_0837_),
    .C(_0838_),
    .D(_0839_),
    .Y(_0840_));
 sg13g2_nor2_1 _3633_ (.A(\charlie_0.memory[0][0] ),
    .B(net1059),
    .Y(_0841_));
 sg13g2_nor2_1 _3634_ (.A(\charlie_0.memory[0][2] ),
    .B(net1068),
    .Y(_0842_));
 sg13g2_nor2_1 _3635_ (.A(\charlie_0.memory[0][1] ),
    .B(net1063),
    .Y(_0843_));
 sg13g2_o21ai_1 _3636_ (.B1(net1123),
    .Y(_0844_),
    .A1(\charlie_0.memory[0][3] ),
    .A2(net1053));
 sg13g2_nor4_1 _3637_ (.A(_0841_),
    .B(_0842_),
    .C(_0843_),
    .D(_0844_),
    .Y(_0845_));
 sg13g2_nor2_1 _3638_ (.A(\charlie_0.memory[1][2] ),
    .B(net1067),
    .Y(_0846_));
 sg13g2_nor2_1 _3639_ (.A(\charlie_0.memory[1][1] ),
    .B(net1063),
    .Y(_0847_));
 sg13g2_nor2_1 _3640_ (.A(\charlie_0.memory[1][3] ),
    .B(net1053),
    .Y(_0848_));
 sg13g2_nor2_1 _3641_ (.A(\charlie_0.memory[1][6] ),
    .B(net1067),
    .Y(_0849_));
 sg13g2_nor2_1 _3642_ (.A(\charlie_0.memory[1][7] ),
    .B(net1053),
    .Y(_0850_));
 sg13g2_nor2_1 _3643_ (.A(\charlie_0.memory[1][4] ),
    .B(net1059),
    .Y(_0851_));
 sg13g2_nor2_1 _3644_ (.A(\charlie_0.memory[6][2] ),
    .B(net1067),
    .Y(_0852_));
 sg13g2_nor2_1 _3645_ (.A(\charlie_0.memory[6][3] ),
    .B(net1053),
    .Y(_0853_));
 sg13g2_nor2_1 _3646_ (.A(\charlie_0.memory[6][0] ),
    .B(net1058),
    .Y(_0854_));
 sg13g2_nor2_1 _3647_ (.A(\charlie_0.memory[6][6] ),
    .B(net1067),
    .Y(_0855_));
 sg13g2_nor2_1 _3648_ (.A(\charlie_0.memory[6][5] ),
    .B(net1063),
    .Y(_0856_));
 sg13g2_nor2_1 _3649_ (.A(\charlie_0.memory[6][4] ),
    .B(net1058),
    .Y(_0857_));
 sg13g2_nor2_1 _3650_ (.A(\charlie_0.memory[7][1] ),
    .B(net1064),
    .Y(_0858_));
 sg13g2_nor2_1 _3651_ (.A(\charlie_0.memory[7][3] ),
    .B(net1054),
    .Y(_0859_));
 sg13g2_nor2_1 _3652_ (.A(\charlie_0.memory[7][2] ),
    .B(net1068),
    .Y(_0860_));
 sg13g2_nor3_1 _3653_ (.A(net1161),
    .B(net1164),
    .C(\charlie_0.memory[7][4] ),
    .Y(_0861_));
 sg13g2_o21ai_1 _3654_ (.B1(net1160),
    .Y(_0862_),
    .A1(\charlie_0.memory[4][6] ),
    .A2(net1067));
 sg13g2_nor2_1 _3655_ (.A(\charlie_0.memory[4][7] ),
    .B(net1053),
    .Y(_0863_));
 sg13g2_nor2_1 _3656_ (.A(\charlie_0.memory[4][5] ),
    .B(net1063),
    .Y(_0864_));
 sg13g2_nor2_1 _3657_ (.A(\charlie_0.memory[4][4] ),
    .B(net1058),
    .Y(_0865_));
 sg13g2_or4_1 _3658_ (.A(_0862_),
    .B(_0863_),
    .C(_0864_),
    .D(_0865_),
    .X(_0866_));
 sg13g2_nor2_1 _3659_ (.A(\charlie_0.memory[4][3] ),
    .B(net1053),
    .Y(_0867_));
 sg13g2_nor2_1 _3660_ (.A(\charlie_0.memory[4][0] ),
    .B(net1058),
    .Y(_0868_));
 sg13g2_nor2_1 _3661_ (.A(\charlie_0.memory[4][1] ),
    .B(net1063),
    .Y(_0869_));
 sg13g2_o21ai_1 _3662_ (.B1(net1122),
    .Y(_0870_),
    .A1(\charlie_0.memory[4][2] ),
    .A2(net1067));
 sg13g2_or4_1 _3663_ (.A(_0867_),
    .B(_0868_),
    .C(_0869_),
    .D(_0870_),
    .X(_0871_));
 sg13g2_nor2_1 _3664_ (.A(\charlie_0.memory[5][3] ),
    .B(net1054),
    .Y(_0872_));
 sg13g2_nor2_1 _3665_ (.A(\charlie_0.memory[5][1] ),
    .B(net1064),
    .Y(_0873_));
 sg13g2_nor2_1 _3666_ (.A(\charlie_0.memory[5][2] ),
    .B(net1068),
    .Y(_0874_));
 sg13g2_nor2_1 _3667_ (.A(\charlie_0.memory[5][6] ),
    .B(net1067),
    .Y(_0875_));
 sg13g2_nor2_1 _3668_ (.A(\charlie_0.memory[5][7] ),
    .B(net1053),
    .Y(_0876_));
 sg13g2_nor2_1 _3669_ (.A(\charlie_0.memory[5][5] ),
    .B(net1063),
    .Y(_0877_));
 sg13g2_nor2_1 _3670_ (.A(\charlie_0.memory[13][2] ),
    .B(net1066),
    .Y(_0878_));
 sg13g2_nor2_1 _3671_ (.A(\charlie_0.memory[13][3] ),
    .B(net1052),
    .Y(_0879_));
 sg13g2_nor2_1 _3672_ (.A(\charlie_0.memory[13][0] ),
    .B(net1056),
    .Y(_0880_));
 sg13g2_nor2_1 _3673_ (.A(\charlie_0.memory[13][4] ),
    .B(net1057),
    .Y(_0881_));
 sg13g2_nor2_1 _3674_ (.A(\charlie_0.memory[13][5] ),
    .B(net1061),
    .Y(_0882_));
 sg13g2_nor2_1 _3675_ (.A(\charlie_0.memory[13][6] ),
    .B(net1065),
    .Y(_0883_));
 sg13g2_nor2_1 _3676_ (.A(\charlie_0.memory[12][1] ),
    .B(net1062),
    .Y(_0884_));
 sg13g2_nor2_1 _3677_ (.A(\charlie_0.memory[12][2] ),
    .B(net1065),
    .Y(_0885_));
 sg13g2_nor2_1 _3678_ (.A(\charlie_0.memory[12][0] ),
    .B(net1060),
    .Y(_0886_));
 sg13g2_nor2_1 _3679_ (.A(\charlie_0.memory[12][6] ),
    .B(net1066),
    .Y(_0887_));
 sg13g2_nor2_1 _3680_ (.A(\charlie_0.memory[12][4] ),
    .B(net1057),
    .Y(_0888_));
 sg13g2_nor2_1 _3681_ (.A(\charlie_0.memory[12][7] ),
    .B(net1052),
    .Y(_0889_));
 sg13g2_nor2_1 _3682_ (.A(\charlie_0.memory[14][1] ),
    .B(net1061),
    .Y(_0890_));
 sg13g2_nor2_1 _3683_ (.A(\charlie_0.memory[14][0] ),
    .B(net1056),
    .Y(_0891_));
 sg13g2_nor2_1 _3684_ (.A(\charlie_0.memory[14][3] ),
    .B(net1051),
    .Y(_0892_));
 sg13g2_o21ai_1 _3685_ (.B1(net1121),
    .Y(_0893_),
    .A1(\charlie_0.memory[14][2] ),
    .A2(net1065));
 sg13g2_or4_1 _3686_ (.A(_0890_),
    .B(_0891_),
    .C(_0892_),
    .D(_0893_),
    .X(_0894_));
 sg13g2_a22oi_1 _3687_ (.Y(_0895_),
    .B1(_0826_),
    .B2(_1792_),
    .A2(_0824_),
    .A1(_1795_));
 sg13g2_a221oi_1 _3688_ (.B2(_1794_),
    .C1(net1121),
    .B1(_0821_),
    .A1(_1793_),
    .Y(_0896_),
    .A2(_0818_));
 sg13g2_nor2_1 _3689_ (.A(\charlie_0.memory[15][1] ),
    .B(net1062),
    .Y(_0897_));
 sg13g2_nor2_1 _3690_ (.A(\charlie_0.memory[15][0] ),
    .B(net1057),
    .Y(_0898_));
 sg13g2_nor2_1 _3691_ (.A(\charlie_0.memory[15][3] ),
    .B(net1052),
    .Y(_0899_));
 sg13g2_nor2_1 _3692_ (.A(\charlie_0.memory[15][6] ),
    .B(net1066),
    .Y(_0900_));
 sg13g2_nor2_1 _3693_ (.A(\charlie_0.memory[15][5] ),
    .B(net1062),
    .Y(_0901_));
 sg13g2_nor2_1 _3694_ (.A(\charlie_0.memory[15][7] ),
    .B(net1052),
    .Y(_0902_));
 sg13g2_nor2_1 _3695_ (.A(\charlie_0.memory[9][2] ),
    .B(net1065),
    .Y(_0903_));
 sg13g2_nor2_1 _3696_ (.A(\charlie_0.memory[9][1] ),
    .B(net1061),
    .Y(_0904_));
 sg13g2_nor2_1 _3697_ (.A(\charlie_0.memory[9][3] ),
    .B(net1051),
    .Y(_0905_));
 sg13g2_nor2_1 _3698_ (.A(\charlie_0.memory[9][7] ),
    .B(net1051),
    .Y(_0906_));
 sg13g2_nor2_1 _3699_ (.A(\charlie_0.memory[9][4] ),
    .B(net1056),
    .Y(_0907_));
 sg13g2_nor2_1 _3700_ (.A(\charlie_0.memory[9][6] ),
    .B(net1065),
    .Y(_0908_));
 sg13g2_nor2_1 _3701_ (.A(\charlie_0.memory[8][3] ),
    .B(net1051),
    .Y(_0909_));
 sg13g2_nor2_1 _3702_ (.A(\charlie_0.memory[8][0] ),
    .B(net1057),
    .Y(_0910_));
 sg13g2_nor2_1 _3703_ (.A(\charlie_0.memory[8][1] ),
    .B(net1061),
    .Y(_0911_));
 sg13g2_nor2_1 _3704_ (.A(\charlie_0.memory[8][7] ),
    .B(net1051),
    .Y(_0912_));
 sg13g2_nor2_1 _3705_ (.A(\charlie_0.memory[8][4] ),
    .B(net1057),
    .Y(_0913_));
 sg13g2_nor2_1 _3706_ (.A(\charlie_0.memory[8][6] ),
    .B(net1069),
    .Y(_0914_));
 sg13g2_a22oi_1 _3707_ (.Y(_0915_),
    .B1(_0824_),
    .B2(_1802_),
    .A2(_0818_),
    .A1(_1800_));
 sg13g2_a221oi_1 _3708_ (.B2(_1799_),
    .C1(net1158),
    .B1(_0826_),
    .A1(_1801_),
    .Y(_0916_),
    .A2(_0821_));
 sg13g2_a21oi_1 _3709_ (.A1(_1796_),
    .A2(_0826_),
    .Y(_0917_),
    .B1(net1121));
 sg13g2_nor2_1 _3710_ (.A(\charlie_0.memory[10][4] ),
    .B(net1056),
    .Y(_0918_));
 sg13g2_a221oi_1 _3711_ (.B2(_1798_),
    .C1(_0918_),
    .B1(_0821_),
    .A1(_1797_),
    .Y(_0919_),
    .A2(_0818_));
 sg13g2_a22oi_1 _3712_ (.Y(_0920_),
    .B1(_0917_),
    .B2(_0919_),
    .A2(_0916_),
    .A1(_0915_));
 sg13g2_nor2_1 _3713_ (.A(\charlie_0.memory[11][1] ),
    .B(net1061),
    .Y(_0921_));
 sg13g2_nor2_1 _3714_ (.A(\charlie_0.memory[11][0] ),
    .B(net1056),
    .Y(_0922_));
 sg13g2_nor2_1 _3715_ (.A(\charlie_0.memory[11][3] ),
    .B(net1051),
    .Y(_0923_));
 sg13g2_nor2_1 _3716_ (.A(\charlie_0.memory[11][4] ),
    .B(net1056),
    .Y(_0924_));
 sg13g2_nor2_1 _3717_ (.A(\charlie_0.memory[11][6] ),
    .B(net1065),
    .Y(_0925_));
 sg13g2_nor2_1 _3718_ (.A(\charlie_0.memory[11][5] ),
    .B(net1061),
    .Y(_0926_));
 sg13g2_o21ai_1 _3719_ (.B1(net1158),
    .Y(_0927_),
    .A1(\charlie_0.memory[8][5] ),
    .A2(net1061));
 sg13g2_nor4_1 _3720_ (.A(_0912_),
    .B(_0913_),
    .C(_0914_),
    .D(_0927_),
    .Y(_0928_));
 sg13g2_o21ai_1 _3721_ (.B1(net1121),
    .Y(_0929_),
    .A1(\charlie_0.memory[8][2] ),
    .A2(net1065));
 sg13g2_nor4_1 _3722_ (.A(_0909_),
    .B(_0910_),
    .C(_0911_),
    .D(_0929_),
    .Y(_0930_));
 sg13g2_nor2_1 _3723_ (.A(_0928_),
    .B(_0930_),
    .Y(_0931_));
 sg13g2_o21ai_1 _3724_ (.B1(net1121),
    .Y(_0932_),
    .A1(\charlie_0.memory[9][0] ),
    .A2(net1056));
 sg13g2_nor4_1 _3725_ (.A(_0903_),
    .B(_0904_),
    .C(_0905_),
    .D(_0932_),
    .Y(_0933_));
 sg13g2_o21ai_1 _3726_ (.B1(net1158),
    .Y(_0934_),
    .A1(\charlie_0.memory[9][5] ),
    .A2(net1061));
 sg13g2_nor4_1 _3727_ (.A(_0906_),
    .B(_0907_),
    .C(_0908_),
    .D(_0934_),
    .Y(_0935_));
 sg13g2_nor2_1 _3728_ (.A(_0933_),
    .B(_0935_),
    .Y(_0936_));
 sg13g2_o21ai_1 _3729_ (.B1(net1158),
    .Y(_0937_),
    .A1(\charlie_0.memory[11][7] ),
    .A2(net1051));
 sg13g2_nor4_1 _3730_ (.A(_0924_),
    .B(_0925_),
    .C(_0926_),
    .D(_0937_),
    .Y(_0938_));
 sg13g2_o21ai_1 _3731_ (.B1(net1121),
    .Y(_0939_),
    .A1(\charlie_0.memory[11][2] ),
    .A2(net1065));
 sg13g2_nor4_1 _3732_ (.A(_0921_),
    .B(_0922_),
    .C(_0923_),
    .D(_0939_),
    .Y(_0940_));
 sg13g2_nor2_1 _3733_ (.A(_0938_),
    .B(_0940_),
    .Y(_0941_));
 sg13g2_mux4_1 _3734_ (.S0(_1780_),
    .A0(_0920_),
    .A1(_0931_),
    .A2(_0941_),
    .A3(_0936_),
    .S1(net1156),
    .X(_0942_));
 sg13g2_o21ai_1 _3735_ (.B1(net1160),
    .Y(_0943_),
    .A1(\charlie_0.memory[12][5] ),
    .A2(net1062));
 sg13g2_nor4_1 _3736_ (.A(_0887_),
    .B(_0888_),
    .C(_0889_),
    .D(_0943_),
    .Y(_0944_));
 sg13g2_o21ai_1 _3737_ (.B1(net1121),
    .Y(_0945_),
    .A1(\charlie_0.memory[12][3] ),
    .A2(net1055));
 sg13g2_nor4_1 _3738_ (.A(_0884_),
    .B(_0885_),
    .C(_0886_),
    .D(_0945_),
    .Y(_0946_));
 sg13g2_nor3_1 _3739_ (.A(net1156),
    .B(_0944_),
    .C(_0946_),
    .Y(_0947_));
 sg13g2_o21ai_1 _3740_ (.B1(net1158),
    .Y(_0948_),
    .A1(\charlie_0.memory[13][7] ),
    .A2(net1051));
 sg13g2_nor4_1 _3741_ (.A(_0881_),
    .B(_0882_),
    .C(_0883_),
    .D(_0948_),
    .Y(_0949_));
 sg13g2_o21ai_1 _3742_ (.B1(net1121),
    .Y(_0950_),
    .A1(\charlie_0.memory[13][1] ),
    .A2(net1062));
 sg13g2_nor4_1 _3743_ (.A(_0878_),
    .B(_0879_),
    .C(_0880_),
    .D(_0950_),
    .Y(_0951_));
 sg13g2_nor3_1 _3744_ (.A(_1781_),
    .B(_0949_),
    .C(_0951_),
    .Y(_0952_));
 sg13g2_or3_1 _3745_ (.A(\charlie_0.memory[17][4] ),
    .B(_0947_),
    .C(_0952_),
    .X(_0953_));
 sg13g2_o21ai_1 _3746_ (.B1(net1158),
    .Y(_0954_),
    .A1(\charlie_0.memory[15][4] ),
    .A2(net1056));
 sg13g2_nor4_1 _3747_ (.A(_0900_),
    .B(_0901_),
    .C(_0902_),
    .D(_0954_),
    .Y(_0955_));
 sg13g2_o21ai_1 _3748_ (.B1(net1124),
    .Y(_0956_),
    .A1(\charlie_0.memory[15][2] ),
    .A2(net1066));
 sg13g2_nor4_1 _3749_ (.A(_0897_),
    .B(_0898_),
    .C(_0899_),
    .D(_0956_),
    .Y(_0957_));
 sg13g2_or3_1 _3750_ (.A(_1781_),
    .B(_0955_),
    .C(_0957_),
    .X(_0958_));
 sg13g2_a21oi_1 _3751_ (.A1(_0895_),
    .A2(_0896_),
    .Y(_0959_),
    .B1(net1156));
 sg13g2_a21oi_1 _3752_ (.A1(_0894_),
    .A2(_0959_),
    .Y(_0960_),
    .B1(_1780_));
 sg13g2_a21oi_1 _3753_ (.A1(_0958_),
    .A2(_0960_),
    .Y(_0961_),
    .B1(_1779_));
 sg13g2_a221oi_1 _3754_ (.B2(_0961_),
    .C1(_1778_),
    .B1(_0953_),
    .A1(_1779_),
    .Y(_0962_),
    .A2(_0942_));
 sg13g2_o21ai_1 _3755_ (.B1(net1159),
    .Y(_0963_),
    .A1(\charlie_0.memory[6][7] ),
    .A2(net1053));
 sg13g2_nor4_1 _3756_ (.A(_0855_),
    .B(_0856_),
    .C(_0857_),
    .D(_0963_),
    .Y(_0964_));
 sg13g2_o21ai_1 _3757_ (.B1(net1122),
    .Y(_0965_),
    .A1(\charlie_0.memory[6][1] ),
    .A2(net1063));
 sg13g2_nor4_1 _3758_ (.A(_0852_),
    .B(_0853_),
    .C(_0854_),
    .D(_0965_),
    .Y(_0966_));
 sg13g2_or3_1 _3759_ (.A(net1157),
    .B(_0964_),
    .C(_0966_),
    .X(_0967_));
 sg13g2_o21ai_1 _3760_ (.B1(net1122),
    .Y(_0968_),
    .A1(\charlie_0.memory[7][0] ),
    .A2(net1058));
 sg13g2_or4_1 _3761_ (.A(_0858_),
    .B(_0859_),
    .C(_0860_),
    .D(_0968_),
    .X(_0969_));
 sg13g2_a21oi_1 _3762_ (.A1(_1804_),
    .A2(_0818_),
    .Y(_0970_),
    .B1(net1122));
 sg13g2_a221oi_1 _3763_ (.B2(_1803_),
    .C1(_0861_),
    .B1(_0826_),
    .A1(_1805_),
    .Y(_0971_),
    .A2(_0821_));
 sg13g2_a21oi_1 _3764_ (.A1(_0970_),
    .A2(_0971_),
    .Y(_0972_),
    .B1(_1781_));
 sg13g2_a21oi_1 _3765_ (.A1(_0969_),
    .A2(_0972_),
    .Y(_0973_),
    .B1(_1780_));
 sg13g2_nand3_1 _3766_ (.B(_0866_),
    .C(_0871_),
    .A(_1781_),
    .Y(_0974_));
 sg13g2_o21ai_1 _3767_ (.B1(net1122),
    .Y(_0975_),
    .A1(\charlie_0.memory[5][0] ),
    .A2(net1058));
 sg13g2_nor4_1 _3768_ (.A(_0872_),
    .B(_0873_),
    .C(_0874_),
    .D(_0975_),
    .Y(_0976_));
 sg13g2_o21ai_1 _3769_ (.B1(net1159),
    .Y(_0977_),
    .A1(\charlie_0.memory[5][4] ),
    .A2(net1058));
 sg13g2_nor4_1 _3770_ (.A(_0875_),
    .B(_0876_),
    .C(_0877_),
    .D(_0977_),
    .Y(_0978_));
 sg13g2_or3_1 _3771_ (.A(_1781_),
    .B(_0976_),
    .C(_0978_),
    .X(_0979_));
 sg13g2_nand3_1 _3772_ (.B(_0974_),
    .C(_0979_),
    .A(_1780_),
    .Y(_0980_));
 sg13g2_a21oi_1 _3773_ (.A1(_0967_),
    .A2(_0973_),
    .Y(_0981_),
    .B1(_1779_));
 sg13g2_o21ai_1 _3774_ (.B1(net1123),
    .Y(_0982_),
    .A1(\charlie_0.memory[1][0] ),
    .A2(net1058));
 sg13g2_nor4_1 _3775_ (.A(_0846_),
    .B(_0847_),
    .C(_0848_),
    .D(_0982_),
    .Y(_0983_));
 sg13g2_o21ai_1 _3776_ (.B1(net1159),
    .Y(_0984_),
    .A1(\charlie_0.memory[1][5] ),
    .A2(net1063));
 sg13g2_nor4_1 _3777_ (.A(_0849_),
    .B(_0850_),
    .C(_0851_),
    .D(_0984_),
    .Y(_0985_));
 sg13g2_nor3_1 _3778_ (.A(_1781_),
    .B(_0983_),
    .C(_0985_),
    .Y(_0986_));
 sg13g2_nor3_1 _3779_ (.A(net1157),
    .B(_0840_),
    .C(_0845_),
    .Y(_0987_));
 sg13g2_or3_1 _3780_ (.A(\charlie_0.memory[17][4] ),
    .B(_0986_),
    .C(_0987_),
    .X(_0988_));
 sg13g2_o21ai_1 _3781_ (.B1(net1159),
    .Y(_0989_),
    .A1(\charlie_0.memory[3][4] ),
    .A2(net1059));
 sg13g2_nor4_1 _3782_ (.A(_0833_),
    .B(_0834_),
    .C(_0835_),
    .D(_0989_),
    .Y(_0990_));
 sg13g2_o21ai_1 _3783_ (.B1(net1123),
    .Y(_0991_),
    .A1(\charlie_0.memory[3][2] ),
    .A2(net1067));
 sg13g2_nor4_1 _3784_ (.A(_0830_),
    .B(_0831_),
    .C(_0832_),
    .D(_0991_),
    .Y(_0992_));
 sg13g2_or3_1 _3785_ (.A(_1781_),
    .B(_0990_),
    .C(_0992_),
    .X(_0993_));
 sg13g2_o21ai_1 _3786_ (.B1(net1122),
    .Y(_0994_),
    .A1(\charlie_0.memory[2][0] ),
    .A2(net1059));
 sg13g2_or4_1 _3787_ (.A(_0820_),
    .B(_0823_),
    .C(_0828_),
    .D(_0994_),
    .X(_0995_));
 sg13g2_a221oi_1 _3788_ (.B2(_1811_),
    .C1(net1122),
    .B1(_0826_),
    .A1(_1812_),
    .Y(_0996_),
    .A2(_0818_));
 sg13g2_a21oi_1 _3789_ (.A1(_0829_),
    .A2(_0996_),
    .Y(_0997_),
    .B1(net1157));
 sg13g2_a21oi_1 _3790_ (.A1(_0995_),
    .A2(_0997_),
    .Y(_0998_),
    .B1(_1780_));
 sg13g2_a21oi_1 _3791_ (.A1(_0993_),
    .A2(_0998_),
    .Y(_0999_),
    .B1(\charlie_0.memory[17][5] ));
 sg13g2_a221oi_1 _3792_ (.B2(_0999_),
    .C1(\charlie_0.memory[17][6] ),
    .B1(_0988_),
    .A1(_0980_),
    .Y(_1000_),
    .A2(_0981_));
 sg13g2_or2_1 _3793_ (.X(_1001_),
    .B(_1000_),
    .A(_0962_));
 sg13g2_o21ai_1 _3794_ (.B1(_0565_),
    .Y(_1002_),
    .A1(_0962_),
    .A2(_1000_));
 sg13g2_nand2_1 _3795_ (.Y(_1003_),
    .A(net383),
    .B(_0564_));
 sg13g2_nand2_1 _3796_ (.Y(_1004_),
    .A(_1002_),
    .B(_1003_));
 sg13g2_a21oi_1 _3797_ (.A1(_1002_),
    .A2(_1003_),
    .Y(_1005_),
    .B1(_0811_));
 sg13g2_nor2_1 _3798_ (.A(\charlie_0.memory[0][0] ),
    .B(net1074),
    .Y(_1006_));
 sg13g2_nor2b_1 _3799_ (.A(\signal_generator_0.index_reg[0] ),
    .B_N(net1182),
    .Y(_1007_));
 sg13g2_nand2b_1 _3800_ (.Y(_1008_),
    .B(\signal_generator_0.index_reg[1] ),
    .A_N(net1183));
 sg13g2_nor2_1 _3801_ (.A(\charlie_0.memory[0][2] ),
    .B(net1047),
    .Y(_1009_));
 sg13g2_nor2b_1 _3802_ (.A(net1182),
    .B_N(net1183),
    .Y(_1010_));
 sg13g2_nand2b_1 _3803_ (.Y(_1011_),
    .B(net1183),
    .A_N(net1182));
 sg13g2_and2_1 _3804_ (.A(net1182),
    .B(net1183),
    .X(_1012_));
 sg13g2_nand2_1 _3805_ (.Y(_1013_),
    .A(net1182),
    .B(net1183));
 sg13g2_nor2_1 _3806_ (.A(\charlie_0.memory[0][3] ),
    .B(net1033),
    .Y(_1014_));
 sg13g2_o21ai_1 _3807_ (.B1(net1117),
    .Y(_1015_),
    .A1(\charlie_0.memory[0][1] ),
    .A2(net1039));
 sg13g2_nor4_1 _3808_ (.A(_1006_),
    .B(_1009_),
    .C(_1014_),
    .D(_1015_),
    .Y(_1016_));
 sg13g2_o21ai_1 _3809_ (.B1(net1179),
    .Y(_1017_),
    .A1(\charlie_0.memory[0][4] ),
    .A2(net1074));
 sg13g2_nor2_1 _3810_ (.A(\charlie_0.memory[0][6] ),
    .B(net1047),
    .Y(_1018_));
 sg13g2_nor2_1 _3811_ (.A(\charlie_0.memory[0][5] ),
    .B(net1040),
    .Y(_1019_));
 sg13g2_nor2_1 _3812_ (.A(\charlie_0.memory[0][7] ),
    .B(net1033),
    .Y(_1020_));
 sg13g2_nor4_1 _3813_ (.A(_1017_),
    .B(_1018_),
    .C(_1019_),
    .D(_1020_),
    .Y(_1021_));
 sg13g2_nor2_1 _3814_ (.A(_1016_),
    .B(_1021_),
    .Y(_1022_));
 sg13g2_nor2_1 _3815_ (.A(\charlie_0.memory[1][3] ),
    .B(net1034),
    .Y(_1023_));
 sg13g2_nor2_1 _3816_ (.A(\charlie_0.memory[1][2] ),
    .B(net1047),
    .Y(_1024_));
 sg13g2_nor2_1 _3817_ (.A(\charlie_0.memory[1][0] ),
    .B(net1075),
    .Y(_1025_));
 sg13g2_o21ai_1 _3818_ (.B1(net1116),
    .Y(_1026_),
    .A1(\charlie_0.memory[1][1] ),
    .A2(net1040));
 sg13g2_nor4_1 _3819_ (.A(_1023_),
    .B(_1024_),
    .C(_1025_),
    .D(_1026_),
    .Y(_1027_));
 sg13g2_o21ai_1 _3820_ (.B1(net1179),
    .Y(_1028_),
    .A1(\charlie_0.memory[1][7] ),
    .A2(net1032));
 sg13g2_nor2_1 _3821_ (.A(\charlie_0.memory[1][6] ),
    .B(net1046),
    .Y(_1029_));
 sg13g2_nor2_1 _3822_ (.A(\charlie_0.memory[1][5] ),
    .B(net1039),
    .Y(_1030_));
 sg13g2_nor2_1 _3823_ (.A(\charlie_0.memory[1][4] ),
    .B(net1075),
    .Y(_1031_));
 sg13g2_nor4_1 _3824_ (.A(_1028_),
    .B(_1029_),
    .C(_1030_),
    .D(_1031_),
    .Y(_1032_));
 sg13g2_nor2_1 _3825_ (.A(_1027_),
    .B(_1032_),
    .Y(_1033_));
 sg13g2_nor2_1 _3826_ (.A(\charlie_0.memory[3][0] ),
    .B(net1074),
    .Y(_1034_));
 sg13g2_nor2_1 _3827_ (.A(\charlie_0.memory[3][2] ),
    .B(net1047),
    .Y(_1035_));
 sg13g2_nor2_1 _3828_ (.A(\charlie_0.memory[3][3] ),
    .B(net1033),
    .Y(_1036_));
 sg13g2_o21ai_1 _3829_ (.B1(net1117),
    .Y(_1037_),
    .A1(\charlie_0.memory[3][1] ),
    .A2(net1039));
 sg13g2_nor4_1 _3830_ (.A(_1034_),
    .B(_1035_),
    .C(_1036_),
    .D(_1037_),
    .Y(_1038_));
 sg13g2_nor2_1 _3831_ (.A(\charlie_0.memory[3][6] ),
    .B(net1047),
    .Y(_1039_));
 sg13g2_nor2_1 _3832_ (.A(\charlie_0.memory[3][5] ),
    .B(net1039),
    .Y(_1040_));
 sg13g2_nor2_1 _3833_ (.A(\charlie_0.memory[3][7] ),
    .B(net1033),
    .Y(_1041_));
 sg13g2_o21ai_1 _3834_ (.B1(net1179),
    .Y(_1042_),
    .A1(\charlie_0.memory[3][4] ),
    .A2(net1074));
 sg13g2_nor4_1 _3835_ (.A(_1039_),
    .B(_1040_),
    .C(_1041_),
    .D(_1042_),
    .Y(_1043_));
 sg13g2_nor2_1 _3836_ (.A(_1038_),
    .B(_1043_),
    .Y(_1044_));
 sg13g2_nand2_2 _3837_ (.Y(_1045_),
    .A(net1176),
    .B(net1118));
 sg13g2_nor2_1 _3838_ (.A(\charlie_0.memory[2][6] ),
    .B(net1047),
    .Y(_1046_));
 sg13g2_a21oi_1 _3839_ (.A1(_1813_),
    .A2(net1042),
    .Y(_1047_),
    .B1(net1116));
 sg13g2_a221oi_1 _3840_ (.B2(_1811_),
    .C1(_1046_),
    .B1(net1035),
    .A1(_1814_),
    .Y(_1048_),
    .A2(net1077));
 sg13g2_nor2_1 _3841_ (.A(\charlie_0.memory[2][2] ),
    .B(net1047),
    .Y(_1049_));
 sg13g2_nor2_1 _3842_ (.A(\charlie_0.memory[2][0] ),
    .B(net1074),
    .Y(_1050_));
 sg13g2_nor2_1 _3843_ (.A(\charlie_0.memory[2][3] ),
    .B(net1033),
    .Y(_1051_));
 sg13g2_o21ai_1 _3844_ (.B1(net1117),
    .Y(_1052_),
    .A1(\charlie_0.memory[2][1] ),
    .A2(net1039));
 sg13g2_nor4_1 _3845_ (.A(_1049_),
    .B(_1050_),
    .C(_1051_),
    .D(_1052_),
    .Y(_1053_));
 sg13g2_a21oi_1 _3846_ (.A1(_1047_),
    .A2(_1048_),
    .Y(_1054_),
    .B1(_1053_));
 sg13g2_mux4_1 _3847_ (.S0(net1177),
    .A0(_1022_),
    .A1(_1033_),
    .A2(_1054_),
    .A3(_1044_),
    .S1(net1176),
    .X(_1055_));
 sg13g2_nor2_1 _3848_ (.A(\signal_generator_0.index_reg[5] ),
    .B(_1055_),
    .Y(_1056_));
 sg13g2_o21ai_1 _3849_ (.B1(_1821_),
    .Y(_1057_),
    .A1(\charlie_0.memory[4][1] ),
    .A2(net1038));
 sg13g2_nor2_1 _3850_ (.A(\charlie_0.memory[4][2] ),
    .B(net1048),
    .Y(_1058_));
 sg13g2_nor2_1 _3851_ (.A(\charlie_0.memory[4][3] ),
    .B(net1032),
    .Y(_1059_));
 sg13g2_nor2_1 _3852_ (.A(\charlie_0.memory[4][0] ),
    .B(net1073),
    .Y(_1060_));
 sg13g2_nor4_1 _3853_ (.A(_1057_),
    .B(_1058_),
    .C(_1059_),
    .D(_1060_),
    .Y(_1061_));
 sg13g2_nor2_1 _3854_ (.A(\charlie_0.memory[5][1] ),
    .B(net1038),
    .Y(_1062_));
 sg13g2_nor2_1 _3855_ (.A(\charlie_0.memory[5][2] ),
    .B(net1046),
    .Y(_1063_));
 sg13g2_nor2_1 _3856_ (.A(\charlie_0.memory[5][3] ),
    .B(net1032),
    .Y(_1064_));
 sg13g2_o21ai_1 _3857_ (.B1(net1177),
    .Y(_1065_),
    .A1(\charlie_0.memory[5][0] ),
    .A2(net1073));
 sg13g2_nor4_1 _3858_ (.A(_1062_),
    .B(_1063_),
    .C(_1064_),
    .D(_1065_),
    .Y(_1066_));
 sg13g2_or3_1 _3859_ (.A(net1179),
    .B(_1061_),
    .C(_1066_),
    .X(_1067_));
 sg13g2_o21ai_1 _3860_ (.B1(net1177),
    .Y(_1068_),
    .A1(\charlie_0.memory[5][4] ),
    .A2(net1073));
 sg13g2_nor2_1 _3861_ (.A(\charlie_0.memory[5][6] ),
    .B(net1046),
    .Y(_1069_));
 sg13g2_nor2_1 _3862_ (.A(\charlie_0.memory[5][7] ),
    .B(net1034),
    .Y(_1070_));
 sg13g2_nor2_1 _3863_ (.A(\charlie_0.memory[5][5] ),
    .B(net1038),
    .Y(_1071_));
 sg13g2_nor4_1 _3864_ (.A(_1068_),
    .B(_1069_),
    .C(_1070_),
    .D(_1071_),
    .Y(_1072_));
 sg13g2_nor2_1 _3865_ (.A(\charlie_0.memory[4][7] ),
    .B(net1032),
    .Y(_1073_));
 sg13g2_nor2_1 _3866_ (.A(\charlie_0.memory[4][4] ),
    .B(net1073),
    .Y(_1074_));
 sg13g2_nor2_1 _3867_ (.A(\charlie_0.memory[4][5] ),
    .B(net1038),
    .Y(_1075_));
 sg13g2_o21ai_1 _3868_ (.B1(_1821_),
    .Y(_1076_),
    .A1(\charlie_0.memory[4][6] ),
    .A2(net1046));
 sg13g2_nor4_1 _3869_ (.A(_1073_),
    .B(_1074_),
    .C(_1075_),
    .D(_1076_),
    .Y(_1077_));
 sg13g2_or3_1 _3870_ (.A(net1116),
    .B(_1072_),
    .C(_1077_),
    .X(_1078_));
 sg13g2_a21oi_2 _3871_ (.B1(net1176),
    .Y(_1079_),
    .A2(_1078_),
    .A1(_1067_));
 sg13g2_o21ai_1 _3872_ (.B1(net1116),
    .Y(_1080_),
    .A1(\charlie_0.memory[7][3] ),
    .A2(net1032));
 sg13g2_nor2_1 _3873_ (.A(\charlie_0.memory[7][2] ),
    .B(net1046),
    .Y(_1081_));
 sg13g2_nor2_1 _3874_ (.A(\charlie_0.memory[7][0] ),
    .B(net1073),
    .Y(_1082_));
 sg13g2_nor2_1 _3875_ (.A(\charlie_0.memory[7][1] ),
    .B(net1038),
    .Y(_1083_));
 sg13g2_nor4_1 _3876_ (.A(_1080_),
    .B(_1081_),
    .C(_1082_),
    .D(_1083_),
    .Y(_1084_));
 sg13g2_nor2_1 _3877_ (.A(\charlie_0.memory[7][6] ),
    .B(net1046),
    .Y(_1085_));
 sg13g2_nor2_1 _3878_ (.A(\charlie_0.memory[7][7] ),
    .B(net1032),
    .Y(_1086_));
 sg13g2_nor2_1 _3879_ (.A(\charlie_0.memory[7][5] ),
    .B(net1038),
    .Y(_1087_));
 sg13g2_o21ai_1 _3880_ (.B1(net1179),
    .Y(_1088_),
    .A1(\charlie_0.memory[7][4] ),
    .A2(net1073));
 sg13g2_nor4_1 _3881_ (.A(_1085_),
    .B(_1086_),
    .C(_1087_),
    .D(_1088_),
    .Y(_1089_));
 sg13g2_nor4_1 _3882_ (.A(_1820_),
    .B(net1118),
    .C(_1084_),
    .D(_1089_),
    .Y(_1090_));
 sg13g2_nor2_1 _3883_ (.A(\charlie_0.memory[6][2] ),
    .B(net1046),
    .Y(_1091_));
 sg13g2_nor2_1 _3884_ (.A(\charlie_0.memory[6][1] ),
    .B(net1038),
    .Y(_1092_));
 sg13g2_nor2_1 _3885_ (.A(\charlie_0.memory[6][0] ),
    .B(net1073),
    .Y(_1093_));
 sg13g2_o21ai_1 _3886_ (.B1(net1116),
    .Y(_1094_),
    .A1(\charlie_0.memory[6][3] ),
    .A2(net1032));
 sg13g2_nor4_1 _3887_ (.A(_1091_),
    .B(_1092_),
    .C(_1093_),
    .D(_1094_),
    .Y(_1095_));
 sg13g2_o21ai_1 _3888_ (.B1(net1179),
    .Y(_1096_),
    .A1(\charlie_0.memory[6][5] ),
    .A2(net1038));
 sg13g2_nor2_1 _3889_ (.A(\charlie_0.memory[6][6] ),
    .B(net1046),
    .Y(_1097_));
 sg13g2_nor2_1 _3890_ (.A(\charlie_0.memory[6][7] ),
    .B(net1032),
    .Y(_1098_));
 sg13g2_nor2_1 _3891_ (.A(\charlie_0.memory[6][4] ),
    .B(net1073),
    .Y(_1099_));
 sg13g2_nor4_1 _3892_ (.A(_1096_),
    .B(_1097_),
    .C(_1098_),
    .D(_1099_),
    .Y(_1100_));
 sg13g2_nor3_1 _3893_ (.A(_1045_),
    .B(_1095_),
    .C(_1100_),
    .Y(_1101_));
 sg13g2_or3_2 _3894_ (.A(_1819_),
    .B(_1090_),
    .C(_1101_),
    .X(_1102_));
 sg13g2_o21ai_1 _3895_ (.B1(_0806_),
    .Y(_1103_),
    .A1(_1079_),
    .A2(_1102_));
 sg13g2_o21ai_1 _3896_ (.B1(_0811_),
    .Y(_1104_),
    .A1(_1056_),
    .A2(_1103_));
 sg13g2_o21ai_1 _3897_ (.B1(net1113),
    .Y(_1105_),
    .A1(\charlie_0.memory[10][2] ),
    .A2(net1043));
 sg13g2_a221oi_1 _3898_ (.B2(_1801_),
    .C1(_1105_),
    .B1(net1041),
    .A1(_1802_),
    .Y(_1106_),
    .A2(net1076));
 sg13g2_o21ai_1 _3899_ (.B1(_1106_),
    .Y(_1107_),
    .A1(\charlie_0.memory[10][3] ),
    .A2(net1029));
 sg13g2_nor2_1 _3900_ (.A(\charlie_0.memory[10][4] ),
    .B(net1070),
    .Y(_1108_));
 sg13g2_a21oi_1 _3901_ (.A1(_1798_),
    .A2(net1041),
    .Y(_1109_),
    .B1(net1113));
 sg13g2_a22oi_1 _3902_ (.Y(_1110_),
    .B1(net1035),
    .B2(_1796_),
    .A2(net1049),
    .A1(_1797_));
 sg13g2_nand3b_1 _3903_ (.B(_1109_),
    .C(_1110_),
    .Y(_1111_),
    .A_N(_1108_));
 sg13g2_nand3_1 _3904_ (.B(_1107_),
    .C(_1111_),
    .A(net1175),
    .Y(_1112_));
 sg13g2_o21ai_1 _3905_ (.B1(net1178),
    .Y(_1113_),
    .A1(\charlie_0.memory[8][4] ),
    .A2(net1070));
 sg13g2_nor2_1 _3906_ (.A(\charlie_0.memory[8][6] ),
    .B(net1043),
    .Y(_1114_));
 sg13g2_nor2_1 _3907_ (.A(\charlie_0.memory[8][7] ),
    .B(net1030),
    .Y(_1115_));
 sg13g2_nor2_1 _3908_ (.A(\charlie_0.memory[8][5] ),
    .B(net1036),
    .Y(_1116_));
 sg13g2_nor4_1 _3909_ (.A(_1113_),
    .B(_1114_),
    .C(_1115_),
    .D(_1116_),
    .Y(_1117_));
 sg13g2_o21ai_1 _3910_ (.B1(net1113),
    .Y(_1118_),
    .A1(\charlie_0.memory[8][0] ),
    .A2(net1070));
 sg13g2_nor2_1 _3911_ (.A(\charlie_0.memory[8][3] ),
    .B(net1030),
    .Y(_1119_));
 sg13g2_nor2_1 _3912_ (.A(\charlie_0.memory[8][2] ),
    .B(net1043),
    .Y(_1120_));
 sg13g2_nor2_1 _3913_ (.A(\charlie_0.memory[8][1] ),
    .B(net1036),
    .Y(_1121_));
 sg13g2_nor4_1 _3914_ (.A(_1118_),
    .B(_1119_),
    .C(_1120_),
    .D(_1121_),
    .Y(_1122_));
 sg13g2_nor3_1 _3915_ (.A(net1175),
    .B(_1117_),
    .C(_1122_),
    .Y(_1123_));
 sg13g2_nor2_1 _3916_ (.A(net1177),
    .B(_1123_),
    .Y(_1124_));
 sg13g2_nor2_1 _3917_ (.A(\charlie_0.memory[11][7] ),
    .B(net1029),
    .Y(_1125_));
 sg13g2_nor2_1 _3918_ (.A(\charlie_0.memory[11][5] ),
    .B(net1037),
    .Y(_1126_));
 sg13g2_o21ai_1 _3919_ (.B1(net1178),
    .Y(_1127_),
    .A1(\charlie_0.memory[11][6] ),
    .A2(net1043));
 sg13g2_nor3_1 _3920_ (.A(_1125_),
    .B(_1126_),
    .C(_1127_),
    .Y(_1128_));
 sg13g2_o21ai_1 _3921_ (.B1(_1128_),
    .Y(_1129_),
    .A1(\charlie_0.memory[11][4] ),
    .A2(net1070));
 sg13g2_nor2_1 _3922_ (.A(\charlie_0.memory[11][0] ),
    .B(net1070),
    .Y(_1130_));
 sg13g2_nor2_1 _3923_ (.A(\charlie_0.memory[11][2] ),
    .B(net1043),
    .Y(_1131_));
 sg13g2_nor2_1 _3924_ (.A(\charlie_0.memory[11][1] ),
    .B(net1036),
    .Y(_1132_));
 sg13g2_o21ai_1 _3925_ (.B1(net1113),
    .Y(_1133_),
    .A1(\charlie_0.memory[11][3] ),
    .A2(net1029));
 sg13g2_or4_1 _3926_ (.A(_1130_),
    .B(_1131_),
    .C(_1132_),
    .D(_1133_),
    .X(_1134_));
 sg13g2_nand3_1 _3927_ (.B(_1129_),
    .C(_1134_),
    .A(net1175),
    .Y(_1135_));
 sg13g2_nor2_1 _3928_ (.A(\charlie_0.memory[9][0] ),
    .B(net1070),
    .Y(_1136_));
 sg13g2_nor2_1 _3929_ (.A(\charlie_0.memory[9][1] ),
    .B(net1036),
    .Y(_1137_));
 sg13g2_nor2_1 _3930_ (.A(\charlie_0.memory[9][2] ),
    .B(net1043),
    .Y(_1138_));
 sg13g2_o21ai_1 _3931_ (.B1(net1113),
    .Y(_1139_),
    .A1(\charlie_0.memory[9][3] ),
    .A2(net1029));
 sg13g2_nor4_1 _3932_ (.A(_1136_),
    .B(_1137_),
    .C(_1138_),
    .D(_1139_),
    .Y(_1140_));
 sg13g2_nor2_1 _3933_ (.A(\charlie_0.memory[9][5] ),
    .B(net1036),
    .Y(_1141_));
 sg13g2_nor2_1 _3934_ (.A(\charlie_0.memory[9][4] ),
    .B(net1070),
    .Y(_1142_));
 sg13g2_nor2_1 _3935_ (.A(\charlie_0.memory[9][7] ),
    .B(net1029),
    .Y(_1143_));
 sg13g2_o21ai_1 _3936_ (.B1(net1178),
    .Y(_1144_),
    .A1(\charlie_0.memory[9][6] ),
    .A2(net1043));
 sg13g2_nor4_1 _3937_ (.A(_1141_),
    .B(_1142_),
    .C(_1143_),
    .D(_1144_),
    .Y(_1145_));
 sg13g2_nor3_1 _3938_ (.A(net1175),
    .B(_1140_),
    .C(_1145_),
    .Y(_1146_));
 sg13g2_nor2_1 _3939_ (.A(net1118),
    .B(_1146_),
    .Y(_1147_));
 sg13g2_a22oi_1 _3940_ (.Y(_1148_),
    .B1(_1135_),
    .B2(_1147_),
    .A2(_1124_),
    .A1(_1112_));
 sg13g2_nor2_1 _3941_ (.A(\charlie_0.memory[12][0] ),
    .B(net1071),
    .Y(_1149_));
 sg13g2_nor2_1 _3942_ (.A(\charlie_0.memory[12][1] ),
    .B(net1037),
    .Y(_1150_));
 sg13g2_nor2_1 _3943_ (.A(\charlie_0.memory[12][3] ),
    .B(net1030),
    .Y(_1151_));
 sg13g2_o21ai_1 _3944_ (.B1(net1114),
    .Y(_1152_),
    .A1(\charlie_0.memory[12][2] ),
    .A2(net1044));
 sg13g2_nor4_1 _3945_ (.A(_1149_),
    .B(_1150_),
    .C(_1151_),
    .D(_1152_),
    .Y(_1153_));
 sg13g2_nor2_1 _3946_ (.A(\charlie_0.memory[12][4] ),
    .B(net1071),
    .Y(_1154_));
 sg13g2_nor2_1 _3947_ (.A(\charlie_0.memory[12][5] ),
    .B(net1037),
    .Y(_1155_));
 sg13g2_nor2_1 _3948_ (.A(\charlie_0.memory[12][6] ),
    .B(net1044),
    .Y(_1156_));
 sg13g2_o21ai_1 _3949_ (.B1(net1178),
    .Y(_1157_),
    .A1(\charlie_0.memory[12][7] ),
    .A2(net1031));
 sg13g2_nor4_1 _3950_ (.A(_1154_),
    .B(_1155_),
    .C(_1156_),
    .D(_1157_),
    .Y(_1158_));
 sg13g2_nor3_1 _3951_ (.A(net1175),
    .B(_1153_),
    .C(_1158_),
    .Y(_1159_));
 sg13g2_a22oi_1 _3952_ (.Y(_1160_),
    .B1(net1049),
    .B2(_1793_),
    .A2(net1076),
    .A1(_1795_));
 sg13g2_a221oi_1 _3953_ (.B2(_1792_),
    .C1(net1113),
    .B1(net1035),
    .A1(_1794_),
    .Y(_1161_),
    .A2(net1041));
 sg13g2_nand2_1 _3954_ (.Y(_1162_),
    .A(_1160_),
    .B(_1161_));
 sg13g2_nor2_1 _3955_ (.A(\charlie_0.memory[14][0] ),
    .B(net1070),
    .Y(_1163_));
 sg13g2_nor2_1 _3956_ (.A(\charlie_0.memory[14][2] ),
    .B(net1043),
    .Y(_1164_));
 sg13g2_o21ai_1 _3957_ (.B1(net1114),
    .Y(_1165_),
    .A1(\charlie_0.memory[14][3] ),
    .A2(net1029));
 sg13g2_nor3_1 _3958_ (.A(_1163_),
    .B(_1164_),
    .C(_1165_),
    .Y(_1166_));
 sg13g2_o21ai_1 _3959_ (.B1(_1166_),
    .Y(_1167_),
    .A1(\charlie_0.memory[14][1] ),
    .A2(net1036));
 sg13g2_nand3_1 _3960_ (.B(_1162_),
    .C(_1167_),
    .A(net1175),
    .Y(_1168_));
 sg13g2_nor2_1 _3961_ (.A(net1177),
    .B(_1159_),
    .Y(_1169_));
 sg13g2_o21ai_1 _3962_ (.B1(net1178),
    .Y(_1170_),
    .A1(\charlie_0.memory[15][4] ),
    .A2(net1071));
 sg13g2_nor2_1 _3963_ (.A(\charlie_0.memory[15][6] ),
    .B(net1044),
    .Y(_1171_));
 sg13g2_nor2_1 _3964_ (.A(\charlie_0.memory[15][7] ),
    .B(net1030),
    .Y(_1172_));
 sg13g2_nor2_1 _3965_ (.A(\charlie_0.memory[15][5] ),
    .B(net1037),
    .Y(_1173_));
 sg13g2_nor4_1 _3966_ (.A(_1170_),
    .B(_1171_),
    .C(_1172_),
    .D(_1173_),
    .Y(_1174_));
 sg13g2_o21ai_1 _3967_ (.B1(net1114),
    .Y(_1175_),
    .A1(\charlie_0.memory[15][2] ),
    .A2(net1044));
 sg13g2_nor2_1 _3968_ (.A(\charlie_0.memory[15][0] ),
    .B(net1071),
    .Y(_1176_));
 sg13g2_nor2_1 _3969_ (.A(\charlie_0.memory[15][1] ),
    .B(net1037),
    .Y(_1177_));
 sg13g2_nor2_1 _3970_ (.A(\charlie_0.memory[15][3] ),
    .B(net1030),
    .Y(_1178_));
 sg13g2_nor4_1 _3971_ (.A(_1175_),
    .B(_1176_),
    .C(_1177_),
    .D(_1178_),
    .Y(_1179_));
 sg13g2_nor3_1 _3972_ (.A(_1820_),
    .B(_1174_),
    .C(_1179_),
    .Y(_1180_));
 sg13g2_nor2_1 _3973_ (.A(\charlie_0.memory[13][1] ),
    .B(net1037),
    .Y(_1181_));
 sg13g2_nor2_1 _3974_ (.A(\charlie_0.memory[13][2] ),
    .B(net1044),
    .Y(_1182_));
 sg13g2_nor2_1 _3975_ (.A(\charlie_0.memory[13][3] ),
    .B(net1030),
    .Y(_1183_));
 sg13g2_o21ai_1 _3976_ (.B1(net1114),
    .Y(_1184_),
    .A1(\charlie_0.memory[13][0] ),
    .A2(net1071));
 sg13g2_nor4_1 _3977_ (.A(_1181_),
    .B(_1182_),
    .C(_1183_),
    .D(_1184_),
    .Y(_1185_));
 sg13g2_nor2_1 _3978_ (.A(\charlie_0.memory[13][5] ),
    .B(net1036),
    .Y(_1186_));
 sg13g2_nor2_1 _3979_ (.A(\charlie_0.memory[13][4] ),
    .B(net1071),
    .Y(_1187_));
 sg13g2_nor2_1 _3980_ (.A(\charlie_0.memory[13][7] ),
    .B(net1030),
    .Y(_1188_));
 sg13g2_o21ai_1 _3981_ (.B1(net1178),
    .Y(_1189_),
    .A1(\charlie_0.memory[13][6] ),
    .A2(net1044));
 sg13g2_nor4_1 _3982_ (.A(_1186_),
    .B(_1187_),
    .C(_1188_),
    .D(_1189_),
    .Y(_1190_));
 sg13g2_or3_1 _3983_ (.A(net1175),
    .B(_1185_),
    .C(_1190_),
    .X(_1191_));
 sg13g2_nor2_1 _3984_ (.A(net1118),
    .B(_1180_),
    .Y(_1192_));
 sg13g2_a221oi_1 _3985_ (.B2(_1192_),
    .C1(_1819_),
    .B1(_1191_),
    .A1(_1168_),
    .Y(_1193_),
    .A2(_1169_));
 sg13g2_o21ai_1 _3986_ (.B1(net1113),
    .Y(_1194_),
    .A1(net1171),
    .A2(net1036));
 sg13g2_a22oi_1 _3987_ (.Y(_1195_),
    .B1(net1049),
    .B2(_1789_),
    .A2(net1076),
    .A1(_1791_));
 sg13g2_o21ai_1 _3988_ (.B1(_1195_),
    .Y(_1196_),
    .A1(\charlie_0.memory[16][3] ),
    .A2(net1029));
 sg13g2_nor2_1 _3989_ (.A(\charlie_0.memory[16][7] ),
    .B(net1029),
    .Y(_1197_));
 sg13g2_a21oi_1 _3990_ (.A1(net1120),
    .A2(net1049),
    .Y(_1198_),
    .B1(net1113));
 sg13g2_a221oi_1 _3991_ (.B2(_1786_),
    .C1(_1197_),
    .B1(net1041),
    .A1(_1787_),
    .Y(_1199_),
    .A2(net1076));
 sg13g2_a21oi_1 _3992_ (.A1(_1198_),
    .A2(_1199_),
    .Y(_1200_),
    .B1(net1177));
 sg13g2_o21ai_1 _3993_ (.B1(_1200_),
    .Y(_1201_),
    .A1(_1194_),
    .A2(_1196_));
 sg13g2_a22oi_1 _3994_ (.Y(_1202_),
    .B1(net1042),
    .B2(_1783_),
    .A2(net1050),
    .A1(net1123));
 sg13g2_a221oi_1 _3995_ (.B2(_1781_),
    .C1(net1179),
    .B1(net1035),
    .A1(_1784_),
    .Y(_1203_),
    .A2(net1077));
 sg13g2_nand2_1 _3996_ (.Y(_1204_),
    .A(_1202_),
    .B(_1203_));
 sg13g2_a21oi_1 _3997_ (.A1(_1779_),
    .A2(net1042),
    .Y(_1205_),
    .B1(net1116));
 sg13g2_nor2_1 _3998_ (.A(\charlie_0.memory[17][7] ),
    .B(net1033),
    .Y(_1206_));
 sg13g2_a221oi_1 _3999_ (.B2(_1778_),
    .C1(_1206_),
    .B1(net1050),
    .A1(_1780_),
    .Y(_1207_),
    .A2(net1077));
 sg13g2_a21oi_1 _4000_ (.A1(_1205_),
    .A2(_1207_),
    .Y(_1208_),
    .B1(net1118));
 sg13g2_a21oi_1 _4001_ (.A1(_1204_),
    .A2(_1208_),
    .Y(_1209_),
    .B1(net1176));
 sg13g2_nor2_1 _4002_ (.A(\charlie_0.memory[18][4] ),
    .B(net1075),
    .Y(_1210_));
 sg13g2_nor2_1 _4003_ (.A(\charlie_0.memory[18][6] ),
    .B(net1048),
    .Y(_1211_));
 sg13g2_nor2_1 _4004_ (.A(\charlie_0.memory[18][7] ),
    .B(net1033),
    .Y(_1212_));
 sg13g2_o21ai_1 _4005_ (.B1(net1180),
    .Y(_1213_),
    .A1(\charlie_0.memory[18][5] ),
    .A2(net1039));
 sg13g2_nor4_1 _4006_ (.A(_1210_),
    .B(_1211_),
    .C(_1212_),
    .D(_1213_),
    .Y(_1214_));
 sg13g2_o21ai_1 _4007_ (.B1(net1116),
    .Y(_1215_),
    .A1(\charlie_0.memory[18][1] ),
    .A2(net1039));
 sg13g2_nor2_1 _4008_ (.A(\charlie_0.memory[18][2] ),
    .B(net1047),
    .Y(_1216_));
 sg13g2_nor2_1 _4009_ (.A(\charlie_0.memory[18][3] ),
    .B(net1034),
    .Y(_1217_));
 sg13g2_nor2_1 _4010_ (.A(\charlie_0.memory[18][0] ),
    .B(net1075),
    .Y(_1218_));
 sg13g2_nor4_1 _4011_ (.A(_1215_),
    .B(_1216_),
    .C(_1217_),
    .D(_1218_),
    .Y(_1219_));
 sg13g2_nor2_1 _4012_ (.A(\charlie_0.memory[19][7] ),
    .B(net1031),
    .Y(_1220_));
 sg13g2_nor2_1 _4013_ (.A(net1148),
    .B(net1072),
    .Y(_1221_));
 sg13g2_nor2_1 _4014_ (.A(\charlie_0.memory[19][6] ),
    .B(net1045),
    .Y(_1222_));
 sg13g2_o21ai_1 _4015_ (.B1(net1181),
    .Y(_1223_),
    .A1(\charlie_0.memory[19][5] ),
    .A2(net1040));
 sg13g2_nor4_1 _4016_ (.A(_1220_),
    .B(_1221_),
    .C(_1222_),
    .D(_1223_),
    .Y(_1224_));
 sg13g2_nor2_1 _4017_ (.A(net1150),
    .B(net1031),
    .Y(_1225_));
 sg13g2_nor2_1 _4018_ (.A(\bi_frame_index[0] ),
    .B(net1072),
    .Y(_1226_));
 sg13g2_nor2_1 _4019_ (.A(net1153),
    .B(net1040),
    .Y(_1227_));
 sg13g2_o21ai_1 _4020_ (.B1(net1115),
    .Y(_1228_),
    .A1(net1151),
    .A2(net1045));
 sg13g2_nor4_1 _4021_ (.A(_1225_),
    .B(_1226_),
    .C(_1227_),
    .D(_1228_),
    .Y(_1229_));
 sg13g2_or3_1 _4022_ (.A(\signal_generator_0.index_reg[3] ),
    .B(_1214_),
    .C(_1219_),
    .X(_1230_));
 sg13g2_nor3_2 _4023_ (.A(net1118),
    .B(_1224_),
    .C(_1229_),
    .Y(_1231_));
 sg13g2_nor2_1 _4024_ (.A(_1820_),
    .B(_1231_),
    .Y(_1232_));
 sg13g2_a22oi_1 _4025_ (.Y(_1233_),
    .B1(_1230_),
    .B2(_1232_),
    .A2(_1209_),
    .A1(_1201_));
 sg13g2_nand2_1 _4026_ (.Y(_1234_),
    .A(\charlie_0.memory[21][4] ),
    .B(net1076));
 sg13g2_a22oi_1 _4027_ (.Y(_1235_),
    .B1(net1041),
    .B2(\charlie_0.memory[20][5] ),
    .A2(net1076),
    .A1(\charlie_0.memory[20][4] ));
 sg13g2_a21oi_1 _4028_ (.A1(\charlie_0.memory[21][7] ),
    .A2(net1035),
    .Y(_1236_),
    .B1(net1115));
 sg13g2_a22oi_1 _4029_ (.Y(_1237_),
    .B1(net1041),
    .B2(\charlie_0.memory[21][5] ),
    .A2(net1050),
    .A1(\charlie_0.memory[21][6] ));
 sg13g2_nand3_1 _4030_ (.B(_1236_),
    .C(_1237_),
    .A(_1234_),
    .Y(_1238_));
 sg13g2_a22oi_1 _4031_ (.Y(_1239_),
    .B1(net1042),
    .B2(\charlie_0.memory[21][1] ),
    .A2(net1049),
    .A1(\charlie_0.memory[21][2] ));
 sg13g2_a221oi_1 _4032_ (.B2(\charlie_0.memory[21][3] ),
    .C1(net1181),
    .B1(net1035),
    .A1(\charlie_0.memory[21][0] ),
    .Y(_1240_),
    .A2(net1077));
 sg13g2_a21oi_1 _4033_ (.A1(_1239_),
    .A2(_1240_),
    .Y(_1241_),
    .B1(net1118));
 sg13g2_nand2_1 _4034_ (.Y(_1242_),
    .A(_1238_),
    .B(_1241_));
 sg13g2_a22oi_1 _4035_ (.Y(_1243_),
    .B1(net1035),
    .B2(\charlie_0.memory[20][3] ),
    .A2(net1041),
    .A1(\charlie_0.memory[20][1] ));
 sg13g2_a221oi_1 _4036_ (.B2(\charlie_0.memory[20][2] ),
    .C1(net1178),
    .B1(net1049),
    .A1(\charlie_0.memory[20][0] ),
    .Y(_1244_),
    .A2(net1076));
 sg13g2_nand2_1 _4037_ (.Y(_1245_),
    .A(_1243_),
    .B(_1244_));
 sg13g2_a22oi_1 _4038_ (.Y(_1246_),
    .B1(net1035),
    .B2(\charlie_0.memory[20][7] ),
    .A2(net1049),
    .A1(\charlie_0.memory[20][6] ));
 sg13g2_nand3_1 _4039_ (.B(_1235_),
    .C(_1246_),
    .A(net1178),
    .Y(_1247_));
 sg13g2_nand3_1 _4040_ (.B(_1245_),
    .C(_1247_),
    .A(net1118),
    .Y(_1248_));
 sg13g2_a21oi_2 _4041_ (.B1(net1175),
    .Y(_1249_),
    .A2(_1248_),
    .A1(_1242_));
 sg13g2_nand2_1 _4042_ (.Y(_1250_),
    .A(\charlie_0.memory[22][5] ),
    .B(net1041));
 sg13g2_a21oi_1 _4043_ (.A1(\charlie_0.memory[22][7] ),
    .A2(_1012_),
    .Y(_1251_),
    .B1(net1115));
 sg13g2_a22oi_1 _4044_ (.Y(_1252_),
    .B1(net1049),
    .B2(\charlie_0.memory[22][6] ),
    .A2(net1076),
    .A1(\charlie_0.memory[22][4] ));
 sg13g2_nand3_1 _4045_ (.B(_1251_),
    .C(_1252_),
    .A(_1250_),
    .Y(_1253_));
 sg13g2_mux4_1 _4046_ (.S0(net1183),
    .A0(net1146),
    .A1(\charlie_0.memory[22][1] ),
    .A2(\charlie_0.memory[22][2] ),
    .A3(\charlie_0.memory[22][3] ),
    .S1(net1182),
    .X(_1254_));
 sg13g2_o21ai_1 _4047_ (.B1(_1253_),
    .Y(_1255_),
    .A1(net1181),
    .A2(_1254_));
 sg13g2_o21ai_1 _4048_ (.B1(\signal_generator_0.index_reg[5] ),
    .Y(_1256_),
    .A1(_1045_),
    .A2(_1255_));
 sg13g2_o21ai_1 _4049_ (.B1(_1818_),
    .Y(_1257_),
    .A1(_1249_),
    .A2(_1256_));
 sg13g2_a21o_1 _4050_ (.A2(_1233_),
    .A1(_1819_),
    .B1(_1257_),
    .X(_1258_));
 sg13g2_a21o_2 _4051_ (.A2(_1148_),
    .A1(_1819_),
    .B1(_1193_),
    .X(_1259_));
 sg13g2_a221oi_1 _4052_ (.B2(\signal_generator_0.index_reg[6] ),
    .C1(_1104_),
    .B1(_1259_),
    .A1(\signal_generator_0.index_reg[7] ),
    .Y(_1260_),
    .A2(_1258_));
 sg13g2_nor2_1 _4053_ (.A(net954),
    .B(_0809_),
    .Y(_1261_));
 sg13g2_o21ai_1 _4054_ (.B1(_1261_),
    .Y(_1262_),
    .A1(_1005_),
    .A2(_1260_));
 sg13g2_a22oi_1 _4055_ (.Y(_1263_),
    .B1(_1004_),
    .B2(net953),
    .A2(_1001_),
    .A1(_0810_));
 sg13g2_a21oi_1 _4056_ (.A1(_1262_),
    .A2(_1263_),
    .Y(_0105_),
    .B1(net1226));
 sg13g2_and2_1 _4057_ (.A(net1240),
    .B(_2122_),
    .X(_0106_));
 sg13g2_nand2_2 _4058_ (.Y(_1264_),
    .A(net1021),
    .B(net953));
 sg13g2_nand2b_2 _4059_ (.Y(_1265_),
    .B(_1264_),
    .A_N(_1261_));
 sg13g2_nor2_1 _4060_ (.A(net278),
    .B(_1265_),
    .Y(_1266_));
 sg13g2_nor2_1 _4061_ (.A(net1183),
    .B(_1264_),
    .Y(_1267_));
 sg13g2_and2_2 _4062_ (.A(_0807_),
    .B(_0811_),
    .X(_1268_));
 sg13g2_nor3_1 _4063_ (.A(_0049_),
    .B(_0809_),
    .C(_1268_),
    .Y(_1269_));
 sg13g2_a21oi_1 _4064_ (.A1(_1836_),
    .A2(_1268_),
    .Y(_1270_),
    .B1(_1269_));
 sg13g2_o21ai_1 _4065_ (.B1(net1257),
    .Y(_1271_),
    .A1(net954),
    .A2(_1270_));
 sg13g2_nor3_1 _4066_ (.A(_1266_),
    .B(_1267_),
    .C(_1271_),
    .Y(_0107_));
 sg13g2_nor3_1 _4067_ (.A(_0824_),
    .B(_0826_),
    .C(_1265_),
    .Y(_1272_));
 sg13g2_xor2_1 _4068_ (.B(\charlie_0.memory[18][0] ),
    .A(\charlie_0.memory[18][1] ),
    .X(_1273_));
 sg13g2_a22oi_1 _4069_ (.Y(_1274_),
    .B1(_1268_),
    .B2(_1273_),
    .A2(net1033),
    .A1(net1074));
 sg13g2_o21ai_1 _4070_ (.B1(net1256),
    .Y(_1275_),
    .A1(net954),
    .A2(_1274_));
 sg13g2_nor2_1 _4071_ (.A(net1182),
    .B(_1264_),
    .Y(_1276_));
 sg13g2_nor3_1 _4072_ (.A(_1272_),
    .B(_1275_),
    .C(_1276_),
    .Y(_0108_));
 sg13g2_nor2_1 _4073_ (.A(net1122),
    .B(_0824_),
    .Y(_1277_));
 sg13g2_nor2_1 _4074_ (.A(net1159),
    .B(net1059),
    .Y(_1278_));
 sg13g2_nor3_1 _4075_ (.A(_1265_),
    .B(_1277_),
    .C(_1278_),
    .Y(_1279_));
 sg13g2_nor2_1 _4076_ (.A(net1180),
    .B(_1264_),
    .Y(_1280_));
 sg13g2_xnor2_1 _4077_ (.Y(_1281_),
    .A(net1116),
    .B(net1077));
 sg13g2_or3_2 _4078_ (.A(\charlie_0.memory[18][2] ),
    .B(\charlie_0.memory[18][1] ),
    .C(\charlie_0.memory[18][0] ),
    .X(_1282_));
 sg13g2_o21ai_1 _4079_ (.B1(\charlie_0.memory[18][2] ),
    .Y(_1283_),
    .A1(\charlie_0.memory[18][1] ),
    .A2(\charlie_0.memory[18][0] ));
 sg13g2_nand3_1 _4080_ (.B(_1282_),
    .C(_1283_),
    .A(_1268_),
    .Y(_1284_));
 sg13g2_a21oi_1 _4081_ (.A1(_1281_),
    .A2(_1284_),
    .Y(_1285_),
    .B1(net954));
 sg13g2_nor4_1 _4082_ (.A(net1226),
    .B(_1279_),
    .C(_1280_),
    .D(_1285_),
    .Y(_0109_));
 sg13g2_nor3_1 _4083_ (.A(net1156),
    .B(net1159),
    .C(net1059),
    .Y(_1286_));
 sg13g2_xnor2_1 _4084_ (.Y(_1287_),
    .A(net1156),
    .B(_1278_));
 sg13g2_o21ai_1 _4085_ (.B1(net1177),
    .Y(_1288_),
    .A1(net1180),
    .A2(net1074));
 sg13g2_nand2b_1 _4086_ (.Y(_1289_),
    .B(_1288_),
    .A_N(_0801_));
 sg13g2_o21ai_1 _4087_ (.B1(_0807_),
    .Y(_1290_),
    .A1(_0795_),
    .A2(_0811_));
 sg13g2_a21oi_1 _4088_ (.A1(_1289_),
    .A2(_1290_),
    .Y(_1291_),
    .B1(net954));
 sg13g2_a21oi_1 _4089_ (.A1(_0565_),
    .A2(_1287_),
    .Y(_1292_),
    .B1(_1291_));
 sg13g2_nand2_1 _4090_ (.Y(_1293_),
    .A(_0795_),
    .B(_0812_));
 sg13g2_xnor2_1 _4091_ (.Y(_1294_),
    .A(\charlie_0.memory[18][3] ),
    .B(_1282_));
 sg13g2_nand2_1 _4092_ (.Y(_1295_),
    .A(_0811_),
    .B(_1294_));
 sg13g2_and2_1 _4093_ (.A(_0813_),
    .B(_1295_),
    .X(_1296_));
 sg13g2_o21ai_1 _4094_ (.B1(_1296_),
    .Y(_1297_),
    .A1(_1287_),
    .A2(_1293_));
 sg13g2_a21oi_1 _4095_ (.A1(_0808_),
    .A2(_1297_),
    .Y(_1298_),
    .B1(_1292_));
 sg13g2_o21ai_1 _4096_ (.B1(net1257),
    .Y(_1299_),
    .A1(net1177),
    .A2(_1264_));
 sg13g2_nor2_1 _4097_ (.A(_1298_),
    .B(_1299_),
    .Y(_0110_));
 sg13g2_xnor2_1 _4098_ (.Y(_1300_),
    .A(_1820_),
    .B(_0801_));
 sg13g2_nor3_2 _4099_ (.A(\charlie_0.memory[18][4] ),
    .B(\charlie_0.memory[18][3] ),
    .C(_1282_),
    .Y(_1301_));
 sg13g2_o21ai_1 _4100_ (.B1(\charlie_0.memory[18][4] ),
    .Y(_1302_),
    .A1(\charlie_0.memory[18][3] ),
    .A2(_1282_));
 sg13g2_nor2b_1 _4101_ (.A(_1301_),
    .B_N(_1302_),
    .Y(_1303_));
 sg13g2_and2_1 _4102_ (.A(_1780_),
    .B(_1286_),
    .X(_1304_));
 sg13g2_xnor2_1 _4103_ (.Y(_1305_),
    .A(\charlie_0.memory[17][4] ),
    .B(_1286_));
 sg13g2_a21o_1 _4104_ (.A2(_1305_),
    .A1(_0809_),
    .B1(_1268_),
    .X(_1306_));
 sg13g2_o21ai_1 _4105_ (.B1(_1306_),
    .Y(_1307_),
    .A1(_0812_),
    .A2(_1303_));
 sg13g2_a21oi_1 _4106_ (.A1(_1300_),
    .A2(_1307_),
    .Y(_1308_),
    .B1(net954));
 sg13g2_nand2_1 _4107_ (.Y(_1309_),
    .A(_0565_),
    .B(_1305_));
 sg13g2_o21ai_1 _4108_ (.B1(_1309_),
    .Y(_1310_),
    .A1(net1176),
    .A2(_1264_));
 sg13g2_nor3_1 _4109_ (.A(net1226),
    .B(_1308_),
    .C(_1310_),
    .Y(_0111_));
 sg13g2_nor2_1 _4110_ (.A(net319),
    .B(_1264_),
    .Y(_1311_));
 sg13g2_nor2b_1 _4111_ (.A(\charlie_0.memory[18][5] ),
    .B_N(_1301_),
    .Y(_1312_));
 sg13g2_xnor2_1 _4112_ (.Y(_1313_),
    .A(\charlie_0.memory[18][5] ),
    .B(_1301_));
 sg13g2_xnor2_1 _4113_ (.Y(_1314_),
    .A(\signal_generator_0.index_reg[5] ),
    .B(_0802_));
 sg13g2_and2_1 _4114_ (.A(_1779_),
    .B(_1304_),
    .X(_1315_));
 sg13g2_xnor2_1 _4115_ (.Y(_1316_),
    .A(_1779_),
    .B(_1304_));
 sg13g2_nand2_1 _4116_ (.Y(_1317_),
    .A(_0795_),
    .B(_1316_));
 sg13g2_a221oi_1 _4117_ (.B2(_0809_),
    .C1(_1314_),
    .B1(_1317_),
    .A1(_1268_),
    .Y(_1318_),
    .A2(_1313_));
 sg13g2_nor2_1 _4118_ (.A(net1021),
    .B(_1316_),
    .Y(_1319_));
 sg13g2_o21ai_1 _4119_ (.B1(net1257),
    .Y(_1320_),
    .A1(net953),
    .A2(_1318_));
 sg13g2_nor3_1 _4120_ (.A(_1311_),
    .B(_1319_),
    .C(_1320_),
    .Y(_0112_));
 sg13g2_nand3_1 _4121_ (.B(net1021),
    .C(net953),
    .A(net308),
    .Y(_1321_));
 sg13g2_and2_1 _4122_ (.A(_1778_),
    .B(_1315_),
    .X(_1322_));
 sg13g2_nand2_1 _4123_ (.Y(_1323_),
    .A(_1778_),
    .B(_1315_));
 sg13g2_xnor2_1 _4124_ (.Y(_1324_),
    .A(\charlie_0.memory[17][6] ),
    .B(_1315_));
 sg13g2_inv_1 _4125_ (.Y(_1325_),
    .A(_1324_));
 sg13g2_nand2_1 _4126_ (.Y(_1326_),
    .A(net308),
    .B(_0803_));
 sg13g2_nand2b_1 _4127_ (.Y(_1327_),
    .B(\charlie_0.memory[18][6] ),
    .A_N(_1312_));
 sg13g2_nor2b_1 _4128_ (.A(\charlie_0.memory[18][6] ),
    .B_N(_1312_),
    .Y(_1328_));
 sg13g2_nor2_1 _4129_ (.A(_0812_),
    .B(_1328_),
    .Y(_1329_));
 sg13g2_a22oi_1 _4130_ (.Y(_1330_),
    .B1(_1327_),
    .B2(_1329_),
    .A2(_1324_),
    .A1(_0796_));
 sg13g2_o21ai_1 _4131_ (.B1(_0804_),
    .Y(_1331_),
    .A1(\signal_generator_0.index_reg[7] ),
    .A2(_1330_));
 sg13g2_a21oi_1 _4132_ (.A1(_1326_),
    .A2(_1331_),
    .Y(_1332_),
    .B1(net953));
 sg13g2_a21oi_1 _4133_ (.A1(_0565_),
    .A2(_1325_),
    .Y(_1333_),
    .B1(_1332_));
 sg13g2_a21oi_1 _4134_ (.A1(_1321_),
    .A2(_1333_),
    .Y(_0113_),
    .B1(net1226));
 sg13g2_xnor2_1 _4135_ (.Y(_1334_),
    .A(\charlie_0.memory[18][7] ),
    .B(_1328_));
 sg13g2_a22oi_1 _4136_ (.Y(_1335_),
    .B1(_1334_),
    .B2(_0811_),
    .A2(_1323_),
    .A1(_0796_));
 sg13g2_and3_1 _4137_ (.X(_1336_),
    .A(net451),
    .B(net1021),
    .C(_0805_));
 sg13g2_a221oi_1 _4138_ (.B2(_0808_),
    .C1(_1336_),
    .B1(_1335_),
    .A1(_0565_),
    .Y(_1337_),
    .A2(_1322_));
 sg13g2_nor2_1 _4139_ (.A(net1226),
    .B(_1337_),
    .Y(_0114_));
 sg13g2_and2_1 _4140_ (.A(net1240),
    .B(_2037_),
    .X(_0115_));
 sg13g2_nor3_2 _4141_ (.A(\spi_address[2] ),
    .B(\spi_address[1] ),
    .C(\spi_address[0] ),
    .Y(_1338_));
 sg13g2_nor3_2 _4142_ (.A(\spi_address[4] ),
    .B(\spi_address[3] ),
    .C(_0571_),
    .Y(_1339_));
 sg13g2_and2_2 _4143_ (.A(_1338_),
    .B(_1339_),
    .X(_1340_));
 sg13g2_o21ai_1 _4144_ (.B1(net1251),
    .Y(_1341_),
    .A1(net318),
    .A2(net996));
 sg13g2_a21oi_1 _4145_ (.A1(net1228),
    .A2(net997),
    .Y(_0116_),
    .B1(_1341_));
 sg13g2_o21ai_1 _4146_ (.B1(net1251),
    .Y(_1342_),
    .A1(net312),
    .A2(net996));
 sg13g2_a21oi_1 _4147_ (.A1(net1126),
    .A2(net996),
    .Y(_0117_),
    .B1(_1342_));
 sg13g2_o21ai_1 _4148_ (.B1(net1253),
    .Y(_1343_),
    .A1(net330),
    .A2(net997));
 sg13g2_a21oi_1 _4149_ (.A1(net1131),
    .A2(net997),
    .Y(_0118_),
    .B1(_1343_));
 sg13g2_o21ai_1 _4150_ (.B1(net1251),
    .Y(_1344_),
    .A1(net327),
    .A2(_1340_));
 sg13g2_a21oi_1 _4151_ (.A1(net1135),
    .A2(net996),
    .Y(_0119_),
    .B1(_1344_));
 sg13g2_o21ai_1 _4152_ (.B1(net1253),
    .Y(_1345_),
    .A1(net317),
    .A2(net996));
 sg13g2_a21oi_1 _4153_ (.A1(net1138),
    .A2(net996),
    .Y(_0120_),
    .B1(_1345_));
 sg13g2_o21ai_1 _4154_ (.B1(net1251),
    .Y(_1346_),
    .A1(net324),
    .A2(net997));
 sg13g2_a21oi_1 _4155_ (.A1(net1141),
    .A2(net997),
    .Y(_0121_),
    .B1(_1346_));
 sg13g2_o21ai_1 _4156_ (.B1(net1251),
    .Y(_1347_),
    .A1(net316),
    .A2(net996));
 sg13g2_a21oi_1 _4157_ (.A1(net1142),
    .A2(net996),
    .Y(_0122_),
    .B1(_1347_));
 sg13g2_o21ai_1 _4158_ (.B1(net1251),
    .Y(_1348_),
    .A1(net329),
    .A2(net997));
 sg13g2_a21oi_1 _4159_ (.A1(net1144),
    .A2(net997),
    .Y(_0123_),
    .B1(_1348_));
 sg13g2_nand2b_1 _4160_ (.Y(_1349_),
    .B(\spi_address[0] ),
    .A_N(\spi_address[1] ));
 sg13g2_nor2_2 _4161_ (.A(\spi_address[2] ),
    .B(_1349_),
    .Y(_1350_));
 sg13g2_and2_1 _4162_ (.A(_1339_),
    .B(_1350_),
    .X(_1351_));
 sg13g2_o21ai_1 _4163_ (.B1(net1248),
    .Y(_1352_),
    .A1(net398),
    .A2(net995));
 sg13g2_a21oi_1 _4164_ (.A1(net1229),
    .A2(net995),
    .Y(_0124_),
    .B1(_1352_));
 sg13g2_o21ai_1 _4165_ (.B1(net1247),
    .Y(_1353_),
    .A1(net401),
    .A2(net994));
 sg13g2_a21oi_1 _4166_ (.A1(net1125),
    .A2(_1351_),
    .Y(_0125_),
    .B1(_1353_));
 sg13g2_o21ai_1 _4167_ (.B1(net1245),
    .Y(_1354_),
    .A1(net392),
    .A2(net995));
 sg13g2_a21oi_1 _4168_ (.A1(net1132),
    .A2(net995),
    .Y(_0126_),
    .B1(_1354_));
 sg13g2_o21ai_1 _4169_ (.B1(net1247),
    .Y(_1355_),
    .A1(net442),
    .A2(net994));
 sg13g2_a21oi_1 _4170_ (.A1(net1134),
    .A2(net995),
    .Y(_0127_),
    .B1(_1355_));
 sg13g2_o21ai_1 _4171_ (.B1(net1247),
    .Y(_1356_),
    .A1(net425),
    .A2(net994));
 sg13g2_a21oi_1 _4172_ (.A1(net1139),
    .A2(net994),
    .Y(_0128_),
    .B1(_1356_));
 sg13g2_o21ai_1 _4173_ (.B1(net1248),
    .Y(_1357_),
    .A1(net422),
    .A2(net995));
 sg13g2_a21oi_1 _4174_ (.A1(net1140),
    .A2(net995),
    .Y(_0129_),
    .B1(_1357_));
 sg13g2_o21ai_1 _4175_ (.B1(net1246),
    .Y(_1358_),
    .A1(net461),
    .A2(net994));
 sg13g2_a21oi_1 _4176_ (.A1(net1143),
    .A2(net994),
    .Y(_0130_),
    .B1(_1358_));
 sg13g2_o21ai_1 _4177_ (.B1(net1246),
    .Y(_1359_),
    .A1(net393),
    .A2(net994));
 sg13g2_a21oi_1 _4178_ (.A1(net1145),
    .A2(net994),
    .Y(_0131_),
    .B1(_1359_));
 sg13g2_nand2b_1 _4179_ (.Y(_1360_),
    .B(\spi_address[1] ),
    .A_N(\spi_address[0] ));
 sg13g2_nor2_2 _4180_ (.A(\spi_address[2] ),
    .B(_1360_),
    .Y(_1361_));
 sg13g2_and2_1 _4181_ (.A(_1339_),
    .B(_1361_),
    .X(_1362_));
 sg13g2_o21ai_1 _4182_ (.B1(net1248),
    .Y(_1363_),
    .A1(net407),
    .A2(net993));
 sg13g2_a21oi_1 _4183_ (.A1(net1229),
    .A2(net993),
    .Y(_0132_),
    .B1(_1363_));
 sg13g2_o21ai_1 _4184_ (.B1(net1245),
    .Y(_1364_),
    .A1(net431),
    .A2(_1362_));
 sg13g2_a21oi_1 _4185_ (.A1(_1775_),
    .A2(net992),
    .Y(_0133_),
    .B1(_1364_));
 sg13g2_o21ai_1 _4186_ (.B1(net1245),
    .Y(_1365_),
    .A1(net426),
    .A2(net993));
 sg13g2_a21oi_1 _4187_ (.A1(net1130),
    .A2(net993),
    .Y(_0134_),
    .B1(_1365_));
 sg13g2_o21ai_1 _4188_ (.B1(net1245),
    .Y(_1366_),
    .A1(net429),
    .A2(net992));
 sg13g2_a21oi_1 _4189_ (.A1(net1134),
    .A2(net992),
    .Y(_0135_),
    .B1(_1366_));
 sg13g2_o21ai_1 _4190_ (.B1(net1245),
    .Y(_1367_),
    .A1(net328),
    .A2(net992));
 sg13g2_a21oi_1 _4191_ (.A1(net1138),
    .A2(net993),
    .Y(_0136_),
    .B1(_1367_));
 sg13g2_o21ai_1 _4192_ (.B1(net1245),
    .Y(_1368_),
    .A1(net385),
    .A2(net993));
 sg13g2_a21oi_1 _4193_ (.A1(net1141),
    .A2(net993),
    .Y(_0137_),
    .B1(_1368_));
 sg13g2_o21ai_1 _4194_ (.B1(net1245),
    .Y(_1369_),
    .A1(net337),
    .A2(net992));
 sg13g2_a21oi_1 _4195_ (.A1(net1142),
    .A2(net992),
    .Y(_0138_),
    .B1(_1369_));
 sg13g2_o21ai_1 _4196_ (.B1(net1245),
    .Y(_1370_),
    .A1(net325),
    .A2(net992));
 sg13g2_a21oi_1 _4197_ (.A1(net1144),
    .A2(net992),
    .Y(_0139_),
    .B1(_1370_));
 sg13g2_nand2_1 _4198_ (.Y(_1371_),
    .A(\spi_address[1] ),
    .B(\spi_address[0] ));
 sg13g2_nor2_2 _4199_ (.A(\spi_address[2] ),
    .B(_1371_),
    .Y(_1372_));
 sg13g2_and2_1 _4200_ (.A(_1339_),
    .B(_1372_),
    .X(_1373_));
 sg13g2_o21ai_1 _4201_ (.B1(net1256),
    .Y(_1374_),
    .A1(net365),
    .A2(net991));
 sg13g2_a21oi_1 _4202_ (.A1(net1228),
    .A2(net991),
    .Y(_0140_),
    .B1(_1374_));
 sg13g2_o21ai_1 _4203_ (.B1(net1254),
    .Y(_1375_),
    .A1(net394),
    .A2(net991));
 sg13g2_a21oi_1 _4204_ (.A1(_1775_),
    .A2(_1373_),
    .Y(_0141_),
    .B1(_1375_));
 sg13g2_o21ai_1 _4205_ (.B1(net1256),
    .Y(_1376_),
    .A1(net448),
    .A2(net991));
 sg13g2_a21oi_1 _4206_ (.A1(net1131),
    .A2(net991),
    .Y(_0142_),
    .B1(_1376_));
 sg13g2_o21ai_1 _4207_ (.B1(net1254),
    .Y(_1377_),
    .A1(net427),
    .A2(net990));
 sg13g2_a21oi_1 _4208_ (.A1(net1135),
    .A2(net990),
    .Y(_0143_),
    .B1(_1377_));
 sg13g2_o21ai_1 _4209_ (.B1(net1254),
    .Y(_1378_),
    .A1(net453),
    .A2(net990));
 sg13g2_a21oi_1 _4210_ (.A1(net1138),
    .A2(net990),
    .Y(_0144_),
    .B1(_1378_));
 sg13g2_o21ai_1 _4211_ (.B1(net1254),
    .Y(_1379_),
    .A1(net400),
    .A2(net991));
 sg13g2_a21oi_1 _4212_ (.A1(net1140),
    .A2(net991),
    .Y(_0145_),
    .B1(_1379_));
 sg13g2_o21ai_1 _4213_ (.B1(net1254),
    .Y(_1380_),
    .A1(net391),
    .A2(net990));
 sg13g2_a21oi_1 _4214_ (.A1(net1142),
    .A2(net990),
    .Y(_0146_),
    .B1(_1380_));
 sg13g2_o21ai_1 _4215_ (.B1(net1254),
    .Y(_1381_),
    .A1(net395),
    .A2(net990));
 sg13g2_a21oi_1 _4216_ (.A1(net1144),
    .A2(net990),
    .Y(_0147_),
    .B1(_1381_));
 sg13g2_and2_1 _4217_ (.A(_0569_),
    .B(_1339_),
    .X(_1382_));
 sg13g2_o21ai_1 _4218_ (.B1(net1249),
    .Y(_1383_),
    .A1(net371),
    .A2(net989));
 sg13g2_a21oi_1 _4219_ (.A1(net1229),
    .A2(net989),
    .Y(_0148_),
    .B1(_1383_));
 sg13g2_o21ai_1 _4220_ (.B1(net1249),
    .Y(_1384_),
    .A1(net437),
    .A2(net988));
 sg13g2_a21oi_1 _4221_ (.A1(net1125),
    .A2(net988),
    .Y(_0149_),
    .B1(_1384_));
 sg13g2_o21ai_1 _4222_ (.B1(net1249),
    .Y(_1385_),
    .A1(net424),
    .A2(net988));
 sg13g2_a21oi_1 _4223_ (.A1(net1130),
    .A2(net988),
    .Y(_0150_),
    .B1(_1385_));
 sg13g2_o21ai_1 _4224_ (.B1(net1249),
    .Y(_1386_),
    .A1(net416),
    .A2(net989));
 sg13g2_a21oi_1 _4225_ (.A1(net1134),
    .A2(net989),
    .Y(_0151_),
    .B1(_1386_));
 sg13g2_o21ai_1 _4226_ (.B1(net1249),
    .Y(_1387_),
    .A1(net352),
    .A2(net989));
 sg13g2_a21oi_1 _4227_ (.A1(net1139),
    .A2(net989),
    .Y(_0152_),
    .B1(_1387_));
 sg13g2_o21ai_1 _4228_ (.B1(net1249),
    .Y(_1388_),
    .A1(net446),
    .A2(net988));
 sg13g2_a21oi_1 _4229_ (.A1(net1140),
    .A2(net988),
    .Y(_0153_),
    .B1(_1388_));
 sg13g2_o21ai_1 _4230_ (.B1(net1249),
    .Y(_1389_),
    .A1(net417),
    .A2(net988));
 sg13g2_a21oi_1 _4231_ (.A1(net1143),
    .A2(net988),
    .Y(_0154_),
    .B1(_1389_));
 sg13g2_o21ai_1 _4232_ (.B1(net1249),
    .Y(_1390_),
    .A1(net389),
    .A2(net989));
 sg13g2_a21oi_1 _4233_ (.A1(net1145),
    .A2(net989),
    .Y(_0155_),
    .B1(_1390_));
 sg13g2_nor2_2 _4234_ (.A(_0074_),
    .B(_1349_),
    .Y(_1391_));
 sg13g2_and2_1 _4235_ (.A(_1339_),
    .B(_1391_),
    .X(_1392_));
 sg13g2_o21ai_1 _4236_ (.B1(net1244),
    .Y(_1393_),
    .A1(net349),
    .A2(net987));
 sg13g2_a21oi_1 _4237_ (.A1(net1229),
    .A2(net987),
    .Y(_0156_),
    .B1(_1393_));
 sg13g2_o21ai_1 _4238_ (.B1(net1244),
    .Y(_1394_),
    .A1(net372),
    .A2(net987));
 sg13g2_a21oi_1 _4239_ (.A1(net1125),
    .A2(net987),
    .Y(_0157_),
    .B1(_1394_));
 sg13g2_o21ai_1 _4240_ (.B1(net1244),
    .Y(_1395_),
    .A1(net428),
    .A2(net986));
 sg13g2_a21oi_1 _4241_ (.A1(net1130),
    .A2(net986),
    .Y(_0158_),
    .B1(_1395_));
 sg13g2_o21ai_1 _4242_ (.B1(net1244),
    .Y(_1396_),
    .A1(net415),
    .A2(net986));
 sg13g2_a21oi_1 _4243_ (.A1(net1134),
    .A2(net986),
    .Y(_0159_),
    .B1(_1396_));
 sg13g2_o21ai_1 _4244_ (.B1(net1244),
    .Y(_1397_),
    .A1(net381),
    .A2(net987));
 sg13g2_a21oi_1 _4245_ (.A1(net1138),
    .A2(net987),
    .Y(_0160_),
    .B1(_1397_));
 sg13g2_o21ai_1 _4246_ (.B1(net1244),
    .Y(_1398_),
    .A1(net399),
    .A2(net986));
 sg13g2_a21oi_1 _4247_ (.A1(net1140),
    .A2(net986),
    .Y(_0161_),
    .B1(_1398_));
 sg13g2_o21ai_1 _4248_ (.B1(net1244),
    .Y(_1399_),
    .A1(net434),
    .A2(net986));
 sg13g2_a21oi_1 _4249_ (.A1(net1142),
    .A2(net986),
    .Y(_0162_),
    .B1(_1399_));
 sg13g2_o21ai_1 _4250_ (.B1(net1244),
    .Y(_1400_),
    .A1(net387),
    .A2(net987));
 sg13g2_a21oi_1 _4251_ (.A1(net1144),
    .A2(net987),
    .Y(_0163_),
    .B1(_1400_));
 sg13g2_nor2_2 _4252_ (.A(_0074_),
    .B(_1360_),
    .Y(_1401_));
 sg13g2_and2_1 _4253_ (.A(_1339_),
    .B(_1401_),
    .X(_1402_));
 sg13g2_o21ai_1 _4254_ (.B1(net1248),
    .Y(_1403_),
    .A1(net364),
    .A2(net985));
 sg13g2_a21oi_1 _4255_ (.A1(net1229),
    .A2(net985),
    .Y(_0164_),
    .B1(_1403_));
 sg13g2_o21ai_1 _4256_ (.B1(net1246),
    .Y(_1404_),
    .A1(net423),
    .A2(net984));
 sg13g2_a21oi_1 _4257_ (.A1(net1125),
    .A2(net985),
    .Y(_0165_),
    .B1(_1404_));
 sg13g2_o21ai_1 _4258_ (.B1(net1248),
    .Y(_1405_),
    .A1(net402),
    .A2(net985));
 sg13g2_a21oi_1 _4259_ (.A1(net1130),
    .A2(net985),
    .Y(_0166_),
    .B1(_1405_));
 sg13g2_o21ai_1 _4260_ (.B1(net1246),
    .Y(_1406_),
    .A1(net450),
    .A2(_1402_));
 sg13g2_a21oi_1 _4261_ (.A1(net1134),
    .A2(net984),
    .Y(_0167_),
    .B1(_1406_));
 sg13g2_o21ai_1 _4262_ (.B1(net1246),
    .Y(_1407_),
    .A1(net382),
    .A2(net984));
 sg13g2_a21oi_1 _4263_ (.A1(net1139),
    .A2(net985),
    .Y(_0168_),
    .B1(_1407_));
 sg13g2_o21ai_1 _4264_ (.B1(net1246),
    .Y(_1408_),
    .A1(net447),
    .A2(net985));
 sg13g2_a21oi_1 _4265_ (.A1(net1140),
    .A2(net984),
    .Y(_0169_),
    .B1(_1408_));
 sg13g2_o21ai_1 _4266_ (.B1(net1246),
    .Y(_1409_),
    .A1(net420),
    .A2(net984));
 sg13g2_a21oi_1 _4267_ (.A1(net1143),
    .A2(net984),
    .Y(_0170_),
    .B1(_1409_));
 sg13g2_o21ai_1 _4268_ (.B1(net1246),
    .Y(_1410_),
    .A1(net356),
    .A2(net984));
 sg13g2_a21oi_1 _4269_ (.A1(net1145),
    .A2(net984),
    .Y(_0171_),
    .B1(_1410_));
 sg13g2_nor2_2 _4270_ (.A(_0074_),
    .B(_1371_),
    .Y(_1411_));
 sg13g2_and2_1 _4271_ (.A(_1339_),
    .B(_1411_),
    .X(_1412_));
 sg13g2_o21ai_1 _4272_ (.B1(net1243),
    .Y(_1413_),
    .A1(net375),
    .A2(net983));
 sg13g2_a21oi_1 _4273_ (.A1(net1228),
    .A2(net983),
    .Y(_0172_),
    .B1(_1413_));
 sg13g2_o21ai_1 _4274_ (.B1(net1243),
    .Y(_1414_),
    .A1(net449),
    .A2(net981));
 sg13g2_a21oi_1 _4275_ (.A1(net1125),
    .A2(net981),
    .Y(_0173_),
    .B1(_1414_));
 sg13g2_o21ai_1 _4276_ (.B1(net1243),
    .Y(_1415_),
    .A1(net374),
    .A2(net982));
 sg13g2_a21oi_1 _4277_ (.A1(net1130),
    .A2(net981),
    .Y(_0174_),
    .B1(_1415_));
 sg13g2_o21ai_1 _4278_ (.B1(net1243),
    .Y(_1416_),
    .A1(net418),
    .A2(net981));
 sg13g2_a21oi_1 _4279_ (.A1(net1134),
    .A2(net982),
    .Y(_0175_),
    .B1(_1416_));
 sg13g2_o21ai_1 _4280_ (.B1(net1243),
    .Y(_1417_),
    .A1(net362),
    .A2(net983));
 sg13g2_a21oi_1 _4281_ (.A1(net1138),
    .A2(net983),
    .Y(_0176_),
    .B1(_1417_));
 sg13g2_o21ai_1 _4282_ (.B1(net1243),
    .Y(_1418_),
    .A1(net336),
    .A2(net981));
 sg13g2_a21oi_1 _4283_ (.A1(net1140),
    .A2(net981),
    .Y(_0177_),
    .B1(_1418_));
 sg13g2_o21ai_1 _4284_ (.B1(net1243),
    .Y(_1419_),
    .A1(net460),
    .A2(net982));
 sg13g2_a21oi_1 _4285_ (.A1(net1142),
    .A2(net982),
    .Y(_0178_),
    .B1(_1419_));
 sg13g2_o21ai_1 _4286_ (.B1(net1243),
    .Y(_1420_),
    .A1(net350),
    .A2(net981));
 sg13g2_a21oi_1 _4287_ (.A1(net1144),
    .A2(net981),
    .Y(_0179_),
    .B1(_1420_));
 sg13g2_nor3_2 _4288_ (.A(\spi_address[4] ),
    .B(net456),
    .C(_0571_),
    .Y(_1421_));
 sg13g2_nand2_1 _4289_ (.Y(_1422_),
    .A(_1338_),
    .B(_1421_));
 sg13g2_and2_1 _4290_ (.A(\charlie_0.memory[20][4] ),
    .B(_0562_),
    .X(_1423_));
 sg13g2_nand2_1 _4291_ (.Y(_1424_),
    .A(\charlie_0.memory[20][4] ),
    .B(_0562_));
 sg13g2_nand2_1 _4292_ (.Y(_1425_),
    .A(\charlie_0.memory[8][0] ),
    .B(net1014));
 sg13g2_nand2_1 _4293_ (.Y(_1426_),
    .A(net1212),
    .B(net1020));
 sg13g2_nand3_1 _4294_ (.B(_1425_),
    .C(_1426_),
    .A(_1422_),
    .Y(_1427_));
 sg13g2_o21ai_1 _4295_ (.B1(_1427_),
    .Y(_1428_),
    .A1(net1231),
    .A2(_1422_));
 sg13g2_nor2_1 _4296_ (.A(net1223),
    .B(_1428_),
    .Y(_0180_));
 sg13g2_nand2_1 _4297_ (.Y(_1429_),
    .A(\charlie_0.memory[8][1] ),
    .B(net1013));
 sg13g2_nand2_1 _4298_ (.Y(_1430_),
    .A(net1209),
    .B(net1016));
 sg13g2_nand3_1 _4299_ (.B(_1429_),
    .C(_1430_),
    .A(net979),
    .Y(_1431_));
 sg13g2_o21ai_1 _4300_ (.B1(_1431_),
    .Y(_1432_),
    .A1(net1198),
    .A2(net979));
 sg13g2_nor2_1 _4301_ (.A(net1215),
    .B(_1432_),
    .Y(_0181_));
 sg13g2_nand2_1 _4302_ (.Y(_1433_),
    .A(\charlie_0.memory[8][2] ),
    .B(net1013));
 sg13g2_nand2_1 _4303_ (.Y(_1434_),
    .A(net1207),
    .B(net1015));
 sg13g2_nand3_1 _4304_ (.B(_1433_),
    .C(_1434_),
    .A(net980),
    .Y(_1435_));
 sg13g2_o21ai_1 _4305_ (.B1(_1435_),
    .Y(_1436_),
    .A1(net1193),
    .A2(net980));
 sg13g2_nor2_1 _4306_ (.A(net1222),
    .B(_1436_),
    .Y(_0182_));
 sg13g2_nand2_1 _4307_ (.Y(_1437_),
    .A(\charlie_0.memory[8][3] ),
    .B(net1013));
 sg13g2_nand2_1 _4308_ (.Y(_1438_),
    .A(net1205),
    .B(net1015));
 sg13g2_nand3_1 _4309_ (.B(_1437_),
    .C(_1438_),
    .A(net980),
    .Y(_1439_));
 sg13g2_o21ai_1 _4310_ (.B1(_1439_),
    .Y(_1440_),
    .A1(net1190),
    .A2(net980));
 sg13g2_nor2_1 _4311_ (.A(net1222),
    .B(_1440_),
    .Y(_0183_));
 sg13g2_nand2_1 _4312_ (.Y(_1441_),
    .A(\charlie_0.memory[8][4] ),
    .B(net1013));
 sg13g2_nand2_1 _4313_ (.Y(_1442_),
    .A(net1203),
    .B(net1015));
 sg13g2_nand3_1 _4314_ (.B(_1441_),
    .C(_1442_),
    .A(net979),
    .Y(_1443_));
 sg13g2_o21ai_1 _4315_ (.B1(_1443_),
    .Y(_1444_),
    .A1(net1188),
    .A2(net979));
 sg13g2_nor2_1 _4316_ (.A(net1222),
    .B(_1444_),
    .Y(_0184_));
 sg13g2_nand2_1 _4317_ (.Y(_1445_),
    .A(\charlie_0.memory[8][5] ),
    .B(net1013));
 sg13g2_nand2_1 _4318_ (.Y(_1446_),
    .A(net1201),
    .B(net1015));
 sg13g2_nand3_1 _4319_ (.B(_1445_),
    .C(_1446_),
    .A(net979),
    .Y(_1447_));
 sg13g2_o21ai_1 _4320_ (.B1(_1447_),
    .Y(_1448_),
    .A1(net1186),
    .A2(net979));
 sg13g2_nor2_1 _4321_ (.A(net1222),
    .B(_1448_),
    .Y(_0185_));
 sg13g2_nand2_1 _4322_ (.Y(_1449_),
    .A(\charlie_0.memory[8][6] ),
    .B(net1012));
 sg13g2_nand2_1 _4323_ (.Y(_1450_),
    .A(net355),
    .B(net1015));
 sg13g2_nand3_1 _4324_ (.B(_1449_),
    .C(_1450_),
    .A(net980),
    .Y(_1451_));
 sg13g2_o21ai_1 _4325_ (.B1(_1451_),
    .Y(_1452_),
    .A1(net1184),
    .A2(net979));
 sg13g2_nor2_1 _4326_ (.A(net1222),
    .B(_1452_),
    .Y(_0186_));
 sg13g2_nand2_1 _4327_ (.Y(_1453_),
    .A(\charlie_0.memory[8][7] ),
    .B(net1012));
 sg13g2_nand2_1 _4328_ (.Y(_1454_),
    .A(net430),
    .B(net1015));
 sg13g2_nand3_1 _4329_ (.B(_1453_),
    .C(_1454_),
    .A(net980),
    .Y(_1455_));
 sg13g2_o21ai_1 _4330_ (.B1(_1455_),
    .Y(_1456_),
    .A1(net1213),
    .A2(net979));
 sg13g2_nor2_1 _4331_ (.A(net1215),
    .B(_1456_),
    .Y(_0187_));
 sg13g2_nand3b_1 _4332_ (.B(net411),
    .C(_1350_),
    .Y(_1457_),
    .A_N(_0072_));
 sg13g2_nor2_2 _4333_ (.A(_0571_),
    .B(net412),
    .Y(_1458_));
 sg13g2_mux2_1 _4334_ (.A0(\charlie_0.memory[9][0] ),
    .A1(net333),
    .S(net1017),
    .X(_1459_));
 sg13g2_nor2_1 _4335_ (.A(_1458_),
    .B(_1459_),
    .Y(_1460_));
 sg13g2_a21oi_1 _4336_ (.A1(net1230),
    .A2(net1001),
    .Y(_1461_),
    .B1(net1219));
 sg13g2_nor2b_1 _4337_ (.A(_1460_),
    .B_N(_1461_),
    .Y(_0188_));
 sg13g2_mux2_1 _4338_ (.A0(\charlie_0.memory[9][1] ),
    .A1(\counter[9] ),
    .S(net1017),
    .X(_1462_));
 sg13g2_nor2_1 _4339_ (.A(net1000),
    .B(_1462_),
    .Y(_1463_));
 sg13g2_a21oi_1 _4340_ (.A1(net1126),
    .A2(net1000),
    .Y(_1464_),
    .B1(net1219));
 sg13g2_nor2b_1 _4341_ (.A(_1463_),
    .B_N(_1464_),
    .Y(_0189_));
 sg13g2_mux2_1 _4342_ (.A0(\charlie_0.memory[9][2] ),
    .A1(net483),
    .S(net1017),
    .X(_1465_));
 sg13g2_nor2_1 _4343_ (.A(net1000),
    .B(_1465_),
    .Y(_1466_));
 sg13g2_a21oi_1 _4344_ (.A1(net1128),
    .A2(net1000),
    .Y(_1467_),
    .B1(net1225));
 sg13g2_nor2b_1 _4345_ (.A(_1466_),
    .B_N(_1467_),
    .Y(_0190_));
 sg13g2_mux2_1 _4346_ (.A0(\charlie_0.memory[9][3] ),
    .A1(net492),
    .S(net1017),
    .X(_1468_));
 sg13g2_nor2_1 _4347_ (.A(net1000),
    .B(_1468_),
    .Y(_1469_));
 sg13g2_a21oi_1 _4348_ (.A1(net1133),
    .A2(net1000),
    .Y(_1470_),
    .B1(net1219));
 sg13g2_nor2b_1 _4349_ (.A(_1469_),
    .B_N(_1470_),
    .Y(_0191_));
 sg13g2_mux2_1 _4350_ (.A0(\charlie_0.memory[9][4] ),
    .A1(\counter[12] ),
    .S(net1017),
    .X(_1471_));
 sg13g2_nor2_1 _4351_ (.A(net1001),
    .B(_1471_),
    .Y(_1472_));
 sg13g2_a21oi_1 _4352_ (.A1(net1136),
    .A2(net1001),
    .Y(_1473_),
    .B1(net1219));
 sg13g2_nor2b_1 _4353_ (.A(_1472_),
    .B_N(_1473_),
    .Y(_0192_));
 sg13g2_mux2_1 _4354_ (.A0(\charlie_0.memory[9][5] ),
    .A1(net440),
    .S(net1017),
    .X(_1474_));
 sg13g2_nor2_1 _4355_ (.A(net1000),
    .B(_1474_),
    .Y(_1475_));
 sg13g2_a21oi_1 _4356_ (.A1(net1141),
    .A2(net1000),
    .Y(_1476_),
    .B1(net1219));
 sg13g2_nor2b_1 _4357_ (.A(_1475_),
    .B_N(_1476_),
    .Y(_0193_));
 sg13g2_nor2_1 _4358_ (.A(\charlie_0.memory[9][6] ),
    .B(net1019),
    .Y(_1477_));
 sg13g2_a21oi_1 _4359_ (.A1(_1830_),
    .A2(net1019),
    .Y(_1478_),
    .B1(_1477_));
 sg13g2_nor2_1 _4360_ (.A(net1001),
    .B(_1478_),
    .Y(_1479_));
 sg13g2_a21oi_1 _4361_ (.A1(net1143),
    .A2(net1001),
    .Y(_1480_),
    .B1(net1218));
 sg13g2_nor2b_1 _4362_ (.A(_1479_),
    .B_N(_1480_),
    .Y(_0194_));
 sg13g2_mux2_1 _4363_ (.A0(\charlie_0.memory[9][7] ),
    .A1(net419),
    .S(net1019),
    .X(_1481_));
 sg13g2_nor2_1 _4364_ (.A(net1001),
    .B(_1481_),
    .Y(_1482_));
 sg13g2_a21oi_1 _4365_ (.A1(net1145),
    .A2(net1001),
    .Y(_1483_),
    .B1(net1218));
 sg13g2_nor2b_1 _4366_ (.A(_1482_),
    .B_N(_1483_),
    .Y(_0195_));
 sg13g2_nand2_1 _4367_ (.Y(_1484_),
    .A(_1361_),
    .B(_1421_));
 sg13g2_nand2_1 _4368_ (.Y(_1485_),
    .A(net479),
    .B(net1014));
 sg13g2_nand2_1 _4369_ (.Y(_1486_),
    .A(\counter[16] ),
    .B(net1019));
 sg13g2_nand3_1 _4370_ (.B(_1485_),
    .C(_1486_),
    .A(net977),
    .Y(_1487_));
 sg13g2_o21ai_1 _4371_ (.B1(net480),
    .Y(_1488_),
    .A1(net1231),
    .A2(net977));
 sg13g2_nor2_1 _4372_ (.A(net1218),
    .B(_1488_),
    .Y(_0196_));
 sg13g2_nand2_1 _4373_ (.Y(_1489_),
    .A(net490),
    .B(net1014));
 sg13g2_nand2_1 _4374_ (.Y(_1490_),
    .A(\counter[17] ),
    .B(net1019));
 sg13g2_nand3_1 _4375_ (.B(_1489_),
    .C(_1490_),
    .A(net977),
    .Y(_1491_));
 sg13g2_o21ai_1 _4376_ (.B1(_1491_),
    .Y(_1492_),
    .A1(net1197),
    .A2(net977));
 sg13g2_nor2_1 _4377_ (.A(net1218),
    .B(_1492_),
    .Y(_0197_));
 sg13g2_nor2_1 _4378_ (.A(_1800_),
    .B(net1018),
    .Y(_1493_));
 sg13g2_a21oi_1 _4379_ (.A1(\counter[18] ),
    .A2(net1018),
    .Y(_1494_),
    .B1(_1493_));
 sg13g2_nand2_1 _4380_ (.Y(_1495_),
    .A(net978),
    .B(_1494_));
 sg13g2_o21ai_1 _4381_ (.B1(_1495_),
    .Y(_1496_),
    .A1(net1194),
    .A2(net978));
 sg13g2_nor2_1 _4382_ (.A(net1220),
    .B(_1496_),
    .Y(_0198_));
 sg13g2_nor2_1 _4383_ (.A(_1799_),
    .B(net1018),
    .Y(_1497_));
 sg13g2_a21oi_1 _4384_ (.A1(\counter[19] ),
    .A2(net1018),
    .Y(_1498_),
    .B1(_1497_));
 sg13g2_nand2_1 _4385_ (.Y(_1499_),
    .A(net978),
    .B(_1498_));
 sg13g2_o21ai_1 _4386_ (.B1(_1499_),
    .Y(_1500_),
    .A1(net1191),
    .A2(net978));
 sg13g2_nor2_1 _4387_ (.A(net1220),
    .B(_1500_),
    .Y(_0199_));
 sg13g2_nand2_1 _4388_ (.Y(_1501_),
    .A(\charlie_0.memory[10][4] ),
    .B(net1014));
 sg13g2_nand2_1 _4389_ (.Y(_1502_),
    .A(net470),
    .B(net1019));
 sg13g2_nand3_1 _4390_ (.B(_1501_),
    .C(_1502_),
    .A(net977),
    .Y(_1503_));
 sg13g2_o21ai_1 _4391_ (.B1(_1503_),
    .Y(_1504_),
    .A1(net1189),
    .A2(net977));
 sg13g2_nor2_1 _4392_ (.A(net1220),
    .B(_1504_),
    .Y(_0200_));
 sg13g2_nor2_1 _4393_ (.A(_1798_),
    .B(net1020),
    .Y(_1505_));
 sg13g2_a21oi_1 _4394_ (.A1(\counter[21] ),
    .A2(net1020),
    .Y(_1506_),
    .B1(_1505_));
 sg13g2_nand2_1 _4395_ (.Y(_1507_),
    .A(_1484_),
    .B(_1506_));
 sg13g2_o21ai_1 _4396_ (.B1(_1507_),
    .Y(_1508_),
    .A1(net1187),
    .A2(net978));
 sg13g2_nor2_1 _4397_ (.A(net1221),
    .B(_1508_),
    .Y(_0201_));
 sg13g2_nor2_1 _4398_ (.A(_1797_),
    .B(net1017),
    .Y(_1509_));
 sg13g2_a21oi_1 _4399_ (.A1(\counter[22] ),
    .A2(net1017),
    .Y(_1510_),
    .B1(_1509_));
 sg13g2_nand2_1 _4400_ (.Y(_1511_),
    .A(net978),
    .B(_1510_));
 sg13g2_o21ai_1 _4401_ (.B1(_1511_),
    .Y(_1512_),
    .A1(net1185),
    .A2(net978));
 sg13g2_nor2_1 _4402_ (.A(net1221),
    .B(_1512_),
    .Y(_0202_));
 sg13g2_nand2_1 _4403_ (.Y(_1513_),
    .A(net444),
    .B(net1014));
 sg13g2_nand2_1 _4404_ (.Y(_1514_),
    .A(\counter[23] ),
    .B(net1019));
 sg13g2_nand3_1 _4405_ (.B(_1513_),
    .C(_1514_),
    .A(net977),
    .Y(_1515_));
 sg13g2_o21ai_1 _4406_ (.B1(net445),
    .Y(_1516_),
    .A1(net1214),
    .A2(net977));
 sg13g2_nor2_1 _4407_ (.A(net1221),
    .B(_1516_),
    .Y(_0203_));
 sg13g2_nand2_1 _4408_ (.Y(_1517_),
    .A(_1372_),
    .B(_1421_));
 sg13g2_nand2_1 _4409_ (.Y(_1518_),
    .A(\charlie_0.memory[11][0] ),
    .B(net1014));
 sg13g2_nand2_1 _4410_ (.Y(_1519_),
    .A(net495),
    .B(net1016));
 sg13g2_nand3_1 _4411_ (.B(_1518_),
    .C(_1519_),
    .A(net976),
    .Y(_1520_));
 sg13g2_o21ai_1 _4412_ (.B1(_1520_),
    .Y(_1521_),
    .A1(net1231),
    .A2(net976));
 sg13g2_nor2_1 _4413_ (.A(net1217),
    .B(_1521_),
    .Y(_0204_));
 sg13g2_nand2_1 _4414_ (.Y(_1522_),
    .A(\charlie_0.memory[11][1] ),
    .B(net1012));
 sg13g2_nand2_1 _4415_ (.Y(_1523_),
    .A(net353),
    .B(net1016));
 sg13g2_nand3_1 _4416_ (.B(_1522_),
    .C(_1523_),
    .A(net974),
    .Y(_1524_));
 sg13g2_o21ai_1 _4417_ (.B1(_1524_),
    .Y(_1525_),
    .A1(net1197),
    .A2(net974));
 sg13g2_nor2_1 _4418_ (.A(net1217),
    .B(_1525_),
    .Y(_0205_));
 sg13g2_nand2_1 _4419_ (.Y(_1526_),
    .A(\charlie_0.memory[11][2] ),
    .B(net1012));
 sg13g2_nand2_1 _4420_ (.Y(_1527_),
    .A(\counter[26] ),
    .B(net1016));
 sg13g2_nand3_1 _4421_ (.B(_1526_),
    .C(_1527_),
    .A(net974),
    .Y(_1528_));
 sg13g2_o21ai_1 _4422_ (.B1(_1528_),
    .Y(_1529_),
    .A1(net1194),
    .A2(net974));
 sg13g2_nor2_1 _4423_ (.A(net1215),
    .B(_1529_),
    .Y(_0206_));
 sg13g2_nand2_1 _4424_ (.Y(_1530_),
    .A(\charlie_0.memory[11][3] ),
    .B(net1012));
 sg13g2_nand2_1 _4425_ (.Y(_1531_),
    .A(net396),
    .B(net1016));
 sg13g2_nand3_1 _4426_ (.B(_1530_),
    .C(_1531_),
    .A(net976),
    .Y(_1532_));
 sg13g2_o21ai_1 _4427_ (.B1(_1532_),
    .Y(_1533_),
    .A1(net1191),
    .A2(net976));
 sg13g2_nor2_1 _4428_ (.A(net1216),
    .B(_1533_),
    .Y(_0207_));
 sg13g2_nand2_1 _4429_ (.Y(_1534_),
    .A(\charlie_0.memory[11][4] ),
    .B(net1012));
 sg13g2_nand2_1 _4430_ (.Y(_1535_),
    .A(net406),
    .B(net1016));
 sg13g2_nand3_1 _4431_ (.B(_1534_),
    .C(_1535_),
    .A(net974),
    .Y(_1536_));
 sg13g2_o21ai_1 _4432_ (.B1(_1536_),
    .Y(_1537_),
    .A1(net1189),
    .A2(net974));
 sg13g2_nor2_1 _4433_ (.A(net1215),
    .B(_1537_),
    .Y(_0208_));
 sg13g2_nand2_1 _4434_ (.Y(_1538_),
    .A(\charlie_0.memory[11][5] ),
    .B(net1012));
 sg13g2_nand2_1 _4435_ (.Y(_1539_),
    .A(net369),
    .B(net1016));
 sg13g2_nand3_1 _4436_ (.B(_1538_),
    .C(_1539_),
    .A(net975),
    .Y(_1540_));
 sg13g2_o21ai_1 _4437_ (.B1(_1540_),
    .Y(_1541_),
    .A1(net1186),
    .A2(net975));
 sg13g2_nor2_1 _4438_ (.A(net1215),
    .B(_1541_),
    .Y(_0209_));
 sg13g2_nand2_1 _4439_ (.Y(_1542_),
    .A(\charlie_0.memory[11][6] ),
    .B(net1012));
 sg13g2_nand2_1 _4440_ (.Y(_1543_),
    .A(net478),
    .B(net1015));
 sg13g2_nand3_1 _4441_ (.B(_1542_),
    .C(_1543_),
    .A(net975),
    .Y(_1544_));
 sg13g2_o21ai_1 _4442_ (.B1(_1544_),
    .Y(_1545_),
    .A1(net1184),
    .A2(net975));
 sg13g2_nor2_1 _4443_ (.A(net1215),
    .B(_1545_),
    .Y(_0210_));
 sg13g2_nand2_1 _4444_ (.Y(_1546_),
    .A(\charlie_0.memory[11][7] ),
    .B(net1013));
 sg13g2_nand2_1 _4445_ (.Y(_1547_),
    .A(\counter[31] ),
    .B(net1015));
 sg13g2_nand3_1 _4446_ (.B(_1546_),
    .C(_1547_),
    .A(net974),
    .Y(_1548_));
 sg13g2_o21ai_1 _4447_ (.B1(_1548_),
    .Y(_1549_),
    .A1(net1213),
    .A2(net974));
 sg13g2_nor2_1 _4448_ (.A(net1216),
    .B(_1549_),
    .Y(_0211_));
 sg13g2_nand2_1 _4449_ (.Y(_1550_),
    .A(_0569_),
    .B(_1421_));
 sg13g2_and2_2 _4450_ (.A(\charlie_0.memory[20][5] ),
    .B(_0563_),
    .X(_1551_));
 sg13g2_nand2_2 _4451_ (.Y(_1552_),
    .A(\charlie_0.memory[20][5] ),
    .B(_0563_));
 sg13g2_nand2_1 _4452_ (.Y(_1553_),
    .A(\charlie_0.memory[12][0] ),
    .B(net1004));
 sg13g2_nand2_1 _4453_ (.Y(_1554_),
    .A(net1212),
    .B(net1007));
 sg13g2_nand3_1 _4454_ (.B(_1553_),
    .C(_1554_),
    .A(net973),
    .Y(_1555_));
 sg13g2_o21ai_1 _4455_ (.B1(_1555_),
    .Y(_1556_),
    .A1(net1231),
    .A2(net973));
 sg13g2_nor2_1 _4456_ (.A(net1216),
    .B(_1556_),
    .Y(_0212_));
 sg13g2_nand2_1 _4457_ (.Y(_1557_),
    .A(\charlie_0.memory[12][1] ),
    .B(_1552_));
 sg13g2_nand2_1 _4458_ (.Y(_1558_),
    .A(net1209),
    .B(_1551_));
 sg13g2_nand3_1 _4459_ (.B(_1557_),
    .C(_1558_),
    .A(net973),
    .Y(_1559_));
 sg13g2_o21ai_1 _4460_ (.B1(_1559_),
    .Y(_1560_),
    .A1(net1198),
    .A2(net972));
 sg13g2_nor2_1 _4461_ (.A(net1216),
    .B(_1560_),
    .Y(_0213_));
 sg13g2_nand2_1 _4462_ (.Y(_1561_),
    .A(\charlie_0.memory[12][2] ),
    .B(net1003));
 sg13g2_nand2_1 _4463_ (.Y(_1562_),
    .A(net1207),
    .B(net1007));
 sg13g2_nand3_1 _4464_ (.B(_1561_),
    .C(_1562_),
    .A(net972),
    .Y(_1563_));
 sg13g2_o21ai_1 _4465_ (.B1(_1563_),
    .Y(_1564_),
    .A1(net1193),
    .A2(net972));
 sg13g2_nor2_1 _4466_ (.A(net1222),
    .B(_1564_),
    .Y(_0214_));
 sg13g2_nand2_1 _4467_ (.Y(_1565_),
    .A(\charlie_0.memory[12][3] ),
    .B(net1003));
 sg13g2_nand2_1 _4468_ (.Y(_1566_),
    .A(net1206),
    .B(net1007));
 sg13g2_nand3_1 _4469_ (.B(_1565_),
    .C(_1566_),
    .A(net973),
    .Y(_1567_));
 sg13g2_o21ai_1 _4470_ (.B1(_1567_),
    .Y(_1568_),
    .A1(net1190),
    .A2(net973));
 sg13g2_nor2_1 _4471_ (.A(net1223),
    .B(_1568_),
    .Y(_0215_));
 sg13g2_nand2_1 _4472_ (.Y(_1569_),
    .A(\charlie_0.memory[12][4] ),
    .B(net1003));
 sg13g2_nand2_1 _4473_ (.Y(_1570_),
    .A(net1203),
    .B(net1007));
 sg13g2_nand3_1 _4474_ (.B(_1569_),
    .C(_1570_),
    .A(net972),
    .Y(_1571_));
 sg13g2_o21ai_1 _4475_ (.B1(_1571_),
    .Y(_1572_),
    .A1(net1188),
    .A2(net972));
 sg13g2_nor2_1 _4476_ (.A(net1222),
    .B(_1572_),
    .Y(_0216_));
 sg13g2_nand2_1 _4477_ (.Y(_1573_),
    .A(\charlie_0.memory[12][5] ),
    .B(net1003));
 sg13g2_nand2_1 _4478_ (.Y(_1574_),
    .A(net1201),
    .B(net1007));
 sg13g2_nand3_1 _4479_ (.B(_1573_),
    .C(_1574_),
    .A(net973),
    .Y(_1575_));
 sg13g2_o21ai_1 _4480_ (.B1(_1575_),
    .Y(_1576_),
    .A1(net1186),
    .A2(net973));
 sg13g2_nor2_1 _4481_ (.A(net1216),
    .B(_1576_),
    .Y(_0217_));
 sg13g2_nand2_1 _4482_ (.Y(_1577_),
    .A(\charlie_0.memory[12][6] ),
    .B(net1003));
 sg13g2_nand2_1 _4483_ (.Y(_1578_),
    .A(net355),
    .B(net1007));
 sg13g2_nand3_1 _4484_ (.B(_1577_),
    .C(_1578_),
    .A(net972),
    .Y(_1579_));
 sg13g2_o21ai_1 _4485_ (.B1(_1579_),
    .Y(_1580_),
    .A1(net1184),
    .A2(net972));
 sg13g2_nor2_1 _4486_ (.A(net1215),
    .B(_1580_),
    .Y(_0218_));
 sg13g2_nand2_1 _4487_ (.Y(_1581_),
    .A(\charlie_0.memory[12][7] ),
    .B(net1003));
 sg13g2_nand2_1 _4488_ (.Y(_1582_),
    .A(net464),
    .B(net1007));
 sg13g2_nand3_1 _4489_ (.B(_1581_),
    .C(_1582_),
    .A(net973),
    .Y(_1583_));
 sg13g2_o21ai_1 _4490_ (.B1(_1583_),
    .Y(_1584_),
    .A1(net1213),
    .A2(net972));
 sg13g2_nor2_1 _4491_ (.A(net1216),
    .B(_1584_),
    .Y(_0219_));
 sg13g2_nand2_1 _4492_ (.Y(_1585_),
    .A(_1391_),
    .B(_1421_));
 sg13g2_nand2_1 _4493_ (.Y(_1586_),
    .A(\charlie_0.memory[13][0] ),
    .B(net1005));
 sg13g2_nand2_1 _4494_ (.Y(_1587_),
    .A(net333),
    .B(net1009));
 sg13g2_nand3_1 _4495_ (.B(_1586_),
    .C(_1587_),
    .A(net970),
    .Y(_1588_));
 sg13g2_o21ai_1 _4496_ (.B1(_1588_),
    .Y(_1589_),
    .A1(net1233),
    .A2(net970));
 sg13g2_nor2_1 _4497_ (.A(net1225),
    .B(_1589_),
    .Y(_0220_));
 sg13g2_nand2_1 _4498_ (.Y(_1590_),
    .A(\charlie_0.memory[13][1] ),
    .B(net1005));
 sg13g2_nand2_1 _4499_ (.Y(_1591_),
    .A(\counter[9] ),
    .B(net1009));
 sg13g2_nand3_1 _4500_ (.B(_1590_),
    .C(_1591_),
    .A(_1585_),
    .Y(_1592_));
 sg13g2_o21ai_1 _4501_ (.B1(_1592_),
    .Y(_1593_),
    .A1(net1199),
    .A2(net971));
 sg13g2_nor2_1 _4502_ (.A(net1225),
    .B(_1593_),
    .Y(_0221_));
 sg13g2_nand2_1 _4503_ (.Y(_1594_),
    .A(\charlie_0.memory[13][2] ),
    .B(net1005));
 sg13g2_nand2_1 _4504_ (.Y(_1595_),
    .A(\counter[10] ),
    .B(net1009));
 sg13g2_nand3_1 _4505_ (.B(_1594_),
    .C(net484),
    .A(net971),
    .Y(_1596_));
 sg13g2_o21ai_1 _4506_ (.B1(_1596_),
    .Y(_1597_),
    .A1(net1195),
    .A2(net970));
 sg13g2_nor2_1 _4507_ (.A(net1225),
    .B(_1597_),
    .Y(_0222_));
 sg13g2_nand2_1 _4508_ (.Y(_1598_),
    .A(\charlie_0.memory[13][3] ),
    .B(net1005));
 sg13g2_nand2_1 _4509_ (.Y(_1599_),
    .A(net486),
    .B(net1009));
 sg13g2_nand3_1 _4510_ (.B(_1598_),
    .C(_1599_),
    .A(net970),
    .Y(_1600_));
 sg13g2_o21ai_1 _4511_ (.B1(_1600_),
    .Y(_1601_),
    .A1(net1191),
    .A2(net970));
 sg13g2_nor2_1 _4512_ (.A(net1225),
    .B(_1601_),
    .Y(_0223_));
 sg13g2_nand2_1 _4513_ (.Y(_1602_),
    .A(\charlie_0.memory[13][4] ),
    .B(net1005));
 sg13g2_nand2_1 _4514_ (.Y(_1603_),
    .A(\counter[12] ),
    .B(net1009));
 sg13g2_nand3_1 _4515_ (.B(_1602_),
    .C(net477),
    .A(net971),
    .Y(_1604_));
 sg13g2_o21ai_1 _4516_ (.B1(_1604_),
    .Y(_1605_),
    .A1(net1189),
    .A2(net970));
 sg13g2_nor2_1 _4517_ (.A(net1219),
    .B(_1605_),
    .Y(_0224_));
 sg13g2_nand2_1 _4518_ (.Y(_1606_),
    .A(\charlie_0.memory[13][5] ),
    .B(net1006));
 sg13g2_nand2_1 _4519_ (.Y(_1607_),
    .A(net440),
    .B(net1009));
 sg13g2_nand3_1 _4520_ (.B(_1606_),
    .C(_1607_),
    .A(net970),
    .Y(_1608_));
 sg13g2_o21ai_1 _4521_ (.B1(_1608_),
    .Y(_1609_),
    .A1(net1187),
    .A2(net970));
 sg13g2_nor2_1 _4522_ (.A(net1219),
    .B(_1609_),
    .Y(_0225_));
 sg13g2_nand2_1 _4523_ (.Y(_1610_),
    .A(\charlie_0.memory[13][6] ),
    .B(net1006));
 sg13g2_nand2_1 _4524_ (.Y(_1611_),
    .A(net360),
    .B(net1011));
 sg13g2_nand3_1 _4525_ (.B(_1610_),
    .C(_1611_),
    .A(net971),
    .Y(_1612_));
 sg13g2_o21ai_1 _4526_ (.B1(_1612_),
    .Y(_1613_),
    .A1(net1185),
    .A2(net971));
 sg13g2_nor2_1 _4527_ (.A(net1218),
    .B(_1613_),
    .Y(_0226_));
 sg13g2_nand2_1 _4528_ (.Y(_1614_),
    .A(\charlie_0.memory[13][7] ),
    .B(net1006));
 sg13g2_nand2_1 _4529_ (.Y(_1615_),
    .A(net419),
    .B(net1011));
 sg13g2_nand3_1 _4530_ (.B(_1614_),
    .C(_1615_),
    .A(net971),
    .Y(_1616_));
 sg13g2_o21ai_1 _4531_ (.B1(_1616_),
    .Y(_1617_),
    .A1(net1214),
    .A2(net971));
 sg13g2_nor2_1 _4532_ (.A(net1218),
    .B(_1617_),
    .Y(_0227_));
 sg13g2_nand2_1 _4533_ (.Y(_1618_),
    .A(_1401_),
    .B(_1421_));
 sg13g2_nand2_1 _4534_ (.Y(_1619_),
    .A(\charlie_0.memory[14][0] ),
    .B(net1005));
 sg13g2_nand2_1 _4535_ (.Y(_1620_),
    .A(net494),
    .B(net1011));
 sg13g2_nand3_1 _4536_ (.B(_1619_),
    .C(_1620_),
    .A(net968),
    .Y(_1621_));
 sg13g2_o21ai_1 _4537_ (.B1(_1621_),
    .Y(_1622_),
    .A1(net1232),
    .A2(net968));
 sg13g2_nor2_1 _4538_ (.A(net1219),
    .B(_1622_),
    .Y(_0228_));
 sg13g2_nand2_1 _4539_ (.Y(_1623_),
    .A(\charlie_0.memory[14][1] ),
    .B(net1005));
 sg13g2_nand2_1 _4540_ (.Y(_1624_),
    .A(\counter[17] ),
    .B(net1009));
 sg13g2_nand3_1 _4541_ (.B(_1623_),
    .C(_1624_),
    .A(net969),
    .Y(_1625_));
 sg13g2_o21ai_1 _4542_ (.B1(_1625_),
    .Y(_1626_),
    .A1(net1199),
    .A2(net969));
 sg13g2_nor2_1 _4543_ (.A(net1225),
    .B(_1626_),
    .Y(_0229_));
 sg13g2_nand2_1 _4544_ (.Y(_1627_),
    .A(\charlie_0.memory[14][2] ),
    .B(net1005));
 sg13g2_nand2_1 _4545_ (.Y(_1628_),
    .A(\counter[18] ),
    .B(net1010));
 sg13g2_nand3_1 _4546_ (.B(_1627_),
    .C(_1628_),
    .A(net969),
    .Y(_1629_));
 sg13g2_o21ai_1 _4547_ (.B1(_1629_),
    .Y(_1630_),
    .A1(net1195),
    .A2(net969));
 sg13g2_nor2_1 _4548_ (.A(net1225),
    .B(_1630_),
    .Y(_0230_));
 sg13g2_nand2_1 _4549_ (.Y(_1631_),
    .A(\charlie_0.memory[14][3] ),
    .B(net1006));
 sg13g2_nand2_1 _4550_ (.Y(_1632_),
    .A(\counter[19] ),
    .B(net1009));
 sg13g2_nand3_1 _4551_ (.B(_1631_),
    .C(_1632_),
    .A(net969),
    .Y(_1633_));
 sg13g2_o21ai_1 _4552_ (.B1(_1633_),
    .Y(_1634_),
    .A1(net1191),
    .A2(net969));
 sg13g2_nor2_1 _4553_ (.A(net1225),
    .B(_1634_),
    .Y(_0231_));
 sg13g2_nand2_1 _4554_ (.Y(_1635_),
    .A(\charlie_0.memory[14][4] ),
    .B(net1006));
 sg13g2_nand2_1 _4555_ (.Y(_1636_),
    .A(net470),
    .B(net1011));
 sg13g2_nand3_1 _4556_ (.B(_1635_),
    .C(_1636_),
    .A(net968),
    .Y(_1637_));
 sg13g2_o21ai_1 _4557_ (.B1(net471),
    .Y(_1638_),
    .A1(net1189),
    .A2(net968));
 sg13g2_nor2_1 _4558_ (.A(net1218),
    .B(_1638_),
    .Y(_0232_));
 sg13g2_nor2_1 _4559_ (.A(_1794_),
    .B(net1010),
    .Y(_1639_));
 sg13g2_a21oi_1 _4560_ (.A1(\counter[21] ),
    .A2(net1010),
    .Y(_1640_),
    .B1(_1639_));
 sg13g2_nand2_1 _4561_ (.Y(_1641_),
    .A(net969),
    .B(_1640_));
 sg13g2_o21ai_1 _4562_ (.B1(_1641_),
    .Y(_1642_),
    .A1(net1187),
    .A2(net969));
 sg13g2_nor2_1 _4563_ (.A(net1226),
    .B(_1642_),
    .Y(_0233_));
 sg13g2_nor2_1 _4564_ (.A(_1793_),
    .B(net1010),
    .Y(_1643_));
 sg13g2_a21oi_1 _4565_ (.A1(\counter[22] ),
    .A2(net1010),
    .Y(_1644_),
    .B1(_1643_));
 sg13g2_nand2_1 _4566_ (.Y(_1645_),
    .A(net968),
    .B(_1644_));
 sg13g2_o21ai_1 _4567_ (.B1(_1645_),
    .Y(_1646_),
    .A1(net1185),
    .A2(net968));
 sg13g2_nor2_1 _4568_ (.A(net1218),
    .B(_1646_),
    .Y(_0234_));
 sg13g2_nor2_1 _4569_ (.A(_1792_),
    .B(net1010),
    .Y(_1647_));
 sg13g2_a21oi_1 _4570_ (.A1(net379),
    .A2(net1010),
    .Y(_1648_),
    .B1(_1647_));
 sg13g2_nand2_1 _4571_ (.Y(_1649_),
    .A(net968),
    .B(_1648_));
 sg13g2_o21ai_1 _4572_ (.B1(_1649_),
    .Y(_1650_),
    .A1(net1214),
    .A2(net968));
 sg13g2_nor2_1 _4573_ (.A(net1221),
    .B(_1650_),
    .Y(_0235_));
 sg13g2_nand2_1 _4574_ (.Y(_1651_),
    .A(_1411_),
    .B(_1421_));
 sg13g2_nand2_1 _4575_ (.Y(_1652_),
    .A(\charlie_0.memory[15][0] ),
    .B(net1004));
 sg13g2_nand2_1 _4576_ (.Y(_1653_),
    .A(net487),
    .B(net1008));
 sg13g2_nand3_1 _4577_ (.B(_1652_),
    .C(_1653_),
    .A(net967),
    .Y(_1654_));
 sg13g2_o21ai_1 _4578_ (.B1(_1654_),
    .Y(_1655_),
    .A1(net1231),
    .A2(net967));
 sg13g2_nor2_1 _4579_ (.A(net1217),
    .B(_1655_),
    .Y(_0236_));
 sg13g2_nand2_1 _4580_ (.Y(_1656_),
    .A(\charlie_0.memory[15][1] ),
    .B(net1004));
 sg13g2_nand2_1 _4581_ (.Y(_1657_),
    .A(net353),
    .B(net1008));
 sg13g2_nand3_1 _4582_ (.B(_1656_),
    .C(_1657_),
    .A(net966),
    .Y(_1658_));
 sg13g2_o21ai_1 _4583_ (.B1(_1658_),
    .Y(_1659_),
    .A1(net1197),
    .A2(net966));
 sg13g2_nor2_1 _4584_ (.A(net1217),
    .B(_1659_),
    .Y(_0237_));
 sg13g2_nand2_1 _4585_ (.Y(_1660_),
    .A(\charlie_0.memory[15][2] ),
    .B(net1004));
 sg13g2_nand2_1 _4586_ (.Y(_1661_),
    .A(\counter[26] ),
    .B(net1008));
 sg13g2_nand3_1 _4587_ (.B(_1660_),
    .C(_1661_),
    .A(net966),
    .Y(_1662_));
 sg13g2_o21ai_1 _4588_ (.B1(_1662_),
    .Y(_1663_),
    .A1(net1194),
    .A2(net966));
 sg13g2_nor2_1 _4589_ (.A(net1217),
    .B(_1663_),
    .Y(_0238_));
 sg13g2_nand2_1 _4590_ (.Y(_1664_),
    .A(net489),
    .B(net1004));
 sg13g2_nand2_1 _4591_ (.Y(_1665_),
    .A(net396),
    .B(net1008));
 sg13g2_nand3_1 _4592_ (.B(_1664_),
    .C(_1665_),
    .A(_1651_),
    .Y(_1666_));
 sg13g2_o21ai_1 _4593_ (.B1(_1666_),
    .Y(_1667_),
    .A1(net1191),
    .A2(net967));
 sg13g2_nor2_1 _4594_ (.A(net1217),
    .B(_1667_),
    .Y(_0239_));
 sg13g2_nand2_1 _4595_ (.Y(_1668_),
    .A(\charlie_0.memory[15][4] ),
    .B(net1004));
 sg13g2_nand2_1 _4596_ (.Y(_1669_),
    .A(net406),
    .B(net1008));
 sg13g2_nand3_1 _4597_ (.B(_1668_),
    .C(_1669_),
    .A(net966),
    .Y(_1670_));
 sg13g2_o21ai_1 _4598_ (.B1(_1670_),
    .Y(_1671_),
    .A1(net1189),
    .A2(net966));
 sg13g2_nor2_1 _4599_ (.A(net1217),
    .B(_1671_),
    .Y(_0240_));
 sg13g2_nand2_1 _4600_ (.Y(_1672_),
    .A(\charlie_0.memory[15][5] ),
    .B(net1004));
 sg13g2_nand2_1 _4601_ (.Y(_1673_),
    .A(net369),
    .B(net1008));
 sg13g2_nand3_1 _4602_ (.B(_1672_),
    .C(_1673_),
    .A(net967),
    .Y(_1674_));
 sg13g2_o21ai_1 _4603_ (.B1(_1674_),
    .Y(_1675_),
    .A1(net1186),
    .A2(net967));
 sg13g2_nor2_1 _4604_ (.A(net1217),
    .B(_1675_),
    .Y(_0241_));
 sg13g2_nand2_1 _4605_ (.Y(_1676_),
    .A(\charlie_0.memory[15][6] ),
    .B(net1003));
 sg13g2_nand2_1 _4606_ (.Y(_1677_),
    .A(net452),
    .B(net1008));
 sg13g2_nand3_1 _4607_ (.B(_1676_),
    .C(_1677_),
    .A(net967),
    .Y(_1678_));
 sg13g2_o21ai_1 _4608_ (.B1(_1678_),
    .Y(_1679_),
    .A1(net1184),
    .A2(net967));
 sg13g2_nor2_1 _4609_ (.A(net1216),
    .B(_1679_),
    .Y(_0242_));
 sg13g2_nand2_1 _4610_ (.Y(_1680_),
    .A(\charlie_0.memory[15][7] ),
    .B(net1003));
 sg13g2_nand2_1 _4611_ (.Y(_1681_),
    .A(\counter[31] ),
    .B(net1007));
 sg13g2_nand3_1 _4612_ (.B(_1680_),
    .C(_1681_),
    .A(net966),
    .Y(_1682_));
 sg13g2_o21ai_1 _4613_ (.B1(_1682_),
    .Y(_1683_),
    .A1(net1213),
    .A2(net966));
 sg13g2_nor2_1 _4614_ (.A(net1215),
    .B(_1683_),
    .Y(_0243_));
 sg13g2_and2_1 _4615_ (.A(_0574_),
    .B(_1338_),
    .X(_1684_));
 sg13g2_o21ai_1 _4616_ (.B1(net1242),
    .Y(_1685_),
    .A1(net1172),
    .A2(net964));
 sg13g2_a21oi_1 _4617_ (.A1(net1230),
    .A2(net964),
    .Y(_0244_),
    .B1(_1685_));
 sg13g2_o21ai_1 _4618_ (.B1(net1242),
    .Y(_1686_),
    .A1(net1170),
    .A2(net964));
 sg13g2_a21oi_1 _4619_ (.A1(net1126),
    .A2(net964),
    .Y(_0245_),
    .B1(_1686_));
 sg13g2_o21ai_1 _4620_ (.B1(net1242),
    .Y(_1687_),
    .A1(net459),
    .A2(net965));
 sg13g2_a21oi_1 _4621_ (.A1(net1128),
    .A2(_1684_),
    .Y(_0246_),
    .B1(_1687_));
 sg13g2_o21ai_1 _4622_ (.B1(net1242),
    .Y(_1688_),
    .A1(net491),
    .A2(net965));
 sg13g2_a21oi_1 _4623_ (.A1(net1133),
    .A2(net965),
    .Y(_0247_),
    .B1(_1688_));
 sg13g2_o21ai_1 _4624_ (.B1(net1242),
    .Y(_1689_),
    .A1(net363),
    .A2(net964));
 sg13g2_a21oi_1 _4625_ (.A1(net1136),
    .A2(net964),
    .Y(_0248_),
    .B1(_1689_));
 sg13g2_o21ai_1 _4626_ (.B1(net1242),
    .Y(_1690_),
    .A1(net463),
    .A2(net965));
 sg13g2_a21oi_1 _4627_ (.A1(net1141),
    .A2(net965),
    .Y(_0249_),
    .B1(_1690_));
 sg13g2_o21ai_1 _4628_ (.B1(net1242),
    .Y(_1691_),
    .A1(net1168),
    .A2(net965));
 sg13g2_a21oi_1 _4629_ (.A1(net1143),
    .A2(net965),
    .Y(_0250_),
    .B1(_1691_));
 sg13g2_o21ai_1 _4630_ (.B1(net1234),
    .Y(_1692_),
    .A1(net314),
    .A2(net964));
 sg13g2_a21oi_1 _4631_ (.A1(net1145),
    .A2(net964),
    .Y(_0251_),
    .B1(_1692_));
 sg13g2_and2_1 _4632_ (.A(_0574_),
    .B(_1350_),
    .X(_1693_));
 sg13g2_o21ai_1 _4633_ (.B1(net1256),
    .Y(_1694_),
    .A1(net1164),
    .A2(net963));
 sg13g2_a21oi_1 _4634_ (.A1(net1228),
    .A2(net963),
    .Y(_0252_),
    .B1(_1694_));
 sg13g2_o21ai_1 _4635_ (.B1(net1256),
    .Y(_1695_),
    .A1(net1161),
    .A2(net963));
 sg13g2_a21oi_1 _4636_ (.A1(net1125),
    .A2(net963),
    .Y(_0253_),
    .B1(_1695_));
 sg13g2_o21ai_1 _4637_ (.B1(net1255),
    .Y(_1696_),
    .A1(net1159),
    .A2(net963));
 sg13g2_a21oi_1 _4638_ (.A1(net1131),
    .A2(net963),
    .Y(_0254_),
    .B1(_1696_));
 sg13g2_o21ai_1 _4639_ (.B1(net1255),
    .Y(_1697_),
    .A1(net1156),
    .A2(net962));
 sg13g2_a21oi_1 _4640_ (.A1(net1134),
    .A2(net962),
    .Y(_0255_),
    .B1(_1697_));
 sg13g2_o21ai_1 _4641_ (.B1(net1255),
    .Y(_1698_),
    .A1(\charlie_0.memory[17][4] ),
    .A2(_1693_));
 sg13g2_a21oi_1 _4642_ (.A1(net1138),
    .A2(net962),
    .Y(_0256_),
    .B1(_1698_));
 sg13g2_o21ai_1 _4643_ (.B1(net1254),
    .Y(_1699_),
    .A1(net468),
    .A2(net962));
 sg13g2_a21oi_1 _4644_ (.A1(net1140),
    .A2(net962),
    .Y(_0257_),
    .B1(_1699_));
 sg13g2_o21ai_1 _4645_ (.B1(net1255),
    .Y(_1700_),
    .A1(\charlie_0.memory[17][6] ),
    .A2(net963));
 sg13g2_a21oi_1 _4646_ (.A1(net1142),
    .A2(net962),
    .Y(_0258_),
    .B1(_1700_));
 sg13g2_o21ai_1 _4647_ (.B1(net1254),
    .Y(_1701_),
    .A1(net357),
    .A2(net962));
 sg13g2_a21oi_1 _4648_ (.A1(net1144),
    .A2(net962),
    .Y(_0259_),
    .B1(_1701_));
 sg13g2_and2_1 _4649_ (.A(_0574_),
    .B(_1361_),
    .X(_1702_));
 sg13g2_o21ai_1 _4650_ (.B1(net1251),
    .Y(_1703_),
    .A1(net458),
    .A2(net960));
 sg13g2_a21oi_1 _4651_ (.A1(net1228),
    .A2(net960),
    .Y(_0260_),
    .B1(_1703_));
 sg13g2_o21ai_1 _4652_ (.B1(net1252),
    .Y(_1704_),
    .A1(net457),
    .A2(net961));
 sg13g2_a21oi_1 _4653_ (.A1(net1125),
    .A2(net961),
    .Y(_0261_),
    .B1(_1704_));
 sg13g2_o21ai_1 _4654_ (.B1(net1253),
    .Y(_1705_),
    .A1(net390),
    .A2(net961));
 sg13g2_a21oi_1 _4655_ (.A1(net1131),
    .A2(net961),
    .Y(_0262_),
    .B1(_1705_));
 sg13g2_o21ai_1 _4656_ (.B1(net1252),
    .Y(_1706_),
    .A1(net473),
    .A2(net961));
 sg13g2_a21oi_1 _4657_ (.A1(net1134),
    .A2(net961),
    .Y(_0263_),
    .B1(_1706_));
 sg13g2_o21ai_1 _4658_ (.B1(net1252),
    .Y(_1707_),
    .A1(net414),
    .A2(net960));
 sg13g2_a21oi_1 _4659_ (.A1(net1138),
    .A2(net960),
    .Y(_0264_),
    .B1(_1707_));
 sg13g2_o21ai_1 _4660_ (.B1(net1252),
    .Y(_1708_),
    .A1(net462),
    .A2(net961));
 sg13g2_a21oi_1 _4661_ (.A1(net1140),
    .A2(net961),
    .Y(_0265_),
    .B1(_1708_));
 sg13g2_o21ai_1 _4662_ (.B1(net1252),
    .Y(_1709_),
    .A1(net469),
    .A2(net960));
 sg13g2_a21oi_1 _4663_ (.A1(net1142),
    .A2(net960),
    .Y(_0266_),
    .B1(_1709_));
 sg13g2_o21ai_1 _4664_ (.B1(net1252),
    .Y(_1710_),
    .A1(net433),
    .A2(net960));
 sg13g2_a21oi_1 _4665_ (.A1(net1144),
    .A2(net960),
    .Y(_0267_),
    .B1(_1710_));
 sg13g2_and2_1 _4666_ (.A(_0574_),
    .B(_1372_),
    .X(_1711_));
 sg13g2_o21ai_1 _4667_ (.B1(net1235),
    .Y(_1712_),
    .A1(net326),
    .A2(net958));
 sg13g2_a21oi_1 _4668_ (.A1(net1230),
    .A2(net958),
    .Y(_0268_),
    .B1(_1712_));
 sg13g2_o21ai_1 _4669_ (.B1(net1236),
    .Y(_1713_),
    .A1(net1154),
    .A2(_1711_));
 sg13g2_a21oi_1 _4670_ (.A1(net1126),
    .A2(net959),
    .Y(_0269_),
    .B1(_1713_));
 sg13g2_o21ai_1 _4671_ (.B1(net1234),
    .Y(_1714_),
    .A1(net315),
    .A2(net958));
 sg13g2_a21oi_1 _4672_ (.A1(net1127),
    .A2(net958),
    .Y(_0270_),
    .B1(_1714_));
 sg13g2_o21ai_1 _4673_ (.B1(net1237),
    .Y(_1715_),
    .A1(net1150),
    .A2(net958));
 sg13g2_a21oi_1 _4674_ (.A1(net1133),
    .A2(net958),
    .Y(_0271_),
    .B1(_1715_));
 sg13g2_o21ai_1 _4675_ (.B1(net1237),
    .Y(_1716_),
    .A1(net1147),
    .A2(net958));
 sg13g2_a21oi_1 _4676_ (.A1(net1136),
    .A2(net958),
    .Y(_0272_),
    .B1(_1716_));
 sg13g2_o21ai_1 _4677_ (.B1(net1239),
    .Y(_1717_),
    .A1(net309),
    .A2(net959));
 sg13g2_a21oi_1 _4678_ (.A1(net1141),
    .A2(net959),
    .Y(_0273_),
    .B1(_1717_));
 sg13g2_o21ai_1 _4679_ (.B1(net1241),
    .Y(_1718_),
    .A1(net332),
    .A2(net959));
 sg13g2_a21oi_1 _4680_ (.A1(net1143),
    .A2(net959),
    .Y(_0274_),
    .B1(_1718_));
 sg13g2_o21ai_1 _4681_ (.B1(net1236),
    .Y(_1719_),
    .A1(net351),
    .A2(net959));
 sg13g2_a21oi_1 _4682_ (.A1(net1145),
    .A2(net959),
    .Y(_0275_),
    .B1(_1719_));
 sg13g2_nand2_1 _4683_ (.Y(_1720_),
    .A(net290),
    .B(_0573_));
 sg13g2_o21ai_1 _4684_ (.B1(_1720_),
    .Y(_1721_),
    .A1(\charlie_0.memory[20][1] ),
    .A2(net999));
 sg13g2_nor2_1 _4685_ (.A(net1223),
    .B(net291),
    .Y(_0276_));
 sg13g2_nand2_1 _4686_ (.Y(_1722_),
    .A(net282),
    .B(_0573_));
 sg13g2_o21ai_1 _4687_ (.B1(_1722_),
    .Y(_1723_),
    .A1(\charlie_0.memory[20][4] ),
    .A2(net998));
 sg13g2_nor2_1 _4688_ (.A(net1223),
    .B(net283),
    .Y(_0277_));
 sg13g2_o21ai_1 _4689_ (.B1(net1237),
    .Y(_1724_),
    .A1(net466),
    .A2(net998));
 sg13g2_a21oi_1 _4690_ (.A1(net1141),
    .A2(net998),
    .Y(_0278_),
    .B1(_1724_));
 sg13g2_o21ai_1 _4691_ (.B1(net1236),
    .Y(_1725_),
    .A1(net341),
    .A2(net998));
 sg13g2_a21oi_1 _4692_ (.A1(net1143),
    .A2(_0573_),
    .Y(_0279_),
    .B1(_1725_));
 sg13g2_o21ai_1 _4693_ (.B1(net1236),
    .Y(_1726_),
    .A1(\charlie_0.memory[20][7] ),
    .A2(net998));
 sg13g2_a21oi_1 _4694_ (.A1(net299),
    .A2(_0573_),
    .Y(_0280_),
    .B1(_1726_));
 sg13g2_nand2_1 _4695_ (.Y(_1727_),
    .A(_0572_),
    .B(_1391_));
 sg13g2_and2_1 _4696_ (.A(_0574_),
    .B(_1391_),
    .X(_1728_));
 sg13g2_nand2_2 _4697_ (.Y(_1729_),
    .A(_0574_),
    .B(_1391_));
 sg13g2_nand3_1 _4698_ (.B(net1021),
    .C(_1729_),
    .A(\charlie_0.memory[21][0] ),
    .Y(_1730_));
 sg13g2_nor2_1 _4699_ (.A(net1021),
    .B(net957),
    .Y(_1731_));
 sg13g2_a22oi_1 _4700_ (.Y(_1732_),
    .B1(_1731_),
    .B2(net276),
    .A2(net957),
    .A1(net1233));
 sg13g2_a21oi_1 _4701_ (.A1(_1730_),
    .A2(_1732_),
    .Y(_0281_),
    .B1(net1227));
 sg13g2_nand3_1 _4702_ (.B(\charlie_0.memory[21][0] ),
    .C(_0565_),
    .A(\charlie_0.memory[21][1] ),
    .Y(_1733_));
 sg13g2_a21o_1 _4703_ (.A2(_0565_),
    .A1(\charlie_0.memory[21][0] ),
    .B1(\charlie_0.memory[21][1] ),
    .X(_1734_));
 sg13g2_and2_1 _4704_ (.A(_1733_),
    .B(_1734_),
    .X(_1735_));
 sg13g2_o21ai_1 _4705_ (.B1(net1239),
    .Y(_1736_),
    .A1(net957),
    .A2(_1735_));
 sg13g2_a21oi_1 _4706_ (.A1(net1126),
    .A2(net957),
    .Y(_0282_),
    .B1(_1736_));
 sg13g2_nand3_1 _4707_ (.B(\charlie_0.memory[21][1] ),
    .C(\charlie_0.memory[21][0] ),
    .A(\charlie_0.memory[21][2] ),
    .Y(_1737_));
 sg13g2_nor2_1 _4708_ (.A(net1021),
    .B(_1737_),
    .Y(_1738_));
 sg13g2_xnor2_1 _4709_ (.Y(_1739_),
    .A(\charlie_0.memory[21][2] ),
    .B(_1733_));
 sg13g2_o21ai_1 _4710_ (.B1(net1239),
    .Y(_1740_),
    .A1(net957),
    .A2(_1739_));
 sg13g2_a21oi_1 _4711_ (.A1(net1127),
    .A2(net957),
    .Y(_0283_),
    .B1(_1740_));
 sg13g2_xor2_1 _4712_ (.B(_1738_),
    .A(\charlie_0.memory[21][3] ),
    .X(_1741_));
 sg13g2_o21ai_1 _4713_ (.B1(net1239),
    .Y(_1742_),
    .A1(net957),
    .A2(_1741_));
 sg13g2_a21oi_1 _4714_ (.A1(net1133),
    .A2(_1728_),
    .Y(_0284_),
    .B1(_1742_));
 sg13g2_a21oi_1 _4715_ (.A1(\charlie_0.memory[21][3] ),
    .A2(_1738_),
    .Y(_1743_),
    .B1(\charlie_0.memory[21][4] ));
 sg13g2_and3_1 _4716_ (.X(_1744_),
    .A(\charlie_0.memory[21][4] ),
    .B(\charlie_0.memory[21][3] ),
    .C(_1738_));
 sg13g2_o21ai_1 _4717_ (.B1(_1729_),
    .Y(_1745_),
    .A1(_1743_),
    .A2(_1744_));
 sg13g2_o21ai_1 _4718_ (.B1(_1745_),
    .Y(_1746_),
    .A1(net1188),
    .A2(_1727_));
 sg13g2_nor2_1 _4719_ (.A(net1223),
    .B(_1746_),
    .Y(_0285_));
 sg13g2_xnor2_1 _4720_ (.Y(_1747_),
    .A(net358),
    .B(_1744_));
 sg13g2_o21ai_1 _4721_ (.B1(net1239),
    .Y(_1748_),
    .A1(net1186),
    .A2(_1727_));
 sg13g2_a21oi_1 _4722_ (.A1(_1729_),
    .A2(_1747_),
    .Y(_0286_),
    .B1(_1748_));
 sg13g2_nand4_1 _4723_ (.B(\charlie_0.memory[21][5] ),
    .C(\charlie_0.memory[21][4] ),
    .A(\charlie_0.memory[21][6] ),
    .Y(_1749_),
    .D(\charlie_0.memory[21][3] ));
 sg13g2_nor2_1 _4724_ (.A(_1737_),
    .B(_1749_),
    .Y(_1750_));
 sg13g2_a21oi_1 _4725_ (.A1(\charlie_0.memory[21][5] ),
    .A2(_1744_),
    .Y(_1751_),
    .B1(net320));
 sg13g2_o21ai_1 _4726_ (.B1(net1239),
    .Y(_1752_),
    .A1(net1184),
    .A2(_1729_));
 sg13g2_a221oi_1 _4727_ (.B2(_1729_),
    .C1(_1752_),
    .B1(net321),
    .A1(_1731_),
    .Y(_0287_),
    .A2(_1750_));
 sg13g2_nand3_1 _4728_ (.B(net1021),
    .C(_1729_),
    .A(net310),
    .Y(_1753_));
 sg13g2_xor2_1 _4729_ (.B(_1750_),
    .A(net310),
    .X(_1754_));
 sg13g2_a22oi_1 _4730_ (.Y(_1755_),
    .B1(_1731_),
    .B2(_1754_),
    .A2(net957),
    .A1(net1213));
 sg13g2_a21oi_1 _4731_ (.A1(_1753_),
    .A2(_1755_),
    .Y(_0288_),
    .B1(net1227));
 sg13g2_o21ai_1 _4732_ (.B1(\charlie_0.memory[20][3] ),
    .Y(_1756_),
    .A1(_0562_),
    .A2(_0567_));
 sg13g2_inv_1 _4733_ (.Y(_1757_),
    .A(_1756_));
 sg13g2_o21ai_1 _4734_ (.B1(net1237),
    .Y(_1758_),
    .A1(net999),
    .A2(_1757_));
 sg13g2_a21oi_1 _4735_ (.A1(net273),
    .A2(net999),
    .Y(_0289_),
    .B1(_1758_));
 sg13g2_and2_1 _4736_ (.A(_0574_),
    .B(_1401_),
    .X(_1759_));
 sg13g2_o21ai_1 _4737_ (.B1(net1239),
    .Y(_1760_),
    .A1(net1146),
    .A2(net955));
 sg13g2_a21oi_1 _4738_ (.A1(net1228),
    .A2(net956),
    .Y(_0290_),
    .B1(_1760_));
 sg13g2_o21ai_1 _4739_ (.B1(net1240),
    .Y(_1761_),
    .A1(net481),
    .A2(net955));
 sg13g2_a21oi_1 _4740_ (.A1(net1126),
    .A2(net955),
    .Y(_0291_),
    .B1(_1761_));
 sg13g2_o21ai_1 _4741_ (.B1(net1240),
    .Y(_1762_),
    .A1(net323),
    .A2(net956));
 sg13g2_a21oi_1 _4742_ (.A1(net1131),
    .A2(net956),
    .Y(_0292_),
    .B1(_1762_));
 sg13g2_o21ai_1 _4743_ (.B1(net1252),
    .Y(_1763_),
    .A1(net366),
    .A2(_1759_));
 sg13g2_a21oi_1 _4744_ (.A1(net1133),
    .A2(net956),
    .Y(_0293_),
    .B1(_1763_));
 sg13g2_o21ai_1 _4745_ (.B1(net1239),
    .Y(_1764_),
    .A1(net388),
    .A2(net955));
 sg13g2_a21oi_1 _4746_ (.A1(net1137),
    .A2(net955),
    .Y(_0294_),
    .B1(_1764_));
 sg13g2_o21ai_1 _4747_ (.B1(net1252),
    .Y(_1765_),
    .A1(net455),
    .A2(net956));
 sg13g2_a21oi_1 _4748_ (.A1(net1141),
    .A2(net956),
    .Y(_0295_),
    .B1(_1765_));
 sg13g2_o21ai_1 _4749_ (.B1(net1240),
    .Y(_1766_),
    .A1(net432),
    .A2(net955));
 sg13g2_a21oi_1 _4750_ (.A1(net1142),
    .A2(net955),
    .Y(_0296_),
    .B1(_1766_));
 sg13g2_o21ai_1 _4751_ (.B1(net1251),
    .Y(_1767_),
    .A1(net386),
    .A2(net956));
 sg13g2_a21oi_1 _4752_ (.A1(net1144),
    .A2(net955),
    .Y(_0297_),
    .B1(_1767_));
 sg13g2_dfrbp_1 _4753_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net11),
    .D(_0081_),
    .Q_N(_0066_),
    .Q(\gen_priority_write_blocks[0].this_priority_write.data_bits[15] ));
 sg13g2_dfrbp_1 _4754_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net265),
    .D(net289),
    .Q_N(_2320_),
    .Q(\charlie_0.memory[20][2] ));
 sg13g2_dfrbp_1 _4755_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net12),
    .D(_0083_),
    .Q_N(_2321_),
    .Q(\spi_slave_0.spi_clk_prev ));
 sg13g2_dfrbp_1 _4756_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net13),
    .D(_0016_),
    .Q_N(_0075_),
    .Q(\charlie_0.charlie_index[0] ));
 sg13g2_dfrbp_1 _4757_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net14),
    .D(_0027_),
    .Q_N(_2322_),
    .Q(\charlie_0.charlie_index[1] ));
 sg13g2_dfrbp_1 _4758_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net15),
    .D(_0038_),
    .Q_N(_0069_),
    .Q(\charlie_0.charlie_index[2] ));
 sg13g2_dfrbp_1 _4759_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net16),
    .D(_0041_),
    .Q_N(_0068_),
    .Q(\charlie_0.charlie_index[3] ));
 sg13g2_dfrbp_1 _4760_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net17),
    .D(_0042_),
    .Q_N(_2323_),
    .Q(\charlie_0.charlie_index[4] ));
 sg13g2_dfrbp_1 _4761_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net18),
    .D(_0043_),
    .Q_N(_0063_),
    .Q(\charlie_0.charlie_index[5] ));
 sg13g2_dfrbp_1 _4762_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net19),
    .D(_0044_),
    .Q_N(_2324_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 _4763_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net20),
    .D(_0045_),
    .Q_N(_2325_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 _4764_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net21),
    .D(net334),
    .Q_N(_2326_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 _4765_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net22),
    .D(_0047_),
    .Q_N(_2327_),
    .Q(\counter[9] ));
 sg13g2_dfrbp_1 _4766_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net23),
    .D(net378),
    .Q_N(_2328_),
    .Q(\counter[10] ));
 sg13g2_dfrbp_1 _4767_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net24),
    .D(_0018_),
    .Q_N(_2329_),
    .Q(\counter[11] ));
 sg13g2_dfrbp_1 _4768_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net25),
    .D(net345),
    .Q_N(_2330_),
    .Q(\counter[12] ));
 sg13g2_dfrbp_1 _4769_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net26),
    .D(_0020_),
    .Q_N(_2331_),
    .Q(\counter[13] ));
 sg13g2_dfrbp_1 _4770_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net27),
    .D(net348),
    .Q_N(_2332_),
    .Q(\counter[14] ));
 sg13g2_dfrbp_1 _4771_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net28),
    .D(net361),
    .Q_N(_2333_),
    .Q(\counter[15] ));
 sg13g2_dfrbp_1 _4772_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net29),
    .D(_0023_),
    .Q_N(_2334_),
    .Q(\counter[16] ));
 sg13g2_dfrbp_1 _4773_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net30),
    .D(_0024_),
    .Q_N(_2335_),
    .Q(\counter[17] ));
 sg13g2_dfrbp_1 _4774_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net31),
    .D(net405),
    .Q_N(_2336_),
    .Q(\counter[18] ));
 sg13g2_dfrbp_1 _4775_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net32),
    .D(_0026_),
    .Q_N(_2337_),
    .Q(\counter[19] ));
 sg13g2_dfrbp_1 _4776_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net33),
    .D(net410),
    .Q_N(_2338_),
    .Q(\counter[20] ));
 sg13g2_dfrbp_1 _4777_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net34),
    .D(_0029_),
    .Q_N(_2339_),
    .Q(\counter[21] ));
 sg13g2_dfrbp_1 _4778_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net35),
    .D(_0030_),
    .Q_N(_2340_),
    .Q(\counter[22] ));
 sg13g2_dfrbp_1 _4779_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net36),
    .D(_0031_),
    .Q_N(_2341_),
    .Q(\counter[23] ));
 sg13g2_dfrbp_1 _4780_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net37),
    .D(net380),
    .Q_N(_2342_),
    .Q(\counter[24] ));
 sg13g2_dfrbp_1 _4781_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net38),
    .D(_0033_),
    .Q_N(_2343_),
    .Q(\counter[25] ));
 sg13g2_dfrbp_1 _4782_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net39),
    .D(net354),
    .Q_N(_2344_),
    .Q(\counter[26] ));
 sg13g2_dfrbp_1 _4783_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net40),
    .D(_0035_),
    .Q_N(_2345_),
    .Q(\counter[27] ));
 sg13g2_dfrbp_1 _4784_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net41),
    .D(net397),
    .Q_N(_2346_),
    .Q(\counter[28] ));
 sg13g2_dfrbp_1 _4785_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net42),
    .D(_0037_),
    .Q_N(_2347_),
    .Q(\counter[29] ));
 sg13g2_dfrbp_1 _4786_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net43),
    .D(net370),
    .Q_N(_2348_),
    .Q(\counter[30] ));
 sg13g2_dfrbp_1 _4787_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net44),
    .D(_0040_),
    .Q_N(_2349_),
    .Q(\counter[31] ));
 sg13g2_dfrbp_1 _4788_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net45),
    .D(_0000_),
    .Q_N(_2350_),
    .Q(\bi_en[0] ));
 sg13g2_dfrbp_1 _4789_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net46),
    .D(_0001_),
    .Q_N(_2351_),
    .Q(\bi_en[1] ));
 sg13g2_dfrbp_1 _4790_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net47),
    .D(_0002_),
    .Q_N(_2352_),
    .Q(\bi_en[2] ));
 sg13g2_dfrbp_1 _4791_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net48),
    .D(_0003_),
    .Q_N(_2353_),
    .Q(\bi_en[3] ));
 sg13g2_dfrbp_1 _4792_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net49),
    .D(_0004_),
    .Q_N(_2354_),
    .Q(\bi_en[4] ));
 sg13g2_dfrbp_1 _4793_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net50),
    .D(_0005_),
    .Q_N(_2355_),
    .Q(\bi_en[5] ));
 sg13g2_dfrbp_1 _4794_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net51),
    .D(_0006_),
    .Q_N(_2356_),
    .Q(\bi_en[6] ));
 sg13g2_dfrbp_1 _4795_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net52),
    .D(_0007_),
    .Q_N(_2357_),
    .Q(\bi_en[7] ));
 sg13g2_dfrbp_1 _4796_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net53),
    .D(_0008_),
    .Q_N(_2358_),
    .Q(\bi_out[0] ));
 sg13g2_dfrbp_1 _4797_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net54),
    .D(_0009_),
    .Q_N(_2359_),
    .Q(\bi_out[1] ));
 sg13g2_dfrbp_1 _4798_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net55),
    .D(_0010_),
    .Q_N(_2360_),
    .Q(\bi_out[2] ));
 sg13g2_dfrbp_1 _4799_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net56),
    .D(_0011_),
    .Q_N(_2361_),
    .Q(\bi_out[3] ));
 sg13g2_dfrbp_1 _4800_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net57),
    .D(_0012_),
    .Q_N(_2362_),
    .Q(\bi_out[4] ));
 sg13g2_dfrbp_1 _4801_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net58),
    .D(_0013_),
    .Q_N(_2363_),
    .Q(\bi_out[5] ));
 sg13g2_dfrbp_1 _4802_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net94),
    .D(_0014_),
    .Q_N(_2364_),
    .Q(\bi_out[6] ));
 sg13g2_dfrbp_1 _4803_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net263),
    .D(_0015_),
    .Q_N(_2319_),
    .Q(\bi_out[7] ));
 sg13g2_dfrbp_1 _4804_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net262),
    .D(_0084_),
    .Q_N(_2318_),
    .Q(\charlie_0.memory[20][0] ));
 sg13g2_dfrbp_1 _4805_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net260),
    .D(_0085_),
    .Q_N(_0079_),
    .Q(\gen_priority_write_blocks[0].this_priority_write.data_bits[9] ));
 sg13g2_dfrbp_1 _4806_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net258),
    .D(_0086_),
    .Q_N(_0078_),
    .Q(\gen_priority_write_blocks[0].this_priority_write.data_bits[10] ));
 sg13g2_dfrbp_1 _4807_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net256),
    .D(_0087_),
    .Q_N(_0077_),
    .Q(\gen_priority_write_blocks[0].this_priority_write.data_bits[11] ));
 sg13g2_dfrbp_1 _4808_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net254),
    .D(_0088_),
    .Q_N(_0076_),
    .Q(\gen_priority_write_blocks[0].this_priority_write.data_bits[12] ));
 sg13g2_dfrbp_1 _4809_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net252),
    .D(_0089_),
    .Q_N(_2317_),
    .Q(\gen_priority_write_blocks[0].this_priority_write.data_bits[13] ));
 sg13g2_dfrbp_1 _4810_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net250),
    .D(_0090_),
    .Q_N(_2316_),
    .Q(\gen_priority_write_blocks[0].this_priority_write.data_bits[14] ));
 sg13g2_dfrbp_1 _4811_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net248),
    .D(_0091_),
    .Q_N(_2315_),
    .Q(\spi_slave_0.reg_data[7] ));
 sg13g2_dfrbp_1 _4812_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net246),
    .D(_0092_),
    .Q_N(_2314_),
    .Q(\spi_address[0] ));
 sg13g2_dfrbp_1 _4813_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net244),
    .D(_0093_),
    .Q_N(_2313_),
    .Q(\spi_address[1] ));
 sg13g2_dfrbp_1 _4814_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net242),
    .D(_0094_),
    .Q_N(_0074_),
    .Q(\spi_address[2] ));
 sg13g2_dfrbp_1 _4815_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net240),
    .D(_0095_),
    .Q_N(_0072_),
    .Q(\spi_address[3] ));
 sg13g2_dfrbp_1 _4816_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net238),
    .D(_0096_),
    .Q_N(_0071_),
    .Q(\spi_address[4] ));
 sg13g2_dfrbp_1 _4817_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net236),
    .D(net287),
    .Q_N(_0073_),
    .Q(\spi_slave_0.is_mosi ));
 sg13g2_dfrbp_1 _4818_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net234),
    .D(net275),
    .Q_N(_0080_),
    .Q(\spi_slave_0.bit_cnt[0] ));
 sg13g2_dfrbp_1 _4819_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net232),
    .D(net294),
    .Q_N(_2312_),
    .Q(\spi_slave_0.bit_cnt[1] ));
 sg13g2_dfrbp_1 _4820_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net230),
    .D(net298),
    .Q_N(_2311_),
    .Q(\spi_slave_0.bit_cnt[2] ));
 sg13g2_dfrbp_1 _4821_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net228),
    .D(net285),
    .Q_N(_2310_),
    .Q(miso));
 sg13g2_dfrbp_1 _4822_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net226),
    .D(_0102_),
    .Q_N(_2309_),
    .Q(\signal_generator_0.state_machine[0] ));
 sg13g2_dfrbp_1 _4823_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net225),
    .D(net339),
    .Q_N(_2308_),
    .Q(\signal_generator_0.state_machine[1] ));
 sg13g2_dfrbp_1 _4824_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net224),
    .D(_0104_),
    .Q_N(_2307_),
    .Q(\spi_slave_0.is_data_phase ));
 sg13g2_dfrbp_1 _4825_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net222),
    .D(net384),
    .Q_N(_0056_),
    .Q(sig_gen_out));
 sg13g2_dfrbp_1 _4826_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net221),
    .D(_0106_),
    .Q_N(_2306_),
    .Q(\signal_generator_0.prev_clk_div ));
 sg13g2_dfrbp_1 _4827_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net220),
    .D(net279),
    .Q_N(_0049_),
    .Q(\signal_generator_0.index_reg[0] ));
 sg13g2_dfrbp_1 _4828_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net218),
    .D(_0108_),
    .Q_N(_2305_),
    .Q(\signal_generator_0.index_reg[1] ));
 sg13g2_dfrbp_1 _4829_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net216),
    .D(_0109_),
    .Q_N(_2304_),
    .Q(\signal_generator_0.index_reg[2] ));
 sg13g2_dfrbp_1 _4830_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net214),
    .D(_0110_),
    .Q_N(_2303_),
    .Q(\signal_generator_0.index_reg[3] ));
 sg13g2_dfrbp_1 _4831_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net212),
    .D(net436),
    .Q_N(_2302_),
    .Q(\signal_generator_0.index_reg[4] ));
 sg13g2_dfrbp_1 _4832_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net210),
    .D(_0112_),
    .Q_N(_2301_),
    .Q(\signal_generator_0.index_reg[5] ));
 sg13g2_dfrbp_1 _4833_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net208),
    .D(_0113_),
    .Q_N(_2300_),
    .Q(\signal_generator_0.index_reg[6] ));
 sg13g2_dfrbp_1 _4834_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net206),
    .D(_0114_),
    .Q_N(_2299_),
    .Q(\signal_generator_0.index_reg[7] ));
 sg13g2_dfrbp_1 _4835_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net204),
    .D(_0115_),
    .Q_N(_0070_),
    .Q(\signal_generator_0.prev_trigger ));
 sg13g2_dfrbp_1 _4836_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net203),
    .D(_0116_),
    .Q_N(_0055_),
    .Q(\charlie_0.memory[0][0] ));
 sg13g2_dfrbp_1 _4837_ (.CLK(clknet_3_6__leaf_clk_regs),
    .RESET_B(net201),
    .D(_0117_),
    .Q_N(_0057_),
    .Q(\charlie_0.memory[0][1] ));
 sg13g2_dfrbp_1 _4838_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net199),
    .D(_0118_),
    .Q_N(_0058_),
    .Q(\charlie_0.memory[0][2] ));
 sg13g2_dfrbp_1 _4839_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net197),
    .D(_0119_),
    .Q_N(_0059_),
    .Q(\charlie_0.memory[0][3] ));
 sg13g2_dfrbp_1 _4840_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net195),
    .D(_0120_),
    .Q_N(_0060_),
    .Q(\charlie_0.memory[0][4] ));
 sg13g2_dfrbp_1 _4841_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net193),
    .D(_0121_),
    .Q_N(_0061_),
    .Q(\charlie_0.memory[0][5] ));
 sg13g2_dfrbp_1 _4842_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net191),
    .D(_0122_),
    .Q_N(_0062_),
    .Q(\charlie_0.memory[0][6] ));
 sg13g2_dfrbp_1 _4843_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net189),
    .D(_0123_),
    .Q_N(_0065_),
    .Q(\charlie_0.memory[0][7] ));
 sg13g2_dfrbp_1 _4844_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net187),
    .D(_0124_),
    .Q_N(_2298_),
    .Q(\charlie_0.memory[1][0] ));
 sg13g2_dfrbp_1 _4845_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net185),
    .D(_0125_),
    .Q_N(_2297_),
    .Q(\charlie_0.memory[1][1] ));
 sg13g2_dfrbp_1 _4846_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net183),
    .D(_0126_),
    .Q_N(_2296_),
    .Q(\charlie_0.memory[1][2] ));
 sg13g2_dfrbp_1 _4847_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net181),
    .D(_0127_),
    .Q_N(_2295_),
    .Q(\charlie_0.memory[1][3] ));
 sg13g2_dfrbp_1 _4848_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net179),
    .D(_0128_),
    .Q_N(_2294_),
    .Q(\charlie_0.memory[1][4] ));
 sg13g2_dfrbp_1 _4849_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net177),
    .D(_0129_),
    .Q_N(_2293_),
    .Q(\charlie_0.memory[1][5] ));
 sg13g2_dfrbp_1 _4850_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net175),
    .D(_0130_),
    .Q_N(_2292_),
    .Q(\charlie_0.memory[1][6] ));
 sg13g2_dfrbp_1 _4851_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net173),
    .D(_0131_),
    .Q_N(_2291_),
    .Q(\charlie_0.memory[1][7] ));
 sg13g2_dfrbp_1 _4852_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net171),
    .D(_0132_),
    .Q_N(_2290_),
    .Q(\charlie_0.memory[2][0] ));
 sg13g2_dfrbp_1 _4853_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net169),
    .D(_0133_),
    .Q_N(_2289_),
    .Q(\charlie_0.memory[2][1] ));
 sg13g2_dfrbp_1 _4854_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net167),
    .D(_0134_),
    .Q_N(_2288_),
    .Q(\charlie_0.memory[2][2] ));
 sg13g2_dfrbp_1 _4855_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net165),
    .D(_0135_),
    .Q_N(_2287_),
    .Q(\charlie_0.memory[2][3] ));
 sg13g2_dfrbp_1 _4856_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net163),
    .D(_0136_),
    .Q_N(_2286_),
    .Q(\charlie_0.memory[2][4] ));
 sg13g2_dfrbp_1 _4857_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net161),
    .D(_0137_),
    .Q_N(_2285_),
    .Q(\charlie_0.memory[2][5] ));
 sg13g2_dfrbp_1 _4858_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net159),
    .D(_0138_),
    .Q_N(_2284_),
    .Q(\charlie_0.memory[2][6] ));
 sg13g2_dfrbp_1 _4859_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net157),
    .D(_0139_),
    .Q_N(_2283_),
    .Q(\charlie_0.memory[2][7] ));
 sg13g2_dfrbp_1 _4860_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net155),
    .D(_0140_),
    .Q_N(_2282_),
    .Q(\charlie_0.memory[3][0] ));
 sg13g2_dfrbp_1 _4861_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net153),
    .D(_0141_),
    .Q_N(_2281_),
    .Q(\charlie_0.memory[3][1] ));
 sg13g2_dfrbp_1 _4862_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net151),
    .D(_0142_),
    .Q_N(_2280_),
    .Q(\charlie_0.memory[3][2] ));
 sg13g2_dfrbp_1 _4863_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net149),
    .D(_0143_),
    .Q_N(_2279_),
    .Q(\charlie_0.memory[3][3] ));
 sg13g2_dfrbp_1 _4864_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net147),
    .D(_0144_),
    .Q_N(_2278_),
    .Q(\charlie_0.memory[3][4] ));
 sg13g2_dfrbp_1 _4865_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net145),
    .D(_0145_),
    .Q_N(_2277_),
    .Q(\charlie_0.memory[3][5] ));
 sg13g2_dfrbp_1 _4866_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net143),
    .D(_0146_),
    .Q_N(_2276_),
    .Q(\charlie_0.memory[3][6] ));
 sg13g2_dfrbp_1 _4867_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net141),
    .D(_0147_),
    .Q_N(_2275_),
    .Q(\charlie_0.memory[3][7] ));
 sg13g2_dfrbp_1 _4868_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net139),
    .D(_0148_),
    .Q_N(_2274_),
    .Q(\charlie_0.memory[4][0] ));
 sg13g2_dfrbp_1 _4869_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net137),
    .D(_0149_),
    .Q_N(_2273_),
    .Q(\charlie_0.memory[4][1] ));
 sg13g2_dfrbp_1 _4870_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net135),
    .D(_0150_),
    .Q_N(_2272_),
    .Q(\charlie_0.memory[4][2] ));
 sg13g2_dfrbp_1 _4871_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net133),
    .D(_0151_),
    .Q_N(_2271_),
    .Q(\charlie_0.memory[4][3] ));
 sg13g2_dfrbp_1 _4872_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net131),
    .D(_0152_),
    .Q_N(_2270_),
    .Q(\charlie_0.memory[4][4] ));
 sg13g2_dfrbp_1 _4873_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net129),
    .D(_0153_),
    .Q_N(_2269_),
    .Q(\charlie_0.memory[4][5] ));
 sg13g2_dfrbp_1 _4874_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net127),
    .D(_0154_),
    .Q_N(_2268_),
    .Q(\charlie_0.memory[4][6] ));
 sg13g2_dfrbp_1 _4875_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net125),
    .D(_0155_),
    .Q_N(_2267_),
    .Q(\charlie_0.memory[4][7] ));
 sg13g2_dfrbp_1 _4876_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net123),
    .D(_0156_),
    .Q_N(_2266_),
    .Q(\charlie_0.memory[5][0] ));
 sg13g2_dfrbp_1 _4877_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net121),
    .D(_0157_),
    .Q_N(_2265_),
    .Q(\charlie_0.memory[5][1] ));
 sg13g2_dfrbp_1 _4878_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net119),
    .D(_0158_),
    .Q_N(_2264_),
    .Q(\charlie_0.memory[5][2] ));
 sg13g2_dfrbp_1 _4879_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net117),
    .D(_0159_),
    .Q_N(_2263_),
    .Q(\charlie_0.memory[5][3] ));
 sg13g2_dfrbp_1 _4880_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net115),
    .D(_0160_),
    .Q_N(_2262_),
    .Q(\charlie_0.memory[5][4] ));
 sg13g2_dfrbp_1 _4881_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net113),
    .D(_0161_),
    .Q_N(_2261_),
    .Q(\charlie_0.memory[5][5] ));
 sg13g2_dfrbp_1 _4882_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net111),
    .D(_0162_),
    .Q_N(_2260_),
    .Q(\charlie_0.memory[5][6] ));
 sg13g2_dfrbp_1 _4883_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net109),
    .D(_0163_),
    .Q_N(_2259_),
    .Q(\charlie_0.memory[5][7] ));
 sg13g2_dfrbp_1 _4884_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net107),
    .D(_0164_),
    .Q_N(_2258_),
    .Q(\charlie_0.memory[6][0] ));
 sg13g2_dfrbp_1 _4885_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net105),
    .D(_0165_),
    .Q_N(_2257_),
    .Q(\charlie_0.memory[6][1] ));
 sg13g2_dfrbp_1 _4886_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net103),
    .D(_0166_),
    .Q_N(_2256_),
    .Q(\charlie_0.memory[6][2] ));
 sg13g2_dfrbp_1 _4887_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net101),
    .D(_0167_),
    .Q_N(_2255_),
    .Q(\charlie_0.memory[6][3] ));
 sg13g2_dfrbp_1 _4888_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net99),
    .D(_0168_),
    .Q_N(_2254_),
    .Q(\charlie_0.memory[6][4] ));
 sg13g2_dfrbp_1 _4889_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net97),
    .D(_0169_),
    .Q_N(_2253_),
    .Q(\charlie_0.memory[6][5] ));
 sg13g2_dfrbp_1 _4890_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net95),
    .D(_0170_),
    .Q_N(_2252_),
    .Q(\charlie_0.memory[6][6] ));
 sg13g2_dfrbp_1 _4891_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net93),
    .D(_0171_),
    .Q_N(_2251_),
    .Q(\charlie_0.memory[6][7] ));
 sg13g2_dfrbp_1 _4892_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net91),
    .D(_0172_),
    .Q_N(_2250_),
    .Q(\charlie_0.memory[7][0] ));
 sg13g2_dfrbp_1 _4893_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net89),
    .D(_0173_),
    .Q_N(_2249_),
    .Q(\charlie_0.memory[7][1] ));
 sg13g2_dfrbp_1 _4894_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net87),
    .D(_0174_),
    .Q_N(_2248_),
    .Q(\charlie_0.memory[7][2] ));
 sg13g2_dfrbp_1 _4895_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net85),
    .D(_0175_),
    .Q_N(_2247_),
    .Q(\charlie_0.memory[7][3] ));
 sg13g2_dfrbp_1 _4896_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net83),
    .D(_0176_),
    .Q_N(_2246_),
    .Q(\charlie_0.memory[7][4] ));
 sg13g2_dfrbp_1 _4897_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net81),
    .D(_0177_),
    .Q_N(_2245_),
    .Q(\charlie_0.memory[7][5] ));
 sg13g2_dfrbp_1 _4898_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net79),
    .D(_0178_),
    .Q_N(_2244_),
    .Q(\charlie_0.memory[7][6] ));
 sg13g2_dfrbp_1 _4899_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net77),
    .D(_0179_),
    .Q_N(_2243_),
    .Q(\charlie_0.memory[7][7] ));
 sg13g2_dfrbp_1 _4900_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net75),
    .D(_0180_),
    .Q_N(_2242_),
    .Q(\charlie_0.memory[8][0] ));
 sg13g2_dfrbp_1 _4901_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net73),
    .D(_0181_),
    .Q_N(_2241_),
    .Q(\charlie_0.memory[8][1] ));
 sg13g2_dfrbp_1 _4902_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net71),
    .D(_0182_),
    .Q_N(_2240_),
    .Q(\charlie_0.memory[8][2] ));
 sg13g2_dfrbp_1 _4903_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net69),
    .D(_0183_),
    .Q_N(_2239_),
    .Q(\charlie_0.memory[8][3] ));
 sg13g2_dfrbp_1 _4904_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net67),
    .D(_0184_),
    .Q_N(_2238_),
    .Q(\charlie_0.memory[8][4] ));
 sg13g2_dfrbp_1 _4905_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net65),
    .D(_0185_),
    .Q_N(_2237_),
    .Q(\charlie_0.memory[8][5] ));
 sg13g2_dfrbp_1 _4906_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net63),
    .D(_0186_),
    .Q_N(_2236_),
    .Q(\charlie_0.memory[8][6] ));
 sg13g2_dfrbp_1 _4907_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net61),
    .D(_0187_),
    .Q_N(_2235_),
    .Q(\charlie_0.memory[8][7] ));
 sg13g2_dfrbp_1 _4908_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net59),
    .D(_0188_),
    .Q_N(_2234_),
    .Q(\charlie_0.memory[9][0] ));
 sg13g2_dfrbp_1 _4909_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net9),
    .D(_0189_),
    .Q_N(_2233_),
    .Q(\charlie_0.memory[9][1] ));
 sg13g2_dfrbp_1 _4910_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net272),
    .D(_0190_),
    .Q_N(_2232_),
    .Q(\charlie_0.memory[9][2] ));
 sg13g2_dfrbp_1 _4911_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net270),
    .D(_0191_),
    .Q_N(_2231_),
    .Q(\charlie_0.memory[9][3] ));
 sg13g2_dfrbp_1 _4912_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net268),
    .D(_0192_),
    .Q_N(_2230_),
    .Q(\charlie_0.memory[9][4] ));
 sg13g2_dfrbp_1 _4913_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net266),
    .D(_0193_),
    .Q_N(_2229_),
    .Q(\charlie_0.memory[9][5] ));
 sg13g2_dfrbp_1 _4914_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net261),
    .D(_0194_),
    .Q_N(_2228_),
    .Q(\charlie_0.memory[9][6] ));
 sg13g2_dfrbp_1 _4915_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net257),
    .D(_0195_),
    .Q_N(_2227_),
    .Q(\charlie_0.memory[9][7] ));
 sg13g2_dfrbp_1 _4916_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net253),
    .D(_0196_),
    .Q_N(_2226_),
    .Q(\charlie_0.memory[10][0] ));
 sg13g2_dfrbp_1 _4917_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net249),
    .D(_0197_),
    .Q_N(_2225_),
    .Q(\charlie_0.memory[10][1] ));
 sg13g2_dfrbp_1 _4918_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net245),
    .D(_0198_),
    .Q_N(_2224_),
    .Q(\charlie_0.memory[10][2] ));
 sg13g2_dfrbp_1 _4919_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net241),
    .D(_0199_),
    .Q_N(_2223_),
    .Q(\charlie_0.memory[10][3] ));
 sg13g2_dfrbp_1 _4920_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net237),
    .D(_0200_),
    .Q_N(_2222_),
    .Q(\charlie_0.memory[10][4] ));
 sg13g2_dfrbp_1 _4921_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net233),
    .D(_0201_),
    .Q_N(_2221_),
    .Q(\charlie_0.memory[10][5] ));
 sg13g2_dfrbp_1 _4922_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net229),
    .D(_0202_),
    .Q_N(_2220_),
    .Q(\charlie_0.memory[10][6] ));
 sg13g2_dfrbp_1 _4923_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net223),
    .D(_0203_),
    .Q_N(_2219_),
    .Q(\charlie_0.memory[10][7] ));
 sg13g2_dfrbp_1 _4924_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net217),
    .D(_0204_),
    .Q_N(_2218_),
    .Q(\charlie_0.memory[11][0] ));
 sg13g2_dfrbp_1 _4925_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net213),
    .D(_0205_),
    .Q_N(_2217_),
    .Q(\charlie_0.memory[11][1] ));
 sg13g2_dfrbp_1 _4926_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net209),
    .D(_0206_),
    .Q_N(_2216_),
    .Q(\charlie_0.memory[11][2] ));
 sg13g2_dfrbp_1 _4927_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net205),
    .D(_0207_),
    .Q_N(_2215_),
    .Q(\charlie_0.memory[11][3] ));
 sg13g2_dfrbp_1 _4928_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net200),
    .D(_0208_),
    .Q_N(_2214_),
    .Q(\charlie_0.memory[11][4] ));
 sg13g2_dfrbp_1 _4929_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net196),
    .D(_0209_),
    .Q_N(_2213_),
    .Q(\charlie_0.memory[11][5] ));
 sg13g2_dfrbp_1 _4930_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net192),
    .D(_0210_),
    .Q_N(_2212_),
    .Q(\charlie_0.memory[11][6] ));
 sg13g2_dfrbp_1 _4931_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net188),
    .D(_0211_),
    .Q_N(_2211_),
    .Q(\charlie_0.memory[11][7] ));
 sg13g2_dfrbp_1 _4932_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net184),
    .D(_0212_),
    .Q_N(_2210_),
    .Q(\charlie_0.memory[12][0] ));
 sg13g2_dfrbp_1 _4933_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net180),
    .D(_0213_),
    .Q_N(_2209_),
    .Q(\charlie_0.memory[12][1] ));
 sg13g2_dfrbp_1 _4934_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net176),
    .D(_0214_),
    .Q_N(_2208_),
    .Q(\charlie_0.memory[12][2] ));
 sg13g2_dfrbp_1 _4935_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net172),
    .D(_0215_),
    .Q_N(_2207_),
    .Q(\charlie_0.memory[12][3] ));
 sg13g2_dfrbp_1 _4936_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net168),
    .D(_0216_),
    .Q_N(_2206_),
    .Q(\charlie_0.memory[12][4] ));
 sg13g2_dfrbp_1 _4937_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net164),
    .D(_0217_),
    .Q_N(_2205_),
    .Q(\charlie_0.memory[12][5] ));
 sg13g2_dfrbp_1 _4938_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net160),
    .D(_0218_),
    .Q_N(_2204_),
    .Q(\charlie_0.memory[12][6] ));
 sg13g2_dfrbp_1 _4939_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net156),
    .D(_0219_),
    .Q_N(_2203_),
    .Q(\charlie_0.memory[12][7] ));
 sg13g2_dfrbp_1 _4940_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net152),
    .D(_0220_),
    .Q_N(_2202_),
    .Q(\charlie_0.memory[13][0] ));
 sg13g2_dfrbp_1 _4941_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net148),
    .D(_0221_),
    .Q_N(_2201_),
    .Q(\charlie_0.memory[13][1] ));
 sg13g2_dfrbp_1 _4942_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net144),
    .D(_0222_),
    .Q_N(_2200_),
    .Q(\charlie_0.memory[13][2] ));
 sg13g2_dfrbp_1 _4943_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net140),
    .D(_0223_),
    .Q_N(_2199_),
    .Q(\charlie_0.memory[13][3] ));
 sg13g2_dfrbp_1 _4944_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net136),
    .D(_0224_),
    .Q_N(_2198_),
    .Q(\charlie_0.memory[13][4] ));
 sg13g2_dfrbp_1 _4945_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net132),
    .D(_0225_),
    .Q_N(_2197_),
    .Q(\charlie_0.memory[13][5] ));
 sg13g2_dfrbp_1 _4946_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net128),
    .D(_0226_),
    .Q_N(_2196_),
    .Q(\charlie_0.memory[13][6] ));
 sg13g2_dfrbp_1 _4947_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net124),
    .D(_0227_),
    .Q_N(_2195_),
    .Q(\charlie_0.memory[13][7] ));
 sg13g2_dfrbp_1 _4948_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net120),
    .D(_0228_),
    .Q_N(_2194_),
    .Q(\charlie_0.memory[14][0] ));
 sg13g2_dfrbp_1 _4949_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net116),
    .D(_0229_),
    .Q_N(_2193_),
    .Q(\charlie_0.memory[14][1] ));
 sg13g2_dfrbp_1 _4950_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net112),
    .D(_0230_),
    .Q_N(_2192_),
    .Q(\charlie_0.memory[14][2] ));
 sg13g2_dfrbp_1 _4951_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net108),
    .D(_0231_),
    .Q_N(_2191_),
    .Q(\charlie_0.memory[14][3] ));
 sg13g2_dfrbp_1 _4952_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net104),
    .D(_0232_),
    .Q_N(_2190_),
    .Q(\charlie_0.memory[14][4] ));
 sg13g2_dfrbp_1 _4953_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net100),
    .D(_0233_),
    .Q_N(_2189_),
    .Q(\charlie_0.memory[14][5] ));
 sg13g2_dfrbp_1 _4954_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net96),
    .D(_0234_),
    .Q_N(_2188_),
    .Q(\charlie_0.memory[14][6] ));
 sg13g2_dfrbp_1 _4955_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net92),
    .D(_0235_),
    .Q_N(_2187_),
    .Q(\charlie_0.memory[14][7] ));
 sg13g2_dfrbp_1 _4956_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net88),
    .D(_0236_),
    .Q_N(_2186_),
    .Q(\charlie_0.memory[15][0] ));
 sg13g2_dfrbp_1 _4957_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net84),
    .D(_0237_),
    .Q_N(_2185_),
    .Q(\charlie_0.memory[15][1] ));
 sg13g2_dfrbp_1 _4958_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net80),
    .D(_0238_),
    .Q_N(_2184_),
    .Q(\charlie_0.memory[15][2] ));
 sg13g2_dfrbp_1 _4959_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net76),
    .D(_0239_),
    .Q_N(_2183_),
    .Q(\charlie_0.memory[15][3] ));
 sg13g2_dfrbp_1 _4960_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net72),
    .D(_0240_),
    .Q_N(_2182_),
    .Q(\charlie_0.memory[15][4] ));
 sg13g2_dfrbp_1 _4961_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net68),
    .D(_0241_),
    .Q_N(_2181_),
    .Q(\charlie_0.memory[15][5] ));
 sg13g2_dfrbp_1 _4962_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net64),
    .D(_0242_),
    .Q_N(_2180_),
    .Q(\charlie_0.memory[15][6] ));
 sg13g2_dfrbp_1 _4963_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net60),
    .D(_0243_),
    .Q_N(_2179_),
    .Q(\charlie_0.memory[15][7] ));
 sg13g2_dfrbp_1 _4964_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net8),
    .D(_0244_),
    .Q_N(_2178_),
    .Q(\charlie_0.memory[16][0] ));
 sg13g2_dfrbp_1 _4965_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net269),
    .D(_0245_),
    .Q_N(_2177_),
    .Q(\charlie_0.memory[16][1] ));
 sg13g2_dfrbp_1 _4966_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net264),
    .D(_0246_),
    .Q_N(_2176_),
    .Q(\charlie_0.memory[16][2] ));
 sg13g2_dfrbp_1 _4967_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net255),
    .D(_0247_),
    .Q_N(_0067_),
    .Q(\charlie_0.memory[16][3] ));
 sg13g2_dfrbp_1 _4968_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net247),
    .D(_0248_),
    .Q_N(_2175_),
    .Q(\charlie_0.memory[16][4] ));
 sg13g2_dfrbp_1 _4969_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net239),
    .D(_0249_),
    .Q_N(_2174_),
    .Q(\charlie_0.memory[16][5] ));
 sg13g2_dfrbp_1 _4970_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net231),
    .D(_0250_),
    .Q_N(_2173_),
    .Q(\charlie_0.memory[16][6] ));
 sg13g2_dfrbp_1 _4971_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net219),
    .D(_0251_),
    .Q_N(_2172_),
    .Q(\charlie_0.memory[16][7] ));
 sg13g2_dfrbp_1 _4972_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net211),
    .D(_0252_),
    .Q_N(_0048_),
    .Q(\charlie_0.memory[17][0] ));
 sg13g2_dfrbp_1 _4973_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net202),
    .D(_0253_),
    .Q_N(_2171_),
    .Q(\charlie_0.memory[17][1] ));
 sg13g2_dfrbp_1 _4974_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net194),
    .D(_0254_),
    .Q_N(_2170_),
    .Q(\charlie_0.memory[17][2] ));
 sg13g2_dfrbp_1 _4975_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net186),
    .D(_0255_),
    .Q_N(_2169_),
    .Q(\charlie_0.memory[17][3] ));
 sg13g2_dfrbp_1 _4976_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net178),
    .D(_0256_),
    .Q_N(_2168_),
    .Q(\charlie_0.memory[17][4] ));
 sg13g2_dfrbp_1 _4977_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net170),
    .D(_0257_),
    .Q_N(_2167_),
    .Q(\charlie_0.memory[17][5] ));
 sg13g2_dfrbp_1 _4978_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net162),
    .D(_0258_),
    .Q_N(_2166_),
    .Q(\charlie_0.memory[17][6] ));
 sg13g2_dfrbp_1 _4979_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net154),
    .D(_0259_),
    .Q_N(_2165_),
    .Q(\charlie_0.memory[17][7] ));
 sg13g2_dfrbp_1 _4980_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net146),
    .D(_0260_),
    .Q_N(_0050_),
    .Q(\charlie_0.memory[18][0] ));
 sg13g2_dfrbp_1 _4981_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net138),
    .D(_0261_),
    .Q_N(_2164_),
    .Q(\charlie_0.memory[18][1] ));
 sg13g2_dfrbp_1 _4982_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net130),
    .D(_0262_),
    .Q_N(_2163_),
    .Q(\charlie_0.memory[18][2] ));
 sg13g2_dfrbp_1 _4983_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net122),
    .D(_0263_),
    .Q_N(_2162_),
    .Q(\charlie_0.memory[18][3] ));
 sg13g2_dfrbp_1 _4984_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net114),
    .D(_0264_),
    .Q_N(_2161_),
    .Q(\charlie_0.memory[18][4] ));
 sg13g2_dfrbp_1 _4985_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net106),
    .D(_0265_),
    .Q_N(_2160_),
    .Q(\charlie_0.memory[18][5] ));
 sg13g2_dfrbp_1 _4986_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net98),
    .D(_0266_),
    .Q_N(_2159_),
    .Q(\charlie_0.memory[18][6] ));
 sg13g2_dfrbp_1 _4987_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net90),
    .D(_0267_),
    .Q_N(_2158_),
    .Q(\charlie_0.memory[18][7] ));
 sg13g2_dfrbp_1 _4988_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net82),
    .D(_0268_),
    .Q_N(_2157_),
    .Q(\bi_frame_index[0] ));
 sg13g2_dfrbp_1 _4989_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net74),
    .D(_0269_),
    .Q_N(_0064_),
    .Q(\bi_frame_index[1] ));
 sg13g2_dfrbp_1 _4990_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net66),
    .D(_0270_),
    .Q_N(_2156_),
    .Q(\charlie_0.is_mirror ));
 sg13g2_dfrbp_1 _4991_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net10),
    .D(_0271_),
    .Q_N(_2155_),
    .Q(\charlie_0.memory[19][3] ));
 sg13g2_dfrbp_1 _4992_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net267),
    .D(_0272_),
    .Q_N(_2154_),
    .Q(\charlie_0.memory[19][4] ));
 sg13g2_dfrbp_1 _4993_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net251),
    .D(_0273_),
    .Q_N(_2153_),
    .Q(\charlie_0.memory[19][5] ));
 sg13g2_dfrbp_1 _4994_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net235),
    .D(_0274_),
    .Q_N(_2152_),
    .Q(\charlie_0.memory[19][6] ));
 sg13g2_dfrbp_1 _4995_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net215),
    .D(_0275_),
    .Q_N(_2151_),
    .Q(\charlie_0.memory[19][7] ));
 sg13g2_dfrbp_1 _4996_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net198),
    .D(_0276_),
    .Q_N(_2150_),
    .Q(\charlie_0.memory[20][1] ));
 sg13g2_dfrbp_1 _4997_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net182),
    .D(_0277_),
    .Q_N(_2149_),
    .Q(\charlie_0.memory[20][4] ));
 sg13g2_dfrbp_1 _4998_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net166),
    .D(_0278_),
    .Q_N(_2148_),
    .Q(\charlie_0.memory[20][5] ));
 sg13g2_dfrbp_1 _4999_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net150),
    .D(_0279_),
    .Q_N(_2147_),
    .Q(\charlie_0.memory[20][6] ));
 sg13g2_dfrbp_1 _5000_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net134),
    .D(net300),
    .Q_N(_2146_),
    .Q(\charlie_0.memory[20][7] ));
 sg13g2_dfrbp_1 _5001_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net118),
    .D(net277),
    .Q_N(_0051_),
    .Q(\charlie_0.memory[21][0] ));
 sg13g2_dfrbp_1 _5002_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net102),
    .D(_0282_),
    .Q_N(_2145_),
    .Q(\charlie_0.memory[21][1] ));
 sg13g2_dfrbp_1 _5003_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net86),
    .D(_0283_),
    .Q_N(_2144_),
    .Q(\charlie_0.memory[21][2] ));
 sg13g2_dfrbp_1 _5004_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net70),
    .D(_0284_),
    .Q_N(_2143_),
    .Q(\charlie_0.memory[21][3] ));
 sg13g2_dfrbp_1 _5005_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net271),
    .D(_0285_),
    .Q_N(_2142_),
    .Q(\charlie_0.memory[21][4] ));
 sg13g2_dfrbp_1 _5006_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net243),
    .D(net359),
    .Q_N(_2141_),
    .Q(\charlie_0.memory[21][5] ));
 sg13g2_dfrbp_1 _5007_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net207),
    .D(net322),
    .Q_N(_2140_),
    .Q(\charlie_0.memory[21][6] ));
 sg13g2_dfrbp_1 _5008_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net174),
    .D(net311),
    .Q_N(_2139_),
    .Q(\charlie_0.memory[21][7] ));
 sg13g2_dfrbp_1 _5009_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net142),
    .D(_0289_),
    .Q_N(_2138_),
    .Q(\charlie_0.memory[20][3] ));
 sg13g2_dfrbp_1 _5010_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net110),
    .D(_0290_),
    .Q_N(_0054_),
    .Q(\charlie_0.memory[22][0] ));
 sg13g2_dfrbp_1 _5011_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net78),
    .D(_0291_),
    .Q_N(_0053_),
    .Q(\charlie_0.memory[22][1] ));
 sg13g2_dfrbp_1 _5012_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net259),
    .D(_0292_),
    .Q_N(_0052_),
    .Q(\charlie_0.memory[22][2] ));
 sg13g2_dfrbp_1 _5013_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net190),
    .D(_0293_),
    .Q_N(_2137_),
    .Q(\charlie_0.memory[22][3] ));
 sg13g2_dfrbp_1 _5014_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net126),
    .D(_0294_),
    .Q_N(_2136_),
    .Q(\charlie_0.memory[22][4] ));
 sg13g2_dfrbp_1 _5015_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net62),
    .D(_0295_),
    .Q_N(_2135_),
    .Q(\charlie_0.memory[22][5] ));
 sg13g2_dfrbp_1 _5016_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net158),
    .D(_0296_),
    .Q_N(_2134_),
    .Q(\charlie_0.memory[22][6] ));
 sg13g2_dfrbp_1 _5017_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net227),
    .D(_0297_),
    .Q_N(_2133_),
    .Q(\charlie_0.memory[22][7] ));
 sg13g2_tiehi _4909__9 (.L_HI(net9));
 sg13g2_tiehi _4991__10 (.L_HI(net10));
 sg13g2_tiehi _4753__11 (.L_HI(net11));
 sg13g2_tiehi _4755__12 (.L_HI(net12));
 sg13g2_tiehi _4756__13 (.L_HI(net13));
 sg13g2_tiehi _4757__14 (.L_HI(net14));
 sg13g2_tiehi _4758__15 (.L_HI(net15));
 sg13g2_tiehi _4759__16 (.L_HI(net16));
 sg13g2_tiehi _4760__17 (.L_HI(net17));
 sg13g2_tiehi _4761__18 (.L_HI(net18));
 sg13g2_tiehi _4762__19 (.L_HI(net19));
 sg13g2_tiehi _4763__20 (.L_HI(net20));
 sg13g2_tiehi _4764__21 (.L_HI(net21));
 sg13g2_tiehi _4765__22 (.L_HI(net22));
 sg13g2_tiehi _4766__23 (.L_HI(net23));
 sg13g2_tiehi _4767__24 (.L_HI(net24));
 sg13g2_tiehi _4768__25 (.L_HI(net25));
 sg13g2_tiehi _4769__26 (.L_HI(net26));
 sg13g2_tiehi _4770__27 (.L_HI(net27));
 sg13g2_tiehi _4771__28 (.L_HI(net28));
 sg13g2_tiehi _4772__29 (.L_HI(net29));
 sg13g2_tiehi _4773__30 (.L_HI(net30));
 sg13g2_tiehi _4774__31 (.L_HI(net31));
 sg13g2_tiehi _4775__32 (.L_HI(net32));
 sg13g2_tiehi _4776__33 (.L_HI(net33));
 sg13g2_tiehi _4777__34 (.L_HI(net34));
 sg13g2_tiehi _4778__35 (.L_HI(net35));
 sg13g2_tiehi _4779__36 (.L_HI(net36));
 sg13g2_tiehi _4780__37 (.L_HI(net37));
 sg13g2_tiehi _4781__38 (.L_HI(net38));
 sg13g2_tiehi _4782__39 (.L_HI(net39));
 sg13g2_tiehi _4783__40 (.L_HI(net40));
 sg13g2_tiehi _4784__41 (.L_HI(net41));
 sg13g2_tiehi _4785__42 (.L_HI(net42));
 sg13g2_tiehi _4786__43 (.L_HI(net43));
 sg13g2_tiehi _4787__44 (.L_HI(net44));
 sg13g2_tiehi _4788__45 (.L_HI(net45));
 sg13g2_tiehi _4789__46 (.L_HI(net46));
 sg13g2_tiehi _4790__47 (.L_HI(net47));
 sg13g2_tiehi _4791__48 (.L_HI(net48));
 sg13g2_tiehi _4792__49 (.L_HI(net49));
 sg13g2_tiehi _4793__50 (.L_HI(net50));
 sg13g2_tiehi _4794__51 (.L_HI(net51));
 sg13g2_tiehi _4795__52 (.L_HI(net52));
 sg13g2_tiehi _4796__53 (.L_HI(net53));
 sg13g2_tiehi _4797__54 (.L_HI(net54));
 sg13g2_tiehi _4798__55 (.L_HI(net55));
 sg13g2_tiehi _4799__56 (.L_HI(net56));
 sg13g2_tiehi _4800__57 (.L_HI(net57));
 sg13g2_tiehi _4801__58 (.L_HI(net58));
 sg13g2_tiehi _4908__59 (.L_HI(net59));
 sg13g2_tiehi _4963__60 (.L_HI(net60));
 sg13g2_tiehi _4907__61 (.L_HI(net61));
 sg13g2_tiehi _5015__62 (.L_HI(net62));
 sg13g2_tiehi _4906__63 (.L_HI(net63));
 sg13g2_tiehi _4962__64 (.L_HI(net64));
 sg13g2_tiehi _4905__65 (.L_HI(net65));
 sg13g2_tiehi _4990__66 (.L_HI(net66));
 sg13g2_tiehi _4904__67 (.L_HI(net67));
 sg13g2_tiehi _4961__68 (.L_HI(net68));
 sg13g2_tiehi _4903__69 (.L_HI(net69));
 sg13g2_tiehi _5004__70 (.L_HI(net70));
 sg13g2_tiehi _4902__71 (.L_HI(net71));
 sg13g2_tiehi _4960__72 (.L_HI(net72));
 sg13g2_tiehi _4901__73 (.L_HI(net73));
 sg13g2_tiehi _4989__74 (.L_HI(net74));
 sg13g2_tiehi _4900__75 (.L_HI(net75));
 sg13g2_tiehi _4959__76 (.L_HI(net76));
 sg13g2_tiehi _4899__77 (.L_HI(net77));
 sg13g2_tiehi _5011__78 (.L_HI(net78));
 sg13g2_tiehi _4898__79 (.L_HI(net79));
 sg13g2_tiehi _4958__80 (.L_HI(net80));
 sg13g2_tiehi _4897__81 (.L_HI(net81));
 sg13g2_tiehi _4988__82 (.L_HI(net82));
 sg13g2_tiehi _4896__83 (.L_HI(net83));
 sg13g2_tiehi _4957__84 (.L_HI(net84));
 sg13g2_tiehi _4895__85 (.L_HI(net85));
 sg13g2_tiehi _5003__86 (.L_HI(net86));
 sg13g2_tiehi _4894__87 (.L_HI(net87));
 sg13g2_tiehi _4956__88 (.L_HI(net88));
 sg13g2_tiehi _4893__89 (.L_HI(net89));
 sg13g2_tiehi _4987__90 (.L_HI(net90));
 sg13g2_tiehi _4892__91 (.L_HI(net91));
 sg13g2_tiehi _4955__92 (.L_HI(net92));
 sg13g2_tiehi _4891__93 (.L_HI(net93));
 sg13g2_tiehi _4802__94 (.L_HI(net94));
 sg13g2_tiehi _4890__95 (.L_HI(net95));
 sg13g2_tiehi _4954__96 (.L_HI(net96));
 sg13g2_tiehi _4889__97 (.L_HI(net97));
 sg13g2_tiehi _4986__98 (.L_HI(net98));
 sg13g2_tiehi _4888__99 (.L_HI(net99));
 sg13g2_tiehi _4953__100 (.L_HI(net100));
 sg13g2_tiehi _4887__101 (.L_HI(net101));
 sg13g2_tiehi _5002__102 (.L_HI(net102));
 sg13g2_tiehi _4886__103 (.L_HI(net103));
 sg13g2_tiehi _4952__104 (.L_HI(net104));
 sg13g2_tiehi _4885__105 (.L_HI(net105));
 sg13g2_tiehi _4985__106 (.L_HI(net106));
 sg13g2_tiehi _4884__107 (.L_HI(net107));
 sg13g2_tiehi _4951__108 (.L_HI(net108));
 sg13g2_tiehi _4883__109 (.L_HI(net109));
 sg13g2_tiehi _5010__110 (.L_HI(net110));
 sg13g2_tiehi _4882__111 (.L_HI(net111));
 sg13g2_tiehi _4950__112 (.L_HI(net112));
 sg13g2_tiehi _4881__113 (.L_HI(net113));
 sg13g2_tiehi _4984__114 (.L_HI(net114));
 sg13g2_tiehi _4880__115 (.L_HI(net115));
 sg13g2_tiehi _4949__116 (.L_HI(net116));
 sg13g2_tiehi _4879__117 (.L_HI(net117));
 sg13g2_tiehi _5001__118 (.L_HI(net118));
 sg13g2_tiehi _4878__119 (.L_HI(net119));
 sg13g2_tiehi _4948__120 (.L_HI(net120));
 sg13g2_tiehi _4877__121 (.L_HI(net121));
 sg13g2_tiehi _4983__122 (.L_HI(net122));
 sg13g2_tiehi _4876__123 (.L_HI(net123));
 sg13g2_tiehi _4947__124 (.L_HI(net124));
 sg13g2_tiehi _4875__125 (.L_HI(net125));
 sg13g2_tiehi _5014__126 (.L_HI(net126));
 sg13g2_tiehi _4874__127 (.L_HI(net127));
 sg13g2_tiehi _4946__128 (.L_HI(net128));
 sg13g2_tiehi _4873__129 (.L_HI(net129));
 sg13g2_tiehi _4982__130 (.L_HI(net130));
 sg13g2_tiehi _4872__131 (.L_HI(net131));
 sg13g2_tiehi _4945__132 (.L_HI(net132));
 sg13g2_tiehi _4871__133 (.L_HI(net133));
 sg13g2_tiehi _5000__134 (.L_HI(net134));
 sg13g2_tiehi _4870__135 (.L_HI(net135));
 sg13g2_tiehi _4944__136 (.L_HI(net136));
 sg13g2_tiehi _4869__137 (.L_HI(net137));
 sg13g2_tiehi _4981__138 (.L_HI(net138));
 sg13g2_tiehi _4868__139 (.L_HI(net139));
 sg13g2_tiehi _4943__140 (.L_HI(net140));
 sg13g2_tiehi _4867__141 (.L_HI(net141));
 sg13g2_tiehi _5009__142 (.L_HI(net142));
 sg13g2_tiehi _4866__143 (.L_HI(net143));
 sg13g2_tiehi _4942__144 (.L_HI(net144));
 sg13g2_tiehi _4865__145 (.L_HI(net145));
 sg13g2_tiehi _4980__146 (.L_HI(net146));
 sg13g2_tiehi _4864__147 (.L_HI(net147));
 sg13g2_tiehi _4941__148 (.L_HI(net148));
 sg13g2_tiehi _4863__149 (.L_HI(net149));
 sg13g2_tiehi _4999__150 (.L_HI(net150));
 sg13g2_tiehi _4862__151 (.L_HI(net151));
 sg13g2_tiehi _4940__152 (.L_HI(net152));
 sg13g2_tiehi _4861__153 (.L_HI(net153));
 sg13g2_tiehi _4979__154 (.L_HI(net154));
 sg13g2_tiehi _4860__155 (.L_HI(net155));
 sg13g2_tiehi _4939__156 (.L_HI(net156));
 sg13g2_tiehi _4859__157 (.L_HI(net157));
 sg13g2_tiehi _5016__158 (.L_HI(net158));
 sg13g2_tiehi _4858__159 (.L_HI(net159));
 sg13g2_tiehi _4938__160 (.L_HI(net160));
 sg13g2_tiehi _4857__161 (.L_HI(net161));
 sg13g2_tiehi _4978__162 (.L_HI(net162));
 sg13g2_tiehi _4856__163 (.L_HI(net163));
 sg13g2_tiehi _4937__164 (.L_HI(net164));
 sg13g2_tiehi _4855__165 (.L_HI(net165));
 sg13g2_tiehi _4998__166 (.L_HI(net166));
 sg13g2_tiehi _4854__167 (.L_HI(net167));
 sg13g2_tiehi _4936__168 (.L_HI(net168));
 sg13g2_tiehi _4853__169 (.L_HI(net169));
 sg13g2_tiehi _4977__170 (.L_HI(net170));
 sg13g2_tiehi _4852__171 (.L_HI(net171));
 sg13g2_tiehi _4935__172 (.L_HI(net172));
 sg13g2_tiehi _4851__173 (.L_HI(net173));
 sg13g2_tiehi _5008__174 (.L_HI(net174));
 sg13g2_tiehi _4850__175 (.L_HI(net175));
 sg13g2_tiehi _4934__176 (.L_HI(net176));
 sg13g2_tiehi _4849__177 (.L_HI(net177));
 sg13g2_tiehi _4976__178 (.L_HI(net178));
 sg13g2_tiehi _4848__179 (.L_HI(net179));
 sg13g2_tiehi _4933__180 (.L_HI(net180));
 sg13g2_tiehi _4847__181 (.L_HI(net181));
 sg13g2_tiehi _4997__182 (.L_HI(net182));
 sg13g2_tiehi _4846__183 (.L_HI(net183));
 sg13g2_tiehi _4932__184 (.L_HI(net184));
 sg13g2_tiehi _4845__185 (.L_HI(net185));
 sg13g2_tiehi _4975__186 (.L_HI(net186));
 sg13g2_tiehi _4844__187 (.L_HI(net187));
 sg13g2_tiehi _4931__188 (.L_HI(net188));
 sg13g2_tiehi _4843__189 (.L_HI(net189));
 sg13g2_tiehi _5013__190 (.L_HI(net190));
 sg13g2_tiehi _4842__191 (.L_HI(net191));
 sg13g2_tiehi _4930__192 (.L_HI(net192));
 sg13g2_tiehi _4841__193 (.L_HI(net193));
 sg13g2_tiehi _4974__194 (.L_HI(net194));
 sg13g2_tiehi _4840__195 (.L_HI(net195));
 sg13g2_tiehi _4929__196 (.L_HI(net196));
 sg13g2_tiehi _4839__197 (.L_HI(net197));
 sg13g2_tiehi _4996__198 (.L_HI(net198));
 sg13g2_tiehi _4838__199 (.L_HI(net199));
 sg13g2_tiehi _4928__200 (.L_HI(net200));
 sg13g2_tiehi _4837__201 (.L_HI(net201));
 sg13g2_tiehi _4973__202 (.L_HI(net202));
 sg13g2_tiehi _4836__203 (.L_HI(net203));
 sg13g2_tiehi _4835__204 (.L_HI(net204));
 sg13g2_tiehi _4927__205 (.L_HI(net205));
 sg13g2_tiehi _4834__206 (.L_HI(net206));
 sg13g2_tiehi _5007__207 (.L_HI(net207));
 sg13g2_tiehi _4833__208 (.L_HI(net208));
 sg13g2_tiehi _4926__209 (.L_HI(net209));
 sg13g2_tiehi _4832__210 (.L_HI(net210));
 sg13g2_tiehi _4972__211 (.L_HI(net211));
 sg13g2_tiehi _4831__212 (.L_HI(net212));
 sg13g2_tiehi _4925__213 (.L_HI(net213));
 sg13g2_tiehi _4830__214 (.L_HI(net214));
 sg13g2_tiehi _4995__215 (.L_HI(net215));
 sg13g2_tiehi _4829__216 (.L_HI(net216));
 sg13g2_tiehi _4924__217 (.L_HI(net217));
 sg13g2_tiehi _4828__218 (.L_HI(net218));
 sg13g2_tiehi _4971__219 (.L_HI(net219));
 sg13g2_tiehi _4827__220 (.L_HI(net220));
 sg13g2_tiehi _4826__221 (.L_HI(net221));
 sg13g2_tiehi _4825__222 (.L_HI(net222));
 sg13g2_tiehi _4923__223 (.L_HI(net223));
 sg13g2_tiehi _4824__224 (.L_HI(net224));
 sg13g2_tiehi _4823__225 (.L_HI(net225));
 sg13g2_tiehi _4822__226 (.L_HI(net226));
 sg13g2_tiehi _5017__227 (.L_HI(net227));
 sg13g2_tiehi _4821__228 (.L_HI(net228));
 sg13g2_tiehi _4922__229 (.L_HI(net229));
 sg13g2_tiehi _4820__230 (.L_HI(net230));
 sg13g2_tiehi _4970__231 (.L_HI(net231));
 sg13g2_tiehi _4819__232 (.L_HI(net232));
 sg13g2_tiehi _4921__233 (.L_HI(net233));
 sg13g2_tiehi _4818__234 (.L_HI(net234));
 sg13g2_tiehi _4994__235 (.L_HI(net235));
 sg13g2_tiehi _4817__236 (.L_HI(net236));
 sg13g2_tiehi _4920__237 (.L_HI(net237));
 sg13g2_tiehi _4816__238 (.L_HI(net238));
 sg13g2_tiehi _4969__239 (.L_HI(net239));
 sg13g2_tiehi _4815__240 (.L_HI(net240));
 sg13g2_tiehi _4919__241 (.L_HI(net241));
 sg13g2_tiehi _4814__242 (.L_HI(net242));
 sg13g2_tiehi _5006__243 (.L_HI(net243));
 sg13g2_tiehi _4813__244 (.L_HI(net244));
 sg13g2_tiehi _4918__245 (.L_HI(net245));
 sg13g2_tiehi _4812__246 (.L_HI(net246));
 sg13g2_tiehi _4968__247 (.L_HI(net247));
 sg13g2_tiehi _4811__248 (.L_HI(net248));
 sg13g2_tiehi _4917__249 (.L_HI(net249));
 sg13g2_tiehi _4810__250 (.L_HI(net250));
 sg13g2_tiehi _4993__251 (.L_HI(net251));
 sg13g2_tiehi _4809__252 (.L_HI(net252));
 sg13g2_tiehi _4916__253 (.L_HI(net253));
 sg13g2_tiehi _4808__254 (.L_HI(net254));
 sg13g2_tiehi _4967__255 (.L_HI(net255));
 sg13g2_tiehi _4807__256 (.L_HI(net256));
 sg13g2_tiehi _4915__257 (.L_HI(net257));
 sg13g2_tiehi _4806__258 (.L_HI(net258));
 sg13g2_tiehi _5012__259 (.L_HI(net259));
 sg13g2_tiehi _4805__260 (.L_HI(net260));
 sg13g2_tiehi _4914__261 (.L_HI(net261));
 sg13g2_tiehi _4804__262 (.L_HI(net262));
 sg13g2_tiehi _4803__263 (.L_HI(net263));
 sg13g2_tiehi _4966__264 (.L_HI(net264));
 sg13g2_tiehi _4754__265 (.L_HI(net265));
 sg13g2_tiehi _4913__266 (.L_HI(net266));
 sg13g2_tiehi _4992__267 (.L_HI(net267));
 sg13g2_tiehi _4912__268 (.L_HI(net268));
 sg13g2_tiehi _4965__269 (.L_HI(net269));
 sg13g2_tiehi _4911__270 (.L_HI(net270));
 sg13g2_tiehi _5005__271 (.L_HI(net271));
 sg13g2_tiehi _4910__272 (.L_HI(net272));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_buf_1 _5283_ (.A(miso),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout952 (.A(_0499_),
    .X(net952));
 sg13g2_buf_2 fanout953 (.A(net954),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(_0798_),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(net956),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(_1759_),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(_1728_),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(net959),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(_1711_),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(_1702_),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(_1702_),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(net963),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(_1693_),
    .X(net963));
 sg13g2_buf_4 fanout964 (.X(net964),
    .A(net965));
 sg13g2_buf_2 fanout965 (.A(_1684_),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(net967),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(_1651_),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(_1618_),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(_1618_),
    .X(net969));
 sg13g2_buf_2 fanout970 (.A(net971),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(_1585_),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(_1550_),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(_1550_),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(net976),
    .X(net974));
 sg13g2_buf_1 fanout975 (.A(net976),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(_1517_),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(net978),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(_1484_),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(net980),
    .X(net979));
 sg13g2_buf_2 fanout980 (.A(_1422_),
    .X(net980));
 sg13g2_buf_2 fanout981 (.A(net983),
    .X(net981));
 sg13g2_buf_1 fanout982 (.A(net983),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(_1412_),
    .X(net983));
 sg13g2_buf_2 fanout984 (.A(net985),
    .X(net984));
 sg13g2_buf_2 fanout985 (.A(_1402_),
    .X(net985));
 sg13g2_buf_2 fanout986 (.A(_1392_),
    .X(net986));
 sg13g2_buf_2 fanout987 (.A(_1392_),
    .X(net987));
 sg13g2_buf_2 fanout988 (.A(_1382_),
    .X(net988));
 sg13g2_buf_2 fanout989 (.A(_1382_),
    .X(net989));
 sg13g2_buf_2 fanout990 (.A(net991),
    .X(net990));
 sg13g2_buf_2 fanout991 (.A(_1373_),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(net993),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(_1362_),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(net995),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(_1351_),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(net997),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(_1340_),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(_0575_),
    .X(net998));
 sg13g2_buf_1 fanout999 (.A(_0575_),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(net1001),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(_1458_),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(_0778_),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(net1004),
    .X(net1003));
 sg13g2_buf_2 fanout1004 (.A(_1552_),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(net1006),
    .X(net1005));
 sg13g2_buf_2 fanout1006 (.A(_1552_),
    .X(net1006));
 sg13g2_buf_2 fanout1007 (.A(net1008),
    .X(net1007));
 sg13g2_buf_2 fanout1008 (.A(_1551_),
    .X(net1008));
 sg13g2_buf_2 fanout1009 (.A(net1010),
    .X(net1009));
 sg13g2_buf_2 fanout1010 (.A(net1011),
    .X(net1010));
 sg13g2_buf_2 fanout1011 (.A(_1551_),
    .X(net1011));
 sg13g2_buf_2 fanout1012 (.A(net1014),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(net1014),
    .X(net1013));
 sg13g2_buf_4 fanout1014 (.X(net1014),
    .A(_1424_));
 sg13g2_buf_2 fanout1015 (.A(net1016),
    .X(net1015));
 sg13g2_buf_4 fanout1016 (.X(net1016),
    .A(_1423_));
 sg13g2_buf_4 fanout1017 (.X(net1017),
    .A(net1020));
 sg13g2_buf_1 fanout1018 (.A(net1019),
    .X(net1018));
 sg13g2_buf_2 fanout1019 (.A(net1020),
    .X(net1019));
 sg13g2_buf_2 fanout1020 (.A(_1423_),
    .X(net1020));
 sg13g2_buf_4 fanout1021 (.X(net1021),
    .A(_0564_));
 sg13g2_buf_2 fanout1022 (.A(net1023),
    .X(net1022));
 sg13g2_buf_2 fanout1023 (.A(_1979_),
    .X(net1023));
 sg13g2_buf_2 fanout1024 (.A(_0516_),
    .X(net1024));
 sg13g2_buf_1 fanout1025 (.A(_0516_),
    .X(net1025));
 sg13g2_buf_2 fanout1026 (.A(_0334_),
    .X(net1026));
 sg13g2_buf_2 fanout1027 (.A(net1028),
    .X(net1027));
 sg13g2_buf_2 fanout1028 (.A(_1850_),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(net1030),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(net1031),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(_1013_),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(net1034),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(net1034),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(_1013_),
    .X(net1034));
 sg13g2_buf_4 fanout1035 (.X(net1035),
    .A(_1012_));
 sg13g2_buf_2 fanout1036 (.A(net1037),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(net1040),
    .X(net1037));
 sg13g2_buf_2 fanout1038 (.A(net1039),
    .X(net1038));
 sg13g2_buf_4 fanout1039 (.X(net1039),
    .A(net1040));
 sg13g2_buf_4 fanout1040 (.X(net1040),
    .A(_1011_));
 sg13g2_buf_4 fanout1041 (.X(net1041),
    .A(net1042));
 sg13g2_buf_2 fanout1042 (.A(_1010_),
    .X(net1042));
 sg13g2_buf_2 fanout1043 (.A(net1045),
    .X(net1043));
 sg13g2_buf_2 fanout1044 (.A(net1045),
    .X(net1044));
 sg13g2_buf_4 fanout1045 (.X(net1045),
    .A(_1008_));
 sg13g2_buf_2 fanout1046 (.A(net1048),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(net1048),
    .X(net1047));
 sg13g2_buf_2 fanout1048 (.A(_1008_),
    .X(net1048));
 sg13g2_buf_4 fanout1049 (.X(net1049),
    .A(net1050));
 sg13g2_buf_2 fanout1050 (.A(_1007_),
    .X(net1050));
 sg13g2_buf_2 fanout1051 (.A(net1055),
    .X(net1051));
 sg13g2_buf_1 fanout1052 (.A(net1055),
    .X(net1052));
 sg13g2_buf_2 fanout1053 (.A(net1054),
    .X(net1053));
 sg13g2_buf_2 fanout1054 (.A(net1055),
    .X(net1054));
 sg13g2_buf_2 fanout1055 (.A(_0827_),
    .X(net1055));
 sg13g2_buf_2 fanout1056 (.A(net1057),
    .X(net1056));
 sg13g2_buf_2 fanout1057 (.A(net1060),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(net1059),
    .X(net1058));
 sg13g2_buf_2 fanout1059 (.A(net1060),
    .X(net1059));
 sg13g2_buf_2 fanout1060 (.A(_0825_),
    .X(net1060));
 sg13g2_buf_2 fanout1061 (.A(_0822_),
    .X(net1061));
 sg13g2_buf_2 fanout1062 (.A(_0822_),
    .X(net1062));
 sg13g2_buf_2 fanout1063 (.A(net1064),
    .X(net1063));
 sg13g2_buf_2 fanout1064 (.A(_0822_),
    .X(net1064));
 sg13g2_buf_2 fanout1065 (.A(net1069),
    .X(net1065));
 sg13g2_buf_1 fanout1066 (.A(net1069),
    .X(net1066));
 sg13g2_buf_2 fanout1067 (.A(net1068),
    .X(net1067));
 sg13g2_buf_2 fanout1068 (.A(net1069),
    .X(net1068));
 sg13g2_buf_2 fanout1069 (.A(_0819_),
    .X(net1069));
 sg13g2_buf_2 fanout1070 (.A(net1072),
    .X(net1070));
 sg13g2_buf_2 fanout1071 (.A(net1072),
    .X(net1071));
 sg13g2_buf_2 fanout1072 (.A(_0800_),
    .X(net1072));
 sg13g2_buf_2 fanout1073 (.A(net1075),
    .X(net1073));
 sg13g2_buf_2 fanout1074 (.A(net1075),
    .X(net1074));
 sg13g2_buf_2 fanout1075 (.A(_0800_),
    .X(net1075));
 sg13g2_buf_4 fanout1076 (.X(net1076),
    .A(net1077));
 sg13g2_buf_2 fanout1077 (.A(_0799_),
    .X(net1077));
 sg13g2_buf_2 fanout1078 (.A(net1079),
    .X(net1078));
 sg13g2_buf_1 fanout1079 (.A(_0520_),
    .X(net1079));
 sg13g2_buf_2 fanout1080 (.A(net1081),
    .X(net1080));
 sg13g2_buf_2 fanout1081 (.A(net1083),
    .X(net1081));
 sg13g2_buf_2 fanout1082 (.A(net1083),
    .X(net1082));
 sg13g2_buf_2 fanout1083 (.A(net1084),
    .X(net1083));
 sg13g2_buf_4 fanout1084 (.X(net1084),
    .A(_0519_));
 sg13g2_buf_2 fanout1085 (.A(_0518_),
    .X(net1085));
 sg13g2_buf_1 fanout1086 (.A(_0518_),
    .X(net1086));
 sg13g2_buf_2 fanout1087 (.A(net1088),
    .X(net1087));
 sg13g2_buf_2 fanout1088 (.A(net1089),
    .X(net1088));
 sg13g2_buf_4 fanout1089 (.X(net1089),
    .A(net1090));
 sg13g2_buf_2 fanout1090 (.A(net1091),
    .X(net1090));
 sg13g2_buf_4 fanout1091 (.X(net1091),
    .A(_0517_));
 sg13g2_buf_2 fanout1092 (.A(net1096),
    .X(net1092));
 sg13g2_buf_2 fanout1093 (.A(net1096),
    .X(net1093));
 sg13g2_buf_2 fanout1094 (.A(net1095),
    .X(net1094));
 sg13g2_buf_1 fanout1095 (.A(net1096),
    .X(net1095));
 sg13g2_buf_2 fanout1096 (.A(net1097),
    .X(net1096));
 sg13g2_buf_4 fanout1097 (.X(net1097),
    .A(_0515_));
 sg13g2_buf_2 fanout1098 (.A(_0513_),
    .X(net1098));
 sg13g2_buf_1 fanout1099 (.A(_0513_),
    .X(net1099));
 sg13g2_buf_2 fanout1100 (.A(net1101),
    .X(net1100));
 sg13g2_buf_2 fanout1101 (.A(net1102),
    .X(net1101));
 sg13g2_buf_1 fanout1102 (.A(net1103),
    .X(net1102));
 sg13g2_buf_4 fanout1103 (.X(net1103),
    .A(net1104));
 sg13g2_buf_2 fanout1104 (.A(_0512_),
    .X(net1104));
 sg13g2_buf_2 fanout1105 (.A(_2006_),
    .X(net1105));
 sg13g2_buf_2 fanout1106 (.A(net1107),
    .X(net1106));
 sg13g2_buf_2 fanout1107 (.A(net1108),
    .X(net1107));
 sg13g2_buf_2 fanout1108 (.A(net1111),
    .X(net1108));
 sg13g2_buf_2 fanout1109 (.A(net1110),
    .X(net1109));
 sg13g2_buf_1 fanout1110 (.A(net1111),
    .X(net1110));
 sg13g2_buf_1 fanout1111 (.A(net1112),
    .X(net1111));
 sg13g2_buf_2 fanout1112 (.A(_1839_),
    .X(net1112));
 sg13g2_buf_2 fanout1113 (.A(net1115),
    .X(net1113));
 sg13g2_buf_2 fanout1114 (.A(net1115),
    .X(net1114));
 sg13g2_buf_4 fanout1115 (.X(net1115),
    .A(net1117));
 sg13g2_buf_4 fanout1116 (.X(net1116),
    .A(net1117));
 sg13g2_buf_2 fanout1117 (.A(_1822_),
    .X(net1117));
 sg13g2_buf_4 fanout1118 (.X(net1118),
    .A(_1821_));
 sg13g2_buf_2 fanout1119 (.A(net1120),
    .X(net1119));
 sg13g2_buf_4 fanout1120 (.X(net1120),
    .A(_1785_));
 sg13g2_buf_2 fanout1121 (.A(net1124),
    .X(net1121));
 sg13g2_buf_4 fanout1122 (.X(net1122),
    .A(net1124));
 sg13g2_buf_2 fanout1123 (.A(net1124),
    .X(net1123));
 sg13g2_buf_2 fanout1124 (.A(_1782_),
    .X(net1124));
 sg13g2_buf_4 fanout1125 (.X(net1125),
    .A(net1126));
 sg13g2_buf_8 fanout1126 (.A(_1775_),
    .X(net1126));
 sg13g2_buf_4 fanout1127 (.X(net1127),
    .A(net1129));
 sg13g2_buf_4 fanout1128 (.X(net1128),
    .A(_1773_));
 sg13g2_buf_2 fanout1129 (.A(_1773_),
    .X(net1129));
 sg13g2_buf_4 fanout1130 (.X(net1130),
    .A(net1132));
 sg13g2_buf_4 fanout1131 (.X(net1131),
    .A(net1132));
 sg13g2_buf_2 fanout1132 (.A(_1773_),
    .X(net1132));
 sg13g2_buf_4 fanout1133 (.X(net1133),
    .A(net1135));
 sg13g2_buf_4 fanout1134 (.X(net1134),
    .A(net1135));
 sg13g2_buf_4 fanout1135 (.X(net1135),
    .A(_1772_));
 sg13g2_buf_4 fanout1136 (.X(net1136),
    .A(net1137));
 sg13g2_buf_2 fanout1137 (.A(net1139),
    .X(net1137));
 sg13g2_buf_4 fanout1138 (.X(net1138),
    .A(net1139));
 sg13g2_buf_4 fanout1139 (.X(net1139),
    .A(_1771_));
 sg13g2_buf_4 fanout1140 (.X(net1140),
    .A(net1141));
 sg13g2_buf_8 fanout1141 (.A(_1770_),
    .X(net1141));
 sg13g2_buf_4 fanout1142 (.X(net1142),
    .A(net1143));
 sg13g2_buf_8 fanout1143 (.A(_1769_),
    .X(net1143));
 sg13g2_buf_4 fanout1144 (.X(net1144),
    .A(net1145));
 sg13g2_buf_8 fanout1145 (.A(_1768_),
    .X(net1145));
 sg13g2_buf_2 fanout1146 (.A(net475),
    .X(net1146));
 sg13g2_buf_4 fanout1147 (.X(net1147),
    .A(net1148));
 sg13g2_buf_4 fanout1148 (.X(net1148),
    .A(\charlie_0.memory[19][4] ));
 sg13g2_buf_4 fanout1149 (.X(net1149),
    .A(net1150));
 sg13g2_buf_4 fanout1150 (.X(net1150),
    .A(net368));
 sg13g2_buf_4 fanout1151 (.X(net1151),
    .A(\charlie_0.is_mirror ));
 sg13g2_buf_4 fanout1152 (.X(net1152),
    .A(net1153));
 sg13g2_buf_2 fanout1153 (.A(net1154),
    .X(net1153));
 sg13g2_buf_2 fanout1154 (.A(net340),
    .X(net1154));
 sg13g2_buf_4 fanout1155 (.X(net1155),
    .A(\bi_frame_index[0] ));
 sg13g2_buf_4 fanout1156 (.X(net1156),
    .A(net467));
 sg13g2_buf_2 fanout1157 (.A(\charlie_0.memory[17][3] ),
    .X(net1157));
 sg13g2_buf_4 fanout1158 (.X(net1158),
    .A(net1160));
 sg13g2_buf_4 fanout1159 (.X(net1159),
    .A(net1160));
 sg13g2_buf_4 fanout1160 (.X(net1160),
    .A(\charlie_0.memory[17][2] ));
 sg13g2_buf_2 fanout1161 (.A(net1162),
    .X(net1161));
 sg13g2_buf_4 fanout1162 (.X(net1162),
    .A(\charlie_0.memory[17][1] ));
 sg13g2_buf_4 fanout1163 (.X(net1163),
    .A(net1164));
 sg13g2_buf_4 fanout1164 (.X(net1164),
    .A(net367));
 sg13g2_buf_2 fanout1165 (.A(net1168),
    .X(net1165));
 sg13g2_buf_2 fanout1166 (.A(net1168),
    .X(net1166));
 sg13g2_buf_2 fanout1167 (.A(net1168),
    .X(net1167));
 sg13g2_buf_2 fanout1168 (.A(net1169),
    .X(net1168));
 sg13g2_buf_4 fanout1169 (.X(net1169),
    .A(net343));
 sg13g2_buf_4 fanout1170 (.X(net1170),
    .A(net1171));
 sg13g2_buf_4 fanout1171 (.X(net1171),
    .A(\charlie_0.memory[16][1] ));
 sg13g2_buf_4 fanout1172 (.X(net1172),
    .A(net1173));
 sg13g2_buf_2 fanout1173 (.A(net1174),
    .X(net1173));
 sg13g2_buf_4 fanout1174 (.X(net1174),
    .A(\charlie_0.memory[16][0] ));
 sg13g2_buf_4 fanout1175 (.X(net1175),
    .A(\signal_generator_0.index_reg[4] ));
 sg13g2_buf_4 fanout1176 (.X(net1176),
    .A(net435));
 sg13g2_buf_4 fanout1177 (.X(net1177),
    .A(\signal_generator_0.index_reg[3] ));
 sg13g2_buf_4 fanout1178 (.X(net1178),
    .A(net1181));
 sg13g2_buf_4 fanout1179 (.X(net1179),
    .A(net1181));
 sg13g2_buf_1 fanout1180 (.A(net1181),
    .X(net1180));
 sg13g2_buf_2 fanout1181 (.A(\signal_generator_0.index_reg[2] ),
    .X(net1181));
 sg13g2_buf_2 fanout1182 (.A(net454),
    .X(net1182));
 sg13g2_buf_4 fanout1183 (.X(net1183),
    .A(\signal_generator_0.index_reg[0] ));
 sg13g2_buf_4 fanout1184 (.X(net1184),
    .A(net443));
 sg13g2_buf_4 fanout1185 (.X(net1185),
    .A(net443));
 sg13g2_buf_4 fanout1186 (.X(net1186),
    .A(net373));
 sg13g2_buf_2 fanout1187 (.A(net373),
    .X(net1187));
 sg13g2_buf_4 fanout1188 (.X(net1188),
    .A(net1189));
 sg13g2_buf_4 fanout1189 (.X(net1189),
    .A(net303));
 sg13g2_buf_4 fanout1190 (.X(net1190),
    .A(net485));
 sg13g2_buf_4 fanout1191 (.X(net1191),
    .A(net485));
 sg13g2_buf_2 fanout1192 (.A(net1193),
    .X(net1192));
 sg13g2_buf_4 fanout1193 (.X(net1193),
    .A(net1194));
 sg13g2_buf_4 fanout1194 (.X(net1194),
    .A(net474));
 sg13g2_buf_4 fanout1195 (.X(net1195),
    .A(net474));
 sg13g2_buf_2 fanout1196 (.A(\gen_priority_write_blocks[0].this_priority_write.data_bits[10] ),
    .X(net1196));
 sg13g2_buf_4 fanout1197 (.X(net1197),
    .A(net1199));
 sg13g2_buf_2 fanout1198 (.A(net1199),
    .X(net1198));
 sg13g2_buf_4 fanout1199 (.X(net1199),
    .A(net441));
 sg13g2_buf_2 fanout1200 (.A(net280),
    .X(net1200));
 sg13g2_buf_4 fanout1201 (.X(net1201),
    .A(net438));
 sg13g2_buf_2 fanout1202 (.A(\charlie_0.charlie_index[5] ),
    .X(net1202));
 sg13g2_buf_2 fanout1203 (.A(net1204),
    .X(net1203));
 sg13g2_buf_2 fanout1204 (.A(\charlie_0.charlie_index[4] ),
    .X(net1204));
 sg13g2_buf_2 fanout1205 (.A(net1206),
    .X(net1205));
 sg13g2_buf_4 fanout1206 (.X(net1206),
    .A(\charlie_0.charlie_index[3] ));
 sg13g2_buf_4 fanout1207 (.X(net1207),
    .A(net1208));
 sg13g2_buf_2 fanout1208 (.A(\charlie_0.charlie_index[2] ),
    .X(net1208));
 sg13g2_buf_4 fanout1209 (.X(net1209),
    .A(net1210));
 sg13g2_buf_4 fanout1210 (.X(net1210),
    .A(\charlie_0.charlie_index[1] ));
 sg13g2_buf_2 fanout1211 (.A(net1212),
    .X(net1211));
 sg13g2_buf_2 fanout1212 (.A(\charlie_0.charlie_index[0] ),
    .X(net1212));
 sg13g2_buf_4 fanout1213 (.X(net1213),
    .A(net413));
 sg13g2_buf_4 fanout1214 (.X(net1214),
    .A(net413));
 sg13g2_buf_2 fanout1215 (.A(net1216),
    .X(net1215));
 sg13g2_buf_2 fanout1216 (.A(net1224),
    .X(net1216));
 sg13g2_buf_2 fanout1217 (.A(net1224),
    .X(net1217));
 sg13g2_buf_2 fanout1218 (.A(net1220),
    .X(net1218));
 sg13g2_buf_2 fanout1219 (.A(net1220),
    .X(net1219));
 sg13g2_buf_2 fanout1220 (.A(net1221),
    .X(net1220));
 sg13g2_buf_2 fanout1221 (.A(net1224),
    .X(net1221));
 sg13g2_buf_2 fanout1222 (.A(net1223),
    .X(net1222));
 sg13g2_buf_4 fanout1223 (.X(net1223),
    .A(net1224));
 sg13g2_buf_2 fanout1224 (.A(net1227),
    .X(net1224));
 sg13g2_buf_2 fanout1225 (.A(net1226),
    .X(net1225));
 sg13g2_buf_4 fanout1226 (.X(net1226),
    .A(net1227));
 sg13g2_buf_2 fanout1227 (.A(_1835_),
    .X(net1227));
 sg13g2_buf_4 fanout1228 (.X(net1228),
    .A(net1230));
 sg13g2_buf_2 fanout1229 (.A(net1230),
    .X(net1229));
 sg13g2_buf_8 fanout1230 (.A(_1776_),
    .X(net1230));
 sg13g2_buf_4 fanout1231 (.X(net1231),
    .A(net1232));
 sg13g2_buf_4 fanout1232 (.X(net1232),
    .A(net1233));
 sg13g2_buf_4 fanout1233 (.X(net1233),
    .A(ui_in[2]));
 sg13g2_buf_2 fanout1234 (.A(net1236),
    .X(net1234));
 sg13g2_buf_2 fanout1235 (.A(net1236),
    .X(net1235));
 sg13g2_buf_2 fanout1236 (.A(net1241),
    .X(net1236));
 sg13g2_buf_2 fanout1237 (.A(net1241),
    .X(net1237));
 sg13g2_buf_2 fanout1238 (.A(net1241),
    .X(net1238));
 sg13g2_buf_2 fanout1239 (.A(net1241),
    .X(net1239));
 sg13g2_buf_2 fanout1240 (.A(net1241),
    .X(net1240));
 sg13g2_buf_2 fanout1241 (.A(net1242),
    .X(net1241));
 sg13g2_buf_4 fanout1242 (.X(net1242),
    .A(net1258));
 sg13g2_buf_2 fanout1243 (.A(net1250),
    .X(net1243));
 sg13g2_buf_2 fanout1244 (.A(net1250),
    .X(net1244));
 sg13g2_buf_2 fanout1245 (.A(net1247),
    .X(net1245));
 sg13g2_buf_2 fanout1246 (.A(net1248),
    .X(net1246));
 sg13g2_buf_1 fanout1247 (.A(net1248),
    .X(net1247));
 sg13g2_buf_2 fanout1248 (.A(net1250),
    .X(net1248));
 sg13g2_buf_2 fanout1249 (.A(net1250),
    .X(net1249));
 sg13g2_buf_2 fanout1250 (.A(net1258),
    .X(net1250));
 sg13g2_buf_2 fanout1251 (.A(net1253),
    .X(net1251));
 sg13g2_buf_2 fanout1252 (.A(net1253),
    .X(net1252));
 sg13g2_buf_2 fanout1253 (.A(net1258),
    .X(net1253));
 sg13g2_buf_2 fanout1254 (.A(net1256),
    .X(net1254));
 sg13g2_buf_1 fanout1255 (.A(net1256),
    .X(net1255));
 sg13g2_buf_2 fanout1256 (.A(net1257),
    .X(net1256));
 sg13g2_buf_2 fanout1257 (.A(net1258),
    .X(net1257));
 sg13g2_buf_2 fanout1258 (.A(rst_n),
    .X(net1258));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[4]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[5]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[6]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[7]),
    .X(net7));
 sg13g2_tiehi _4964__8 (.L_HI(net8));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_leaf_0_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_0_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_1_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_1_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_2_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_2_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_3_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_3_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_4_clk_regs (.A(clknet_3_1__leaf_clk_regs),
    .X(clknet_leaf_4_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_5_clk_regs (.A(clknet_3_3__leaf_clk_regs),
    .X(clknet_leaf_5_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_6_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_6_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_7_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_7_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_8_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_8_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_9_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_9_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_10_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_10_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_11_clk_regs (.A(clknet_3_3__leaf_clk_regs),
    .X(clknet_leaf_11_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_12_clk_regs (.A(clknet_3_3__leaf_clk_regs),
    .X(clknet_leaf_12_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_13_clk_regs (.A(clknet_3_6__leaf_clk_regs),
    .X(clknet_leaf_13_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_14_clk_regs (.A(clknet_3_3__leaf_clk_regs),
    .X(clknet_leaf_14_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_15_clk_regs (.A(clknet_3_6__leaf_clk_regs),
    .X(clknet_leaf_15_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_16_clk_regs (.A(clknet_3_6__leaf_clk_regs),
    .X(clknet_leaf_16_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_17_clk_regs (.A(clknet_3_6__leaf_clk_regs),
    .X(clknet_leaf_17_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_18_clk_regs (.A(clknet_3_7__leaf_clk_regs),
    .X(clknet_leaf_18_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_19_clk_regs (.A(clknet_3_7__leaf_clk_regs),
    .X(clknet_leaf_19_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_20_clk_regs (.A(clknet_3_7__leaf_clk_regs),
    .X(clknet_leaf_20_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_21_clk_regs (.A(clknet_3_5__leaf_clk_regs),
    .X(clknet_leaf_21_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_22_clk_regs (.A(clknet_3_7__leaf_clk_regs),
    .X(clknet_leaf_22_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_24_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_24_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_25_clk_regs (.A(clknet_3_5__leaf_clk_regs),
    .X(clknet_leaf_25_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_26_clk_regs (.A(clknet_3_5__leaf_clk_regs),
    .X(clknet_leaf_26_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_27_clk_regs (.A(clknet_3_5__leaf_clk_regs),
    .X(clknet_leaf_27_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_28_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_28_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_29_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_29_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_30_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_30_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_31_clk_regs (.A(clknet_3_1__leaf_clk_regs),
    .X(clknet_leaf_31_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_32_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_32_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_33_clk_regs (.A(clknet_3_1__leaf_clk_regs),
    .X(clknet_leaf_33_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_34_clk_regs (.A(clknet_3_1__leaf_clk_regs),
    .X(clknet_leaf_34_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_35_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_35_clk_regs));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_3_0__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_1__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_1__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_2__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_2__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_3__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_3__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_4__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_4__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_5__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_5__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_6__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_6__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_7__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_7__leaf_clk_regs));
 sg13g2_buf_1 clkload0 (.A(clknet_3_0__leaf_clk_regs));
 sg13g2_inv_1 clkload1 (.A(clknet_3_1__leaf_clk_regs));
 sg13g2_buf_1 clkload2 (.A(clknet_3_2__leaf_clk_regs));
 sg13g2_inv_1 clkload3 (.A(clknet_3_3__leaf_clk_regs));
 sg13g2_buf_1 clkload4 (.A(clknet_3_4__leaf_clk_regs));
 sg13g2_inv_1 clkload5 (.A(clknet_3_5__leaf_clk_regs));
 sg13g2_inv_1 clkload6 (.A(clknet_3_7__leaf_clk_regs));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_14_clk_regs));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_24_clk_regs));
 sg13g2_inv_2 clkload9 (.A(clknet_leaf_28_clk_regs));
 sg13g2_inv_2 clkload10 (.A(clknet_leaf_30_clk_regs));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_18_clk_regs));
 sg13g2_inv_4 clkload12 (.A(clknet_leaf_22_clk_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0077_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0080_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0098_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0051_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0281_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0048_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0107_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0063_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0309_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0076_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold11 (.A(_1723_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold12 (.A(\spi_slave_0.reg_data[7] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0101_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold14 (.A(\spi_slave_0.is_mosi ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0097_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0078_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0082_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0079_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold19 (.A(_1721_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold20 (.A(\spi_slave_0.bit_cnt[1] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0790_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0099_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0075_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold24 (.A(\spi_slave_0.bit_cnt[2] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0792_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0100_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0066_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0280_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0066_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0775_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold31 (.A(\gen_priority_write_blocks[0].this_priority_write.data_bits[12] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0068_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold33 (.A(\spi_slave_0.is_data_phase ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0817_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0069_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold36 (.A(\signal_generator_0.index_reg[6] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold37 (.A(\charlie_0.memory[19][5] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold38 (.A(\charlie_0.memory[21][7] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0288_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold40 (.A(\charlie_0.memory[0][1] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold41 (.A(\spi_address[4] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold42 (.A(\charlie_0.memory[16][7] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold43 (.A(\charlie_0.is_mirror ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold44 (.A(\charlie_0.memory[0][6] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold45 (.A(\charlie_0.memory[0][4] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold46 (.A(\charlie_0.memory[0][0] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold47 (.A(\signal_generator_0.index_reg[5] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold48 (.A(\charlie_0.memory[21][6] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold49 (.A(_1751_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0287_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold51 (.A(\charlie_0.memory[22][2] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold52 (.A(\charlie_0.memory[0][5] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold53 (.A(\charlie_0.memory[2][7] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold54 (.A(\bi_frame_index[0] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold55 (.A(\charlie_0.memory[0][3] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold56 (.A(\charlie_0.memory[2][4] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold57 (.A(\charlie_0.memory[0][7] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold58 (.A(\charlie_0.memory[0][2] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold59 (.A(\spi_address[3] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold60 (.A(\charlie_0.memory[19][6] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold61 (.A(\counter[8] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0046_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold63 (.A(\spi_address[0] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold64 (.A(\charlie_0.memory[7][5] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold65 (.A(\charlie_0.memory[2][6] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold66 (.A(\signal_generator_0.state_machine[1] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0103_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold68 (.A(\bi_frame_index[1] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold69 (.A(\charlie_0.memory[20][6] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold70 (.A(\spi_address[1] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold71 (.A(\charlie_0.memory[16][6] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold72 (.A(_1892_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0019_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold74 (.A(\spi_address[2] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold75 (.A(\counter[13] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0021_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold77 (.A(\charlie_0.memory[5][0] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold78 (.A(\charlie_0.memory[7][7] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold79 (.A(\charlie_0.memory[19][7] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold80 (.A(\charlie_0.memory[4][4] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold81 (.A(\counter[25] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0034_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold83 (.A(\counter[6] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold84 (.A(\charlie_0.memory[6][7] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold85 (.A(\charlie_0.memory[17][7] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold86 (.A(\charlie_0.memory[21][5] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0286_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold88 (.A(\counter[14] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0022_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold90 (.A(\charlie_0.memory[7][4] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold91 (.A(\charlie_0.memory[16][4] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold92 (.A(\charlie_0.memory[6][0] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold93 (.A(\charlie_0.memory[3][0] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold94 (.A(\charlie_0.memory[22][3] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold95 (.A(\charlie_0.memory[17][0] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold96 (.A(\charlie_0.memory[19][3] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold97 (.A(\counter[29] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0039_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold99 (.A(\charlie_0.memory[4][0] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold100 (.A(\charlie_0.memory[5][1] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold101 (.A(\gen_priority_write_blocks[0].this_priority_write.data_bits[13] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold102 (.A(\charlie_0.memory[7][2] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold103 (.A(\charlie_0.memory[7][0] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold104 (.A(\counter[10] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold105 (.A(_1884_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0017_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold107 (.A(\counter[23] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0032_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold109 (.A(\charlie_0.memory[5][4] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold110 (.A(\charlie_0.memory[6][4] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold111 (.A(sig_gen_out),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0105_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold113 (.A(\charlie_0.memory[2][5] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold114 (.A(\charlie_0.memory[22][7] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold115 (.A(\charlie_0.memory[5][7] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold116 (.A(\charlie_0.memory[22][4] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold117 (.A(\charlie_0.memory[4][7] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold118 (.A(\charlie_0.memory[18][2] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold119 (.A(\charlie_0.memory[3][6] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold120 (.A(\charlie_0.memory[1][2] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold121 (.A(\charlie_0.memory[1][7] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold122 (.A(\charlie_0.memory[3][1] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold123 (.A(\charlie_0.memory[3][7] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold124 (.A(\counter[27] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0036_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold126 (.A(\charlie_0.memory[1][0] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold127 (.A(\charlie_0.memory[5][5] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold128 (.A(\charlie_0.memory[3][5] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold129 (.A(\charlie_0.memory[1][1] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold130 (.A(\charlie_0.memory[6][2] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold131 (.A(\counter[18] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold132 (.A(_1911_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0025_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold134 (.A(\counter[28] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold135 (.A(\charlie_0.memory[2][0] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold136 (.A(\counter[20] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold137 (.A(_1921_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0028_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0071_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold140 (.A(_1457_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold141 (.A(\gen_priority_write_blocks[0].this_priority_write.data_bits[15] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold142 (.A(\charlie_0.memory[18][4] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold143 (.A(\charlie_0.memory[5][3] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold144 (.A(\charlie_0.memory[4][3] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold145 (.A(\charlie_0.memory[4][6] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold146 (.A(\charlie_0.memory[7][3] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold147 (.A(\counter[15] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold148 (.A(\charlie_0.memory[6][6] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold149 (.A(\counter[22] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold150 (.A(\charlie_0.memory[1][5] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold151 (.A(\charlie_0.memory[6][1] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold152 (.A(\charlie_0.memory[4][2] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold153 (.A(\charlie_0.memory[1][4] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold154 (.A(\charlie_0.memory[2][2] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold155 (.A(\charlie_0.memory[3][3] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold156 (.A(\charlie_0.memory[5][2] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold157 (.A(\charlie_0.memory[2][3] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold158 (.A(\counter[7] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold159 (.A(\charlie_0.memory[2][1] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold160 (.A(\charlie_0.memory[22][6] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold161 (.A(\charlie_0.memory[18][7] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold162 (.A(\charlie_0.memory[5][6] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold163 (.A(\signal_generator_0.index_reg[4] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0111_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold165 (.A(\charlie_0.memory[4][1] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold166 (.A(\charlie_0.charlie_index[5] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0073_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold168 (.A(\counter[13] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold169 (.A(\gen_priority_write_blocks[0].this_priority_write.data_bits[9] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold170 (.A(\charlie_0.memory[1][3] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold171 (.A(\gen_priority_write_blocks[0].this_priority_write.data_bits[14] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold172 (.A(\charlie_0.memory[10][7] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold173 (.A(_1515_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold174 (.A(\charlie_0.memory[4][5] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold175 (.A(\charlie_0.memory[6][5] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold176 (.A(\charlie_0.memory[3][2] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold177 (.A(\charlie_0.memory[7][1] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold178 (.A(\charlie_0.memory[6][3] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold179 (.A(\signal_generator_0.index_reg[7] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold180 (.A(\counter[30] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold181 (.A(\charlie_0.memory[3][4] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold182 (.A(\signal_generator_0.index_reg[1] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold183 (.A(\charlie_0.memory[22][5] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0072_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold185 (.A(\charlie_0.memory[18][1] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold186 (.A(\charlie_0.memory[18][0] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold187 (.A(\charlie_0.memory[16][2] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold188 (.A(\charlie_0.memory[7][6] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold189 (.A(\charlie_0.memory[1][6] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold190 (.A(\charlie_0.memory[18][5] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold191 (.A(\charlie_0.memory[16][5] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold192 (.A(\counter[7] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold193 (.A(\counter[16] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold194 (.A(\charlie_0.memory[20][5] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold195 (.A(\charlie_0.memory[17][3] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold196 (.A(\charlie_0.memory[17][5] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold197 (.A(\charlie_0.memory[18][6] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold198 (.A(\counter[20] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold199 (.A(_1637_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold200 (.A(\counter[9] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold201 (.A(\charlie_0.memory[18][3] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold202 (.A(\gen_priority_write_blocks[0].this_priority_write.data_bits[10] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold203 (.A(\charlie_0.memory[22][0] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold204 (.A(\counter[12] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold205 (.A(_1603_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold206 (.A(\counter[30] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold207 (.A(\charlie_0.memory[10][0] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold208 (.A(_1487_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold209 (.A(\charlie_0.memory[22][1] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold210 (.A(\counter[18] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold211 (.A(\counter[10] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold212 (.A(_1595_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold213 (.A(\gen_priority_write_blocks[0].this_priority_write.data_bits[11] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold214 (.A(\counter[11] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold215 (.A(\counter[24] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold216 (.A(\counter[20] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold217 (.A(\charlie_0.memory[15][3] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold218 (.A(\charlie_0.memory[10][1] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold219 (.A(\charlie_0.memory[16][3] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold220 (.A(\counter[11] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold221 (.A(\counter[7] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold222 (.A(\counter[16] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold223 (.A(\counter[24] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold224 (.A(\counter[24] ),
    .X(net496));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_decap_8 FILLER_13_588 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_decap_8 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_637 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_8 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_decap_8 FILLER_13_798 ();
 sg13g2_decap_8 FILLER_13_805 ();
 sg13g2_decap_8 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_833 ();
 sg13g2_decap_8 FILLER_13_840 ();
 sg13g2_decap_8 FILLER_13_847 ();
 sg13g2_decap_8 FILLER_13_854 ();
 sg13g2_fill_1 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_8 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_511 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_574 ();
 sg13g2_decap_8 FILLER_14_581 ();
 sg13g2_decap_8 FILLER_14_588 ();
 sg13g2_decap_8 FILLER_14_595 ();
 sg13g2_decap_8 FILLER_14_602 ();
 sg13g2_decap_8 FILLER_14_609 ();
 sg13g2_decap_8 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_623 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_decap_8 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_decap_8 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_658 ();
 sg13g2_decap_8 FILLER_14_665 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_decap_8 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_decap_8 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_14_840 ();
 sg13g2_decap_8 FILLER_14_847 ();
 sg13g2_decap_8 FILLER_14_854 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_434 ();
 sg13g2_decap_8 FILLER_15_441 ();
 sg13g2_decap_8 FILLER_15_448 ();
 sg13g2_decap_8 FILLER_15_455 ();
 sg13g2_decap_8 FILLER_15_462 ();
 sg13g2_decap_8 FILLER_15_469 ();
 sg13g2_decap_8 FILLER_15_476 ();
 sg13g2_decap_8 FILLER_15_483 ();
 sg13g2_decap_8 FILLER_15_490 ();
 sg13g2_decap_8 FILLER_15_497 ();
 sg13g2_decap_8 FILLER_15_504 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_518 ();
 sg13g2_decap_8 FILLER_15_525 ();
 sg13g2_decap_8 FILLER_15_532 ();
 sg13g2_decap_8 FILLER_15_539 ();
 sg13g2_decap_8 FILLER_15_546 ();
 sg13g2_decap_8 FILLER_15_553 ();
 sg13g2_decap_8 FILLER_15_560 ();
 sg13g2_decap_8 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_574 ();
 sg13g2_decap_8 FILLER_15_581 ();
 sg13g2_decap_8 FILLER_15_588 ();
 sg13g2_decap_8 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_602 ();
 sg13g2_decap_8 FILLER_15_609 ();
 sg13g2_decap_8 FILLER_15_616 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_8 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_644 ();
 sg13g2_decap_8 FILLER_15_651 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_decap_8 FILLER_15_665 ();
 sg13g2_decap_8 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_679 ();
 sg13g2_decap_8 FILLER_15_686 ();
 sg13g2_decap_8 FILLER_15_693 ();
 sg13g2_decap_8 FILLER_15_700 ();
 sg13g2_decap_8 FILLER_15_707 ();
 sg13g2_decap_8 FILLER_15_714 ();
 sg13g2_decap_8 FILLER_15_721 ();
 sg13g2_decap_8 FILLER_15_728 ();
 sg13g2_decap_8 FILLER_15_735 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_decap_8 FILLER_15_749 ();
 sg13g2_decap_8 FILLER_15_756 ();
 sg13g2_decap_8 FILLER_15_763 ();
 sg13g2_decap_8 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_777 ();
 sg13g2_decap_8 FILLER_15_784 ();
 sg13g2_decap_8 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_798 ();
 sg13g2_decap_8 FILLER_15_805 ();
 sg13g2_decap_8 FILLER_15_812 ();
 sg13g2_decap_8 FILLER_15_819 ();
 sg13g2_decap_8 FILLER_15_826 ();
 sg13g2_decap_8 FILLER_15_833 ();
 sg13g2_decap_8 FILLER_15_840 ();
 sg13g2_decap_8 FILLER_15_847 ();
 sg13g2_decap_8 FILLER_15_854 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_8 FILLER_16_455 ();
 sg13g2_decap_8 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_469 ();
 sg13g2_decap_8 FILLER_16_476 ();
 sg13g2_decap_8 FILLER_16_483 ();
 sg13g2_decap_8 FILLER_16_490 ();
 sg13g2_decap_8 FILLER_16_497 ();
 sg13g2_decap_8 FILLER_16_504 ();
 sg13g2_decap_8 FILLER_16_511 ();
 sg13g2_decap_8 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_525 ();
 sg13g2_decap_8 FILLER_16_532 ();
 sg13g2_decap_8 FILLER_16_539 ();
 sg13g2_decap_8 FILLER_16_546 ();
 sg13g2_decap_8 FILLER_16_553 ();
 sg13g2_decap_8 FILLER_16_560 ();
 sg13g2_decap_8 FILLER_16_567 ();
 sg13g2_decap_8 FILLER_16_574 ();
 sg13g2_decap_8 FILLER_16_581 ();
 sg13g2_decap_8 FILLER_16_588 ();
 sg13g2_decap_8 FILLER_16_595 ();
 sg13g2_decap_8 FILLER_16_602 ();
 sg13g2_decap_8 FILLER_16_609 ();
 sg13g2_decap_8 FILLER_16_616 ();
 sg13g2_decap_8 FILLER_16_623 ();
 sg13g2_decap_8 FILLER_16_630 ();
 sg13g2_decap_8 FILLER_16_637 ();
 sg13g2_decap_8 FILLER_16_644 ();
 sg13g2_decap_8 FILLER_16_651 ();
 sg13g2_decap_8 FILLER_16_658 ();
 sg13g2_decap_8 FILLER_16_665 ();
 sg13g2_decap_8 FILLER_16_672 ();
 sg13g2_decap_8 FILLER_16_679 ();
 sg13g2_decap_8 FILLER_16_686 ();
 sg13g2_decap_8 FILLER_16_693 ();
 sg13g2_decap_8 FILLER_16_700 ();
 sg13g2_decap_8 FILLER_16_707 ();
 sg13g2_decap_8 FILLER_16_714 ();
 sg13g2_decap_8 FILLER_16_721 ();
 sg13g2_decap_8 FILLER_16_728 ();
 sg13g2_decap_8 FILLER_16_735 ();
 sg13g2_decap_8 FILLER_16_742 ();
 sg13g2_decap_8 FILLER_16_749 ();
 sg13g2_decap_8 FILLER_16_756 ();
 sg13g2_decap_8 FILLER_16_763 ();
 sg13g2_decap_8 FILLER_16_770 ();
 sg13g2_decap_8 FILLER_16_777 ();
 sg13g2_decap_8 FILLER_16_784 ();
 sg13g2_decap_8 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_798 ();
 sg13g2_decap_8 FILLER_16_805 ();
 sg13g2_decap_8 FILLER_16_812 ();
 sg13g2_decap_8 FILLER_16_819 ();
 sg13g2_decap_8 FILLER_16_826 ();
 sg13g2_decap_8 FILLER_16_833 ();
 sg13g2_decap_8 FILLER_16_840 ();
 sg13g2_decap_8 FILLER_16_847 ();
 sg13g2_decap_8 FILLER_16_854 ();
 sg13g2_fill_1 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_427 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_448 ();
 sg13g2_decap_8 FILLER_17_455 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_497 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_fill_1 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_decap_8 FILLER_18_427 ();
 sg13g2_decap_8 FILLER_18_434 ();
 sg13g2_decap_8 FILLER_18_441 ();
 sg13g2_decap_8 FILLER_18_448 ();
 sg13g2_decap_8 FILLER_18_455 ();
 sg13g2_decap_8 FILLER_18_462 ();
 sg13g2_decap_8 FILLER_18_469 ();
 sg13g2_decap_8 FILLER_18_476 ();
 sg13g2_decap_8 FILLER_18_483 ();
 sg13g2_decap_8 FILLER_18_490 ();
 sg13g2_decap_8 FILLER_18_497 ();
 sg13g2_decap_8 FILLER_18_504 ();
 sg13g2_decap_8 FILLER_18_511 ();
 sg13g2_decap_8 FILLER_18_518 ();
 sg13g2_decap_8 FILLER_18_525 ();
 sg13g2_decap_8 FILLER_18_532 ();
 sg13g2_decap_8 FILLER_18_539 ();
 sg13g2_decap_8 FILLER_18_546 ();
 sg13g2_decap_8 FILLER_18_553 ();
 sg13g2_decap_8 FILLER_18_560 ();
 sg13g2_decap_8 FILLER_18_567 ();
 sg13g2_decap_8 FILLER_18_574 ();
 sg13g2_decap_8 FILLER_18_581 ();
 sg13g2_decap_8 FILLER_18_588 ();
 sg13g2_decap_8 FILLER_18_595 ();
 sg13g2_decap_8 FILLER_18_602 ();
 sg13g2_decap_8 FILLER_18_609 ();
 sg13g2_decap_8 FILLER_18_616 ();
 sg13g2_decap_8 FILLER_18_623 ();
 sg13g2_decap_8 FILLER_18_630 ();
 sg13g2_decap_8 FILLER_18_637 ();
 sg13g2_decap_8 FILLER_18_644 ();
 sg13g2_decap_8 FILLER_18_651 ();
 sg13g2_decap_8 FILLER_18_658 ();
 sg13g2_decap_8 FILLER_18_665 ();
 sg13g2_decap_8 FILLER_18_672 ();
 sg13g2_decap_8 FILLER_18_679 ();
 sg13g2_decap_8 FILLER_18_686 ();
 sg13g2_decap_8 FILLER_18_693 ();
 sg13g2_decap_8 FILLER_18_700 ();
 sg13g2_decap_8 FILLER_18_707 ();
 sg13g2_decap_8 FILLER_18_714 ();
 sg13g2_decap_8 FILLER_18_721 ();
 sg13g2_decap_8 FILLER_18_728 ();
 sg13g2_decap_8 FILLER_18_735 ();
 sg13g2_decap_8 FILLER_18_742 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_decap_8 FILLER_18_756 ();
 sg13g2_decap_8 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_770 ();
 sg13g2_decap_8 FILLER_18_777 ();
 sg13g2_decap_8 FILLER_18_784 ();
 sg13g2_decap_8 FILLER_18_791 ();
 sg13g2_decap_8 FILLER_18_798 ();
 sg13g2_decap_8 FILLER_18_805 ();
 sg13g2_decap_8 FILLER_18_812 ();
 sg13g2_decap_8 FILLER_18_819 ();
 sg13g2_decap_8 FILLER_18_826 ();
 sg13g2_decap_8 FILLER_18_833 ();
 sg13g2_decap_8 FILLER_18_840 ();
 sg13g2_decap_8 FILLER_18_847 ();
 sg13g2_decap_8 FILLER_18_854 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_decap_8 FILLER_19_427 ();
 sg13g2_decap_8 FILLER_19_434 ();
 sg13g2_decap_8 FILLER_19_441 ();
 sg13g2_decap_8 FILLER_19_448 ();
 sg13g2_decap_8 FILLER_19_455 ();
 sg13g2_decap_8 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_490 ();
 sg13g2_decap_8 FILLER_19_497 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_532 ();
 sg13g2_decap_8 FILLER_19_539 ();
 sg13g2_decap_8 FILLER_19_546 ();
 sg13g2_decap_8 FILLER_19_553 ();
 sg13g2_decap_8 FILLER_19_560 ();
 sg13g2_decap_8 FILLER_19_567 ();
 sg13g2_decap_8 FILLER_19_574 ();
 sg13g2_decap_8 FILLER_19_581 ();
 sg13g2_decap_8 FILLER_19_588 ();
 sg13g2_decap_8 FILLER_19_595 ();
 sg13g2_decap_8 FILLER_19_602 ();
 sg13g2_decap_8 FILLER_19_609 ();
 sg13g2_decap_8 FILLER_19_616 ();
 sg13g2_decap_8 FILLER_19_623 ();
 sg13g2_decap_8 FILLER_19_630 ();
 sg13g2_decap_8 FILLER_19_637 ();
 sg13g2_decap_8 FILLER_19_644 ();
 sg13g2_decap_8 FILLER_19_651 ();
 sg13g2_decap_8 FILLER_19_658 ();
 sg13g2_decap_8 FILLER_19_665 ();
 sg13g2_decap_8 FILLER_19_672 ();
 sg13g2_decap_8 FILLER_19_679 ();
 sg13g2_decap_8 FILLER_19_686 ();
 sg13g2_decap_8 FILLER_19_693 ();
 sg13g2_decap_8 FILLER_19_700 ();
 sg13g2_decap_8 FILLER_19_707 ();
 sg13g2_decap_8 FILLER_19_714 ();
 sg13g2_decap_8 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_784 ();
 sg13g2_decap_8 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_798 ();
 sg13g2_decap_8 FILLER_19_805 ();
 sg13g2_decap_8 FILLER_19_812 ();
 sg13g2_decap_8 FILLER_19_819 ();
 sg13g2_decap_8 FILLER_19_826 ();
 sg13g2_decap_8 FILLER_19_833 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_decap_8 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_854 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_decap_8 FILLER_20_427 ();
 sg13g2_decap_8 FILLER_20_434 ();
 sg13g2_decap_8 FILLER_20_441 ();
 sg13g2_decap_8 FILLER_20_448 ();
 sg13g2_decap_8 FILLER_20_455 ();
 sg13g2_decap_8 FILLER_20_462 ();
 sg13g2_decap_8 FILLER_20_469 ();
 sg13g2_decap_8 FILLER_20_476 ();
 sg13g2_decap_8 FILLER_20_483 ();
 sg13g2_decap_8 FILLER_20_490 ();
 sg13g2_decap_8 FILLER_20_497 ();
 sg13g2_decap_8 FILLER_20_504 ();
 sg13g2_decap_8 FILLER_20_511 ();
 sg13g2_decap_8 FILLER_20_518 ();
 sg13g2_decap_8 FILLER_20_525 ();
 sg13g2_decap_8 FILLER_20_532 ();
 sg13g2_decap_8 FILLER_20_539 ();
 sg13g2_decap_8 FILLER_20_546 ();
 sg13g2_decap_8 FILLER_20_553 ();
 sg13g2_decap_8 FILLER_20_560 ();
 sg13g2_decap_8 FILLER_20_567 ();
 sg13g2_decap_8 FILLER_20_574 ();
 sg13g2_decap_8 FILLER_20_581 ();
 sg13g2_decap_8 FILLER_20_588 ();
 sg13g2_decap_8 FILLER_20_595 ();
 sg13g2_decap_8 FILLER_20_602 ();
 sg13g2_decap_8 FILLER_20_609 ();
 sg13g2_decap_8 FILLER_20_616 ();
 sg13g2_decap_8 FILLER_20_623 ();
 sg13g2_decap_8 FILLER_20_630 ();
 sg13g2_decap_8 FILLER_20_637 ();
 sg13g2_decap_8 FILLER_20_644 ();
 sg13g2_decap_8 FILLER_20_651 ();
 sg13g2_decap_8 FILLER_20_658 ();
 sg13g2_decap_8 FILLER_20_665 ();
 sg13g2_decap_8 FILLER_20_672 ();
 sg13g2_decap_8 FILLER_20_679 ();
 sg13g2_decap_8 FILLER_20_686 ();
 sg13g2_decap_8 FILLER_20_693 ();
 sg13g2_decap_8 FILLER_20_700 ();
 sg13g2_decap_8 FILLER_20_707 ();
 sg13g2_decap_8 FILLER_20_714 ();
 sg13g2_decap_8 FILLER_20_721 ();
 sg13g2_decap_8 FILLER_20_728 ();
 sg13g2_decap_8 FILLER_20_735 ();
 sg13g2_decap_8 FILLER_20_742 ();
 sg13g2_decap_8 FILLER_20_749 ();
 sg13g2_decap_8 FILLER_20_756 ();
 sg13g2_decap_8 FILLER_20_763 ();
 sg13g2_decap_8 FILLER_20_770 ();
 sg13g2_decap_8 FILLER_20_777 ();
 sg13g2_decap_8 FILLER_20_784 ();
 sg13g2_decap_8 FILLER_20_791 ();
 sg13g2_decap_8 FILLER_20_798 ();
 sg13g2_decap_8 FILLER_20_805 ();
 sg13g2_decap_8 FILLER_20_812 ();
 sg13g2_decap_8 FILLER_20_819 ();
 sg13g2_decap_8 FILLER_20_826 ();
 sg13g2_decap_8 FILLER_20_833 ();
 sg13g2_decap_8 FILLER_20_840 ();
 sg13g2_decap_8 FILLER_20_847 ();
 sg13g2_decap_8 FILLER_20_854 ();
 sg13g2_fill_1 FILLER_20_861 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_decap_8 FILLER_21_427 ();
 sg13g2_decap_8 FILLER_21_434 ();
 sg13g2_decap_8 FILLER_21_441 ();
 sg13g2_decap_8 FILLER_21_448 ();
 sg13g2_decap_8 FILLER_21_455 ();
 sg13g2_decap_8 FILLER_21_462 ();
 sg13g2_decap_8 FILLER_21_469 ();
 sg13g2_decap_8 FILLER_21_476 ();
 sg13g2_decap_8 FILLER_21_483 ();
 sg13g2_decap_8 FILLER_21_490 ();
 sg13g2_decap_8 FILLER_21_497 ();
 sg13g2_decap_8 FILLER_21_504 ();
 sg13g2_decap_8 FILLER_21_511 ();
 sg13g2_decap_8 FILLER_21_518 ();
 sg13g2_decap_8 FILLER_21_525 ();
 sg13g2_decap_8 FILLER_21_532 ();
 sg13g2_decap_8 FILLER_21_539 ();
 sg13g2_decap_8 FILLER_21_546 ();
 sg13g2_decap_8 FILLER_21_553 ();
 sg13g2_decap_8 FILLER_21_560 ();
 sg13g2_decap_8 FILLER_21_567 ();
 sg13g2_decap_8 FILLER_21_574 ();
 sg13g2_decap_8 FILLER_21_581 ();
 sg13g2_decap_8 FILLER_21_588 ();
 sg13g2_decap_8 FILLER_21_595 ();
 sg13g2_decap_8 FILLER_21_602 ();
 sg13g2_decap_8 FILLER_21_609 ();
 sg13g2_decap_8 FILLER_21_616 ();
 sg13g2_decap_8 FILLER_21_623 ();
 sg13g2_decap_8 FILLER_21_630 ();
 sg13g2_decap_8 FILLER_21_637 ();
 sg13g2_decap_8 FILLER_21_644 ();
 sg13g2_decap_8 FILLER_21_651 ();
 sg13g2_decap_8 FILLER_21_658 ();
 sg13g2_decap_8 FILLER_21_665 ();
 sg13g2_decap_8 FILLER_21_672 ();
 sg13g2_decap_8 FILLER_21_679 ();
 sg13g2_decap_8 FILLER_21_686 ();
 sg13g2_decap_8 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_700 ();
 sg13g2_decap_8 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_714 ();
 sg13g2_decap_8 FILLER_21_721 ();
 sg13g2_decap_8 FILLER_21_728 ();
 sg13g2_decap_8 FILLER_21_735 ();
 sg13g2_decap_8 FILLER_21_742 ();
 sg13g2_decap_8 FILLER_21_749 ();
 sg13g2_decap_8 FILLER_21_756 ();
 sg13g2_decap_8 FILLER_21_763 ();
 sg13g2_decap_8 FILLER_21_770 ();
 sg13g2_decap_8 FILLER_21_777 ();
 sg13g2_decap_8 FILLER_21_784 ();
 sg13g2_decap_8 FILLER_21_791 ();
 sg13g2_decap_8 FILLER_21_798 ();
 sg13g2_decap_8 FILLER_21_805 ();
 sg13g2_decap_8 FILLER_21_812 ();
 sg13g2_decap_8 FILLER_21_819 ();
 sg13g2_decap_8 FILLER_21_826 ();
 sg13g2_decap_8 FILLER_21_833 ();
 sg13g2_decap_8 FILLER_21_840 ();
 sg13g2_decap_8 FILLER_21_847 ();
 sg13g2_decap_8 FILLER_21_854 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_22_406 ();
 sg13g2_decap_8 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_decap_8 FILLER_22_427 ();
 sg13g2_decap_8 FILLER_22_434 ();
 sg13g2_decap_8 FILLER_22_441 ();
 sg13g2_decap_8 FILLER_22_448 ();
 sg13g2_decap_8 FILLER_22_455 ();
 sg13g2_decap_8 FILLER_22_462 ();
 sg13g2_decap_8 FILLER_22_469 ();
 sg13g2_decap_8 FILLER_22_476 ();
 sg13g2_decap_8 FILLER_22_483 ();
 sg13g2_decap_8 FILLER_22_490 ();
 sg13g2_decap_8 FILLER_22_497 ();
 sg13g2_decap_8 FILLER_22_504 ();
 sg13g2_decap_8 FILLER_22_511 ();
 sg13g2_decap_8 FILLER_22_518 ();
 sg13g2_decap_8 FILLER_22_525 ();
 sg13g2_decap_8 FILLER_22_532 ();
 sg13g2_decap_8 FILLER_22_539 ();
 sg13g2_decap_8 FILLER_22_546 ();
 sg13g2_decap_8 FILLER_22_553 ();
 sg13g2_decap_8 FILLER_22_560 ();
 sg13g2_decap_8 FILLER_22_567 ();
 sg13g2_decap_8 FILLER_22_574 ();
 sg13g2_decap_8 FILLER_22_581 ();
 sg13g2_decap_8 FILLER_22_588 ();
 sg13g2_decap_8 FILLER_22_595 ();
 sg13g2_decap_8 FILLER_22_602 ();
 sg13g2_decap_8 FILLER_22_609 ();
 sg13g2_decap_8 FILLER_22_616 ();
 sg13g2_decap_8 FILLER_22_623 ();
 sg13g2_decap_8 FILLER_22_630 ();
 sg13g2_decap_8 FILLER_22_637 ();
 sg13g2_decap_8 FILLER_22_644 ();
 sg13g2_decap_8 FILLER_22_651 ();
 sg13g2_decap_8 FILLER_22_658 ();
 sg13g2_decap_8 FILLER_22_665 ();
 sg13g2_decap_8 FILLER_22_672 ();
 sg13g2_decap_8 FILLER_22_679 ();
 sg13g2_decap_8 FILLER_22_686 ();
 sg13g2_decap_8 FILLER_22_693 ();
 sg13g2_decap_8 FILLER_22_700 ();
 sg13g2_decap_8 FILLER_22_707 ();
 sg13g2_decap_8 FILLER_22_714 ();
 sg13g2_decap_8 FILLER_22_721 ();
 sg13g2_decap_8 FILLER_22_728 ();
 sg13g2_decap_8 FILLER_22_735 ();
 sg13g2_decap_8 FILLER_22_742 ();
 sg13g2_decap_8 FILLER_22_749 ();
 sg13g2_decap_8 FILLER_22_756 ();
 sg13g2_decap_8 FILLER_22_763 ();
 sg13g2_decap_8 FILLER_22_770 ();
 sg13g2_decap_8 FILLER_22_777 ();
 sg13g2_decap_8 FILLER_22_784 ();
 sg13g2_decap_8 FILLER_22_791 ();
 sg13g2_decap_8 FILLER_22_798 ();
 sg13g2_decap_8 FILLER_22_805 ();
 sg13g2_decap_8 FILLER_22_812 ();
 sg13g2_decap_8 FILLER_22_819 ();
 sg13g2_decap_8 FILLER_22_826 ();
 sg13g2_decap_8 FILLER_22_833 ();
 sg13g2_decap_8 FILLER_22_840 ();
 sg13g2_decap_8 FILLER_22_847 ();
 sg13g2_decap_8 FILLER_22_854 ();
 sg13g2_fill_1 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_decap_8 FILLER_23_406 ();
 sg13g2_decap_8 FILLER_23_413 ();
 sg13g2_decap_8 FILLER_23_420 ();
 sg13g2_decap_8 FILLER_23_427 ();
 sg13g2_decap_8 FILLER_23_434 ();
 sg13g2_decap_8 FILLER_23_441 ();
 sg13g2_decap_8 FILLER_23_448 ();
 sg13g2_decap_8 FILLER_23_455 ();
 sg13g2_decap_8 FILLER_23_462 ();
 sg13g2_decap_8 FILLER_23_469 ();
 sg13g2_decap_8 FILLER_23_476 ();
 sg13g2_decap_8 FILLER_23_483 ();
 sg13g2_decap_8 FILLER_23_490 ();
 sg13g2_decap_8 FILLER_23_497 ();
 sg13g2_decap_8 FILLER_23_504 ();
 sg13g2_decap_8 FILLER_23_511 ();
 sg13g2_decap_8 FILLER_23_518 ();
 sg13g2_decap_8 FILLER_23_525 ();
 sg13g2_decap_8 FILLER_23_532 ();
 sg13g2_decap_8 FILLER_23_539 ();
 sg13g2_decap_8 FILLER_23_546 ();
 sg13g2_decap_8 FILLER_23_553 ();
 sg13g2_decap_8 FILLER_23_560 ();
 sg13g2_decap_8 FILLER_23_567 ();
 sg13g2_decap_8 FILLER_23_574 ();
 sg13g2_decap_8 FILLER_23_581 ();
 sg13g2_decap_8 FILLER_23_588 ();
 sg13g2_decap_8 FILLER_23_595 ();
 sg13g2_decap_8 FILLER_23_602 ();
 sg13g2_decap_8 FILLER_23_609 ();
 sg13g2_decap_8 FILLER_23_616 ();
 sg13g2_decap_8 FILLER_23_623 ();
 sg13g2_decap_8 FILLER_23_630 ();
 sg13g2_decap_8 FILLER_23_637 ();
 sg13g2_decap_8 FILLER_23_644 ();
 sg13g2_decap_8 FILLER_23_651 ();
 sg13g2_decap_8 FILLER_23_658 ();
 sg13g2_decap_8 FILLER_23_665 ();
 sg13g2_decap_8 FILLER_23_672 ();
 sg13g2_decap_8 FILLER_23_679 ();
 sg13g2_decap_8 FILLER_23_686 ();
 sg13g2_decap_8 FILLER_23_693 ();
 sg13g2_decap_8 FILLER_23_700 ();
 sg13g2_decap_8 FILLER_23_707 ();
 sg13g2_decap_8 FILLER_23_714 ();
 sg13g2_decap_8 FILLER_23_721 ();
 sg13g2_decap_8 FILLER_23_728 ();
 sg13g2_decap_8 FILLER_23_735 ();
 sg13g2_decap_8 FILLER_23_742 ();
 sg13g2_decap_8 FILLER_23_749 ();
 sg13g2_decap_8 FILLER_23_756 ();
 sg13g2_decap_8 FILLER_23_763 ();
 sg13g2_decap_8 FILLER_23_770 ();
 sg13g2_decap_8 FILLER_23_777 ();
 sg13g2_decap_8 FILLER_23_784 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_798 ();
 sg13g2_decap_8 FILLER_23_805 ();
 sg13g2_decap_8 FILLER_23_812 ();
 sg13g2_decap_8 FILLER_23_819 ();
 sg13g2_decap_8 FILLER_23_826 ();
 sg13g2_decap_8 FILLER_23_833 ();
 sg13g2_decap_8 FILLER_23_840 ();
 sg13g2_decap_8 FILLER_23_847 ();
 sg13g2_decap_8 FILLER_23_854 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_decap_8 FILLER_24_406 ();
 sg13g2_decap_8 FILLER_24_413 ();
 sg13g2_decap_8 FILLER_24_420 ();
 sg13g2_decap_8 FILLER_24_427 ();
 sg13g2_decap_8 FILLER_24_434 ();
 sg13g2_decap_8 FILLER_24_441 ();
 sg13g2_decap_8 FILLER_24_448 ();
 sg13g2_decap_8 FILLER_24_455 ();
 sg13g2_decap_8 FILLER_24_462 ();
 sg13g2_decap_8 FILLER_24_469 ();
 sg13g2_decap_8 FILLER_24_476 ();
 sg13g2_decap_8 FILLER_24_483 ();
 sg13g2_decap_8 FILLER_24_490 ();
 sg13g2_decap_8 FILLER_24_497 ();
 sg13g2_decap_8 FILLER_24_504 ();
 sg13g2_decap_8 FILLER_24_511 ();
 sg13g2_decap_8 FILLER_24_518 ();
 sg13g2_decap_8 FILLER_24_525 ();
 sg13g2_decap_8 FILLER_24_532 ();
 sg13g2_decap_8 FILLER_24_539 ();
 sg13g2_decap_8 FILLER_24_546 ();
 sg13g2_decap_8 FILLER_24_553 ();
 sg13g2_decap_8 FILLER_24_560 ();
 sg13g2_decap_8 FILLER_24_567 ();
 sg13g2_decap_8 FILLER_24_574 ();
 sg13g2_decap_8 FILLER_24_581 ();
 sg13g2_decap_8 FILLER_24_588 ();
 sg13g2_decap_8 FILLER_24_595 ();
 sg13g2_decap_8 FILLER_24_602 ();
 sg13g2_decap_8 FILLER_24_609 ();
 sg13g2_decap_8 FILLER_24_616 ();
 sg13g2_decap_8 FILLER_24_623 ();
 sg13g2_decap_8 FILLER_24_630 ();
 sg13g2_decap_8 FILLER_24_637 ();
 sg13g2_decap_8 FILLER_24_644 ();
 sg13g2_decap_8 FILLER_24_651 ();
 sg13g2_decap_8 FILLER_24_658 ();
 sg13g2_decap_8 FILLER_24_665 ();
 sg13g2_decap_8 FILLER_24_672 ();
 sg13g2_decap_8 FILLER_24_679 ();
 sg13g2_decap_8 FILLER_24_686 ();
 sg13g2_decap_8 FILLER_24_693 ();
 sg13g2_decap_8 FILLER_24_700 ();
 sg13g2_decap_8 FILLER_24_707 ();
 sg13g2_decap_8 FILLER_24_714 ();
 sg13g2_decap_8 FILLER_24_721 ();
 sg13g2_decap_8 FILLER_24_728 ();
 sg13g2_decap_8 FILLER_24_735 ();
 sg13g2_decap_8 FILLER_24_742 ();
 sg13g2_decap_8 FILLER_24_749 ();
 sg13g2_decap_8 FILLER_24_756 ();
 sg13g2_decap_8 FILLER_24_763 ();
 sg13g2_decap_8 FILLER_24_770 ();
 sg13g2_decap_8 FILLER_24_777 ();
 sg13g2_decap_8 FILLER_24_784 ();
 sg13g2_decap_8 FILLER_24_791 ();
 sg13g2_decap_8 FILLER_24_798 ();
 sg13g2_decap_8 FILLER_24_805 ();
 sg13g2_decap_8 FILLER_24_812 ();
 sg13g2_decap_8 FILLER_24_819 ();
 sg13g2_decap_8 FILLER_24_826 ();
 sg13g2_decap_8 FILLER_24_833 ();
 sg13g2_decap_8 FILLER_24_840 ();
 sg13g2_decap_8 FILLER_24_847 ();
 sg13g2_decap_8 FILLER_24_854 ();
 sg13g2_fill_1 FILLER_24_861 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_decap_8 FILLER_25_406 ();
 sg13g2_decap_8 FILLER_25_413 ();
 sg13g2_decap_8 FILLER_25_420 ();
 sg13g2_decap_8 FILLER_25_427 ();
 sg13g2_decap_8 FILLER_25_434 ();
 sg13g2_decap_8 FILLER_25_441 ();
 sg13g2_decap_8 FILLER_25_448 ();
 sg13g2_decap_8 FILLER_25_455 ();
 sg13g2_decap_8 FILLER_25_462 ();
 sg13g2_decap_8 FILLER_25_469 ();
 sg13g2_decap_8 FILLER_25_476 ();
 sg13g2_decap_8 FILLER_25_483 ();
 sg13g2_decap_8 FILLER_25_490 ();
 sg13g2_decap_8 FILLER_25_497 ();
 sg13g2_decap_8 FILLER_25_504 ();
 sg13g2_decap_8 FILLER_25_511 ();
 sg13g2_decap_8 FILLER_25_518 ();
 sg13g2_decap_8 FILLER_25_525 ();
 sg13g2_decap_8 FILLER_25_532 ();
 sg13g2_decap_8 FILLER_25_539 ();
 sg13g2_decap_8 FILLER_25_546 ();
 sg13g2_decap_8 FILLER_25_553 ();
 sg13g2_decap_8 FILLER_25_560 ();
 sg13g2_decap_8 FILLER_25_567 ();
 sg13g2_decap_8 FILLER_25_574 ();
 sg13g2_decap_8 FILLER_25_581 ();
 sg13g2_decap_8 FILLER_25_588 ();
 sg13g2_decap_8 FILLER_25_595 ();
 sg13g2_decap_8 FILLER_25_602 ();
 sg13g2_decap_8 FILLER_25_609 ();
 sg13g2_decap_8 FILLER_25_616 ();
 sg13g2_decap_8 FILLER_25_623 ();
 sg13g2_decap_8 FILLER_25_630 ();
 sg13g2_decap_8 FILLER_25_637 ();
 sg13g2_decap_8 FILLER_25_644 ();
 sg13g2_decap_8 FILLER_25_651 ();
 sg13g2_decap_8 FILLER_25_658 ();
 sg13g2_decap_8 FILLER_25_665 ();
 sg13g2_decap_8 FILLER_25_672 ();
 sg13g2_decap_8 FILLER_25_679 ();
 sg13g2_decap_8 FILLER_25_686 ();
 sg13g2_decap_8 FILLER_25_693 ();
 sg13g2_decap_8 FILLER_25_700 ();
 sg13g2_decap_8 FILLER_25_707 ();
 sg13g2_decap_8 FILLER_25_714 ();
 sg13g2_decap_8 FILLER_25_721 ();
 sg13g2_decap_8 FILLER_25_728 ();
 sg13g2_decap_8 FILLER_25_735 ();
 sg13g2_decap_8 FILLER_25_742 ();
 sg13g2_decap_8 FILLER_25_749 ();
 sg13g2_decap_8 FILLER_25_756 ();
 sg13g2_decap_8 FILLER_25_763 ();
 sg13g2_decap_8 FILLER_25_770 ();
 sg13g2_decap_8 FILLER_25_777 ();
 sg13g2_decap_8 FILLER_25_784 ();
 sg13g2_decap_8 FILLER_25_791 ();
 sg13g2_decap_8 FILLER_25_798 ();
 sg13g2_decap_8 FILLER_25_805 ();
 sg13g2_decap_8 FILLER_25_812 ();
 sg13g2_decap_8 FILLER_25_819 ();
 sg13g2_decap_8 FILLER_25_826 ();
 sg13g2_decap_8 FILLER_25_833 ();
 sg13g2_decap_8 FILLER_25_840 ();
 sg13g2_decap_8 FILLER_25_847 ();
 sg13g2_decap_8 FILLER_25_854 ();
 sg13g2_fill_1 FILLER_25_861 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_decap_8 FILLER_26_406 ();
 sg13g2_decap_8 FILLER_26_413 ();
 sg13g2_decap_8 FILLER_26_420 ();
 sg13g2_decap_8 FILLER_26_427 ();
 sg13g2_decap_8 FILLER_26_434 ();
 sg13g2_decap_8 FILLER_26_441 ();
 sg13g2_decap_8 FILLER_26_448 ();
 sg13g2_decap_8 FILLER_26_455 ();
 sg13g2_decap_8 FILLER_26_462 ();
 sg13g2_decap_8 FILLER_26_469 ();
 sg13g2_decap_8 FILLER_26_476 ();
 sg13g2_decap_8 FILLER_26_483 ();
 sg13g2_decap_8 FILLER_26_490 ();
 sg13g2_decap_8 FILLER_26_497 ();
 sg13g2_decap_8 FILLER_26_504 ();
 sg13g2_decap_8 FILLER_26_511 ();
 sg13g2_decap_8 FILLER_26_518 ();
 sg13g2_decap_8 FILLER_26_525 ();
 sg13g2_decap_8 FILLER_26_532 ();
 sg13g2_decap_8 FILLER_26_539 ();
 sg13g2_decap_8 FILLER_26_546 ();
 sg13g2_decap_8 FILLER_26_553 ();
 sg13g2_decap_8 FILLER_26_560 ();
 sg13g2_decap_8 FILLER_26_567 ();
 sg13g2_decap_8 FILLER_26_574 ();
 sg13g2_decap_8 FILLER_26_581 ();
 sg13g2_decap_8 FILLER_26_588 ();
 sg13g2_decap_8 FILLER_26_595 ();
 sg13g2_decap_8 FILLER_26_602 ();
 sg13g2_decap_8 FILLER_26_609 ();
 sg13g2_decap_8 FILLER_26_616 ();
 sg13g2_decap_8 FILLER_26_623 ();
 sg13g2_decap_8 FILLER_26_630 ();
 sg13g2_decap_8 FILLER_26_637 ();
 sg13g2_decap_8 FILLER_26_644 ();
 sg13g2_decap_8 FILLER_26_651 ();
 sg13g2_decap_8 FILLER_26_658 ();
 sg13g2_decap_8 FILLER_26_665 ();
 sg13g2_decap_8 FILLER_26_672 ();
 sg13g2_decap_8 FILLER_26_679 ();
 sg13g2_decap_8 FILLER_26_686 ();
 sg13g2_decap_8 FILLER_26_693 ();
 sg13g2_decap_8 FILLER_26_700 ();
 sg13g2_decap_8 FILLER_26_707 ();
 sg13g2_decap_8 FILLER_26_714 ();
 sg13g2_decap_8 FILLER_26_721 ();
 sg13g2_decap_8 FILLER_26_728 ();
 sg13g2_decap_8 FILLER_26_735 ();
 sg13g2_decap_8 FILLER_26_742 ();
 sg13g2_decap_8 FILLER_26_749 ();
 sg13g2_decap_8 FILLER_26_756 ();
 sg13g2_decap_8 FILLER_26_763 ();
 sg13g2_decap_8 FILLER_26_770 ();
 sg13g2_decap_8 FILLER_26_777 ();
 sg13g2_decap_8 FILLER_26_784 ();
 sg13g2_decap_8 FILLER_26_791 ();
 sg13g2_decap_8 FILLER_26_798 ();
 sg13g2_decap_8 FILLER_26_805 ();
 sg13g2_decap_8 FILLER_26_812 ();
 sg13g2_decap_8 FILLER_26_819 ();
 sg13g2_decap_8 FILLER_26_826 ();
 sg13g2_decap_8 FILLER_26_833 ();
 sg13g2_decap_8 FILLER_26_840 ();
 sg13g2_decap_8 FILLER_26_847 ();
 sg13g2_decap_8 FILLER_26_854 ();
 sg13g2_fill_1 FILLER_26_861 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_decap_8 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_294 ();
 sg13g2_decap_8 FILLER_27_301 ();
 sg13g2_decap_8 FILLER_27_308 ();
 sg13g2_decap_8 FILLER_27_315 ();
 sg13g2_decap_8 FILLER_27_322 ();
 sg13g2_decap_8 FILLER_27_329 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_decap_8 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_decap_8 FILLER_27_406 ();
 sg13g2_decap_8 FILLER_27_413 ();
 sg13g2_decap_8 FILLER_27_420 ();
 sg13g2_decap_8 FILLER_27_427 ();
 sg13g2_decap_8 FILLER_27_434 ();
 sg13g2_decap_8 FILLER_27_441 ();
 sg13g2_decap_8 FILLER_27_448 ();
 sg13g2_decap_8 FILLER_27_455 ();
 sg13g2_decap_8 FILLER_27_462 ();
 sg13g2_decap_8 FILLER_27_469 ();
 sg13g2_decap_8 FILLER_27_476 ();
 sg13g2_decap_8 FILLER_27_483 ();
 sg13g2_decap_8 FILLER_27_490 ();
 sg13g2_decap_8 FILLER_27_497 ();
 sg13g2_decap_8 FILLER_27_504 ();
 sg13g2_decap_8 FILLER_27_511 ();
 sg13g2_decap_8 FILLER_27_518 ();
 sg13g2_decap_8 FILLER_27_525 ();
 sg13g2_decap_8 FILLER_27_532 ();
 sg13g2_decap_8 FILLER_27_539 ();
 sg13g2_decap_8 FILLER_27_546 ();
 sg13g2_decap_8 FILLER_27_553 ();
 sg13g2_decap_8 FILLER_27_560 ();
 sg13g2_decap_8 FILLER_27_567 ();
 sg13g2_decap_8 FILLER_27_574 ();
 sg13g2_decap_8 FILLER_27_581 ();
 sg13g2_decap_8 FILLER_27_588 ();
 sg13g2_decap_8 FILLER_27_595 ();
 sg13g2_decap_8 FILLER_27_602 ();
 sg13g2_decap_8 FILLER_27_609 ();
 sg13g2_decap_8 FILLER_27_616 ();
 sg13g2_decap_8 FILLER_27_623 ();
 sg13g2_decap_8 FILLER_27_630 ();
 sg13g2_decap_8 FILLER_27_637 ();
 sg13g2_decap_8 FILLER_27_644 ();
 sg13g2_decap_8 FILLER_27_651 ();
 sg13g2_decap_8 FILLER_27_658 ();
 sg13g2_decap_8 FILLER_27_665 ();
 sg13g2_decap_8 FILLER_27_672 ();
 sg13g2_decap_8 FILLER_27_679 ();
 sg13g2_decap_8 FILLER_27_686 ();
 sg13g2_decap_8 FILLER_27_693 ();
 sg13g2_decap_8 FILLER_27_700 ();
 sg13g2_decap_8 FILLER_27_707 ();
 sg13g2_decap_8 FILLER_27_714 ();
 sg13g2_decap_8 FILLER_27_721 ();
 sg13g2_decap_8 FILLER_27_728 ();
 sg13g2_decap_8 FILLER_27_735 ();
 sg13g2_decap_8 FILLER_27_742 ();
 sg13g2_decap_8 FILLER_27_749 ();
 sg13g2_decap_8 FILLER_27_756 ();
 sg13g2_decap_8 FILLER_27_763 ();
 sg13g2_decap_8 FILLER_27_770 ();
 sg13g2_decap_8 FILLER_27_777 ();
 sg13g2_decap_8 FILLER_27_784 ();
 sg13g2_decap_8 FILLER_27_791 ();
 sg13g2_decap_8 FILLER_27_798 ();
 sg13g2_decap_8 FILLER_27_805 ();
 sg13g2_decap_8 FILLER_27_812 ();
 sg13g2_decap_8 FILLER_27_819 ();
 sg13g2_decap_8 FILLER_27_826 ();
 sg13g2_decap_8 FILLER_27_833 ();
 sg13g2_decap_8 FILLER_27_840 ();
 sg13g2_decap_8 FILLER_27_847 ();
 sg13g2_decap_8 FILLER_27_854 ();
 sg13g2_fill_1 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_8 FILLER_28_245 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_decap_8 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_266 ();
 sg13g2_decap_8 FILLER_28_273 ();
 sg13g2_decap_8 FILLER_28_280 ();
 sg13g2_decap_8 FILLER_28_287 ();
 sg13g2_decap_8 FILLER_28_294 ();
 sg13g2_decap_8 FILLER_28_301 ();
 sg13g2_decap_8 FILLER_28_308 ();
 sg13g2_decap_8 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_322 ();
 sg13g2_decap_8 FILLER_28_329 ();
 sg13g2_decap_8 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_343 ();
 sg13g2_decap_8 FILLER_28_350 ();
 sg13g2_decap_8 FILLER_28_357 ();
 sg13g2_decap_8 FILLER_28_364 ();
 sg13g2_decap_8 FILLER_28_371 ();
 sg13g2_decap_8 FILLER_28_378 ();
 sg13g2_decap_8 FILLER_28_385 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_decap_8 FILLER_28_406 ();
 sg13g2_decap_8 FILLER_28_413 ();
 sg13g2_decap_8 FILLER_28_420 ();
 sg13g2_decap_8 FILLER_28_427 ();
 sg13g2_decap_8 FILLER_28_434 ();
 sg13g2_decap_8 FILLER_28_441 ();
 sg13g2_decap_8 FILLER_28_448 ();
 sg13g2_decap_8 FILLER_28_455 ();
 sg13g2_decap_8 FILLER_28_462 ();
 sg13g2_decap_8 FILLER_28_469 ();
 sg13g2_decap_8 FILLER_28_476 ();
 sg13g2_decap_8 FILLER_28_483 ();
 sg13g2_decap_8 FILLER_28_490 ();
 sg13g2_decap_8 FILLER_28_497 ();
 sg13g2_decap_8 FILLER_28_504 ();
 sg13g2_decap_8 FILLER_28_511 ();
 sg13g2_decap_8 FILLER_28_518 ();
 sg13g2_decap_8 FILLER_28_525 ();
 sg13g2_decap_8 FILLER_28_532 ();
 sg13g2_decap_8 FILLER_28_539 ();
 sg13g2_decap_8 FILLER_28_546 ();
 sg13g2_decap_8 FILLER_28_553 ();
 sg13g2_decap_8 FILLER_28_560 ();
 sg13g2_decap_8 FILLER_28_567 ();
 sg13g2_decap_8 FILLER_28_574 ();
 sg13g2_decap_8 FILLER_28_581 ();
 sg13g2_decap_8 FILLER_28_588 ();
 sg13g2_decap_8 FILLER_28_595 ();
 sg13g2_decap_8 FILLER_28_602 ();
 sg13g2_decap_8 FILLER_28_609 ();
 sg13g2_decap_8 FILLER_28_616 ();
 sg13g2_decap_8 FILLER_28_623 ();
 sg13g2_decap_8 FILLER_28_630 ();
 sg13g2_decap_8 FILLER_28_637 ();
 sg13g2_decap_8 FILLER_28_644 ();
 sg13g2_decap_8 FILLER_28_651 ();
 sg13g2_decap_8 FILLER_28_658 ();
 sg13g2_decap_8 FILLER_28_665 ();
 sg13g2_decap_8 FILLER_28_672 ();
 sg13g2_decap_8 FILLER_28_679 ();
 sg13g2_decap_8 FILLER_28_686 ();
 sg13g2_decap_8 FILLER_28_693 ();
 sg13g2_decap_8 FILLER_28_700 ();
 sg13g2_decap_8 FILLER_28_707 ();
 sg13g2_decap_8 FILLER_28_714 ();
 sg13g2_decap_8 FILLER_28_721 ();
 sg13g2_decap_8 FILLER_28_728 ();
 sg13g2_decap_8 FILLER_28_735 ();
 sg13g2_decap_8 FILLER_28_742 ();
 sg13g2_decap_8 FILLER_28_749 ();
 sg13g2_decap_8 FILLER_28_756 ();
 sg13g2_decap_8 FILLER_28_763 ();
 sg13g2_decap_8 FILLER_28_770 ();
 sg13g2_decap_8 FILLER_28_777 ();
 sg13g2_decap_8 FILLER_28_784 ();
 sg13g2_decap_8 FILLER_28_791 ();
 sg13g2_decap_8 FILLER_28_798 ();
 sg13g2_decap_8 FILLER_28_805 ();
 sg13g2_decap_8 FILLER_28_812 ();
 sg13g2_decap_8 FILLER_28_819 ();
 sg13g2_decap_8 FILLER_28_826 ();
 sg13g2_decap_8 FILLER_28_833 ();
 sg13g2_decap_8 FILLER_28_840 ();
 sg13g2_decap_8 FILLER_28_847 ();
 sg13g2_decap_8 FILLER_28_854 ();
 sg13g2_fill_1 FILLER_28_861 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_231 ();
 sg13g2_decap_8 FILLER_29_238 ();
 sg13g2_decap_8 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_252 ();
 sg13g2_decap_8 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_decap_8 FILLER_29_280 ();
 sg13g2_decap_8 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_29_294 ();
 sg13g2_decap_8 FILLER_29_301 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_decap_8 FILLER_29_322 ();
 sg13g2_decap_8 FILLER_29_329 ();
 sg13g2_decap_8 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_343 ();
 sg13g2_decap_8 FILLER_29_350 ();
 sg13g2_decap_8 FILLER_29_357 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_decap_8 FILLER_29_406 ();
 sg13g2_decap_8 FILLER_29_413 ();
 sg13g2_decap_8 FILLER_29_420 ();
 sg13g2_decap_8 FILLER_29_427 ();
 sg13g2_decap_8 FILLER_29_434 ();
 sg13g2_decap_8 FILLER_29_441 ();
 sg13g2_decap_8 FILLER_29_448 ();
 sg13g2_decap_8 FILLER_29_455 ();
 sg13g2_decap_8 FILLER_29_462 ();
 sg13g2_decap_8 FILLER_29_469 ();
 sg13g2_decap_8 FILLER_29_476 ();
 sg13g2_decap_8 FILLER_29_483 ();
 sg13g2_decap_8 FILLER_29_490 ();
 sg13g2_decap_8 FILLER_29_497 ();
 sg13g2_decap_8 FILLER_29_504 ();
 sg13g2_decap_8 FILLER_29_511 ();
 sg13g2_decap_8 FILLER_29_518 ();
 sg13g2_decap_8 FILLER_29_525 ();
 sg13g2_decap_8 FILLER_29_532 ();
 sg13g2_decap_8 FILLER_29_539 ();
 sg13g2_decap_8 FILLER_29_546 ();
 sg13g2_decap_8 FILLER_29_553 ();
 sg13g2_decap_8 FILLER_29_560 ();
 sg13g2_decap_8 FILLER_29_567 ();
 sg13g2_decap_8 FILLER_29_574 ();
 sg13g2_decap_8 FILLER_29_581 ();
 sg13g2_decap_8 FILLER_29_588 ();
 sg13g2_decap_8 FILLER_29_595 ();
 sg13g2_decap_8 FILLER_29_602 ();
 sg13g2_decap_8 FILLER_29_609 ();
 sg13g2_decap_8 FILLER_29_616 ();
 sg13g2_decap_8 FILLER_29_623 ();
 sg13g2_decap_8 FILLER_29_630 ();
 sg13g2_decap_8 FILLER_29_637 ();
 sg13g2_decap_8 FILLER_29_644 ();
 sg13g2_decap_8 FILLER_29_651 ();
 sg13g2_decap_8 FILLER_29_658 ();
 sg13g2_decap_8 FILLER_29_665 ();
 sg13g2_decap_8 FILLER_29_672 ();
 sg13g2_decap_8 FILLER_29_679 ();
 sg13g2_decap_8 FILLER_29_686 ();
 sg13g2_decap_8 FILLER_29_693 ();
 sg13g2_decap_8 FILLER_29_700 ();
 sg13g2_decap_8 FILLER_29_707 ();
 sg13g2_decap_8 FILLER_29_714 ();
 sg13g2_decap_8 FILLER_29_721 ();
 sg13g2_decap_8 FILLER_29_728 ();
 sg13g2_decap_8 FILLER_29_735 ();
 sg13g2_decap_8 FILLER_29_742 ();
 sg13g2_decap_8 FILLER_29_749 ();
 sg13g2_decap_8 FILLER_29_756 ();
 sg13g2_decap_8 FILLER_29_763 ();
 sg13g2_decap_8 FILLER_29_770 ();
 sg13g2_decap_8 FILLER_29_777 ();
 sg13g2_decap_8 FILLER_29_784 ();
 sg13g2_decap_8 FILLER_29_791 ();
 sg13g2_decap_8 FILLER_29_798 ();
 sg13g2_decap_8 FILLER_29_805 ();
 sg13g2_decap_8 FILLER_29_812 ();
 sg13g2_decap_8 FILLER_29_819 ();
 sg13g2_decap_8 FILLER_29_826 ();
 sg13g2_decap_8 FILLER_29_833 ();
 sg13g2_decap_8 FILLER_29_840 ();
 sg13g2_decap_8 FILLER_29_847 ();
 sg13g2_decap_8 FILLER_29_854 ();
 sg13g2_fill_1 FILLER_29_861 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_266 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_350 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_decap_8 FILLER_30_406 ();
 sg13g2_decap_8 FILLER_30_413 ();
 sg13g2_decap_8 FILLER_30_420 ();
 sg13g2_decap_8 FILLER_30_427 ();
 sg13g2_decap_8 FILLER_30_434 ();
 sg13g2_decap_8 FILLER_30_441 ();
 sg13g2_decap_8 FILLER_30_448 ();
 sg13g2_decap_8 FILLER_30_455 ();
 sg13g2_decap_8 FILLER_30_462 ();
 sg13g2_decap_8 FILLER_30_469 ();
 sg13g2_decap_8 FILLER_30_476 ();
 sg13g2_decap_8 FILLER_30_483 ();
 sg13g2_decap_8 FILLER_30_490 ();
 sg13g2_decap_8 FILLER_30_497 ();
 sg13g2_decap_8 FILLER_30_504 ();
 sg13g2_decap_8 FILLER_30_511 ();
 sg13g2_decap_8 FILLER_30_518 ();
 sg13g2_decap_8 FILLER_30_525 ();
 sg13g2_decap_8 FILLER_30_532 ();
 sg13g2_decap_8 FILLER_30_539 ();
 sg13g2_decap_8 FILLER_30_546 ();
 sg13g2_decap_8 FILLER_30_553 ();
 sg13g2_decap_8 FILLER_30_560 ();
 sg13g2_decap_8 FILLER_30_567 ();
 sg13g2_decap_8 FILLER_30_574 ();
 sg13g2_decap_8 FILLER_30_581 ();
 sg13g2_decap_8 FILLER_30_588 ();
 sg13g2_decap_8 FILLER_30_595 ();
 sg13g2_decap_8 FILLER_30_602 ();
 sg13g2_decap_8 FILLER_30_609 ();
 sg13g2_decap_8 FILLER_30_616 ();
 sg13g2_decap_8 FILLER_30_623 ();
 sg13g2_decap_8 FILLER_30_630 ();
 sg13g2_decap_8 FILLER_30_637 ();
 sg13g2_decap_8 FILLER_30_644 ();
 sg13g2_decap_8 FILLER_30_651 ();
 sg13g2_decap_8 FILLER_30_658 ();
 sg13g2_decap_8 FILLER_30_665 ();
 sg13g2_decap_8 FILLER_30_672 ();
 sg13g2_decap_8 FILLER_30_679 ();
 sg13g2_decap_8 FILLER_30_686 ();
 sg13g2_decap_8 FILLER_30_693 ();
 sg13g2_decap_8 FILLER_30_700 ();
 sg13g2_decap_8 FILLER_30_707 ();
 sg13g2_decap_8 FILLER_30_714 ();
 sg13g2_decap_8 FILLER_30_721 ();
 sg13g2_decap_8 FILLER_30_728 ();
 sg13g2_decap_8 FILLER_30_735 ();
 sg13g2_decap_8 FILLER_30_742 ();
 sg13g2_decap_8 FILLER_30_749 ();
 sg13g2_decap_8 FILLER_30_756 ();
 sg13g2_decap_8 FILLER_30_763 ();
 sg13g2_decap_8 FILLER_30_770 ();
 sg13g2_decap_8 FILLER_30_777 ();
 sg13g2_decap_8 FILLER_30_784 ();
 sg13g2_decap_8 FILLER_30_791 ();
 sg13g2_decap_8 FILLER_30_798 ();
 sg13g2_decap_8 FILLER_30_805 ();
 sg13g2_decap_8 FILLER_30_812 ();
 sg13g2_decap_8 FILLER_30_819 ();
 sg13g2_decap_8 FILLER_30_826 ();
 sg13g2_decap_8 FILLER_30_833 ();
 sg13g2_decap_8 FILLER_30_840 ();
 sg13g2_decap_8 FILLER_30_847 ();
 sg13g2_decap_8 FILLER_30_854 ();
 sg13g2_fill_1 FILLER_30_861 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_252 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_266 ();
 sg13g2_decap_8 FILLER_31_273 ();
 sg13g2_decap_8 FILLER_31_280 ();
 sg13g2_decap_8 FILLER_31_287 ();
 sg13g2_decap_8 FILLER_31_294 ();
 sg13g2_decap_8 FILLER_31_301 ();
 sg13g2_decap_8 FILLER_31_308 ();
 sg13g2_decap_8 FILLER_31_315 ();
 sg13g2_decap_8 FILLER_31_322 ();
 sg13g2_decap_8 FILLER_31_329 ();
 sg13g2_decap_8 FILLER_31_336 ();
 sg13g2_decap_8 FILLER_31_343 ();
 sg13g2_decap_8 FILLER_31_350 ();
 sg13g2_decap_8 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_371 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_decap_8 FILLER_31_406 ();
 sg13g2_decap_8 FILLER_31_413 ();
 sg13g2_decap_8 FILLER_31_420 ();
 sg13g2_decap_8 FILLER_31_427 ();
 sg13g2_decap_8 FILLER_31_434 ();
 sg13g2_decap_8 FILLER_31_441 ();
 sg13g2_decap_8 FILLER_31_448 ();
 sg13g2_decap_8 FILLER_31_455 ();
 sg13g2_decap_8 FILLER_31_462 ();
 sg13g2_decap_8 FILLER_31_469 ();
 sg13g2_decap_8 FILLER_31_476 ();
 sg13g2_decap_8 FILLER_31_483 ();
 sg13g2_decap_8 FILLER_31_490 ();
 sg13g2_decap_8 FILLER_31_497 ();
 sg13g2_decap_8 FILLER_31_504 ();
 sg13g2_decap_8 FILLER_31_511 ();
 sg13g2_decap_8 FILLER_31_518 ();
 sg13g2_decap_8 FILLER_31_525 ();
 sg13g2_decap_8 FILLER_31_532 ();
 sg13g2_decap_8 FILLER_31_539 ();
 sg13g2_decap_8 FILLER_31_546 ();
 sg13g2_decap_8 FILLER_31_553 ();
 sg13g2_decap_8 FILLER_31_560 ();
 sg13g2_decap_8 FILLER_31_567 ();
 sg13g2_decap_8 FILLER_31_574 ();
 sg13g2_decap_8 FILLER_31_581 ();
 sg13g2_decap_8 FILLER_31_588 ();
 sg13g2_decap_8 FILLER_31_595 ();
 sg13g2_decap_8 FILLER_31_602 ();
 sg13g2_decap_8 FILLER_31_609 ();
 sg13g2_decap_8 FILLER_31_616 ();
 sg13g2_decap_8 FILLER_31_623 ();
 sg13g2_decap_8 FILLER_31_630 ();
 sg13g2_decap_8 FILLER_31_637 ();
 sg13g2_decap_8 FILLER_31_644 ();
 sg13g2_decap_8 FILLER_31_651 ();
 sg13g2_decap_8 FILLER_31_658 ();
 sg13g2_decap_8 FILLER_31_665 ();
 sg13g2_decap_8 FILLER_31_672 ();
 sg13g2_decap_8 FILLER_31_679 ();
 sg13g2_decap_8 FILLER_31_686 ();
 sg13g2_decap_8 FILLER_31_693 ();
 sg13g2_decap_8 FILLER_31_700 ();
 sg13g2_decap_8 FILLER_31_707 ();
 sg13g2_decap_8 FILLER_31_714 ();
 sg13g2_decap_8 FILLER_31_721 ();
 sg13g2_decap_8 FILLER_31_728 ();
 sg13g2_decap_8 FILLER_31_735 ();
 sg13g2_decap_8 FILLER_31_742 ();
 sg13g2_decap_8 FILLER_31_749 ();
 sg13g2_decap_8 FILLER_31_756 ();
 sg13g2_decap_8 FILLER_31_763 ();
 sg13g2_decap_8 FILLER_31_770 ();
 sg13g2_decap_8 FILLER_31_777 ();
 sg13g2_decap_8 FILLER_31_784 ();
 sg13g2_decap_8 FILLER_31_791 ();
 sg13g2_decap_8 FILLER_31_798 ();
 sg13g2_decap_8 FILLER_31_805 ();
 sg13g2_decap_8 FILLER_31_812 ();
 sg13g2_decap_8 FILLER_31_819 ();
 sg13g2_decap_8 FILLER_31_826 ();
 sg13g2_decap_8 FILLER_31_833 ();
 sg13g2_decap_8 FILLER_31_840 ();
 sg13g2_decap_8 FILLER_31_847 ();
 sg13g2_decap_8 FILLER_31_854 ();
 sg13g2_fill_1 FILLER_31_861 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_245 ();
 sg13g2_decap_8 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_259 ();
 sg13g2_decap_8 FILLER_32_266 ();
 sg13g2_decap_8 FILLER_32_273 ();
 sg13g2_decap_8 FILLER_32_280 ();
 sg13g2_decap_8 FILLER_32_287 ();
 sg13g2_decap_8 FILLER_32_294 ();
 sg13g2_decap_8 FILLER_32_301 ();
 sg13g2_decap_8 FILLER_32_308 ();
 sg13g2_decap_8 FILLER_32_315 ();
 sg13g2_decap_8 FILLER_32_322 ();
 sg13g2_decap_8 FILLER_32_329 ();
 sg13g2_decap_8 FILLER_32_336 ();
 sg13g2_decap_8 FILLER_32_343 ();
 sg13g2_decap_8 FILLER_32_350 ();
 sg13g2_decap_8 FILLER_32_357 ();
 sg13g2_decap_8 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_decap_8 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_decap_8 FILLER_32_406 ();
 sg13g2_decap_8 FILLER_32_413 ();
 sg13g2_decap_8 FILLER_32_420 ();
 sg13g2_decap_8 FILLER_32_427 ();
 sg13g2_decap_8 FILLER_32_434 ();
 sg13g2_decap_8 FILLER_32_441 ();
 sg13g2_decap_8 FILLER_32_448 ();
 sg13g2_decap_8 FILLER_32_455 ();
 sg13g2_decap_8 FILLER_32_462 ();
 sg13g2_decap_8 FILLER_32_469 ();
 sg13g2_decap_8 FILLER_32_476 ();
 sg13g2_decap_8 FILLER_32_483 ();
 sg13g2_decap_8 FILLER_32_490 ();
 sg13g2_decap_8 FILLER_32_497 ();
 sg13g2_decap_8 FILLER_32_504 ();
 sg13g2_decap_8 FILLER_32_511 ();
 sg13g2_decap_8 FILLER_32_518 ();
 sg13g2_decap_8 FILLER_32_525 ();
 sg13g2_decap_8 FILLER_32_532 ();
 sg13g2_decap_8 FILLER_32_539 ();
 sg13g2_decap_8 FILLER_32_546 ();
 sg13g2_decap_8 FILLER_32_553 ();
 sg13g2_decap_8 FILLER_32_560 ();
 sg13g2_decap_8 FILLER_32_567 ();
 sg13g2_decap_8 FILLER_32_574 ();
 sg13g2_decap_8 FILLER_32_581 ();
 sg13g2_decap_8 FILLER_32_588 ();
 sg13g2_decap_8 FILLER_32_595 ();
 sg13g2_decap_8 FILLER_32_602 ();
 sg13g2_decap_8 FILLER_32_609 ();
 sg13g2_decap_8 FILLER_32_616 ();
 sg13g2_decap_8 FILLER_32_623 ();
 sg13g2_decap_8 FILLER_32_630 ();
 sg13g2_decap_8 FILLER_32_637 ();
 sg13g2_decap_8 FILLER_32_644 ();
 sg13g2_decap_8 FILLER_32_651 ();
 sg13g2_decap_8 FILLER_32_658 ();
 sg13g2_decap_8 FILLER_32_665 ();
 sg13g2_decap_8 FILLER_32_672 ();
 sg13g2_decap_8 FILLER_32_679 ();
 sg13g2_decap_8 FILLER_32_686 ();
 sg13g2_decap_8 FILLER_32_693 ();
 sg13g2_decap_8 FILLER_32_700 ();
 sg13g2_decap_8 FILLER_32_707 ();
 sg13g2_decap_8 FILLER_32_714 ();
 sg13g2_decap_8 FILLER_32_721 ();
 sg13g2_decap_8 FILLER_32_728 ();
 sg13g2_decap_8 FILLER_32_735 ();
 sg13g2_decap_8 FILLER_32_742 ();
 sg13g2_decap_8 FILLER_32_749 ();
 sg13g2_decap_8 FILLER_32_756 ();
 sg13g2_decap_8 FILLER_32_763 ();
 sg13g2_decap_8 FILLER_32_770 ();
 sg13g2_decap_8 FILLER_32_777 ();
 sg13g2_decap_8 FILLER_32_784 ();
 sg13g2_decap_8 FILLER_32_791 ();
 sg13g2_decap_8 FILLER_32_798 ();
 sg13g2_decap_8 FILLER_32_805 ();
 sg13g2_decap_8 FILLER_32_812 ();
 sg13g2_decap_8 FILLER_32_819 ();
 sg13g2_decap_8 FILLER_32_826 ();
 sg13g2_decap_8 FILLER_32_833 ();
 sg13g2_decap_8 FILLER_32_840 ();
 sg13g2_decap_8 FILLER_32_847 ();
 sg13g2_decap_8 FILLER_32_854 ();
 sg13g2_fill_1 FILLER_32_861 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_273 ();
 sg13g2_decap_8 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_287 ();
 sg13g2_decap_8 FILLER_33_294 ();
 sg13g2_decap_8 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_308 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_decap_8 FILLER_33_322 ();
 sg13g2_decap_8 FILLER_33_329 ();
 sg13g2_decap_8 FILLER_33_336 ();
 sg13g2_decap_8 FILLER_33_343 ();
 sg13g2_decap_8 FILLER_33_350 ();
 sg13g2_decap_8 FILLER_33_357 ();
 sg13g2_decap_8 FILLER_33_364 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_decap_8 FILLER_33_406 ();
 sg13g2_decap_8 FILLER_33_413 ();
 sg13g2_decap_8 FILLER_33_420 ();
 sg13g2_decap_8 FILLER_33_427 ();
 sg13g2_decap_8 FILLER_33_434 ();
 sg13g2_decap_8 FILLER_33_441 ();
 sg13g2_decap_8 FILLER_33_448 ();
 sg13g2_decap_8 FILLER_33_455 ();
 sg13g2_decap_8 FILLER_33_462 ();
 sg13g2_decap_8 FILLER_33_469 ();
 sg13g2_decap_8 FILLER_33_476 ();
 sg13g2_decap_8 FILLER_33_483 ();
 sg13g2_decap_8 FILLER_33_490 ();
 sg13g2_decap_8 FILLER_33_497 ();
 sg13g2_decap_8 FILLER_33_504 ();
 sg13g2_decap_8 FILLER_33_511 ();
 sg13g2_decap_8 FILLER_33_518 ();
 sg13g2_decap_8 FILLER_33_525 ();
 sg13g2_decap_8 FILLER_33_532 ();
 sg13g2_decap_8 FILLER_33_539 ();
 sg13g2_decap_8 FILLER_33_546 ();
 sg13g2_decap_8 FILLER_33_553 ();
 sg13g2_decap_8 FILLER_33_560 ();
 sg13g2_decap_8 FILLER_33_567 ();
 sg13g2_decap_8 FILLER_33_574 ();
 sg13g2_decap_8 FILLER_33_581 ();
 sg13g2_decap_8 FILLER_33_588 ();
 sg13g2_decap_8 FILLER_33_595 ();
 sg13g2_decap_8 FILLER_33_602 ();
 sg13g2_decap_8 FILLER_33_609 ();
 sg13g2_decap_8 FILLER_33_616 ();
 sg13g2_decap_8 FILLER_33_623 ();
 sg13g2_decap_8 FILLER_33_630 ();
 sg13g2_decap_8 FILLER_33_637 ();
 sg13g2_decap_8 FILLER_33_644 ();
 sg13g2_decap_8 FILLER_33_651 ();
 sg13g2_decap_8 FILLER_33_658 ();
 sg13g2_decap_8 FILLER_33_665 ();
 sg13g2_decap_8 FILLER_33_672 ();
 sg13g2_decap_8 FILLER_33_679 ();
 sg13g2_decap_8 FILLER_33_686 ();
 sg13g2_decap_8 FILLER_33_693 ();
 sg13g2_decap_8 FILLER_33_700 ();
 sg13g2_decap_8 FILLER_33_707 ();
 sg13g2_decap_8 FILLER_33_714 ();
 sg13g2_decap_8 FILLER_33_721 ();
 sg13g2_decap_8 FILLER_33_728 ();
 sg13g2_decap_8 FILLER_33_735 ();
 sg13g2_decap_8 FILLER_33_742 ();
 sg13g2_decap_8 FILLER_33_749 ();
 sg13g2_decap_8 FILLER_33_756 ();
 sg13g2_decap_8 FILLER_33_763 ();
 sg13g2_decap_8 FILLER_33_770 ();
 sg13g2_decap_8 FILLER_33_777 ();
 sg13g2_decap_8 FILLER_33_784 ();
 sg13g2_decap_8 FILLER_33_791 ();
 sg13g2_decap_8 FILLER_33_798 ();
 sg13g2_decap_8 FILLER_33_805 ();
 sg13g2_decap_8 FILLER_33_812 ();
 sg13g2_decap_8 FILLER_33_819 ();
 sg13g2_decap_8 FILLER_33_826 ();
 sg13g2_decap_8 FILLER_33_833 ();
 sg13g2_decap_8 FILLER_33_840 ();
 sg13g2_decap_8 FILLER_33_847 ();
 sg13g2_decap_8 FILLER_33_854 ();
 sg13g2_fill_1 FILLER_33_861 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_280 ();
 sg13g2_decap_8 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_294 ();
 sg13g2_decap_8 FILLER_34_301 ();
 sg13g2_decap_8 FILLER_34_308 ();
 sg13g2_decap_8 FILLER_34_315 ();
 sg13g2_decap_8 FILLER_34_322 ();
 sg13g2_decap_8 FILLER_34_329 ();
 sg13g2_decap_8 FILLER_34_336 ();
 sg13g2_decap_8 FILLER_34_343 ();
 sg13g2_decap_8 FILLER_34_350 ();
 sg13g2_decap_8 FILLER_34_357 ();
 sg13g2_decap_8 FILLER_34_364 ();
 sg13g2_decap_8 FILLER_34_371 ();
 sg13g2_decap_8 FILLER_34_378 ();
 sg13g2_decap_8 FILLER_34_385 ();
 sg13g2_decap_8 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_decap_8 FILLER_34_406 ();
 sg13g2_decap_8 FILLER_34_413 ();
 sg13g2_decap_8 FILLER_34_420 ();
 sg13g2_decap_8 FILLER_34_427 ();
 sg13g2_decap_8 FILLER_34_434 ();
 sg13g2_decap_8 FILLER_34_441 ();
 sg13g2_decap_8 FILLER_34_448 ();
 sg13g2_decap_8 FILLER_34_455 ();
 sg13g2_decap_8 FILLER_34_462 ();
 sg13g2_decap_8 FILLER_34_469 ();
 sg13g2_decap_8 FILLER_34_476 ();
 sg13g2_decap_8 FILLER_34_483 ();
 sg13g2_decap_8 FILLER_34_490 ();
 sg13g2_decap_8 FILLER_34_497 ();
 sg13g2_decap_8 FILLER_34_504 ();
 sg13g2_decap_8 FILLER_34_511 ();
 sg13g2_decap_8 FILLER_34_518 ();
 sg13g2_decap_8 FILLER_34_525 ();
 sg13g2_decap_8 FILLER_34_532 ();
 sg13g2_decap_8 FILLER_34_539 ();
 sg13g2_decap_8 FILLER_34_546 ();
 sg13g2_decap_8 FILLER_34_553 ();
 sg13g2_decap_8 FILLER_34_560 ();
 sg13g2_decap_8 FILLER_34_567 ();
 sg13g2_decap_8 FILLER_34_574 ();
 sg13g2_decap_8 FILLER_34_581 ();
 sg13g2_decap_8 FILLER_34_588 ();
 sg13g2_decap_8 FILLER_34_595 ();
 sg13g2_decap_8 FILLER_34_602 ();
 sg13g2_decap_8 FILLER_34_609 ();
 sg13g2_decap_8 FILLER_34_616 ();
 sg13g2_decap_8 FILLER_34_623 ();
 sg13g2_decap_8 FILLER_34_630 ();
 sg13g2_decap_8 FILLER_34_637 ();
 sg13g2_decap_8 FILLER_34_644 ();
 sg13g2_decap_8 FILLER_34_651 ();
 sg13g2_decap_8 FILLER_34_658 ();
 sg13g2_decap_8 FILLER_34_665 ();
 sg13g2_decap_8 FILLER_34_672 ();
 sg13g2_decap_8 FILLER_34_679 ();
 sg13g2_decap_8 FILLER_34_686 ();
 sg13g2_decap_8 FILLER_34_693 ();
 sg13g2_decap_8 FILLER_34_700 ();
 sg13g2_decap_8 FILLER_34_707 ();
 sg13g2_decap_8 FILLER_34_714 ();
 sg13g2_decap_8 FILLER_34_721 ();
 sg13g2_decap_8 FILLER_34_728 ();
 sg13g2_decap_8 FILLER_34_735 ();
 sg13g2_decap_8 FILLER_34_742 ();
 sg13g2_decap_8 FILLER_34_749 ();
 sg13g2_decap_8 FILLER_34_756 ();
 sg13g2_decap_8 FILLER_34_763 ();
 sg13g2_decap_8 FILLER_34_770 ();
 sg13g2_decap_8 FILLER_34_777 ();
 sg13g2_decap_8 FILLER_34_784 ();
 sg13g2_decap_8 FILLER_34_791 ();
 sg13g2_decap_8 FILLER_34_798 ();
 sg13g2_decap_8 FILLER_34_805 ();
 sg13g2_decap_8 FILLER_34_812 ();
 sg13g2_decap_8 FILLER_34_819 ();
 sg13g2_decap_8 FILLER_34_826 ();
 sg13g2_decap_8 FILLER_34_833 ();
 sg13g2_decap_8 FILLER_34_840 ();
 sg13g2_decap_8 FILLER_34_847 ();
 sg13g2_decap_8 FILLER_34_854 ();
 sg13g2_fill_1 FILLER_34_861 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_245 ();
 sg13g2_decap_8 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_266 ();
 sg13g2_decap_8 FILLER_35_273 ();
 sg13g2_decap_8 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_decap_8 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_decap_8 FILLER_35_322 ();
 sg13g2_decap_8 FILLER_35_329 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_decap_8 FILLER_35_406 ();
 sg13g2_decap_8 FILLER_35_413 ();
 sg13g2_decap_8 FILLER_35_420 ();
 sg13g2_decap_8 FILLER_35_427 ();
 sg13g2_decap_8 FILLER_35_434 ();
 sg13g2_decap_8 FILLER_35_441 ();
 sg13g2_decap_8 FILLER_35_448 ();
 sg13g2_decap_8 FILLER_35_455 ();
 sg13g2_decap_8 FILLER_35_462 ();
 sg13g2_decap_8 FILLER_35_469 ();
 sg13g2_decap_8 FILLER_35_476 ();
 sg13g2_decap_8 FILLER_35_483 ();
 sg13g2_decap_8 FILLER_35_490 ();
 sg13g2_decap_8 FILLER_35_497 ();
 sg13g2_decap_8 FILLER_35_504 ();
 sg13g2_decap_8 FILLER_35_511 ();
 sg13g2_decap_8 FILLER_35_518 ();
 sg13g2_decap_8 FILLER_35_525 ();
 sg13g2_decap_8 FILLER_35_532 ();
 sg13g2_decap_8 FILLER_35_539 ();
 sg13g2_decap_8 FILLER_35_546 ();
 sg13g2_decap_8 FILLER_35_553 ();
 sg13g2_decap_8 FILLER_35_560 ();
 sg13g2_decap_8 FILLER_35_567 ();
 sg13g2_decap_8 FILLER_35_574 ();
 sg13g2_decap_8 FILLER_35_581 ();
 sg13g2_decap_8 FILLER_35_588 ();
 sg13g2_decap_8 FILLER_35_595 ();
 sg13g2_decap_8 FILLER_35_602 ();
 sg13g2_decap_8 FILLER_35_609 ();
 sg13g2_decap_8 FILLER_35_616 ();
 sg13g2_decap_8 FILLER_35_623 ();
 sg13g2_decap_8 FILLER_35_630 ();
 sg13g2_decap_8 FILLER_35_637 ();
 sg13g2_decap_8 FILLER_35_644 ();
 sg13g2_decap_8 FILLER_35_651 ();
 sg13g2_decap_8 FILLER_35_658 ();
 sg13g2_decap_8 FILLER_35_665 ();
 sg13g2_decap_8 FILLER_35_672 ();
 sg13g2_decap_8 FILLER_35_679 ();
 sg13g2_decap_8 FILLER_35_686 ();
 sg13g2_decap_8 FILLER_35_693 ();
 sg13g2_decap_8 FILLER_35_700 ();
 sg13g2_decap_8 FILLER_35_707 ();
 sg13g2_decap_8 FILLER_35_714 ();
 sg13g2_decap_8 FILLER_35_721 ();
 sg13g2_decap_8 FILLER_35_728 ();
 sg13g2_decap_8 FILLER_35_735 ();
 sg13g2_decap_8 FILLER_35_742 ();
 sg13g2_decap_8 FILLER_35_749 ();
 sg13g2_decap_8 FILLER_35_756 ();
 sg13g2_decap_8 FILLER_35_763 ();
 sg13g2_decap_8 FILLER_35_770 ();
 sg13g2_decap_8 FILLER_35_777 ();
 sg13g2_decap_8 FILLER_35_784 ();
 sg13g2_decap_8 FILLER_35_791 ();
 sg13g2_decap_8 FILLER_35_798 ();
 sg13g2_decap_8 FILLER_35_805 ();
 sg13g2_decap_8 FILLER_35_812 ();
 sg13g2_decap_8 FILLER_35_819 ();
 sg13g2_decap_8 FILLER_35_826 ();
 sg13g2_decap_8 FILLER_35_833 ();
 sg13g2_decap_8 FILLER_35_840 ();
 sg13g2_decap_8 FILLER_35_847 ();
 sg13g2_decap_8 FILLER_35_854 ();
 sg13g2_fill_1 FILLER_35_861 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_4 FILLER_36_126 ();
 sg13g2_fill_2 FILLER_36_130 ();
 sg13g2_decap_4 FILLER_36_136 ();
 sg13g2_decap_4 FILLER_36_144 ();
 sg13g2_fill_2 FILLER_36_153 ();
 sg13g2_decap_8 FILLER_36_159 ();
 sg13g2_decap_4 FILLER_36_166 ();
 sg13g2_fill_2 FILLER_36_170 ();
 sg13g2_decap_8 FILLER_36_177 ();
 sg13g2_decap_8 FILLER_36_184 ();
 sg13g2_decap_8 FILLER_36_191 ();
 sg13g2_decap_8 FILLER_36_198 ();
 sg13g2_decap_8 FILLER_36_205 ();
 sg13g2_decap_8 FILLER_36_212 ();
 sg13g2_decap_8 FILLER_36_219 ();
 sg13g2_decap_8 FILLER_36_226 ();
 sg13g2_decap_8 FILLER_36_233 ();
 sg13g2_decap_8 FILLER_36_240 ();
 sg13g2_decap_8 FILLER_36_247 ();
 sg13g2_decap_8 FILLER_36_254 ();
 sg13g2_decap_8 FILLER_36_261 ();
 sg13g2_decap_8 FILLER_36_268 ();
 sg13g2_decap_8 FILLER_36_275 ();
 sg13g2_decap_8 FILLER_36_282 ();
 sg13g2_decap_8 FILLER_36_289 ();
 sg13g2_decap_8 FILLER_36_296 ();
 sg13g2_decap_8 FILLER_36_303 ();
 sg13g2_decap_8 FILLER_36_310 ();
 sg13g2_decap_8 FILLER_36_317 ();
 sg13g2_decap_8 FILLER_36_324 ();
 sg13g2_decap_8 FILLER_36_331 ();
 sg13g2_decap_8 FILLER_36_338 ();
 sg13g2_decap_8 FILLER_36_345 ();
 sg13g2_decap_8 FILLER_36_352 ();
 sg13g2_decap_8 FILLER_36_359 ();
 sg13g2_decap_8 FILLER_36_366 ();
 sg13g2_decap_8 FILLER_36_373 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_decap_8 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_36_415 ();
 sg13g2_decap_8 FILLER_36_422 ();
 sg13g2_decap_8 FILLER_36_429 ();
 sg13g2_decap_8 FILLER_36_436 ();
 sg13g2_decap_8 FILLER_36_443 ();
 sg13g2_decap_8 FILLER_36_450 ();
 sg13g2_decap_8 FILLER_36_457 ();
 sg13g2_decap_8 FILLER_36_464 ();
 sg13g2_decap_8 FILLER_36_471 ();
 sg13g2_decap_8 FILLER_36_478 ();
 sg13g2_decap_8 FILLER_36_485 ();
 sg13g2_decap_8 FILLER_36_492 ();
 sg13g2_decap_8 FILLER_36_499 ();
 sg13g2_decap_8 FILLER_36_506 ();
 sg13g2_decap_8 FILLER_36_513 ();
 sg13g2_decap_8 FILLER_36_520 ();
 sg13g2_decap_8 FILLER_36_527 ();
 sg13g2_decap_8 FILLER_36_534 ();
 sg13g2_decap_8 FILLER_36_541 ();
 sg13g2_decap_8 FILLER_36_548 ();
 sg13g2_decap_8 FILLER_36_555 ();
 sg13g2_decap_8 FILLER_36_562 ();
 sg13g2_decap_8 FILLER_36_569 ();
 sg13g2_decap_8 FILLER_36_576 ();
 sg13g2_decap_8 FILLER_36_583 ();
 sg13g2_decap_8 FILLER_36_590 ();
 sg13g2_decap_8 FILLER_36_597 ();
 sg13g2_decap_8 FILLER_36_604 ();
 sg13g2_decap_8 FILLER_36_611 ();
 sg13g2_decap_8 FILLER_36_618 ();
 sg13g2_decap_8 FILLER_36_625 ();
 sg13g2_decap_8 FILLER_36_632 ();
 sg13g2_decap_8 FILLER_36_639 ();
 sg13g2_decap_8 FILLER_36_646 ();
 sg13g2_decap_8 FILLER_36_653 ();
 sg13g2_decap_8 FILLER_36_660 ();
 sg13g2_decap_8 FILLER_36_667 ();
 sg13g2_decap_8 FILLER_36_674 ();
 sg13g2_decap_8 FILLER_36_681 ();
 sg13g2_decap_8 FILLER_36_688 ();
 sg13g2_decap_8 FILLER_36_695 ();
 sg13g2_decap_8 FILLER_36_702 ();
 sg13g2_decap_8 FILLER_36_709 ();
 sg13g2_decap_8 FILLER_36_716 ();
 sg13g2_decap_8 FILLER_36_723 ();
 sg13g2_decap_8 FILLER_36_730 ();
 sg13g2_decap_8 FILLER_36_737 ();
 sg13g2_decap_8 FILLER_36_744 ();
 sg13g2_decap_8 FILLER_36_751 ();
 sg13g2_decap_8 FILLER_36_758 ();
 sg13g2_decap_8 FILLER_36_765 ();
 sg13g2_decap_8 FILLER_36_772 ();
 sg13g2_decap_8 FILLER_36_779 ();
 sg13g2_decap_8 FILLER_36_786 ();
 sg13g2_decap_8 FILLER_36_793 ();
 sg13g2_decap_8 FILLER_36_800 ();
 sg13g2_decap_8 FILLER_36_807 ();
 sg13g2_decap_8 FILLER_36_814 ();
 sg13g2_decap_8 FILLER_36_821 ();
 sg13g2_decap_8 FILLER_36_828 ();
 sg13g2_decap_8 FILLER_36_835 ();
 sg13g2_decap_8 FILLER_36_842 ();
 sg13g2_decap_8 FILLER_36_849 ();
 sg13g2_decap_4 FILLER_36_856 ();
 sg13g2_fill_2 FILLER_36_860 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_4 FILLER_37_84 ();
 sg13g2_fill_1 FILLER_37_88 ();
 sg13g2_decap_8 FILLER_37_97 ();
 sg13g2_decap_8 FILLER_37_104 ();
 sg13g2_decap_8 FILLER_37_111 ();
 sg13g2_fill_2 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_193 ();
 sg13g2_decap_8 FILLER_37_204 ();
 sg13g2_decap_8 FILLER_37_211 ();
 sg13g2_decap_8 FILLER_37_218 ();
 sg13g2_decap_8 FILLER_37_225 ();
 sg13g2_decap_8 FILLER_37_232 ();
 sg13g2_decap_8 FILLER_37_239 ();
 sg13g2_decap_8 FILLER_37_246 ();
 sg13g2_decap_4 FILLER_37_253 ();
 sg13g2_fill_2 FILLER_37_257 ();
 sg13g2_decap_8 FILLER_37_263 ();
 sg13g2_fill_2 FILLER_37_270 ();
 sg13g2_fill_1 FILLER_37_272 ();
 sg13g2_decap_8 FILLER_37_304 ();
 sg13g2_fill_2 FILLER_37_311 ();
 sg13g2_decap_8 FILLER_37_317 ();
 sg13g2_decap_8 FILLER_37_324 ();
 sg13g2_decap_8 FILLER_37_331 ();
 sg13g2_decap_8 FILLER_37_338 ();
 sg13g2_decap_8 FILLER_37_345 ();
 sg13g2_decap_8 FILLER_37_352 ();
 sg13g2_decap_8 FILLER_37_359 ();
 sg13g2_decap_8 FILLER_37_366 ();
 sg13g2_decap_8 FILLER_37_373 ();
 sg13g2_decap_8 FILLER_37_380 ();
 sg13g2_decap_8 FILLER_37_387 ();
 sg13g2_decap_8 FILLER_37_394 ();
 sg13g2_decap_8 FILLER_37_401 ();
 sg13g2_decap_8 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_37_415 ();
 sg13g2_decap_8 FILLER_37_422 ();
 sg13g2_decap_8 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_37_436 ();
 sg13g2_decap_8 FILLER_37_443 ();
 sg13g2_decap_8 FILLER_37_450 ();
 sg13g2_decap_8 FILLER_37_457 ();
 sg13g2_decap_8 FILLER_37_464 ();
 sg13g2_decap_8 FILLER_37_471 ();
 sg13g2_decap_8 FILLER_37_478 ();
 sg13g2_decap_8 FILLER_37_485 ();
 sg13g2_decap_8 FILLER_37_492 ();
 sg13g2_decap_8 FILLER_37_499 ();
 sg13g2_decap_8 FILLER_37_506 ();
 sg13g2_decap_8 FILLER_37_513 ();
 sg13g2_decap_8 FILLER_37_520 ();
 sg13g2_decap_8 FILLER_37_527 ();
 sg13g2_decap_8 FILLER_37_534 ();
 sg13g2_decap_8 FILLER_37_541 ();
 sg13g2_decap_8 FILLER_37_548 ();
 sg13g2_decap_8 FILLER_37_555 ();
 sg13g2_decap_8 FILLER_37_562 ();
 sg13g2_decap_8 FILLER_37_569 ();
 sg13g2_decap_8 FILLER_37_576 ();
 sg13g2_decap_8 FILLER_37_583 ();
 sg13g2_decap_8 FILLER_37_590 ();
 sg13g2_decap_8 FILLER_37_597 ();
 sg13g2_decap_8 FILLER_37_604 ();
 sg13g2_decap_8 FILLER_37_611 ();
 sg13g2_decap_8 FILLER_37_618 ();
 sg13g2_decap_8 FILLER_37_625 ();
 sg13g2_decap_8 FILLER_37_632 ();
 sg13g2_decap_8 FILLER_37_639 ();
 sg13g2_decap_8 FILLER_37_646 ();
 sg13g2_decap_8 FILLER_37_653 ();
 sg13g2_decap_8 FILLER_37_660 ();
 sg13g2_decap_8 FILLER_37_667 ();
 sg13g2_decap_8 FILLER_37_674 ();
 sg13g2_decap_8 FILLER_37_681 ();
 sg13g2_decap_8 FILLER_37_688 ();
 sg13g2_decap_8 FILLER_37_695 ();
 sg13g2_decap_8 FILLER_37_702 ();
 sg13g2_decap_8 FILLER_37_709 ();
 sg13g2_decap_8 FILLER_37_716 ();
 sg13g2_decap_8 FILLER_37_723 ();
 sg13g2_decap_8 FILLER_37_730 ();
 sg13g2_decap_8 FILLER_37_737 ();
 sg13g2_decap_8 FILLER_37_744 ();
 sg13g2_decap_8 FILLER_37_751 ();
 sg13g2_decap_8 FILLER_37_758 ();
 sg13g2_decap_8 FILLER_37_765 ();
 sg13g2_decap_8 FILLER_37_772 ();
 sg13g2_decap_8 FILLER_37_779 ();
 sg13g2_decap_8 FILLER_37_786 ();
 sg13g2_decap_8 FILLER_37_793 ();
 sg13g2_decap_8 FILLER_37_800 ();
 sg13g2_decap_8 FILLER_37_807 ();
 sg13g2_decap_8 FILLER_37_814 ();
 sg13g2_decap_8 FILLER_37_821 ();
 sg13g2_decap_8 FILLER_37_828 ();
 sg13g2_decap_8 FILLER_37_835 ();
 sg13g2_decap_8 FILLER_37_842 ();
 sg13g2_decap_8 FILLER_37_849 ();
 sg13g2_decap_4 FILLER_37_856 ();
 sg13g2_fill_2 FILLER_37_860 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_fill_1 FILLER_38_77 ();
 sg13g2_decap_4 FILLER_38_104 ();
 sg13g2_fill_1 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_113 ();
 sg13g2_fill_2 FILLER_38_117 ();
 sg13g2_fill_1 FILLER_38_132 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_fill_2 FILLER_38_222 ();
 sg13g2_fill_1 FILLER_38_224 ();
 sg13g2_fill_2 FILLER_38_235 ();
 sg13g2_fill_1 FILLER_38_237 ();
 sg13g2_decap_4 FILLER_38_242 ();
 sg13g2_fill_2 FILLER_38_246 ();
 sg13g2_decap_4 FILLER_38_278 ();
 sg13g2_fill_2 FILLER_38_282 ();
 sg13g2_fill_2 FILLER_38_288 ();
 sg13g2_fill_2 FILLER_38_300 ();
 sg13g2_decap_4 FILLER_38_328 ();
 sg13g2_decap_8 FILLER_38_336 ();
 sg13g2_decap_8 FILLER_38_343 ();
 sg13g2_decap_4 FILLER_38_350 ();
 sg13g2_fill_1 FILLER_38_354 ();
 sg13g2_fill_1 FILLER_38_359 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_decap_8 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_38_414 ();
 sg13g2_decap_8 FILLER_38_421 ();
 sg13g2_decap_8 FILLER_38_428 ();
 sg13g2_decap_8 FILLER_38_435 ();
 sg13g2_decap_8 FILLER_38_442 ();
 sg13g2_decap_8 FILLER_38_449 ();
 sg13g2_decap_8 FILLER_38_456 ();
 sg13g2_decap_8 FILLER_38_463 ();
 sg13g2_decap_8 FILLER_38_470 ();
 sg13g2_decap_8 FILLER_38_477 ();
 sg13g2_decap_8 FILLER_38_484 ();
 sg13g2_decap_8 FILLER_38_491 ();
 sg13g2_decap_8 FILLER_38_498 ();
 sg13g2_decap_8 FILLER_38_505 ();
 sg13g2_decap_8 FILLER_38_512 ();
 sg13g2_decap_8 FILLER_38_519 ();
 sg13g2_decap_8 FILLER_38_526 ();
 sg13g2_decap_8 FILLER_38_533 ();
 sg13g2_decap_8 FILLER_38_540 ();
 sg13g2_decap_8 FILLER_38_547 ();
 sg13g2_decap_8 FILLER_38_554 ();
 sg13g2_decap_8 FILLER_38_561 ();
 sg13g2_decap_8 FILLER_38_568 ();
 sg13g2_decap_8 FILLER_38_575 ();
 sg13g2_decap_8 FILLER_38_582 ();
 sg13g2_decap_8 FILLER_38_589 ();
 sg13g2_decap_8 FILLER_38_596 ();
 sg13g2_decap_8 FILLER_38_603 ();
 sg13g2_decap_8 FILLER_38_610 ();
 sg13g2_decap_8 FILLER_38_617 ();
 sg13g2_decap_8 FILLER_38_624 ();
 sg13g2_decap_8 FILLER_38_631 ();
 sg13g2_decap_8 FILLER_38_638 ();
 sg13g2_decap_8 FILLER_38_645 ();
 sg13g2_decap_8 FILLER_38_652 ();
 sg13g2_decap_8 FILLER_38_659 ();
 sg13g2_decap_8 FILLER_38_666 ();
 sg13g2_decap_8 FILLER_38_673 ();
 sg13g2_decap_8 FILLER_38_680 ();
 sg13g2_decap_8 FILLER_38_687 ();
 sg13g2_decap_8 FILLER_38_694 ();
 sg13g2_decap_8 FILLER_38_701 ();
 sg13g2_decap_8 FILLER_38_708 ();
 sg13g2_decap_8 FILLER_38_715 ();
 sg13g2_decap_8 FILLER_38_722 ();
 sg13g2_decap_8 FILLER_38_729 ();
 sg13g2_decap_8 FILLER_38_736 ();
 sg13g2_decap_8 FILLER_38_743 ();
 sg13g2_decap_8 FILLER_38_750 ();
 sg13g2_decap_8 FILLER_38_757 ();
 sg13g2_decap_8 FILLER_38_764 ();
 sg13g2_decap_8 FILLER_38_771 ();
 sg13g2_decap_8 FILLER_38_778 ();
 sg13g2_decap_8 FILLER_38_785 ();
 sg13g2_decap_8 FILLER_38_792 ();
 sg13g2_decap_8 FILLER_38_799 ();
 sg13g2_decap_8 FILLER_38_806 ();
 sg13g2_decap_8 FILLER_38_813 ();
 sg13g2_decap_8 FILLER_38_820 ();
 sg13g2_decap_8 FILLER_38_827 ();
 sg13g2_decap_8 FILLER_38_834 ();
 sg13g2_decap_8 FILLER_38_841 ();
 sg13g2_decap_8 FILLER_38_848 ();
 sg13g2_decap_8 FILLER_38_855 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_fill_1 FILLER_39_70 ();
 sg13g2_fill_2 FILLER_39_89 ();
 sg13g2_fill_2 FILLER_39_96 ();
 sg13g2_fill_2 FILLER_39_124 ();
 sg13g2_fill_1 FILLER_39_126 ();
 sg13g2_fill_1 FILLER_39_132 ();
 sg13g2_fill_1 FILLER_39_147 ();
 sg13g2_fill_1 FILLER_39_180 ();
 sg13g2_fill_1 FILLER_39_226 ();
 sg13g2_fill_2 FILLER_39_266 ();
 sg13g2_fill_1 FILLER_39_268 ();
 sg13g2_decap_8 FILLER_39_284 ();
 sg13g2_fill_2 FILLER_39_291 ();
 sg13g2_fill_2 FILLER_39_327 ();
 sg13g2_fill_1 FILLER_39_343 ();
 sg13g2_fill_1 FILLER_39_370 ();
 sg13g2_fill_1 FILLER_39_375 ();
 sg13g2_decap_8 FILLER_39_402 ();
 sg13g2_decap_8 FILLER_39_409 ();
 sg13g2_decap_8 FILLER_39_416 ();
 sg13g2_decap_8 FILLER_39_423 ();
 sg13g2_decap_8 FILLER_39_430 ();
 sg13g2_decap_8 FILLER_39_437 ();
 sg13g2_decap_8 FILLER_39_444 ();
 sg13g2_decap_8 FILLER_39_451 ();
 sg13g2_decap_8 FILLER_39_458 ();
 sg13g2_decap_8 FILLER_39_465 ();
 sg13g2_decap_8 FILLER_39_472 ();
 sg13g2_decap_8 FILLER_39_479 ();
 sg13g2_decap_8 FILLER_39_486 ();
 sg13g2_decap_8 FILLER_39_493 ();
 sg13g2_decap_8 FILLER_39_500 ();
 sg13g2_decap_8 FILLER_39_507 ();
 sg13g2_decap_8 FILLER_39_514 ();
 sg13g2_decap_8 FILLER_39_521 ();
 sg13g2_decap_8 FILLER_39_528 ();
 sg13g2_decap_8 FILLER_39_535 ();
 sg13g2_decap_8 FILLER_39_542 ();
 sg13g2_decap_8 FILLER_39_549 ();
 sg13g2_decap_8 FILLER_39_556 ();
 sg13g2_decap_8 FILLER_39_563 ();
 sg13g2_decap_8 FILLER_39_570 ();
 sg13g2_decap_8 FILLER_39_577 ();
 sg13g2_decap_8 FILLER_39_584 ();
 sg13g2_decap_8 FILLER_39_591 ();
 sg13g2_decap_8 FILLER_39_598 ();
 sg13g2_decap_8 FILLER_39_605 ();
 sg13g2_decap_8 FILLER_39_612 ();
 sg13g2_decap_8 FILLER_39_619 ();
 sg13g2_decap_8 FILLER_39_626 ();
 sg13g2_decap_8 FILLER_39_633 ();
 sg13g2_decap_8 FILLER_39_640 ();
 sg13g2_decap_8 FILLER_39_647 ();
 sg13g2_decap_8 FILLER_39_654 ();
 sg13g2_decap_8 FILLER_39_661 ();
 sg13g2_decap_8 FILLER_39_668 ();
 sg13g2_decap_8 FILLER_39_675 ();
 sg13g2_decap_8 FILLER_39_682 ();
 sg13g2_decap_8 FILLER_39_689 ();
 sg13g2_decap_8 FILLER_39_696 ();
 sg13g2_decap_8 FILLER_39_703 ();
 sg13g2_decap_8 FILLER_39_710 ();
 sg13g2_decap_8 FILLER_39_717 ();
 sg13g2_decap_8 FILLER_39_724 ();
 sg13g2_decap_8 FILLER_39_731 ();
 sg13g2_decap_8 FILLER_39_738 ();
 sg13g2_decap_8 FILLER_39_745 ();
 sg13g2_decap_8 FILLER_39_752 ();
 sg13g2_decap_8 FILLER_39_759 ();
 sg13g2_decap_8 FILLER_39_766 ();
 sg13g2_decap_8 FILLER_39_773 ();
 sg13g2_decap_8 FILLER_39_780 ();
 sg13g2_decap_8 FILLER_39_787 ();
 sg13g2_decap_8 FILLER_39_794 ();
 sg13g2_decap_8 FILLER_39_801 ();
 sg13g2_decap_8 FILLER_39_808 ();
 sg13g2_decap_8 FILLER_39_815 ();
 sg13g2_decap_8 FILLER_39_822 ();
 sg13g2_decap_8 FILLER_39_829 ();
 sg13g2_decap_8 FILLER_39_836 ();
 sg13g2_decap_8 FILLER_39_843 ();
 sg13g2_decap_8 FILLER_39_850 ();
 sg13g2_decap_4 FILLER_39_857 ();
 sg13g2_fill_1 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_4 FILLER_40_42 ();
 sg13g2_fill_1 FILLER_40_80 ();
 sg13g2_fill_2 FILLER_40_171 ();
 sg13g2_fill_1 FILLER_40_195 ();
 sg13g2_fill_1 FILLER_40_221 ();
 sg13g2_fill_2 FILLER_40_259 ();
 sg13g2_fill_1 FILLER_40_275 ();
 sg13g2_decap_4 FILLER_40_302 ();
 sg13g2_fill_2 FILLER_40_306 ();
 sg13g2_decap_8 FILLER_40_354 ();
 sg13g2_decap_8 FILLER_40_365 ();
 sg13g2_decap_8 FILLER_40_372 ();
 sg13g2_fill_1 FILLER_40_384 ();
 sg13g2_decap_8 FILLER_40_415 ();
 sg13g2_decap_8 FILLER_40_422 ();
 sg13g2_decap_8 FILLER_40_429 ();
 sg13g2_decap_8 FILLER_40_436 ();
 sg13g2_decap_8 FILLER_40_443 ();
 sg13g2_decap_8 FILLER_40_450 ();
 sg13g2_decap_8 FILLER_40_457 ();
 sg13g2_decap_8 FILLER_40_464 ();
 sg13g2_decap_8 FILLER_40_471 ();
 sg13g2_decap_8 FILLER_40_478 ();
 sg13g2_decap_8 FILLER_40_485 ();
 sg13g2_decap_8 FILLER_40_492 ();
 sg13g2_decap_8 FILLER_40_499 ();
 sg13g2_decap_8 FILLER_40_506 ();
 sg13g2_decap_8 FILLER_40_513 ();
 sg13g2_decap_8 FILLER_40_520 ();
 sg13g2_decap_8 FILLER_40_527 ();
 sg13g2_decap_8 FILLER_40_534 ();
 sg13g2_decap_8 FILLER_40_541 ();
 sg13g2_decap_8 FILLER_40_548 ();
 sg13g2_decap_8 FILLER_40_555 ();
 sg13g2_decap_8 FILLER_40_562 ();
 sg13g2_decap_8 FILLER_40_569 ();
 sg13g2_decap_8 FILLER_40_576 ();
 sg13g2_decap_8 FILLER_40_583 ();
 sg13g2_decap_8 FILLER_40_590 ();
 sg13g2_decap_8 FILLER_40_597 ();
 sg13g2_decap_8 FILLER_40_604 ();
 sg13g2_decap_8 FILLER_40_611 ();
 sg13g2_decap_8 FILLER_40_618 ();
 sg13g2_decap_8 FILLER_40_625 ();
 sg13g2_decap_8 FILLER_40_632 ();
 sg13g2_decap_8 FILLER_40_639 ();
 sg13g2_decap_8 FILLER_40_646 ();
 sg13g2_decap_8 FILLER_40_653 ();
 sg13g2_decap_8 FILLER_40_660 ();
 sg13g2_decap_8 FILLER_40_667 ();
 sg13g2_decap_8 FILLER_40_674 ();
 sg13g2_decap_8 FILLER_40_681 ();
 sg13g2_decap_8 FILLER_40_688 ();
 sg13g2_decap_8 FILLER_40_695 ();
 sg13g2_decap_8 FILLER_40_702 ();
 sg13g2_decap_8 FILLER_40_709 ();
 sg13g2_decap_8 FILLER_40_716 ();
 sg13g2_decap_8 FILLER_40_723 ();
 sg13g2_decap_8 FILLER_40_730 ();
 sg13g2_decap_8 FILLER_40_737 ();
 sg13g2_decap_8 FILLER_40_744 ();
 sg13g2_decap_8 FILLER_40_751 ();
 sg13g2_decap_8 FILLER_40_758 ();
 sg13g2_decap_8 FILLER_40_765 ();
 sg13g2_decap_8 FILLER_40_772 ();
 sg13g2_decap_8 FILLER_40_779 ();
 sg13g2_decap_8 FILLER_40_786 ();
 sg13g2_decap_8 FILLER_40_793 ();
 sg13g2_decap_8 FILLER_40_800 ();
 sg13g2_decap_8 FILLER_40_807 ();
 sg13g2_decap_8 FILLER_40_814 ();
 sg13g2_decap_8 FILLER_40_821 ();
 sg13g2_decap_8 FILLER_40_828 ();
 sg13g2_decap_8 FILLER_40_835 ();
 sg13g2_decap_8 FILLER_40_842 ();
 sg13g2_decap_8 FILLER_40_849 ();
 sg13g2_decap_4 FILLER_40_856 ();
 sg13g2_fill_2 FILLER_40_860 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_fill_2 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_fill_1 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_48 ();
 sg13g2_fill_2 FILLER_41_55 ();
 sg13g2_fill_1 FILLER_41_57 ();
 sg13g2_fill_1 FILLER_41_67 ();
 sg13g2_fill_1 FILLER_41_72 ();
 sg13g2_fill_1 FILLER_41_86 ();
 sg13g2_fill_1 FILLER_41_150 ();
 sg13g2_fill_1 FILLER_41_176 ();
 sg13g2_fill_2 FILLER_41_244 ();
 sg13g2_fill_1 FILLER_41_246 ();
 sg13g2_decap_8 FILLER_41_252 ();
 sg13g2_fill_2 FILLER_41_284 ();
 sg13g2_fill_1 FILLER_41_286 ();
 sg13g2_fill_2 FILLER_41_291 ();
 sg13g2_fill_2 FILLER_41_302 ();
 sg13g2_fill_2 FILLER_41_308 ();
 sg13g2_fill_1 FILLER_41_310 ();
 sg13g2_fill_2 FILLER_41_315 ();
 sg13g2_decap_4 FILLER_41_324 ();
 sg13g2_fill_2 FILLER_41_333 ();
 sg13g2_fill_1 FILLER_41_335 ();
 sg13g2_decap_4 FILLER_41_376 ();
 sg13g2_fill_2 FILLER_41_380 ();
 sg13g2_decap_8 FILLER_41_386 ();
 sg13g2_decap_8 FILLER_41_393 ();
 sg13g2_decap_4 FILLER_41_400 ();
 sg13g2_fill_2 FILLER_41_430 ();
 sg13g2_fill_1 FILLER_41_432 ();
 sg13g2_decap_8 FILLER_41_437 ();
 sg13g2_decap_8 FILLER_41_444 ();
 sg13g2_decap_8 FILLER_41_451 ();
 sg13g2_decap_8 FILLER_41_458 ();
 sg13g2_decap_8 FILLER_41_465 ();
 sg13g2_decap_8 FILLER_41_472 ();
 sg13g2_decap_8 FILLER_41_479 ();
 sg13g2_decap_8 FILLER_41_486 ();
 sg13g2_decap_8 FILLER_41_493 ();
 sg13g2_decap_8 FILLER_41_500 ();
 sg13g2_decap_8 FILLER_41_507 ();
 sg13g2_decap_8 FILLER_41_514 ();
 sg13g2_decap_8 FILLER_41_521 ();
 sg13g2_decap_8 FILLER_41_528 ();
 sg13g2_decap_8 FILLER_41_535 ();
 sg13g2_decap_8 FILLER_41_542 ();
 sg13g2_decap_8 FILLER_41_549 ();
 sg13g2_decap_8 FILLER_41_556 ();
 sg13g2_decap_8 FILLER_41_563 ();
 sg13g2_decap_8 FILLER_41_570 ();
 sg13g2_decap_8 FILLER_41_577 ();
 sg13g2_decap_8 FILLER_41_584 ();
 sg13g2_decap_8 FILLER_41_591 ();
 sg13g2_decap_8 FILLER_41_598 ();
 sg13g2_decap_8 FILLER_41_605 ();
 sg13g2_decap_8 FILLER_41_612 ();
 sg13g2_decap_8 FILLER_41_619 ();
 sg13g2_decap_8 FILLER_41_626 ();
 sg13g2_decap_8 FILLER_41_633 ();
 sg13g2_decap_8 FILLER_41_640 ();
 sg13g2_decap_8 FILLER_41_647 ();
 sg13g2_decap_8 FILLER_41_654 ();
 sg13g2_decap_8 FILLER_41_661 ();
 sg13g2_decap_8 FILLER_41_668 ();
 sg13g2_decap_8 FILLER_41_675 ();
 sg13g2_decap_8 FILLER_41_682 ();
 sg13g2_decap_8 FILLER_41_689 ();
 sg13g2_decap_8 FILLER_41_696 ();
 sg13g2_decap_8 FILLER_41_703 ();
 sg13g2_decap_8 FILLER_41_710 ();
 sg13g2_decap_8 FILLER_41_717 ();
 sg13g2_decap_8 FILLER_41_724 ();
 sg13g2_decap_8 FILLER_41_731 ();
 sg13g2_decap_8 FILLER_41_738 ();
 sg13g2_decap_8 FILLER_41_745 ();
 sg13g2_decap_8 FILLER_41_752 ();
 sg13g2_decap_8 FILLER_41_759 ();
 sg13g2_decap_8 FILLER_41_766 ();
 sg13g2_decap_8 FILLER_41_773 ();
 sg13g2_decap_8 FILLER_41_780 ();
 sg13g2_decap_8 FILLER_41_787 ();
 sg13g2_decap_8 FILLER_41_794 ();
 sg13g2_decap_8 FILLER_41_801 ();
 sg13g2_decap_8 FILLER_41_808 ();
 sg13g2_decap_8 FILLER_41_815 ();
 sg13g2_decap_8 FILLER_41_822 ();
 sg13g2_decap_8 FILLER_41_829 ();
 sg13g2_decap_8 FILLER_41_836 ();
 sg13g2_decap_8 FILLER_41_843 ();
 sg13g2_decap_8 FILLER_41_850 ();
 sg13g2_decap_4 FILLER_41_857 ();
 sg13g2_fill_1 FILLER_41_861 ();
 sg13g2_fill_1 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_41 ();
 sg13g2_fill_2 FILLER_42_69 ();
 sg13g2_fill_1 FILLER_42_79 ();
 sg13g2_fill_2 FILLER_42_87 ();
 sg13g2_fill_1 FILLER_42_100 ();
 sg13g2_decap_4 FILLER_42_114 ();
 sg13g2_fill_2 FILLER_42_140 ();
 sg13g2_fill_1 FILLER_42_142 ();
 sg13g2_decap_4 FILLER_42_159 ();
 sg13g2_fill_2 FILLER_42_163 ();
 sg13g2_fill_1 FILLER_42_175 ();
 sg13g2_fill_2 FILLER_42_195 ();
 sg13g2_fill_1 FILLER_42_197 ();
 sg13g2_decap_8 FILLER_42_202 ();
 sg13g2_fill_1 FILLER_42_209 ();
 sg13g2_decap_4 FILLER_42_263 ();
 sg13g2_fill_1 FILLER_42_267 ();
 sg13g2_decap_4 FILLER_42_276 ();
 sg13g2_fill_2 FILLER_42_303 ();
 sg13g2_fill_1 FILLER_42_310 ();
 sg13g2_fill_2 FILLER_42_316 ();
 sg13g2_fill_2 FILLER_42_337 ();
 sg13g2_fill_1 FILLER_42_339 ();
 sg13g2_fill_1 FILLER_42_345 ();
 sg13g2_fill_2 FILLER_42_356 ();
 sg13g2_decap_4 FILLER_42_366 ();
 sg13g2_fill_1 FILLER_42_370 ();
 sg13g2_fill_2 FILLER_42_397 ();
 sg13g2_fill_1 FILLER_42_399 ();
 sg13g2_decap_8 FILLER_42_404 ();
 sg13g2_decap_4 FILLER_42_411 ();
 sg13g2_fill_2 FILLER_42_419 ();
 sg13g2_fill_1 FILLER_42_421 ();
 sg13g2_decap_8 FILLER_42_448 ();
 sg13g2_decap_8 FILLER_42_455 ();
 sg13g2_decap_8 FILLER_42_462 ();
 sg13g2_decap_8 FILLER_42_469 ();
 sg13g2_decap_8 FILLER_42_476 ();
 sg13g2_decap_8 FILLER_42_483 ();
 sg13g2_decap_8 FILLER_42_490 ();
 sg13g2_decap_8 FILLER_42_497 ();
 sg13g2_decap_8 FILLER_42_504 ();
 sg13g2_decap_8 FILLER_42_511 ();
 sg13g2_decap_8 FILLER_42_518 ();
 sg13g2_decap_8 FILLER_42_525 ();
 sg13g2_decap_8 FILLER_42_532 ();
 sg13g2_decap_8 FILLER_42_539 ();
 sg13g2_decap_8 FILLER_42_546 ();
 sg13g2_decap_8 FILLER_42_553 ();
 sg13g2_decap_8 FILLER_42_560 ();
 sg13g2_decap_8 FILLER_42_567 ();
 sg13g2_decap_8 FILLER_42_574 ();
 sg13g2_decap_8 FILLER_42_581 ();
 sg13g2_decap_8 FILLER_42_588 ();
 sg13g2_decap_8 FILLER_42_595 ();
 sg13g2_decap_8 FILLER_42_602 ();
 sg13g2_decap_8 FILLER_42_609 ();
 sg13g2_decap_8 FILLER_42_616 ();
 sg13g2_decap_8 FILLER_42_623 ();
 sg13g2_decap_8 FILLER_42_630 ();
 sg13g2_decap_8 FILLER_42_637 ();
 sg13g2_decap_8 FILLER_42_644 ();
 sg13g2_decap_8 FILLER_42_651 ();
 sg13g2_decap_8 FILLER_42_658 ();
 sg13g2_decap_8 FILLER_42_665 ();
 sg13g2_decap_8 FILLER_42_672 ();
 sg13g2_decap_8 FILLER_42_679 ();
 sg13g2_decap_8 FILLER_42_686 ();
 sg13g2_decap_8 FILLER_42_693 ();
 sg13g2_decap_8 FILLER_42_700 ();
 sg13g2_decap_8 FILLER_42_707 ();
 sg13g2_decap_8 FILLER_42_714 ();
 sg13g2_decap_8 FILLER_42_721 ();
 sg13g2_decap_8 FILLER_42_728 ();
 sg13g2_decap_8 FILLER_42_735 ();
 sg13g2_decap_8 FILLER_42_742 ();
 sg13g2_decap_8 FILLER_42_749 ();
 sg13g2_decap_8 FILLER_42_756 ();
 sg13g2_decap_8 FILLER_42_763 ();
 sg13g2_decap_8 FILLER_42_770 ();
 sg13g2_decap_8 FILLER_42_777 ();
 sg13g2_decap_8 FILLER_42_784 ();
 sg13g2_decap_8 FILLER_42_791 ();
 sg13g2_decap_8 FILLER_42_798 ();
 sg13g2_decap_8 FILLER_42_805 ();
 sg13g2_decap_8 FILLER_42_812 ();
 sg13g2_decap_8 FILLER_42_819 ();
 sg13g2_decap_8 FILLER_42_826 ();
 sg13g2_decap_8 FILLER_42_833 ();
 sg13g2_decap_8 FILLER_42_840 ();
 sg13g2_decap_8 FILLER_42_847 ();
 sg13g2_decap_8 FILLER_42_854 ();
 sg13g2_fill_1 FILLER_42_861 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_7 ();
 sg13g2_fill_2 FILLER_43_16 ();
 sg13g2_fill_2 FILLER_43_35 ();
 sg13g2_fill_1 FILLER_43_37 ();
 sg13g2_fill_1 FILLER_43_61 ();
 sg13g2_fill_2 FILLER_43_115 ();
 sg13g2_decap_4 FILLER_43_152 ();
 sg13g2_fill_2 FILLER_43_156 ();
 sg13g2_fill_2 FILLER_43_218 ();
 sg13g2_fill_1 FILLER_43_220 ();
 sg13g2_fill_2 FILLER_43_255 ();
 sg13g2_fill_1 FILLER_43_257 ();
 sg13g2_fill_2 FILLER_43_293 ();
 sg13g2_fill_1 FILLER_43_295 ();
 sg13g2_decap_4 FILLER_43_325 ();
 sg13g2_decap_4 FILLER_43_333 ();
 sg13g2_decap_8 FILLER_43_341 ();
 sg13g2_decap_4 FILLER_43_348 ();
 sg13g2_decap_4 FILLER_43_360 ();
 sg13g2_fill_2 FILLER_43_364 ();
 sg13g2_decap_4 FILLER_43_375 ();
 sg13g2_fill_2 FILLER_43_379 ();
 sg13g2_decap_4 FILLER_43_407 ();
 sg13g2_decap_8 FILLER_43_415 ();
 sg13g2_decap_4 FILLER_43_431 ();
 sg13g2_fill_1 FILLER_43_435 ();
 sg13g2_decap_8 FILLER_43_462 ();
 sg13g2_decap_8 FILLER_43_469 ();
 sg13g2_decap_8 FILLER_43_476 ();
 sg13g2_decap_8 FILLER_43_483 ();
 sg13g2_decap_4 FILLER_43_490 ();
 sg13g2_decap_8 FILLER_43_498 ();
 sg13g2_decap_8 FILLER_43_505 ();
 sg13g2_decap_8 FILLER_43_512 ();
 sg13g2_decap_8 FILLER_43_545 ();
 sg13g2_decap_8 FILLER_43_552 ();
 sg13g2_fill_2 FILLER_43_559 ();
 sg13g2_fill_1 FILLER_43_561 ();
 sg13g2_fill_1 FILLER_43_566 ();
 sg13g2_decap_8 FILLER_43_572 ();
 sg13g2_fill_2 FILLER_43_579 ();
 sg13g2_decap_8 FILLER_43_607 ();
 sg13g2_decap_8 FILLER_43_614 ();
 sg13g2_decap_8 FILLER_43_621 ();
 sg13g2_decap_8 FILLER_43_628 ();
 sg13g2_decap_8 FILLER_43_635 ();
 sg13g2_decap_8 FILLER_43_642 ();
 sg13g2_decap_8 FILLER_43_649 ();
 sg13g2_decap_8 FILLER_43_656 ();
 sg13g2_decap_8 FILLER_43_663 ();
 sg13g2_decap_8 FILLER_43_670 ();
 sg13g2_decap_8 FILLER_43_677 ();
 sg13g2_decap_8 FILLER_43_684 ();
 sg13g2_decap_8 FILLER_43_691 ();
 sg13g2_decap_8 FILLER_43_698 ();
 sg13g2_decap_8 FILLER_43_705 ();
 sg13g2_decap_8 FILLER_43_712 ();
 sg13g2_decap_8 FILLER_43_719 ();
 sg13g2_decap_8 FILLER_43_726 ();
 sg13g2_decap_8 FILLER_43_733 ();
 sg13g2_decap_8 FILLER_43_740 ();
 sg13g2_decap_8 FILLER_43_747 ();
 sg13g2_decap_8 FILLER_43_754 ();
 sg13g2_decap_8 FILLER_43_761 ();
 sg13g2_decap_8 FILLER_43_768 ();
 sg13g2_decap_8 FILLER_43_775 ();
 sg13g2_decap_8 FILLER_43_782 ();
 sg13g2_decap_8 FILLER_43_789 ();
 sg13g2_decap_8 FILLER_43_796 ();
 sg13g2_decap_8 FILLER_43_803 ();
 sg13g2_decap_8 FILLER_43_810 ();
 sg13g2_decap_8 FILLER_43_817 ();
 sg13g2_decap_8 FILLER_43_824 ();
 sg13g2_decap_8 FILLER_43_831 ();
 sg13g2_decap_8 FILLER_43_838 ();
 sg13g2_decap_8 FILLER_43_845 ();
 sg13g2_decap_8 FILLER_43_852 ();
 sg13g2_fill_2 FILLER_43_859 ();
 sg13g2_fill_1 FILLER_43_861 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_33 ();
 sg13g2_fill_2 FILLER_44_40 ();
 sg13g2_fill_2 FILLER_44_63 ();
 sg13g2_fill_1 FILLER_44_65 ();
 sg13g2_decap_8 FILLER_44_109 ();
 sg13g2_decap_4 FILLER_44_116 ();
 sg13g2_fill_1 FILLER_44_120 ();
 sg13g2_decap_4 FILLER_44_126 ();
 sg13g2_fill_1 FILLER_44_130 ();
 sg13g2_fill_2 FILLER_44_144 ();
 sg13g2_decap_8 FILLER_44_150 ();
 sg13g2_decap_4 FILLER_44_157 ();
 sg13g2_fill_2 FILLER_44_161 ();
 sg13g2_decap_4 FILLER_44_193 ();
 sg13g2_fill_2 FILLER_44_227 ();
 sg13g2_fill_1 FILLER_44_229 ();
 sg13g2_fill_1 FILLER_44_235 ();
 sg13g2_decap_8 FILLER_44_269 ();
 sg13g2_decap_8 FILLER_44_276 ();
 sg13g2_fill_2 FILLER_44_292 ();
 sg13g2_fill_1 FILLER_44_299 ();
 sg13g2_fill_1 FILLER_44_305 ();
 sg13g2_fill_2 FILLER_44_311 ();
 sg13g2_fill_1 FILLER_44_313 ();
 sg13g2_fill_2 FILLER_44_353 ();
 sg13g2_decap_8 FILLER_44_385 ();
 sg13g2_decap_4 FILLER_44_396 ();
 sg13g2_fill_2 FILLER_44_426 ();
 sg13g2_decap_8 FILLER_44_458 ();
 sg13g2_fill_2 FILLER_44_465 ();
 sg13g2_fill_1 FILLER_44_467 ();
 sg13g2_decap_8 FILLER_44_472 ();
 sg13g2_decap_4 FILLER_44_479 ();
 sg13g2_decap_8 FILLER_44_539 ();
 sg13g2_decap_4 FILLER_44_546 ();
 sg13g2_fill_1 FILLER_44_550 ();
 sg13g2_fill_2 FILLER_44_591 ();
 sg13g2_decap_8 FILLER_44_615 ();
 sg13g2_decap_4 FILLER_44_627 ();
 sg13g2_decap_8 FILLER_44_635 ();
 sg13g2_decap_8 FILLER_44_642 ();
 sg13g2_decap_8 FILLER_44_649 ();
 sg13g2_decap_8 FILLER_44_656 ();
 sg13g2_decap_8 FILLER_44_663 ();
 sg13g2_decap_8 FILLER_44_670 ();
 sg13g2_decap_8 FILLER_44_677 ();
 sg13g2_decap_8 FILLER_44_684 ();
 sg13g2_decap_8 FILLER_44_691 ();
 sg13g2_decap_8 FILLER_44_698 ();
 sg13g2_decap_8 FILLER_44_705 ();
 sg13g2_decap_8 FILLER_44_712 ();
 sg13g2_decap_8 FILLER_44_719 ();
 sg13g2_decap_8 FILLER_44_726 ();
 sg13g2_decap_8 FILLER_44_733 ();
 sg13g2_decap_8 FILLER_44_740 ();
 sg13g2_decap_8 FILLER_44_747 ();
 sg13g2_decap_8 FILLER_44_754 ();
 sg13g2_decap_8 FILLER_44_761 ();
 sg13g2_decap_8 FILLER_44_768 ();
 sg13g2_decap_8 FILLER_44_775 ();
 sg13g2_decap_8 FILLER_44_782 ();
 sg13g2_decap_8 FILLER_44_789 ();
 sg13g2_decap_8 FILLER_44_796 ();
 sg13g2_decap_8 FILLER_44_803 ();
 sg13g2_decap_8 FILLER_44_810 ();
 sg13g2_decap_8 FILLER_44_817 ();
 sg13g2_decap_8 FILLER_44_824 ();
 sg13g2_decap_8 FILLER_44_831 ();
 sg13g2_decap_8 FILLER_44_838 ();
 sg13g2_decap_8 FILLER_44_845 ();
 sg13g2_decap_8 FILLER_44_852 ();
 sg13g2_fill_2 FILLER_44_859 ();
 sg13g2_fill_1 FILLER_44_861 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_37 ();
 sg13g2_fill_1 FILLER_45_39 ();
 sg13g2_fill_1 FILLER_45_57 ();
 sg13g2_fill_1 FILLER_45_108 ();
 sg13g2_decap_4 FILLER_45_120 ();
 sg13g2_decap_8 FILLER_45_185 ();
 sg13g2_fill_2 FILLER_45_192 ();
 sg13g2_fill_1 FILLER_45_194 ();
 sg13g2_decap_8 FILLER_45_199 ();
 sg13g2_decap_8 FILLER_45_206 ();
 sg13g2_fill_1 FILLER_45_227 ();
 sg13g2_fill_2 FILLER_45_246 ();
 sg13g2_decap_4 FILLER_45_301 ();
 sg13g2_fill_2 FILLER_45_305 ();
 sg13g2_fill_1 FILLER_45_321 ();
 sg13g2_decap_8 FILLER_45_326 ();
 sg13g2_decap_4 FILLER_45_333 ();
 sg13g2_decap_4 FILLER_45_341 ();
 sg13g2_fill_1 FILLER_45_345 ();
 sg13g2_fill_1 FILLER_45_354 ();
 sg13g2_fill_2 FILLER_45_367 ();
 sg13g2_fill_1 FILLER_45_369 ();
 sg13g2_fill_1 FILLER_45_374 ();
 sg13g2_decap_8 FILLER_45_379 ();
 sg13g2_decap_8 FILLER_45_386 ();
 sg13g2_decap_8 FILLER_45_393 ();
 sg13g2_fill_2 FILLER_45_412 ();
 sg13g2_fill_1 FILLER_45_430 ();
 sg13g2_decap_4 FILLER_45_435 ();
 sg13g2_decap_8 FILLER_45_443 ();
 sg13g2_decap_8 FILLER_45_450 ();
 sg13g2_decap_4 FILLER_45_483 ();
 sg13g2_fill_1 FILLER_45_487 ();
 sg13g2_fill_2 FILLER_45_517 ();
 sg13g2_fill_1 FILLER_45_528 ();
 sg13g2_fill_2 FILLER_45_542 ();
 sg13g2_fill_1 FILLER_45_615 ();
 sg13g2_fill_1 FILLER_45_642 ();
 sg13g2_decap_8 FILLER_45_661 ();
 sg13g2_decap_8 FILLER_45_668 ();
 sg13g2_decap_8 FILLER_45_675 ();
 sg13g2_decap_8 FILLER_45_682 ();
 sg13g2_decap_8 FILLER_45_689 ();
 sg13g2_decap_8 FILLER_45_696 ();
 sg13g2_decap_8 FILLER_45_703 ();
 sg13g2_decap_8 FILLER_45_710 ();
 sg13g2_decap_8 FILLER_45_717 ();
 sg13g2_decap_8 FILLER_45_724 ();
 sg13g2_decap_8 FILLER_45_731 ();
 sg13g2_decap_8 FILLER_45_738 ();
 sg13g2_decap_8 FILLER_45_745 ();
 sg13g2_decap_8 FILLER_45_752 ();
 sg13g2_decap_8 FILLER_45_759 ();
 sg13g2_decap_8 FILLER_45_766 ();
 sg13g2_decap_8 FILLER_45_773 ();
 sg13g2_decap_8 FILLER_45_780 ();
 sg13g2_decap_8 FILLER_45_787 ();
 sg13g2_decap_8 FILLER_45_794 ();
 sg13g2_decap_8 FILLER_45_801 ();
 sg13g2_decap_8 FILLER_45_808 ();
 sg13g2_decap_8 FILLER_45_815 ();
 sg13g2_decap_8 FILLER_45_822 ();
 sg13g2_decap_8 FILLER_45_829 ();
 sg13g2_decap_8 FILLER_45_836 ();
 sg13g2_decap_8 FILLER_45_843 ();
 sg13g2_decap_8 FILLER_45_850 ();
 sg13g2_decap_4 FILLER_45_857 ();
 sg13g2_fill_1 FILLER_45_861 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_decap_4 FILLER_46_57 ();
 sg13g2_fill_2 FILLER_46_69 ();
 sg13g2_fill_1 FILLER_46_81 ();
 sg13g2_fill_1 FILLER_46_87 ();
 sg13g2_fill_2 FILLER_46_146 ();
 sg13g2_decap_8 FILLER_46_152 ();
 sg13g2_decap_4 FILLER_46_169 ();
 sg13g2_fill_1 FILLER_46_173 ();
 sg13g2_fill_2 FILLER_46_218 ();
 sg13g2_decap_8 FILLER_46_250 ();
 sg13g2_fill_1 FILLER_46_257 ();
 sg13g2_fill_2 FILLER_46_266 ();
 sg13g2_fill_1 FILLER_46_268 ();
 sg13g2_decap_4 FILLER_46_272 ();
 sg13g2_fill_2 FILLER_46_276 ();
 sg13g2_decap_8 FILLER_46_282 ();
 sg13g2_decap_8 FILLER_46_289 ();
 sg13g2_fill_2 FILLER_46_308 ();
 sg13g2_fill_1 FILLER_46_310 ();
 sg13g2_fill_1 FILLER_46_341 ();
 sg13g2_fill_2 FILLER_46_348 ();
 sg13g2_fill_1 FILLER_46_360 ();
 sg13g2_fill_2 FILLER_46_385 ();
 sg13g2_fill_1 FILLER_46_387 ();
 sg13g2_fill_1 FILLER_46_414 ();
 sg13g2_decap_4 FILLER_46_447 ();
 sg13g2_fill_1 FILLER_46_451 ();
 sg13g2_fill_2 FILLER_46_457 ();
 sg13g2_fill_2 FILLER_46_469 ();
 sg13g2_fill_1 FILLER_46_471 ();
 sg13g2_fill_2 FILLER_46_481 ();
 sg13g2_fill_2 FILLER_46_505 ();
 sg13g2_decap_4 FILLER_46_552 ();
 sg13g2_fill_1 FILLER_46_561 ();
 sg13g2_decap_4 FILLER_46_593 ();
 sg13g2_fill_2 FILLER_46_597 ();
 sg13g2_decap_4 FILLER_46_608 ();
 sg13g2_fill_1 FILLER_46_644 ();
 sg13g2_decap_8 FILLER_46_671 ();
 sg13g2_decap_8 FILLER_46_678 ();
 sg13g2_decap_8 FILLER_46_685 ();
 sg13g2_decap_8 FILLER_46_692 ();
 sg13g2_decap_8 FILLER_46_699 ();
 sg13g2_decap_8 FILLER_46_706 ();
 sg13g2_decap_8 FILLER_46_713 ();
 sg13g2_decap_8 FILLER_46_720 ();
 sg13g2_decap_8 FILLER_46_727 ();
 sg13g2_decap_8 FILLER_46_734 ();
 sg13g2_decap_8 FILLER_46_741 ();
 sg13g2_decap_8 FILLER_46_748 ();
 sg13g2_decap_8 FILLER_46_755 ();
 sg13g2_decap_8 FILLER_46_762 ();
 sg13g2_decap_8 FILLER_46_769 ();
 sg13g2_decap_8 FILLER_46_776 ();
 sg13g2_decap_8 FILLER_46_783 ();
 sg13g2_decap_8 FILLER_46_790 ();
 sg13g2_decap_8 FILLER_46_797 ();
 sg13g2_decap_8 FILLER_46_804 ();
 sg13g2_decap_8 FILLER_46_811 ();
 sg13g2_decap_8 FILLER_46_818 ();
 sg13g2_decap_8 FILLER_46_825 ();
 sg13g2_decap_8 FILLER_46_832 ();
 sg13g2_decap_8 FILLER_46_839 ();
 sg13g2_decap_8 FILLER_46_846 ();
 sg13g2_decap_8 FILLER_46_853 ();
 sg13g2_fill_2 FILLER_46_860 ();
 sg13g2_fill_2 FILLER_47_26 ();
 sg13g2_fill_2 FILLER_47_37 ();
 sg13g2_fill_1 FILLER_47_62 ();
 sg13g2_fill_1 FILLER_47_68 ();
 sg13g2_decap_8 FILLER_47_92 ();
 sg13g2_decap_4 FILLER_47_99 ();
 sg13g2_fill_2 FILLER_47_103 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_fill_1 FILLER_47_126 ();
 sg13g2_decap_4 FILLER_47_152 ();
 sg13g2_fill_2 FILLER_47_176 ();
 sg13g2_fill_2 FILLER_47_183 ();
 sg13g2_decap_8 FILLER_47_198 ();
 sg13g2_decap_4 FILLER_47_205 ();
 sg13g2_fill_2 FILLER_47_234 ();
 sg13g2_fill_1 FILLER_47_236 ();
 sg13g2_fill_1 FILLER_47_249 ();
 sg13g2_fill_2 FILLER_47_284 ();
 sg13g2_fill_1 FILLER_47_286 ();
 sg13g2_decap_4 FILLER_47_291 ();
 sg13g2_fill_1 FILLER_47_295 ();
 sg13g2_decap_4 FILLER_47_319 ();
 sg13g2_decap_8 FILLER_47_330 ();
 sg13g2_decap_4 FILLER_47_337 ();
 sg13g2_fill_1 FILLER_47_341 ();
 sg13g2_fill_2 FILLER_47_354 ();
 sg13g2_fill_2 FILLER_47_366 ();
 sg13g2_fill_1 FILLER_47_368 ();
 sg13g2_decap_8 FILLER_47_373 ();
 sg13g2_fill_2 FILLER_47_380 ();
 sg13g2_decap_4 FILLER_47_394 ();
 sg13g2_fill_1 FILLER_47_402 ();
 sg13g2_fill_1 FILLER_47_407 ();
 sg13g2_decap_8 FILLER_47_412 ();
 sg13g2_fill_2 FILLER_47_419 ();
 sg13g2_fill_2 FILLER_47_426 ();
 sg13g2_fill_1 FILLER_47_428 ();
 sg13g2_fill_2 FILLER_47_448 ();
 sg13g2_fill_2 FILLER_47_459 ();
 sg13g2_fill_2 FILLER_47_476 ();
 sg13g2_fill_2 FILLER_47_550 ();
 sg13g2_fill_1 FILLER_47_552 ();
 sg13g2_fill_1 FILLER_47_579 ();
 sg13g2_fill_2 FILLER_47_611 ();
 sg13g2_fill_1 FILLER_47_613 ();
 sg13g2_fill_2 FILLER_47_645 ();
 sg13g2_fill_2 FILLER_47_652 ();
 sg13g2_decap_8 FILLER_47_680 ();
 sg13g2_decap_8 FILLER_47_687 ();
 sg13g2_decap_8 FILLER_47_694 ();
 sg13g2_decap_8 FILLER_47_701 ();
 sg13g2_decap_8 FILLER_47_708 ();
 sg13g2_decap_8 FILLER_47_715 ();
 sg13g2_decap_8 FILLER_47_722 ();
 sg13g2_decap_8 FILLER_47_729 ();
 sg13g2_decap_8 FILLER_47_736 ();
 sg13g2_decap_8 FILLER_47_743 ();
 sg13g2_decap_8 FILLER_47_750 ();
 sg13g2_decap_8 FILLER_47_757 ();
 sg13g2_decap_8 FILLER_47_764 ();
 sg13g2_decap_8 FILLER_47_771 ();
 sg13g2_decap_8 FILLER_47_778 ();
 sg13g2_decap_8 FILLER_47_785 ();
 sg13g2_decap_8 FILLER_47_792 ();
 sg13g2_decap_8 FILLER_47_799 ();
 sg13g2_decap_8 FILLER_47_806 ();
 sg13g2_decap_8 FILLER_47_813 ();
 sg13g2_decap_8 FILLER_47_820 ();
 sg13g2_decap_8 FILLER_47_827 ();
 sg13g2_decap_8 FILLER_47_834 ();
 sg13g2_decap_8 FILLER_47_841 ();
 sg13g2_decap_8 FILLER_47_848 ();
 sg13g2_decap_8 FILLER_47_855 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_7 ();
 sg13g2_fill_2 FILLER_48_17 ();
 sg13g2_fill_2 FILLER_48_39 ();
 sg13g2_fill_1 FILLER_48_59 ();
 sg13g2_fill_1 FILLER_48_70 ();
 sg13g2_fill_2 FILLER_48_97 ();
 sg13g2_fill_1 FILLER_48_99 ();
 sg13g2_decap_4 FILLER_48_130 ();
 sg13g2_fill_2 FILLER_48_134 ();
 sg13g2_fill_1 FILLER_48_142 ();
 sg13g2_fill_2 FILLER_48_148 ();
 sg13g2_fill_2 FILLER_48_168 ();
 sg13g2_fill_1 FILLER_48_170 ();
 sg13g2_fill_2 FILLER_48_176 ();
 sg13g2_fill_1 FILLER_48_178 ();
 sg13g2_fill_1 FILLER_48_203 ();
 sg13g2_fill_1 FILLER_48_235 ();
 sg13g2_decap_8 FILLER_48_318 ();
 sg13g2_fill_1 FILLER_48_325 ();
 sg13g2_decap_8 FILLER_48_342 ();
 sg13g2_fill_2 FILLER_48_363 ();
 sg13g2_fill_1 FILLER_48_365 ();
 sg13g2_fill_2 FILLER_48_371 ();
 sg13g2_fill_2 FILLER_48_381 ();
 sg13g2_fill_1 FILLER_48_389 ();
 sg13g2_decap_8 FILLER_48_413 ();
 sg13g2_decap_8 FILLER_48_425 ();
 sg13g2_decap_4 FILLER_48_432 ();
 sg13g2_fill_2 FILLER_48_436 ();
 sg13g2_fill_2 FILLER_48_446 ();
 sg13g2_decap_4 FILLER_48_471 ();
 sg13g2_fill_1 FILLER_48_475 ();
 sg13g2_decap_8 FILLER_48_503 ();
 sg13g2_fill_1 FILLER_48_510 ();
 sg13g2_fill_2 FILLER_48_562 ();
 sg13g2_fill_1 FILLER_48_564 ();
 sg13g2_fill_2 FILLER_48_579 ();
 sg13g2_fill_1 FILLER_48_595 ();
 sg13g2_decap_8 FILLER_48_600 ();
 sg13g2_fill_2 FILLER_48_607 ();
 sg13g2_fill_1 FILLER_48_645 ();
 sg13g2_decap_8 FILLER_48_681 ();
 sg13g2_decap_8 FILLER_48_688 ();
 sg13g2_fill_2 FILLER_48_695 ();
 sg13g2_decap_8 FILLER_48_701 ();
 sg13g2_decap_8 FILLER_48_708 ();
 sg13g2_decap_8 FILLER_48_715 ();
 sg13g2_decap_8 FILLER_48_722 ();
 sg13g2_decap_8 FILLER_48_729 ();
 sg13g2_decap_8 FILLER_48_736 ();
 sg13g2_decap_8 FILLER_48_743 ();
 sg13g2_decap_8 FILLER_48_750 ();
 sg13g2_decap_8 FILLER_48_757 ();
 sg13g2_decap_8 FILLER_48_764 ();
 sg13g2_decap_8 FILLER_48_771 ();
 sg13g2_decap_8 FILLER_48_778 ();
 sg13g2_decap_8 FILLER_48_785 ();
 sg13g2_decap_8 FILLER_48_792 ();
 sg13g2_decap_8 FILLER_48_799 ();
 sg13g2_decap_8 FILLER_48_806 ();
 sg13g2_decap_8 FILLER_48_813 ();
 sg13g2_decap_8 FILLER_48_820 ();
 sg13g2_decap_8 FILLER_48_827 ();
 sg13g2_decap_8 FILLER_48_834 ();
 sg13g2_decap_8 FILLER_48_841 ();
 sg13g2_decap_8 FILLER_48_848 ();
 sg13g2_decap_8 FILLER_48_855 ();
 sg13g2_decap_4 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_4 ();
 sg13g2_fill_2 FILLER_49_80 ();
 sg13g2_fill_2 FILLER_49_108 ();
 sg13g2_fill_1 FILLER_49_110 ();
 sg13g2_decap_4 FILLER_49_137 ();
 sg13g2_fill_2 FILLER_49_145 ();
 sg13g2_fill_1 FILLER_49_147 ();
 sg13g2_decap_8 FILLER_49_152 ();
 sg13g2_fill_2 FILLER_49_159 ();
 sg13g2_decap_4 FILLER_49_166 ();
 sg13g2_fill_1 FILLER_49_170 ();
 sg13g2_decap_8 FILLER_49_175 ();
 sg13g2_fill_2 FILLER_49_182 ();
 sg13g2_fill_1 FILLER_49_184 ();
 sg13g2_fill_2 FILLER_49_240 ();
 sg13g2_fill_2 FILLER_49_247 ();
 sg13g2_fill_1 FILLER_49_275 ();
 sg13g2_decap_8 FILLER_49_280 ();
 sg13g2_decap_8 FILLER_49_287 ();
 sg13g2_decap_8 FILLER_49_294 ();
 sg13g2_fill_2 FILLER_49_301 ();
 sg13g2_decap_4 FILLER_49_365 ();
 sg13g2_fill_2 FILLER_49_382 ();
 sg13g2_fill_2 FILLER_49_406 ();
 sg13g2_fill_2 FILLER_49_429 ();
 sg13g2_fill_1 FILLER_49_441 ();
 sg13g2_fill_2 FILLER_49_452 ();
 sg13g2_fill_1 FILLER_49_454 ();
 sg13g2_fill_1 FILLER_49_468 ();
 sg13g2_fill_2 FILLER_49_479 ();
 sg13g2_decap_8 FILLER_49_502 ();
 sg13g2_fill_2 FILLER_49_514 ();
 sg13g2_decap_4 FILLER_49_547 ();
 sg13g2_fill_1 FILLER_49_582 ();
 sg13g2_decap_4 FILLER_49_609 ();
 sg13g2_fill_1 FILLER_49_613 ();
 sg13g2_fill_2 FILLER_49_629 ();
 sg13g2_fill_1 FILLER_49_631 ();
 sg13g2_fill_2 FILLER_49_650 ();
 sg13g2_decap_8 FILLER_49_679 ();
 sg13g2_fill_2 FILLER_49_686 ();
 sg13g2_decap_4 FILLER_49_714 ();
 sg13g2_fill_1 FILLER_49_718 ();
 sg13g2_decap_8 FILLER_49_723 ();
 sg13g2_decap_8 FILLER_49_730 ();
 sg13g2_decap_8 FILLER_49_737 ();
 sg13g2_decap_8 FILLER_49_744 ();
 sg13g2_decap_8 FILLER_49_751 ();
 sg13g2_decap_8 FILLER_49_758 ();
 sg13g2_decap_8 FILLER_49_765 ();
 sg13g2_decap_8 FILLER_49_772 ();
 sg13g2_decap_8 FILLER_49_779 ();
 sg13g2_decap_8 FILLER_49_786 ();
 sg13g2_decap_8 FILLER_49_793 ();
 sg13g2_decap_8 FILLER_49_800 ();
 sg13g2_decap_8 FILLER_49_807 ();
 sg13g2_decap_8 FILLER_49_814 ();
 sg13g2_decap_8 FILLER_49_821 ();
 sg13g2_decap_8 FILLER_49_828 ();
 sg13g2_decap_8 FILLER_49_835 ();
 sg13g2_decap_8 FILLER_49_842 ();
 sg13g2_decap_8 FILLER_49_849 ();
 sg13g2_decap_4 FILLER_49_856 ();
 sg13g2_fill_2 FILLER_49_860 ();
 sg13g2_fill_1 FILLER_50_57 ();
 sg13g2_fill_2 FILLER_50_76 ();
 sg13g2_fill_1 FILLER_50_86 ();
 sg13g2_fill_2 FILLER_50_91 ();
 sg13g2_fill_2 FILLER_50_97 ();
 sg13g2_fill_1 FILLER_50_99 ();
 sg13g2_fill_1 FILLER_50_108 ();
 sg13g2_fill_2 FILLER_50_113 ();
 sg13g2_fill_1 FILLER_50_115 ();
 sg13g2_fill_1 FILLER_50_146 ();
 sg13g2_decap_8 FILLER_50_173 ();
 sg13g2_decap_8 FILLER_50_180 ();
 sg13g2_fill_2 FILLER_50_213 ();
 sg13g2_fill_1 FILLER_50_225 ();
 sg13g2_fill_2 FILLER_50_235 ();
 sg13g2_fill_2 FILLER_50_251 ();
 sg13g2_fill_2 FILLER_50_262 ();
 sg13g2_fill_1 FILLER_50_264 ();
 sg13g2_fill_2 FILLER_50_280 ();
 sg13g2_fill_1 FILLER_50_282 ();
 sg13g2_decap_4 FILLER_50_309 ();
 sg13g2_decap_8 FILLER_50_320 ();
 sg13g2_decap_4 FILLER_50_327 ();
 sg13g2_fill_2 FILLER_50_331 ();
 sg13g2_decap_8 FILLER_50_362 ();
 sg13g2_decap_8 FILLER_50_369 ();
 sg13g2_fill_2 FILLER_50_376 ();
 sg13g2_fill_1 FILLER_50_381 ();
 sg13g2_decap_4 FILLER_50_385 ();
 sg13g2_fill_1 FILLER_50_389 ();
 sg13g2_fill_1 FILLER_50_401 ();
 sg13g2_decap_8 FILLER_50_406 ();
 sg13g2_decap_8 FILLER_50_413 ();
 sg13g2_decap_8 FILLER_50_420 ();
 sg13g2_decap_8 FILLER_50_427 ();
 sg13g2_decap_4 FILLER_50_434 ();
 sg13g2_decap_4 FILLER_50_456 ();
 sg13g2_fill_1 FILLER_50_460 ();
 sg13g2_decap_4 FILLER_50_481 ();
 sg13g2_fill_2 FILLER_50_485 ();
 sg13g2_decap_4 FILLER_50_494 ();
 sg13g2_fill_1 FILLER_50_498 ();
 sg13g2_decap_8 FILLER_50_504 ();
 sg13g2_fill_2 FILLER_50_511 ();
 sg13g2_fill_1 FILLER_50_513 ();
 sg13g2_decap_4 FILLER_50_551 ();
 sg13g2_fill_1 FILLER_50_555 ();
 sg13g2_fill_1 FILLER_50_565 ();
 sg13g2_fill_2 FILLER_50_579 ();
 sg13g2_fill_2 FILLER_50_627 ();
 sg13g2_fill_2 FILLER_50_638 ();
 sg13g2_fill_1 FILLER_50_669 ();
 sg13g2_fill_2 FILLER_50_701 ();
 sg13g2_decap_8 FILLER_50_734 ();
 sg13g2_decap_8 FILLER_50_741 ();
 sg13g2_decap_8 FILLER_50_748 ();
 sg13g2_decap_8 FILLER_50_755 ();
 sg13g2_decap_8 FILLER_50_762 ();
 sg13g2_decap_8 FILLER_50_769 ();
 sg13g2_decap_8 FILLER_50_776 ();
 sg13g2_decap_8 FILLER_50_783 ();
 sg13g2_decap_8 FILLER_50_790 ();
 sg13g2_decap_8 FILLER_50_797 ();
 sg13g2_decap_8 FILLER_50_804 ();
 sg13g2_decap_8 FILLER_50_811 ();
 sg13g2_decap_8 FILLER_50_818 ();
 sg13g2_decap_8 FILLER_50_825 ();
 sg13g2_decap_8 FILLER_50_832 ();
 sg13g2_decap_8 FILLER_50_839 ();
 sg13g2_decap_8 FILLER_50_846 ();
 sg13g2_decap_8 FILLER_50_853 ();
 sg13g2_fill_2 FILLER_50_860 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_28 ();
 sg13g2_fill_1 FILLER_51_34 ();
 sg13g2_fill_2 FILLER_51_92 ();
 sg13g2_fill_1 FILLER_51_94 ();
 sg13g2_fill_1 FILLER_51_105 ();
 sg13g2_decap_4 FILLER_51_142 ();
 sg13g2_fill_1 FILLER_51_146 ();
 sg13g2_fill_1 FILLER_51_169 ();
 sg13g2_decap_4 FILLER_51_204 ();
 sg13g2_fill_1 FILLER_51_208 ();
 sg13g2_fill_2 FILLER_51_266 ();
 sg13g2_fill_1 FILLER_51_268 ();
 sg13g2_fill_1 FILLER_51_281 ();
 sg13g2_decap_8 FILLER_51_286 ();
 sg13g2_fill_1 FILLER_51_293 ();
 sg13g2_decap_8 FILLER_51_298 ();
 sg13g2_fill_2 FILLER_51_305 ();
 sg13g2_fill_2 FILLER_51_312 ();
 sg13g2_fill_1 FILLER_51_314 ();
 sg13g2_fill_2 FILLER_51_323 ();
 sg13g2_fill_1 FILLER_51_325 ();
 sg13g2_fill_1 FILLER_51_348 ();
 sg13g2_fill_2 FILLER_51_374 ();
 sg13g2_fill_1 FILLER_51_376 ();
 sg13g2_decap_4 FILLER_51_382 ();
 sg13g2_fill_1 FILLER_51_402 ();
 sg13g2_fill_2 FILLER_51_418 ();
 sg13g2_fill_1 FILLER_51_420 ();
 sg13g2_decap_8 FILLER_51_432 ();
 sg13g2_decap_4 FILLER_51_439 ();
 sg13g2_fill_2 FILLER_51_443 ();
 sg13g2_decap_4 FILLER_51_455 ();
 sg13g2_fill_1 FILLER_51_475 ();
 sg13g2_fill_1 FILLER_51_481 ();
 sg13g2_fill_1 FILLER_51_500 ();
 sg13g2_fill_1 FILLER_51_514 ();
 sg13g2_fill_1 FILLER_51_525 ();
 sg13g2_fill_1 FILLER_51_542 ();
 sg13g2_fill_2 FILLER_51_549 ();
 sg13g2_fill_1 FILLER_51_551 ();
 sg13g2_fill_2 FILLER_51_575 ();
 sg13g2_fill_1 FILLER_51_577 ();
 sg13g2_fill_2 FILLER_51_589 ();
 sg13g2_fill_2 FILLER_51_600 ();
 sg13g2_fill_1 FILLER_51_602 ();
 sg13g2_fill_2 FILLER_51_614 ();
 sg13g2_fill_2 FILLER_51_642 ();
 sg13g2_fill_2 FILLER_51_684 ();
 sg13g2_fill_1 FILLER_51_686 ();
 sg13g2_decap_8 FILLER_51_740 ();
 sg13g2_decap_8 FILLER_51_747 ();
 sg13g2_decap_8 FILLER_51_754 ();
 sg13g2_decap_8 FILLER_51_761 ();
 sg13g2_decap_8 FILLER_51_768 ();
 sg13g2_decap_8 FILLER_51_775 ();
 sg13g2_decap_8 FILLER_51_782 ();
 sg13g2_decap_8 FILLER_51_789 ();
 sg13g2_decap_8 FILLER_51_796 ();
 sg13g2_decap_8 FILLER_51_803 ();
 sg13g2_decap_8 FILLER_51_810 ();
 sg13g2_decap_8 FILLER_51_817 ();
 sg13g2_decap_8 FILLER_51_824 ();
 sg13g2_decap_8 FILLER_51_831 ();
 sg13g2_decap_8 FILLER_51_838 ();
 sg13g2_decap_8 FILLER_51_845 ();
 sg13g2_decap_8 FILLER_51_852 ();
 sg13g2_fill_2 FILLER_51_859 ();
 sg13g2_fill_1 FILLER_51_861 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_7 ();
 sg13g2_fill_1 FILLER_52_35 ();
 sg13g2_decap_4 FILLER_52_62 ();
 sg13g2_fill_1 FILLER_52_66 ();
 sg13g2_fill_2 FILLER_52_84 ();
 sg13g2_fill_1 FILLER_52_86 ();
 sg13g2_fill_2 FILLER_52_109 ();
 sg13g2_fill_1 FILLER_52_111 ();
 sg13g2_fill_2 FILLER_52_121 ();
 sg13g2_fill_1 FILLER_52_123 ();
 sg13g2_fill_2 FILLER_52_136 ();
 sg13g2_fill_1 FILLER_52_138 ();
 sg13g2_decap_8 FILLER_52_160 ();
 sg13g2_fill_1 FILLER_52_167 ();
 sg13g2_fill_1 FILLER_52_196 ();
 sg13g2_fill_2 FILLER_52_206 ();
 sg13g2_fill_2 FILLER_52_229 ();
 sg13g2_fill_1 FILLER_52_231 ();
 sg13g2_fill_2 FILLER_52_236 ();
 sg13g2_fill_1 FILLER_52_238 ();
 sg13g2_fill_1 FILLER_52_249 ();
 sg13g2_fill_2 FILLER_52_255 ();
 sg13g2_decap_4 FILLER_52_262 ();
 sg13g2_fill_2 FILLER_52_266 ();
 sg13g2_fill_2 FILLER_52_281 ();
 sg13g2_decap_4 FILLER_52_297 ();
 sg13g2_decap_8 FILLER_52_317 ();
 sg13g2_decap_8 FILLER_52_324 ();
 sg13g2_decap_4 FILLER_52_331 ();
 sg13g2_fill_1 FILLER_52_335 ();
 sg13g2_fill_2 FILLER_52_383 ();
 sg13g2_fill_2 FILLER_52_394 ();
 sg13g2_fill_1 FILLER_52_434 ();
 sg13g2_fill_2 FILLER_52_444 ();
 sg13g2_fill_1 FILLER_52_461 ();
 sg13g2_decap_4 FILLER_52_492 ();
 sg13g2_decap_8 FILLER_52_510 ();
 sg13g2_decap_8 FILLER_52_517 ();
 sg13g2_fill_2 FILLER_52_524 ();
 sg13g2_fill_1 FILLER_52_526 ();
 sg13g2_decap_4 FILLER_52_535 ();
 sg13g2_decap_8 FILLER_52_566 ();
 sg13g2_fill_1 FILLER_52_573 ();
 sg13g2_fill_2 FILLER_52_590 ();
 sg13g2_fill_1 FILLER_52_592 ();
 sg13g2_fill_2 FILLER_52_599 ();
 sg13g2_fill_1 FILLER_52_607 ();
 sg13g2_fill_2 FILLER_52_612 ();
 sg13g2_fill_2 FILLER_52_624 ();
 sg13g2_fill_1 FILLER_52_626 ();
 sg13g2_fill_1 FILLER_52_640 ();
 sg13g2_fill_2 FILLER_52_646 ();
 sg13g2_fill_1 FILLER_52_658 ();
 sg13g2_decap_4 FILLER_52_664 ();
 sg13g2_decap_8 FILLER_52_745 ();
 sg13g2_decap_8 FILLER_52_752 ();
 sg13g2_decap_8 FILLER_52_759 ();
 sg13g2_decap_8 FILLER_52_766 ();
 sg13g2_decap_8 FILLER_52_773 ();
 sg13g2_decap_8 FILLER_52_780 ();
 sg13g2_decap_8 FILLER_52_787 ();
 sg13g2_decap_8 FILLER_52_794 ();
 sg13g2_decap_8 FILLER_52_801 ();
 sg13g2_decap_8 FILLER_52_808 ();
 sg13g2_decap_8 FILLER_52_815 ();
 sg13g2_decap_8 FILLER_52_822 ();
 sg13g2_decap_8 FILLER_52_829 ();
 sg13g2_decap_8 FILLER_52_836 ();
 sg13g2_decap_8 FILLER_52_843 ();
 sg13g2_decap_8 FILLER_52_850 ();
 sg13g2_decap_4 FILLER_52_857 ();
 sg13g2_fill_1 FILLER_52_861 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_7 ();
 sg13g2_fill_2 FILLER_53_17 ();
 sg13g2_fill_1 FILLER_53_19 ();
 sg13g2_decap_4 FILLER_53_24 ();
 sg13g2_fill_2 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_34 ();
 sg13g2_decap_4 FILLER_53_41 ();
 sg13g2_fill_2 FILLER_53_45 ();
 sg13g2_decap_4 FILLER_53_51 ();
 sg13g2_fill_2 FILLER_53_55 ();
 sg13g2_fill_2 FILLER_53_79 ();
 sg13g2_fill_1 FILLER_53_81 ();
 sg13g2_fill_2 FILLER_53_96 ();
 sg13g2_fill_1 FILLER_53_98 ();
 sg13g2_decap_4 FILLER_53_103 ();
 sg13g2_fill_1 FILLER_53_107 ();
 sg13g2_fill_2 FILLER_53_132 ();
 sg13g2_fill_1 FILLER_53_134 ();
 sg13g2_fill_1 FILLER_53_165 ();
 sg13g2_decap_8 FILLER_53_170 ();
 sg13g2_decap_8 FILLER_53_177 ();
 sg13g2_fill_1 FILLER_53_184 ();
 sg13g2_fill_1 FILLER_53_189 ();
 sg13g2_fill_2 FILLER_53_257 ();
 sg13g2_fill_1 FILLER_53_259 ();
 sg13g2_fill_2 FILLER_53_271 ();
 sg13g2_fill_1 FILLER_53_273 ();
 sg13g2_fill_1 FILLER_53_280 ();
 sg13g2_decap_8 FILLER_53_323 ();
 sg13g2_decap_8 FILLER_53_330 ();
 sg13g2_decap_4 FILLER_53_337 ();
 sg13g2_fill_1 FILLER_53_341 ();
 sg13g2_decap_4 FILLER_53_360 ();
 sg13g2_fill_2 FILLER_53_369 ();
 sg13g2_fill_1 FILLER_53_371 ();
 sg13g2_decap_4 FILLER_53_377 ();
 sg13g2_decap_8 FILLER_53_386 ();
 sg13g2_fill_2 FILLER_53_393 ();
 sg13g2_decap_8 FILLER_53_399 ();
 sg13g2_decap_8 FILLER_53_406 ();
 sg13g2_fill_2 FILLER_53_413 ();
 sg13g2_fill_1 FILLER_53_415 ();
 sg13g2_decap_8 FILLER_53_424 ();
 sg13g2_decap_8 FILLER_53_431 ();
 sg13g2_decap_4 FILLER_53_438 ();
 sg13g2_fill_1 FILLER_53_442 ();
 sg13g2_fill_2 FILLER_53_460 ();
 sg13g2_fill_1 FILLER_53_462 ();
 sg13g2_decap_8 FILLER_53_482 ();
 sg13g2_decap_4 FILLER_53_489 ();
 sg13g2_fill_1 FILLER_53_493 ();
 sg13g2_decap_8 FILLER_53_498 ();
 sg13g2_fill_2 FILLER_53_505 ();
 sg13g2_decap_8 FILLER_53_532 ();
 sg13g2_fill_1 FILLER_53_539 ();
 sg13g2_fill_1 FILLER_53_564 ();
 sg13g2_fill_1 FILLER_53_576 ();
 sg13g2_fill_2 FILLER_53_595 ();
 sg13g2_fill_1 FILLER_53_597 ();
 sg13g2_fill_1 FILLER_53_651 ();
 sg13g2_fill_2 FILLER_53_704 ();
 sg13g2_fill_2 FILLER_53_721 ();
 sg13g2_decap_8 FILLER_53_745 ();
 sg13g2_decap_8 FILLER_53_752 ();
 sg13g2_decap_8 FILLER_53_759 ();
 sg13g2_decap_8 FILLER_53_766 ();
 sg13g2_decap_8 FILLER_53_773 ();
 sg13g2_decap_8 FILLER_53_780 ();
 sg13g2_decap_8 FILLER_53_787 ();
 sg13g2_decap_8 FILLER_53_794 ();
 sg13g2_decap_8 FILLER_53_801 ();
 sg13g2_decap_8 FILLER_53_808 ();
 sg13g2_decap_8 FILLER_53_815 ();
 sg13g2_decap_8 FILLER_53_822 ();
 sg13g2_decap_8 FILLER_53_829 ();
 sg13g2_decap_8 FILLER_53_836 ();
 sg13g2_decap_8 FILLER_53_843 ();
 sg13g2_decap_8 FILLER_53_850 ();
 sg13g2_decap_4 FILLER_53_857 ();
 sg13g2_fill_1 FILLER_53_861 ();
 sg13g2_fill_1 FILLER_54_0 ();
 sg13g2_decap_4 FILLER_54_53 ();
 sg13g2_fill_2 FILLER_54_57 ();
 sg13g2_fill_2 FILLER_54_68 ();
 sg13g2_fill_1 FILLER_54_70 ();
 sg13g2_fill_2 FILLER_54_81 ();
 sg13g2_fill_1 FILLER_54_83 ();
 sg13g2_decap_8 FILLER_54_88 ();
 sg13g2_fill_2 FILLER_54_95 ();
 sg13g2_fill_1 FILLER_54_106 ();
 sg13g2_decap_8 FILLER_54_121 ();
 sg13g2_decap_4 FILLER_54_132 ();
 sg13g2_fill_2 FILLER_54_144 ();
 sg13g2_fill_2 FILLER_54_160 ();
 sg13g2_fill_1 FILLER_54_172 ();
 sg13g2_decap_4 FILLER_54_199 ();
 sg13g2_decap_8 FILLER_54_221 ();
 sg13g2_decap_8 FILLER_54_228 ();
 sg13g2_decap_4 FILLER_54_235 ();
 sg13g2_fill_1 FILLER_54_239 ();
 sg13g2_fill_1 FILLER_54_244 ();
 sg13g2_decap_4 FILLER_54_254 ();
 sg13g2_decap_8 FILLER_54_263 ();
 sg13g2_decap_4 FILLER_54_270 ();
 sg13g2_fill_1 FILLER_54_279 ();
 sg13g2_decap_4 FILLER_54_286 ();
 sg13g2_fill_2 FILLER_54_290 ();
 sg13g2_fill_1 FILLER_54_303 ();
 sg13g2_decap_8 FILLER_54_315 ();
 sg13g2_decap_4 FILLER_54_322 ();
 sg13g2_fill_1 FILLER_54_326 ();
 sg13g2_decap_8 FILLER_54_339 ();
 sg13g2_fill_2 FILLER_54_346 ();
 sg13g2_decap_8 FILLER_54_360 ();
 sg13g2_fill_2 FILLER_54_367 ();
 sg13g2_fill_2 FILLER_54_381 ();
 sg13g2_decap_8 FILLER_54_389 ();
 sg13g2_decap_4 FILLER_54_425 ();
 sg13g2_fill_1 FILLER_54_429 ();
 sg13g2_fill_2 FILLER_54_441 ();
 sg13g2_fill_1 FILLER_54_449 ();
 sg13g2_decap_8 FILLER_54_456 ();
 sg13g2_decap_4 FILLER_54_463 ();
 sg13g2_decap_8 FILLER_54_475 ();
 sg13g2_decap_4 FILLER_54_482 ();
 sg13g2_fill_2 FILLER_54_486 ();
 sg13g2_decap_4 FILLER_54_507 ();
 sg13g2_fill_1 FILLER_54_511 ();
 sg13g2_decap_8 FILLER_54_537 ();
 sg13g2_decap_4 FILLER_54_544 ();
 sg13g2_fill_1 FILLER_54_548 ();
 sg13g2_decap_8 FILLER_54_558 ();
 sg13g2_decap_8 FILLER_54_565 ();
 sg13g2_fill_1 FILLER_54_572 ();
 sg13g2_fill_2 FILLER_54_595 ();
 sg13g2_fill_1 FILLER_54_597 ();
 sg13g2_decap_8 FILLER_54_618 ();
 sg13g2_fill_1 FILLER_54_625 ();
 sg13g2_fill_2 FILLER_54_638 ();
 sg13g2_fill_1 FILLER_54_640 ();
 sg13g2_fill_1 FILLER_54_651 ();
 sg13g2_decap_8 FILLER_54_678 ();
 sg13g2_fill_2 FILLER_54_685 ();
 sg13g2_fill_2 FILLER_54_692 ();
 sg13g2_fill_1 FILLER_54_694 ();
 sg13g2_fill_1 FILLER_54_705 ();
 sg13g2_decap_8 FILLER_54_758 ();
 sg13g2_decap_8 FILLER_54_765 ();
 sg13g2_decap_8 FILLER_54_772 ();
 sg13g2_decap_8 FILLER_54_779 ();
 sg13g2_decap_8 FILLER_54_786 ();
 sg13g2_decap_8 FILLER_54_793 ();
 sg13g2_decap_8 FILLER_54_800 ();
 sg13g2_decap_8 FILLER_54_807 ();
 sg13g2_decap_8 FILLER_54_814 ();
 sg13g2_decap_8 FILLER_54_821 ();
 sg13g2_decap_8 FILLER_54_828 ();
 sg13g2_decap_8 FILLER_54_835 ();
 sg13g2_decap_8 FILLER_54_842 ();
 sg13g2_decap_8 FILLER_54_849 ();
 sg13g2_decap_4 FILLER_54_856 ();
 sg13g2_fill_2 FILLER_54_860 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_4 FILLER_55_7 ();
 sg13g2_fill_2 FILLER_55_11 ();
 sg13g2_decap_8 FILLER_55_25 ();
 sg13g2_decap_4 FILLER_55_32 ();
 sg13g2_fill_1 FILLER_55_36 ();
 sg13g2_decap_8 FILLER_55_41 ();
 sg13g2_fill_2 FILLER_55_48 ();
 sg13g2_fill_1 FILLER_55_50 ();
 sg13g2_fill_2 FILLER_55_92 ();
 sg13g2_fill_1 FILLER_55_94 ();
 sg13g2_fill_2 FILLER_55_126 ();
 sg13g2_fill_1 FILLER_55_128 ();
 sg13g2_decap_4 FILLER_55_155 ();
 sg13g2_fill_2 FILLER_55_159 ();
 sg13g2_fill_1 FILLER_55_170 ();
 sg13g2_fill_2 FILLER_55_175 ();
 sg13g2_fill_2 FILLER_55_182 ();
 sg13g2_fill_1 FILLER_55_192 ();
 sg13g2_decap_8 FILLER_55_223 ();
 sg13g2_decap_4 FILLER_55_230 ();
 sg13g2_fill_2 FILLER_55_234 ();
 sg13g2_decap_8 FILLER_55_261 ();
 sg13g2_fill_1 FILLER_55_268 ();
 sg13g2_decap_4 FILLER_55_320 ();
 sg13g2_fill_1 FILLER_55_330 ();
 sg13g2_fill_2 FILLER_55_343 ();
 sg13g2_fill_1 FILLER_55_345 ();
 sg13g2_decap_4 FILLER_55_400 ();
 sg13g2_decap_4 FILLER_55_410 ();
 sg13g2_fill_2 FILLER_55_426 ();
 sg13g2_fill_1 FILLER_55_428 ();
 sg13g2_fill_2 FILLER_55_447 ();
 sg13g2_fill_2 FILLER_55_473 ();
 sg13g2_decap_4 FILLER_55_481 ();
 sg13g2_fill_1 FILLER_55_485 ();
 sg13g2_decap_8 FILLER_55_510 ();
 sg13g2_fill_2 FILLER_55_517 ();
 sg13g2_fill_1 FILLER_55_519 ();
 sg13g2_fill_2 FILLER_55_542 ();
 sg13g2_fill_1 FILLER_55_560 ();
 sg13g2_decap_8 FILLER_55_574 ();
 sg13g2_decap_4 FILLER_55_599 ();
 sg13g2_fill_2 FILLER_55_609 ();
 sg13g2_decap_8 FILLER_55_615 ();
 sg13g2_decap_4 FILLER_55_622 ();
 sg13g2_fill_1 FILLER_55_691 ();
 sg13g2_fill_1 FILLER_55_725 ();
 sg13g2_decap_8 FILLER_55_756 ();
 sg13g2_decap_8 FILLER_55_763 ();
 sg13g2_decap_8 FILLER_55_770 ();
 sg13g2_decap_8 FILLER_55_777 ();
 sg13g2_decap_8 FILLER_55_784 ();
 sg13g2_decap_8 FILLER_55_791 ();
 sg13g2_decap_8 FILLER_55_798 ();
 sg13g2_decap_8 FILLER_55_805 ();
 sg13g2_decap_8 FILLER_55_812 ();
 sg13g2_decap_8 FILLER_55_819 ();
 sg13g2_decap_8 FILLER_55_826 ();
 sg13g2_decap_8 FILLER_55_833 ();
 sg13g2_decap_8 FILLER_55_840 ();
 sg13g2_decap_8 FILLER_55_847 ();
 sg13g2_decap_8 FILLER_55_854 ();
 sg13g2_fill_1 FILLER_55_861 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_33 ();
 sg13g2_fill_1 FILLER_56_60 ();
 sg13g2_fill_2 FILLER_56_70 ();
 sg13g2_fill_1 FILLER_56_72 ();
 sg13g2_fill_1 FILLER_56_104 ();
 sg13g2_decap_4 FILLER_56_109 ();
 sg13g2_fill_1 FILLER_56_113 ();
 sg13g2_fill_1 FILLER_56_128 ();
 sg13g2_fill_2 FILLER_56_161 ();
 sg13g2_decap_4 FILLER_56_171 ();
 sg13g2_fill_2 FILLER_56_175 ();
 sg13g2_fill_1 FILLER_56_187 ();
 sg13g2_fill_1 FILLER_56_192 ();
 sg13g2_decap_8 FILLER_56_232 ();
 sg13g2_fill_1 FILLER_56_265 ();
 sg13g2_decap_8 FILLER_56_287 ();
 sg13g2_fill_1 FILLER_56_294 ();
 sg13g2_fill_2 FILLER_56_302 ();
 sg13g2_fill_1 FILLER_56_304 ();
 sg13g2_decap_8 FILLER_56_316 ();
 sg13g2_decap_8 FILLER_56_323 ();
 sg13g2_fill_2 FILLER_56_330 ();
 sg13g2_decap_4 FILLER_56_350 ();
 sg13g2_fill_1 FILLER_56_354 ();
 sg13g2_decap_8 FILLER_56_391 ();
 sg13g2_decap_4 FILLER_56_398 ();
 sg13g2_fill_2 FILLER_56_402 ();
 sg13g2_fill_1 FILLER_56_432 ();
 sg13g2_decap_4 FILLER_56_439 ();
 sg13g2_fill_1 FILLER_56_443 ();
 sg13g2_fill_2 FILLER_56_478 ();
 sg13g2_fill_1 FILLER_56_480 ();
 sg13g2_decap_8 FILLER_56_487 ();
 sg13g2_fill_2 FILLER_56_494 ();
 sg13g2_decap_4 FILLER_56_500 ();
 sg13g2_fill_1 FILLER_56_504 ();
 sg13g2_fill_2 FILLER_56_562 ();
 sg13g2_fill_1 FILLER_56_564 ();
 sg13g2_fill_2 FILLER_56_593 ();
 sg13g2_fill_1 FILLER_56_595 ();
 sg13g2_decap_4 FILLER_56_626 ();
 sg13g2_fill_1 FILLER_56_630 ();
 sg13g2_fill_1 FILLER_56_636 ();
 sg13g2_fill_2 FILLER_56_656 ();
 sg13g2_fill_1 FILLER_56_684 ();
 sg13g2_fill_2 FILLER_56_689 ();
 sg13g2_fill_1 FILLER_56_691 ();
 sg13g2_fill_2 FILLER_56_706 ();
 sg13g2_decap_8 FILLER_56_760 ();
 sg13g2_decap_8 FILLER_56_767 ();
 sg13g2_decap_8 FILLER_56_774 ();
 sg13g2_decap_8 FILLER_56_781 ();
 sg13g2_decap_8 FILLER_56_788 ();
 sg13g2_decap_8 FILLER_56_795 ();
 sg13g2_decap_8 FILLER_56_802 ();
 sg13g2_decap_8 FILLER_56_809 ();
 sg13g2_decap_8 FILLER_56_816 ();
 sg13g2_decap_8 FILLER_56_823 ();
 sg13g2_decap_8 FILLER_56_830 ();
 sg13g2_decap_8 FILLER_56_837 ();
 sg13g2_decap_8 FILLER_56_844 ();
 sg13g2_decap_8 FILLER_56_851 ();
 sg13g2_decap_4 FILLER_56_858 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_2 ();
 sg13g2_fill_1 FILLER_57_29 ();
 sg13g2_fill_2 FILLER_57_35 ();
 sg13g2_fill_1 FILLER_57_37 ();
 sg13g2_fill_2 FILLER_57_42 ();
 sg13g2_fill_1 FILLER_57_44 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_4 FILLER_57_56 ();
 sg13g2_fill_2 FILLER_57_60 ();
 sg13g2_decap_4 FILLER_57_75 ();
 sg13g2_fill_2 FILLER_57_96 ();
 sg13g2_fill_1 FILLER_57_98 ();
 sg13g2_fill_2 FILLER_57_103 ();
 sg13g2_fill_1 FILLER_57_105 ();
 sg13g2_decap_8 FILLER_57_140 ();
 sg13g2_decap_8 FILLER_57_147 ();
 sg13g2_fill_2 FILLER_57_215 ();
 sg13g2_decap_8 FILLER_57_221 ();
 sg13g2_decap_4 FILLER_57_228 ();
 sg13g2_fill_2 FILLER_57_245 ();
 sg13g2_fill_1 FILLER_57_252 ();
 sg13g2_decap_4 FILLER_57_261 ();
 sg13g2_fill_1 FILLER_57_265 ();
 sg13g2_decap_4 FILLER_57_271 ();
 sg13g2_fill_2 FILLER_57_275 ();
 sg13g2_fill_2 FILLER_57_283 ();
 sg13g2_decap_8 FILLER_57_290 ();
 sg13g2_fill_1 FILLER_57_315 ();
 sg13g2_decap_4 FILLER_57_322 ();
 sg13g2_fill_2 FILLER_57_326 ();
 sg13g2_fill_2 FILLER_57_346 ();
 sg13g2_fill_2 FILLER_57_354 ();
 sg13g2_fill_1 FILLER_57_356 ();
 sg13g2_decap_4 FILLER_57_363 ();
 sg13g2_fill_1 FILLER_57_367 ();
 sg13g2_fill_2 FILLER_57_438 ();
 sg13g2_fill_1 FILLER_57_440 ();
 sg13g2_decap_4 FILLER_57_451 ();
 sg13g2_fill_1 FILLER_57_455 ();
 sg13g2_decap_4 FILLER_57_480 ();
 sg13g2_fill_1 FILLER_57_484 ();
 sg13g2_fill_1 FILLER_57_493 ();
 sg13g2_fill_2 FILLER_57_509 ();
 sg13g2_fill_1 FILLER_57_511 ();
 sg13g2_decap_4 FILLER_57_521 ();
 sg13g2_fill_1 FILLER_57_525 ();
 sg13g2_decap_8 FILLER_57_541 ();
 sg13g2_fill_2 FILLER_57_548 ();
 sg13g2_fill_1 FILLER_57_562 ();
 sg13g2_fill_2 FILLER_57_599 ();
 sg13g2_fill_2 FILLER_57_606 ();
 sg13g2_fill_1 FILLER_57_608 ();
 sg13g2_decap_8 FILLER_57_614 ();
 sg13g2_fill_2 FILLER_57_621 ();
 sg13g2_fill_2 FILLER_57_628 ();
 sg13g2_fill_1 FILLER_57_630 ();
 sg13g2_fill_1 FILLER_57_640 ();
 sg13g2_fill_1 FILLER_57_655 ();
 sg13g2_decap_4 FILLER_57_661 ();
 sg13g2_fill_1 FILLER_57_670 ();
 sg13g2_fill_2 FILLER_57_735 ();
 sg13g2_decap_8 FILLER_57_763 ();
 sg13g2_decap_8 FILLER_57_770 ();
 sg13g2_decap_8 FILLER_57_777 ();
 sg13g2_decap_8 FILLER_57_784 ();
 sg13g2_decap_8 FILLER_57_791 ();
 sg13g2_decap_8 FILLER_57_798 ();
 sg13g2_decap_8 FILLER_57_805 ();
 sg13g2_decap_8 FILLER_57_812 ();
 sg13g2_decap_8 FILLER_57_819 ();
 sg13g2_decap_8 FILLER_57_826 ();
 sg13g2_decap_8 FILLER_57_833 ();
 sg13g2_decap_8 FILLER_57_840 ();
 sg13g2_decap_8 FILLER_57_847 ();
 sg13g2_decap_8 FILLER_57_854 ();
 sg13g2_fill_1 FILLER_57_861 ();
 sg13g2_fill_1 FILLER_58_26 ();
 sg13g2_fill_2 FILLER_58_57 ();
 sg13g2_fill_1 FILLER_58_78 ();
 sg13g2_decap_8 FILLER_58_109 ();
 sg13g2_decap_4 FILLER_58_116 ();
 sg13g2_fill_2 FILLER_58_120 ();
 sg13g2_decap_4 FILLER_58_130 ();
 sg13g2_fill_2 FILLER_58_134 ();
 sg13g2_fill_1 FILLER_58_140 ();
 sg13g2_fill_1 FILLER_58_151 ();
 sg13g2_fill_1 FILLER_58_170 ();
 sg13g2_decap_8 FILLER_58_189 ();
 sg13g2_decap_4 FILLER_58_196 ();
 sg13g2_fill_2 FILLER_58_204 ();
 sg13g2_fill_1 FILLER_58_206 ();
 sg13g2_fill_2 FILLER_58_227 ();
 sg13g2_fill_1 FILLER_58_229 ();
 sg13g2_decap_8 FILLER_58_294 ();
 sg13g2_decap_4 FILLER_58_318 ();
 sg13g2_decap_8 FILLER_58_346 ();
 sg13g2_fill_1 FILLER_58_353 ();
 sg13g2_decap_8 FILLER_58_361 ();
 sg13g2_fill_1 FILLER_58_368 ();
 sg13g2_fill_2 FILLER_58_375 ();
 sg13g2_decap_8 FILLER_58_396 ();
 sg13g2_fill_1 FILLER_58_403 ();
 sg13g2_decap_8 FILLER_58_435 ();
 sg13g2_decap_8 FILLER_58_442 ();
 sg13g2_fill_2 FILLER_58_449 ();
 sg13g2_fill_1 FILLER_58_457 ();
 sg13g2_decap_8 FILLER_58_476 ();
 sg13g2_fill_1 FILLER_58_483 ();
 sg13g2_decap_4 FILLER_58_504 ();
 sg13g2_fill_2 FILLER_58_517 ();
 sg13g2_fill_1 FILLER_58_519 ();
 sg13g2_decap_4 FILLER_58_525 ();
 sg13g2_decap_8 FILLER_58_546 ();
 sg13g2_fill_1 FILLER_58_560 ();
 sg13g2_decap_8 FILLER_58_569 ();
 sg13g2_fill_2 FILLER_58_576 ();
 sg13g2_decap_4 FILLER_58_582 ();
 sg13g2_fill_2 FILLER_58_601 ();
 sg13g2_fill_1 FILLER_58_603 ();
 sg13g2_fill_2 FILLER_58_608 ();
 sg13g2_fill_2 FILLER_58_623 ();
 sg13g2_fill_1 FILLER_58_625 ();
 sg13g2_fill_2 FILLER_58_642 ();
 sg13g2_decap_4 FILLER_58_655 ();
 sg13g2_fill_2 FILLER_58_690 ();
 sg13g2_fill_1 FILLER_58_697 ();
 sg13g2_fill_1 FILLER_58_703 ();
 sg13g2_fill_2 FILLER_58_709 ();
 sg13g2_fill_2 FILLER_58_746 ();
 sg13g2_decap_8 FILLER_58_756 ();
 sg13g2_decap_8 FILLER_58_763 ();
 sg13g2_decap_8 FILLER_58_770 ();
 sg13g2_decap_8 FILLER_58_777 ();
 sg13g2_decap_8 FILLER_58_784 ();
 sg13g2_decap_8 FILLER_58_791 ();
 sg13g2_decap_8 FILLER_58_798 ();
 sg13g2_decap_8 FILLER_58_805 ();
 sg13g2_decap_8 FILLER_58_812 ();
 sg13g2_decap_8 FILLER_58_819 ();
 sg13g2_decap_8 FILLER_58_826 ();
 sg13g2_decap_8 FILLER_58_833 ();
 sg13g2_decap_8 FILLER_58_840 ();
 sg13g2_decap_8 FILLER_58_847 ();
 sg13g2_decap_8 FILLER_58_854 ();
 sg13g2_fill_1 FILLER_58_861 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_fill_2 FILLER_59_7 ();
 sg13g2_fill_1 FILLER_59_13 ();
 sg13g2_fill_1 FILLER_59_18 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_4 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_4 FILLER_59_84 ();
 sg13g2_fill_2 FILLER_59_88 ();
 sg13g2_decap_4 FILLER_59_108 ();
 sg13g2_decap_8 FILLER_59_116 ();
 sg13g2_decap_8 FILLER_59_123 ();
 sg13g2_decap_8 FILLER_59_156 ();
 sg13g2_fill_1 FILLER_59_163 ();
 sg13g2_decap_8 FILLER_59_172 ();
 sg13g2_fill_1 FILLER_59_179 ();
 sg13g2_fill_1 FILLER_59_193 ();
 sg13g2_decap_8 FILLER_59_202 ();
 sg13g2_fill_2 FILLER_59_209 ();
 sg13g2_fill_2 FILLER_59_215 ();
 sg13g2_decap_8 FILLER_59_222 ();
 sg13g2_decap_8 FILLER_59_229 ();
 sg13g2_decap_4 FILLER_59_236 ();
 sg13g2_fill_1 FILLER_59_259 ();
 sg13g2_decap_8 FILLER_59_265 ();
 sg13g2_decap_4 FILLER_59_272 ();
 sg13g2_fill_1 FILLER_59_276 ();
 sg13g2_decap_8 FILLER_59_285 ();
 sg13g2_fill_1 FILLER_59_292 ();
 sg13g2_fill_2 FILLER_59_302 ();
 sg13g2_fill_2 FILLER_59_328 ();
 sg13g2_fill_2 FILLER_59_336 ();
 sg13g2_decap_4 FILLER_59_362 ();
 sg13g2_decap_8 FILLER_59_384 ();
 sg13g2_decap_4 FILLER_59_391 ();
 sg13g2_fill_2 FILLER_59_401 ();
 sg13g2_fill_2 FILLER_59_434 ();
 sg13g2_decap_8 FILLER_59_440 ();
 sg13g2_decap_4 FILLER_59_453 ();
 sg13g2_fill_1 FILLER_59_457 ();
 sg13g2_decap_8 FILLER_59_476 ();
 sg13g2_decap_8 FILLER_59_483 ();
 sg13g2_decap_8 FILLER_59_490 ();
 sg13g2_decap_4 FILLER_59_497 ();
 sg13g2_fill_2 FILLER_59_501 ();
 sg13g2_fill_2 FILLER_59_520 ();
 sg13g2_fill_1 FILLER_59_522 ();
 sg13g2_fill_2 FILLER_59_528 ();
 sg13g2_fill_1 FILLER_59_530 ();
 sg13g2_decap_8 FILLER_59_543 ();
 sg13g2_decap_4 FILLER_59_550 ();
 sg13g2_fill_2 FILLER_59_565 ();
 sg13g2_fill_1 FILLER_59_567 ();
 sg13g2_fill_2 FILLER_59_577 ();
 sg13g2_fill_1 FILLER_59_579 ();
 sg13g2_decap_8 FILLER_59_591 ();
 sg13g2_fill_2 FILLER_59_618 ();
 sg13g2_decap_4 FILLER_59_629 ();
 sg13g2_fill_1 FILLER_59_633 ();
 sg13g2_decap_4 FILLER_59_651 ();
 sg13g2_fill_1 FILLER_59_655 ();
 sg13g2_fill_2 FILLER_59_661 ();
 sg13g2_fill_1 FILLER_59_663 ();
 sg13g2_fill_1 FILLER_59_692 ();
 sg13g2_fill_2 FILLER_59_708 ();
 sg13g2_fill_2 FILLER_59_734 ();
 sg13g2_fill_1 FILLER_59_736 ();
 sg13g2_decap_8 FILLER_59_763 ();
 sg13g2_decap_8 FILLER_59_770 ();
 sg13g2_decap_8 FILLER_59_777 ();
 sg13g2_decap_8 FILLER_59_784 ();
 sg13g2_decap_8 FILLER_59_791 ();
 sg13g2_decap_8 FILLER_59_798 ();
 sg13g2_decap_8 FILLER_59_805 ();
 sg13g2_decap_8 FILLER_59_812 ();
 sg13g2_decap_8 FILLER_59_819 ();
 sg13g2_decap_8 FILLER_59_826 ();
 sg13g2_decap_8 FILLER_59_833 ();
 sg13g2_decap_8 FILLER_59_840 ();
 sg13g2_decap_8 FILLER_59_847 ();
 sg13g2_decap_8 FILLER_59_854 ();
 sg13g2_fill_1 FILLER_59_861 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_7 ();
 sg13g2_fill_1 FILLER_60_9 ();
 sg13g2_fill_2 FILLER_60_52 ();
 sg13g2_fill_1 FILLER_60_74 ();
 sg13g2_fill_2 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_122 ();
 sg13g2_fill_1 FILLER_60_129 ();
 sg13g2_decap_4 FILLER_60_148 ();
 sg13g2_fill_2 FILLER_60_157 ();
 sg13g2_fill_1 FILLER_60_159 ();
 sg13g2_fill_2 FILLER_60_180 ();
 sg13g2_decap_4 FILLER_60_213 ();
 sg13g2_decap_8 FILLER_60_234 ();
 sg13g2_fill_2 FILLER_60_241 ();
 sg13g2_fill_2 FILLER_60_256 ();
 sg13g2_fill_1 FILLER_60_287 ();
 sg13g2_fill_2 FILLER_60_330 ();
 sg13g2_decap_4 FILLER_60_338 ();
 sg13g2_fill_1 FILLER_60_361 ();
 sg13g2_fill_2 FILLER_60_391 ();
 sg13g2_fill_1 FILLER_60_393 ();
 sg13g2_fill_2 FILLER_60_406 ();
 sg13g2_fill_1 FILLER_60_444 ();
 sg13g2_decap_4 FILLER_60_487 ();
 sg13g2_fill_1 FILLER_60_504 ();
 sg13g2_fill_2 FILLER_60_520 ();
 sg13g2_fill_1 FILLER_60_527 ();
 sg13g2_fill_2 FILLER_60_533 ();
 sg13g2_decap_4 FILLER_60_543 ();
 sg13g2_fill_1 FILLER_60_547 ();
 sg13g2_fill_1 FILLER_60_551 ();
 sg13g2_fill_2 FILLER_60_575 ();
 sg13g2_decap_8 FILLER_60_585 ();
 sg13g2_decap_8 FILLER_60_592 ();
 sg13g2_fill_2 FILLER_60_599 ();
 sg13g2_fill_2 FILLER_60_617 ();
 sg13g2_decap_8 FILLER_60_637 ();
 sg13g2_fill_2 FILLER_60_729 ();
 sg13g2_fill_1 FILLER_60_731 ();
 sg13g2_fill_2 FILLER_60_737 ();
 sg13g2_fill_1 FILLER_60_739 ();
 sg13g2_decap_8 FILLER_60_775 ();
 sg13g2_decap_8 FILLER_60_782 ();
 sg13g2_decap_8 FILLER_60_789 ();
 sg13g2_decap_8 FILLER_60_796 ();
 sg13g2_decap_8 FILLER_60_803 ();
 sg13g2_decap_8 FILLER_60_810 ();
 sg13g2_decap_8 FILLER_60_817 ();
 sg13g2_decap_8 FILLER_60_824 ();
 sg13g2_decap_8 FILLER_60_831 ();
 sg13g2_decap_8 FILLER_60_838 ();
 sg13g2_decap_8 FILLER_60_845 ();
 sg13g2_decap_8 FILLER_60_852 ();
 sg13g2_fill_2 FILLER_60_859 ();
 sg13g2_fill_1 FILLER_60_861 ();
 sg13g2_decap_4 FILLER_61_26 ();
 sg13g2_fill_2 FILLER_61_64 ();
 sg13g2_decap_8 FILLER_61_75 ();
 sg13g2_fill_2 FILLER_61_82 ();
 sg13g2_fill_1 FILLER_61_88 ();
 sg13g2_fill_1 FILLER_61_94 ();
 sg13g2_decap_4 FILLER_61_99 ();
 sg13g2_fill_1 FILLER_61_103 ();
 sg13g2_fill_2 FILLER_61_108 ();
 sg13g2_fill_2 FILLER_61_119 ();
 sg13g2_fill_1 FILLER_61_121 ();
 sg13g2_decap_4 FILLER_61_126 ();
 sg13g2_fill_1 FILLER_61_130 ();
 sg13g2_fill_2 FILLER_61_141 ();
 sg13g2_decap_8 FILLER_61_173 ();
 sg13g2_fill_2 FILLER_61_180 ();
 sg13g2_fill_1 FILLER_61_182 ();
 sg13g2_decap_4 FILLER_61_197 ();
 sg13g2_fill_1 FILLER_61_201 ();
 sg13g2_fill_2 FILLER_61_212 ();
 sg13g2_decap_8 FILLER_61_227 ();
 sg13g2_fill_1 FILLER_61_234 ();
 sg13g2_fill_1 FILLER_61_243 ();
 sg13g2_fill_2 FILLER_61_266 ();
 sg13g2_fill_1 FILLER_61_268 ();
 sg13g2_fill_1 FILLER_61_278 ();
 sg13g2_fill_2 FILLER_61_284 ();
 sg13g2_fill_1 FILLER_61_286 ();
 sg13g2_fill_2 FILLER_61_293 ();
 sg13g2_fill_1 FILLER_61_295 ();
 sg13g2_decap_8 FILLER_61_308 ();
 sg13g2_fill_1 FILLER_61_315 ();
 sg13g2_fill_2 FILLER_61_322 ();
 sg13g2_fill_2 FILLER_61_333 ();
 sg13g2_fill_1 FILLER_61_335 ();
 sg13g2_decap_8 FILLER_61_343 ();
 sg13g2_fill_1 FILLER_61_350 ();
 sg13g2_fill_1 FILLER_61_357 ();
 sg13g2_decap_4 FILLER_61_364 ();
 sg13g2_fill_1 FILLER_61_368 ();
 sg13g2_decap_4 FILLER_61_375 ();
 sg13g2_fill_2 FILLER_61_379 ();
 sg13g2_decap_8 FILLER_61_387 ();
 sg13g2_fill_1 FILLER_61_394 ();
 sg13g2_decap_4 FILLER_61_401 ();
 sg13g2_fill_2 FILLER_61_411 ();
 sg13g2_decap_8 FILLER_61_436 ();
 sg13g2_decap_8 FILLER_61_443 ();
 sg13g2_decap_4 FILLER_61_480 ();
 sg13g2_fill_1 FILLER_61_484 ();
 sg13g2_fill_1 FILLER_61_506 ();
 sg13g2_decap_4 FILLER_61_512 ();
 sg13g2_fill_2 FILLER_61_516 ();
 sg13g2_decap_4 FILLER_61_546 ();
 sg13g2_fill_2 FILLER_61_550 ();
 sg13g2_fill_2 FILLER_61_567 ();
 sg13g2_fill_1 FILLER_61_588 ();
 sg13g2_decap_8 FILLER_61_599 ();
 sg13g2_fill_1 FILLER_61_616 ();
 sg13g2_decap_8 FILLER_61_636 ();
 sg13g2_decap_4 FILLER_61_643 ();
 sg13g2_fill_2 FILLER_61_647 ();
 sg13g2_fill_2 FILLER_61_657 ();
 sg13g2_fill_1 FILLER_61_659 ();
 sg13g2_fill_2 FILLER_61_664 ();
 sg13g2_fill_2 FILLER_61_697 ();
 sg13g2_fill_2 FILLER_61_725 ();
 sg13g2_decap_8 FILLER_61_766 ();
 sg13g2_decap_8 FILLER_61_773 ();
 sg13g2_decap_8 FILLER_61_780 ();
 sg13g2_decap_8 FILLER_61_787 ();
 sg13g2_decap_8 FILLER_61_794 ();
 sg13g2_decap_8 FILLER_61_801 ();
 sg13g2_decap_8 FILLER_61_808 ();
 sg13g2_decap_8 FILLER_61_815 ();
 sg13g2_decap_8 FILLER_61_822 ();
 sg13g2_decap_8 FILLER_61_829 ();
 sg13g2_decap_8 FILLER_61_836 ();
 sg13g2_decap_8 FILLER_61_843 ();
 sg13g2_decap_8 FILLER_61_850 ();
 sg13g2_decap_4 FILLER_61_857 ();
 sg13g2_fill_1 FILLER_61_861 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_4 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_15 ();
 sg13g2_decap_8 FILLER_62_22 ();
 sg13g2_decap_8 FILLER_62_38 ();
 sg13g2_decap_4 FILLER_62_45 ();
 sg13g2_decap_4 FILLER_62_53 ();
 sg13g2_fill_2 FILLER_62_57 ();
 sg13g2_fill_1 FILLER_62_80 ();
 sg13g2_decap_4 FILLER_62_107 ();
 sg13g2_decap_4 FILLER_62_150 ();
 sg13g2_fill_1 FILLER_62_154 ();
 sg13g2_fill_2 FILLER_62_163 ();
 sg13g2_fill_1 FILLER_62_191 ();
 sg13g2_decap_4 FILLER_62_252 ();
 sg13g2_fill_2 FILLER_62_256 ();
 sg13g2_fill_2 FILLER_62_263 ();
 sg13g2_fill_1 FILLER_62_265 ();
 sg13g2_decap_8 FILLER_62_275 ();
 sg13g2_fill_1 FILLER_62_282 ();
 sg13g2_fill_2 FILLER_62_299 ();
 sg13g2_fill_1 FILLER_62_301 ();
 sg13g2_fill_2 FILLER_62_323 ();
 sg13g2_fill_2 FILLER_62_331 ();
 sg13g2_decap_4 FILLER_62_345 ();
 sg13g2_decap_4 FILLER_62_382 ();
 sg13g2_fill_1 FILLER_62_386 ();
 sg13g2_fill_1 FILLER_62_405 ();
 sg13g2_decap_8 FILLER_62_410 ();
 sg13g2_decap_4 FILLER_62_417 ();
 sg13g2_fill_1 FILLER_62_421 ();
 sg13g2_decap_8 FILLER_62_427 ();
 sg13g2_decap_8 FILLER_62_440 ();
 sg13g2_fill_2 FILLER_62_447 ();
 sg13g2_decap_8 FILLER_62_476 ();
 sg13g2_fill_2 FILLER_62_514 ();
 sg13g2_fill_1 FILLER_62_516 ();
 sg13g2_decap_8 FILLER_62_547 ();
 sg13g2_fill_2 FILLER_62_554 ();
 sg13g2_fill_2 FILLER_62_566 ();
 sg13g2_fill_1 FILLER_62_568 ();
 sg13g2_fill_2 FILLER_62_582 ();
 sg13g2_fill_1 FILLER_62_584 ();
 sg13g2_fill_2 FILLER_62_599 ();
 sg13g2_fill_1 FILLER_62_606 ();
 sg13g2_fill_2 FILLER_62_613 ();
 sg13g2_fill_1 FILLER_62_615 ();
 sg13g2_decap_4 FILLER_62_637 ();
 sg13g2_decap_8 FILLER_62_645 ();
 sg13g2_fill_1 FILLER_62_652 ();
 sg13g2_fill_1 FILLER_62_661 ();
 sg13g2_decap_8 FILLER_62_667 ();
 sg13g2_fill_2 FILLER_62_674 ();
 sg13g2_decap_4 FILLER_62_689 ();
 sg13g2_fill_1 FILLER_62_693 ();
 sg13g2_fill_1 FILLER_62_708 ();
 sg13g2_fill_2 FILLER_62_721 ();
 sg13g2_fill_1 FILLER_62_723 ();
 sg13g2_decap_8 FILLER_62_756 ();
 sg13g2_decap_8 FILLER_62_763 ();
 sg13g2_decap_8 FILLER_62_770 ();
 sg13g2_decap_8 FILLER_62_777 ();
 sg13g2_decap_8 FILLER_62_784 ();
 sg13g2_decap_8 FILLER_62_791 ();
 sg13g2_decap_8 FILLER_62_798 ();
 sg13g2_decap_8 FILLER_62_805 ();
 sg13g2_decap_8 FILLER_62_812 ();
 sg13g2_decap_8 FILLER_62_819 ();
 sg13g2_decap_8 FILLER_62_826 ();
 sg13g2_decap_8 FILLER_62_833 ();
 sg13g2_decap_8 FILLER_62_840 ();
 sg13g2_decap_8 FILLER_62_847 ();
 sg13g2_decap_8 FILLER_62_854 ();
 sg13g2_fill_1 FILLER_62_861 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_4 FILLER_63_7 ();
 sg13g2_fill_1 FILLER_63_11 ();
 sg13g2_decap_8 FILLER_63_16 ();
 sg13g2_fill_1 FILLER_63_33 ();
 sg13g2_fill_1 FILLER_63_60 ();
 sg13g2_fill_2 FILLER_63_67 ();
 sg13g2_fill_1 FILLER_63_69 ();
 sg13g2_decap_4 FILLER_63_87 ();
 sg13g2_fill_2 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_102 ();
 sg13g2_decap_4 FILLER_63_109 ();
 sg13g2_decap_4 FILLER_63_117 ();
 sg13g2_fill_2 FILLER_63_121 ();
 sg13g2_decap_8 FILLER_63_138 ();
 sg13g2_decap_8 FILLER_63_145 ();
 sg13g2_decap_4 FILLER_63_152 ();
 sg13g2_decap_8 FILLER_63_161 ();
 sg13g2_decap_8 FILLER_63_168 ();
 sg13g2_fill_1 FILLER_63_175 ();
 sg13g2_decap_4 FILLER_63_180 ();
 sg13g2_fill_1 FILLER_63_184 ();
 sg13g2_decap_4 FILLER_63_200 ();
 sg13g2_decap_8 FILLER_63_209 ();
 sg13g2_decap_8 FILLER_63_216 ();
 sg13g2_fill_2 FILLER_63_223 ();
 sg13g2_decap_4 FILLER_63_233 ();
 sg13g2_fill_1 FILLER_63_237 ();
 sg13g2_decap_4 FILLER_63_243 ();
 sg13g2_fill_2 FILLER_63_247 ();
 sg13g2_decap_4 FILLER_63_286 ();
 sg13g2_fill_2 FILLER_63_290 ();
 sg13g2_decap_8 FILLER_63_303 ();
 sg13g2_decap_8 FILLER_63_310 ();
 sg13g2_decap_4 FILLER_63_317 ();
 sg13g2_fill_1 FILLER_63_321 ();
 sg13g2_fill_2 FILLER_63_343 ();
 sg13g2_fill_1 FILLER_63_345 ();
 sg13g2_fill_2 FILLER_63_352 ();
 sg13g2_decap_8 FILLER_63_360 ();
 sg13g2_decap_4 FILLER_63_367 ();
 sg13g2_fill_2 FILLER_63_371 ();
 sg13g2_fill_1 FILLER_63_379 ();
 sg13g2_decap_8 FILLER_63_387 ();
 sg13g2_decap_8 FILLER_63_400 ();
 sg13g2_decap_8 FILLER_63_407 ();
 sg13g2_decap_4 FILLER_63_437 ();
 sg13g2_fill_1 FILLER_63_441 ();
 sg13g2_fill_2 FILLER_63_458 ();
 sg13g2_fill_1 FILLER_63_460 ();
 sg13g2_decap_8 FILLER_63_481 ();
 sg13g2_decap_8 FILLER_63_488 ();
 sg13g2_decap_8 FILLER_63_499 ();
 sg13g2_fill_1 FILLER_63_506 ();
 sg13g2_fill_2 FILLER_63_513 ();
 sg13g2_fill_1 FILLER_63_515 ();
 sg13g2_decap_4 FILLER_63_542 ();
 sg13g2_fill_1 FILLER_63_546 ();
 sg13g2_fill_1 FILLER_63_566 ();
 sg13g2_decap_4 FILLER_63_577 ();
 sg13g2_fill_2 FILLER_63_581 ();
 sg13g2_fill_1 FILLER_63_589 ();
 sg13g2_fill_2 FILLER_63_603 ();
 sg13g2_decap_8 FILLER_63_615 ();
 sg13g2_fill_2 FILLER_63_622 ();
 sg13g2_fill_1 FILLER_63_624 ();
 sg13g2_fill_1 FILLER_63_661 ();
 sg13g2_fill_2 FILLER_63_723 ();
 sg13g2_fill_1 FILLER_63_725 ();
 sg13g2_fill_2 FILLER_63_731 ();
 sg13g2_fill_1 FILLER_63_733 ();
 sg13g2_fill_1 FILLER_63_739 ();
 sg13g2_decap_8 FILLER_63_766 ();
 sg13g2_decap_8 FILLER_63_773 ();
 sg13g2_decap_8 FILLER_63_780 ();
 sg13g2_decap_8 FILLER_63_787 ();
 sg13g2_decap_8 FILLER_63_794 ();
 sg13g2_decap_8 FILLER_63_801 ();
 sg13g2_decap_8 FILLER_63_808 ();
 sg13g2_decap_8 FILLER_63_815 ();
 sg13g2_decap_8 FILLER_63_822 ();
 sg13g2_decap_8 FILLER_63_829 ();
 sg13g2_decap_8 FILLER_63_836 ();
 sg13g2_decap_8 FILLER_63_843 ();
 sg13g2_decap_8 FILLER_63_850 ();
 sg13g2_decap_4 FILLER_63_857 ();
 sg13g2_fill_1 FILLER_63_861 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_33 ();
 sg13g2_fill_2 FILLER_64_43 ();
 sg13g2_decap_8 FILLER_64_53 ();
 sg13g2_fill_2 FILLER_64_60 ();
 sg13g2_fill_1 FILLER_64_62 ();
 sg13g2_fill_2 FILLER_64_74 ();
 sg13g2_fill_2 FILLER_64_81 ();
 sg13g2_fill_1 FILLER_64_83 ();
 sg13g2_fill_2 FILLER_64_100 ();
 sg13g2_fill_1 FILLER_64_133 ();
 sg13g2_fill_2 FILLER_64_231 ();
 sg13g2_fill_1 FILLER_64_233 ();
 sg13g2_fill_1 FILLER_64_242 ();
 sg13g2_decap_8 FILLER_64_267 ();
 sg13g2_decap_4 FILLER_64_274 ();
 sg13g2_fill_2 FILLER_64_301 ();
 sg13g2_decap_4 FILLER_64_341 ();
 sg13g2_fill_1 FILLER_64_345 ();
 sg13g2_fill_2 FILLER_64_389 ();
 sg13g2_fill_1 FILLER_64_391 ();
 sg13g2_fill_1 FILLER_64_398 ();
 sg13g2_decap_8 FILLER_64_403 ();
 sg13g2_fill_2 FILLER_64_410 ();
 sg13g2_fill_2 FILLER_64_436 ();
 sg13g2_fill_1 FILLER_64_438 ();
 sg13g2_decap_8 FILLER_64_444 ();
 sg13g2_fill_1 FILLER_64_451 ();
 sg13g2_fill_1 FILLER_64_506 ();
 sg13g2_decap_4 FILLER_64_512 ();
 sg13g2_fill_2 FILLER_64_516 ();
 sg13g2_decap_8 FILLER_64_522 ();
 sg13g2_decap_8 FILLER_64_534 ();
 sg13g2_fill_1 FILLER_64_541 ();
 sg13g2_decap_8 FILLER_64_560 ();
 sg13g2_decap_8 FILLER_64_567 ();
 sg13g2_decap_8 FILLER_64_620 ();
 sg13g2_fill_2 FILLER_64_627 ();
 sg13g2_fill_1 FILLER_64_629 ();
 sg13g2_decap_8 FILLER_64_635 ();
 sg13g2_decap_8 FILLER_64_642 ();
 sg13g2_fill_1 FILLER_64_649 ();
 sg13g2_fill_1 FILLER_64_655 ();
 sg13g2_fill_2 FILLER_64_688 ();
 sg13g2_fill_2 FILLER_64_719 ();
 sg13g2_fill_2 FILLER_64_726 ();
 sg13g2_decap_8 FILLER_64_768 ();
 sg13g2_decap_8 FILLER_64_775 ();
 sg13g2_decap_8 FILLER_64_782 ();
 sg13g2_decap_8 FILLER_64_789 ();
 sg13g2_decap_8 FILLER_64_796 ();
 sg13g2_decap_8 FILLER_64_803 ();
 sg13g2_decap_8 FILLER_64_810 ();
 sg13g2_decap_8 FILLER_64_817 ();
 sg13g2_decap_8 FILLER_64_824 ();
 sg13g2_decap_8 FILLER_64_831 ();
 sg13g2_decap_8 FILLER_64_838 ();
 sg13g2_decap_8 FILLER_64_845 ();
 sg13g2_decap_8 FILLER_64_852 ();
 sg13g2_fill_2 FILLER_64_859 ();
 sg13g2_fill_1 FILLER_64_861 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_4 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_15 ();
 sg13g2_fill_1 FILLER_65_40 ();
 sg13g2_decap_8 FILLER_65_81 ();
 sg13g2_fill_1 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_111 ();
 sg13g2_decap_8 FILLER_65_118 ();
 sg13g2_fill_1 FILLER_65_125 ();
 sg13g2_fill_1 FILLER_65_139 ();
 sg13g2_fill_2 FILLER_65_163 ();
 sg13g2_fill_1 FILLER_65_170 ();
 sg13g2_fill_2 FILLER_65_175 ();
 sg13g2_fill_2 FILLER_65_186 ();
 sg13g2_fill_1 FILLER_65_188 ();
 sg13g2_fill_2 FILLER_65_193 ();
 sg13g2_fill_1 FILLER_65_195 ();
 sg13g2_decap_8 FILLER_65_216 ();
 sg13g2_fill_2 FILLER_65_223 ();
 sg13g2_fill_1 FILLER_65_225 ();
 sg13g2_fill_2 FILLER_65_247 ();
 sg13g2_decap_8 FILLER_65_268 ();
 sg13g2_decap_8 FILLER_65_275 ();
 sg13g2_fill_1 FILLER_65_282 ();
 sg13g2_decap_8 FILLER_65_300 ();
 sg13g2_decap_4 FILLER_65_307 ();
 sg13g2_decap_4 FILLER_65_320 ();
 sg13g2_fill_2 FILLER_65_353 ();
 sg13g2_decap_8 FILLER_65_361 ();
 sg13g2_fill_2 FILLER_65_368 ();
 sg13g2_fill_1 FILLER_65_382 ();
 sg13g2_fill_2 FILLER_65_389 ();
 sg13g2_fill_1 FILLER_65_391 ();
 sg13g2_fill_2 FILLER_65_405 ();
 sg13g2_fill_2 FILLER_65_422 ();
 sg13g2_fill_2 FILLER_65_429 ();
 sg13g2_decap_4 FILLER_65_439 ();
 sg13g2_decap_4 FILLER_65_477 ();
 sg13g2_fill_2 FILLER_65_481 ();
 sg13g2_fill_1 FILLER_65_488 ();
 sg13g2_decap_8 FILLER_65_559 ();
 sg13g2_decap_4 FILLER_65_581 ();
 sg13g2_decap_8 FILLER_65_599 ();
 sg13g2_fill_1 FILLER_65_620 ();
 sg13g2_fill_2 FILLER_65_661 ();
 sg13g2_fill_1 FILLER_65_663 ();
 sg13g2_decap_8 FILLER_65_690 ();
 sg13g2_fill_1 FILLER_65_741 ();
 sg13g2_decap_8 FILLER_65_755 ();
 sg13g2_decap_8 FILLER_65_762 ();
 sg13g2_decap_8 FILLER_65_769 ();
 sg13g2_decap_8 FILLER_65_776 ();
 sg13g2_decap_8 FILLER_65_783 ();
 sg13g2_decap_8 FILLER_65_790 ();
 sg13g2_decap_8 FILLER_65_797 ();
 sg13g2_decap_8 FILLER_65_804 ();
 sg13g2_decap_8 FILLER_65_811 ();
 sg13g2_decap_8 FILLER_65_818 ();
 sg13g2_decap_8 FILLER_65_825 ();
 sg13g2_decap_8 FILLER_65_832 ();
 sg13g2_decap_8 FILLER_65_839 ();
 sg13g2_decap_8 FILLER_65_846 ();
 sg13g2_decap_8 FILLER_65_853 ();
 sg13g2_fill_2 FILLER_65_860 ();
 sg13g2_fill_1 FILLER_66_26 ();
 sg13g2_fill_2 FILLER_66_41 ();
 sg13g2_fill_1 FILLER_66_43 ();
 sg13g2_decap_8 FILLER_66_52 ();
 sg13g2_decap_4 FILLER_66_59 ();
 sg13g2_fill_1 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_69 ();
 sg13g2_decap_8 FILLER_66_76 ();
 sg13g2_fill_2 FILLER_66_83 ();
 sg13g2_fill_1 FILLER_66_85 ();
 sg13g2_decap_4 FILLER_66_112 ();
 sg13g2_fill_1 FILLER_66_147 ();
 sg13g2_decap_4 FILLER_66_168 ();
 sg13g2_fill_1 FILLER_66_172 ();
 sg13g2_decap_8 FILLER_66_181 ();
 sg13g2_fill_2 FILLER_66_188 ();
 sg13g2_fill_1 FILLER_66_199 ();
 sg13g2_decap_4 FILLER_66_218 ();
 sg13g2_decap_4 FILLER_66_227 ();
 sg13g2_fill_1 FILLER_66_231 ();
 sg13g2_decap_8 FILLER_66_243 ();
 sg13g2_fill_1 FILLER_66_271 ();
 sg13g2_decap_8 FILLER_66_299 ();
 sg13g2_fill_1 FILLER_66_306 ();
 sg13g2_decap_8 FILLER_66_346 ();
 sg13g2_decap_8 FILLER_66_365 ();
 sg13g2_decap_8 FILLER_66_380 ();
 sg13g2_fill_1 FILLER_66_393 ();
 sg13g2_fill_2 FILLER_66_409 ();
 sg13g2_decap_4 FILLER_66_430 ();
 sg13g2_decap_8 FILLER_66_439 ();
 sg13g2_decap_4 FILLER_66_468 ();
 sg13g2_fill_1 FILLER_66_472 ();
 sg13g2_fill_1 FILLER_66_501 ();
 sg13g2_fill_2 FILLER_66_521 ();
 sg13g2_fill_2 FILLER_66_528 ();
 sg13g2_fill_1 FILLER_66_530 ();
 sg13g2_fill_2 FILLER_66_536 ();
 sg13g2_fill_1 FILLER_66_538 ();
 sg13g2_decap_4 FILLER_66_548 ();
 sg13g2_decap_4 FILLER_66_563 ();
 sg13g2_fill_1 FILLER_66_567 ();
 sg13g2_fill_1 FILLER_66_572 ();
 sg13g2_fill_1 FILLER_66_590 ();
 sg13g2_decap_8 FILLER_66_612 ();
 sg13g2_decap_4 FILLER_66_619 ();
 sg13g2_decap_4 FILLER_66_651 ();
 sg13g2_fill_2 FILLER_66_655 ();
 sg13g2_decap_4 FILLER_66_667 ();
 sg13g2_fill_1 FILLER_66_671 ();
 sg13g2_decap_4 FILLER_66_706 ();
 sg13g2_decap_8 FILLER_66_745 ();
 sg13g2_decap_8 FILLER_66_752 ();
 sg13g2_decap_8 FILLER_66_759 ();
 sg13g2_decap_8 FILLER_66_766 ();
 sg13g2_decap_8 FILLER_66_773 ();
 sg13g2_decap_8 FILLER_66_780 ();
 sg13g2_decap_8 FILLER_66_787 ();
 sg13g2_decap_8 FILLER_66_794 ();
 sg13g2_decap_8 FILLER_66_801 ();
 sg13g2_decap_8 FILLER_66_808 ();
 sg13g2_decap_8 FILLER_66_815 ();
 sg13g2_decap_8 FILLER_66_822 ();
 sg13g2_decap_8 FILLER_66_829 ();
 sg13g2_decap_8 FILLER_66_836 ();
 sg13g2_decap_8 FILLER_66_843 ();
 sg13g2_decap_8 FILLER_66_850 ();
 sg13g2_decap_4 FILLER_66_857 ();
 sg13g2_fill_1 FILLER_66_861 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_7 ();
 sg13g2_decap_4 FILLER_67_105 ();
 sg13g2_fill_1 FILLER_67_109 ();
 sg13g2_fill_2 FILLER_67_115 ();
 sg13g2_fill_1 FILLER_67_117 ();
 sg13g2_fill_2 FILLER_67_160 ();
 sg13g2_fill_1 FILLER_67_188 ();
 sg13g2_fill_2 FILLER_67_214 ();
 sg13g2_fill_1 FILLER_67_216 ();
 sg13g2_decap_8 FILLER_67_233 ();
 sg13g2_decap_8 FILLER_67_240 ();
 sg13g2_fill_1 FILLER_67_264 ();
 sg13g2_fill_2 FILLER_67_270 ();
 sg13g2_fill_1 FILLER_67_272 ();
 sg13g2_decap_8 FILLER_67_301 ();
 sg13g2_fill_1 FILLER_67_322 ();
 sg13g2_decap_8 FILLER_67_343 ();
 sg13g2_fill_1 FILLER_67_396 ();
 sg13g2_fill_1 FILLER_67_405 ();
 sg13g2_fill_2 FILLER_67_416 ();
 sg13g2_fill_1 FILLER_67_418 ();
 sg13g2_decap_8 FILLER_67_423 ();
 sg13g2_decap_8 FILLER_67_430 ();
 sg13g2_decap_4 FILLER_67_468 ();
 sg13g2_fill_1 FILLER_67_472 ();
 sg13g2_fill_1 FILLER_67_499 ();
 sg13g2_fill_2 FILLER_67_552 ();
 sg13g2_fill_2 FILLER_67_567 ();
 sg13g2_fill_2 FILLER_67_593 ();
 sg13g2_fill_1 FILLER_67_612 ();
 sg13g2_decap_8 FILLER_67_618 ();
 sg13g2_fill_2 FILLER_67_625 ();
 sg13g2_fill_1 FILLER_67_637 ();
 sg13g2_fill_2 FILLER_67_642 ();
 sg13g2_fill_1 FILLER_67_672 ();
 sg13g2_fill_1 FILLER_67_687 ();
 sg13g2_fill_1 FILLER_67_697 ();
 sg13g2_fill_2 FILLER_67_706 ();
 sg13g2_decap_8 FILLER_67_741 ();
 sg13g2_decap_8 FILLER_67_748 ();
 sg13g2_decap_8 FILLER_67_755 ();
 sg13g2_decap_8 FILLER_67_762 ();
 sg13g2_decap_8 FILLER_67_769 ();
 sg13g2_decap_8 FILLER_67_776 ();
 sg13g2_decap_8 FILLER_67_783 ();
 sg13g2_decap_8 FILLER_67_790 ();
 sg13g2_decap_8 FILLER_67_797 ();
 sg13g2_decap_8 FILLER_67_804 ();
 sg13g2_decap_8 FILLER_67_811 ();
 sg13g2_decap_8 FILLER_67_818 ();
 sg13g2_decap_8 FILLER_67_825 ();
 sg13g2_decap_8 FILLER_67_832 ();
 sg13g2_decap_8 FILLER_67_839 ();
 sg13g2_decap_8 FILLER_67_846 ();
 sg13g2_decap_8 FILLER_67_853 ();
 sg13g2_fill_2 FILLER_67_860 ();
 sg13g2_decap_4 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_4 ();
 sg13g2_decap_8 FILLER_68_31 ();
 sg13g2_fill_1 FILLER_68_38 ();
 sg13g2_fill_1 FILLER_68_76 ();
 sg13g2_fill_1 FILLER_68_131 ();
 sg13g2_fill_2 FILLER_68_137 ();
 sg13g2_fill_2 FILLER_68_148 ();
 sg13g2_fill_1 FILLER_68_150 ();
 sg13g2_decap_4 FILLER_68_205 ();
 sg13g2_fill_1 FILLER_68_230 ();
 sg13g2_fill_1 FILLER_68_292 ();
 sg13g2_fill_2 FILLER_68_331 ();
 sg13g2_fill_1 FILLER_68_333 ();
 sg13g2_fill_1 FILLER_68_362 ();
 sg13g2_fill_1 FILLER_68_367 ();
 sg13g2_decap_8 FILLER_68_376 ();
 sg13g2_fill_2 FILLER_68_383 ();
 sg13g2_decap_4 FILLER_68_400 ();
 sg13g2_decap_4 FILLER_68_409 ();
 sg13g2_fill_2 FILLER_68_413 ();
 sg13g2_fill_1 FILLER_68_425 ();
 sg13g2_decap_4 FILLER_68_431 ();
 sg13g2_fill_2 FILLER_68_440 ();
 sg13g2_decap_8 FILLER_68_457 ();
 sg13g2_decap_4 FILLER_68_464 ();
 sg13g2_fill_1 FILLER_68_468 ();
 sg13g2_fill_1 FILLER_68_473 ();
 sg13g2_decap_4 FILLER_68_493 ();
 sg13g2_fill_2 FILLER_68_515 ();
 sg13g2_fill_1 FILLER_68_517 ();
 sg13g2_decap_4 FILLER_68_532 ();
 sg13g2_decap_4 FILLER_68_540 ();
 sg13g2_fill_2 FILLER_68_544 ();
 sg13g2_decap_4 FILLER_68_568 ();
 sg13g2_fill_2 FILLER_68_582 ();
 sg13g2_fill_1 FILLER_68_584 ();
 sg13g2_fill_2 FILLER_68_590 ();
 sg13g2_fill_2 FILLER_68_609 ();
 sg13g2_fill_2 FILLER_68_624 ();
 sg13g2_fill_1 FILLER_68_626 ();
 sg13g2_decap_4 FILLER_68_653 ();
 sg13g2_decap_4 FILLER_68_674 ();
 sg13g2_fill_1 FILLER_68_704 ();
 sg13g2_decap_8 FILLER_68_740 ();
 sg13g2_decap_8 FILLER_68_747 ();
 sg13g2_decap_8 FILLER_68_754 ();
 sg13g2_decap_8 FILLER_68_761 ();
 sg13g2_decap_8 FILLER_68_768 ();
 sg13g2_decap_8 FILLER_68_775 ();
 sg13g2_decap_8 FILLER_68_782 ();
 sg13g2_decap_8 FILLER_68_789 ();
 sg13g2_decap_8 FILLER_68_796 ();
 sg13g2_decap_8 FILLER_68_803 ();
 sg13g2_decap_8 FILLER_68_810 ();
 sg13g2_decap_8 FILLER_68_817 ();
 sg13g2_decap_8 FILLER_68_824 ();
 sg13g2_decap_8 FILLER_68_831 ();
 sg13g2_decap_8 FILLER_68_838 ();
 sg13g2_decap_8 FILLER_68_845 ();
 sg13g2_decap_8 FILLER_68_852 ();
 sg13g2_fill_2 FILLER_68_859 ();
 sg13g2_fill_1 FILLER_68_861 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_4 FILLER_69_37 ();
 sg13g2_fill_1 FILLER_69_41 ();
 sg13g2_fill_1 FILLER_69_71 ();
 sg13g2_fill_2 FILLER_69_87 ();
 sg13g2_fill_1 FILLER_69_89 ();
 sg13g2_fill_2 FILLER_69_109 ();
 sg13g2_fill_1 FILLER_69_111 ();
 sg13g2_fill_2 FILLER_69_138 ();
 sg13g2_fill_2 FILLER_69_191 ();
 sg13g2_fill_1 FILLER_69_193 ();
 sg13g2_decap_4 FILLER_69_203 ();
 sg13g2_decap_8 FILLER_69_233 ();
 sg13g2_fill_2 FILLER_69_240 ();
 sg13g2_decap_8 FILLER_69_246 ();
 sg13g2_decap_8 FILLER_69_253 ();
 sg13g2_fill_2 FILLER_69_260 ();
 sg13g2_fill_1 FILLER_69_262 ();
 sg13g2_fill_2 FILLER_69_268 ();
 sg13g2_fill_1 FILLER_69_270 ();
 sg13g2_decap_8 FILLER_69_279 ();
 sg13g2_fill_2 FILLER_69_286 ();
 sg13g2_fill_1 FILLER_69_288 ();
 sg13g2_fill_1 FILLER_69_307 ();
 sg13g2_fill_2 FILLER_69_312 ();
 sg13g2_decap_4 FILLER_69_322 ();
 sg13g2_decap_4 FILLER_69_332 ();
 sg13g2_fill_1 FILLER_69_336 ();
 sg13g2_decap_8 FILLER_69_345 ();
 sg13g2_fill_2 FILLER_69_352 ();
 sg13g2_fill_1 FILLER_69_354 ();
 sg13g2_decap_8 FILLER_69_388 ();
 sg13g2_decap_8 FILLER_69_395 ();
 sg13g2_decap_8 FILLER_69_402 ();
 sg13g2_fill_1 FILLER_69_409 ();
 sg13g2_fill_1 FILLER_69_426 ();
 sg13g2_decap_4 FILLER_69_437 ();
 sg13g2_fill_2 FILLER_69_441 ();
 sg13g2_fill_1 FILLER_69_457 ();
 sg13g2_fill_2 FILLER_69_489 ();
 sg13g2_decap_4 FILLER_69_522 ();
 sg13g2_fill_1 FILLER_69_526 ();
 sg13g2_fill_1 FILLER_69_540 ();
 sg13g2_fill_1 FILLER_69_552 ();
 sg13g2_decap_4 FILLER_69_558 ();
 sg13g2_fill_2 FILLER_69_595 ();
 sg13g2_decap_8 FILLER_69_646 ();
 sg13g2_decap_4 FILLER_69_653 ();
 sg13g2_fill_1 FILLER_69_682 ();
 sg13g2_fill_1 FILLER_69_692 ();
 sg13g2_decap_8 FILLER_69_719 ();
 sg13g2_decap_8 FILLER_69_726 ();
 sg13g2_decap_8 FILLER_69_733 ();
 sg13g2_decap_8 FILLER_69_740 ();
 sg13g2_decap_8 FILLER_69_747 ();
 sg13g2_decap_8 FILLER_69_754 ();
 sg13g2_decap_8 FILLER_69_761 ();
 sg13g2_decap_8 FILLER_69_768 ();
 sg13g2_decap_8 FILLER_69_775 ();
 sg13g2_decap_8 FILLER_69_782 ();
 sg13g2_decap_8 FILLER_69_789 ();
 sg13g2_decap_8 FILLER_69_796 ();
 sg13g2_decap_8 FILLER_69_803 ();
 sg13g2_decap_8 FILLER_69_810 ();
 sg13g2_decap_8 FILLER_69_817 ();
 sg13g2_decap_8 FILLER_69_824 ();
 sg13g2_decap_8 FILLER_69_831 ();
 sg13g2_decap_8 FILLER_69_838 ();
 sg13g2_decap_8 FILLER_69_845 ();
 sg13g2_decap_8 FILLER_69_852 ();
 sg13g2_fill_2 FILLER_69_859 ();
 sg13g2_fill_1 FILLER_69_861 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_4 FILLER_70_7 ();
 sg13g2_fill_1 FILLER_70_23 ();
 sg13g2_fill_2 FILLER_70_37 ();
 sg13g2_fill_2 FILLER_70_54 ();
 sg13g2_decap_8 FILLER_70_62 ();
 sg13g2_fill_2 FILLER_70_74 ();
 sg13g2_decap_8 FILLER_70_89 ();
 sg13g2_fill_1 FILLER_70_96 ();
 sg13g2_decap_8 FILLER_70_109 ();
 sg13g2_fill_1 FILLER_70_116 ();
 sg13g2_fill_2 FILLER_70_168 ();
 sg13g2_fill_1 FILLER_70_231 ();
 sg13g2_fill_1 FILLER_70_258 ();
 sg13g2_fill_2 FILLER_70_316 ();
 sg13g2_fill_2 FILLER_70_326 ();
 sg13g2_fill_1 FILLER_70_348 ();
 sg13g2_fill_1 FILLER_70_354 ();
 sg13g2_fill_1 FILLER_70_359 ();
 sg13g2_fill_1 FILLER_70_365 ();
 sg13g2_decap_8 FILLER_70_376 ();
 sg13g2_fill_2 FILLER_70_383 ();
 sg13g2_fill_2 FILLER_70_427 ();
 sg13g2_decap_4 FILLER_70_448 ();
 sg13g2_fill_2 FILLER_70_452 ();
 sg13g2_decap_4 FILLER_70_480 ();
 sg13g2_fill_1 FILLER_70_484 ();
 sg13g2_decap_8 FILLER_70_489 ();
 sg13g2_fill_1 FILLER_70_496 ();
 sg13g2_fill_2 FILLER_70_502 ();
 sg13g2_fill_2 FILLER_70_509 ();
 sg13g2_fill_1 FILLER_70_511 ();
 sg13g2_fill_1 FILLER_70_536 ();
 sg13g2_fill_2 FILLER_70_560 ();
 sg13g2_fill_1 FILLER_70_579 ();
 sg13g2_decap_8 FILLER_70_585 ();
 sg13g2_fill_2 FILLER_70_592 ();
 sg13g2_fill_1 FILLER_70_594 ();
 sg13g2_decap_4 FILLER_70_599 ();
 sg13g2_fill_2 FILLER_70_603 ();
 sg13g2_fill_1 FILLER_70_654 ();
 sg13g2_decap_4 FILLER_70_698 ();
 sg13g2_fill_2 FILLER_70_702 ();
 sg13g2_decap_8 FILLER_70_708 ();
 sg13g2_decap_8 FILLER_70_715 ();
 sg13g2_decap_8 FILLER_70_722 ();
 sg13g2_decap_8 FILLER_70_729 ();
 sg13g2_decap_8 FILLER_70_736 ();
 sg13g2_decap_8 FILLER_70_743 ();
 sg13g2_decap_8 FILLER_70_750 ();
 sg13g2_decap_8 FILLER_70_757 ();
 sg13g2_decap_8 FILLER_70_764 ();
 sg13g2_decap_8 FILLER_70_771 ();
 sg13g2_decap_8 FILLER_70_778 ();
 sg13g2_decap_8 FILLER_70_785 ();
 sg13g2_decap_8 FILLER_70_792 ();
 sg13g2_decap_8 FILLER_70_799 ();
 sg13g2_decap_8 FILLER_70_806 ();
 sg13g2_decap_8 FILLER_70_813 ();
 sg13g2_decap_8 FILLER_70_820 ();
 sg13g2_decap_8 FILLER_70_827 ();
 sg13g2_decap_8 FILLER_70_834 ();
 sg13g2_decap_8 FILLER_70_841 ();
 sg13g2_decap_8 FILLER_70_848 ();
 sg13g2_decap_8 FILLER_70_855 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_2 ();
 sg13g2_fill_2 FILLER_71_26 ();
 sg13g2_fill_1 FILLER_71_28 ();
 sg13g2_fill_1 FILLER_71_43 ();
 sg13g2_fill_2 FILLER_71_57 ();
 sg13g2_fill_1 FILLER_71_59 ();
 sg13g2_decap_4 FILLER_71_74 ();
 sg13g2_decap_8 FILLER_71_83 ();
 sg13g2_fill_2 FILLER_71_124 ();
 sg13g2_fill_1 FILLER_71_148 ();
 sg13g2_fill_1 FILLER_71_164 ();
 sg13g2_fill_2 FILLER_71_174 ();
 sg13g2_fill_1 FILLER_71_180 ();
 sg13g2_fill_2 FILLER_71_202 ();
 sg13g2_fill_1 FILLER_71_230 ();
 sg13g2_decap_4 FILLER_71_238 ();
 sg13g2_fill_1 FILLER_71_250 ();
 sg13g2_fill_2 FILLER_71_256 ();
 sg13g2_fill_1 FILLER_71_258 ();
 sg13g2_fill_1 FILLER_71_274 ();
 sg13g2_decap_4 FILLER_71_282 ();
 sg13g2_fill_1 FILLER_71_286 ();
 sg13g2_decap_4 FILLER_71_328 ();
 sg13g2_fill_2 FILLER_71_362 ();
 sg13g2_fill_2 FILLER_71_369 ();
 sg13g2_decap_8 FILLER_71_379 ();
 sg13g2_fill_1 FILLER_71_386 ();
 sg13g2_fill_2 FILLER_71_406 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_fill_1 FILLER_71_418 ();
 sg13g2_decap_8 FILLER_71_457 ();
 sg13g2_fill_2 FILLER_71_464 ();
 sg13g2_fill_1 FILLER_71_466 ();
 sg13g2_fill_2 FILLER_71_472 ();
 sg13g2_decap_4 FILLER_71_505 ();
 sg13g2_fill_1 FILLER_71_514 ();
 sg13g2_decap_4 FILLER_71_545 ();
 sg13g2_fill_1 FILLER_71_549 ();
 sg13g2_fill_2 FILLER_71_556 ();
 sg13g2_decap_4 FILLER_71_582 ();
 sg13g2_fill_1 FILLER_71_586 ();
 sg13g2_fill_2 FILLER_71_591 ();
 sg13g2_fill_2 FILLER_71_610 ();
 sg13g2_fill_1 FILLER_71_612 ();
 sg13g2_fill_2 FILLER_71_628 ();
 sg13g2_fill_2 FILLER_71_639 ();
 sg13g2_fill_1 FILLER_71_641 ();
 sg13g2_decap_8 FILLER_71_677 ();
 sg13g2_decap_8 FILLER_71_692 ();
 sg13g2_decap_8 FILLER_71_699 ();
 sg13g2_decap_8 FILLER_71_706 ();
 sg13g2_decap_8 FILLER_71_713 ();
 sg13g2_decap_8 FILLER_71_720 ();
 sg13g2_decap_8 FILLER_71_727 ();
 sg13g2_decap_8 FILLER_71_734 ();
 sg13g2_decap_8 FILLER_71_741 ();
 sg13g2_decap_8 FILLER_71_748 ();
 sg13g2_decap_8 FILLER_71_755 ();
 sg13g2_decap_8 FILLER_71_762 ();
 sg13g2_decap_8 FILLER_71_769 ();
 sg13g2_decap_8 FILLER_71_776 ();
 sg13g2_decap_8 FILLER_71_783 ();
 sg13g2_decap_8 FILLER_71_790 ();
 sg13g2_decap_8 FILLER_71_797 ();
 sg13g2_decap_8 FILLER_71_804 ();
 sg13g2_decap_8 FILLER_71_811 ();
 sg13g2_decap_8 FILLER_71_818 ();
 sg13g2_decap_8 FILLER_71_825 ();
 sg13g2_decap_8 FILLER_71_832 ();
 sg13g2_decap_8 FILLER_71_839 ();
 sg13g2_decap_8 FILLER_71_846 ();
 sg13g2_decap_8 FILLER_71_853 ();
 sg13g2_fill_2 FILLER_71_860 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_22 ();
 sg13g2_fill_2 FILLER_72_33 ();
 sg13g2_fill_1 FILLER_72_35 ();
 sg13g2_fill_2 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_fill_2 FILLER_72_98 ();
 sg13g2_fill_1 FILLER_72_100 ();
 sg13g2_fill_2 FILLER_72_105 ();
 sg13g2_fill_1 FILLER_72_107 ();
 sg13g2_decap_4 FILLER_72_120 ();
 sg13g2_fill_2 FILLER_72_124 ();
 sg13g2_fill_2 FILLER_72_183 ();
 sg13g2_fill_2 FILLER_72_268 ();
 sg13g2_fill_1 FILLER_72_283 ();
 sg13g2_fill_1 FILLER_72_356 ();
 sg13g2_decap_8 FILLER_72_365 ();
 sg13g2_decap_8 FILLER_72_372 ();
 sg13g2_decap_8 FILLER_72_379 ();
 sg13g2_fill_2 FILLER_72_394 ();
 sg13g2_fill_2 FILLER_72_431 ();
 sg13g2_decap_4 FILLER_72_438 ();
 sg13g2_decap_8 FILLER_72_447 ();
 sg13g2_fill_2 FILLER_72_454 ();
 sg13g2_fill_2 FILLER_72_488 ();
 sg13g2_fill_1 FILLER_72_504 ();
 sg13g2_fill_2 FILLER_72_520 ();
 sg13g2_fill_1 FILLER_72_522 ();
 sg13g2_decap_8 FILLER_72_551 ();
 sg13g2_decap_4 FILLER_72_562 ();
 sg13g2_decap_8 FILLER_72_576 ();
 sg13g2_fill_2 FILLER_72_583 ();
 sg13g2_fill_1 FILLER_72_585 ();
 sg13g2_decap_4 FILLER_72_600 ();
 sg13g2_fill_2 FILLER_72_604 ();
 sg13g2_fill_2 FILLER_72_649 ();
 sg13g2_fill_1 FILLER_72_651 ();
 sg13g2_decap_8 FILLER_72_683 ();
 sg13g2_decap_8 FILLER_72_690 ();
 sg13g2_decap_8 FILLER_72_697 ();
 sg13g2_decap_8 FILLER_72_704 ();
 sg13g2_decap_8 FILLER_72_711 ();
 sg13g2_decap_8 FILLER_72_718 ();
 sg13g2_decap_8 FILLER_72_725 ();
 sg13g2_decap_8 FILLER_72_732 ();
 sg13g2_decap_8 FILLER_72_739 ();
 sg13g2_decap_8 FILLER_72_746 ();
 sg13g2_decap_8 FILLER_72_753 ();
 sg13g2_decap_8 FILLER_72_760 ();
 sg13g2_decap_8 FILLER_72_767 ();
 sg13g2_decap_8 FILLER_72_774 ();
 sg13g2_decap_8 FILLER_72_781 ();
 sg13g2_decap_8 FILLER_72_788 ();
 sg13g2_decap_8 FILLER_72_795 ();
 sg13g2_decap_8 FILLER_72_802 ();
 sg13g2_decap_8 FILLER_72_809 ();
 sg13g2_decap_8 FILLER_72_816 ();
 sg13g2_decap_8 FILLER_72_823 ();
 sg13g2_decap_8 FILLER_72_830 ();
 sg13g2_decap_8 FILLER_72_837 ();
 sg13g2_decap_8 FILLER_72_844 ();
 sg13g2_decap_8 FILLER_72_851 ();
 sg13g2_decap_4 FILLER_72_858 ();
 sg13g2_fill_1 FILLER_73_26 ();
 sg13g2_decap_4 FILLER_73_39 ();
 sg13g2_fill_2 FILLER_73_43 ();
 sg13g2_decap_8 FILLER_73_96 ();
 sg13g2_fill_2 FILLER_73_103 ();
 sg13g2_fill_1 FILLER_73_131 ();
 sg13g2_decap_4 FILLER_73_159 ();
 sg13g2_fill_1 FILLER_73_197 ();
 sg13g2_fill_2 FILLER_73_243 ();
 sg13g2_fill_1 FILLER_73_245 ();
 sg13g2_fill_1 FILLER_73_260 ();
 sg13g2_fill_2 FILLER_73_287 ();
 sg13g2_fill_2 FILLER_73_303 ();
 sg13g2_fill_1 FILLER_73_314 ();
 sg13g2_fill_2 FILLER_73_354 ();
 sg13g2_fill_1 FILLER_73_356 ();
 sg13g2_decap_8 FILLER_73_393 ();
 sg13g2_fill_1 FILLER_73_400 ();
 sg13g2_fill_2 FILLER_73_411 ();
 sg13g2_fill_1 FILLER_73_413 ();
 sg13g2_fill_2 FILLER_73_427 ();
 sg13g2_fill_1 FILLER_73_438 ();
 sg13g2_decap_4 FILLER_73_470 ();
 sg13g2_fill_1 FILLER_73_474 ();
 sg13g2_decap_4 FILLER_73_555 ();
 sg13g2_fill_1 FILLER_73_559 ();
 sg13g2_fill_2 FILLER_73_575 ();
 sg13g2_fill_1 FILLER_73_577 ();
 sg13g2_fill_2 FILLER_73_600 ();
 sg13g2_fill_1 FILLER_73_617 ();
 sg13g2_fill_1 FILLER_73_627 ();
 sg13g2_decap_8 FILLER_73_653 ();
 sg13g2_fill_2 FILLER_73_660 ();
 sg13g2_decap_8 FILLER_73_666 ();
 sg13g2_decap_8 FILLER_73_673 ();
 sg13g2_decap_8 FILLER_73_680 ();
 sg13g2_fill_2 FILLER_73_687 ();
 sg13g2_fill_1 FILLER_73_689 ();
 sg13g2_decap_8 FILLER_73_698 ();
 sg13g2_decap_8 FILLER_73_705 ();
 sg13g2_decap_8 FILLER_73_712 ();
 sg13g2_decap_8 FILLER_73_719 ();
 sg13g2_decap_8 FILLER_73_726 ();
 sg13g2_decap_8 FILLER_73_733 ();
 sg13g2_decap_8 FILLER_73_740 ();
 sg13g2_decap_8 FILLER_73_747 ();
 sg13g2_decap_8 FILLER_73_754 ();
 sg13g2_decap_8 FILLER_73_761 ();
 sg13g2_decap_8 FILLER_73_768 ();
 sg13g2_decap_8 FILLER_73_775 ();
 sg13g2_decap_8 FILLER_73_782 ();
 sg13g2_decap_8 FILLER_73_789 ();
 sg13g2_decap_8 FILLER_73_796 ();
 sg13g2_decap_8 FILLER_73_803 ();
 sg13g2_decap_8 FILLER_73_810 ();
 sg13g2_decap_8 FILLER_73_817 ();
 sg13g2_decap_8 FILLER_73_824 ();
 sg13g2_decap_8 FILLER_73_831 ();
 sg13g2_decap_8 FILLER_73_838 ();
 sg13g2_decap_8 FILLER_73_845 ();
 sg13g2_decap_8 FILLER_73_852 ();
 sg13g2_fill_2 FILLER_73_859 ();
 sg13g2_fill_1 FILLER_73_861 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_7 ();
 sg13g2_fill_2 FILLER_74_15 ();
 sg13g2_decap_8 FILLER_74_51 ();
 sg13g2_fill_2 FILLER_74_118 ();
 sg13g2_fill_1 FILLER_74_120 ();
 sg13g2_decap_4 FILLER_74_151 ();
 sg13g2_fill_2 FILLER_74_199 ();
 sg13g2_fill_1 FILLER_74_201 ();
 sg13g2_fill_2 FILLER_74_211 ();
 sg13g2_fill_2 FILLER_74_232 ();
 sg13g2_fill_2 FILLER_74_261 ();
 sg13g2_fill_1 FILLER_74_272 ();
 sg13g2_fill_2 FILLER_74_282 ();
 sg13g2_fill_1 FILLER_74_315 ();
 sg13g2_fill_2 FILLER_74_325 ();
 sg13g2_fill_2 FILLER_74_340 ();
 sg13g2_fill_2 FILLER_74_347 ();
 sg13g2_decap_4 FILLER_74_353 ();
 sg13g2_fill_2 FILLER_74_357 ();
 sg13g2_fill_2 FILLER_74_364 ();
 sg13g2_fill_1 FILLER_74_405 ();
 sg13g2_fill_1 FILLER_74_416 ();
 sg13g2_decap_4 FILLER_74_448 ();
 sg13g2_fill_1 FILLER_74_452 ();
 sg13g2_decap_4 FILLER_74_462 ();
 sg13g2_fill_1 FILLER_74_466 ();
 sg13g2_fill_2 FILLER_74_512 ();
 sg13g2_fill_1 FILLER_74_514 ();
 sg13g2_decap_8 FILLER_74_585 ();
 sg13g2_fill_1 FILLER_74_592 ();
 sg13g2_fill_2 FILLER_74_613 ();
 sg13g2_decap_8 FILLER_74_667 ();
 sg13g2_decap_8 FILLER_74_674 ();
 sg13g2_decap_8 FILLER_74_681 ();
 sg13g2_decap_8 FILLER_74_688 ();
 sg13g2_decap_8 FILLER_74_695 ();
 sg13g2_decap_8 FILLER_74_702 ();
 sg13g2_decap_8 FILLER_74_709 ();
 sg13g2_decap_8 FILLER_74_716 ();
 sg13g2_decap_8 FILLER_74_723 ();
 sg13g2_decap_8 FILLER_74_730 ();
 sg13g2_decap_8 FILLER_74_737 ();
 sg13g2_decap_8 FILLER_74_744 ();
 sg13g2_decap_8 FILLER_74_751 ();
 sg13g2_decap_8 FILLER_74_758 ();
 sg13g2_decap_8 FILLER_74_765 ();
 sg13g2_decap_8 FILLER_74_772 ();
 sg13g2_decap_8 FILLER_74_779 ();
 sg13g2_decap_8 FILLER_74_786 ();
 sg13g2_decap_8 FILLER_74_793 ();
 sg13g2_decap_8 FILLER_74_800 ();
 sg13g2_decap_8 FILLER_74_807 ();
 sg13g2_decap_8 FILLER_74_814 ();
 sg13g2_decap_8 FILLER_74_821 ();
 sg13g2_decap_8 FILLER_74_828 ();
 sg13g2_decap_8 FILLER_74_835 ();
 sg13g2_decap_8 FILLER_74_842 ();
 sg13g2_decap_8 FILLER_74_849 ();
 sg13g2_decap_4 FILLER_74_856 ();
 sg13g2_fill_2 FILLER_74_860 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_4 FILLER_75_60 ();
 sg13g2_fill_1 FILLER_75_64 ();
 sg13g2_decap_8 FILLER_75_73 ();
 sg13g2_fill_2 FILLER_75_80 ();
 sg13g2_decap_4 FILLER_75_90 ();
 sg13g2_fill_2 FILLER_75_94 ();
 sg13g2_fill_1 FILLER_75_112 ();
 sg13g2_fill_2 FILLER_75_139 ();
 sg13g2_fill_1 FILLER_75_172 ();
 sg13g2_fill_1 FILLER_75_187 ();
 sg13g2_fill_2 FILLER_75_289 ();
 sg13g2_fill_1 FILLER_75_291 ();
 sg13g2_fill_2 FILLER_75_297 ();
 sg13g2_fill_1 FILLER_75_299 ();
 sg13g2_fill_2 FILLER_75_335 ();
 sg13g2_fill_1 FILLER_75_337 ();
 sg13g2_decap_8 FILLER_75_364 ();
 sg13g2_fill_2 FILLER_75_371 ();
 sg13g2_fill_1 FILLER_75_373 ();
 sg13g2_decap_4 FILLER_75_379 ();
 sg13g2_fill_1 FILLER_75_386 ();
 sg13g2_fill_2 FILLER_75_412 ();
 sg13g2_decap_4 FILLER_75_429 ();
 sg13g2_fill_2 FILLER_75_433 ();
 sg13g2_decap_4 FILLER_75_444 ();
 sg13g2_fill_2 FILLER_75_448 ();
 sg13g2_fill_2 FILLER_75_465 ();
 sg13g2_decap_4 FILLER_75_493 ();
 sg13g2_fill_1 FILLER_75_497 ();
 sg13g2_fill_1 FILLER_75_524 ();
 sg13g2_decap_8 FILLER_75_545 ();
 sg13g2_decap_8 FILLER_75_552 ();
 sg13g2_fill_1 FILLER_75_585 ();
 sg13g2_decap_4 FILLER_75_607 ();
 sg13g2_fill_2 FILLER_75_611 ();
 sg13g2_decap_8 FILLER_75_627 ();
 sg13g2_fill_1 FILLER_75_634 ();
 sg13g2_decap_8 FILLER_75_639 ();
 sg13g2_decap_8 FILLER_75_646 ();
 sg13g2_decap_8 FILLER_75_653 ();
 sg13g2_decap_8 FILLER_75_660 ();
 sg13g2_decap_8 FILLER_75_667 ();
 sg13g2_decap_8 FILLER_75_674 ();
 sg13g2_decap_8 FILLER_75_681 ();
 sg13g2_decap_8 FILLER_75_688 ();
 sg13g2_decap_8 FILLER_75_695 ();
 sg13g2_decap_8 FILLER_75_702 ();
 sg13g2_decap_8 FILLER_75_709 ();
 sg13g2_decap_8 FILLER_75_716 ();
 sg13g2_decap_8 FILLER_75_723 ();
 sg13g2_decap_8 FILLER_75_730 ();
 sg13g2_decap_8 FILLER_75_737 ();
 sg13g2_decap_8 FILLER_75_744 ();
 sg13g2_decap_8 FILLER_75_751 ();
 sg13g2_decap_8 FILLER_75_758 ();
 sg13g2_decap_8 FILLER_75_765 ();
 sg13g2_decap_8 FILLER_75_772 ();
 sg13g2_decap_8 FILLER_75_779 ();
 sg13g2_decap_8 FILLER_75_786 ();
 sg13g2_decap_8 FILLER_75_793 ();
 sg13g2_decap_8 FILLER_75_800 ();
 sg13g2_decap_8 FILLER_75_807 ();
 sg13g2_decap_8 FILLER_75_814 ();
 sg13g2_decap_8 FILLER_75_821 ();
 sg13g2_decap_8 FILLER_75_828 ();
 sg13g2_decap_8 FILLER_75_835 ();
 sg13g2_decap_8 FILLER_75_842 ();
 sg13g2_decap_8 FILLER_75_849 ();
 sg13g2_decap_4 FILLER_75_856 ();
 sg13g2_fill_2 FILLER_75_860 ();
 sg13g2_fill_2 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_2 ();
 sg13g2_fill_1 FILLER_76_29 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_fill_2 FILLER_76_42 ();
 sg13g2_fill_1 FILLER_76_44 ();
 sg13g2_fill_1 FILLER_76_49 ();
 sg13g2_fill_1 FILLER_76_115 ();
 sg13g2_decap_4 FILLER_76_136 ();
 sg13g2_fill_2 FILLER_76_140 ();
 sg13g2_fill_2 FILLER_76_146 ();
 sg13g2_fill_1 FILLER_76_148 ();
 sg13g2_fill_2 FILLER_76_166 ();
 sg13g2_fill_2 FILLER_76_187 ();
 sg13g2_fill_2 FILLER_76_219 ();
 sg13g2_fill_1 FILLER_76_221 ();
 sg13g2_fill_2 FILLER_76_254 ();
 sg13g2_fill_2 FILLER_76_270 ();
 sg13g2_fill_1 FILLER_76_272 ();
 sg13g2_decap_4 FILLER_76_281 ();
 sg13g2_decap_4 FILLER_76_300 ();
 sg13g2_fill_2 FILLER_76_340 ();
 sg13g2_fill_1 FILLER_76_342 ();
 sg13g2_fill_1 FILLER_76_352 ();
 sg13g2_fill_2 FILLER_76_406 ();
 sg13g2_fill_2 FILLER_76_435 ();
 sg13g2_decap_8 FILLER_76_446 ();
 sg13g2_fill_2 FILLER_76_479 ();
 sg13g2_fill_2 FILLER_76_520 ();
 sg13g2_fill_1 FILLER_76_522 ();
 sg13g2_decap_4 FILLER_76_548 ();
 sg13g2_fill_2 FILLER_76_552 ();
 sg13g2_fill_1 FILLER_76_559 ();
 sg13g2_fill_1 FILLER_76_571 ();
 sg13g2_fill_1 FILLER_76_576 ();
 sg13g2_fill_2 FILLER_76_582 ();
 sg13g2_fill_1 FILLER_76_584 ();
 sg13g2_fill_1 FILLER_76_594 ();
 sg13g2_fill_2 FILLER_76_599 ();
 sg13g2_fill_1 FILLER_76_601 ();
 sg13g2_decap_4 FILLER_76_627 ();
 sg13g2_fill_1 FILLER_76_631 ();
 sg13g2_decap_8 FILLER_76_636 ();
 sg13g2_decap_8 FILLER_76_643 ();
 sg13g2_decap_8 FILLER_76_650 ();
 sg13g2_decap_8 FILLER_76_657 ();
 sg13g2_decap_8 FILLER_76_664 ();
 sg13g2_decap_8 FILLER_76_671 ();
 sg13g2_decap_8 FILLER_76_678 ();
 sg13g2_decap_8 FILLER_76_685 ();
 sg13g2_decap_8 FILLER_76_692 ();
 sg13g2_decap_8 FILLER_76_699 ();
 sg13g2_decap_8 FILLER_76_706 ();
 sg13g2_decap_8 FILLER_76_713 ();
 sg13g2_decap_8 FILLER_76_720 ();
 sg13g2_decap_8 FILLER_76_727 ();
 sg13g2_decap_8 FILLER_76_734 ();
 sg13g2_decap_8 FILLER_76_741 ();
 sg13g2_decap_8 FILLER_76_748 ();
 sg13g2_decap_8 FILLER_76_755 ();
 sg13g2_decap_8 FILLER_76_762 ();
 sg13g2_decap_8 FILLER_76_769 ();
 sg13g2_decap_8 FILLER_76_776 ();
 sg13g2_decap_8 FILLER_76_783 ();
 sg13g2_decap_8 FILLER_76_790 ();
 sg13g2_decap_8 FILLER_76_797 ();
 sg13g2_decap_8 FILLER_76_804 ();
 sg13g2_decap_8 FILLER_76_811 ();
 sg13g2_decap_8 FILLER_76_818 ();
 sg13g2_decap_8 FILLER_76_825 ();
 sg13g2_decap_8 FILLER_76_832 ();
 sg13g2_decap_8 FILLER_76_839 ();
 sg13g2_decap_8 FILLER_76_846 ();
 sg13g2_decap_8 FILLER_76_853 ();
 sg13g2_fill_2 FILLER_76_860 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_4 FILLER_77_7 ();
 sg13g2_fill_2 FILLER_77_11 ();
 sg13g2_fill_2 FILLER_77_17 ();
 sg13g2_fill_2 FILLER_77_23 ();
 sg13g2_fill_1 FILLER_77_33 ();
 sg13g2_fill_2 FILLER_77_68 ();
 sg13g2_fill_1 FILLER_77_70 ();
 sg13g2_fill_2 FILLER_77_79 ();
 sg13g2_fill_1 FILLER_77_81 ();
 sg13g2_fill_1 FILLER_77_157 ();
 sg13g2_fill_2 FILLER_77_187 ();
 sg13g2_fill_2 FILLER_77_200 ();
 sg13g2_fill_2 FILLER_77_226 ();
 sg13g2_fill_2 FILLER_77_242 ();
 sg13g2_fill_2 FILLER_77_274 ();
 sg13g2_fill_1 FILLER_77_311 ();
 sg13g2_fill_2 FILLER_77_336 ();
 sg13g2_fill_1 FILLER_77_462 ();
 sg13g2_fill_2 FILLER_77_480 ();
 sg13g2_fill_1 FILLER_77_491 ();
 sg13g2_fill_2 FILLER_77_554 ();
 sg13g2_fill_2 FILLER_77_586 ();
 sg13g2_fill_2 FILLER_77_598 ();
 sg13g2_fill_2 FILLER_77_620 ();
 sg13g2_decap_8 FILLER_77_648 ();
 sg13g2_decap_8 FILLER_77_655 ();
 sg13g2_decap_8 FILLER_77_662 ();
 sg13g2_decap_8 FILLER_77_669 ();
 sg13g2_decap_8 FILLER_77_676 ();
 sg13g2_decap_8 FILLER_77_683 ();
 sg13g2_decap_8 FILLER_77_690 ();
 sg13g2_decap_8 FILLER_77_697 ();
 sg13g2_decap_8 FILLER_77_704 ();
 sg13g2_decap_8 FILLER_77_711 ();
 sg13g2_decap_8 FILLER_77_718 ();
 sg13g2_decap_8 FILLER_77_725 ();
 sg13g2_decap_8 FILLER_77_732 ();
 sg13g2_decap_8 FILLER_77_739 ();
 sg13g2_decap_8 FILLER_77_746 ();
 sg13g2_decap_8 FILLER_77_753 ();
 sg13g2_decap_8 FILLER_77_760 ();
 sg13g2_decap_8 FILLER_77_767 ();
 sg13g2_decap_8 FILLER_77_774 ();
 sg13g2_decap_8 FILLER_77_781 ();
 sg13g2_decap_8 FILLER_77_788 ();
 sg13g2_decap_8 FILLER_77_795 ();
 sg13g2_decap_8 FILLER_77_802 ();
 sg13g2_decap_8 FILLER_77_809 ();
 sg13g2_decap_8 FILLER_77_816 ();
 sg13g2_decap_8 FILLER_77_823 ();
 sg13g2_decap_8 FILLER_77_830 ();
 sg13g2_decap_8 FILLER_77_837 ();
 sg13g2_decap_8 FILLER_77_844 ();
 sg13g2_decap_8 FILLER_77_851 ();
 sg13g2_decap_4 FILLER_77_858 ();
 sg13g2_fill_1 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_4 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_54 ();
 sg13g2_fill_2 FILLER_78_65 ();
 sg13g2_fill_1 FILLER_78_67 ();
 sg13g2_fill_2 FILLER_78_118 ();
 sg13g2_fill_2 FILLER_78_129 ();
 sg13g2_fill_1 FILLER_78_131 ();
 sg13g2_fill_2 FILLER_78_182 ();
 sg13g2_fill_1 FILLER_78_184 ();
 sg13g2_fill_2 FILLER_78_191 ();
 sg13g2_fill_1 FILLER_78_193 ();
 sg13g2_fill_2 FILLER_78_261 ();
 sg13g2_fill_2 FILLER_78_268 ();
 sg13g2_fill_1 FILLER_78_270 ();
 sg13g2_decap_4 FILLER_78_275 ();
 sg13g2_decap_4 FILLER_78_305 ();
 sg13g2_decap_4 FILLER_78_369 ();
 sg13g2_fill_1 FILLER_78_373 ();
 sg13g2_decap_8 FILLER_78_382 ();
 sg13g2_fill_2 FILLER_78_389 ();
 sg13g2_decap_8 FILLER_78_395 ();
 sg13g2_decap_8 FILLER_78_402 ();
 sg13g2_decap_8 FILLER_78_409 ();
 sg13g2_fill_2 FILLER_78_416 ();
 sg13g2_fill_1 FILLER_78_418 ();
 sg13g2_decap_8 FILLER_78_423 ();
 sg13g2_decap_8 FILLER_78_430 ();
 sg13g2_fill_1 FILLER_78_437 ();
 sg13g2_decap_4 FILLER_78_442 ();
 sg13g2_decap_4 FILLER_78_476 ();
 sg13g2_fill_1 FILLER_78_480 ();
 sg13g2_fill_2 FILLER_78_485 ();
 sg13g2_fill_1 FILLER_78_487 ();
 sg13g2_fill_2 FILLER_78_497 ();
 sg13g2_fill_1 FILLER_78_499 ();
 sg13g2_decap_8 FILLER_78_521 ();
 sg13g2_decap_8 FILLER_78_528 ();
 sg13g2_fill_2 FILLER_78_550 ();
 sg13g2_decap_8 FILLER_78_578 ();
 sg13g2_fill_2 FILLER_78_585 ();
 sg13g2_fill_1 FILLER_78_587 ();
 sg13g2_fill_2 FILLER_78_593 ();
 sg13g2_fill_1 FILLER_78_595 ();
 sg13g2_decap_8 FILLER_78_632 ();
 sg13g2_decap_8 FILLER_78_639 ();
 sg13g2_decap_8 FILLER_78_646 ();
 sg13g2_decap_8 FILLER_78_653 ();
 sg13g2_decap_8 FILLER_78_660 ();
 sg13g2_decap_8 FILLER_78_667 ();
 sg13g2_decap_8 FILLER_78_674 ();
 sg13g2_decap_8 FILLER_78_681 ();
 sg13g2_decap_8 FILLER_78_688 ();
 sg13g2_decap_8 FILLER_78_695 ();
 sg13g2_decap_8 FILLER_78_702 ();
 sg13g2_decap_8 FILLER_78_709 ();
 sg13g2_decap_8 FILLER_78_716 ();
 sg13g2_decap_8 FILLER_78_723 ();
 sg13g2_decap_8 FILLER_78_730 ();
 sg13g2_decap_8 FILLER_78_737 ();
 sg13g2_decap_8 FILLER_78_744 ();
 sg13g2_decap_8 FILLER_78_751 ();
 sg13g2_decap_8 FILLER_78_758 ();
 sg13g2_decap_8 FILLER_78_765 ();
 sg13g2_decap_8 FILLER_78_772 ();
 sg13g2_decap_8 FILLER_78_779 ();
 sg13g2_decap_8 FILLER_78_786 ();
 sg13g2_decap_8 FILLER_78_793 ();
 sg13g2_decap_8 FILLER_78_800 ();
 sg13g2_decap_8 FILLER_78_807 ();
 sg13g2_decap_8 FILLER_78_814 ();
 sg13g2_decap_8 FILLER_78_821 ();
 sg13g2_decap_8 FILLER_78_828 ();
 sg13g2_decap_8 FILLER_78_835 ();
 sg13g2_decap_8 FILLER_78_842 ();
 sg13g2_decap_8 FILLER_78_849 ();
 sg13g2_decap_4 FILLER_78_856 ();
 sg13g2_fill_2 FILLER_78_860 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_4 FILLER_79_7 ();
 sg13g2_fill_1 FILLER_79_11 ();
 sg13g2_fill_2 FILLER_79_112 ();
 sg13g2_fill_1 FILLER_79_114 ();
 sg13g2_fill_2 FILLER_79_151 ();
 sg13g2_fill_1 FILLER_79_166 ();
 sg13g2_decap_4 FILLER_79_206 ();
 sg13g2_fill_1 FILLER_79_210 ();
 sg13g2_fill_2 FILLER_79_224 ();
 sg13g2_fill_1 FILLER_79_226 ();
 sg13g2_fill_2 FILLER_79_231 ();
 sg13g2_decap_4 FILLER_79_289 ();
 sg13g2_decap_8 FILLER_79_362 ();
 sg13g2_decap_8 FILLER_79_369 ();
 sg13g2_decap_8 FILLER_79_376 ();
 sg13g2_decap_8 FILLER_79_383 ();
 sg13g2_decap_8 FILLER_79_390 ();
 sg13g2_decap_8 FILLER_79_397 ();
 sg13g2_decap_8 FILLER_79_404 ();
 sg13g2_decap_8 FILLER_79_411 ();
 sg13g2_decap_8 FILLER_79_418 ();
 sg13g2_decap_8 FILLER_79_425 ();
 sg13g2_decap_8 FILLER_79_432 ();
 sg13g2_decap_8 FILLER_79_439 ();
 sg13g2_decap_8 FILLER_79_446 ();
 sg13g2_decap_4 FILLER_79_453 ();
 sg13g2_decap_8 FILLER_79_461 ();
 sg13g2_decap_8 FILLER_79_468 ();
 sg13g2_fill_1 FILLER_79_475 ();
 sg13g2_fill_2 FILLER_79_519 ();
 sg13g2_fill_1 FILLER_79_521 ();
 sg13g2_fill_2 FILLER_79_535 ();
 sg13g2_fill_1 FILLER_79_537 ();
 sg13g2_fill_1 FILLER_79_542 ();
 sg13g2_fill_2 FILLER_79_548 ();
 sg13g2_fill_2 FILLER_79_559 ();
 sg13g2_fill_1 FILLER_79_561 ();
 sg13g2_decap_8 FILLER_79_590 ();
 sg13g2_decap_4 FILLER_79_597 ();
 sg13g2_decap_4 FILLER_79_606 ();
 sg13g2_fill_1 FILLER_79_610 ();
 sg13g2_decap_8 FILLER_79_624 ();
 sg13g2_decap_8 FILLER_79_631 ();
 sg13g2_decap_8 FILLER_79_638 ();
 sg13g2_decap_8 FILLER_79_645 ();
 sg13g2_decap_8 FILLER_79_652 ();
 sg13g2_decap_8 FILLER_79_659 ();
 sg13g2_decap_8 FILLER_79_666 ();
 sg13g2_decap_8 FILLER_79_673 ();
 sg13g2_decap_8 FILLER_79_680 ();
 sg13g2_decap_8 FILLER_79_687 ();
 sg13g2_decap_8 FILLER_79_694 ();
 sg13g2_decap_8 FILLER_79_701 ();
 sg13g2_decap_8 FILLER_79_708 ();
 sg13g2_decap_8 FILLER_79_715 ();
 sg13g2_decap_8 FILLER_79_722 ();
 sg13g2_decap_8 FILLER_79_729 ();
 sg13g2_decap_8 FILLER_79_736 ();
 sg13g2_decap_8 FILLER_79_743 ();
 sg13g2_decap_8 FILLER_79_750 ();
 sg13g2_decap_8 FILLER_79_757 ();
 sg13g2_decap_8 FILLER_79_764 ();
 sg13g2_decap_8 FILLER_79_771 ();
 sg13g2_decap_8 FILLER_79_778 ();
 sg13g2_decap_8 FILLER_79_785 ();
 sg13g2_decap_8 FILLER_79_792 ();
 sg13g2_decap_8 FILLER_79_799 ();
 sg13g2_decap_8 FILLER_79_806 ();
 sg13g2_decap_8 FILLER_79_813 ();
 sg13g2_decap_8 FILLER_79_820 ();
 sg13g2_decap_8 FILLER_79_827 ();
 sg13g2_decap_8 FILLER_79_834 ();
 sg13g2_decap_8 FILLER_79_841 ();
 sg13g2_decap_8 FILLER_79_848 ();
 sg13g2_decap_8 FILLER_79_855 ();
 sg13g2_fill_2 FILLER_80_0 ();
 sg13g2_fill_1 FILLER_80_2 ();
 sg13g2_decap_8 FILLER_80_41 ();
 sg13g2_decap_8 FILLER_80_48 ();
 sg13g2_fill_2 FILLER_80_55 ();
 sg13g2_decap_4 FILLER_80_61 ();
 sg13g2_fill_1 FILLER_80_65 ();
 sg13g2_fill_2 FILLER_80_96 ();
 sg13g2_fill_2 FILLER_80_138 ();
 sg13g2_decap_8 FILLER_80_205 ();
 sg13g2_decap_8 FILLER_80_212 ();
 sg13g2_fill_1 FILLER_80_245 ();
 sg13g2_decap_8 FILLER_80_262 ();
 sg13g2_decap_4 FILLER_80_269 ();
 sg13g2_fill_1 FILLER_80_273 ();
 sg13g2_decap_8 FILLER_80_278 ();
 sg13g2_decap_4 FILLER_80_285 ();
 sg13g2_fill_1 FILLER_80_289 ();
 sg13g2_decap_8 FILLER_80_294 ();
 sg13g2_decap_8 FILLER_80_301 ();
 sg13g2_fill_1 FILLER_80_317 ();
 sg13g2_fill_2 FILLER_80_338 ();
 sg13g2_fill_1 FILLER_80_340 ();
 sg13g2_fill_2 FILLER_80_346 ();
 sg13g2_decap_4 FILLER_80_356 ();
 sg13g2_fill_2 FILLER_80_365 ();
 sg13g2_fill_1 FILLER_80_367 ();
 sg13g2_decap_8 FILLER_80_373 ();
 sg13g2_decap_8 FILLER_80_380 ();
 sg13g2_decap_8 FILLER_80_387 ();
 sg13g2_decap_8 FILLER_80_394 ();
 sg13g2_decap_8 FILLER_80_401 ();
 sg13g2_decap_8 FILLER_80_408 ();
 sg13g2_decap_8 FILLER_80_415 ();
 sg13g2_decap_8 FILLER_80_422 ();
 sg13g2_decap_8 FILLER_80_429 ();
 sg13g2_decap_8 FILLER_80_436 ();
 sg13g2_decap_8 FILLER_80_443 ();
 sg13g2_decap_8 FILLER_80_450 ();
 sg13g2_decap_8 FILLER_80_457 ();
 sg13g2_decap_8 FILLER_80_464 ();
 sg13g2_decap_8 FILLER_80_471 ();
 sg13g2_decap_8 FILLER_80_478 ();
 sg13g2_decap_8 FILLER_80_485 ();
 sg13g2_decap_8 FILLER_80_492 ();
 sg13g2_fill_2 FILLER_80_525 ();
 sg13g2_decap_8 FILLER_80_553 ();
 sg13g2_fill_2 FILLER_80_560 ();
 sg13g2_decap_8 FILLER_80_588 ();
 sg13g2_decap_8 FILLER_80_595 ();
 sg13g2_decap_8 FILLER_80_602 ();
 sg13g2_decap_8 FILLER_80_609 ();
 sg13g2_decap_8 FILLER_80_616 ();
 sg13g2_decap_8 FILLER_80_623 ();
 sg13g2_decap_8 FILLER_80_630 ();
 sg13g2_decap_8 FILLER_80_637 ();
 sg13g2_decap_8 FILLER_80_644 ();
 sg13g2_decap_8 FILLER_80_651 ();
 sg13g2_decap_8 FILLER_80_658 ();
 sg13g2_decap_8 FILLER_80_665 ();
 sg13g2_decap_8 FILLER_80_672 ();
 sg13g2_decap_8 FILLER_80_679 ();
 sg13g2_decap_8 FILLER_80_686 ();
 sg13g2_decap_8 FILLER_80_693 ();
 sg13g2_decap_8 FILLER_80_700 ();
 sg13g2_decap_8 FILLER_80_707 ();
 sg13g2_decap_8 FILLER_80_714 ();
 sg13g2_decap_8 FILLER_80_721 ();
 sg13g2_decap_8 FILLER_80_728 ();
 sg13g2_decap_8 FILLER_80_735 ();
 sg13g2_decap_8 FILLER_80_742 ();
 sg13g2_decap_8 FILLER_80_749 ();
 sg13g2_decap_8 FILLER_80_756 ();
 sg13g2_decap_8 FILLER_80_763 ();
 sg13g2_decap_8 FILLER_80_770 ();
 sg13g2_decap_8 FILLER_80_777 ();
 sg13g2_decap_8 FILLER_80_784 ();
 sg13g2_decap_8 FILLER_80_791 ();
 sg13g2_decap_8 FILLER_80_798 ();
 sg13g2_decap_8 FILLER_80_805 ();
 sg13g2_decap_8 FILLER_80_812 ();
 sg13g2_decap_8 FILLER_80_819 ();
 sg13g2_decap_8 FILLER_80_826 ();
 sg13g2_decap_8 FILLER_80_833 ();
 sg13g2_decap_8 FILLER_80_840 ();
 sg13g2_decap_8 FILLER_80_847 ();
 sg13g2_decap_8 FILLER_80_854 ();
 sg13g2_fill_1 FILLER_80_861 ();
endmodule

module tt_um_jayjaywong12 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[10][0] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[11][0] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[12][0] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[13][0] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[14][0] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[15][0] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[16][0] ;
 wire \mem[16][1] ;
 wire \mem[16][2] ;
 wire \mem[16][3] ;
 wire \mem[17][0] ;
 wire \mem[17][1] ;
 wire \mem[17][2] ;
 wire \mem[17][3] ;
 wire \mem[18][0] ;
 wire \mem[18][1] ;
 wire \mem[18][2] ;
 wire \mem[18][3] ;
 wire \mem[19][0] ;
 wire \mem[19][1] ;
 wire \mem[19][2] ;
 wire \mem[19][3] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[20][0] ;
 wire \mem[20][1] ;
 wire \mem[20][2] ;
 wire \mem[20][3] ;
 wire \mem[21][0] ;
 wire \mem[21][1] ;
 wire \mem[21][2] ;
 wire \mem[21][3] ;
 wire \mem[22][0] ;
 wire \mem[22][1] ;
 wire \mem[22][2] ;
 wire \mem[22][3] ;
 wire \mem[23][0] ;
 wire \mem[23][1] ;
 wire \mem[23][2] ;
 wire \mem[23][3] ;
 wire \mem[24][0] ;
 wire \mem[24][1] ;
 wire \mem[24][2] ;
 wire \mem[24][3] ;
 wire \mem[25][0] ;
 wire \mem[25][1] ;
 wire \mem[25][2] ;
 wire \mem[25][3] ;
 wire \mem[26][0] ;
 wire \mem[26][1] ;
 wire \mem[26][2] ;
 wire \mem[26][3] ;
 wire \mem[27][0] ;
 wire \mem[27][1] ;
 wire \mem[27][2] ;
 wire \mem[27][3] ;
 wire \mem[28][0] ;
 wire \mem[28][1] ;
 wire \mem[28][2] ;
 wire \mem[28][3] ;
 wire \mem[29][0] ;
 wire \mem[29][1] ;
 wire \mem[29][2] ;
 wire \mem[29][3] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[30][0] ;
 wire \mem[30][1] ;
 wire \mem[30][2] ;
 wire \mem[30][3] ;
 wire \mem[31][0] ;
 wire \mem[31][1] ;
 wire \mem[31][2] ;
 wire \mem[31][3] ;
 wire \mem[32][0] ;
 wire \mem[32][1] ;
 wire \mem[32][2] ;
 wire \mem[32][3] ;
 wire \mem[35][0] ;
 wire \mem[35][1] ;
 wire \mem[35][2] ;
 wire \mem[35][3] ;
 wire \mem[36][0] ;
 wire \mem[36][1] ;
 wire \mem[36][2] ;
 wire \mem[36][3] ;
 wire \mem[37][0] ;
 wire \mem[37][1] ;
 wire \mem[37][2] ;
 wire \mem[37][3] ;
 wire \mem[38][0] ;
 wire \mem[38][1] ;
 wire \mem[38][2] ;
 wire \mem[38][3] ;
 wire \mem[39][0] ;
 wire \mem[39][1] ;
 wire \mem[39][2] ;
 wire \mem[39][3] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[40][0] ;
 wire \mem[40][1] ;
 wire \mem[40][2] ;
 wire \mem[40][3] ;
 wire \mem[41][0] ;
 wire \mem[41][1] ;
 wire \mem[41][2] ;
 wire \mem[41][3] ;
 wire \mem[42][0] ;
 wire \mem[42][1] ;
 wire \mem[42][2] ;
 wire \mem[42][3] ;
 wire \mem[43][0] ;
 wire \mem[43][1] ;
 wire \mem[43][2] ;
 wire \mem[43][3] ;
 wire \mem[44][0] ;
 wire \mem[44][1] ;
 wire \mem[44][2] ;
 wire \mem[44][3] ;
 wire \mem[45][0] ;
 wire \mem[45][1] ;
 wire \mem[45][2] ;
 wire \mem[45][3] ;
 wire \mem[46][0] ;
 wire \mem[46][1] ;
 wire \mem[46][2] ;
 wire \mem[46][3] ;
 wire \mem[47][0] ;
 wire \mem[47][1] ;
 wire \mem[47][2] ;
 wire \mem[47][3] ;
 wire \mem[48][0] ;
 wire \mem[48][1] ;
 wire \mem[48][2] ;
 wire \mem[48][3] ;
 wire \mem[49][0] ;
 wire \mem[49][1] ;
 wire \mem[49][2] ;
 wire \mem[49][3] ;
 wire \mem[4][0] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[50][0] ;
 wire \mem[50][1] ;
 wire \mem[50][2] ;
 wire \mem[50][3] ;
 wire \mem[51][0] ;
 wire \mem[51][1] ;
 wire \mem[51][2] ;
 wire \mem[51][3] ;
 wire \mem[52][0] ;
 wire \mem[52][1] ;
 wire \mem[52][2] ;
 wire \mem[52][3] ;
 wire \mem[53][0] ;
 wire \mem[53][1] ;
 wire \mem[53][2] ;
 wire \mem[53][3] ;
 wire \mem[54][0] ;
 wire \mem[54][1] ;
 wire \mem[54][2] ;
 wire \mem[54][3] ;
 wire \mem[55][0] ;
 wire \mem[55][1] ;
 wire \mem[55][2] ;
 wire \mem[55][3] ;
 wire \mem[56][0] ;
 wire \mem[56][1] ;
 wire \mem[56][2] ;
 wire \mem[56][3] ;
 wire \mem[57][0] ;
 wire \mem[57][1] ;
 wire \mem[57][2] ;
 wire \mem[57][3] ;
 wire \mem[58][0] ;
 wire \mem[58][1] ;
 wire \mem[58][2] ;
 wire \mem[58][3] ;
 wire \mem[59][0] ;
 wire \mem[59][1] ;
 wire \mem[59][2] ;
 wire \mem[59][3] ;
 wire \mem[5][0] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[60][0] ;
 wire \mem[60][1] ;
 wire \mem[60][2] ;
 wire \mem[60][3] ;
 wire \mem[61][0] ;
 wire \mem[61][1] ;
 wire \mem[61][2] ;
 wire \mem[61][3] ;
 wire \mem[62][0] ;
 wire \mem[62][1] ;
 wire \mem[62][2] ;
 wire \mem[62][3] ;
 wire \mem[63][0] ;
 wire \mem[63][1] ;
 wire \mem[63][2] ;
 wire \mem[63][3] ;
 wire \mem[6][0] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[7][0] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[8][0] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[9][0] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \prev_acc[0] ;
 wire \prev_acc[1] ;
 wire \prev_acc[2] ;
 wire \prev_acc[3] ;
 wire \prev_acc[4] ;
 wire \prev_acc[5] ;
 wire \prev_acc[6] ;
 wire \prev_acc[7] ;
 wire \products[0][0] ;
 wire \products[0][1] ;
 wire \products[0][2] ;
 wire \products[0][3] ;
 wire \products[0][4] ;
 wire \products[0][5] ;
 wire \products[0][6] ;
 wire \products[0][7] ;
 wire \products[10][0] ;
 wire \products[10][1] ;
 wire \products[10][2] ;
 wire \products[10][3] ;
 wire \products[10][4] ;
 wire \products[10][5] ;
 wire \products[10][6] ;
 wire \products[10][7] ;
 wire \products[11][0] ;
 wire \products[11][1] ;
 wire \products[11][2] ;
 wire \products[11][3] ;
 wire \products[11][4] ;
 wire \products[11][5] ;
 wire \products[11][6] ;
 wire \products[11][7] ;
 wire \products[12][0] ;
 wire \products[12][1] ;
 wire \products[12][2] ;
 wire \products[12][3] ;
 wire \products[12][4] ;
 wire \products[12][5] ;
 wire \products[12][6] ;
 wire \products[12][7] ;
 wire \products[13][0] ;
 wire \products[13][1] ;
 wire \products[13][2] ;
 wire \products[13][3] ;
 wire \products[13][4] ;
 wire \products[13][5] ;
 wire \products[13][6] ;
 wire \products[13][7] ;
 wire \products[14][0] ;
 wire \products[14][1] ;
 wire \products[14][2] ;
 wire \products[14][3] ;
 wire \products[14][4] ;
 wire \products[14][5] ;
 wire \products[14][6] ;
 wire \products[14][7] ;
 wire \products[15][0] ;
 wire \products[15][1] ;
 wire \products[15][2] ;
 wire \products[15][3] ;
 wire \products[15][4] ;
 wire \products[15][5] ;
 wire \products[15][6] ;
 wire \products[15][7] ;
 wire \products[1][0] ;
 wire \products[1][1] ;
 wire \products[1][2] ;
 wire \products[1][3] ;
 wire \products[1][4] ;
 wire \products[1][5] ;
 wire \products[1][6] ;
 wire \products[1][7] ;
 wire \products[2][0] ;
 wire \products[2][1] ;
 wire \products[2][2] ;
 wire \products[2][3] ;
 wire \products[2][4] ;
 wire \products[2][5] ;
 wire \products[2][6] ;
 wire \products[2][7] ;
 wire \products[3][0] ;
 wire \products[3][1] ;
 wire \products[3][2] ;
 wire \products[3][3] ;
 wire \products[3][4] ;
 wire \products[3][5] ;
 wire \products[3][6] ;
 wire \products[3][7] ;
 wire \products[4][0] ;
 wire \products[4][1] ;
 wire \products[4][2] ;
 wire \products[4][3] ;
 wire \products[4][4] ;
 wire \products[4][5] ;
 wire \products[4][6] ;
 wire \products[4][7] ;
 wire \products[5][0] ;
 wire \products[5][1] ;
 wire \products[5][2] ;
 wire \products[5][3] ;
 wire \products[5][4] ;
 wire \products[5][5] ;
 wire \products[5][6] ;
 wire \products[5][7] ;
 wire \products[6][0] ;
 wire \products[6][1] ;
 wire \products[6][2] ;
 wire \products[6][3] ;
 wire \products[6][4] ;
 wire \products[6][5] ;
 wire \products[6][6] ;
 wire \products[6][7] ;
 wire \products[7][0] ;
 wire \products[7][1] ;
 wire \products[7][2] ;
 wire \products[7][3] ;
 wire \products[7][4] ;
 wire \products[7][5] ;
 wire \products[7][6] ;
 wire \products[7][7] ;
 wire \products[8][0] ;
 wire \products[8][1] ;
 wire \products[8][2] ;
 wire \products[8][3] ;
 wire \products[8][4] ;
 wire \products[8][5] ;
 wire \products[8][6] ;
 wire \products[8][7] ;
 wire \products[9][0] ;
 wire \products[9][1] ;
 wire \products[9][2] ;
 wire \products[9][3] ;
 wire \products[9][4] ;
 wire \products[9][5] ;
 wire \products[9][6] ;
 wire \products[9][7] ;
 wire read_operation;
 wire net406;
 wire clknet_leaf_0_clk;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;

 sg13g2_inv_1 _3058_ (.Y(_2082_),
    .A(uo_out[7]));
 sg13g2_inv_1 _3059_ (.Y(_2083_),
    .A(uo_out[6]));
 sg13g2_inv_1 _3060_ (.Y(_2084_),
    .A(net703));
 sg13g2_inv_1 _3061_ (.Y(_2085_),
    .A(net822));
 sg13g2_inv_1 _3062_ (.Y(_2086_),
    .A(net693));
 sg13g2_inv_1 _3063_ (.Y(_2087_),
    .A(net691));
 sg13g2_inv_1 _3064_ (.Y(_2088_),
    .A(net721));
 sg13g2_inv_1 _3065_ (.Y(_2089_),
    .A(net711));
 sg13g2_inv_1 _3066_ (.Y(_2090_),
    .A(net407));
 sg13g2_inv_1 _3067_ (.Y(_2091_),
    .A(net2));
 sg13g2_inv_1 _3068_ (.Y(_2092_),
    .A(net552));
 sg13g2_inv_2 _3069_ (.Y(_2093_),
    .A(net536));
 sg13g2_inv_2 _3070_ (.Y(_2094_),
    .A(net531));
 sg13g2_inv_1 _3071_ (.Y(_2095_),
    .A(net528));
 sg13g2_inv_1 _3072_ (.Y(_2096_),
    .A(net680));
 sg13g2_inv_1 _3073_ (.Y(_2097_),
    .A(net674));
 sg13g2_inv_1 _3074_ (.Y(_2098_),
    .A(net745));
 sg13g2_inv_1 _3075_ (.Y(_2099_),
    .A(net796));
 sg13g2_inv_1 _3076_ (.Y(_2100_),
    .A(net688));
 sg13g2_inv_1 _3077_ (.Y(_2101_),
    .A(net632));
 sg13g2_inv_2 _3078_ (.Y(_2102_),
    .A(net732));
 sg13g2_inv_1 _3079_ (.Y(_2103_),
    .A(net840));
 sg13g2_inv_1 _3080_ (.Y(_2104_),
    .A(net831));
 sg13g2_inv_1 _3081_ (.Y(_2105_),
    .A(net729));
 sg13g2_nor2_1 _3082_ (.A(net2),
    .B(net1),
    .Y(read_operation));
 sg13g2_nand2_1 _3083_ (.Y(_2106_),
    .A(net515),
    .B(\mem[44][0] ));
 sg13g2_a21oi_1 _3084_ (.A1(net559),
    .A2(\mem[45][0] ),
    .Y(_2107_),
    .B1(net539));
 sg13g2_nor2b_1 _3085_ (.A(net557),
    .B_N(\mem[46][0] ),
    .Y(_2108_));
 sg13g2_a21oi_1 _3086_ (.A1(net558),
    .A2(\mem[47][0] ),
    .Y(_2109_),
    .B1(_2108_));
 sg13g2_a221oi_1 _3087_ (.B2(net537),
    .C1(net506),
    .B1(_2109_),
    .A1(_2106_),
    .Y(_2110_),
    .A2(_2107_));
 sg13g2_mux4_1 _3088_ (.S0(net558),
    .A0(\mem[40][0] ),
    .A1(\mem[41][0] ),
    .A2(\mem[42][0] ),
    .A3(\mem[43][0] ),
    .S1(net539),
    .X(_2111_));
 sg13g2_and2_1 _3089_ (.A(net506),
    .B(_2111_),
    .X(_2112_));
 sg13g2_o21ai_1 _3090_ (.B1(net528),
    .Y(_2113_),
    .A1(_2110_),
    .A2(_2112_));
 sg13g2_nand2_1 _3091_ (.Y(_2114_),
    .A(net515),
    .B(\mem[36][0] ));
 sg13g2_a21oi_1 _3092_ (.A1(net560),
    .A2(\mem[37][0] ),
    .Y(_2115_),
    .B1(net541));
 sg13g2_nor2b_1 _3093_ (.A(net560),
    .B_N(\mem[38][0] ),
    .Y(_2116_));
 sg13g2_a21oi_1 _3094_ (.A1(net560),
    .A2(\mem[39][0] ),
    .Y(_2117_),
    .B1(_2116_));
 sg13g2_a221oi_1 _3095_ (.B2(net541),
    .C1(net507),
    .B1(_2117_),
    .A1(_2114_),
    .Y(_2118_),
    .A2(_2115_));
 sg13g2_nand2_1 _3096_ (.Y(_2119_),
    .A(net521),
    .B(\mem[32][0] ));
 sg13g2_a21oi_1 _3097_ (.A1(uo_out[0]),
    .A2(net561),
    .Y(_2120_),
    .B1(net542));
 sg13g2_nor2_1 _3098_ (.A(_2085_),
    .B(net561),
    .Y(_2121_));
 sg13g2_a21oi_1 _3099_ (.A1(net561),
    .A2(\mem[35][0] ),
    .Y(_2122_),
    .B1(_2121_));
 sg13g2_a221oi_1 _3100_ (.B2(net541),
    .C1(net532),
    .B1(_2122_),
    .A1(_2119_),
    .Y(_2123_),
    .A2(_2120_));
 sg13g2_o21ai_1 _3101_ (.B1(net503),
    .Y(_2124_),
    .A1(_2118_),
    .A2(_2123_));
 sg13g2_nand3b_1 _3102_ (.B(_2113_),
    .C(_2124_),
    .Y(_2125_),
    .A_N(net526));
 sg13g2_nand2_1 _3103_ (.Y(_2126_),
    .A(net518),
    .B(\mem[60][0] ));
 sg13g2_a21oi_1 _3104_ (.A1(net552),
    .A2(\mem[61][0] ),
    .Y(_2127_),
    .B1(net533));
 sg13g2_nor2b_1 _3105_ (.A(net551),
    .B_N(\mem[62][0] ),
    .Y(_2128_));
 sg13g2_a21oi_1 _3106_ (.A1(net551),
    .A2(\mem[63][0] ),
    .Y(_2129_),
    .B1(_2128_));
 sg13g2_a221oi_1 _3107_ (.B2(net533),
    .C1(net505),
    .B1(_2129_),
    .A1(_2126_),
    .Y(_2130_),
    .A2(_2127_));
 sg13g2_mux4_1 _3108_ (.S0(net553),
    .A0(\mem[56][0] ),
    .A1(\mem[57][0] ),
    .A2(\mem[58][0] ),
    .A3(\mem[59][0] ),
    .S1(net536),
    .X(_2131_));
 sg13g2_and2_1 _3109_ (.A(net509),
    .B(_2131_),
    .X(_2132_));
 sg13g2_o21ai_1 _3110_ (.B1(net527),
    .Y(_2133_),
    .A1(_2130_),
    .A2(_2132_));
 sg13g2_nand2_1 _3111_ (.Y(_2134_),
    .A(net516),
    .B(\mem[52][0] ));
 sg13g2_a21oi_1 _3112_ (.A1(net557),
    .A2(\mem[53][0] ),
    .Y(_2135_),
    .B1(net538));
 sg13g2_nor2b_1 _3113_ (.A(net554),
    .B_N(\mem[54][0] ),
    .Y(_2136_));
 sg13g2_a21oi_1 _3114_ (.A1(net554),
    .A2(\mem[55][0] ),
    .Y(_2137_),
    .B1(_2136_));
 sg13g2_a221oi_1 _3115_ (.B2(net538),
    .C1(net507),
    .B1(_2137_),
    .A1(_2134_),
    .Y(_2138_),
    .A2(_2135_));
 sg13g2_mux4_1 _3116_ (.S0(net556),
    .A0(\mem[48][0] ),
    .A1(\mem[49][0] ),
    .A2(\mem[50][0] ),
    .A3(\mem[51][0] ),
    .S1(net537),
    .X(_2139_));
 sg13g2_and2_1 _3117_ (.A(net507),
    .B(_2139_),
    .X(_2140_));
 sg13g2_o21ai_1 _3118_ (.B1(net502),
    .Y(_2141_),
    .A1(_2138_),
    .A2(_2140_));
 sg13g2_nand3_1 _3119_ (.B(_2133_),
    .C(_2141_),
    .A(net524),
    .Y(_2142_));
 sg13g2_nand3_1 _3120_ (.B(_2125_),
    .C(_2142_),
    .A(net522),
    .Y(_2143_));
 sg13g2_nand2_1 _3121_ (.Y(_2144_),
    .A(net520),
    .B(\mem[28][0] ));
 sg13g2_a21oi_1 _3122_ (.A1(net564),
    .A2(\mem[29][0] ),
    .Y(_2145_),
    .B1(net543));
 sg13g2_nor2b_1 _3123_ (.A(net564),
    .B_N(\mem[30][0] ),
    .Y(_2146_));
 sg13g2_a21oi_1 _3124_ (.A1(net564),
    .A2(\mem[31][0] ),
    .Y(_2147_),
    .B1(_2146_));
 sg13g2_a221oi_1 _3125_ (.B2(net544),
    .C1(net510),
    .B1(_2147_),
    .A1(_2144_),
    .Y(_2148_),
    .A2(_2145_));
 sg13g2_nand2_1 _3126_ (.Y(_2149_),
    .A(net518),
    .B(\mem[24][0] ));
 sg13g2_a21oi_1 _3127_ (.A1(net568),
    .A2(\mem[25][0] ),
    .Y(_2150_),
    .B1(net545));
 sg13g2_nor2b_1 _3128_ (.A(net568),
    .B_N(\mem[26][0] ),
    .Y(_2151_));
 sg13g2_a21oi_1 _3129_ (.A1(net568),
    .A2(\mem[27][0] ),
    .Y(_2152_),
    .B1(_2151_));
 sg13g2_a221oi_1 _3130_ (.B2(net545),
    .C1(net532),
    .B1(_2152_),
    .A1(_2149_),
    .Y(_2153_),
    .A2(_2150_));
 sg13g2_o21ai_1 _3131_ (.B1(net530),
    .Y(_2154_),
    .A1(_2148_),
    .A2(_2153_));
 sg13g2_a21oi_1 _3132_ (.A1(net575),
    .A2(\mem[21][0] ),
    .Y(_2155_),
    .B1(net549));
 sg13g2_o21ai_1 _3133_ (.B1(_2155_),
    .Y(_2156_),
    .A1(net575),
    .A2(_2098_));
 sg13g2_nand2_1 _3134_ (.Y(_2157_),
    .A(net519),
    .B(\mem[22][0] ));
 sg13g2_a21oi_1 _3135_ (.A1(net575),
    .A2(\mem[23][0] ),
    .Y(_2158_),
    .B1(_2093_));
 sg13g2_a21oi_1 _3136_ (.A1(_2157_),
    .A2(_2158_),
    .Y(_2159_),
    .B1(net513));
 sg13g2_mux4_1 _3137_ (.S0(net575),
    .A0(\mem[16][0] ),
    .A1(\mem[17][0] ),
    .A2(\mem[18][0] ),
    .A3(\mem[19][0] ),
    .S1(net549),
    .X(_2160_));
 sg13g2_a22oi_1 _3138_ (.Y(_2161_),
    .B1(_2160_),
    .B2(net513),
    .A2(_2159_),
    .A1(_2156_));
 sg13g2_o21ai_1 _3139_ (.B1(net525),
    .Y(_2162_),
    .A1(net530),
    .A2(_2161_));
 sg13g2_nand2b_1 _3140_ (.Y(_2163_),
    .B(_2154_),
    .A_N(_2162_));
 sg13g2_a21oi_1 _3141_ (.A1(net564),
    .A2(\mem[13][0] ),
    .Y(_2164_),
    .B1(net544));
 sg13g2_o21ai_1 _3142_ (.B1(_2164_),
    .Y(_2165_),
    .A1(net564),
    .A2(_2097_));
 sg13g2_nor2b_1 _3143_ (.A(net567),
    .B_N(net497),
    .Y(_2166_));
 sg13g2_a21oi_1 _3144_ (.A1(net564),
    .A2(net499),
    .Y(_2167_),
    .B1(_2166_));
 sg13g2_a21oi_1 _3145_ (.A1(net544),
    .A2(_2167_),
    .Y(_2168_),
    .B1(net510));
 sg13g2_mux4_1 _3146_ (.S0(net568),
    .A0(\mem[8][0] ),
    .A1(\mem[9][0] ),
    .A2(\mem[10][0] ),
    .A3(\mem[11][0] ),
    .S1(net545),
    .X(_2169_));
 sg13g2_a22oi_1 _3147_ (.Y(_2170_),
    .B1(_2169_),
    .B2(net510),
    .A2(_2168_),
    .A1(_2165_));
 sg13g2_nor2_1 _3148_ (.A(net504),
    .B(_2170_),
    .Y(_2171_));
 sg13g2_a21oi_1 _3149_ (.A1(net572),
    .A2(net495),
    .Y(_2172_),
    .B1(net547));
 sg13g2_o21ai_1 _3150_ (.B1(_2172_),
    .Y(_2173_),
    .A1(net572),
    .A2(_2096_));
 sg13g2_nand2_1 _3151_ (.Y(_2174_),
    .A(net521),
    .B(\mem[6][0] ));
 sg13g2_a21oi_1 _3152_ (.A1(net571),
    .A2(\mem[7][0] ),
    .Y(_2175_),
    .B1(_2093_));
 sg13g2_a21oi_1 _3153_ (.A1(_2174_),
    .A2(_2175_),
    .Y(_2176_),
    .B1(net512));
 sg13g2_mux4_1 _3154_ (.S0(net569),
    .A0(\mem[0][0] ),
    .A1(\mem[1][0] ),
    .A2(\mem[2][0] ),
    .A3(\mem[3][0] ),
    .S1(net547),
    .X(_2177_));
 sg13g2_a22oi_1 _3155_ (.Y(_2178_),
    .B1(_2177_),
    .B2(net512),
    .A2(_2176_),
    .A1(_2173_));
 sg13g2_nor2_1 _3156_ (.A(net529),
    .B(_2178_),
    .Y(_2179_));
 sg13g2_nor3_1 _3157_ (.A(net526),
    .B(_2171_),
    .C(_2179_),
    .Y(_2180_));
 sg13g2_nand2b_1 _3158_ (.Y(_2181_),
    .B(_2163_),
    .A_N(net523));
 sg13g2_o21ai_1 _3159_ (.B1(_2143_),
    .Y(uio_out[0]),
    .A1(_2180_),
    .A2(_2181_));
 sg13g2_nand2_1 _3160_ (.Y(_2182_),
    .A(net515),
    .B(\mem[44][1] ));
 sg13g2_a21oi_1 _3161_ (.A1(net558),
    .A2(\mem[45][1] ),
    .Y(_2183_),
    .B1(net539));
 sg13g2_nor2b_1 _3162_ (.A(net557),
    .B_N(\mem[46][1] ),
    .Y(_2184_));
 sg13g2_a21oi_1 _3163_ (.A1(net558),
    .A2(\mem[47][1] ),
    .Y(_2185_),
    .B1(_2184_));
 sg13g2_a221oi_1 _3164_ (.B2(net537),
    .C1(net506),
    .B1(_2185_),
    .A1(_2182_),
    .Y(_2186_),
    .A2(_2183_));
 sg13g2_mux4_1 _3165_ (.S0(net558),
    .A0(\mem[40][1] ),
    .A1(\mem[41][1] ),
    .A2(\mem[42][1] ),
    .A3(\mem[43][1] ),
    .S1(net539),
    .X(_2187_));
 sg13g2_a21oi_1 _3166_ (.A1(net506),
    .A2(_2187_),
    .Y(_2188_),
    .B1(_2186_));
 sg13g2_nor2_1 _3167_ (.A(net503),
    .B(_2188_),
    .Y(_2189_));
 sg13g2_nand2_1 _3168_ (.Y(_2190_),
    .A(net517),
    .B(\mem[36][1] ));
 sg13g2_a21oi_1 _3169_ (.A1(net560),
    .A2(\mem[37][1] ),
    .Y(_2191_),
    .B1(net541));
 sg13g2_nor2b_1 _3170_ (.A(net560),
    .B_N(\mem[38][1] ),
    .Y(_2192_));
 sg13g2_a21oi_1 _3171_ (.A1(net560),
    .A2(\mem[39][1] ),
    .Y(_2193_),
    .B1(_2192_));
 sg13g2_a221oi_1 _3172_ (.B2(net541),
    .C1(net508),
    .B1(_2193_),
    .A1(_2190_),
    .Y(_2194_),
    .A2(_2191_));
 sg13g2_nand2_1 _3173_ (.Y(_2195_),
    .A(net517),
    .B(\mem[32][1] ));
 sg13g2_a21oi_1 _3174_ (.A1(uo_out[1]),
    .A2(net561),
    .Y(_2196_),
    .B1(net541));
 sg13g2_a21oi_1 _3175_ (.A1(net561),
    .A2(\mem[35][1] ),
    .Y(_2197_),
    .B1(net514));
 sg13g2_o21ai_1 _3176_ (.B1(_2197_),
    .Y(_2198_),
    .A1(_2084_),
    .A2(net561));
 sg13g2_a21oi_1 _3177_ (.A1(_2195_),
    .A2(_2196_),
    .Y(_2199_),
    .B1(net532));
 sg13g2_a21oi_1 _3178_ (.A1(_2198_),
    .A2(_2199_),
    .Y(_2200_),
    .B1(_2194_));
 sg13g2_nor2_1 _3179_ (.A(net528),
    .B(_2200_),
    .Y(_2201_));
 sg13g2_nor3_1 _3180_ (.A(net524),
    .B(_2189_),
    .C(_2201_),
    .Y(_2202_));
 sg13g2_nand2_1 _3181_ (.Y(_2203_),
    .A(net518),
    .B(\mem[60][1] ));
 sg13g2_a21oi_1 _3182_ (.A1(net554),
    .A2(\mem[61][1] ),
    .Y(_2204_),
    .B1(net534));
 sg13g2_nor2b_1 _3183_ (.A(net552),
    .B_N(\mem[62][1] ),
    .Y(_2205_));
 sg13g2_a21oi_1 _3184_ (.A1(net551),
    .A2(\mem[63][1] ),
    .Y(_2206_),
    .B1(_2205_));
 sg13g2_a221oi_1 _3185_ (.B2(net534),
    .C1(net505),
    .B1(_2206_),
    .A1(_2203_),
    .Y(_2207_),
    .A2(_2204_));
 sg13g2_mux4_1 _3186_ (.S0(net554),
    .A0(\mem[56][1] ),
    .A1(\mem[57][1] ),
    .A2(\mem[58][1] ),
    .A3(\mem[59][1] ),
    .S1(net534),
    .X(_2208_));
 sg13g2_a21oi_1 _3187_ (.A1(net505),
    .A2(_2208_),
    .Y(_2209_),
    .B1(_2207_));
 sg13g2_nor2_1 _3188_ (.A(net502),
    .B(_2209_),
    .Y(_2210_));
 sg13g2_a21oi_1 _3189_ (.A1(net562),
    .A2(\mem[53][1] ),
    .Y(_2211_),
    .B1(net542));
 sg13g2_o21ai_1 _3190_ (.B1(_2211_),
    .Y(_2212_),
    .A1(net562),
    .A2(_2101_));
 sg13g2_nand2_1 _3191_ (.Y(_2213_),
    .A(net516),
    .B(\mem[54][1] ));
 sg13g2_a21oi_1 _3192_ (.A1(net555),
    .A2(\mem[55][1] ),
    .Y(_2214_),
    .B1(net514));
 sg13g2_a21oi_1 _3193_ (.A1(_2213_),
    .A2(_2214_),
    .Y(_2215_),
    .B1(net507));
 sg13g2_mux4_1 _3194_ (.S0(net556),
    .A0(\mem[48][1] ),
    .A1(\mem[49][1] ),
    .A2(\mem[50][1] ),
    .A3(\mem[51][1] ),
    .S1(net537),
    .X(_2216_));
 sg13g2_a22oi_1 _3195_ (.Y(_2217_),
    .B1(_2216_),
    .B2(net507),
    .A2(_2215_),
    .A1(_2212_));
 sg13g2_o21ai_1 _3196_ (.B1(net524),
    .Y(_2218_),
    .A1(net528),
    .A2(_2217_));
 sg13g2_o21ai_1 _3197_ (.B1(net522),
    .Y(_2219_),
    .A1(_2210_),
    .A2(_2218_));
 sg13g2_nand2_1 _3198_ (.Y(_2220_),
    .A(net520),
    .B(\mem[28][1] ));
 sg13g2_a21oi_1 _3199_ (.A1(net565),
    .A2(\mem[29][1] ),
    .Y(_2221_),
    .B1(net543));
 sg13g2_nor2b_1 _3200_ (.A(net566),
    .B_N(\mem[30][1] ),
    .Y(_2222_));
 sg13g2_a21oi_1 _3201_ (.A1(net566),
    .A2(\mem[31][1] ),
    .Y(_2223_),
    .B1(_2222_));
 sg13g2_a221oi_1 _3202_ (.B2(net544),
    .C1(net510),
    .B1(_2223_),
    .A1(_2220_),
    .Y(_2224_),
    .A2(_2221_));
 sg13g2_mux4_1 _3203_ (.S0(net568),
    .A0(\mem[24][1] ),
    .A1(\mem[25][1] ),
    .A2(\mem[26][1] ),
    .A3(\mem[27][1] ),
    .S1(net545),
    .X(_2225_));
 sg13g2_a21oi_2 _3204_ (.B1(_2224_),
    .Y(_2226_),
    .A2(_2225_),
    .A1(net511));
 sg13g2_nor2_1 _3205_ (.A(net504),
    .B(_2226_),
    .Y(_2227_));
 sg13g2_a21oi_1 _3206_ (.A1(net570),
    .A2(\mem[21][1] ),
    .Y(_2228_),
    .B1(net546));
 sg13g2_o21ai_1 _3207_ (.B1(_2228_),
    .Y(_2229_),
    .A1(net570),
    .A2(_2100_));
 sg13g2_nand2_1 _3208_ (.Y(_2230_),
    .A(net519),
    .B(\mem[22][1] ));
 sg13g2_a21oi_1 _3209_ (.A1(net569),
    .A2(\mem[23][1] ),
    .Y(_2231_),
    .B1(_2093_));
 sg13g2_a21oi_1 _3210_ (.A1(_2230_),
    .A2(_2231_),
    .Y(_2232_),
    .B1(net512));
 sg13g2_mux4_1 _3211_ (.S0(net575),
    .A0(\mem[16][1] ),
    .A1(\mem[17][1] ),
    .A2(\mem[18][1] ),
    .A3(\mem[19][1] ),
    .S1(net549),
    .X(_2233_));
 sg13g2_a22oi_1 _3212_ (.Y(_2234_),
    .B1(_2233_),
    .B2(net513),
    .A2(_2232_),
    .A1(_2229_));
 sg13g2_o21ai_1 _3213_ (.B1(net525),
    .Y(_2235_),
    .A1(net529),
    .A2(_2234_));
 sg13g2_nand2_1 _3214_ (.Y(_2236_),
    .A(net520),
    .B(\mem[12][1] ));
 sg13g2_a21oi_1 _3215_ (.A1(net566),
    .A2(\mem[13][1] ),
    .Y(_2237_),
    .B1(net543));
 sg13g2_nor2b_1 _3216_ (.A(net566),
    .B_N(net496),
    .Y(_2238_));
 sg13g2_a21oi_1 _3217_ (.A1(net566),
    .A2(net498),
    .Y(_2239_),
    .B1(_2238_));
 sg13g2_a221oi_1 _3218_ (.B2(net543),
    .C1(net511),
    .B1(_2239_),
    .A1(_2236_),
    .Y(_2240_),
    .A2(_2237_));
 sg13g2_mux4_1 _3219_ (.S0(net568),
    .A0(net490),
    .A1(\mem[9][1] ),
    .A2(\mem[10][1] ),
    .A3(\mem[11][1] ),
    .S1(net545),
    .X(_2241_));
 sg13g2_and2_1 _3220_ (.A(net511),
    .B(_2241_),
    .X(_2242_));
 sg13g2_o21ai_1 _3221_ (.B1(net530),
    .Y(_2243_),
    .A1(_2240_),
    .A2(_2242_));
 sg13g2_nand2_1 _3222_ (.Y(_2244_),
    .A(net519),
    .B(\mem[4][1] ));
 sg13g2_a21oi_1 _3223_ (.A1(net571),
    .A2(net494),
    .Y(_2245_),
    .B1(net548));
 sg13g2_nor2b_1 _3224_ (.A(net571),
    .B_N(\mem[6][1] ),
    .Y(_2246_));
 sg13g2_a21oi_1 _3225_ (.A1(net571),
    .A2(\mem[7][1] ),
    .Y(_2247_),
    .B1(_2246_));
 sg13g2_a221oi_1 _3226_ (.B2(net547),
    .C1(net512),
    .B1(_2247_),
    .A1(_2244_),
    .Y(_2248_),
    .A2(_2245_));
 sg13g2_nand2_1 _3227_ (.Y(_2249_),
    .A(\mem[0][1] ),
    .B(net519));
 sg13g2_a21oi_1 _3228_ (.A1(net569),
    .A2(\mem[1][1] ),
    .Y(_2250_),
    .B1(net546));
 sg13g2_nor2b_1 _3229_ (.A(net574),
    .B_N(\mem[2][1] ),
    .Y(_2251_));
 sg13g2_a21oi_1 _3230_ (.A1(net574),
    .A2(\mem[3][1] ),
    .Y(_2252_),
    .B1(_2251_));
 sg13g2_a221oi_1 _3231_ (.B2(net546),
    .C1(net532),
    .B1(_2252_),
    .A1(_2249_),
    .Y(_2253_),
    .A2(_2250_));
 sg13g2_o21ai_1 _3232_ (.B1(net504),
    .Y(_2254_),
    .A1(_2248_),
    .A2(_2253_));
 sg13g2_nor2b_1 _3233_ (.A(net525),
    .B_N(_2254_),
    .Y(_2255_));
 sg13g2_a21oi_1 _3234_ (.A1(_2243_),
    .A2(_2255_),
    .Y(_2256_),
    .B1(net523));
 sg13g2_o21ai_1 _3235_ (.B1(_2256_),
    .Y(_2257_),
    .A1(_2227_),
    .A2(_2235_));
 sg13g2_o21ai_1 _3236_ (.B1(_2257_),
    .Y(uio_out[1]),
    .A1(_2202_),
    .A2(_2219_));
 sg13g2_nand2_1 _3237_ (.Y(_2258_),
    .A(net515),
    .B(\mem[44][2] ));
 sg13g2_a21oi_1 _3238_ (.A1(net556),
    .A2(\mem[45][2] ),
    .Y(_2259_),
    .B1(net537));
 sg13g2_nor2b_1 _3239_ (.A(net556),
    .B_N(\mem[46][2] ),
    .Y(_2260_));
 sg13g2_a21oi_1 _3240_ (.A1(net556),
    .A2(\mem[47][2] ),
    .Y(_2261_),
    .B1(_2260_));
 sg13g2_a221oi_1 _3241_ (.B2(net537),
    .C1(net506),
    .B1(_2261_),
    .A1(_2258_),
    .Y(_2262_),
    .A2(_2259_));
 sg13g2_mux4_1 _3242_ (.S0(net558),
    .A0(\mem[40][2] ),
    .A1(\mem[41][2] ),
    .A2(\mem[42][2] ),
    .A3(\mem[43][2] ),
    .S1(net539),
    .X(_2263_));
 sg13g2_and2_1 _3243_ (.A(net506),
    .B(_2263_),
    .X(_2264_));
 sg13g2_o21ai_1 _3244_ (.B1(net527),
    .Y(_2265_),
    .A1(_2262_),
    .A2(_2264_));
 sg13g2_nand2_1 _3245_ (.Y(_2266_),
    .A(net515),
    .B(\mem[36][2] ));
 sg13g2_a21oi_1 _3246_ (.A1(net560),
    .A2(\mem[37][2] ),
    .Y(_2267_),
    .B1(net539));
 sg13g2_nor2b_1 _3247_ (.A(net559),
    .B_N(\mem[38][2] ),
    .Y(_2268_));
 sg13g2_a21oi_1 _3248_ (.A1(net560),
    .A2(\mem[39][2] ),
    .Y(_2269_),
    .B1(_2268_));
 sg13g2_a221oi_1 _3249_ (.B2(net540),
    .C1(net508),
    .B1(_2269_),
    .A1(_2266_),
    .Y(_2270_),
    .A2(_2267_));
 sg13g2_nand2_1 _3250_ (.Y(_0395_),
    .A(net517),
    .B(\mem[32][2] ));
 sg13g2_a21oi_1 _3251_ (.A1(uo_out[2]),
    .A2(net561),
    .Y(_0396_),
    .B1(net541));
 sg13g2_nand2_1 _3252_ (.Y(_0397_),
    .A(uo_out[6]),
    .B(net517));
 sg13g2_a21oi_1 _3253_ (.A1(net562),
    .A2(\mem[35][2] ),
    .Y(_0398_),
    .B1(net514));
 sg13g2_a221oi_1 _3254_ (.B2(_0398_),
    .C1(net531),
    .B1(_0397_),
    .A1(_0395_),
    .Y(_0399_),
    .A2(_0396_));
 sg13g2_o21ai_1 _3255_ (.B1(net503),
    .Y(_0400_),
    .A1(_2270_),
    .A2(_0399_));
 sg13g2_nand3b_1 _3256_ (.B(_2265_),
    .C(_0400_),
    .Y(_0401_),
    .A_N(net524));
 sg13g2_nand2_1 _3257_ (.Y(_0402_),
    .A(net518),
    .B(\mem[60][2] ));
 sg13g2_a21oi_1 _3258_ (.A1(net552),
    .A2(\mem[61][2] ),
    .Y(_0403_),
    .B1(net533));
 sg13g2_nor2b_1 _3259_ (.A(net551),
    .B_N(\mem[62][2] ),
    .Y(_0404_));
 sg13g2_a21oi_1 _3260_ (.A1(net551),
    .A2(\mem[63][2] ),
    .Y(_0405_),
    .B1(_0404_));
 sg13g2_a221oi_1 _3261_ (.B2(net533),
    .C1(net505),
    .B1(_0405_),
    .A1(_0402_),
    .Y(_0406_),
    .A2(_0403_));
 sg13g2_mux4_1 _3262_ (.S0(net553),
    .A0(\mem[56][2] ),
    .A1(\mem[57][2] ),
    .A2(\mem[58][2] ),
    .A3(\mem[59][2] ),
    .S1(net533),
    .X(_0407_));
 sg13g2_and2_1 _3263_ (.A(net505),
    .B(_0407_),
    .X(_0408_));
 sg13g2_o21ai_1 _3264_ (.B1(net527),
    .Y(_0409_),
    .A1(_0406_),
    .A2(_0408_));
 sg13g2_nand2_1 _3265_ (.Y(_0410_),
    .A(net516),
    .B(\mem[52][2] ));
 sg13g2_a21oi_1 _3266_ (.A1(net577),
    .A2(\mem[53][2] ),
    .Y(_0411_),
    .B1(net535));
 sg13g2_nor2b_1 _3267_ (.A(net553),
    .B_N(\mem[54][2] ),
    .Y(_0412_));
 sg13g2_a21oi_1 _3268_ (.A1(net553),
    .A2(\mem[55][2] ),
    .Y(_0413_),
    .B1(_0412_));
 sg13g2_a221oi_1 _3269_ (.B2(net535),
    .C1(net507),
    .B1(_0413_),
    .A1(_0410_),
    .Y(_0414_),
    .A2(_0411_));
 sg13g2_mux4_1 _3270_ (.S0(net553),
    .A0(\mem[48][2] ),
    .A1(\mem[49][2] ),
    .A2(\mem[50][2] ),
    .A3(\mem[51][2] ),
    .S1(net535),
    .X(_0415_));
 sg13g2_and2_1 _3271_ (.A(net507),
    .B(_0415_),
    .X(_0416_));
 sg13g2_o21ai_1 _3272_ (.B1(net502),
    .Y(_0417_),
    .A1(_0414_),
    .A2(_0416_));
 sg13g2_nand3_1 _3273_ (.B(_0409_),
    .C(_0417_),
    .A(net524),
    .Y(_0418_));
 sg13g2_nand3_1 _3274_ (.B(_0401_),
    .C(_0418_),
    .A(net522),
    .Y(_0419_));
 sg13g2_nor2_1 _3275_ (.A(net565),
    .B(_2104_),
    .Y(_0420_));
 sg13g2_a21oi_1 _3276_ (.A1(net565),
    .A2(\mem[29][2] ),
    .Y(_0421_),
    .B1(_0420_));
 sg13g2_nand2_1 _3277_ (.Y(_0422_),
    .A(net520),
    .B(\mem[30][2] ));
 sg13g2_a21oi_1 _3278_ (.A1(net567),
    .A2(\mem[31][2] ),
    .Y(_0423_),
    .B1(net514));
 sg13g2_a221oi_1 _3279_ (.B2(_0423_),
    .C1(net510),
    .B1(_0422_),
    .A1(net514),
    .Y(_0424_),
    .A2(_0421_));
 sg13g2_mux4_1 _3280_ (.S0(net555),
    .A0(\mem[24][2] ),
    .A1(\mem[25][2] ),
    .A2(\mem[26][2] ),
    .A3(\mem[27][2] ),
    .S1(net536),
    .X(_0425_));
 sg13g2_a21o_1 _3281_ (.A2(_0425_),
    .A1(net511),
    .B1(_0424_),
    .X(_0426_));
 sg13g2_a21oi_1 _3282_ (.A1(net570),
    .A2(\mem[21][2] ),
    .Y(_0427_),
    .B1(net546));
 sg13g2_o21ai_1 _3283_ (.B1(_0427_),
    .Y(_0428_),
    .A1(net569),
    .A2(_2103_));
 sg13g2_nor2b_1 _3284_ (.A(net569),
    .B_N(\mem[22][2] ),
    .Y(_0429_));
 sg13g2_a21oi_1 _3285_ (.A1(net569),
    .A2(\mem[23][2] ),
    .Y(_0430_),
    .B1(_0429_));
 sg13g2_a21oi_1 _3286_ (.A1(net547),
    .A2(_0430_),
    .Y(_0431_),
    .B1(net512));
 sg13g2_mux4_1 _3287_ (.S0(net575),
    .A0(\mem[16][2] ),
    .A1(\mem[17][2] ),
    .A2(\mem[18][2] ),
    .A3(\mem[19][2] ),
    .S1(net548),
    .X(_0432_));
 sg13g2_a22oi_1 _3288_ (.Y(_0433_),
    .B1(_0432_),
    .B2(net513),
    .A2(_0431_),
    .A1(_0428_));
 sg13g2_o21ai_1 _3289_ (.B1(net525),
    .Y(_0434_),
    .A1(net529),
    .A2(_0433_));
 sg13g2_a21oi_1 _3290_ (.A1(net529),
    .A2(_0426_),
    .Y(_0435_),
    .B1(_0434_));
 sg13g2_nand2_1 _3291_ (.Y(_0436_),
    .A(net520),
    .B(\mem[12][2] ));
 sg13g2_a21oi_1 _3292_ (.A1(net565),
    .A2(\mem[13][2] ),
    .Y(_0437_),
    .B1(net543));
 sg13g2_nor2b_1 _3293_ (.A(net565),
    .B_N(\mem[14][2] ),
    .Y(_0438_));
 sg13g2_a21oi_1 _3294_ (.A1(net565),
    .A2(\mem[15][2] ),
    .Y(_0439_),
    .B1(_0438_));
 sg13g2_a221oi_1 _3295_ (.B2(net543),
    .C1(net510),
    .B1(_0439_),
    .A1(_0436_),
    .Y(_0440_),
    .A2(_0437_));
 sg13g2_mux4_1 _3296_ (.S0(net555),
    .A0(\mem[8][2] ),
    .A1(\mem[9][2] ),
    .A2(\mem[10][2] ),
    .A3(\mem[11][2] ),
    .S1(net536),
    .X(_0441_));
 sg13g2_and2_1 _3297_ (.A(net511),
    .B(_0441_),
    .X(_0442_));
 sg13g2_o21ai_1 _3298_ (.B1(net530),
    .Y(_0443_),
    .A1(_0440_),
    .A2(_0442_));
 sg13g2_nand2_1 _3299_ (.Y(_0444_),
    .A(net521),
    .B(\mem[4][2] ));
 sg13g2_a21oi_1 _3300_ (.A1(net572),
    .A2(\mem[5][2] ),
    .Y(_0445_),
    .B1(net548));
 sg13g2_nor2_1 _3301_ (.A(net571),
    .B(_2102_),
    .Y(_0446_));
 sg13g2_a21oi_1 _3302_ (.A1(net571),
    .A2(\mem[7][2] ),
    .Y(_0447_),
    .B1(_0446_));
 sg13g2_a221oi_1 _3303_ (.B2(net547),
    .C1(net512),
    .B1(_0447_),
    .A1(_0444_),
    .Y(_0448_),
    .A2(_0445_));
 sg13g2_nand2_1 _3304_ (.Y(_0449_),
    .A(\mem[0][2] ),
    .B(net519));
 sg13g2_a21oi_1 _3305_ (.A1(net574),
    .A2(\mem[1][2] ),
    .Y(_0450_),
    .B1(net546));
 sg13g2_nor2b_1 _3306_ (.A(net576),
    .B_N(\mem[2][2] ),
    .Y(_0451_));
 sg13g2_a21oi_1 _3307_ (.A1(net574),
    .A2(\mem[3][2] ),
    .Y(_0452_),
    .B1(_0451_));
 sg13g2_a221oi_1 _3308_ (.B2(net546),
    .C1(net532),
    .B1(_0452_),
    .A1(_0449_),
    .Y(_0453_),
    .A2(_0450_));
 sg13g2_o21ai_1 _3309_ (.B1(net504),
    .Y(_0454_),
    .A1(_0448_),
    .A2(_0453_));
 sg13g2_nand3b_1 _3310_ (.B(_0443_),
    .C(_0454_),
    .Y(_0455_),
    .A_N(net525));
 sg13g2_nand2b_1 _3311_ (.Y(_0456_),
    .B(_0455_),
    .A_N(net523));
 sg13g2_o21ai_1 _3312_ (.B1(_0419_),
    .Y(uio_out[2]),
    .A1(_0435_),
    .A2(_0456_));
 sg13g2_nand2_1 _3313_ (.Y(_0457_),
    .A(net515),
    .B(\mem[44][3] ));
 sg13g2_a21oi_1 _3314_ (.A1(net556),
    .A2(\mem[45][3] ),
    .Y(_0458_),
    .B1(net537));
 sg13g2_nor2b_1 _3315_ (.A(net556),
    .B_N(\mem[46][3] ),
    .Y(_0459_));
 sg13g2_a21oi_1 _3316_ (.A1(net556),
    .A2(\mem[47][3] ),
    .Y(_0460_),
    .B1(_0459_));
 sg13g2_a221oi_1 _3317_ (.B2(net537),
    .C1(net506),
    .B1(_0460_),
    .A1(_0457_),
    .Y(_0461_),
    .A2(_0458_));
 sg13g2_mux4_1 _3318_ (.S0(net558),
    .A0(\mem[40][3] ),
    .A1(\mem[41][3] ),
    .A2(\mem[42][3] ),
    .A3(\mem[43][3] ),
    .S1(net539),
    .X(_0462_));
 sg13g2_and2_1 _3319_ (.A(net506),
    .B(_0462_),
    .X(_0463_));
 sg13g2_o21ai_1 _3320_ (.B1(net527),
    .Y(_0464_),
    .A1(_0461_),
    .A2(_0463_));
 sg13g2_nand2_1 _3321_ (.Y(_0465_),
    .A(net516),
    .B(\mem[36][3] ));
 sg13g2_a21oi_1 _3322_ (.A1(net558),
    .A2(\mem[37][3] ),
    .Y(_0466_),
    .B1(net539));
 sg13g2_nor2b_1 _3323_ (.A(net559),
    .B_N(\mem[38][3] ),
    .Y(_0467_));
 sg13g2_a21oi_1 _3324_ (.A1(net559),
    .A2(\mem[39][3] ),
    .Y(_0468_),
    .B1(_0467_));
 sg13g2_a221oi_1 _3325_ (.B2(net540),
    .C1(net508),
    .B1(_0468_),
    .A1(_0465_),
    .Y(_0469_),
    .A2(_0466_));
 sg13g2_nand2_1 _3326_ (.Y(_0470_),
    .A(net517),
    .B(\mem[32][3] ));
 sg13g2_a21oi_1 _3327_ (.A1(uo_out[3]),
    .A2(net561),
    .Y(_0471_),
    .B1(net541));
 sg13g2_nand2_1 _3328_ (.Y(_0472_),
    .A(uo_out[7]),
    .B(net517));
 sg13g2_a21oi_1 _3329_ (.A1(net562),
    .A2(\mem[35][3] ),
    .Y(_0473_),
    .B1(net514));
 sg13g2_a221oi_1 _3330_ (.B2(_0473_),
    .C1(net531),
    .B1(_0472_),
    .A1(_0470_),
    .Y(_0474_),
    .A2(_0471_));
 sg13g2_o21ai_1 _3331_ (.B1(net503),
    .Y(_0475_),
    .A1(_0469_),
    .A2(_0474_));
 sg13g2_nand3b_1 _3332_ (.B(_0464_),
    .C(_0475_),
    .Y(_0476_),
    .A_N(net524));
 sg13g2_nand2_1 _3333_ (.Y(_0477_),
    .A(net518),
    .B(\mem[60][3] ));
 sg13g2_a21oi_1 _3334_ (.A1(net552),
    .A2(\mem[61][3] ),
    .Y(_0478_),
    .B1(net533));
 sg13g2_nor2b_1 _3335_ (.A(net551),
    .B_N(\mem[62][3] ),
    .Y(_0479_));
 sg13g2_a21oi_1 _3336_ (.A1(net551),
    .A2(\mem[63][3] ),
    .Y(_0480_),
    .B1(_0479_));
 sg13g2_a221oi_1 _3337_ (.B2(net533),
    .C1(net505),
    .B1(_0480_),
    .A1(_0477_),
    .Y(_0481_),
    .A2(_0478_));
 sg13g2_mux4_1 _3338_ (.S0(net551),
    .A0(\mem[56][3] ),
    .A1(\mem[57][3] ),
    .A2(\mem[58][3] ),
    .A3(\mem[59][3] ),
    .S1(net533),
    .X(_0482_));
 sg13g2_and2_1 _3339_ (.A(net505),
    .B(_0482_),
    .X(_0483_));
 sg13g2_o21ai_1 _3340_ (.B1(net527),
    .Y(_0484_),
    .A1(_0481_),
    .A2(_0483_));
 sg13g2_nand2_1 _3341_ (.Y(_0485_),
    .A(net516),
    .B(\mem[52][3] ));
 sg13g2_a21oi_1 _3342_ (.A1(net555),
    .A2(\mem[53][3] ),
    .Y(_0486_),
    .B1(net535));
 sg13g2_nor2b_1 _3343_ (.A(net553),
    .B_N(\mem[54][3] ),
    .Y(_0487_));
 sg13g2_a21oi_1 _3344_ (.A1(net553),
    .A2(\mem[55][3] ),
    .Y(_0488_),
    .B1(_0487_));
 sg13g2_a221oi_1 _3345_ (.B2(net535),
    .C1(net509),
    .B1(_0488_),
    .A1(_0485_),
    .Y(_0489_),
    .A2(_0486_));
 sg13g2_mux4_1 _3346_ (.S0(net553),
    .A0(\mem[48][3] ),
    .A1(\mem[49][3] ),
    .A2(\mem[50][3] ),
    .A3(\mem[51][3] ),
    .S1(net535),
    .X(_0490_));
 sg13g2_and2_1 _3347_ (.A(net505),
    .B(_0490_),
    .X(_0491_));
 sg13g2_o21ai_1 _3348_ (.B1(net502),
    .Y(_0492_),
    .A1(_0489_),
    .A2(_0491_));
 sg13g2_nand3_1 _3349_ (.B(_0484_),
    .C(_0492_),
    .A(net524),
    .Y(_0493_));
 sg13g2_nand3_1 _3350_ (.B(_0476_),
    .C(_0493_),
    .A(net522),
    .Y(_0494_));
 sg13g2_nor2_1 _3351_ (.A(net564),
    .B(_2105_),
    .Y(_0495_));
 sg13g2_a21oi_1 _3352_ (.A1(net564),
    .A2(\mem[29][3] ),
    .Y(_0496_),
    .B1(_0495_));
 sg13g2_nand2_1 _3353_ (.Y(_0497_),
    .A(net520),
    .B(\mem[30][3] ));
 sg13g2_a21oi_1 _3354_ (.A1(net567),
    .A2(\mem[31][3] ),
    .Y(_0498_),
    .B1(net514));
 sg13g2_a221oi_1 _3355_ (.B2(_0498_),
    .C1(net510),
    .B1(_0497_),
    .A1(net514),
    .Y(_0499_),
    .A2(_0496_));
 sg13g2_mux4_1 _3356_ (.S0(net555),
    .A0(\mem[24][3] ),
    .A1(\mem[25][3] ),
    .A2(\mem[26][3] ),
    .A3(\mem[27][3] ),
    .S1(net536),
    .X(_0500_));
 sg13g2_a21o_1 _3357_ (.A2(_0500_),
    .A1(net511),
    .B1(_0499_),
    .X(_0501_));
 sg13g2_nand2_1 _3358_ (.Y(_0502_),
    .A(net519),
    .B(\mem[20][3] ));
 sg13g2_a21oi_1 _3359_ (.A1(net570),
    .A2(\mem[21][3] ),
    .Y(_0503_),
    .B1(net547));
 sg13g2_nor2b_1 _3360_ (.A(net569),
    .B_N(\mem[22][3] ),
    .Y(_0504_));
 sg13g2_a21oi_1 _3361_ (.A1(net569),
    .A2(\mem[23][3] ),
    .Y(_0505_),
    .B1(_0504_));
 sg13g2_a221oi_1 _3362_ (.B2(net546),
    .C1(net512),
    .B1(_0505_),
    .A1(_0502_),
    .Y(_0506_),
    .A2(_0503_));
 sg13g2_mux4_1 _3363_ (.S0(net575),
    .A0(\mem[16][3] ),
    .A1(\mem[17][3] ),
    .A2(\mem[18][3] ),
    .A3(\mem[19][3] ),
    .S1(net549),
    .X(_0507_));
 sg13g2_a21oi_1 _3364_ (.A1(net513),
    .A2(_0507_),
    .Y(_0508_),
    .B1(_0506_));
 sg13g2_o21ai_1 _3365_ (.B1(net525),
    .Y(_0509_),
    .A1(net529),
    .A2(_0508_));
 sg13g2_a21oi_1 _3366_ (.A1(net529),
    .A2(_0501_),
    .Y(_0510_),
    .B1(_0509_));
 sg13g2_nand2_1 _3367_ (.Y(_0511_),
    .A(net520),
    .B(\mem[12][3] ));
 sg13g2_a21oi_1 _3368_ (.A1(net566),
    .A2(\mem[13][3] ),
    .Y(_0512_),
    .B1(net543));
 sg13g2_nor2b_1 _3369_ (.A(net565),
    .B_N(\mem[14][3] ),
    .Y(_0513_));
 sg13g2_a21oi_1 _3370_ (.A1(net565),
    .A2(\mem[15][3] ),
    .Y(_0514_),
    .B1(_0513_));
 sg13g2_a221oi_1 _3371_ (.B2(net543),
    .C1(net510),
    .B1(_0514_),
    .A1(_0511_),
    .Y(_0515_),
    .A2(_0512_));
 sg13g2_mux4_1 _3372_ (.S0(net555),
    .A0(\mem[8][3] ),
    .A1(\mem[9][3] ),
    .A2(\mem[10][3] ),
    .A3(\mem[11][3] ),
    .S1(net536),
    .X(_0516_));
 sg13g2_and2_1 _3373_ (.A(net511),
    .B(_0516_),
    .X(_0517_));
 sg13g2_o21ai_1 _3374_ (.B1(net530),
    .Y(_0518_),
    .A1(_0515_),
    .A2(_0517_));
 sg13g2_nand2_1 _3375_ (.Y(_0519_),
    .A(net519),
    .B(\mem[4][3] ));
 sg13g2_a21oi_1 _3376_ (.A1(net572),
    .A2(\mem[5][3] ),
    .Y(_0520_),
    .B1(net548));
 sg13g2_nor2b_1 _3377_ (.A(net571),
    .B_N(\mem[6][3] ),
    .Y(_0521_));
 sg13g2_a21oi_1 _3378_ (.A1(net571),
    .A2(\mem[7][3] ),
    .Y(_0522_),
    .B1(_0521_));
 sg13g2_a221oi_1 _3379_ (.B2(net547),
    .C1(net512),
    .B1(_0522_),
    .A1(_0519_),
    .Y(_0523_),
    .A2(_0520_));
 sg13g2_nand2_1 _3380_ (.Y(_0524_),
    .A(\mem[0][3] ),
    .B(net519));
 sg13g2_a21oi_1 _3381_ (.A1(net574),
    .A2(\mem[1][3] ),
    .Y(_0525_),
    .B1(net548));
 sg13g2_nor2b_1 _3382_ (.A(net574),
    .B_N(\mem[2][3] ),
    .Y(_0526_));
 sg13g2_a21oi_1 _3383_ (.A1(net574),
    .A2(\mem[3][3] ),
    .Y(_0527_),
    .B1(_0526_));
 sg13g2_a221oi_1 _3384_ (.B2(net546),
    .C1(net532),
    .B1(_0527_),
    .A1(_0524_),
    .Y(_0528_),
    .A2(_0525_));
 sg13g2_o21ai_1 _3385_ (.B1(net504),
    .Y(_0529_),
    .A1(_0523_),
    .A2(_0528_));
 sg13g2_nand3b_1 _3386_ (.B(_0518_),
    .C(_0529_),
    .Y(_0530_),
    .A_N(net525));
 sg13g2_nand2b_1 _3387_ (.Y(_0531_),
    .B(_0530_),
    .A_N(net523));
 sg13g2_o21ai_1 _3388_ (.B1(_0494_),
    .Y(uio_out[3]),
    .A1(_0510_),
    .A2(_0531_));
 sg13g2_nand2_1 _3389_ (.Y(_0532_),
    .A(uio_out[5]),
    .B(uio_out[4]));
 sg13g2_and4_2 _3390_ (.A(net578),
    .B(_2091_),
    .C(net1),
    .D(_0532_),
    .X(_0533_));
 sg13g2_nand4_1 _3391_ (.B(_2091_),
    .C(net1),
    .A(net578),
    .Y(_0534_),
    .D(_0532_));
 sg13g2_nand2_2 _3392_ (.Y(_0535_),
    .A(net531),
    .B(net488));
 sg13g2_nor2_1 _3393_ (.A(net538),
    .B(_0535_),
    .Y(_0536_));
 sg13g2_nor3_2 _3394_ (.A(net518),
    .B(net534),
    .C(_0535_),
    .Y(_0537_));
 sg13g2_nand2_2 _3395_ (.Y(_0538_),
    .A(net557),
    .B(_0536_));
 sg13g2_nor3_2 _3396_ (.A(net525),
    .B(net523),
    .C(_0534_),
    .Y(_0539_));
 sg13g2_and2_2 _3397_ (.A(net530),
    .B(_0539_),
    .X(_0540_));
 sg13g2_nand2_2 _3398_ (.Y(_0541_),
    .A(net530),
    .B(_0539_));
 sg13g2_nand2_2 _3399_ (.Y(_0542_),
    .A(_0537_),
    .B(_0540_));
 sg13g2_and2_1 _3400_ (.A(\products[6][0] ),
    .B(\products[5][0] ),
    .X(_0543_));
 sg13g2_xor2_1 _3401_ (.B(\products[5][0] ),
    .A(\products[6][0] ),
    .X(_0544_));
 sg13g2_xnor2_1 _3402_ (.Y(_0545_),
    .A(\products[7][0] ),
    .B(_0544_));
 sg13g2_and2_1 _3403_ (.A(\prev_acc[0] ),
    .B(\products[0][0] ),
    .X(_0546_));
 sg13g2_xor2_1 _3404_ (.B(\products[0][0] ),
    .A(\prev_acc[0] ),
    .X(_0547_));
 sg13g2_xnor2_1 _3405_ (.Y(_0548_),
    .A(\products[1][0] ),
    .B(_0547_));
 sg13g2_and2_1 _3406_ (.A(\products[3][0] ),
    .B(\products[2][0] ),
    .X(_0549_));
 sg13g2_xor2_1 _3407_ (.B(\products[2][0] ),
    .A(\products[3][0] ),
    .X(_0550_));
 sg13g2_xnor2_1 _3408_ (.Y(_0551_),
    .A(\products[4][0] ),
    .B(_0550_));
 sg13g2_nor2_1 _3409_ (.A(_0548_),
    .B(_0551_),
    .Y(_0552_));
 sg13g2_xor2_1 _3410_ (.B(_0551_),
    .A(_0548_),
    .X(_0553_));
 sg13g2_nand2b_1 _3411_ (.Y(_0554_),
    .B(_0553_),
    .A_N(_0545_));
 sg13g2_xnor2_1 _3412_ (.Y(_0555_),
    .A(_0545_),
    .B(_0553_));
 sg13g2_and2_1 _3413_ (.A(\products[9][0] ),
    .B(\products[8][0] ),
    .X(_0556_));
 sg13g2_xor2_1 _3414_ (.B(\products[8][0] ),
    .A(\products[9][0] ),
    .X(_0557_));
 sg13g2_xnor2_1 _3415_ (.Y(_0558_),
    .A(\products[10][0] ),
    .B(_0557_));
 sg13g2_and2_1 _3416_ (.A(\products[12][0] ),
    .B(\products[11][0] ),
    .X(_0559_));
 sg13g2_xor2_1 _3417_ (.B(\products[11][0] ),
    .A(\products[12][0] ),
    .X(_0560_));
 sg13g2_xnor2_1 _3418_ (.Y(_0561_),
    .A(\products[13][0] ),
    .B(_0560_));
 sg13g2_nor2_1 _3419_ (.A(_0558_),
    .B(_0561_),
    .Y(_0562_));
 sg13g2_xor2_1 _3420_ (.B(_0561_),
    .A(_0558_),
    .X(_0563_));
 sg13g2_nand2_1 _3421_ (.Y(_0564_),
    .A(_0555_),
    .B(_0563_));
 sg13g2_xnor2_1 _3422_ (.Y(_0565_),
    .A(_0555_),
    .B(_0563_));
 sg13g2_nand2_1 _3423_ (.Y(_0566_),
    .A(\products[14][0] ),
    .B(\products[15][0] ));
 sg13g2_xnor2_1 _3424_ (.Y(_0567_),
    .A(\products[14][0] ),
    .B(\products[15][0] ));
 sg13g2_nor2_1 _3425_ (.A(_0565_),
    .B(_0567_),
    .Y(_0568_));
 sg13g2_a21o_1 _3426_ (.A2(_0567_),
    .A1(_0565_),
    .B1(net487),
    .X(_0569_));
 sg13g2_nand2_1 _3427_ (.Y(_0570_),
    .A(net3),
    .B(net487));
 sg13g2_o21ai_1 _3428_ (.B1(_0570_),
    .Y(_0571_),
    .A1(_0568_),
    .A2(_0569_));
 sg13g2_mux2_1 _3429_ (.A0(net479),
    .A1(net794),
    .S(_0542_),
    .X(_0001_));
 sg13g2_a21oi_1 _3430_ (.A1(\products[13][0] ),
    .A2(_0560_),
    .Y(_0572_),
    .B1(_0559_));
 sg13g2_nor2b_1 _3431_ (.A(_0572_),
    .B_N(\products[14][1] ),
    .Y(_0573_));
 sg13g2_xnor2_1 _3432_ (.Y(_0574_),
    .A(\products[14][1] ),
    .B(_0572_));
 sg13g2_xnor2_1 _3433_ (.Y(_0575_),
    .A(\products[15][1] ),
    .B(_0574_));
 sg13g2_nor2_1 _3434_ (.A(_0566_),
    .B(_0575_),
    .Y(_0576_));
 sg13g2_xor2_1 _3435_ (.B(_0575_),
    .A(_0566_),
    .X(_0577_));
 sg13g2_and2_1 _3436_ (.A(\products[12][1] ),
    .B(\products[11][1] ),
    .X(_0578_));
 sg13g2_xor2_1 _3437_ (.B(\products[11][1] ),
    .A(\products[12][1] ),
    .X(_0579_));
 sg13g2_xnor2_1 _3438_ (.Y(_0580_),
    .A(\products[13][1] ),
    .B(_0579_));
 sg13g2_inv_1 _3439_ (.Y(_0581_),
    .A(_0580_));
 sg13g2_a21oi_1 _3440_ (.A1(\products[10][0] ),
    .A2(_0557_),
    .Y(_0582_),
    .B1(_0556_));
 sg13g2_and2_1 _3441_ (.A(\products[9][1] ),
    .B(\products[8][1] ),
    .X(_0583_));
 sg13g2_xor2_1 _3442_ (.B(\products[8][1] ),
    .A(\products[9][1] ),
    .X(_0584_));
 sg13g2_xnor2_1 _3443_ (.Y(_0585_),
    .A(\products[10][1] ),
    .B(_0584_));
 sg13g2_nor2_1 _3444_ (.A(_0582_),
    .B(_0585_),
    .Y(_0586_));
 sg13g2_xor2_1 _3445_ (.B(_0585_),
    .A(_0582_),
    .X(_0587_));
 sg13g2_xnor2_1 _3446_ (.Y(_0588_),
    .A(_0580_),
    .B(_0587_));
 sg13g2_nand2_1 _3447_ (.Y(_0589_),
    .A(_0562_),
    .B(_0588_));
 sg13g2_xnor2_1 _3448_ (.Y(_0590_),
    .A(_0562_),
    .B(_0588_));
 sg13g2_a21oi_1 _3449_ (.A1(\products[7][0] ),
    .A2(_0544_),
    .Y(_0591_),
    .B1(_0543_));
 sg13g2_inv_1 _3450_ (.Y(_0592_),
    .A(_0591_));
 sg13g2_a21oi_2 _3451_ (.B1(_0549_),
    .Y(_0593_),
    .A2(_0550_),
    .A1(\products[4][0] ));
 sg13g2_and2_1 _3452_ (.A(\products[6][1] ),
    .B(\products[5][1] ),
    .X(_0594_));
 sg13g2_xor2_1 _3453_ (.B(\products[5][1] ),
    .A(\products[6][1] ),
    .X(_0595_));
 sg13g2_xnor2_1 _3454_ (.Y(_0596_),
    .A(\products[7][1] ),
    .B(_0595_));
 sg13g2_nor2_1 _3455_ (.A(_0593_),
    .B(_0596_),
    .Y(_0597_));
 sg13g2_xor2_1 _3456_ (.B(_0596_),
    .A(_0593_),
    .X(_0598_));
 sg13g2_xnor2_1 _3457_ (.Y(_0599_),
    .A(_0591_),
    .B(_0598_));
 sg13g2_inv_1 _3458_ (.Y(_0600_),
    .A(_0599_));
 sg13g2_and2_1 _3459_ (.A(\products[3][1] ),
    .B(\products[2][1] ),
    .X(_0601_));
 sg13g2_xor2_1 _3460_ (.B(\products[2][1] ),
    .A(\products[3][1] ),
    .X(_0602_));
 sg13g2_xor2_1 _3461_ (.B(_0602_),
    .A(\products[4][1] ),
    .X(_0603_));
 sg13g2_a21oi_1 _3462_ (.A1(\products[1][0] ),
    .A2(_0547_),
    .Y(_0604_),
    .B1(_0546_));
 sg13g2_and2_1 _3463_ (.A(\prev_acc[1] ),
    .B(\products[0][1] ),
    .X(_0605_));
 sg13g2_xor2_1 _3464_ (.B(\products[0][1] ),
    .A(\prev_acc[1] ),
    .X(_0606_));
 sg13g2_xnor2_1 _3465_ (.Y(_0607_),
    .A(\products[1][1] ),
    .B(_0606_));
 sg13g2_nor2_1 _3466_ (.A(_0604_),
    .B(_0607_),
    .Y(_0608_));
 sg13g2_xor2_1 _3467_ (.B(_0607_),
    .A(_0604_),
    .X(_0609_));
 sg13g2_xor2_1 _3468_ (.B(_0609_),
    .A(_0603_),
    .X(_0610_));
 sg13g2_nand2_1 _3469_ (.Y(_0611_),
    .A(_0552_),
    .B(_0610_));
 sg13g2_xnor2_1 _3470_ (.Y(_0612_),
    .A(_0552_),
    .B(_0610_));
 sg13g2_xnor2_1 _3471_ (.Y(_0613_),
    .A(_0600_),
    .B(_0612_));
 sg13g2_or2_1 _3472_ (.X(_0614_),
    .B(_0613_),
    .A(_0554_));
 sg13g2_xnor2_1 _3473_ (.Y(_0615_),
    .A(_0554_),
    .B(_0613_));
 sg13g2_xnor2_1 _3474_ (.Y(_0616_),
    .A(_0590_),
    .B(_0615_));
 sg13g2_nor2_1 _3475_ (.A(_0564_),
    .B(_0616_),
    .Y(_0617_));
 sg13g2_xor2_1 _3476_ (.B(_0616_),
    .A(_0564_),
    .X(_0618_));
 sg13g2_xor2_1 _3477_ (.B(_0618_),
    .A(_0577_),
    .X(_0619_));
 sg13g2_nand2_1 _3478_ (.Y(_0620_),
    .A(_0568_),
    .B(_0619_));
 sg13g2_o21ai_1 _3479_ (.B1(_0534_),
    .Y(_0621_),
    .A1(_0568_),
    .A2(_0619_));
 sg13g2_nor2b_1 _3480_ (.A(_0621_),
    .B_N(_0620_),
    .Y(_0622_));
 sg13g2_a21o_1 _3481_ (.A2(net487),
    .A1(net4),
    .B1(_0622_),
    .X(_0623_));
 sg13g2_mux2_1 _3482_ (.A0(net467),
    .A1(net842),
    .S(_0542_),
    .X(_0002_));
 sg13g2_a21oi_1 _3483_ (.A1(_0577_),
    .A2(_0618_),
    .Y(_0624_),
    .B1(_0617_));
 sg13g2_a21o_1 _3484_ (.A2(_0574_),
    .A1(\products[15][1] ),
    .B1(_0573_),
    .X(_0625_));
 sg13g2_a21oi_2 _3485_ (.B1(_0578_),
    .Y(_0626_),
    .A2(_0579_),
    .A1(\products[13][1] ));
 sg13g2_nor2b_1 _3486_ (.A(_0626_),
    .B_N(\products[14][2] ),
    .Y(_0627_));
 sg13g2_xnor2_1 _3487_ (.Y(_0628_),
    .A(\products[14][2] ),
    .B(_0626_));
 sg13g2_xnor2_1 _3488_ (.Y(_0629_),
    .A(\products[15][2] ),
    .B(_0628_));
 sg13g2_xor2_1 _3489_ (.B(_0629_),
    .A(_0589_),
    .X(_0630_));
 sg13g2_nand2_1 _3490_ (.Y(_0631_),
    .A(_0625_),
    .B(_0630_));
 sg13g2_xnor2_1 _3491_ (.Y(_0632_),
    .A(_0625_),
    .B(_0630_));
 sg13g2_o21ai_1 _3492_ (.B1(_0614_),
    .Y(_0633_),
    .A1(_0590_),
    .A2(_0615_));
 sg13g2_a21oi_2 _3493_ (.B1(_0586_),
    .Y(_0634_),
    .A2(_0587_),
    .A1(_0581_));
 sg13g2_a21oi_2 _3494_ (.B1(_0597_),
    .Y(_0635_),
    .A2(_0598_),
    .A1(_0592_));
 sg13g2_and2_1 _3495_ (.A(\products[12][2] ),
    .B(\products[11][2] ),
    .X(_0636_));
 sg13g2_xor2_1 _3496_ (.B(\products[11][2] ),
    .A(\products[12][2] ),
    .X(_0637_));
 sg13g2_xnor2_1 _3497_ (.Y(_0638_),
    .A(\products[13][2] ),
    .B(_0637_));
 sg13g2_inv_1 _3498_ (.Y(_0639_),
    .A(_0638_));
 sg13g2_a21oi_1 _3499_ (.A1(\products[10][1] ),
    .A2(_0584_),
    .Y(_0640_),
    .B1(_0583_));
 sg13g2_and2_1 _3500_ (.A(\products[9][2] ),
    .B(\products[8][2] ),
    .X(_0641_));
 sg13g2_xor2_1 _3501_ (.B(\products[8][2] ),
    .A(\products[9][2] ),
    .X(_0642_));
 sg13g2_xnor2_1 _3502_ (.Y(_0643_),
    .A(\products[10][2] ),
    .B(_0642_));
 sg13g2_nor2_1 _3503_ (.A(_0640_),
    .B(_0643_),
    .Y(_0644_));
 sg13g2_xor2_1 _3504_ (.B(_0643_),
    .A(_0640_),
    .X(_0645_));
 sg13g2_xnor2_1 _3505_ (.Y(_0646_),
    .A(_0638_),
    .B(_0645_));
 sg13g2_nor2b_1 _3506_ (.A(_0635_),
    .B_N(_0646_),
    .Y(_0647_));
 sg13g2_xnor2_1 _3507_ (.Y(_0648_),
    .A(_0635_),
    .B(_0646_));
 sg13g2_nor2b_1 _3508_ (.A(_0634_),
    .B_N(_0648_),
    .Y(_0649_));
 sg13g2_xnor2_1 _3509_ (.Y(_0650_),
    .A(_0634_),
    .B(_0648_));
 sg13g2_inv_1 _3510_ (.Y(_0651_),
    .A(_0650_));
 sg13g2_o21ai_1 _3511_ (.B1(_0611_),
    .Y(_0652_),
    .A1(_0600_),
    .A2(_0612_));
 sg13g2_a21o_1 _3512_ (.A2(_0595_),
    .A1(\products[7][1] ),
    .B1(_0594_),
    .X(_0653_));
 sg13g2_a21oi_2 _3513_ (.B1(_0601_),
    .Y(_0654_),
    .A2(_0602_),
    .A1(\products[4][1] ));
 sg13g2_and2_1 _3514_ (.A(\products[6][2] ),
    .B(\products[5][2] ),
    .X(_0655_));
 sg13g2_xor2_1 _3515_ (.B(\products[5][2] ),
    .A(\products[6][2] ),
    .X(_0656_));
 sg13g2_xnor2_1 _3516_ (.Y(_0657_),
    .A(\products[7][2] ),
    .B(_0656_));
 sg13g2_nor2_1 _3517_ (.A(_0654_),
    .B(_0657_),
    .Y(_0658_));
 sg13g2_xor2_1 _3518_ (.B(_0657_),
    .A(_0654_),
    .X(_0659_));
 sg13g2_xor2_1 _3519_ (.B(_0659_),
    .A(_0653_),
    .X(_0660_));
 sg13g2_a21oi_1 _3520_ (.A1(_0603_),
    .A2(_0609_),
    .Y(_0661_),
    .B1(_0608_));
 sg13g2_and2_1 _3521_ (.A(\products[3][2] ),
    .B(\products[2][2] ),
    .X(_0662_));
 sg13g2_xor2_1 _3522_ (.B(\products[2][2] ),
    .A(\products[3][2] ),
    .X(_0663_));
 sg13g2_xor2_1 _3523_ (.B(_0663_),
    .A(\products[4][2] ),
    .X(_0664_));
 sg13g2_a21oi_1 _3524_ (.A1(\products[1][1] ),
    .A2(_0606_),
    .Y(_0665_),
    .B1(_0605_));
 sg13g2_and2_1 _3525_ (.A(\prev_acc[2] ),
    .B(\products[0][2] ),
    .X(_0666_));
 sg13g2_xor2_1 _3526_ (.B(\products[0][2] ),
    .A(\prev_acc[2] ),
    .X(_0667_));
 sg13g2_xnor2_1 _3527_ (.Y(_0668_),
    .A(\products[1][2] ),
    .B(_0667_));
 sg13g2_nor2_1 _3528_ (.A(_0665_),
    .B(_0668_),
    .Y(_0669_));
 sg13g2_xor2_1 _3529_ (.B(_0668_),
    .A(_0665_),
    .X(_0670_));
 sg13g2_xor2_1 _3530_ (.B(_0670_),
    .A(_0664_),
    .X(_0671_));
 sg13g2_nor2b_1 _3531_ (.A(_0661_),
    .B_N(_0671_),
    .Y(_0672_));
 sg13g2_xnor2_1 _3532_ (.Y(_0673_),
    .A(_0661_),
    .B(_0671_));
 sg13g2_xnor2_1 _3533_ (.Y(_0674_),
    .A(_0660_),
    .B(_0673_));
 sg13g2_nand2b_1 _3534_ (.Y(_0675_),
    .B(_0652_),
    .A_N(_0674_));
 sg13g2_xor2_1 _3535_ (.B(_0674_),
    .A(_0652_),
    .X(_0676_));
 sg13g2_xnor2_1 _3536_ (.Y(_0677_),
    .A(_0651_),
    .B(_0676_));
 sg13g2_nand2b_1 _3537_ (.Y(_0678_),
    .B(_0633_),
    .A_N(_0677_));
 sg13g2_xor2_1 _3538_ (.B(_0677_),
    .A(_0633_),
    .X(_0679_));
 sg13g2_xnor2_1 _3539_ (.Y(_0680_),
    .A(_0632_),
    .B(_0679_));
 sg13g2_nor2_1 _3540_ (.A(_0624_),
    .B(_0680_),
    .Y(_0681_));
 sg13g2_xor2_1 _3541_ (.B(_0680_),
    .A(_0624_),
    .X(_0682_));
 sg13g2_xnor2_1 _3542_ (.Y(_0683_),
    .A(_0576_),
    .B(_0682_));
 sg13g2_nor2_2 _3543_ (.A(_0620_),
    .B(_0683_),
    .Y(_0684_));
 sg13g2_nand2_1 _3544_ (.Y(_0685_),
    .A(net5),
    .B(net487));
 sg13g2_a21o_1 _3545_ (.A2(_0683_),
    .A1(_0620_),
    .B1(net487),
    .X(_0686_));
 sg13g2_o21ai_1 _3546_ (.B1(_0685_),
    .Y(_0687_),
    .A1(_0684_),
    .A2(_0686_));
 sg13g2_mux2_1 _3547_ (.A0(net457),
    .A1(net843),
    .S(_0542_),
    .X(_0003_));
 sg13g2_nand2_1 _3548_ (.Y(_0688_),
    .A(net6),
    .B(net487));
 sg13g2_a21oi_1 _3549_ (.A1(_0576_),
    .A2(_0682_),
    .Y(_0689_),
    .B1(_0681_));
 sg13g2_o21ai_1 _3550_ (.B1(_0631_),
    .Y(_0690_),
    .A1(_0589_),
    .A2(_0629_));
 sg13g2_o21ai_1 _3551_ (.B1(_0678_),
    .Y(_0691_),
    .A1(_0632_),
    .A2(_0679_));
 sg13g2_a21oi_1 _3552_ (.A1(\products[15][2] ),
    .A2(_0628_),
    .Y(_0692_),
    .B1(_0627_));
 sg13g2_nor2_1 _3553_ (.A(_0647_),
    .B(_0649_),
    .Y(_0693_));
 sg13g2_a21oi_2 _3554_ (.B1(_0636_),
    .Y(_0694_),
    .A2(_0637_),
    .A1(\products[13][2] ));
 sg13g2_nor2b_1 _3555_ (.A(_0694_),
    .B_N(\products[14][3] ),
    .Y(_0695_));
 sg13g2_xnor2_1 _3556_ (.Y(_0696_),
    .A(\products[14][3] ),
    .B(_0694_));
 sg13g2_xnor2_1 _3557_ (.Y(_0697_),
    .A(\products[15][3] ),
    .B(_0696_));
 sg13g2_or2_1 _3558_ (.X(_0698_),
    .B(_0697_),
    .A(_0693_));
 sg13g2_xnor2_1 _3559_ (.Y(_0699_),
    .A(_0693_),
    .B(_0697_));
 sg13g2_xor2_1 _3560_ (.B(_0699_),
    .A(_0692_),
    .X(_0700_));
 sg13g2_o21ai_1 _3561_ (.B1(_0675_),
    .Y(_0701_),
    .A1(_0651_),
    .A2(_0676_));
 sg13g2_a21oi_2 _3562_ (.B1(_0644_),
    .Y(_0702_),
    .A2(_0645_),
    .A1(_0639_));
 sg13g2_a21oi_2 _3563_ (.B1(_0658_),
    .Y(_0703_),
    .A2(_0659_),
    .A1(_0653_));
 sg13g2_inv_1 _3564_ (.Y(_0704_),
    .A(_0703_));
 sg13g2_and2_1 _3565_ (.A(\products[12][3] ),
    .B(\products[11][3] ),
    .X(_0705_));
 sg13g2_xor2_1 _3566_ (.B(\products[11][3] ),
    .A(\products[12][3] ),
    .X(_0706_));
 sg13g2_xnor2_1 _3567_ (.Y(_0707_),
    .A(\products[13][3] ),
    .B(_0706_));
 sg13g2_inv_1 _3568_ (.Y(_0708_),
    .A(_0707_));
 sg13g2_a21oi_2 _3569_ (.B1(_0641_),
    .Y(_0709_),
    .A2(_0642_),
    .A1(\products[10][2] ));
 sg13g2_and2_1 _3570_ (.A(\products[9][3] ),
    .B(\products[8][3] ),
    .X(_0710_));
 sg13g2_xor2_1 _3571_ (.B(\products[8][3] ),
    .A(\products[9][3] ),
    .X(_0711_));
 sg13g2_xnor2_1 _3572_ (.Y(_0712_),
    .A(\products[10][3] ),
    .B(_0711_));
 sg13g2_nor2_1 _3573_ (.A(_0709_),
    .B(_0712_),
    .Y(_0713_));
 sg13g2_xor2_1 _3574_ (.B(_0712_),
    .A(_0709_),
    .X(_0714_));
 sg13g2_xnor2_1 _3575_ (.Y(_0715_),
    .A(_0707_),
    .B(_0714_));
 sg13g2_xnor2_1 _3576_ (.Y(_0716_),
    .A(_0703_),
    .B(_0715_));
 sg13g2_nor2b_1 _3577_ (.A(_0702_),
    .B_N(_0716_),
    .Y(_0717_));
 sg13g2_xnor2_1 _3578_ (.Y(_0718_),
    .A(_0702_),
    .B(_0716_));
 sg13g2_a21oi_1 _3579_ (.A1(_0660_),
    .A2(_0673_),
    .Y(_0719_),
    .B1(_0672_));
 sg13g2_a21o_1 _3580_ (.A2(_0656_),
    .A1(\products[7][2] ),
    .B1(_0655_),
    .X(_0720_));
 sg13g2_a21oi_2 _3581_ (.B1(_0662_),
    .Y(_0721_),
    .A2(_0663_),
    .A1(\products[4][2] ));
 sg13g2_and2_1 _3582_ (.A(\products[6][3] ),
    .B(\products[5][3] ),
    .X(_0722_));
 sg13g2_xor2_1 _3583_ (.B(\products[5][3] ),
    .A(\products[6][3] ),
    .X(_0723_));
 sg13g2_xnor2_1 _3584_ (.Y(_0724_),
    .A(\products[7][3] ),
    .B(_0723_));
 sg13g2_nor2_1 _3585_ (.A(_0721_),
    .B(_0724_),
    .Y(_0725_));
 sg13g2_xor2_1 _3586_ (.B(_0724_),
    .A(_0721_),
    .X(_0726_));
 sg13g2_xor2_1 _3587_ (.B(_0726_),
    .A(_0720_),
    .X(_0727_));
 sg13g2_a21oi_2 _3588_ (.B1(_0669_),
    .Y(_0728_),
    .A2(_0670_),
    .A1(_0664_));
 sg13g2_and2_1 _3589_ (.A(\products[3][3] ),
    .B(\products[2][3] ),
    .X(_0729_));
 sg13g2_xor2_1 _3590_ (.B(\products[2][3] ),
    .A(\products[3][3] ),
    .X(_0730_));
 sg13g2_xnor2_1 _3591_ (.Y(_0731_),
    .A(\products[4][3] ),
    .B(_0730_));
 sg13g2_inv_1 _3592_ (.Y(_0732_),
    .A(_0731_));
 sg13g2_a21oi_2 _3593_ (.B1(_0666_),
    .Y(_0733_),
    .A2(_0667_),
    .A1(\products[1][2] ));
 sg13g2_and2_1 _3594_ (.A(\prev_acc[3] ),
    .B(\products[0][3] ),
    .X(_0734_));
 sg13g2_xor2_1 _3595_ (.B(\products[0][3] ),
    .A(\prev_acc[3] ),
    .X(_0735_));
 sg13g2_xnor2_1 _3596_ (.Y(_0736_),
    .A(\products[1][3] ),
    .B(_0735_));
 sg13g2_nor2_2 _3597_ (.A(_0733_),
    .B(_0736_),
    .Y(_0737_));
 sg13g2_xor2_1 _3598_ (.B(_0736_),
    .A(_0733_),
    .X(_0738_));
 sg13g2_xnor2_1 _3599_ (.Y(_0739_),
    .A(_0732_),
    .B(_0738_));
 sg13g2_nor2_1 _3600_ (.A(_0728_),
    .B(_0739_),
    .Y(_0740_));
 sg13g2_xor2_1 _3601_ (.B(_0739_),
    .A(_0728_),
    .X(_0741_));
 sg13g2_xnor2_1 _3602_ (.Y(_0742_),
    .A(_0727_),
    .B(_0741_));
 sg13g2_nor2_1 _3603_ (.A(_0719_),
    .B(_0742_),
    .Y(_0743_));
 sg13g2_xor2_1 _3604_ (.B(_0742_),
    .A(_0719_),
    .X(_0744_));
 sg13g2_xnor2_1 _3605_ (.Y(_0745_),
    .A(_0718_),
    .B(_0744_));
 sg13g2_nor2b_1 _3606_ (.A(_0745_),
    .B_N(_0701_),
    .Y(_0746_));
 sg13g2_xnor2_1 _3607_ (.Y(_0747_),
    .A(_0701_),
    .B(_0745_));
 sg13g2_xnor2_1 _3608_ (.Y(_0748_),
    .A(_0700_),
    .B(_0747_));
 sg13g2_nor2b_1 _3609_ (.A(_0748_),
    .B_N(_0691_),
    .Y(_0749_));
 sg13g2_xnor2_1 _3610_ (.Y(_0750_),
    .A(_0691_),
    .B(_0748_));
 sg13g2_xnor2_1 _3611_ (.Y(_0751_),
    .A(_0690_),
    .B(_0750_));
 sg13g2_nor2_1 _3612_ (.A(_0689_),
    .B(_0751_),
    .Y(_0752_));
 sg13g2_xor2_1 _3613_ (.B(_0751_),
    .A(_0689_),
    .X(_0753_));
 sg13g2_xnor2_1 _3614_ (.Y(_0754_),
    .A(_0684_),
    .B(_0753_));
 sg13g2_o21ai_1 _3615_ (.B1(_0688_),
    .Y(_0755_),
    .A1(net487),
    .A2(_0754_));
 sg13g2_mux2_1 _3616_ (.A0(net449),
    .A1(net829),
    .S(_0542_),
    .X(_0004_));
 sg13g2_nand2_2 _3617_ (.Y(_0756_),
    .A(net542),
    .B(net488));
 sg13g2_nor2_1 _3618_ (.A(net531),
    .B(_0756_),
    .Y(_0757_));
 sg13g2_nor3_2 _3619_ (.A(net518),
    .B(net531),
    .C(_0756_),
    .Y(_0758_));
 sg13g2_nand2_2 _3620_ (.Y(_0759_),
    .A(net562),
    .B(_0757_));
 sg13g2_nand2_2 _3621_ (.Y(_0760_),
    .A(net526),
    .B(net488));
 sg13g2_nor2_2 _3622_ (.A(net522),
    .B(_0760_),
    .Y(_0761_));
 sg13g2_nor3_2 _3623_ (.A(net529),
    .B(net523),
    .C(_0760_),
    .Y(_0762_));
 sg13g2_nand2_2 _3624_ (.Y(_0763_),
    .A(net503),
    .B(_0761_));
 sg13g2_nand2_2 _3625_ (.Y(_0764_),
    .A(_0758_),
    .B(_0762_));
 sg13g2_mux2_1 _3626_ (.A0(net481),
    .A1(net818),
    .S(_0764_),
    .X(_0005_));
 sg13g2_mux2_1 _3627_ (.A0(net468),
    .A1(net701),
    .S(_0764_),
    .X(_0006_));
 sg13g2_mux2_1 _3628_ (.A0(net459),
    .A1(net808),
    .S(_0764_),
    .X(_0007_));
 sg13g2_mux2_1 _3629_ (.A0(net447),
    .A1(net821),
    .S(_0764_),
    .X(_0008_));
 sg13g2_nand2_2 _3630_ (.Y(_0765_),
    .A(_0540_),
    .B(_0758_));
 sg13g2_mux2_1 _3631_ (.A0(net474),
    .A1(net769),
    .S(_0765_),
    .X(_0009_));
 sg13g2_mux2_1 _3632_ (.A0(net462),
    .A1(net798),
    .S(_0765_),
    .X(_0010_));
 sg13g2_mux2_1 _3633_ (.A0(net452),
    .A1(net761),
    .S(_0765_),
    .X(_0011_));
 sg13g2_mux2_1 _3634_ (.A0(net443),
    .A1(net719),
    .S(_0765_),
    .X(_0012_));
 sg13g2_nor3_2 _3635_ (.A(net502),
    .B(net522),
    .C(_0760_),
    .Y(_0766_));
 sg13g2_nand2_2 _3636_ (.Y(_0767_),
    .A(net527),
    .B(_0761_));
 sg13g2_nand2_2 _3637_ (.Y(_0768_),
    .A(_0537_),
    .B(_0766_));
 sg13g2_mux2_1 _3638_ (.A0(net479),
    .A1(net716),
    .S(_0768_),
    .X(_0013_));
 sg13g2_mux2_1 _3639_ (.A0(net467),
    .A1(net835),
    .S(_0768_),
    .X(_0014_));
 sg13g2_mux2_1 _3640_ (.A0(net457),
    .A1(net838),
    .S(_0768_),
    .X(_0015_));
 sg13g2_mux2_1 _3641_ (.A0(net449),
    .A1(net810),
    .S(_0768_),
    .X(_0016_));
 sg13g2_nor3_2 _3642_ (.A(net555),
    .B(net531),
    .C(_0756_),
    .Y(_0769_));
 sg13g2_nand2_2 _3643_ (.Y(_0770_),
    .A(net516),
    .B(_0757_));
 sg13g2_nand2_2 _3644_ (.Y(_0771_),
    .A(_0540_),
    .B(_0769_));
 sg13g2_mux2_1 _3645_ (.A0(net472),
    .A1(net730),
    .S(_0771_),
    .X(_0017_));
 sg13g2_mux2_1 _3646_ (.A0(net461),
    .A1(net809),
    .S(_0771_),
    .X(_0018_));
 sg13g2_mux2_1 _3647_ (.A0(net451),
    .A1(net833),
    .S(_0771_),
    .X(_0019_));
 sg13g2_mux2_1 _3648_ (.A0(net450),
    .A1(net776),
    .S(_0771_),
    .X(_0020_));
 sg13g2_o21ai_1 _3649_ (.B1(net488),
    .Y(_0772_),
    .A1(net549),
    .A2(net532));
 sg13g2_o21ai_1 _3650_ (.B1(_0772_),
    .Y(_0773_),
    .A1(net575),
    .A2(_0534_));
 sg13g2_nand3_1 _3651_ (.B(net522),
    .C(net488),
    .A(net524),
    .Y(_0774_));
 sg13g2_nor2_2 _3652_ (.A(net527),
    .B(_0774_),
    .Y(_0775_));
 sg13g2_nand2b_2 _3653_ (.Y(_0776_),
    .B(net502),
    .A_N(_0774_));
 sg13g2_nor2_2 _3654_ (.A(_0773_),
    .B(_0776_),
    .Y(_0777_));
 sg13g2_mux2_1 _3655_ (.A0(net608),
    .A1(net475),
    .S(_0777_),
    .X(_0021_));
 sg13g2_mux2_1 _3656_ (.A0(net618),
    .A1(net463),
    .S(_0777_),
    .X(_0022_));
 sg13g2_mux2_1 _3657_ (.A0(net629),
    .A1(net453),
    .S(_0777_),
    .X(_0023_));
 sg13g2_mux2_1 _3658_ (.A0(net633),
    .A1(net441),
    .S(_0777_),
    .X(_0024_));
 sg13g2_nor2_2 _3659_ (.A(net502),
    .B(_0774_),
    .Y(_0778_));
 sg13g2_nand2_2 _3660_ (.Y(_0779_),
    .A(_0758_),
    .B(_0778_));
 sg13g2_mux2_1 _3661_ (.A0(net473),
    .A1(net673),
    .S(_0779_),
    .X(_0025_));
 sg13g2_mux2_1 _3662_ (.A0(net462),
    .A1(net641),
    .S(_0779_),
    .X(_0026_));
 sg13g2_mux2_1 _3663_ (.A0(net452),
    .A1(net642),
    .S(_0779_),
    .X(_0027_));
 sg13g2_mux2_1 _3664_ (.A0(net441),
    .A1(net651),
    .S(_0779_),
    .X(_0028_));
 sg13g2_nor2b_1 _3665_ (.A(uio_out[5]),
    .B_N(uio_out[4]),
    .Y(_0780_));
 sg13g2_and2_2 _3666_ (.A(net580),
    .B(_0780_),
    .X(_0781_));
 sg13g2_nand2_1 _3667_ (.Y(_0782_),
    .A(net579),
    .B(net489));
 sg13g2_nand2_1 _3668_ (.Y(_0783_),
    .A(net765),
    .B(net713));
 sg13g2_nor2_1 _3669_ (.A(net485),
    .B(net714),
    .Y(_0029_));
 sg13g2_a22oi_1 _3670_ (.Y(_0784_),
    .B1(net727),
    .B2(\mem[1][0] ),
    .A2(\mem[1][1] ),
    .A1(net713));
 sg13g2_nand2_1 _3671_ (.Y(_0785_),
    .A(\mem[1][1] ),
    .B(\mem[17][1] ));
 sg13g2_or2_1 _3672_ (.X(_0786_),
    .B(_0785_),
    .A(_0783_));
 sg13g2_inv_1 _3673_ (.Y(_0787_),
    .A(_0786_));
 sg13g2_nor3_1 _3674_ (.A(net485),
    .B(net728),
    .C(_0787_),
    .Y(_0030_));
 sg13g2_nand2_1 _3675_ (.Y(_0788_),
    .A(\mem[1][0] ),
    .B(\mem[17][2] ));
 sg13g2_nand2_2 _3676_ (.Y(_0789_),
    .A(\mem[17][1] ),
    .B(\mem[1][2] ));
 sg13g2_nand2_1 _3677_ (.Y(_0790_),
    .A(\mem[17][0] ),
    .B(\mem[1][2] ));
 sg13g2_or2_1 _3678_ (.X(_0791_),
    .B(_0790_),
    .A(_0785_));
 sg13g2_xnor2_1 _3679_ (.Y(_0792_),
    .A(_0785_),
    .B(_0790_));
 sg13g2_xnor2_1 _3680_ (.Y(_0793_),
    .A(_0788_),
    .B(_0792_));
 sg13g2_or2_1 _3681_ (.X(_0794_),
    .B(_0793_),
    .A(_0786_));
 sg13g2_nand2_1 _3682_ (.Y(_0795_),
    .A(_0781_),
    .B(_0794_));
 sg13g2_a21oi_1 _3683_ (.A1(_0786_),
    .A2(_0793_),
    .Y(_0031_),
    .B1(_0795_));
 sg13g2_nand2_1 _3684_ (.Y(_0796_),
    .A(\mem[1][0] ),
    .B(\mem[17][3] ));
 sg13g2_o21ai_1 _3685_ (.B1(_0791_),
    .Y(_0797_),
    .A1(_0788_),
    .A2(_0792_));
 sg13g2_nand2_1 _3686_ (.Y(_0798_),
    .A(\mem[1][1] ),
    .B(\mem[17][2] ));
 sg13g2_nand2_1 _3687_ (.Y(_0799_),
    .A(\mem[17][1] ),
    .B(\mem[1][3] ));
 sg13g2_nand2_1 _3688_ (.Y(_0800_),
    .A(\mem[17][0] ),
    .B(\mem[1][3] ));
 sg13g2_xor2_1 _3689_ (.B(_0800_),
    .A(_0789_),
    .X(_0801_));
 sg13g2_nand2b_1 _3690_ (.Y(_0802_),
    .B(_0801_),
    .A_N(_0798_));
 sg13g2_xnor2_1 _3691_ (.Y(_0803_),
    .A(_0798_),
    .B(_0801_));
 sg13g2_nand2_1 _3692_ (.Y(_0804_),
    .A(_0797_),
    .B(_0803_));
 sg13g2_xnor2_1 _3693_ (.Y(_0805_),
    .A(_0797_),
    .B(_0803_));
 sg13g2_xnor2_1 _3694_ (.Y(_0806_),
    .A(_0796_),
    .B(_0805_));
 sg13g2_and2_1 _3695_ (.A(_0794_),
    .B(_0806_),
    .X(_0807_));
 sg13g2_nor2_1 _3696_ (.A(_0794_),
    .B(_0806_),
    .Y(_0808_));
 sg13g2_nor3_1 _3697_ (.A(net485),
    .B(_0807_),
    .C(_0808_),
    .Y(_0032_));
 sg13g2_nand2_1 _3698_ (.Y(_0809_),
    .A(\mem[1][1] ),
    .B(\mem[17][3] ));
 sg13g2_o21ai_1 _3699_ (.B1(_0802_),
    .Y(_0810_),
    .A1(_0789_),
    .A2(_0800_));
 sg13g2_nand2_1 _3700_ (.Y(_0811_),
    .A(\mem[1][2] ),
    .B(\mem[17][2] ));
 sg13g2_nand2_1 _3701_ (.Y(_0812_),
    .A(\mem[17][2] ),
    .B(\mem[1][3] ));
 sg13g2_xor2_1 _3702_ (.B(_0811_),
    .A(_0799_),
    .X(_0813_));
 sg13g2_nand2_1 _3703_ (.Y(_0814_),
    .A(_0810_),
    .B(_0813_));
 sg13g2_xor2_1 _3704_ (.B(_0813_),
    .A(_0810_),
    .X(_0815_));
 sg13g2_nand2b_1 _3705_ (.Y(_0816_),
    .B(_0815_),
    .A_N(_0809_));
 sg13g2_xnor2_1 _3706_ (.Y(_0817_),
    .A(_0809_),
    .B(_0815_));
 sg13g2_o21ai_1 _3707_ (.B1(_0804_),
    .Y(_0818_),
    .A1(_0796_),
    .A2(_0805_));
 sg13g2_nand2_1 _3708_ (.Y(_0819_),
    .A(_0817_),
    .B(_0818_));
 sg13g2_xor2_1 _3709_ (.B(_0818_),
    .A(_0817_),
    .X(_0820_));
 sg13g2_or2_1 _3710_ (.X(_0821_),
    .B(_0820_),
    .A(_0808_));
 sg13g2_nand2_1 _3711_ (.Y(_0822_),
    .A(_0808_),
    .B(_0820_));
 sg13g2_and3_1 _3712_ (.X(_0033_),
    .A(_0781_),
    .B(_0821_),
    .C(_0822_));
 sg13g2_nand2b_1 _3713_ (.Y(_0823_),
    .B(_0789_),
    .A_N(_0812_));
 sg13g2_nand2_1 _3714_ (.Y(_0824_),
    .A(\mem[1][2] ),
    .B(\mem[17][3] ));
 sg13g2_xnor2_1 _3715_ (.Y(_0825_),
    .A(_0823_),
    .B(_0824_));
 sg13g2_nand3_1 _3716_ (.B(_0816_),
    .C(_0825_),
    .A(_0814_),
    .Y(_0826_));
 sg13g2_inv_1 _3717_ (.Y(_0827_),
    .A(_0826_));
 sg13g2_a21o_1 _3718_ (.A2(_0816_),
    .A1(_0814_),
    .B1(_0825_),
    .X(_0828_));
 sg13g2_nand2_1 _3719_ (.Y(_0829_),
    .A(_0826_),
    .B(_0828_));
 sg13g2_nand2_1 _3720_ (.Y(_0830_),
    .A(_0819_),
    .B(_0822_));
 sg13g2_xor2_1 _3721_ (.B(_0830_),
    .A(_0829_),
    .X(_0831_));
 sg13g2_nor2_1 _3722_ (.A(net485),
    .B(_0831_),
    .Y(_0034_));
 sg13g2_a21oi_1 _3723_ (.A1(_0789_),
    .A2(_0824_),
    .Y(_0832_),
    .B1(_0812_));
 sg13g2_nand2_1 _3724_ (.Y(_0833_),
    .A(\mem[1][3] ),
    .B(\mem[17][3] ));
 sg13g2_nand2b_1 _3725_ (.Y(_0834_),
    .B(_0832_),
    .A_N(_0833_));
 sg13g2_xnor2_1 _3726_ (.Y(_0835_),
    .A(_0832_),
    .B(_0833_));
 sg13g2_o21ai_1 _3727_ (.B1(_0828_),
    .Y(_0836_),
    .A1(_0819_),
    .A2(_0827_));
 sg13g2_or2_1 _3728_ (.X(_0837_),
    .B(_0836_),
    .A(_0835_));
 sg13g2_nand2_1 _3729_ (.Y(_0838_),
    .A(_0835_),
    .B(_0836_));
 sg13g2_nand3_1 _3730_ (.B(_0837_),
    .C(_0838_),
    .A(_0781_),
    .Y(_0839_));
 sg13g2_inv_1 _3731_ (.Y(_0035_),
    .A(_0839_));
 sg13g2_a21oi_1 _3732_ (.A1(_0834_),
    .A2(_0838_),
    .Y(_0036_),
    .B1(net485));
 sg13g2_nand3_1 _3733_ (.B(net531),
    .C(net488),
    .A(net538),
    .Y(_0840_));
 sg13g2_nor2_2 _3734_ (.A(net518),
    .B(_0840_),
    .Y(_0841_));
 sg13g2_or2_2 _3735_ (.X(_0842_),
    .B(_0840_),
    .A(net515));
 sg13g2_nand2_2 _3736_ (.Y(_0843_),
    .A(_0778_),
    .B(_0841_));
 sg13g2_mux2_1 _3737_ (.A0(net472),
    .A1(net664),
    .S(_0843_),
    .X(_0037_));
 sg13g2_mux2_1 _3738_ (.A0(net461),
    .A1(net638),
    .S(_0843_),
    .X(_0038_));
 sg13g2_mux2_1 _3739_ (.A0(net451),
    .A1(net636),
    .S(_0843_),
    .X(_0039_));
 sg13g2_mux2_1 _3740_ (.A0(net442),
    .A1(net653),
    .S(_0843_),
    .X(_0040_));
 sg13g2_and2_2 _3741_ (.A(net504),
    .B(_0539_),
    .X(_0844_));
 sg13g2_nand2_2 _3742_ (.Y(_0845_),
    .A(net504),
    .B(_0539_));
 sg13g2_nor2_2 _3743_ (.A(net552),
    .B(_0840_),
    .Y(_0846_));
 sg13g2_nand2b_2 _3744_ (.Y(_0847_),
    .B(net516),
    .A_N(_0840_));
 sg13g2_nor2_2 _3745_ (.A(_0845_),
    .B(_0847_),
    .Y(_0848_));
 sg13g2_mux2_1 _3746_ (.A0(net725),
    .A1(net481),
    .S(_0848_),
    .X(_0041_));
 sg13g2_mux2_1 _3747_ (.A0(net762),
    .A1(net469),
    .S(_0848_),
    .X(_0042_));
 sg13g2_nand2_1 _3748_ (.Y(_0849_),
    .A(net458),
    .B(_0848_));
 sg13g2_o21ai_1 _3749_ (.B1(_0849_),
    .Y(_0043_),
    .A1(_2102_),
    .A2(_0848_));
 sg13g2_mux2_1 _3750_ (.A0(net752),
    .A1(net448),
    .S(_0848_),
    .X(_0044_));
 sg13g2_nand2_2 _3751_ (.Y(_0850_),
    .A(_0841_),
    .B(_0844_));
 sg13g2_mux2_1 _3752_ (.A0(net481),
    .A1(net707),
    .S(_0850_),
    .X(_0045_));
 sg13g2_mux2_1 _3753_ (.A0(net469),
    .A1(net763),
    .S(_0850_),
    .X(_0046_));
 sg13g2_mux2_1 _3754_ (.A0(net458),
    .A1(net766),
    .S(_0850_),
    .X(_0047_));
 sg13g2_mux2_1 _3755_ (.A0(net448),
    .A1(net756),
    .S(_0850_),
    .X(_0048_));
 sg13g2_nor2_2 _3756_ (.A(_0770_),
    .B(_0845_),
    .Y(_0851_));
 sg13g2_mux2_1 _3757_ (.A0(net684),
    .A1(net481),
    .S(_0851_),
    .X(_0049_));
 sg13g2_mux2_1 _3758_ (.A0(net749),
    .A1(net469),
    .S(_0851_),
    .X(_0050_));
 sg13g2_mux2_1 _3759_ (.A0(net767),
    .A1(net458),
    .S(_0851_),
    .X(_0051_));
 sg13g2_mux2_1 _3760_ (.A0(net724),
    .A1(net448),
    .S(_0851_),
    .X(_0052_));
 sg13g2_and3_2 _3761_ (.X(_0852_),
    .A(uio_out[5]),
    .B(uio_out[4]),
    .C(net578));
 sg13g2_nand3_1 _3762_ (.B(net733),
    .C(net578),
    .A(uio_out[5]),
    .Y(_0853_));
 sg13g2_a21oi_2 _3763_ (.B1(_0752_),
    .Y(_0854_),
    .A2(_0753_),
    .A1(_0684_));
 sg13g2_o21ai_1 _3764_ (.B1(_0698_),
    .Y(_0855_),
    .A1(_0692_),
    .A2(_0699_));
 sg13g2_a21oi_1 _3765_ (.A1(_0700_),
    .A2(_0747_),
    .Y(_0856_),
    .B1(_0746_));
 sg13g2_a21oi_1 _3766_ (.A1(\products[15][3] ),
    .A2(_0696_),
    .Y(_0857_),
    .B1(_0695_));
 sg13g2_a21oi_1 _3767_ (.A1(_0704_),
    .A2(_0715_),
    .Y(_0858_),
    .B1(_0717_));
 sg13g2_a21oi_2 _3768_ (.B1(_0705_),
    .Y(_0859_),
    .A2(_0706_),
    .A1(\products[13][3] ));
 sg13g2_nor2b_1 _3769_ (.A(_0859_),
    .B_N(\products[14][4] ),
    .Y(_0860_));
 sg13g2_xnor2_1 _3770_ (.Y(_0861_),
    .A(\products[14][4] ),
    .B(_0859_));
 sg13g2_xnor2_1 _3771_ (.Y(_0862_),
    .A(\products[15][4] ),
    .B(_0861_));
 sg13g2_or2_1 _3772_ (.X(_0863_),
    .B(_0862_),
    .A(_0858_));
 sg13g2_xnor2_1 _3773_ (.Y(_0864_),
    .A(_0858_),
    .B(_0862_));
 sg13g2_xor2_1 _3774_ (.B(_0864_),
    .A(_0857_),
    .X(_0865_));
 sg13g2_a21oi_1 _3775_ (.A1(_0718_),
    .A2(_0744_),
    .Y(_0866_),
    .B1(_0743_));
 sg13g2_a21oi_2 _3776_ (.B1(_0713_),
    .Y(_0867_),
    .A2(_0714_),
    .A1(_0708_));
 sg13g2_a21oi_1 _3777_ (.A1(_0720_),
    .A2(_0726_),
    .Y(_0868_),
    .B1(_0725_));
 sg13g2_and2_1 _3778_ (.A(\products[12][4] ),
    .B(\products[11][4] ),
    .X(_0869_));
 sg13g2_xor2_1 _3779_ (.B(\products[11][4] ),
    .A(\products[12][4] ),
    .X(_0870_));
 sg13g2_xnor2_1 _3780_ (.Y(_0871_),
    .A(\products[13][4] ),
    .B(_0870_));
 sg13g2_inv_1 _3781_ (.Y(_0872_),
    .A(_0871_));
 sg13g2_a21oi_2 _3782_ (.B1(_0710_),
    .Y(_0873_),
    .A2(_0711_),
    .A1(\products[10][3] ));
 sg13g2_and2_1 _3783_ (.A(\products[9][4] ),
    .B(\products[8][4] ),
    .X(_0874_));
 sg13g2_xor2_1 _3784_ (.B(\products[8][4] ),
    .A(\products[9][4] ),
    .X(_0875_));
 sg13g2_xnor2_1 _3785_ (.Y(_0876_),
    .A(\products[10][4] ),
    .B(_0875_));
 sg13g2_nor2_1 _3786_ (.A(_0873_),
    .B(_0876_),
    .Y(_0877_));
 sg13g2_xor2_1 _3787_ (.B(_0876_),
    .A(_0873_),
    .X(_0878_));
 sg13g2_xnor2_1 _3788_ (.Y(_0879_),
    .A(_0871_),
    .B(_0878_));
 sg13g2_nand2b_1 _3789_ (.Y(_0880_),
    .B(_0879_),
    .A_N(_0868_));
 sg13g2_xnor2_1 _3790_ (.Y(_0881_),
    .A(_0868_),
    .B(_0879_));
 sg13g2_nand2b_1 _3791_ (.Y(_0882_),
    .B(_0881_),
    .A_N(_0867_));
 sg13g2_xnor2_1 _3792_ (.Y(_0883_),
    .A(_0867_),
    .B(_0881_));
 sg13g2_a21oi_1 _3793_ (.A1(_0727_),
    .A2(_0741_),
    .Y(_0884_),
    .B1(_0740_));
 sg13g2_a21oi_1 _3794_ (.A1(\products[7][3] ),
    .A2(_0723_),
    .Y(_0885_),
    .B1(_0722_));
 sg13g2_a21oi_2 _3795_ (.B1(_0729_),
    .Y(_0886_),
    .A2(_0730_),
    .A1(\products[4][3] ));
 sg13g2_and2_1 _3796_ (.A(\products[6][4] ),
    .B(\products[5][4] ),
    .X(_0887_));
 sg13g2_xor2_1 _3797_ (.B(\products[5][4] ),
    .A(\products[6][4] ),
    .X(_0888_));
 sg13g2_xnor2_1 _3798_ (.Y(_0889_),
    .A(\products[7][4] ),
    .B(_0888_));
 sg13g2_nor2_1 _3799_ (.A(_0886_),
    .B(_0889_),
    .Y(_0890_));
 sg13g2_xnor2_1 _3800_ (.Y(_0891_),
    .A(_0886_),
    .B(_0889_));
 sg13g2_nor2_1 _3801_ (.A(_0885_),
    .B(_0891_),
    .Y(_0892_));
 sg13g2_xor2_1 _3802_ (.B(_0891_),
    .A(_0885_),
    .X(_0893_));
 sg13g2_a21oi_2 _3803_ (.B1(_0737_),
    .Y(_0894_),
    .A2(_0738_),
    .A1(_0732_));
 sg13g2_and2_1 _3804_ (.A(\products[3][4] ),
    .B(\products[2][4] ),
    .X(_0895_));
 sg13g2_xor2_1 _3805_ (.B(\products[2][4] ),
    .A(\products[3][4] ),
    .X(_0896_));
 sg13g2_xnor2_1 _3806_ (.Y(_0897_),
    .A(\products[4][4] ),
    .B(_0896_));
 sg13g2_inv_1 _3807_ (.Y(_0898_),
    .A(_0897_));
 sg13g2_a21oi_2 _3808_ (.B1(_0734_),
    .Y(_0899_),
    .A2(_0735_),
    .A1(\products[1][3] ));
 sg13g2_and2_1 _3809_ (.A(\prev_acc[4] ),
    .B(\products[0][4] ),
    .X(_0900_));
 sg13g2_xor2_1 _3810_ (.B(\products[0][4] ),
    .A(\prev_acc[4] ),
    .X(_0901_));
 sg13g2_xnor2_1 _3811_ (.Y(_0902_),
    .A(\products[1][4] ),
    .B(_0901_));
 sg13g2_nor2_1 _3812_ (.A(_0899_),
    .B(_0902_),
    .Y(_0903_));
 sg13g2_xor2_1 _3813_ (.B(_0902_),
    .A(_0899_),
    .X(_0904_));
 sg13g2_xnor2_1 _3814_ (.Y(_0905_),
    .A(_0898_),
    .B(_0904_));
 sg13g2_nor2_1 _3815_ (.A(_0894_),
    .B(_0905_),
    .Y(_0906_));
 sg13g2_xor2_1 _3816_ (.B(_0905_),
    .A(_0894_),
    .X(_0907_));
 sg13g2_xnor2_1 _3817_ (.Y(_0908_),
    .A(_0893_),
    .B(_0907_));
 sg13g2_nor2_1 _3818_ (.A(_0884_),
    .B(_0908_),
    .Y(_0909_));
 sg13g2_xor2_1 _3819_ (.B(_0908_),
    .A(_0884_),
    .X(_0910_));
 sg13g2_xnor2_1 _3820_ (.Y(_0911_),
    .A(_0883_),
    .B(_0910_));
 sg13g2_nor2_1 _3821_ (.A(_0866_),
    .B(_0911_),
    .Y(_0912_));
 sg13g2_xor2_1 _3822_ (.B(_0911_),
    .A(_0866_),
    .X(_0913_));
 sg13g2_xnor2_1 _3823_ (.Y(_0914_),
    .A(_0865_),
    .B(_0913_));
 sg13g2_nor2_1 _3824_ (.A(_0856_),
    .B(_0914_),
    .Y(_0915_));
 sg13g2_xor2_1 _3825_ (.B(_0914_),
    .A(_0856_),
    .X(_0916_));
 sg13g2_xnor2_1 _3826_ (.Y(_0917_),
    .A(_0855_),
    .B(_0916_));
 sg13g2_a21oi_1 _3827_ (.A1(_0690_),
    .A2(_0750_),
    .Y(_0918_),
    .B1(_0749_));
 sg13g2_nor2_1 _3828_ (.A(_0917_),
    .B(_0918_),
    .Y(_0919_));
 sg13g2_xnor2_1 _3829_ (.Y(_0920_),
    .A(_0917_),
    .B(_0918_));
 sg13g2_nor2_1 _3830_ (.A(_0854_),
    .B(_0920_),
    .Y(_0921_));
 sg13g2_xnor2_1 _3831_ (.Y(_0922_),
    .A(_0854_),
    .B(_0920_));
 sg13g2_o21ai_1 _3832_ (.B1(_0760_),
    .Y(_0923_),
    .A1(net523),
    .A2(_0534_));
 sg13g2_a21o_2 _3833_ (.A2(net487),
    .A1(net529),
    .B1(_0923_),
    .X(_0924_));
 sg13g2_nor2_2 _3834_ (.A(_0770_),
    .B(_0924_),
    .Y(_0925_));
 sg13g2_nor2b_1 _3835_ (.A(net477),
    .B_N(_0925_),
    .Y(_0926_));
 sg13g2_nor2_2 _3836_ (.A(_0852_),
    .B(_0925_),
    .Y(_0927_));
 sg13g2_a221oi_1 _3837_ (.B2(_2085_),
    .C1(_0926_),
    .B1(_0927_),
    .A1(_0852_),
    .Y(_0053_),
    .A2(_0922_));
 sg13g2_a21oi_2 _3838_ (.B1(_0915_),
    .Y(_0928_),
    .A2(_0916_),
    .A1(_0855_));
 sg13g2_o21ai_1 _3839_ (.B1(_0863_),
    .Y(_0929_),
    .A1(_0857_),
    .A2(_0864_));
 sg13g2_a21oi_1 _3840_ (.A1(_0865_),
    .A2(_0913_),
    .Y(_0930_),
    .B1(_0912_));
 sg13g2_a21oi_1 _3841_ (.A1(\products[15][4] ),
    .A2(_0861_),
    .Y(_0931_),
    .B1(_0860_));
 sg13g2_nand2_1 _3842_ (.Y(_0932_),
    .A(_0880_),
    .B(_0882_));
 sg13g2_a21oi_2 _3843_ (.B1(_0869_),
    .Y(_0933_),
    .A2(_0870_),
    .A1(\products[13][4] ));
 sg13g2_nor2b_1 _3844_ (.A(_0933_),
    .B_N(\products[14][5] ),
    .Y(_0934_));
 sg13g2_xnor2_1 _3845_ (.Y(_0935_),
    .A(\products[14][5] ),
    .B(_0933_));
 sg13g2_xnor2_1 _3846_ (.Y(_0936_),
    .A(\products[15][5] ),
    .B(_0935_));
 sg13g2_nand2b_1 _3847_ (.Y(_0937_),
    .B(_0932_),
    .A_N(_0936_));
 sg13g2_xor2_1 _3848_ (.B(_0936_),
    .A(_0932_),
    .X(_0938_));
 sg13g2_xor2_1 _3849_ (.B(_0938_),
    .A(_0931_),
    .X(_0939_));
 sg13g2_a21oi_1 _3850_ (.A1(_0883_),
    .A2(_0910_),
    .Y(_0940_),
    .B1(_0909_));
 sg13g2_a21oi_2 _3851_ (.B1(_0877_),
    .Y(_0941_),
    .A2(_0878_),
    .A1(_0872_));
 sg13g2_nor2_2 _3852_ (.A(_0890_),
    .B(_0892_),
    .Y(_0942_));
 sg13g2_and2_1 _3853_ (.A(\products[12][5] ),
    .B(\products[11][5] ),
    .X(_0943_));
 sg13g2_xor2_1 _3854_ (.B(\products[11][5] ),
    .A(\products[12][5] ),
    .X(_0944_));
 sg13g2_xnor2_1 _3855_ (.Y(_0945_),
    .A(\products[13][5] ),
    .B(_0944_));
 sg13g2_inv_1 _3856_ (.Y(_0946_),
    .A(_0945_));
 sg13g2_a21oi_2 _3857_ (.B1(_0874_),
    .Y(_0947_),
    .A2(_0875_),
    .A1(\products[10][4] ));
 sg13g2_and2_1 _3858_ (.A(\products[9][5] ),
    .B(\products[8][5] ),
    .X(_0948_));
 sg13g2_xor2_1 _3859_ (.B(\products[8][5] ),
    .A(\products[9][5] ),
    .X(_0949_));
 sg13g2_xnor2_1 _3860_ (.Y(_0950_),
    .A(\products[10][5] ),
    .B(_0949_));
 sg13g2_nor2_1 _3861_ (.A(_0947_),
    .B(_0950_),
    .Y(_0951_));
 sg13g2_xor2_1 _3862_ (.B(_0950_),
    .A(_0947_),
    .X(_0952_));
 sg13g2_xnor2_1 _3863_ (.Y(_0953_),
    .A(_0945_),
    .B(_0952_));
 sg13g2_nor2b_1 _3864_ (.A(_0942_),
    .B_N(_0953_),
    .Y(_0954_));
 sg13g2_xnor2_1 _3865_ (.Y(_0955_),
    .A(_0942_),
    .B(_0953_));
 sg13g2_nor2b_1 _3866_ (.A(_0941_),
    .B_N(_0955_),
    .Y(_0956_));
 sg13g2_xnor2_1 _3867_ (.Y(_0957_),
    .A(_0941_),
    .B(_0955_));
 sg13g2_a21oi_1 _3868_ (.A1(_0893_),
    .A2(_0907_),
    .Y(_0958_),
    .B1(_0906_));
 sg13g2_a21oi_1 _3869_ (.A1(\products[7][4] ),
    .A2(_0888_),
    .Y(_0959_),
    .B1(_0887_));
 sg13g2_a21oi_2 _3870_ (.B1(_0895_),
    .Y(_0960_),
    .A2(_0896_),
    .A1(\products[4][4] ));
 sg13g2_and2_1 _3871_ (.A(\products[6][5] ),
    .B(\products[5][5] ),
    .X(_0961_));
 sg13g2_xor2_1 _3872_ (.B(\products[5][5] ),
    .A(\products[6][5] ),
    .X(_0962_));
 sg13g2_xnor2_1 _3873_ (.Y(_0963_),
    .A(\products[7][5] ),
    .B(_0962_));
 sg13g2_nor2_1 _3874_ (.A(_0960_),
    .B(_0963_),
    .Y(_0964_));
 sg13g2_xor2_1 _3875_ (.B(_0963_),
    .A(_0960_),
    .X(_0965_));
 sg13g2_nor2b_1 _3876_ (.A(_0959_),
    .B_N(_0965_),
    .Y(_0966_));
 sg13g2_xnor2_1 _3877_ (.Y(_0967_),
    .A(_0959_),
    .B(_0965_));
 sg13g2_a21oi_2 _3878_ (.B1(_0903_),
    .Y(_0968_),
    .A2(_0904_),
    .A1(_0898_));
 sg13g2_and2_1 _3879_ (.A(\products[3][5] ),
    .B(\products[2][5] ),
    .X(_0969_));
 sg13g2_xor2_1 _3880_ (.B(\products[2][5] ),
    .A(\products[3][5] ),
    .X(_0970_));
 sg13g2_xnor2_1 _3881_ (.Y(_0971_),
    .A(\products[4][5] ),
    .B(_0970_));
 sg13g2_inv_1 _3882_ (.Y(_0972_),
    .A(_0971_));
 sg13g2_a21oi_2 _3883_ (.B1(_0900_),
    .Y(_0973_),
    .A2(_0901_),
    .A1(\products[1][4] ));
 sg13g2_and2_1 _3884_ (.A(\prev_acc[5] ),
    .B(\products[0][5] ),
    .X(_0974_));
 sg13g2_xor2_1 _3885_ (.B(\products[0][5] ),
    .A(\prev_acc[5] ),
    .X(_0975_));
 sg13g2_xnor2_1 _3886_ (.Y(_0976_),
    .A(\products[1][5] ),
    .B(_0975_));
 sg13g2_nor2_1 _3887_ (.A(_0973_),
    .B(_0976_),
    .Y(_0977_));
 sg13g2_xor2_1 _3888_ (.B(_0976_),
    .A(_0973_),
    .X(_0978_));
 sg13g2_xnor2_1 _3889_ (.Y(_0979_),
    .A(_0971_),
    .B(_0978_));
 sg13g2_nor2b_1 _3890_ (.A(_0968_),
    .B_N(_0979_),
    .Y(_0980_));
 sg13g2_xnor2_1 _3891_ (.Y(_0981_),
    .A(_0968_),
    .B(_0979_));
 sg13g2_xnor2_1 _3892_ (.Y(_0982_),
    .A(_0967_),
    .B(_0981_));
 sg13g2_nor2_1 _3893_ (.A(_0958_),
    .B(_0982_),
    .Y(_0983_));
 sg13g2_xor2_1 _3894_ (.B(_0982_),
    .A(_0958_),
    .X(_0984_));
 sg13g2_xnor2_1 _3895_ (.Y(_0985_),
    .A(_0957_),
    .B(_0984_));
 sg13g2_nor2_1 _3896_ (.A(_0940_),
    .B(_0985_),
    .Y(_0986_));
 sg13g2_xor2_1 _3897_ (.B(_0985_),
    .A(_0940_),
    .X(_0987_));
 sg13g2_xnor2_1 _3898_ (.Y(_0988_),
    .A(_0939_),
    .B(_0987_));
 sg13g2_nor2_1 _3899_ (.A(_0930_),
    .B(_0988_),
    .Y(_0989_));
 sg13g2_xor2_1 _3900_ (.B(_0988_),
    .A(_0930_),
    .X(_0990_));
 sg13g2_xnor2_1 _3901_ (.Y(_0991_),
    .A(_0929_),
    .B(_0990_));
 sg13g2_nor2_1 _3902_ (.A(_0928_),
    .B(_0991_),
    .Y(_0992_));
 sg13g2_nand2_1 _3903_ (.Y(_0993_),
    .A(_0928_),
    .B(_0991_));
 sg13g2_xor2_1 _3904_ (.B(_0991_),
    .A(_0928_),
    .X(_0994_));
 sg13g2_nor2_1 _3905_ (.A(_0919_),
    .B(_0921_),
    .Y(_0995_));
 sg13g2_xor2_1 _3906_ (.B(_0995_),
    .A(_0994_),
    .X(_0996_));
 sg13g2_a22oi_1 _3907_ (.Y(_0997_),
    .B1(_0927_),
    .B2(net703),
    .A2(_0925_),
    .A1(net465));
 sg13g2_o21ai_1 _3908_ (.B1(_0997_),
    .Y(_0054_),
    .A1(_0853_),
    .A2(_0996_));
 sg13g2_nand2b_1 _3909_ (.Y(_0998_),
    .B(_0994_),
    .A_N(_0920_));
 sg13g2_a21oi_1 _3910_ (.A1(_0919_),
    .A2(_0993_),
    .Y(_0999_),
    .B1(_0992_));
 sg13g2_o21ai_1 _3911_ (.B1(_0999_),
    .Y(_1000_),
    .A1(_0854_),
    .A2(_0998_));
 sg13g2_o21ai_1 _3912_ (.B1(_0937_),
    .Y(_1001_),
    .A1(_0931_),
    .A2(_0938_));
 sg13g2_a21oi_1 _3913_ (.A1(_0939_),
    .A2(_0987_),
    .Y(_1002_),
    .B1(_0986_));
 sg13g2_a21oi_1 _3914_ (.A1(\products[15][5] ),
    .A2(_0935_),
    .Y(_1003_),
    .B1(_0934_));
 sg13g2_nor2_1 _3915_ (.A(_0954_),
    .B(_0956_),
    .Y(_1004_));
 sg13g2_a21oi_2 _3916_ (.B1(_0943_),
    .Y(_1005_),
    .A2(_0944_),
    .A1(\products[13][5] ));
 sg13g2_nor2b_1 _3917_ (.A(_1005_),
    .B_N(\products[14][6] ),
    .Y(_1006_));
 sg13g2_xnor2_1 _3918_ (.Y(_1007_),
    .A(\products[14][6] ),
    .B(_1005_));
 sg13g2_xnor2_1 _3919_ (.Y(_1008_),
    .A(\products[15][6] ),
    .B(_1007_));
 sg13g2_or2_1 _3920_ (.X(_1009_),
    .B(_1008_),
    .A(_1004_));
 sg13g2_xnor2_1 _3921_ (.Y(_1010_),
    .A(_1004_),
    .B(_1008_));
 sg13g2_xor2_1 _3922_ (.B(_1010_),
    .A(_1003_),
    .X(_1011_));
 sg13g2_a21oi_1 _3923_ (.A1(_0957_),
    .A2(_0984_),
    .Y(_1012_),
    .B1(_0983_));
 sg13g2_a21oi_1 _3924_ (.A1(_0967_),
    .A2(_0981_),
    .Y(_1013_),
    .B1(_0980_));
 sg13g2_a21oi_2 _3925_ (.B1(_0977_),
    .Y(_1014_),
    .A2(_0978_),
    .A1(_0972_));
 sg13g2_a21oi_1 _3926_ (.A1(\products[1][5] ),
    .A2(_0975_),
    .Y(_1015_),
    .B1(_0974_));
 sg13g2_and2_1 _3927_ (.A(\prev_acc[6] ),
    .B(\products[0][6] ),
    .X(_1016_));
 sg13g2_xor2_1 _3928_ (.B(\products[0][6] ),
    .A(\prev_acc[6] ),
    .X(_1017_));
 sg13g2_xnor2_1 _3929_ (.Y(_1018_),
    .A(\products[1][6] ),
    .B(_1017_));
 sg13g2_or2_1 _3930_ (.X(_1019_),
    .B(_1018_),
    .A(_1015_));
 sg13g2_xnor2_1 _3931_ (.Y(_1020_),
    .A(_1015_),
    .B(_1018_));
 sg13g2_and2_1 _3932_ (.A(\products[3][6] ),
    .B(\products[2][6] ),
    .X(_1021_));
 sg13g2_xor2_1 _3933_ (.B(\products[2][6] ),
    .A(\products[3][6] ),
    .X(_1022_));
 sg13g2_xnor2_1 _3934_ (.Y(_1023_),
    .A(\products[4][6] ),
    .B(_1022_));
 sg13g2_xnor2_1 _3935_ (.Y(_1024_),
    .A(_1020_),
    .B(_1023_));
 sg13g2_nor2_1 _3936_ (.A(_1014_),
    .B(_1024_),
    .Y(_1025_));
 sg13g2_xor2_1 _3937_ (.B(_1024_),
    .A(_1014_),
    .X(_1026_));
 sg13g2_a21oi_1 _3938_ (.A1(\products[7][5] ),
    .A2(_0962_),
    .Y(_1027_),
    .B1(_0961_));
 sg13g2_a21oi_2 _3939_ (.B1(_0969_),
    .Y(_1028_),
    .A2(_0970_),
    .A1(\products[4][5] ));
 sg13g2_and2_1 _3940_ (.A(\products[6][6] ),
    .B(\products[5][6] ),
    .X(_1029_));
 sg13g2_xor2_1 _3941_ (.B(\products[5][6] ),
    .A(\products[6][6] ),
    .X(_1030_));
 sg13g2_xnor2_1 _3942_ (.Y(_1031_),
    .A(\products[7][6] ),
    .B(_1030_));
 sg13g2_xor2_1 _3943_ (.B(_1031_),
    .A(_1028_),
    .X(_1032_));
 sg13g2_nand2b_1 _3944_ (.Y(_1033_),
    .B(_1032_),
    .A_N(_1027_));
 sg13g2_xnor2_1 _3945_ (.Y(_1034_),
    .A(_1027_),
    .B(_1032_));
 sg13g2_xnor2_1 _3946_ (.Y(_1035_),
    .A(_1026_),
    .B(_1034_));
 sg13g2_nor2_1 _3947_ (.A(_1013_),
    .B(_1035_),
    .Y(_1036_));
 sg13g2_xor2_1 _3948_ (.B(_1035_),
    .A(_1013_),
    .X(_1037_));
 sg13g2_a21oi_2 _3949_ (.B1(_0951_),
    .Y(_1038_),
    .A2(_0952_),
    .A1(_0946_));
 sg13g2_and2_1 _3950_ (.A(\products[12][6] ),
    .B(\products[11][6] ),
    .X(_1039_));
 sg13g2_xor2_1 _3951_ (.B(\products[11][6] ),
    .A(\products[12][6] ),
    .X(_1040_));
 sg13g2_xnor2_1 _3952_ (.Y(_1041_),
    .A(\products[13][6] ),
    .B(_1040_));
 sg13g2_a21oi_2 _3953_ (.B1(_0948_),
    .Y(_1042_),
    .A2(_0949_),
    .A1(\products[10][5] ));
 sg13g2_and2_1 _3954_ (.A(\products[9][6] ),
    .B(\products[8][6] ),
    .X(_1043_));
 sg13g2_xor2_1 _3955_ (.B(\products[8][6] ),
    .A(\products[9][6] ),
    .X(_1044_));
 sg13g2_xnor2_1 _3956_ (.Y(_1045_),
    .A(\products[10][6] ),
    .B(_1044_));
 sg13g2_xor2_1 _3957_ (.B(_1045_),
    .A(_1042_),
    .X(_1046_));
 sg13g2_nand2b_1 _3958_ (.Y(_1047_),
    .B(_1046_),
    .A_N(_1041_));
 sg13g2_xnor2_1 _3959_ (.Y(_1048_),
    .A(_1041_),
    .B(_1046_));
 sg13g2_o21ai_1 _3960_ (.B1(_1048_),
    .Y(_1049_),
    .A1(_0964_),
    .A2(_0966_));
 sg13g2_or3_1 _3961_ (.A(_0964_),
    .B(_0966_),
    .C(_1048_),
    .X(_1050_));
 sg13g2_and2_1 _3962_ (.A(_1049_),
    .B(_1050_),
    .X(_1051_));
 sg13g2_inv_1 _3963_ (.Y(_1052_),
    .A(_1051_));
 sg13g2_xnor2_1 _3964_ (.Y(_1053_),
    .A(_1038_),
    .B(_1051_));
 sg13g2_xnor2_1 _3965_ (.Y(_1054_),
    .A(_1037_),
    .B(_1053_));
 sg13g2_nor2_1 _3966_ (.A(_1012_),
    .B(_1054_),
    .Y(_1055_));
 sg13g2_xor2_1 _3967_ (.B(_1054_),
    .A(_1012_),
    .X(_1056_));
 sg13g2_xnor2_1 _3968_ (.Y(_1057_),
    .A(_1011_),
    .B(_1056_));
 sg13g2_xnor2_1 _3969_ (.Y(_1058_),
    .A(_1002_),
    .B(_1057_));
 sg13g2_nand2b_1 _3970_ (.Y(_1059_),
    .B(_1001_),
    .A_N(_1058_));
 sg13g2_xor2_1 _3971_ (.B(_1058_),
    .A(_1001_),
    .X(_1060_));
 sg13g2_a21oi_1 _3972_ (.A1(_0929_),
    .A2(_0990_),
    .Y(_1061_),
    .B1(_0989_));
 sg13g2_nor2_1 _3973_ (.A(_1060_),
    .B(_1061_),
    .Y(_1062_));
 sg13g2_xor2_1 _3974_ (.B(_1061_),
    .A(_1060_),
    .X(_1063_));
 sg13g2_and2_1 _3975_ (.A(_1000_),
    .B(_1063_),
    .X(_1064_));
 sg13g2_o21ai_1 _3976_ (.B1(_0852_),
    .Y(_1065_),
    .A1(_1000_),
    .A2(_1063_));
 sg13g2_a22oi_1 _3977_ (.Y(_1066_),
    .B1(_0927_),
    .B2(net741),
    .A2(_0925_),
    .A1(net455));
 sg13g2_o21ai_1 _3978_ (.B1(_1066_),
    .Y(_0055_),
    .A1(_1064_),
    .A2(_1065_));
 sg13g2_a21oi_1 _3979_ (.A1(_1000_),
    .A2(_1063_),
    .Y(_1067_),
    .B1(_1062_));
 sg13g2_o21ai_1 _3980_ (.B1(_1059_),
    .Y(_1068_),
    .A1(_1002_),
    .A2(_1057_));
 sg13g2_a21oi_1 _3981_ (.A1(_1011_),
    .A2(_1056_),
    .Y(_1069_),
    .B1(_1055_));
 sg13g2_o21ai_1 _3982_ (.B1(_1009_),
    .Y(_1070_),
    .A1(_1003_),
    .A2(_1010_));
 sg13g2_a21oi_2 _3983_ (.B1(_1025_),
    .Y(_1071_),
    .A2(_1034_),
    .A1(_1026_));
 sg13g2_o21ai_1 _3984_ (.B1(_1047_),
    .Y(_1072_),
    .A1(_1042_),
    .A2(_1045_));
 sg13g2_xnor2_1 _3985_ (.Y(_1073_),
    .A(_1071_),
    .B(_1072_));
 sg13g2_a21oi_1 _3986_ (.A1(\products[15][6] ),
    .A2(_1007_),
    .Y(_1074_),
    .B1(_1006_));
 sg13g2_a21oi_2 _3987_ (.B1(_1039_),
    .Y(_1075_),
    .A2(_1040_),
    .A1(\products[13][6] ));
 sg13g2_xor2_1 _3988_ (.B(\products[15][7] ),
    .A(\products[14][7] ),
    .X(_1076_));
 sg13g2_xnor2_1 _3989_ (.Y(_1077_),
    .A(_1075_),
    .B(_1076_));
 sg13g2_xnor2_1 _3990_ (.Y(_1078_),
    .A(_1074_),
    .B(_1077_));
 sg13g2_o21ai_1 _3991_ (.B1(_1049_),
    .Y(_1079_),
    .A1(_1038_),
    .A2(_1052_));
 sg13g2_xnor2_1 _3992_ (.Y(_1080_),
    .A(_1078_),
    .B(_1079_));
 sg13g2_xnor2_1 _3993_ (.Y(_1081_),
    .A(_1073_),
    .B(_1080_));
 sg13g2_xnor2_1 _3994_ (.Y(_1082_),
    .A(_1070_),
    .B(_1081_));
 sg13g2_a21oi_1 _3995_ (.A1(\products[4][6] ),
    .A2(_1022_),
    .Y(_1083_),
    .B1(_1021_));
 sg13g2_xnor2_1 _3996_ (.Y(_1084_),
    .A(\prev_acc[7] ),
    .B(\products[2][7] ));
 sg13g2_xnor2_1 _3997_ (.Y(_1085_),
    .A(_1083_),
    .B(_1084_));
 sg13g2_xor2_1 _3998_ (.B(\products[7][7] ),
    .A(\products[5][7] ),
    .X(_1086_));
 sg13g2_xnor2_1 _3999_ (.Y(_1087_),
    .A(\products[6][7] ),
    .B(_1086_));
 sg13g2_xor2_1 _4000_ (.B(\products[1][7] ),
    .A(\products[0][7] ),
    .X(_1088_));
 sg13g2_xnor2_1 _4001_ (.Y(_1089_),
    .A(\products[4][7] ),
    .B(_1088_));
 sg13g2_xnor2_1 _4002_ (.Y(_1090_),
    .A(_1087_),
    .B(_1089_));
 sg13g2_a21oi_1 _4003_ (.A1(\products[1][6] ),
    .A2(_1017_),
    .Y(_1091_),
    .B1(_1016_));
 sg13g2_xnor2_1 _4004_ (.Y(_1092_),
    .A(\products[3][7] ),
    .B(_1091_));
 sg13g2_xnor2_1 _4005_ (.Y(_1093_),
    .A(_1090_),
    .B(_1092_));
 sg13g2_xnor2_1 _4006_ (.Y(_1094_),
    .A(_1085_),
    .B(_1093_));
 sg13g2_o21ai_1 _4007_ (.B1(_1033_),
    .Y(_1095_),
    .A1(_1028_),
    .A2(_1031_));
 sg13g2_a21oi_2 _4008_ (.B1(_1043_),
    .Y(_1096_),
    .A2(_1044_),
    .A1(\products[10][6] ));
 sg13g2_xnor2_1 _4009_ (.Y(_1097_),
    .A(\products[12][7] ),
    .B(_1096_));
 sg13g2_xor2_1 _4010_ (.B(\products[8][7] ),
    .A(\products[9][7] ),
    .X(_1098_));
 sg13g2_xor2_1 _4011_ (.B(\products[13][7] ),
    .A(\products[10][7] ),
    .X(_1099_));
 sg13g2_xnor2_1 _4012_ (.Y(_1100_),
    .A(\products[11][7] ),
    .B(_1099_));
 sg13g2_xnor2_1 _4013_ (.Y(_1101_),
    .A(_1098_),
    .B(_1100_));
 sg13g2_xnor2_1 _4014_ (.Y(_1102_),
    .A(_1097_),
    .B(_1101_));
 sg13g2_xnor2_1 _4015_ (.Y(_1103_),
    .A(_1095_),
    .B(_1102_));
 sg13g2_a21oi_2 _4016_ (.B1(_1029_),
    .Y(_1104_),
    .A2(_1030_),
    .A1(\products[7][6] ));
 sg13g2_o21ai_1 _4017_ (.B1(_1019_),
    .Y(_1105_),
    .A1(_1020_),
    .A2(_1023_));
 sg13g2_xnor2_1 _4018_ (.Y(_1106_),
    .A(_1104_),
    .B(_1105_));
 sg13g2_xnor2_1 _4019_ (.Y(_1107_),
    .A(_1094_),
    .B(_1106_));
 sg13g2_xnor2_1 _4020_ (.Y(_1108_),
    .A(_1103_),
    .B(_1107_));
 sg13g2_a21oi_1 _4021_ (.A1(_1037_),
    .A2(_1053_),
    .Y(_1109_),
    .B1(_1036_));
 sg13g2_xnor2_1 _4022_ (.Y(_1110_),
    .A(_1108_),
    .B(_1109_));
 sg13g2_xnor2_1 _4023_ (.Y(_1111_),
    .A(_1082_),
    .B(_1110_));
 sg13g2_xnor2_1 _4024_ (.Y(_1112_),
    .A(_1069_),
    .B(_1111_));
 sg13g2_xnor2_1 _4025_ (.Y(_1113_),
    .A(_1068_),
    .B(_1112_));
 sg13g2_xnor2_1 _4026_ (.Y(_1114_),
    .A(_1067_),
    .B(_1113_));
 sg13g2_a22oi_1 _4027_ (.Y(_1115_),
    .B1(_0927_),
    .B2(net772),
    .A2(_0925_),
    .A1(net446));
 sg13g2_o21ai_1 _4028_ (.B1(_1115_),
    .Y(_0056_),
    .A1(_0853_),
    .A2(_1114_));
 sg13g2_nor2_2 _4029_ (.A(_0767_),
    .B(_0773_),
    .Y(_1116_));
 sg13g2_mux2_1 _4030_ (.A0(net782),
    .A1(net474),
    .S(_1116_),
    .X(_0057_));
 sg13g2_mux2_1 _4031_ (.A0(net806),
    .A1(net462),
    .S(_1116_),
    .X(_0058_));
 sg13g2_mux2_1 _4032_ (.A0(net800),
    .A1(net456),
    .S(_1116_),
    .X(_0059_));
 sg13g2_mux2_1 _4033_ (.A0(net718),
    .A1(net443),
    .S(_1116_),
    .X(_0060_));
 sg13g2_nor3_2 _4034_ (.A(net552),
    .B(net534),
    .C(_0535_),
    .Y(_1117_));
 sg13g2_nand2_2 _4035_ (.Y(_1118_),
    .A(net515),
    .B(_0536_));
 sg13g2_nor2_2 _4036_ (.A(_0763_),
    .B(_1118_),
    .Y(_1119_));
 sg13g2_nand2_1 _4037_ (.Y(_1120_),
    .A(net480),
    .B(_1119_));
 sg13g2_o21ai_1 _4038_ (.B1(_1120_),
    .Y(_0061_),
    .A1(_2098_),
    .A2(_1119_));
 sg13g2_nand2_1 _4039_ (.Y(_1121_),
    .A(net469),
    .B(_1119_));
 sg13g2_o21ai_1 _4040_ (.B1(_1121_),
    .Y(_0062_),
    .A1(_2100_),
    .A2(_1119_));
 sg13g2_nand2_1 _4041_ (.Y(_1122_),
    .A(net458),
    .B(_1119_));
 sg13g2_o21ai_1 _4042_ (.B1(_1122_),
    .Y(_0063_),
    .A1(_2103_),
    .A2(_1119_));
 sg13g2_mux2_1 _4043_ (.A0(net775),
    .A1(net447),
    .S(_1119_),
    .X(_0064_));
 sg13g2_nand2_2 _4044_ (.Y(_1123_),
    .A(_0766_),
    .B(_0846_));
 sg13g2_mux2_1 _4045_ (.A0(net479),
    .A1(net735),
    .S(_1123_),
    .X(_0065_));
 sg13g2_mux2_1 _4046_ (.A0(net467),
    .A1(net827),
    .S(_1123_),
    .X(_0066_));
 sg13g2_mux2_1 _4047_ (.A0(net457),
    .A1(net849),
    .S(_1123_),
    .X(_0067_));
 sg13g2_mux2_1 _4048_ (.A0(net449),
    .A1(net828),
    .S(_1123_),
    .X(_0068_));
 sg13g2_nor2_2 _4049_ (.A(_0759_),
    .B(_0924_),
    .Y(_1124_));
 sg13g2_mux2_1 _4050_ (.A0(net427),
    .A1(net477),
    .S(_1124_),
    .X(_0069_));
 sg13g2_mux2_1 _4051_ (.A0(net600),
    .A1(net466),
    .S(_1124_),
    .X(_0070_));
 sg13g2_mux2_1 _4052_ (.A0(net626),
    .A1(net455),
    .S(_1124_),
    .X(_0071_));
 sg13g2_mux2_1 _4053_ (.A0(net616),
    .A1(net446),
    .S(_1124_),
    .X(_0072_));
 sg13g2_nand2_2 _4054_ (.Y(_1125_),
    .A(_0766_),
    .B(_0769_));
 sg13g2_mux2_1 _4055_ (.A0(net472),
    .A1(net826),
    .S(_1125_),
    .X(_0073_));
 sg13g2_mux2_1 _4056_ (.A0(net462),
    .A1(net788),
    .S(_1125_),
    .X(_0074_));
 sg13g2_mux2_1 _4057_ (.A0(net456),
    .A1(net793),
    .S(_1125_),
    .X(_0075_));
 sg13g2_mux2_1 _4058_ (.A0(net443),
    .A1(net760),
    .S(_1125_),
    .X(_0076_));
 sg13g2_nand2_2 _4059_ (.Y(_1126_),
    .A(_0537_),
    .B(_0762_));
 sg13g2_mux2_1 _4060_ (.A0(net480),
    .A1(net846),
    .S(_1126_),
    .X(_0077_));
 sg13g2_mux2_1 _4061_ (.A0(net468),
    .A1(net815),
    .S(_1126_),
    .X(_0078_));
 sg13g2_mux2_1 _4062_ (.A0(net458),
    .A1(net848),
    .S(_1126_),
    .X(_0079_));
 sg13g2_mux2_1 _4063_ (.A0(net448),
    .A1(net845),
    .S(_1126_),
    .X(_0080_));
 sg13g2_nor2_2 _4064_ (.A(_0842_),
    .B(_0924_),
    .Y(_1127_));
 sg13g2_mux2_1 _4065_ (.A0(net426),
    .A1(net477),
    .S(_1127_),
    .X(_0081_));
 sg13g2_mux2_1 _4066_ (.A0(net582),
    .A1(net465),
    .S(_1127_),
    .X(_0082_));
 sg13g2_mux2_1 _4067_ (.A0(net431),
    .A1(net454),
    .S(_1127_),
    .X(_0083_));
 sg13g2_mux2_1 _4068_ (.A0(net418),
    .A1(net444),
    .S(_1127_),
    .X(_0084_));
 sg13g2_nand2_2 _4069_ (.Y(_1128_),
    .A(_0766_),
    .B(_0841_));
 sg13g2_mux2_1 _4070_ (.A0(net479),
    .A1(net690),
    .S(_1128_),
    .X(_0085_));
 sg13g2_mux2_1 _4071_ (.A0(net467),
    .A1(net780),
    .S(_1128_),
    .X(_0086_));
 sg13g2_mux2_1 _4072_ (.A0(net457),
    .A1(net812),
    .S(_1128_),
    .X(_0087_));
 sg13g2_mux2_1 _4073_ (.A0(net449),
    .A1(net777),
    .S(_1128_),
    .X(_0088_));
 sg13g2_nand2_2 _4074_ (.Y(_1129_),
    .A(_0758_),
    .B(_0766_));
 sg13g2_mux2_1 _4075_ (.A0(net479),
    .A1(net737),
    .S(_1129_),
    .X(_0089_));
 sg13g2_mux2_1 _4076_ (.A0(net467),
    .A1(net799),
    .S(_1129_),
    .X(_0090_));
 sg13g2_mux2_1 _4077_ (.A0(net457),
    .A1(net811),
    .S(_1129_),
    .X(_0091_));
 sg13g2_mux2_1 _4078_ (.A0(net443),
    .A1(net743),
    .S(_1129_),
    .X(_0092_));
 sg13g2_nor2_2 _4079_ (.A(_0763_),
    .B(_0847_),
    .Y(_1130_));
 sg13g2_mux2_1 _4080_ (.A0(net783),
    .A1(net480),
    .S(_1130_),
    .X(_0093_));
 sg13g2_mux2_1 _4081_ (.A0(net787),
    .A1(net468),
    .S(_1130_),
    .X(_0094_));
 sg13g2_mux2_1 _4082_ (.A0(net747),
    .A1(net459),
    .S(_1130_),
    .X(_0095_));
 sg13g2_mux2_1 _4083_ (.A0(net823),
    .A1(net447),
    .S(_1130_),
    .X(_0096_));
 sg13g2_nor2_2 _4084_ (.A(_0763_),
    .B(_0773_),
    .Y(_1131_));
 sg13g2_mux2_1 _4085_ (.A0(net713),
    .A1(net480),
    .S(_1131_),
    .X(_0097_));
 sg13g2_mux2_1 _4086_ (.A0(net727),
    .A1(net468),
    .S(_1131_),
    .X(_0098_));
 sg13g2_mux2_1 _4087_ (.A0(net750),
    .A1(net459),
    .S(_1131_),
    .X(_0099_));
 sg13g2_mux2_1 _4088_ (.A0(net746),
    .A1(net447),
    .S(_1131_),
    .X(_0100_));
 sg13g2_nand3_1 _4089_ (.B(_0533_),
    .C(_0772_),
    .A(net517),
    .Y(_1132_));
 sg13g2_nor2_2 _4090_ (.A(_0924_),
    .B(_1132_),
    .Y(_1133_));
 sg13g2_mux2_1 _4091_ (.A0(net781),
    .A1(net477),
    .S(_1133_),
    .X(_0101_));
 sg13g2_mux2_1 _4092_ (.A0(net803),
    .A1(net465),
    .S(_1133_),
    .X(_0102_));
 sg13g2_mux2_1 _4093_ (.A0(net814),
    .A1(net455),
    .S(_1133_),
    .X(_0103_));
 sg13g2_mux2_1 _4094_ (.A0(net744),
    .A1(net446),
    .S(_1133_),
    .X(_0104_));
 sg13g2_nand2_2 _4095_ (.Y(_1134_),
    .A(_0762_),
    .B(_0841_));
 sg13g2_mux2_1 _4096_ (.A0(net480),
    .A1(net837),
    .S(_1134_),
    .X(_0105_));
 sg13g2_mux2_1 _4097_ (.A0(net468),
    .A1(net836),
    .S(_1134_),
    .X(_0106_));
 sg13g2_mux2_1 _4098_ (.A0(net458),
    .A1(net807),
    .S(_1134_),
    .X(_0107_));
 sg13g2_mux2_1 _4099_ (.A0(net448),
    .A1(net758),
    .S(_1134_),
    .X(_0108_));
 sg13g2_nor2_2 _4100_ (.A(_0763_),
    .B(_0770_),
    .Y(_1135_));
 sg13g2_mux2_1 _4101_ (.A0(net797),
    .A1(net480),
    .S(_1135_),
    .X(_0109_));
 sg13g2_mux2_1 _4102_ (.A0(net722),
    .A1(net468),
    .S(_1135_),
    .X(_0110_));
 sg13g2_mux2_1 _4103_ (.A0(net841),
    .A1(net459),
    .S(_1135_),
    .X(_0111_));
 sg13g2_mux2_1 _4104_ (.A0(net786),
    .A1(net447),
    .S(_1135_),
    .X(_0112_));
 sg13g2_nor2_1 _4105_ (.A(_0773_),
    .B(_0924_),
    .Y(_1136_));
 sg13g2_o21ai_1 _4106_ (.B1(_1136_),
    .Y(_1137_),
    .A1(_0533_),
    .A2(_0852_));
 sg13g2_nor2_1 _4107_ (.A(net477),
    .B(_1137_),
    .Y(_1138_));
 sg13g2_a21oi_1 _4108_ (.A1(_2089_),
    .A2(_1137_),
    .Y(_0113_),
    .B1(_1138_));
 sg13g2_nor2_1 _4109_ (.A(net465),
    .B(_1137_),
    .Y(_1139_));
 sg13g2_a21oi_1 _4110_ (.A1(_2088_),
    .A2(_1137_),
    .Y(_0114_),
    .B1(_1139_));
 sg13g2_nor2_1 _4111_ (.A(net455),
    .B(_1137_),
    .Y(_1140_));
 sg13g2_a21oi_1 _4112_ (.A1(_2087_),
    .A2(_1137_),
    .Y(_0115_),
    .B1(_1140_));
 sg13g2_nor2_1 _4113_ (.A(net446),
    .B(_1137_),
    .Y(_1141_));
 sg13g2_a21oi_1 _4114_ (.A1(_2086_),
    .A2(_1137_),
    .Y(_0116_),
    .B1(_1141_));
 sg13g2_nand2_2 _4115_ (.Y(_1142_),
    .A(_0766_),
    .B(_1117_));
 sg13g2_mux2_1 _4116_ (.A0(net479),
    .A1(net699),
    .S(_1142_),
    .X(_0117_));
 sg13g2_mux2_1 _4117_ (.A0(net467),
    .A1(net824),
    .S(_1142_),
    .X(_0118_));
 sg13g2_nor2_1 _4118_ (.A(net460),
    .B(_1142_),
    .Y(_1143_));
 sg13g2_a21oi_1 _4119_ (.A1(_2104_),
    .A2(_1142_),
    .Y(_0119_),
    .B1(_1143_));
 sg13g2_nor2_1 _4120_ (.A(net449),
    .B(_1142_),
    .Y(_1144_));
 sg13g2_a21oi_1 _4121_ (.A1(_2105_),
    .A2(_1142_),
    .Y(_0120_),
    .B1(_1144_));
 sg13g2_nor2_2 _4122_ (.A(_0767_),
    .B(_1132_),
    .Y(_1145_));
 sg13g2_mux2_1 _4123_ (.A0(net705),
    .A1(net474),
    .S(_1145_),
    .X(_0121_));
 sg13g2_mux2_1 _4124_ (.A0(net792),
    .A1(net462),
    .S(_1145_),
    .X(_0122_));
 sg13g2_mux2_1 _4125_ (.A0(net813),
    .A1(net452),
    .S(_1145_),
    .X(_0123_));
 sg13g2_mux2_1 _4126_ (.A0(net751),
    .A1(net443),
    .S(_1145_),
    .X(_0124_));
 sg13g2_nor2_2 _4127_ (.A(_0773_),
    .B(_0845_),
    .Y(_1146_));
 sg13g2_mux2_1 _4128_ (.A0(net765),
    .A1(net480),
    .S(_1146_),
    .X(_0125_));
 sg13g2_mux2_1 _4129_ (.A0(net757),
    .A1(net468),
    .S(_1146_),
    .X(_0126_));
 sg13g2_mux2_1 _4130_ (.A0(net778),
    .A1(net459),
    .S(_1146_),
    .X(_0127_));
 sg13g2_mux2_1 _4131_ (.A0(net759),
    .A1(net447),
    .S(_1146_),
    .X(_0128_));
 sg13g2_nand4_1 _4132_ (.B(net522),
    .C(net488),
    .A(net527),
    .Y(_1147_),
    .D(_0760_));
 sg13g2_nor2_2 _4133_ (.A(_1132_),
    .B(_1147_),
    .Y(_1148_));
 sg13g2_mux2_1 _4134_ (.A0(net639),
    .A1(net476),
    .S(_1148_),
    .X(_0129_));
 sg13g2_mux2_1 _4135_ (.A0(net624),
    .A1(net464),
    .S(_1148_),
    .X(_0130_));
 sg13g2_mux2_1 _4136_ (.A0(net613),
    .A1(net454),
    .S(_1148_),
    .X(_0131_));
 sg13g2_mux2_1 _4137_ (.A0(net631),
    .A1(net444),
    .S(_1148_),
    .X(_0132_));
 sg13g2_nand2_2 _4138_ (.Y(_1149_),
    .A(_0758_),
    .B(_0844_));
 sg13g2_mux2_1 _4139_ (.A0(net481),
    .A1(net676),
    .S(_1149_),
    .X(_0133_));
 sg13g2_mux2_1 _4140_ (.A0(net469),
    .A1(net748),
    .S(_1149_),
    .X(_0134_));
 sg13g2_mux2_1 _4141_ (.A0(net459),
    .A1(net819),
    .S(_1149_),
    .X(_0135_));
 sg13g2_mux2_1 _4142_ (.A0(net448),
    .A1(net755),
    .S(_1149_),
    .X(_0136_));
 sg13g2_nor2_2 _4143_ (.A(_0847_),
    .B(_0924_),
    .Y(_1150_));
 sg13g2_mux2_1 _4144_ (.A0(net610),
    .A1(net476),
    .S(_1150_),
    .X(_0137_));
 sg13g2_mux2_1 _4145_ (.A0(net416),
    .A1(net465),
    .S(_1150_),
    .X(_0138_));
 sg13g2_mux2_1 _4146_ (.A0(net420),
    .A1(net454),
    .S(_1150_),
    .X(_0139_));
 sg13g2_mux2_1 _4147_ (.A0(net414),
    .A1(net445),
    .S(_1150_),
    .X(_0140_));
 sg13g2_nor2_2 _4148_ (.A(_0538_),
    .B(_0924_),
    .Y(_1151_));
 sg13g2_mux2_1 _4149_ (.A0(net627),
    .A1(net477),
    .S(_1151_),
    .X(_0141_));
 sg13g2_mux2_1 _4150_ (.A0(net649),
    .A1(net465),
    .S(_1151_),
    .X(_0142_));
 sg13g2_mux2_1 _4151_ (.A0(net628),
    .A1(net454),
    .S(_1151_),
    .X(_0143_));
 sg13g2_mux2_1 _4152_ (.A0(net607),
    .A1(net444),
    .S(_1151_),
    .X(_0144_));
 sg13g2_nor2_2 _4153_ (.A(_0924_),
    .B(_1118_),
    .Y(_1152_));
 sg13g2_mux2_1 _4154_ (.A0(net591),
    .A1(net478),
    .S(_1152_),
    .X(_0145_));
 sg13g2_mux2_1 _4155_ (.A0(net602),
    .A1(net466),
    .S(_1152_),
    .X(_0146_));
 sg13g2_mux2_1 _4156_ (.A0(net609),
    .A1(net455),
    .S(_1152_),
    .X(_0147_));
 sg13g2_mux2_1 _4157_ (.A0(net617),
    .A1(net444),
    .S(_1152_),
    .X(_0148_));
 sg13g2_nand3b_1 _4158_ (.B(net578),
    .C(net2),
    .Y(_1153_),
    .A_N(net854));
 sg13g2_o21ai_1 _4159_ (.B1(net484),
    .Y(_0149_),
    .A1(net1),
    .A2(_1153_));
 sg13g2_nor2_2 _4160_ (.A(_0763_),
    .B(_1132_),
    .Y(_1154_));
 sg13g2_mux2_1 _4161_ (.A0(net501),
    .A1(net477),
    .S(_1154_),
    .X(_0150_));
 sg13g2_mux2_1 _4162_ (.A0(net500),
    .A1(net465),
    .S(_1154_),
    .X(_0151_));
 sg13g2_mux2_1 _4163_ (.A0(net839),
    .A1(net455),
    .S(_1154_),
    .X(_0152_));
 sg13g2_mux2_1 _4164_ (.A0(net736),
    .A1(net446),
    .S(_1154_),
    .X(_0153_));
 sg13g2_nand2_2 _4165_ (.Y(_1155_),
    .A(_0540_),
    .B(_0841_));
 sg13g2_mux2_1 _4166_ (.A0(net482),
    .A1(net635),
    .S(_1155_),
    .X(_0154_));
 sg13g2_mux2_1 _4167_ (.A0(net467),
    .A1(net658),
    .S(_1155_),
    .X(_0155_));
 sg13g2_mux2_1 _4168_ (.A0(net457),
    .A1(net779),
    .S(_1155_),
    .X(_0156_));
 sg13g2_mux2_1 _4169_ (.A0(net449),
    .A1(net739),
    .S(_1155_),
    .X(_0157_));
 sg13g2_nand2_2 _4170_ (.Y(_1156_),
    .A(_0540_),
    .B(_0846_));
 sg13g2_mux2_1 _4171_ (.A0(net479),
    .A1(net497),
    .S(_1156_),
    .X(_0158_));
 sg13g2_mux2_1 _4172_ (.A0(net467),
    .A1(net496),
    .S(_1156_),
    .X(_0159_));
 sg13g2_mux2_1 _4173_ (.A0(net457),
    .A1(net830),
    .S(_1156_),
    .X(_0160_));
 sg13g2_mux2_1 _4174_ (.A0(net449),
    .A1(net774),
    .S(_1156_),
    .X(_0161_));
 sg13g2_nand2_2 _4175_ (.Y(_1157_),
    .A(_0778_),
    .B(_0846_));
 sg13g2_mux2_1 _4176_ (.A0(net472),
    .A1(net663),
    .S(_1157_),
    .X(_0162_));
 sg13g2_mux2_1 _4177_ (.A0(net461),
    .A1(net650),
    .S(_1157_),
    .X(_0163_));
 sg13g2_mux2_1 _4178_ (.A0(net451),
    .A1(net648),
    .S(_1157_),
    .X(_0164_));
 sg13g2_mux2_1 _4179_ (.A0(net442),
    .A1(net634),
    .S(_1157_),
    .X(_0165_));
 sg13g2_nand2_2 _4180_ (.Y(_1158_),
    .A(_0537_),
    .B(_0778_));
 sg13g2_mux2_1 _4181_ (.A0(net472),
    .A1(net646),
    .S(_1158_),
    .X(_0166_));
 sg13g2_mux2_1 _4182_ (.A0(net461),
    .A1(net662),
    .S(_1158_),
    .X(_0167_));
 sg13g2_mux2_1 _4183_ (.A0(net451),
    .A1(net672),
    .S(_1158_),
    .X(_0168_));
 sg13g2_mux2_1 _4184_ (.A0(net442),
    .A1(net667),
    .S(_1158_),
    .X(_0169_));
 sg13g2_nand2_2 _4185_ (.Y(_1159_),
    .A(_0778_),
    .B(_1117_));
 sg13g2_mux2_1 _4186_ (.A0(net472),
    .A1(net668),
    .S(_1159_),
    .X(_0170_));
 sg13g2_mux2_1 _4187_ (.A0(net461),
    .A1(net671),
    .S(_1159_),
    .X(_0171_));
 sg13g2_mux2_1 _4188_ (.A0(net451),
    .A1(net652),
    .S(_1159_),
    .X(_0172_));
 sg13g2_mux2_1 _4189_ (.A0(net442),
    .A1(net665),
    .S(_1159_),
    .X(_0173_));
 sg13g2_nand2_2 _4190_ (.Y(_1160_),
    .A(_0537_),
    .B(_0844_));
 sg13g2_mux2_1 _4191_ (.A0(net481),
    .A1(net495),
    .S(_1160_),
    .X(_0174_));
 sg13g2_mux2_1 _4192_ (.A0(net469),
    .A1(net494),
    .S(_1160_),
    .X(_0175_));
 sg13g2_mux2_1 _4193_ (.A0(net458),
    .A1(net832),
    .S(_1160_),
    .X(_0176_));
 sg13g2_mux2_1 _4194_ (.A0(net448),
    .A1(net805),
    .S(_1160_),
    .X(_0177_));
 sg13g2_nand2_2 _4195_ (.Y(_1161_),
    .A(_0769_),
    .B(_0778_));
 sg13g2_mux2_1 _4196_ (.A0(net473),
    .A1(net637),
    .S(_1161_),
    .X(_0178_));
 sg13g2_mux2_1 _4197_ (.A0(net461),
    .A1(net645),
    .S(_1161_),
    .X(_0179_));
 sg13g2_mux2_1 _4198_ (.A0(net452),
    .A1(net660),
    .S(_1161_),
    .X(_0180_));
 sg13g2_mux2_1 _4199_ (.A0(net441),
    .A1(net647),
    .S(_1161_),
    .X(_0181_));
 sg13g2_nor2b_2 _4200_ (.A(_0773_),
    .B_N(_0778_),
    .Y(_1162_));
 sg13g2_mux2_1 _4201_ (.A0(net581),
    .A1(net472),
    .S(_1162_),
    .X(_0182_));
 sg13g2_mux2_1 _4202_ (.A0(net423),
    .A1(net461),
    .S(_1162_),
    .X(_0183_));
 sg13g2_mux2_1 _4203_ (.A0(net625),
    .A1(net452),
    .S(_1162_),
    .X(_0184_));
 sg13g2_mux2_1 _4204_ (.A0(net605),
    .A1(net441),
    .S(_1162_),
    .X(_0185_));
 sg13g2_nor3_2 _4205_ (.A(net502),
    .B(_0774_),
    .C(_1132_),
    .Y(_1163_));
 sg13g2_mux2_1 _4206_ (.A0(net615),
    .A1(net472),
    .S(_1163_),
    .X(_0186_));
 sg13g2_mux2_1 _4207_ (.A0(net435),
    .A1(net461),
    .S(_1163_),
    .X(_0187_));
 sg13g2_mux2_1 _4208_ (.A0(net606),
    .A1(net451),
    .S(_1163_),
    .X(_0188_));
 sg13g2_mux2_1 _4209_ (.A0(net611),
    .A1(net441),
    .S(_1163_),
    .X(_0189_));
 sg13g2_nand2_2 _4210_ (.Y(_1164_),
    .A(_0775_),
    .B(_0841_));
 sg13g2_mux2_1 _4211_ (.A0(net473),
    .A1(net670),
    .S(_1164_),
    .X(_0190_));
 sg13g2_mux2_1 _4212_ (.A0(net471),
    .A1(net656),
    .S(_1164_),
    .X(_0191_));
 sg13g2_mux2_1 _4213_ (.A0(net451),
    .A1(net659),
    .S(_1164_),
    .X(_0192_));
 sg13g2_mux2_1 _4214_ (.A0(net442),
    .A1(net666),
    .S(_1164_),
    .X(_0193_));
 sg13g2_nor2_2 _4215_ (.A(_0776_),
    .B(_0847_),
    .Y(_1165_));
 sg13g2_mux2_1 _4216_ (.A0(net415),
    .A1(net473),
    .S(_1165_),
    .X(_0194_));
 sg13g2_mux2_1 _4217_ (.A0(net583),
    .A1(net463),
    .S(_1165_),
    .X(_0195_));
 sg13g2_mux2_1 _4218_ (.A0(net584),
    .A1(net451),
    .S(_1165_),
    .X(_0196_));
 sg13g2_mux2_1 _4219_ (.A0(net421),
    .A1(net442),
    .S(_1165_),
    .X(_0197_));
 sg13g2_nand2_2 _4220_ (.Y(_1166_),
    .A(_0537_),
    .B(_0775_));
 sg13g2_mux2_1 _4221_ (.A0(net477),
    .A1(net643),
    .S(_1166_),
    .X(_0198_));
 sg13g2_mux2_1 _4222_ (.A0(net465),
    .A1(net657),
    .S(_1166_),
    .X(_0199_));
 sg13g2_mux2_1 _4223_ (.A0(net456),
    .A1(net655),
    .S(_1166_),
    .X(_0200_));
 sg13g2_mux2_1 _4224_ (.A0(net446),
    .A1(net654),
    .S(_1166_),
    .X(_0201_));
 sg13g2_nor2_2 _4225_ (.A(_0776_),
    .B(_1118_),
    .Y(_1167_));
 sg13g2_mux2_1 _4226_ (.A0(net434),
    .A1(net475),
    .S(_1167_),
    .X(_0202_));
 sg13g2_nand2_1 _4227_ (.Y(_1168_),
    .A(net463),
    .B(_1167_));
 sg13g2_o21ai_1 _4228_ (.B1(_1168_),
    .Y(_0203_),
    .A1(_2101_),
    .A2(_1167_));
 sg13g2_mux2_1 _4229_ (.A0(net588),
    .A1(net453),
    .S(_1167_),
    .X(_0204_));
 sg13g2_mux2_1 _4230_ (.A0(net590),
    .A1(net445),
    .S(_1167_),
    .X(_0205_));
 sg13g2_nand2_2 _4231_ (.Y(_1169_),
    .A(_0758_),
    .B(_0775_));
 sg13g2_mux2_1 _4232_ (.A0(net475),
    .A1(net661),
    .S(_1169_),
    .X(_0206_));
 sg13g2_mux2_1 _4233_ (.A0(net463),
    .A1(net669),
    .S(_1169_),
    .X(_0207_));
 sg13g2_mux2_1 _4234_ (.A0(net453),
    .A1(net640),
    .S(_1169_),
    .X(_0208_));
 sg13g2_mux2_1 _4235_ (.A0(net441),
    .A1(net644),
    .S(_1169_),
    .X(_0209_));
 sg13g2_nor2_2 _4236_ (.A(_0770_),
    .B(_0776_),
    .Y(_1170_));
 sg13g2_mux2_1 _4237_ (.A0(net428),
    .A1(net475),
    .S(_1170_),
    .X(_0210_));
 sg13g2_mux2_1 _4238_ (.A0(net440),
    .A1(net463),
    .S(_1170_),
    .X(_0211_));
 sg13g2_mux2_1 _4239_ (.A0(net589),
    .A1(net453),
    .S(_1170_),
    .X(_0212_));
 sg13g2_mux2_1 _4240_ (.A0(net438),
    .A1(net441),
    .S(_1170_),
    .X(_0213_));
 sg13g2_nor2_2 _4241_ (.A(_0845_),
    .B(_1118_),
    .Y(_1171_));
 sg13g2_nand2_1 _4242_ (.Y(_1172_),
    .A(net481),
    .B(_1171_));
 sg13g2_o21ai_1 _4243_ (.B1(_1172_),
    .Y(_0214_),
    .A1(_2096_),
    .A2(_1171_));
 sg13g2_nand2_1 _4244_ (.Y(_1173_),
    .A(net469),
    .B(_1171_));
 sg13g2_o21ai_1 _4245_ (.B1(_1173_),
    .Y(_0215_),
    .A1(_2099_),
    .A2(_1171_));
 sg13g2_mux2_1 _4246_ (.A0(net768),
    .A1(net458),
    .S(_1171_),
    .X(_0216_));
 sg13g2_mux2_1 _4247_ (.A0(net742),
    .A1(net447),
    .S(_1171_),
    .X(_0217_));
 sg13g2_nor2_2 _4248_ (.A(_0776_),
    .B(_1132_),
    .Y(_1174_));
 sg13g2_mux2_1 _4249_ (.A0(net619),
    .A1(net475),
    .S(_1174_),
    .X(_0218_));
 sg13g2_mux2_1 _4250_ (.A0(net596),
    .A1(net463),
    .S(_1174_),
    .X(_0219_));
 sg13g2_mux2_1 _4251_ (.A0(net586),
    .A1(net453),
    .S(_1174_),
    .X(_0220_));
 sg13g2_mux2_1 _4252_ (.A0(net614),
    .A1(net441),
    .S(_1174_),
    .X(_0221_));
 sg13g2_nor2_2 _4253_ (.A(_0842_),
    .B(_1147_),
    .Y(_1175_));
 sg13g2_mux2_1 _4254_ (.A0(net597),
    .A1(net476),
    .S(_1175_),
    .X(_0222_));
 sg13g2_mux2_1 _4255_ (.A0(net439),
    .A1(net464),
    .S(_1175_),
    .X(_0223_));
 sg13g2_mux2_1 _4256_ (.A0(net595),
    .A1(net453),
    .S(_1175_),
    .X(_0224_));
 sg13g2_mux2_1 _4257_ (.A0(net594),
    .A1(net445),
    .S(_1175_),
    .X(_0225_));
 sg13g2_nor2_2 _4258_ (.A(_0847_),
    .B(_1147_),
    .Y(_1176_));
 sg13g2_mux2_1 _4259_ (.A0(net417),
    .A1(net475),
    .S(_1176_),
    .X(_0226_));
 sg13g2_mux2_1 _4260_ (.A0(net433),
    .A1(net463),
    .S(_1176_),
    .X(_0227_));
 sg13g2_mux2_1 _4261_ (.A0(net620),
    .A1(net453),
    .S(_1176_),
    .X(_0228_));
 sg13g2_mux2_1 _4262_ (.A0(net422),
    .A1(net445),
    .S(_1176_),
    .X(_0229_));
 sg13g2_nor2_2 _4263_ (.A(_0538_),
    .B(_1147_),
    .Y(_1177_));
 sg13g2_mux2_1 _4264_ (.A0(net592),
    .A1(net475),
    .S(_1177_),
    .X(_0230_));
 sg13g2_mux2_1 _4265_ (.A0(net585),
    .A1(net464),
    .S(_1177_),
    .X(_0231_));
 sg13g2_mux2_1 _4266_ (.A0(net621),
    .A1(net454),
    .S(_1177_),
    .X(_0232_));
 sg13g2_mux2_1 _4267_ (.A0(net598),
    .A1(net444),
    .S(_1177_),
    .X(_0233_));
 sg13g2_nor2_2 _4268_ (.A(_1118_),
    .B(_1147_),
    .Y(_1178_));
 sg13g2_mux2_1 _4269_ (.A0(net430),
    .A1(net475),
    .S(_1178_),
    .X(_0234_));
 sg13g2_mux2_1 _4270_ (.A0(net593),
    .A1(net463),
    .S(_1178_),
    .X(_0235_));
 sg13g2_mux2_1 _4271_ (.A0(net603),
    .A1(net453),
    .S(_1178_),
    .X(_0236_));
 sg13g2_mux2_1 _4272_ (.A0(net612),
    .A1(net445),
    .S(_1178_),
    .X(_0237_));
 sg13g2_nor2_2 _4273_ (.A(_0759_),
    .B(_1147_),
    .Y(_1179_));
 sg13g2_mux2_1 _4274_ (.A0(net436),
    .A1(net476),
    .S(_1179_),
    .X(_0238_));
 sg13g2_mux2_1 _4275_ (.A0(net604),
    .A1(net464),
    .S(_1179_),
    .X(_0239_));
 sg13g2_mux2_1 _4276_ (.A0(net587),
    .A1(net454),
    .S(_1179_),
    .X(_0240_));
 sg13g2_mux2_1 _4277_ (.A0(net437),
    .A1(net444),
    .S(_1179_),
    .X(_0241_));
 sg13g2_nor2_2 _4278_ (.A(_0770_),
    .B(_1147_),
    .Y(_1180_));
 sg13g2_mux2_1 _4279_ (.A0(net432),
    .A1(net476),
    .S(_1180_),
    .X(_0242_));
 sg13g2_mux2_1 _4280_ (.A0(net429),
    .A1(net464),
    .S(_1180_),
    .X(_0243_));
 sg13g2_mux2_1 _4281_ (.A0(net599),
    .A1(net454),
    .S(_1180_),
    .X(_0244_));
 sg13g2_mux2_1 _4282_ (.A0(net419),
    .A1(net444),
    .S(_1180_),
    .X(_0245_));
 sg13g2_nor2_2 _4283_ (.A(_0845_),
    .B(_1132_),
    .Y(_1181_));
 sg13g2_mux2_1 _4284_ (.A0(net804),
    .A1(net480),
    .S(_1181_),
    .X(_0246_));
 sg13g2_mux2_1 _4285_ (.A0(net771),
    .A1(net468),
    .S(_1181_),
    .X(_0247_));
 sg13g2_mux2_1 _4286_ (.A0(net493),
    .A1(net459),
    .S(_1181_),
    .X(_0248_));
 sg13g2_mux2_1 _4287_ (.A0(net492),
    .A1(net447),
    .S(_1181_),
    .X(_0249_));
 sg13g2_nor2_2 _4288_ (.A(_0773_),
    .B(_1147_),
    .Y(_1182_));
 sg13g2_mux2_1 _4289_ (.A0(net623),
    .A1(net476),
    .S(_1182_),
    .X(_0250_));
 sg13g2_mux2_1 _4290_ (.A0(net622),
    .A1(net464),
    .S(_1182_),
    .X(_0251_));
 sg13g2_mux2_1 _4291_ (.A0(net630),
    .A1(net454),
    .S(_1182_),
    .X(_0252_));
 sg13g2_mux2_1 _4292_ (.A0(net601),
    .A1(net444),
    .S(_1182_),
    .X(_0253_));
 sg13g2_nor2_2 _4293_ (.A(_0541_),
    .B(_1132_),
    .Y(_1183_));
 sg13g2_mux2_1 _4294_ (.A0(net491),
    .A1(net474),
    .S(_1183_),
    .X(_0254_));
 sg13g2_mux2_1 _4295_ (.A0(net490),
    .A1(net462),
    .S(_1183_),
    .X(_0255_));
 sg13g2_mux2_1 _4296_ (.A0(net801),
    .A1(net452),
    .S(_1183_),
    .X(_0256_));
 sg13g2_mux2_1 _4297_ (.A0(net712),
    .A1(net443),
    .S(_1183_),
    .X(_0257_));
 sg13g2_nand2_2 _4298_ (.Y(_1184_),
    .A(_0540_),
    .B(_1117_));
 sg13g2_nor2_1 _4299_ (.A(net479),
    .B(_1184_),
    .Y(_1185_));
 sg13g2_a21oi_1 _4300_ (.A1(_2097_),
    .A2(_1184_),
    .Y(_0258_),
    .B1(_1185_));
 sg13g2_mux2_1 _4301_ (.A0(net470),
    .A1(net790),
    .S(_1184_),
    .X(_0259_));
 sg13g2_mux2_1 _4302_ (.A0(net457),
    .A1(net834),
    .S(_1184_),
    .X(_0260_));
 sg13g2_mux2_1 _4303_ (.A0(net449),
    .A1(net785),
    .S(_1184_),
    .X(_0261_));
 sg13g2_nor2_2 _4304_ (.A(_0541_),
    .B(_0773_),
    .Y(_1186_));
 sg13g2_mux2_1 _4305_ (.A0(net697),
    .A1(net474),
    .S(_1186_),
    .X(_0262_));
 sg13g2_mux2_1 _4306_ (.A0(net753),
    .A1(net462),
    .S(_1186_),
    .X(_0263_));
 sg13g2_mux2_1 _4307_ (.A0(net740),
    .A1(net452),
    .S(_1186_),
    .X(_0264_));
 sg13g2_mux2_1 _4308_ (.A0(net720),
    .A1(net443),
    .S(_1186_),
    .X(_0265_));
 sg13g2_nor2_1 _4309_ (.A(\mem[0][1] ),
    .B(\mem[0][0] ),
    .Y(_1187_));
 sg13g2_or2_2 _4310_ (.X(_1188_),
    .B(\mem[0][0] ),
    .A(\mem[0][1] ));
 sg13g2_nor2_2 _4311_ (.A(net493),
    .B(net492),
    .Y(_1189_));
 sg13g2_nor4_2 _4312_ (.A(net493),
    .B(net492),
    .C(net486),
    .Y(_1190_),
    .D(_1188_));
 sg13g2_nand3_1 _4313_ (.B(_1187_),
    .C(_1189_),
    .A(_0781_),
    .Y(_1191_));
 sg13g2_and3_1 _4314_ (.X(_0266_),
    .A(net501),
    .B(net781),
    .C(net483));
 sg13g2_and4_1 _4315_ (.A(net501),
    .B(\mem[32][0] ),
    .C(net500),
    .D(\mem[32][1] ),
    .X(_1192_));
 sg13g2_a22oi_1 _4316_ (.Y(_1193_),
    .B1(net803),
    .B2(net501),
    .A2(net500),
    .A1(net781));
 sg13g2_nor3_1 _4317_ (.A(_1191_),
    .B(_1192_),
    .C(_1193_),
    .Y(_0267_));
 sg13g2_a22oi_1 _4318_ (.Y(_1194_),
    .B1(\mem[32][2] ),
    .B2(net501),
    .A2(\mem[32][1] ),
    .A1(net500));
 sg13g2_nand4_1 _4319_ (.B(net500),
    .C(\mem[32][1] ),
    .A(net501),
    .Y(_1195_),
    .D(\mem[32][2] ));
 sg13g2_nor2b_1 _4320_ (.A(_1194_),
    .B_N(_1195_),
    .Y(_1196_));
 sg13g2_and3_1 _4321_ (.X(_1197_),
    .A(\mem[32][0] ),
    .B(\mem[16][2] ),
    .C(_1196_));
 sg13g2_a21oi_1 _4322_ (.A1(\mem[32][0] ),
    .A2(\mem[16][2] ),
    .Y(_1198_),
    .B1(_1196_));
 sg13g2_nor2_1 _4323_ (.A(_1197_),
    .B(_1198_),
    .Y(_1199_));
 sg13g2_and2_1 _4324_ (.A(_1192_),
    .B(_1199_),
    .X(_1200_));
 sg13g2_o21ai_1 _4325_ (.B1(net483),
    .Y(_1201_),
    .A1(_1192_),
    .A2(_1199_));
 sg13g2_nor2_1 _4326_ (.A(_1200_),
    .B(_1201_),
    .Y(_0268_));
 sg13g2_and2_1 _4327_ (.A(\mem[32][0] ),
    .B(\mem[16][3] ),
    .X(_1202_));
 sg13g2_nand2_1 _4328_ (.Y(_1203_),
    .A(\mem[32][1] ),
    .B(\mem[16][2] ));
 sg13g2_nand2_1 _4329_ (.Y(_1204_),
    .A(net500),
    .B(\mem[32][3] ));
 sg13g2_and4_1 _4330_ (.A(net501),
    .B(net500),
    .C(\mem[32][2] ),
    .D(\mem[32][3] ),
    .X(_1205_));
 sg13g2_a22oi_1 _4331_ (.Y(_1206_),
    .B1(\mem[32][3] ),
    .B2(net501),
    .A2(\mem[32][2] ),
    .A1(net500));
 sg13g2_nor3_1 _4332_ (.A(_1203_),
    .B(_1205_),
    .C(_1206_),
    .Y(_1207_));
 sg13g2_o21ai_1 _4333_ (.B1(_1203_),
    .Y(_1208_),
    .A1(_1205_),
    .A2(_1206_));
 sg13g2_nor2b_1 _4334_ (.A(_1207_),
    .B_N(_1208_),
    .Y(_1209_));
 sg13g2_nor2b_1 _4335_ (.A(_1195_),
    .B_N(_1209_),
    .Y(_1210_));
 sg13g2_xnor2_1 _4336_ (.Y(_1211_),
    .A(_1195_),
    .B(_1209_));
 sg13g2_xor2_1 _4337_ (.B(_1211_),
    .A(_1202_),
    .X(_1212_));
 sg13g2_and2_1 _4338_ (.A(_1197_),
    .B(_1212_),
    .X(_1213_));
 sg13g2_xor2_1 _4339_ (.B(_1212_),
    .A(_1197_),
    .X(_1214_));
 sg13g2_o21ai_1 _4340_ (.B1(net483),
    .Y(_1215_),
    .A1(_1200_),
    .A2(_1214_));
 sg13g2_a21oi_2 _4341_ (.B1(_1215_),
    .Y(_0269_),
    .A2(_1214_),
    .A1(_1200_));
 sg13g2_a21o_1 _4342_ (.A2(_1214_),
    .A1(_1200_),
    .B1(_1213_),
    .X(_1216_));
 sg13g2_or2_1 _4343_ (.X(_1217_),
    .B(_1207_),
    .A(_1205_));
 sg13g2_nand2_1 _4344_ (.Y(_1218_),
    .A(\mem[32][1] ),
    .B(\mem[16][3] ));
 sg13g2_nand2_1 _4345_ (.Y(_1219_),
    .A(\mem[16][2] ),
    .B(\mem[32][3] ));
 sg13g2_nand2_2 _4346_ (.Y(_1220_),
    .A(\mem[16][2] ),
    .B(\mem[32][2] ));
 sg13g2_xor2_1 _4347_ (.B(_1220_),
    .A(_1204_),
    .X(_1221_));
 sg13g2_nand2b_1 _4348_ (.Y(_1222_),
    .B(_1221_),
    .A_N(_1218_));
 sg13g2_xnor2_1 _4349_ (.Y(_1223_),
    .A(_1218_),
    .B(_1221_));
 sg13g2_nand2_1 _4350_ (.Y(_1224_),
    .A(_1217_),
    .B(_1223_));
 sg13g2_xor2_1 _4351_ (.B(_1223_),
    .A(_1217_),
    .X(_1225_));
 sg13g2_a21oi_1 _4352_ (.A1(_1202_),
    .A2(_1211_),
    .Y(_1226_),
    .B1(_1210_));
 sg13g2_nand2b_1 _4353_ (.Y(_1227_),
    .B(_1225_),
    .A_N(_1226_));
 sg13g2_xnor2_1 _4354_ (.Y(_1228_),
    .A(_1225_),
    .B(_1226_));
 sg13g2_or2_1 _4355_ (.X(_1229_),
    .B(_1228_),
    .A(_1216_));
 sg13g2_nand2_1 _4356_ (.Y(_1230_),
    .A(_1216_),
    .B(_1228_));
 sg13g2_and3_2 _4357_ (.X(_0270_),
    .A(net483),
    .B(_1229_),
    .C(_1230_));
 sg13g2_nor2b_1 _4358_ (.A(_1216_),
    .B_N(_1227_),
    .Y(_1231_));
 sg13g2_o21ai_1 _4359_ (.B1(_1222_),
    .Y(_1232_),
    .A1(_1204_),
    .A2(_1220_));
 sg13g2_nand2_1 _4360_ (.Y(_1233_),
    .A(\mem[32][2] ),
    .B(\mem[16][3] ));
 sg13g2_nand2_1 _4361_ (.Y(_1234_),
    .A(\mem[16][3] ),
    .B(\mem[32][3] ));
 sg13g2_xor2_1 _4362_ (.B(_1233_),
    .A(_1219_),
    .X(_1235_));
 sg13g2_nand2_1 _4363_ (.Y(_1236_),
    .A(_1232_),
    .B(_1235_));
 sg13g2_xnor2_1 _4364_ (.Y(_1237_),
    .A(_1232_),
    .B(_1235_));
 sg13g2_xnor2_1 _4365_ (.Y(_1238_),
    .A(_1224_),
    .B(_1237_));
 sg13g2_and3_1 _4366_ (.X(_1239_),
    .A(_1227_),
    .B(_1230_),
    .C(_1238_));
 sg13g2_a21oi_1 _4367_ (.A1(_1227_),
    .A2(_1230_),
    .Y(_1240_),
    .B1(_1238_));
 sg13g2_nor3_2 _4368_ (.A(_1191_),
    .B(_1239_),
    .C(_1240_),
    .Y(_0271_));
 sg13g2_a21oi_1 _4369_ (.A1(_1224_),
    .A2(_1231_),
    .Y(_1241_),
    .B1(_1237_));
 sg13g2_nand2b_1 _4370_ (.Y(_1242_),
    .B(_1220_),
    .A_N(_1234_));
 sg13g2_xor2_1 _4371_ (.B(_1242_),
    .A(_1236_),
    .X(_1243_));
 sg13g2_or2_1 _4372_ (.X(_1244_),
    .B(_1243_),
    .A(_1241_));
 sg13g2_nand2_1 _4373_ (.Y(_1245_),
    .A(_1241_),
    .B(_1243_));
 sg13g2_and3_2 _4374_ (.X(_0272_),
    .A(net483),
    .B(_1244_),
    .C(_1245_));
 sg13g2_a21o_1 _4375_ (.A2(_1236_),
    .A1(_1220_),
    .B1(_1234_),
    .X(_1246_));
 sg13g2_a21oi_2 _4376_ (.B1(_1191_),
    .Y(_0273_),
    .A2(_1246_),
    .A1(_1245_));
 sg13g2_and2_1 _4377_ (.A(net411),
    .B(_0781_),
    .X(_1247_));
 sg13g2_nand2_1 _4378_ (.Y(_1248_),
    .A(net492),
    .B(_0781_));
 sg13g2_nand2_2 _4379_ (.Y(_1249_),
    .A(\mem[0][1] ),
    .B(\mem[0][0] ));
 sg13g2_nor2_2 _4380_ (.A(net486),
    .B(_1249_),
    .Y(_1250_));
 sg13g2_and3_1 _4381_ (.X(_1251_),
    .A(\mem[0][1] ),
    .B(net493),
    .C(_0781_));
 sg13g2_a21oi_2 _4382_ (.B1(_1190_),
    .Y(_1252_),
    .A2(_1251_),
    .A1(net492));
 sg13g2_inv_2 _4383_ (.Y(_1253_),
    .A(_1252_));
 sg13g2_o21ai_1 _4384_ (.B1(_1253_),
    .Y(_1254_),
    .A1(\mem[0][0] ),
    .A2(_1190_));
 sg13g2_nand2_1 _4385_ (.Y(_1255_),
    .A(net499),
    .B(net690));
 sg13g2_nor2_1 _4386_ (.A(_1254_),
    .B(_1255_),
    .Y(_0274_));
 sg13g2_a22oi_1 _4387_ (.Y(_1256_),
    .B1(net780),
    .B2(net499),
    .A2(net498),
    .A1(net690));
 sg13g2_and4_1 _4388_ (.A(net499),
    .B(net802),
    .C(net498),
    .D(\mem[31][1] ),
    .X(_1257_));
 sg13g2_nor3_1 _4389_ (.A(_1254_),
    .B(_1256_),
    .C(_1257_),
    .Y(_0275_));
 sg13g2_a22oi_1 _4390_ (.Y(_1258_),
    .B1(\mem[31][2] ),
    .B2(net499),
    .A2(\mem[31][1] ),
    .A1(net498));
 sg13g2_and4_2 _4391_ (.A(net499),
    .B(net498),
    .C(\mem[31][1] ),
    .D(\mem[31][2] ),
    .X(_1259_));
 sg13g2_nor2_1 _4392_ (.A(_1258_),
    .B(_1259_),
    .Y(_1260_));
 sg13g2_nand2_1 _4393_ (.Y(_1261_),
    .A(\mem[31][0] ),
    .B(\mem[15][2] ));
 sg13g2_nor3_1 _4394_ (.A(_1258_),
    .B(_1259_),
    .C(_1261_),
    .Y(_1262_));
 sg13g2_xnor2_1 _4395_ (.Y(_1263_),
    .A(_1260_),
    .B(_1261_));
 sg13g2_nand2_1 _4396_ (.Y(_1264_),
    .A(_1257_),
    .B(_1263_));
 sg13g2_xnor2_1 _4397_ (.Y(_1265_),
    .A(_1257_),
    .B(_1263_));
 sg13g2_nor2_1 _4398_ (.A(_1254_),
    .B(_1265_),
    .Y(_0276_));
 sg13g2_nand2_1 _4399_ (.Y(_1266_),
    .A(\mem[31][0] ),
    .B(\mem[15][3] ));
 sg13g2_nand2_1 _4400_ (.Y(_1267_),
    .A(\mem[31][1] ),
    .B(\mem[15][2] ));
 sg13g2_nand2_1 _4401_ (.Y(_1268_),
    .A(net498),
    .B(\mem[31][3] ));
 sg13g2_and4_1 _4402_ (.A(net499),
    .B(net498),
    .C(\mem[31][2] ),
    .D(\mem[31][3] ),
    .X(_1269_));
 sg13g2_a22oi_1 _4403_ (.Y(_1270_),
    .B1(\mem[31][3] ),
    .B2(net499),
    .A2(\mem[31][2] ),
    .A1(net498));
 sg13g2_nor3_1 _4404_ (.A(_1267_),
    .B(_1269_),
    .C(_1270_),
    .Y(_1271_));
 sg13g2_o21ai_1 _4405_ (.B1(_1267_),
    .Y(_1272_),
    .A1(_1269_),
    .A2(_1270_));
 sg13g2_nor2b_1 _4406_ (.A(_1271_),
    .B_N(_1272_),
    .Y(_1273_));
 sg13g2_nand2_1 _4407_ (.Y(_1274_),
    .A(_1259_),
    .B(_1273_));
 sg13g2_xor2_1 _4408_ (.B(_1273_),
    .A(_1259_),
    .X(_1275_));
 sg13g2_nand2b_1 _4409_ (.Y(_1276_),
    .B(_1275_),
    .A_N(_1266_));
 sg13g2_xnor2_1 _4410_ (.Y(_1277_),
    .A(_1266_),
    .B(_1275_));
 sg13g2_nand2_1 _4411_ (.Y(_1278_),
    .A(_1262_),
    .B(_1277_));
 sg13g2_xnor2_1 _4412_ (.Y(_1279_),
    .A(_1262_),
    .B(_1277_));
 sg13g2_xnor2_1 _4413_ (.Y(_1280_),
    .A(_1264_),
    .B(_1279_));
 sg13g2_nor2_1 _4414_ (.A(_1254_),
    .B(_1280_),
    .Y(_0277_));
 sg13g2_o21ai_1 _4415_ (.B1(_1278_),
    .Y(_1281_),
    .A1(_1264_),
    .A2(_1279_));
 sg13g2_or2_1 _4416_ (.X(_1282_),
    .B(_1271_),
    .A(_1269_));
 sg13g2_nand2_1 _4417_ (.Y(_1283_),
    .A(\mem[31][1] ),
    .B(\mem[15][3] ));
 sg13g2_nand2_1 _4418_ (.Y(_1284_),
    .A(\mem[15][2] ),
    .B(\mem[31][3] ));
 sg13g2_nand2_2 _4419_ (.Y(_1285_),
    .A(net779),
    .B(\mem[31][2] ));
 sg13g2_xor2_1 _4420_ (.B(_1285_),
    .A(_1268_),
    .X(_1286_));
 sg13g2_nand2b_1 _4421_ (.Y(_1287_),
    .B(_1286_),
    .A_N(_1283_));
 sg13g2_xnor2_1 _4422_ (.Y(_1288_),
    .A(_1283_),
    .B(_1286_));
 sg13g2_nand2_1 _4423_ (.Y(_1289_),
    .A(_1282_),
    .B(_1288_));
 sg13g2_xnor2_1 _4424_ (.Y(_1290_),
    .A(_1282_),
    .B(_1288_));
 sg13g2_a21o_1 _4425_ (.A2(_1276_),
    .A1(_1274_),
    .B1(_1290_),
    .X(_1291_));
 sg13g2_inv_1 _4426_ (.Y(_1292_),
    .A(_1291_));
 sg13g2_nand3_1 _4427_ (.B(_1276_),
    .C(_1290_),
    .A(_1274_),
    .Y(_1293_));
 sg13g2_nand2_1 _4428_ (.Y(_1294_),
    .A(_1291_),
    .B(_1293_));
 sg13g2_xor2_1 _4429_ (.B(_1294_),
    .A(_1281_),
    .X(_1295_));
 sg13g2_nor2_1 _4430_ (.A(_1254_),
    .B(_1295_),
    .Y(_0278_));
 sg13g2_nor2_1 _4431_ (.A(_1281_),
    .B(_1292_),
    .Y(_1296_));
 sg13g2_a21oi_1 _4432_ (.A1(_1281_),
    .A2(_1293_),
    .Y(_1297_),
    .B1(_1292_));
 sg13g2_o21ai_1 _4433_ (.B1(_1287_),
    .Y(_1298_),
    .A1(_1268_),
    .A2(_1285_));
 sg13g2_nand2_1 _4434_ (.Y(_1299_),
    .A(\mem[31][2] ),
    .B(\mem[15][3] ));
 sg13g2_nand2_1 _4435_ (.Y(_1300_),
    .A(net739),
    .B(net777));
 sg13g2_xor2_1 _4436_ (.B(_1299_),
    .A(_1284_),
    .X(_1301_));
 sg13g2_nand2_1 _4437_ (.Y(_1302_),
    .A(_1298_),
    .B(_1301_));
 sg13g2_xnor2_1 _4438_ (.Y(_1303_),
    .A(_1298_),
    .B(_1301_));
 sg13g2_xnor2_1 _4439_ (.Y(_1304_),
    .A(_1289_),
    .B(_1303_));
 sg13g2_xnor2_1 _4440_ (.Y(_1305_),
    .A(_1297_),
    .B(_1304_));
 sg13g2_nor2_1 _4441_ (.A(_1254_),
    .B(_1305_),
    .Y(_0279_));
 sg13g2_nand2b_1 _4442_ (.Y(_1306_),
    .B(_1285_),
    .A_N(_1300_));
 sg13g2_xor2_1 _4443_ (.B(_1306_),
    .A(_1302_),
    .X(_1307_));
 sg13g2_a21oi_1 _4444_ (.A1(_1289_),
    .A2(_1296_),
    .Y(_1308_),
    .B1(_1303_));
 sg13g2_xnor2_1 _4445_ (.Y(_1309_),
    .A(_1307_),
    .B(_1308_));
 sg13g2_nor2_1 _4446_ (.A(_1254_),
    .B(_1309_),
    .Y(_0280_));
 sg13g2_a21oi_1 _4447_ (.A1(_1285_),
    .A2(_1302_),
    .Y(_1310_),
    .B1(_1300_));
 sg13g2_a21oi_1 _4448_ (.A1(_1307_),
    .A2(_1308_),
    .Y(_1311_),
    .B1(_1310_));
 sg13g2_nor2_1 _4449_ (.A(_1254_),
    .B(_1311_),
    .Y(_0281_));
 sg13g2_and3_1 _4450_ (.X(_0282_),
    .A(net497),
    .B(net735),
    .C(_1253_));
 sg13g2_a22oi_1 _4451_ (.Y(_1312_),
    .B1(\mem[30][1] ),
    .B2(net424),
    .A2(\mem[14][1] ),
    .A1(\mem[30][0] ));
 sg13g2_and4_1 _4452_ (.A(net497),
    .B(\mem[30][0] ),
    .C(net496),
    .D(\mem[30][1] ),
    .X(_1313_));
 sg13g2_nor3_1 _4453_ (.A(_1252_),
    .B(net425),
    .C(_1313_),
    .Y(_0283_));
 sg13g2_a22oi_1 _4454_ (.Y(_1314_),
    .B1(\mem[30][2] ),
    .B2(net497),
    .A2(\mem[30][1] ),
    .A1(net496));
 sg13g2_nand4_1 _4455_ (.B(net496),
    .C(\mem[30][1] ),
    .A(net497),
    .Y(_1315_),
    .D(\mem[30][2] ));
 sg13g2_nor2b_1 _4456_ (.A(_1314_),
    .B_N(_1315_),
    .Y(_1316_));
 sg13g2_and3_1 _4457_ (.X(_1317_),
    .A(\mem[30][0] ),
    .B(\mem[14][2] ),
    .C(_1316_));
 sg13g2_a21oi_1 _4458_ (.A1(\mem[30][0] ),
    .A2(\mem[14][2] ),
    .Y(_1318_),
    .B1(_1316_));
 sg13g2_nor2_1 _4459_ (.A(_1317_),
    .B(_1318_),
    .Y(_1319_));
 sg13g2_and2_1 _4460_ (.A(_1313_),
    .B(_1319_),
    .X(_1320_));
 sg13g2_nor2_1 _4461_ (.A(_1313_),
    .B(_1319_),
    .Y(_1321_));
 sg13g2_nor3_1 _4462_ (.A(_1252_),
    .B(_1320_),
    .C(_1321_),
    .Y(_0284_));
 sg13g2_nand2_1 _4463_ (.Y(_1322_),
    .A(\mem[30][0] ),
    .B(\mem[14][3] ));
 sg13g2_nand2_1 _4464_ (.Y(_1323_),
    .A(\mem[30][1] ),
    .B(\mem[14][2] ));
 sg13g2_nand2_1 _4465_ (.Y(_1324_),
    .A(net496),
    .B(\mem[30][3] ));
 sg13g2_and4_1 _4466_ (.A(net497),
    .B(net496),
    .C(\mem[30][2] ),
    .D(\mem[30][3] ),
    .X(_1325_));
 sg13g2_a22oi_1 _4467_ (.Y(_1326_),
    .B1(\mem[30][3] ),
    .B2(net497),
    .A2(\mem[30][2] ),
    .A1(net496));
 sg13g2_nor3_1 _4468_ (.A(_1323_),
    .B(_1325_),
    .C(_1326_),
    .Y(_1327_));
 sg13g2_o21ai_1 _4469_ (.B1(_1323_),
    .Y(_1328_),
    .A1(_1325_),
    .A2(_1326_));
 sg13g2_nor2b_1 _4470_ (.A(_1327_),
    .B_N(_1328_),
    .Y(_1329_));
 sg13g2_inv_1 _4471_ (.Y(_1330_),
    .A(_1329_));
 sg13g2_xnor2_1 _4472_ (.Y(_1331_),
    .A(_1315_),
    .B(_1329_));
 sg13g2_nand2b_1 _4473_ (.Y(_1332_),
    .B(_1331_),
    .A_N(_1322_));
 sg13g2_xnor2_1 _4474_ (.Y(_1333_),
    .A(_1322_),
    .B(_1331_));
 sg13g2_and2_1 _4475_ (.A(_1317_),
    .B(_1333_),
    .X(_1334_));
 sg13g2_xor2_1 _4476_ (.B(_1333_),
    .A(_1317_),
    .X(_1335_));
 sg13g2_o21ai_1 _4477_ (.B1(_1253_),
    .Y(_1336_),
    .A1(_1320_),
    .A2(_1335_));
 sg13g2_a21oi_1 _4478_ (.A1(_1320_),
    .A2(_1335_),
    .Y(_0285_),
    .B1(_1336_));
 sg13g2_or2_1 _4479_ (.X(_1337_),
    .B(_1327_),
    .A(_1325_));
 sg13g2_nand2_1 _4480_ (.Y(_1338_),
    .A(\mem[30][1] ),
    .B(\mem[14][3] ));
 sg13g2_nand2_1 _4481_ (.Y(_1339_),
    .A(\mem[14][2] ),
    .B(\mem[30][3] ));
 sg13g2_nand2_2 _4482_ (.Y(_1340_),
    .A(\mem[14][2] ),
    .B(\mem[30][2] ));
 sg13g2_xor2_1 _4483_ (.B(_1340_),
    .A(_1324_),
    .X(_1341_));
 sg13g2_nand2b_1 _4484_ (.Y(_1342_),
    .B(_1341_),
    .A_N(_1338_));
 sg13g2_xnor2_1 _4485_ (.Y(_1343_),
    .A(_1338_),
    .B(_1341_));
 sg13g2_nand2_1 _4486_ (.Y(_1344_),
    .A(_1337_),
    .B(_1343_));
 sg13g2_xnor2_1 _4487_ (.Y(_1345_),
    .A(_1337_),
    .B(_1343_));
 sg13g2_o21ai_1 _4488_ (.B1(_1332_),
    .Y(_1346_),
    .A1(_1315_),
    .A2(_1330_));
 sg13g2_nand2b_1 _4489_ (.Y(_1347_),
    .B(_1346_),
    .A_N(_1345_));
 sg13g2_xor2_1 _4490_ (.B(_1346_),
    .A(_1345_),
    .X(_1348_));
 sg13g2_a21o_1 _4491_ (.A2(_1335_),
    .A1(_1320_),
    .B1(_1334_),
    .X(_1349_));
 sg13g2_inv_1 _4492_ (.Y(_1350_),
    .A(_1349_));
 sg13g2_nand2b_1 _4493_ (.Y(_1351_),
    .B(_1349_),
    .A_N(_1348_));
 sg13g2_a21oi_1 _4494_ (.A1(_1348_),
    .A2(_1350_),
    .Y(_1352_),
    .B1(_1252_));
 sg13g2_and2_1 _4495_ (.A(_1351_),
    .B(_1352_),
    .X(_0286_));
 sg13g2_nand2_1 _4496_ (.Y(_1353_),
    .A(_1347_),
    .B(_1351_));
 sg13g2_o21ai_1 _4497_ (.B1(_1342_),
    .Y(_1354_),
    .A1(_1324_),
    .A2(_1340_));
 sg13g2_nand2_1 _4498_ (.Y(_1355_),
    .A(\mem[30][2] ),
    .B(\mem[14][3] ));
 sg13g2_nand2_1 _4499_ (.Y(_1356_),
    .A(net774),
    .B(net852));
 sg13g2_xor2_1 _4500_ (.B(_1355_),
    .A(_1339_),
    .X(_1357_));
 sg13g2_nand2_1 _4501_ (.Y(_1358_),
    .A(_1354_),
    .B(_1357_));
 sg13g2_xnor2_1 _4502_ (.Y(_1359_),
    .A(_1354_),
    .B(_1357_));
 sg13g2_xor2_1 _4503_ (.B(_1359_),
    .A(_1344_),
    .X(_1360_));
 sg13g2_xnor2_1 _4504_ (.Y(_1361_),
    .A(_1353_),
    .B(_1360_));
 sg13g2_nor2_1 _4505_ (.A(_1252_),
    .B(_1361_),
    .Y(_0287_));
 sg13g2_and2_1 _4506_ (.A(_1344_),
    .B(_1347_),
    .X(_1362_));
 sg13g2_a21oi_1 _4507_ (.A1(_1350_),
    .A2(_1362_),
    .Y(_1363_),
    .B1(_1359_));
 sg13g2_nand2b_1 _4508_ (.Y(_1364_),
    .B(_1340_),
    .A_N(_1356_));
 sg13g2_xor2_1 _4509_ (.B(_1364_),
    .A(_1358_),
    .X(_1365_));
 sg13g2_xnor2_1 _4510_ (.Y(_1366_),
    .A(_1363_),
    .B(_1365_));
 sg13g2_nor2_1 _4511_ (.A(_1252_),
    .B(_1366_),
    .Y(_0288_));
 sg13g2_a21oi_1 _4512_ (.A1(_1340_),
    .A2(_1358_),
    .Y(_1367_),
    .B1(_1356_));
 sg13g2_a21oi_1 _4513_ (.A1(_1363_),
    .A2(_1365_),
    .Y(_1368_),
    .B1(_1367_));
 sg13g2_nor2_1 _4514_ (.A(_1252_),
    .B(_1368_),
    .Y(_0289_));
 sg13g2_a21oi_2 _4515_ (.B1(net483),
    .Y(_1369_),
    .A2(_1247_),
    .A1(net493));
 sg13g2_a21o_2 _4516_ (.A2(_1247_),
    .A1(net493),
    .B1(_1190_),
    .X(_1370_));
 sg13g2_o21ai_1 _4517_ (.B1(_1370_),
    .Y(_1371_),
    .A1(_1188_),
    .A2(_1189_));
 sg13g2_inv_1 _4518_ (.Y(_1372_),
    .A(_1371_));
 sg13g2_and3_1 _4519_ (.X(_0290_),
    .A(\mem[13][0] ),
    .B(net716),
    .C(_1372_));
 sg13g2_nand4_1 _4520_ (.B(net860),
    .C(\mem[13][1] ),
    .A(\mem[13][0] ),
    .Y(_1373_),
    .D(\mem[29][1] ));
 sg13g2_inv_1 _4521_ (.Y(_1374_),
    .A(_1373_));
 sg13g2_a22oi_1 _4522_ (.Y(_1375_),
    .B1(\mem[29][1] ),
    .B2(net794),
    .A2(\mem[13][1] ),
    .A1(net716));
 sg13g2_nor3_1 _4523_ (.A(_1371_),
    .B(_1374_),
    .C(net795),
    .Y(_0291_));
 sg13g2_a22oi_1 _4524_ (.Y(_1376_),
    .B1(\mem[29][2] ),
    .B2(\mem[13][0] ),
    .A2(\mem[29][1] ),
    .A1(\mem[13][1] ));
 sg13g2_nand2_1 _4525_ (.Y(_1377_),
    .A(\mem[13][1] ),
    .B(\mem[29][2] ));
 sg13g2_and4_2 _4526_ (.A(\mem[13][0] ),
    .B(\mem[13][1] ),
    .C(\mem[29][1] ),
    .D(\mem[29][2] ),
    .X(_1378_));
 sg13g2_nor2_1 _4527_ (.A(_1376_),
    .B(_1378_),
    .Y(_1379_));
 sg13g2_nand2_1 _4528_ (.Y(_1380_),
    .A(\mem[29][0] ),
    .B(\mem[13][2] ));
 sg13g2_nor3_1 _4529_ (.A(_1376_),
    .B(_1378_),
    .C(_1380_),
    .Y(_1381_));
 sg13g2_xor2_1 _4530_ (.B(_1380_),
    .A(_1379_),
    .X(_1382_));
 sg13g2_and2_1 _4531_ (.A(_1373_),
    .B(_1382_),
    .X(_1383_));
 sg13g2_nor2_2 _4532_ (.A(_1373_),
    .B(_1382_),
    .Y(_1384_));
 sg13g2_nor3_1 _4533_ (.A(_1371_),
    .B(_1383_),
    .C(_1384_),
    .Y(_0292_));
 sg13g2_nand2_1 _4534_ (.Y(_1385_),
    .A(\mem[29][0] ),
    .B(\mem[13][3] ));
 sg13g2_nand2_1 _4535_ (.Y(_1386_),
    .A(\mem[29][1] ),
    .B(\mem[13][2] ));
 sg13g2_nand2_1 _4536_ (.Y(_1387_),
    .A(\mem[13][1] ),
    .B(\mem[29][3] ));
 sg13g2_nand2_1 _4537_ (.Y(_1388_),
    .A(\mem[13][0] ),
    .B(\mem[29][3] ));
 sg13g2_xor2_1 _4538_ (.B(_1388_),
    .A(_1377_),
    .X(_1389_));
 sg13g2_nand2b_1 _4539_ (.Y(_1390_),
    .B(_1389_),
    .A_N(_1386_));
 sg13g2_xnor2_1 _4540_ (.Y(_1391_),
    .A(_1386_),
    .B(_1389_));
 sg13g2_nand2_1 _4541_ (.Y(_1392_),
    .A(_1378_),
    .B(_1391_));
 sg13g2_xor2_1 _4542_ (.B(_1391_),
    .A(_1378_),
    .X(_1393_));
 sg13g2_nand2b_1 _4543_ (.Y(_1394_),
    .B(_1393_),
    .A_N(_1385_));
 sg13g2_xnor2_1 _4544_ (.Y(_1395_),
    .A(_1385_),
    .B(_1393_));
 sg13g2_and2_1 _4545_ (.A(_1381_),
    .B(_1395_),
    .X(_1396_));
 sg13g2_xor2_1 _4546_ (.B(_1395_),
    .A(_1381_),
    .X(_1397_));
 sg13g2_o21ai_1 _4547_ (.B1(_1372_),
    .Y(_1398_),
    .A1(_1384_),
    .A2(_1397_));
 sg13g2_a21oi_1 _4548_ (.A1(_1384_),
    .A2(_1397_),
    .Y(_0293_),
    .B1(_1398_));
 sg13g2_a21oi_1 _4549_ (.A1(_1384_),
    .A2(_1397_),
    .Y(_1399_),
    .B1(_1396_));
 sg13g2_o21ai_1 _4550_ (.B1(_1390_),
    .Y(_1400_),
    .A1(_1377_),
    .A2(_1388_));
 sg13g2_nand2_1 _4551_ (.Y(_1401_),
    .A(\mem[29][1] ),
    .B(\mem[13][3] ));
 sg13g2_nand2_1 _4552_ (.Y(_1402_),
    .A(\mem[13][2] ),
    .B(\mem[29][3] ));
 sg13g2_nand2_2 _4553_ (.Y(_1403_),
    .A(\mem[13][2] ),
    .B(\mem[29][2] ));
 sg13g2_or2_1 _4554_ (.X(_1404_),
    .B(_1403_),
    .A(_1387_));
 sg13g2_xnor2_1 _4555_ (.Y(_1405_),
    .A(_1387_),
    .B(_1403_));
 sg13g2_xor2_1 _4556_ (.B(_1405_),
    .A(_1401_),
    .X(_1406_));
 sg13g2_nand2_1 _4557_ (.Y(_1407_),
    .A(_1400_),
    .B(_1406_));
 sg13g2_xnor2_1 _4558_ (.Y(_1408_),
    .A(_1400_),
    .B(_1406_));
 sg13g2_a21o_1 _4559_ (.A2(_1394_),
    .A1(_1392_),
    .B1(_1408_),
    .X(_1409_));
 sg13g2_nand3_1 _4560_ (.B(_1394_),
    .C(_1408_),
    .A(_1392_),
    .Y(_1410_));
 sg13g2_nand2_1 _4561_ (.Y(_1411_),
    .A(_1409_),
    .B(_1410_));
 sg13g2_or2_1 _4562_ (.X(_1412_),
    .B(_1411_),
    .A(_1399_));
 sg13g2_nand2_1 _4563_ (.Y(_1413_),
    .A(_1372_),
    .B(_1412_));
 sg13g2_a21oi_1 _4564_ (.A1(_1399_),
    .A2(_1411_),
    .Y(_0294_),
    .B1(_1413_));
 sg13g2_nand2_1 _4565_ (.Y(_1414_),
    .A(_1409_),
    .B(_1412_));
 sg13g2_o21ai_1 _4566_ (.B1(_1404_),
    .Y(_1415_),
    .A1(_1401_),
    .A2(_1405_));
 sg13g2_nand2_1 _4567_ (.Y(_1416_),
    .A(\mem[29][2] ),
    .B(\mem[13][3] ));
 sg13g2_nand2_1 _4568_ (.Y(_1417_),
    .A(net829),
    .B(net810));
 sg13g2_xor2_1 _4569_ (.B(_1416_),
    .A(_1402_),
    .X(_1418_));
 sg13g2_nand2_1 _4570_ (.Y(_1419_),
    .A(_1415_),
    .B(_1418_));
 sg13g2_xnor2_1 _4571_ (.Y(_1420_),
    .A(_1415_),
    .B(_1418_));
 sg13g2_xor2_1 _4572_ (.B(_1420_),
    .A(_1407_),
    .X(_1421_));
 sg13g2_xnor2_1 _4573_ (.Y(_1422_),
    .A(_1414_),
    .B(_1421_));
 sg13g2_nor2_1 _4574_ (.A(_1371_),
    .B(_1422_),
    .Y(_0295_));
 sg13g2_nand2b_1 _4575_ (.Y(_1423_),
    .B(_1403_),
    .A_N(_1417_));
 sg13g2_xor2_1 _4576_ (.B(_1423_),
    .A(_1419_),
    .X(_1424_));
 sg13g2_and2_1 _4577_ (.A(_1407_),
    .B(_1409_),
    .X(_1425_));
 sg13g2_a21oi_1 _4578_ (.A1(_1399_),
    .A2(_1425_),
    .Y(_1426_),
    .B1(_1420_));
 sg13g2_or2_1 _4579_ (.X(_1427_),
    .B(_1426_),
    .A(_1424_));
 sg13g2_nand2_1 _4580_ (.Y(_1428_),
    .A(_1424_),
    .B(_1426_));
 sg13g2_and3_1 _4581_ (.X(_0296_),
    .A(_1372_),
    .B(_1427_),
    .C(_1428_));
 sg13g2_a21o_1 _4582_ (.A2(_1419_),
    .A1(_1403_),
    .B1(_1417_),
    .X(_1429_));
 sg13g2_a21oi_1 _4583_ (.A1(_1428_),
    .A2(_1429_),
    .Y(_0297_),
    .B1(_1371_));
 sg13g2_and3_1 _4584_ (.X(_0298_),
    .A(net674),
    .B(\mem[28][0] ),
    .C(_1370_));
 sg13g2_a22oi_1 _4585_ (.Y(_1430_),
    .B1(\mem[28][1] ),
    .B2(net674),
    .A2(\mem[12][1] ),
    .A1(net699));
 sg13g2_nand4_1 _4586_ (.B(net699),
    .C(net853),
    .A(net674),
    .Y(_1431_),
    .D(\mem[28][1] ));
 sg13g2_inv_1 _4587_ (.Y(_1432_),
    .A(_1431_));
 sg13g2_nor3_1 _4588_ (.A(_1369_),
    .B(net700),
    .C(_1432_),
    .Y(_0299_));
 sg13g2_a22oi_1 _4589_ (.Y(_1433_),
    .B1(\mem[28][2] ),
    .B2(\mem[12][0] ),
    .A2(\mem[28][1] ),
    .A1(\mem[12][1] ));
 sg13g2_nand4_1 _4590_ (.B(\mem[12][1] ),
    .C(\mem[28][1] ),
    .A(\mem[12][0] ),
    .Y(_1434_),
    .D(\mem[28][2] ));
 sg13g2_nor2b_1 _4591_ (.A(_1433_),
    .B_N(_1434_),
    .Y(_1435_));
 sg13g2_and3_1 _4592_ (.X(_1436_),
    .A(\mem[28][0] ),
    .B(\mem[12][2] ),
    .C(_1435_));
 sg13g2_inv_1 _4593_ (.Y(_1437_),
    .A(_1436_));
 sg13g2_a21oi_1 _4594_ (.A1(\mem[28][0] ),
    .A2(\mem[12][2] ),
    .Y(_1438_),
    .B1(_1435_));
 sg13g2_or2_1 _4595_ (.X(_1439_),
    .B(_1438_),
    .A(_1436_));
 sg13g2_and2_1 _4596_ (.A(_1431_),
    .B(_1439_),
    .X(_1440_));
 sg13g2_nor2_1 _4597_ (.A(_1431_),
    .B(_1439_),
    .Y(_1441_));
 sg13g2_nor3_1 _4598_ (.A(_1369_),
    .B(_1440_),
    .C(_1441_),
    .Y(_0300_));
 sg13g2_and2_1 _4599_ (.A(\mem[28][0] ),
    .B(\mem[12][3] ),
    .X(_1442_));
 sg13g2_nand2_1 _4600_ (.Y(_1443_),
    .A(\mem[28][1] ),
    .B(\mem[12][2] ));
 sg13g2_nand2_1 _4601_ (.Y(_1444_),
    .A(\mem[12][1] ),
    .B(\mem[28][3] ));
 sg13g2_nor3_1 _4602_ (.A(_2097_),
    .B(_2104_),
    .C(_1444_),
    .Y(_1445_));
 sg13g2_a22oi_1 _4603_ (.Y(_1446_),
    .B1(\mem[28][3] ),
    .B2(\mem[12][0] ),
    .A2(\mem[28][2] ),
    .A1(\mem[12][1] ));
 sg13g2_nor3_1 _4604_ (.A(_1443_),
    .B(_1445_),
    .C(_1446_),
    .Y(_1447_));
 sg13g2_o21ai_1 _4605_ (.B1(_1443_),
    .Y(_1448_),
    .A1(_1445_),
    .A2(_1446_));
 sg13g2_nor2b_1 _4606_ (.A(_1447_),
    .B_N(_1448_),
    .Y(_1449_));
 sg13g2_nor2b_1 _4607_ (.A(_1434_),
    .B_N(_1449_),
    .Y(_1450_));
 sg13g2_xnor2_1 _4608_ (.Y(_1451_),
    .A(_1434_),
    .B(_1449_));
 sg13g2_xnor2_1 _4609_ (.Y(_1452_),
    .A(_1442_),
    .B(_1451_));
 sg13g2_nor2_1 _4610_ (.A(_1437_),
    .B(_1452_),
    .Y(_1453_));
 sg13g2_xnor2_1 _4611_ (.Y(_1454_),
    .A(_1436_),
    .B(_1452_));
 sg13g2_xnor2_1 _4612_ (.Y(_1455_),
    .A(_1441_),
    .B(_1454_));
 sg13g2_nor2_1 _4613_ (.A(_1369_),
    .B(_1455_),
    .Y(_0301_));
 sg13g2_a21o_1 _4614_ (.A2(_1454_),
    .A1(_1441_),
    .B1(_1453_),
    .X(_1456_));
 sg13g2_or2_1 _4615_ (.X(_1457_),
    .B(_1447_),
    .A(_1445_));
 sg13g2_nand2_1 _4616_ (.Y(_1458_),
    .A(\mem[28][1] ),
    .B(\mem[12][3] ));
 sg13g2_nand2_1 _4617_ (.Y(_1459_),
    .A(\mem[12][2] ),
    .B(\mem[28][3] ));
 sg13g2_nand2_2 _4618_ (.Y(_1460_),
    .A(net861),
    .B(net831));
 sg13g2_xor2_1 _4619_ (.B(_1460_),
    .A(_1444_),
    .X(_1461_));
 sg13g2_nand2b_1 _4620_ (.Y(_1462_),
    .B(_1461_),
    .A_N(_1458_));
 sg13g2_xnor2_1 _4621_ (.Y(_1463_),
    .A(_1458_),
    .B(_1461_));
 sg13g2_nand2_1 _4622_ (.Y(_1464_),
    .A(_1457_),
    .B(_1463_));
 sg13g2_xor2_1 _4623_ (.B(_1463_),
    .A(_1457_),
    .X(_1465_));
 sg13g2_a21oi_1 _4624_ (.A1(_1442_),
    .A2(_1451_),
    .Y(_1466_),
    .B1(_1450_));
 sg13g2_nand2b_1 _4625_ (.Y(_1467_),
    .B(_1465_),
    .A_N(_1466_));
 sg13g2_xnor2_1 _4626_ (.Y(_1468_),
    .A(_1465_),
    .B(_1466_));
 sg13g2_or2_1 _4627_ (.X(_1469_),
    .B(_1468_),
    .A(_1456_));
 sg13g2_nand2_1 _4628_ (.Y(_1470_),
    .A(_1456_),
    .B(_1468_));
 sg13g2_and3_1 _4629_ (.X(_0302_),
    .A(_1370_),
    .B(_1469_),
    .C(_1470_));
 sg13g2_nor2b_1 _4630_ (.A(_1456_),
    .B_N(_1467_),
    .Y(_1471_));
 sg13g2_o21ai_1 _4631_ (.B1(_1462_),
    .Y(_1472_),
    .A1(_1444_),
    .A2(_1460_));
 sg13g2_nand2_1 _4632_ (.Y(_1473_),
    .A(\mem[28][2] ),
    .B(\mem[12][3] ));
 sg13g2_nand2_1 _4633_ (.Y(_1474_),
    .A(net785),
    .B(net729));
 sg13g2_xor2_1 _4634_ (.B(_1473_),
    .A(_1459_),
    .X(_1475_));
 sg13g2_nand2_1 _4635_ (.Y(_1476_),
    .A(_1472_),
    .B(_1475_));
 sg13g2_xnor2_1 _4636_ (.Y(_1477_),
    .A(_1472_),
    .B(_1475_));
 sg13g2_xnor2_1 _4637_ (.Y(_1478_),
    .A(_1464_),
    .B(_1477_));
 sg13g2_and3_1 _4638_ (.X(_1479_),
    .A(_1467_),
    .B(_1470_),
    .C(_1478_));
 sg13g2_a21oi_1 _4639_ (.A1(_1467_),
    .A2(_1470_),
    .Y(_1480_),
    .B1(_1478_));
 sg13g2_nor3_2 _4640_ (.A(_1369_),
    .B(_1479_),
    .C(_1480_),
    .Y(_0303_));
 sg13g2_a21oi_1 _4641_ (.A1(_1464_),
    .A2(_1471_),
    .Y(_1481_),
    .B1(_1477_));
 sg13g2_nand2b_1 _4642_ (.Y(_1482_),
    .B(_1460_),
    .A_N(_1474_));
 sg13g2_xor2_1 _4643_ (.B(_1482_),
    .A(_1476_),
    .X(_1483_));
 sg13g2_xnor2_1 _4644_ (.Y(_1484_),
    .A(_1481_),
    .B(_1483_));
 sg13g2_nor2_1 _4645_ (.A(_1369_),
    .B(_1484_),
    .Y(_0304_));
 sg13g2_a21oi_1 _4646_ (.A1(_1460_),
    .A2(_1476_),
    .Y(_1485_),
    .B1(_1474_));
 sg13g2_a21oi_1 _4647_ (.A1(_1481_),
    .A2(_1483_),
    .Y(_1486_),
    .B1(_1485_));
 sg13g2_nor2_1 _4648_ (.A(_1369_),
    .B(_1486_),
    .Y(_0305_));
 sg13g2_a21oi_2 _4649_ (.B1(_1370_),
    .Y(_1487_),
    .A2(_1250_),
    .A1(net492));
 sg13g2_o21ai_1 _4650_ (.B1(_1369_),
    .Y(_1488_),
    .A1(_1248_),
    .A2(_1249_));
 sg13g2_and3_1 _4651_ (.X(_0306_),
    .A(\mem[11][0] ),
    .B(net737),
    .C(_1488_));
 sg13g2_a22oi_1 _4652_ (.Y(_1489_),
    .B1(\mem[27][1] ),
    .B2(net769),
    .A2(\mem[11][1] ),
    .A1(net737));
 sg13g2_nand4_1 _4653_ (.B(net737),
    .C(net798),
    .A(net769),
    .Y(_1490_),
    .D(net799));
 sg13g2_nand2_1 _4654_ (.Y(_1491_),
    .A(_1488_),
    .B(_1490_));
 sg13g2_nor2_1 _4655_ (.A(net770),
    .B(_1491_),
    .Y(_0307_));
 sg13g2_a22oi_1 _4656_ (.Y(_1492_),
    .B1(\mem[27][2] ),
    .B2(\mem[11][0] ),
    .A2(\mem[27][1] ),
    .A1(\mem[11][1] ));
 sg13g2_nand2_1 _4657_ (.Y(_1493_),
    .A(\mem[11][1] ),
    .B(\mem[27][2] ));
 sg13g2_and4_2 _4658_ (.A(\mem[11][0] ),
    .B(\mem[11][1] ),
    .C(\mem[27][1] ),
    .D(\mem[27][2] ),
    .X(_1494_));
 sg13g2_nor2_1 _4659_ (.A(_1492_),
    .B(_1494_),
    .Y(_1495_));
 sg13g2_nand2_1 _4660_ (.Y(_1496_),
    .A(\mem[27][0] ),
    .B(\mem[11][2] ));
 sg13g2_nor3_1 _4661_ (.A(_1492_),
    .B(_1494_),
    .C(_1496_),
    .Y(_1497_));
 sg13g2_xor2_1 _4662_ (.B(_1496_),
    .A(_1495_),
    .X(_1498_));
 sg13g2_or2_1 _4663_ (.X(_1499_),
    .B(_1498_),
    .A(_1490_));
 sg13g2_nand2_1 _4664_ (.Y(_1500_),
    .A(_1488_),
    .B(_1499_));
 sg13g2_a21oi_1 _4665_ (.A1(_1490_),
    .A2(_1498_),
    .Y(_0308_),
    .B1(_1500_));
 sg13g2_nand2_1 _4666_ (.Y(_1501_),
    .A(\mem[27][0] ),
    .B(\mem[11][3] ));
 sg13g2_nand2_1 _4667_ (.Y(_1502_),
    .A(\mem[27][1] ),
    .B(\mem[11][2] ));
 sg13g2_nand2_1 _4668_ (.Y(_1503_),
    .A(\mem[11][1] ),
    .B(\mem[27][3] ));
 sg13g2_nand2_1 _4669_ (.Y(_1504_),
    .A(\mem[11][0] ),
    .B(\mem[27][3] ));
 sg13g2_xor2_1 _4670_ (.B(_1504_),
    .A(_1493_),
    .X(_1505_));
 sg13g2_nand2b_1 _4671_ (.Y(_1506_),
    .B(_1505_),
    .A_N(_1502_));
 sg13g2_xnor2_1 _4672_ (.Y(_1507_),
    .A(_1502_),
    .B(_1505_));
 sg13g2_nand2_1 _4673_ (.Y(_1508_),
    .A(_1494_),
    .B(_1507_));
 sg13g2_xor2_1 _4674_ (.B(_1507_),
    .A(_1494_),
    .X(_1509_));
 sg13g2_nand2b_1 _4675_ (.Y(_1510_),
    .B(_1509_),
    .A_N(_1501_));
 sg13g2_xnor2_1 _4676_ (.Y(_1511_),
    .A(_1501_),
    .B(_1509_));
 sg13g2_xnor2_1 _4677_ (.Y(_1512_),
    .A(_1497_),
    .B(_1511_));
 sg13g2_nor2_1 _4678_ (.A(_1499_),
    .B(_1512_),
    .Y(_1513_));
 sg13g2_a21oi_1 _4679_ (.A1(_1499_),
    .A2(_1512_),
    .Y(_1514_),
    .B1(_1487_));
 sg13g2_nor2b_1 _4680_ (.A(_1513_),
    .B_N(_1514_),
    .Y(_0309_));
 sg13g2_a21oi_1 _4681_ (.A1(_1497_),
    .A2(_1511_),
    .Y(_1515_),
    .B1(_1513_));
 sg13g2_o21ai_1 _4682_ (.B1(_1506_),
    .Y(_1516_),
    .A1(_1493_),
    .A2(_1504_));
 sg13g2_nand2_1 _4683_ (.Y(_1517_),
    .A(\mem[27][1] ),
    .B(\mem[11][3] ));
 sg13g2_nand2_1 _4684_ (.Y(_1518_),
    .A(\mem[11][2] ),
    .B(\mem[27][3] ));
 sg13g2_nand2_2 _4685_ (.Y(_1519_),
    .A(\mem[11][2] ),
    .B(\mem[27][2] ));
 sg13g2_or2_1 _4686_ (.X(_1520_),
    .B(_1519_),
    .A(_1503_));
 sg13g2_xnor2_1 _4687_ (.Y(_1521_),
    .A(_1503_),
    .B(_1519_));
 sg13g2_xor2_1 _4688_ (.B(_1521_),
    .A(_1517_),
    .X(_1522_));
 sg13g2_nand2_1 _4689_ (.Y(_1523_),
    .A(_1516_),
    .B(_1522_));
 sg13g2_xnor2_1 _4690_ (.Y(_1524_),
    .A(_1516_),
    .B(_1522_));
 sg13g2_a21o_1 _4691_ (.A2(_1510_),
    .A1(_1508_),
    .B1(_1524_),
    .X(_1525_));
 sg13g2_nand3_1 _4692_ (.B(_1510_),
    .C(_1524_),
    .A(_1508_),
    .Y(_1526_));
 sg13g2_nand2_1 _4693_ (.Y(_1527_),
    .A(_1525_),
    .B(_1526_));
 sg13g2_or2_1 _4694_ (.X(_1528_),
    .B(_1527_),
    .A(_1515_));
 sg13g2_nand2_1 _4695_ (.Y(_1529_),
    .A(_1488_),
    .B(_1528_));
 sg13g2_a21oi_1 _4696_ (.A1(_1515_),
    .A2(_1527_),
    .Y(_0310_),
    .B1(_1529_));
 sg13g2_nand2_1 _4697_ (.Y(_1530_),
    .A(_1525_),
    .B(_1528_));
 sg13g2_o21ai_1 _4698_ (.B1(_1520_),
    .Y(_1531_),
    .A1(_1517_),
    .A2(_1521_));
 sg13g2_nand2_1 _4699_ (.Y(_1532_),
    .A(\mem[27][2] ),
    .B(\mem[11][3] ));
 sg13g2_nand2_1 _4700_ (.Y(_1533_),
    .A(net719),
    .B(net743));
 sg13g2_xor2_1 _4701_ (.B(_1532_),
    .A(_1518_),
    .X(_1534_));
 sg13g2_nand2_1 _4702_ (.Y(_1535_),
    .A(_1531_),
    .B(_1534_));
 sg13g2_xnor2_1 _4703_ (.Y(_1536_),
    .A(_1531_),
    .B(_1534_));
 sg13g2_xor2_1 _4704_ (.B(_1536_),
    .A(_1523_),
    .X(_1537_));
 sg13g2_xnor2_1 _4705_ (.Y(_1538_),
    .A(_1530_),
    .B(_1537_));
 sg13g2_nor2_1 _4706_ (.A(_1487_),
    .B(_1538_),
    .Y(_0311_));
 sg13g2_nand2b_1 _4707_ (.Y(_1539_),
    .B(_1519_),
    .A_N(_1533_));
 sg13g2_xor2_1 _4708_ (.B(_1539_),
    .A(_1535_),
    .X(_1540_));
 sg13g2_and2_1 _4709_ (.A(_1523_),
    .B(_1525_),
    .X(_1541_));
 sg13g2_a21oi_1 _4710_ (.A1(_1515_),
    .A2(_1541_),
    .Y(_1542_),
    .B1(_1536_));
 sg13g2_or2_1 _4711_ (.X(_1543_),
    .B(_1542_),
    .A(_1540_));
 sg13g2_nand2_1 _4712_ (.Y(_1544_),
    .A(_1540_),
    .B(_1542_));
 sg13g2_and3_1 _4713_ (.X(_0312_),
    .A(_1488_),
    .B(_1543_),
    .C(_1544_));
 sg13g2_a21o_1 _4714_ (.A2(_1535_),
    .A1(_1519_),
    .B1(_1533_),
    .X(_1545_));
 sg13g2_a21oi_1 _4715_ (.A1(_1544_),
    .A2(_1545_),
    .Y(_0313_),
    .B1(_1487_));
 sg13g2_nor2_1 _4716_ (.A(\mem[0][1] ),
    .B(net493),
    .Y(_1546_));
 sg13g2_nor2_2 _4717_ (.A(net486),
    .B(_1546_),
    .Y(_1547_));
 sg13g2_a21oi_2 _4718_ (.B1(net483),
    .Y(_1548_),
    .A2(_1547_),
    .A1(net492));
 sg13g2_nand2_2 _4719_ (.Y(_1549_),
    .A(net730),
    .B(\mem[26][0] ));
 sg13g2_nor2_1 _4720_ (.A(_1548_),
    .B(net731),
    .Y(_0314_));
 sg13g2_a22oi_1 _4721_ (.Y(_1550_),
    .B1(net788),
    .B2(net730),
    .A2(\mem[10][1] ),
    .A1(\mem[26][0] ));
 sg13g2_nand2_1 _4722_ (.Y(_1551_),
    .A(\mem[10][1] ),
    .B(\mem[26][1] ));
 sg13g2_or2_1 _4723_ (.X(_1552_),
    .B(_1551_),
    .A(_1549_));
 sg13g2_inv_1 _4724_ (.Y(_1553_),
    .A(_1552_));
 sg13g2_nor3_1 _4725_ (.A(_1548_),
    .B(net789),
    .C(_1553_),
    .Y(_0315_));
 sg13g2_nand2_1 _4726_ (.Y(_1554_),
    .A(\mem[10][0] ),
    .B(\mem[26][2] ));
 sg13g2_nand2_2 _4727_ (.Y(_1555_),
    .A(\mem[26][1] ),
    .B(\mem[10][2] ));
 sg13g2_nand2_1 _4728_ (.Y(_1556_),
    .A(\mem[26][0] ),
    .B(\mem[10][2] ));
 sg13g2_or2_1 _4729_ (.X(_1557_),
    .B(_1556_),
    .A(_1551_));
 sg13g2_xnor2_1 _4730_ (.Y(_1558_),
    .A(_1551_),
    .B(_1556_));
 sg13g2_xnor2_1 _4731_ (.Y(_1559_),
    .A(_1554_),
    .B(_1558_));
 sg13g2_or2_1 _4732_ (.X(_1560_),
    .B(_1559_),
    .A(_1552_));
 sg13g2_nand2b_1 _4733_ (.Y(_1561_),
    .B(_1560_),
    .A_N(_1548_));
 sg13g2_a21oi_1 _4734_ (.A1(_1552_),
    .A2(_1559_),
    .Y(_0316_),
    .B1(_1561_));
 sg13g2_nand2_1 _4735_ (.Y(_1562_),
    .A(\mem[26][3] ),
    .B(\mem[10][0] ));
 sg13g2_o21ai_1 _4736_ (.B1(_1557_),
    .Y(_1563_),
    .A1(_1554_),
    .A2(_1558_));
 sg13g2_nand2_1 _4737_ (.Y(_1564_),
    .A(\mem[10][1] ),
    .B(\mem[26][2] ));
 sg13g2_nand2_1 _4738_ (.Y(_1565_),
    .A(\mem[10][3] ),
    .B(\mem[26][1] ));
 sg13g2_nand2_1 _4739_ (.Y(_1566_),
    .A(\mem[10][3] ),
    .B(\mem[26][0] ));
 sg13g2_xor2_1 _4740_ (.B(_1566_),
    .A(_1555_),
    .X(_1567_));
 sg13g2_nand2b_1 _4741_ (.Y(_1568_),
    .B(_1567_),
    .A_N(_1564_));
 sg13g2_xnor2_1 _4742_ (.Y(_1569_),
    .A(_1564_),
    .B(_1567_));
 sg13g2_nand2_1 _4743_ (.Y(_1570_),
    .A(_1563_),
    .B(_1569_));
 sg13g2_xnor2_1 _4744_ (.Y(_1571_),
    .A(_1563_),
    .B(_1569_));
 sg13g2_xnor2_1 _4745_ (.Y(_1572_),
    .A(_1562_),
    .B(_1571_));
 sg13g2_and2_1 _4746_ (.A(_1560_),
    .B(_1572_),
    .X(_1573_));
 sg13g2_nor2_1 _4747_ (.A(_1560_),
    .B(_1572_),
    .Y(_1574_));
 sg13g2_nor3_1 _4748_ (.A(_1548_),
    .B(_1573_),
    .C(_1574_),
    .Y(_0317_));
 sg13g2_o21ai_1 _4749_ (.B1(_1570_),
    .Y(_1575_),
    .A1(_1562_),
    .A2(_1571_));
 sg13g2_nand2_1 _4750_ (.Y(_1576_),
    .A(\mem[26][3] ),
    .B(\mem[10][1] ));
 sg13g2_o21ai_1 _4751_ (.B1(_1568_),
    .Y(_1577_),
    .A1(_1555_),
    .A2(_1566_));
 sg13g2_nand2_1 _4752_ (.Y(_1578_),
    .A(\mem[10][2] ),
    .B(\mem[26][2] ));
 sg13g2_nand2_1 _4753_ (.Y(_1579_),
    .A(net776),
    .B(net793));
 sg13g2_xor2_1 _4754_ (.B(_1578_),
    .A(_1565_),
    .X(_1580_));
 sg13g2_and2_1 _4755_ (.A(_1577_),
    .B(_1580_),
    .X(_1581_));
 sg13g2_xor2_1 _4756_ (.B(_1580_),
    .A(_1577_),
    .X(_1582_));
 sg13g2_nor2b_1 _4757_ (.A(_1576_),
    .B_N(_1582_),
    .Y(_1583_));
 sg13g2_xnor2_1 _4758_ (.Y(_1584_),
    .A(_1576_),
    .B(_1582_));
 sg13g2_nand2_1 _4759_ (.Y(_1585_),
    .A(_1575_),
    .B(_1584_));
 sg13g2_xor2_1 _4760_ (.B(_1584_),
    .A(_1575_),
    .X(_1586_));
 sg13g2_nand2_1 _4761_ (.Y(_1587_),
    .A(_1574_),
    .B(_1586_));
 sg13g2_a21oi_1 _4762_ (.A1(_1574_),
    .A2(_1586_),
    .Y(_1588_),
    .B1(_1548_));
 sg13g2_o21ai_1 _4763_ (.B1(_1588_),
    .Y(_1589_),
    .A1(_1574_),
    .A2(_1586_));
 sg13g2_inv_1 _4764_ (.Y(_0318_),
    .A(_1589_));
 sg13g2_nand2_1 _4765_ (.Y(_1590_),
    .A(\mem[26][3] ),
    .B(\mem[10][2] ));
 sg13g2_nand2b_1 _4766_ (.Y(_1591_),
    .B(_1555_),
    .A_N(_1579_));
 sg13g2_xor2_1 _4767_ (.B(_1591_),
    .A(_1590_),
    .X(_1592_));
 sg13g2_o21ai_1 _4768_ (.B1(_1592_),
    .Y(_1593_),
    .A1(_1581_),
    .A2(_1583_));
 sg13g2_or3_1 _4769_ (.A(_1581_),
    .B(_1583_),
    .C(_1592_),
    .X(_1594_));
 sg13g2_nand2_1 _4770_ (.Y(_1595_),
    .A(_1593_),
    .B(_1594_));
 sg13g2_and3_1 _4771_ (.X(_1596_),
    .A(_1585_),
    .B(_1587_),
    .C(_1595_));
 sg13g2_a21oi_1 _4772_ (.A1(_1585_),
    .A2(_1587_),
    .Y(_1597_),
    .B1(_1595_));
 sg13g2_nor3_1 _4773_ (.A(_1548_),
    .B(_1596_),
    .C(_1597_),
    .Y(_0319_));
 sg13g2_a21oi_2 _4774_ (.B1(_1579_),
    .Y(_1598_),
    .A2(_1590_),
    .A1(_1555_));
 sg13g2_nand2_1 _4775_ (.Y(_1599_),
    .A(net760),
    .B(net776));
 sg13g2_nand2b_1 _4776_ (.Y(_1600_),
    .B(_1598_),
    .A_N(_1599_));
 sg13g2_xor2_1 _4777_ (.B(_1599_),
    .A(_1598_),
    .X(_1601_));
 sg13g2_nand2_1 _4778_ (.Y(_1602_),
    .A(_1585_),
    .B(_1593_));
 sg13g2_nand2_1 _4779_ (.Y(_1603_),
    .A(_1594_),
    .B(_1602_));
 sg13g2_or2_1 _4780_ (.X(_1604_),
    .B(_1603_),
    .A(_1601_));
 sg13g2_nand2b_1 _4781_ (.Y(_1605_),
    .B(_1604_),
    .A_N(_1548_));
 sg13g2_a21oi_1 _4782_ (.A1(_1601_),
    .A2(_1603_),
    .Y(_0320_),
    .B1(_1605_));
 sg13g2_a21oi_1 _4783_ (.A1(_1600_),
    .A2(_1604_),
    .Y(_0321_),
    .B1(_1548_));
 sg13g2_a21oi_2 _4784_ (.B1(_1370_),
    .Y(_1606_),
    .A2(_1247_),
    .A1(_1188_));
 sg13g2_o21ai_1 _4785_ (.B1(_1369_),
    .Y(_1607_),
    .A1(_1187_),
    .A2(_1248_));
 sg13g2_and3_1 _4786_ (.X(_0322_),
    .A(net697),
    .B(\mem[25][0] ),
    .C(_1607_));
 sg13g2_a22oi_1 _4787_ (.Y(_1608_),
    .B1(\mem[25][1] ),
    .B2(net697),
    .A2(net753),
    .A1(\mem[25][0] ));
 sg13g2_nand4_1 _4788_ (.B(net782),
    .C(net753),
    .A(net697),
    .Y(_1609_),
    .D(\mem[25][1] ));
 sg13g2_inv_1 _4789_ (.Y(_1610_),
    .A(_1609_));
 sg13g2_nor3_1 _4790_ (.A(_1606_),
    .B(net754),
    .C(_1610_),
    .Y(_0323_));
 sg13g2_a22oi_1 _4791_ (.Y(_1611_),
    .B1(\mem[25][2] ),
    .B2(\mem[9][0] ),
    .A2(\mem[25][1] ),
    .A1(\mem[9][1] ));
 sg13g2_nand2_1 _4792_ (.Y(_1612_),
    .A(\mem[9][1] ),
    .B(\mem[25][2] ));
 sg13g2_and4_2 _4793_ (.A(\mem[9][0] ),
    .B(\mem[9][1] ),
    .C(\mem[25][1] ),
    .D(\mem[25][2] ),
    .X(_1613_));
 sg13g2_nor2_1 _4794_ (.A(_1611_),
    .B(_1613_),
    .Y(_1614_));
 sg13g2_nand2_1 _4795_ (.Y(_1615_),
    .A(\mem[25][0] ),
    .B(\mem[9][2] ));
 sg13g2_nor3_1 _4796_ (.A(_1611_),
    .B(_1613_),
    .C(_1615_),
    .Y(_1616_));
 sg13g2_xor2_1 _4797_ (.B(_1615_),
    .A(_1614_),
    .X(_1617_));
 sg13g2_and2_1 _4798_ (.A(_1609_),
    .B(_1617_),
    .X(_1618_));
 sg13g2_nor2_1 _4799_ (.A(_1609_),
    .B(_1617_),
    .Y(_1619_));
 sg13g2_nor3_1 _4800_ (.A(_1606_),
    .B(_1618_),
    .C(_1619_),
    .Y(_0324_));
 sg13g2_nand2_1 _4801_ (.Y(_1620_),
    .A(\mem[25][0] ),
    .B(\mem[9][3] ));
 sg13g2_nand2_1 _4802_ (.Y(_1621_),
    .A(\mem[25][1] ),
    .B(\mem[9][2] ));
 sg13g2_nand2_1 _4803_ (.Y(_1622_),
    .A(\mem[9][1] ),
    .B(\mem[25][3] ));
 sg13g2_nand2_1 _4804_ (.Y(_1623_),
    .A(\mem[9][0] ),
    .B(\mem[25][3] ));
 sg13g2_xor2_1 _4805_ (.B(_1623_),
    .A(_1612_),
    .X(_1624_));
 sg13g2_nand2b_1 _4806_ (.Y(_1625_),
    .B(_1624_),
    .A_N(_1621_));
 sg13g2_xnor2_1 _4807_ (.Y(_1626_),
    .A(_1621_),
    .B(_1624_));
 sg13g2_nand2_1 _4808_ (.Y(_1627_),
    .A(_1613_),
    .B(_1626_));
 sg13g2_xor2_1 _4809_ (.B(_1626_),
    .A(_1613_),
    .X(_1628_));
 sg13g2_nand2b_1 _4810_ (.Y(_1629_),
    .B(_1628_),
    .A_N(_1620_));
 sg13g2_xnor2_1 _4811_ (.Y(_1630_),
    .A(_1620_),
    .B(_1628_));
 sg13g2_and2_1 _4812_ (.A(_1616_),
    .B(_1630_),
    .X(_1631_));
 sg13g2_xor2_1 _4813_ (.B(_1630_),
    .A(_1616_),
    .X(_1632_));
 sg13g2_o21ai_1 _4814_ (.B1(_1607_),
    .Y(_1633_),
    .A1(_1619_),
    .A2(_1632_));
 sg13g2_a21oi_1 _4815_ (.A1(_1619_),
    .A2(_1632_),
    .Y(_0325_),
    .B1(_1633_));
 sg13g2_a21oi_1 _4816_ (.A1(_1619_),
    .A2(_1632_),
    .Y(_1634_),
    .B1(_1631_));
 sg13g2_o21ai_1 _4817_ (.B1(_1625_),
    .Y(_1635_),
    .A1(_1612_),
    .A2(_1623_));
 sg13g2_nand2_1 _4818_ (.Y(_1636_),
    .A(\mem[25][1] ),
    .B(\mem[9][3] ));
 sg13g2_nand2_1 _4819_ (.Y(_1637_),
    .A(\mem[9][2] ),
    .B(\mem[25][3] ));
 sg13g2_nand2_2 _4820_ (.Y(_1638_),
    .A(net740),
    .B(\mem[25][2] ));
 sg13g2_xor2_1 _4821_ (.B(_1638_),
    .A(_1622_),
    .X(_1639_));
 sg13g2_nand2b_1 _4822_ (.Y(_1640_),
    .B(_1639_),
    .A_N(_1636_));
 sg13g2_xnor2_1 _4823_ (.Y(_1641_),
    .A(_1636_),
    .B(_1639_));
 sg13g2_nand2_1 _4824_ (.Y(_1642_),
    .A(_1635_),
    .B(_1641_));
 sg13g2_xnor2_1 _4825_ (.Y(_1643_),
    .A(_1635_),
    .B(_1641_));
 sg13g2_a21o_1 _4826_ (.A2(_1629_),
    .A1(_1627_),
    .B1(_1643_),
    .X(_1644_));
 sg13g2_nand3_1 _4827_ (.B(_1629_),
    .C(_1643_),
    .A(_1627_),
    .Y(_1645_));
 sg13g2_nand2_1 _4828_ (.Y(_1646_),
    .A(_1644_),
    .B(_1645_));
 sg13g2_or2_1 _4829_ (.X(_1647_),
    .B(_1646_),
    .A(_1634_));
 sg13g2_nand2_1 _4830_ (.Y(_1648_),
    .A(_1607_),
    .B(_1647_));
 sg13g2_a21oi_1 _4831_ (.A1(_1634_),
    .A2(_1646_),
    .Y(_0326_),
    .B1(_1648_));
 sg13g2_nand2_1 _4832_ (.Y(_1649_),
    .A(_1644_),
    .B(_1647_));
 sg13g2_o21ai_1 _4833_ (.B1(_1640_),
    .Y(_1650_),
    .A1(_1622_),
    .A2(_1638_));
 sg13g2_nand2_1 _4834_ (.Y(_1651_),
    .A(\mem[25][2] ),
    .B(\mem[9][3] ));
 sg13g2_nand2_1 _4835_ (.Y(_1652_),
    .A(net720),
    .B(net718));
 sg13g2_xor2_1 _4836_ (.B(_1651_),
    .A(_1637_),
    .X(_1653_));
 sg13g2_nand2_1 _4837_ (.Y(_1654_),
    .A(_1650_),
    .B(_1653_));
 sg13g2_xnor2_1 _4838_ (.Y(_1655_),
    .A(_1650_),
    .B(_1653_));
 sg13g2_xor2_1 _4839_ (.B(_1655_),
    .A(_1642_),
    .X(_1656_));
 sg13g2_xnor2_1 _4840_ (.Y(_1657_),
    .A(_1649_),
    .B(_1656_));
 sg13g2_nor2_1 _4841_ (.A(_1606_),
    .B(_1657_),
    .Y(_0327_));
 sg13g2_nand2b_1 _4842_ (.Y(_1658_),
    .B(_1638_),
    .A_N(_1652_));
 sg13g2_xor2_1 _4843_ (.B(_1658_),
    .A(_1654_),
    .X(_1659_));
 sg13g2_and2_1 _4844_ (.A(_1642_),
    .B(_1644_),
    .X(_1660_));
 sg13g2_a21oi_1 _4845_ (.A1(_1634_),
    .A2(_1660_),
    .Y(_1661_),
    .B1(_1655_));
 sg13g2_xnor2_1 _4846_ (.Y(_1662_),
    .A(_1659_),
    .B(_1661_));
 sg13g2_nor2_1 _4847_ (.A(_1606_),
    .B(_1662_),
    .Y(_0328_));
 sg13g2_a21oi_1 _4848_ (.A1(_1638_),
    .A2(_1654_),
    .Y(_1663_),
    .B1(_1652_));
 sg13g2_a21oi_1 _4849_ (.A1(_1659_),
    .A2(_1661_),
    .Y(_1664_),
    .B1(_1663_));
 sg13g2_nor2_1 _4850_ (.A(_1606_),
    .B(_1664_),
    .Y(_0329_));
 sg13g2_a21oi_2 _4851_ (.B1(net483),
    .Y(_1665_),
    .A2(_0781_),
    .A1(_2090_));
 sg13g2_o21ai_1 _4852_ (.B1(_1191_),
    .Y(_1666_),
    .A1(net407),
    .A2(net486));
 sg13g2_and3_1 _4853_ (.X(_0330_),
    .A(net491),
    .B(net705),
    .C(_1666_));
 sg13g2_a22oi_1 _4854_ (.Y(_1667_),
    .B1(\mem[24][1] ),
    .B2(net491),
    .A2(net412),
    .A1(\mem[24][0] ));
 sg13g2_and4_1 _4855_ (.A(net491),
    .B(\mem[24][0] ),
    .C(net490),
    .D(\mem[24][1] ),
    .X(_1668_));
 sg13g2_nor3_2 _4856_ (.A(_1665_),
    .B(net413),
    .C(_1668_),
    .Y(_0331_));
 sg13g2_a22oi_1 _4857_ (.Y(_1669_),
    .B1(\mem[24][2] ),
    .B2(net491),
    .A2(\mem[24][1] ),
    .A1(net490));
 sg13g2_nand4_1 _4858_ (.B(net490),
    .C(\mem[24][1] ),
    .A(net491),
    .Y(_1670_),
    .D(\mem[24][2] ));
 sg13g2_nor2b_1 _4859_ (.A(_1669_),
    .B_N(_1670_),
    .Y(_1671_));
 sg13g2_and3_1 _4860_ (.X(_1672_),
    .A(\mem[24][0] ),
    .B(\mem[8][2] ),
    .C(_1671_));
 sg13g2_a21oi_1 _4861_ (.A1(\mem[24][0] ),
    .A2(\mem[8][2] ),
    .Y(_1673_),
    .B1(_1671_));
 sg13g2_nor2_1 _4862_ (.A(_1672_),
    .B(_1673_),
    .Y(_1674_));
 sg13g2_nor2_1 _4863_ (.A(_1668_),
    .B(_1674_),
    .Y(_1675_));
 sg13g2_nand2_2 _4864_ (.Y(_1676_),
    .A(_1668_),
    .B(_1674_));
 sg13g2_nand2_1 _4865_ (.Y(_1677_),
    .A(_1666_),
    .B(_1676_));
 sg13g2_nor2_2 _4866_ (.A(_1675_),
    .B(_1677_),
    .Y(_0332_));
 sg13g2_and2_1 _4867_ (.A(\mem[24][0] ),
    .B(\mem[8][3] ),
    .X(_1678_));
 sg13g2_nand2_1 _4868_ (.Y(_1679_),
    .A(\mem[24][1] ),
    .B(\mem[8][2] ));
 sg13g2_nand2_1 _4869_ (.Y(_1680_),
    .A(net490),
    .B(\mem[24][3] ));
 sg13g2_and4_1 _4870_ (.A(net491),
    .B(net490),
    .C(\mem[24][2] ),
    .D(\mem[24][3] ),
    .X(_1681_));
 sg13g2_a22oi_1 _4871_ (.Y(_1682_),
    .B1(\mem[24][3] ),
    .B2(net491),
    .A2(\mem[24][2] ),
    .A1(net490));
 sg13g2_nor3_1 _4872_ (.A(_1679_),
    .B(_1681_),
    .C(_1682_),
    .Y(_1683_));
 sg13g2_o21ai_1 _4873_ (.B1(_1679_),
    .Y(_1684_),
    .A1(_1681_),
    .A2(_1682_));
 sg13g2_nor2b_1 _4874_ (.A(_1683_),
    .B_N(_1684_),
    .Y(_1685_));
 sg13g2_nor2b_1 _4875_ (.A(_1670_),
    .B_N(_1685_),
    .Y(_1686_));
 sg13g2_xnor2_1 _4876_ (.Y(_1687_),
    .A(_1670_),
    .B(_1685_));
 sg13g2_xor2_1 _4877_ (.B(_1687_),
    .A(_1678_),
    .X(_1688_));
 sg13g2_nand2_1 _4878_ (.Y(_1689_),
    .A(_1672_),
    .B(_1688_));
 sg13g2_xnor2_1 _4879_ (.Y(_1690_),
    .A(_1672_),
    .B(_1688_));
 sg13g2_o21ai_1 _4880_ (.B1(_1666_),
    .Y(_1691_),
    .A1(_1676_),
    .A2(_1690_));
 sg13g2_a21oi_2 _4881_ (.B1(_1691_),
    .Y(_0333_),
    .A2(_1690_),
    .A1(_1676_));
 sg13g2_o21ai_1 _4882_ (.B1(_1689_),
    .Y(_1692_),
    .A1(_1676_),
    .A2(_1690_));
 sg13g2_or2_1 _4883_ (.X(_1693_),
    .B(_1683_),
    .A(_1681_));
 sg13g2_nand2_1 _4884_ (.Y(_1694_),
    .A(\mem[24][1] ),
    .B(\mem[8][3] ));
 sg13g2_nand2_1 _4885_ (.Y(_1695_),
    .A(\mem[8][2] ),
    .B(\mem[24][3] ));
 sg13g2_nand2_2 _4886_ (.Y(_1696_),
    .A(\mem[8][2] ),
    .B(\mem[24][2] ));
 sg13g2_xor2_1 _4887_ (.B(_1696_),
    .A(_1680_),
    .X(_1697_));
 sg13g2_nand2b_1 _4888_ (.Y(_1698_),
    .B(_1697_),
    .A_N(_1694_));
 sg13g2_xnor2_1 _4889_ (.Y(_1699_),
    .A(_1694_),
    .B(_1697_));
 sg13g2_nand2_1 _4890_ (.Y(_1700_),
    .A(_1693_),
    .B(_1699_));
 sg13g2_xor2_1 _4891_ (.B(_1699_),
    .A(_1693_),
    .X(_1701_));
 sg13g2_a21oi_1 _4892_ (.A1(_1678_),
    .A2(_1687_),
    .Y(_1702_),
    .B1(_1686_));
 sg13g2_nand2b_1 _4893_ (.Y(_1703_),
    .B(_1701_),
    .A_N(_1702_));
 sg13g2_xnor2_1 _4894_ (.Y(_1704_),
    .A(_1701_),
    .B(_1702_));
 sg13g2_or2_1 _4895_ (.X(_1705_),
    .B(_1704_),
    .A(_1692_));
 sg13g2_nand2_1 _4896_ (.Y(_1706_),
    .A(_1692_),
    .B(_1704_));
 sg13g2_and3_2 _4897_ (.X(_0334_),
    .A(_1666_),
    .B(_1705_),
    .C(_1706_));
 sg13g2_nor2b_1 _4898_ (.A(_1692_),
    .B_N(_1703_),
    .Y(_1707_));
 sg13g2_and2_1 _4899_ (.A(_1703_),
    .B(_1706_),
    .X(_1708_));
 sg13g2_o21ai_1 _4900_ (.B1(_1698_),
    .Y(_1709_),
    .A1(_1680_),
    .A2(_1696_));
 sg13g2_nand2_1 _4901_ (.Y(_1710_),
    .A(\mem[24][2] ),
    .B(\mem[8][3] ));
 sg13g2_nand2_1 _4902_ (.Y(_1711_),
    .A(\mem[8][3] ),
    .B(\mem[24][3] ));
 sg13g2_xor2_1 _4903_ (.B(_1710_),
    .A(_1695_),
    .X(_1712_));
 sg13g2_nand2_1 _4904_ (.Y(_1713_),
    .A(_1709_),
    .B(_1712_));
 sg13g2_xnor2_1 _4905_ (.Y(_1714_),
    .A(_1709_),
    .B(_1712_));
 sg13g2_xnor2_1 _4906_ (.Y(_1715_),
    .A(_1700_),
    .B(_1714_));
 sg13g2_o21ai_1 _4907_ (.B1(_1666_),
    .Y(_1716_),
    .A1(_1708_),
    .A2(_1715_));
 sg13g2_a21oi_2 _4908_ (.B1(_1716_),
    .Y(_0335_),
    .A2(_1715_),
    .A1(_1708_));
 sg13g2_a21oi_1 _4909_ (.A1(_1700_),
    .A2(_1707_),
    .Y(_1717_),
    .B1(_1714_));
 sg13g2_nand2b_1 _4910_ (.Y(_1718_),
    .B(_1696_),
    .A_N(_1711_));
 sg13g2_xor2_1 _4911_ (.B(_1718_),
    .A(_1713_),
    .X(_1719_));
 sg13g2_xnor2_1 _4912_ (.Y(_1720_),
    .A(_1717_),
    .B(_1719_));
 sg13g2_nor2_2 _4913_ (.A(_1665_),
    .B(_1720_),
    .Y(_0336_));
 sg13g2_a21oi_1 _4914_ (.A1(_1696_),
    .A2(_1713_),
    .Y(_1721_),
    .B1(_1711_));
 sg13g2_a21oi_1 _4915_ (.A1(_1717_),
    .A2(_1719_),
    .Y(_1722_),
    .B1(_1721_));
 sg13g2_nor2_2 _4916_ (.A(_1665_),
    .B(_1722_),
    .Y(_0337_));
 sg13g2_nor2b_1 _4917_ (.A(net492),
    .B_N(net493),
    .Y(_1723_));
 sg13g2_a21oi_2 _4918_ (.B1(net486),
    .Y(_1724_),
    .A2(_1189_),
    .A1(_1188_));
 sg13g2_a21o_2 _4919_ (.A2(_1189_),
    .A1(_1188_),
    .B1(net486),
    .X(_1725_));
 sg13g2_a21oi_2 _4920_ (.B1(_1725_),
    .Y(_1726_),
    .A2(_1723_),
    .A1(_1249_));
 sg13g2_a21o_2 _4921_ (.A2(_1723_),
    .A1(_1249_),
    .B1(_1725_),
    .X(_1727_));
 sg13g2_and3_1 _4922_ (.X(_0338_),
    .A(net707),
    .B(\mem[23][0] ),
    .C(_1726_));
 sg13g2_nand4_1 _4923_ (.B(\mem[23][0] ),
    .C(net791),
    .A(net859),
    .Y(_1728_),
    .D(\mem[23][1] ));
 sg13g2_inv_1 _4924_ (.Y(_1729_),
    .A(_1728_));
 sg13g2_a22oi_1 _4925_ (.Y(_1730_),
    .B1(\mem[23][1] ),
    .B2(net707),
    .A2(net763),
    .A1(\mem[23][0] ));
 sg13g2_nor3_1 _4926_ (.A(_1727_),
    .B(_1729_),
    .C(net764),
    .Y(_0339_));
 sg13g2_nand2_1 _4927_ (.Y(_1731_),
    .A(\mem[23][0] ),
    .B(\mem[7][2] ));
 sg13g2_a22oi_1 _4928_ (.Y(_1732_),
    .B1(\mem[23][2] ),
    .B2(\mem[7][0] ),
    .A2(\mem[23][1] ),
    .A1(\mem[7][1] ));
 sg13g2_nand2_1 _4929_ (.Y(_1733_),
    .A(\mem[7][1] ),
    .B(\mem[23][2] ));
 sg13g2_and4_1 _4930_ (.A(\mem[7][0] ),
    .B(\mem[7][1] ),
    .C(\mem[23][1] ),
    .D(\mem[23][2] ),
    .X(_1734_));
 sg13g2_nor2_1 _4931_ (.A(_1732_),
    .B(_1734_),
    .Y(_1735_));
 sg13g2_nor3_1 _4932_ (.A(_1731_),
    .B(_1732_),
    .C(_1734_),
    .Y(_1736_));
 sg13g2_xor2_1 _4933_ (.B(_1735_),
    .A(_1731_),
    .X(_1737_));
 sg13g2_and2_1 _4934_ (.A(_1728_),
    .B(_1737_),
    .X(_1738_));
 sg13g2_nor2_1 _4935_ (.A(_1728_),
    .B(_1737_),
    .Y(_1739_));
 sg13g2_nor3_1 _4936_ (.A(_1727_),
    .B(_1738_),
    .C(_1739_),
    .Y(_0340_));
 sg13g2_nand2_1 _4937_ (.Y(_1740_),
    .A(\mem[23][0] ),
    .B(\mem[7][3] ));
 sg13g2_nand2_1 _4938_ (.Y(_1741_),
    .A(\mem[23][1] ),
    .B(\mem[7][2] ));
 sg13g2_nand2_1 _4939_ (.Y(_1742_),
    .A(\mem[7][1] ),
    .B(\mem[23][3] ));
 sg13g2_nand2_1 _4940_ (.Y(_1743_),
    .A(\mem[7][0] ),
    .B(\mem[23][3] ));
 sg13g2_xor2_1 _4941_ (.B(_1743_),
    .A(_1733_),
    .X(_1744_));
 sg13g2_nand2b_1 _4942_ (.Y(_1745_),
    .B(_1744_),
    .A_N(_1741_));
 sg13g2_xnor2_1 _4943_ (.Y(_1746_),
    .A(_1741_),
    .B(_1744_));
 sg13g2_nand2_1 _4944_ (.Y(_1747_),
    .A(_1734_),
    .B(_1746_));
 sg13g2_xor2_1 _4945_ (.B(_1746_),
    .A(_1734_),
    .X(_1748_));
 sg13g2_nand2b_1 _4946_ (.Y(_1749_),
    .B(_1748_),
    .A_N(_1740_));
 sg13g2_xnor2_1 _4947_ (.Y(_1750_),
    .A(_1740_),
    .B(_1748_));
 sg13g2_and2_1 _4948_ (.A(_1736_),
    .B(_1750_),
    .X(_1751_));
 sg13g2_xor2_1 _4949_ (.B(_1750_),
    .A(_1736_),
    .X(_1752_));
 sg13g2_xnor2_1 _4950_ (.Y(_1753_),
    .A(_1739_),
    .B(_1752_));
 sg13g2_nor2_1 _4951_ (.A(_1727_),
    .B(_1753_),
    .Y(_0341_));
 sg13g2_a21oi_1 _4952_ (.A1(_1739_),
    .A2(_1752_),
    .Y(_1754_),
    .B1(_1751_));
 sg13g2_o21ai_1 _4953_ (.B1(_1745_),
    .Y(_1755_),
    .A1(_1733_),
    .A2(_1743_));
 sg13g2_nand2_1 _4954_ (.Y(_1756_),
    .A(\mem[23][1] ),
    .B(\mem[7][3] ));
 sg13g2_nand2_1 _4955_ (.Y(_1757_),
    .A(\mem[7][2] ),
    .B(\mem[23][3] ));
 sg13g2_nand2_2 _4956_ (.Y(_1758_),
    .A(\mem[7][2] ),
    .B(\mem[23][2] ));
 sg13g2_or2_1 _4957_ (.X(_1759_),
    .B(_1758_),
    .A(_1742_));
 sg13g2_xnor2_1 _4958_ (.Y(_1760_),
    .A(_1742_),
    .B(_1758_));
 sg13g2_xor2_1 _4959_ (.B(_1760_),
    .A(_1756_),
    .X(_1761_));
 sg13g2_nand2_1 _4960_ (.Y(_1762_),
    .A(_1755_),
    .B(_1761_));
 sg13g2_xnor2_1 _4961_ (.Y(_1763_),
    .A(_1755_),
    .B(_1761_));
 sg13g2_a21o_1 _4962_ (.A2(_1749_),
    .A1(_1747_),
    .B1(_1763_),
    .X(_1764_));
 sg13g2_nand3_1 _4963_ (.B(_1749_),
    .C(_1763_),
    .A(_1747_),
    .Y(_1765_));
 sg13g2_nand2_1 _4964_ (.Y(_1766_),
    .A(_1764_),
    .B(_1765_));
 sg13g2_or2_1 _4965_ (.X(_1767_),
    .B(_1766_),
    .A(_1754_));
 sg13g2_nand2_1 _4966_ (.Y(_1768_),
    .A(_1726_),
    .B(_1767_));
 sg13g2_a21oi_1 _4967_ (.A1(_1754_),
    .A2(_1766_),
    .Y(_0342_),
    .B1(_1768_));
 sg13g2_nand2_1 _4968_ (.Y(_1769_),
    .A(_1764_),
    .B(_1767_));
 sg13g2_o21ai_1 _4969_ (.B1(_1759_),
    .Y(_1770_),
    .A1(_1756_),
    .A2(_1760_));
 sg13g2_nand2_1 _4970_ (.Y(_1771_),
    .A(\mem[23][2] ),
    .B(\mem[7][3] ));
 sg13g2_nand2_1 _4971_ (.Y(_1772_),
    .A(net756),
    .B(net758));
 sg13g2_xor2_1 _4972_ (.B(_1771_),
    .A(_1757_),
    .X(_1773_));
 sg13g2_nand2_1 _4973_ (.Y(_1774_),
    .A(_1770_),
    .B(_1773_));
 sg13g2_xnor2_1 _4974_ (.Y(_1775_),
    .A(_1770_),
    .B(_1773_));
 sg13g2_xor2_1 _4975_ (.B(_1775_),
    .A(_1762_),
    .X(_1776_));
 sg13g2_xnor2_1 _4976_ (.Y(_1777_),
    .A(_1769_),
    .B(_1776_));
 sg13g2_nor2_1 _4977_ (.A(_1727_),
    .B(_1777_),
    .Y(_0343_));
 sg13g2_nand2b_1 _4978_ (.Y(_1778_),
    .B(_1758_),
    .A_N(_1772_));
 sg13g2_xor2_1 _4979_ (.B(_1778_),
    .A(_1774_),
    .X(_1779_));
 sg13g2_and2_1 _4980_ (.A(_1762_),
    .B(_1764_),
    .X(_1780_));
 sg13g2_a21oi_1 _4981_ (.A1(_1754_),
    .A2(_1780_),
    .Y(_1781_),
    .B1(_1775_));
 sg13g2_or2_1 _4982_ (.X(_1782_),
    .B(_1781_),
    .A(_1779_));
 sg13g2_nand2_1 _4983_ (.Y(_1783_),
    .A(_1779_),
    .B(_1781_));
 sg13g2_and3_1 _4984_ (.X(_0344_),
    .A(_1726_),
    .B(_1782_),
    .C(_1783_));
 sg13g2_a21o_1 _4985_ (.A2(_1774_),
    .A1(_1758_),
    .B1(_1772_),
    .X(_1784_));
 sg13g2_a21oi_1 _4986_ (.A1(_1783_),
    .A2(_1784_),
    .Y(_0345_),
    .B1(_1727_));
 sg13g2_nor2_2 _4987_ (.A(_1251_),
    .B(_1666_),
    .Y(_1785_));
 sg13g2_inv_1 _4988_ (.Y(_1786_),
    .A(_1785_));
 sg13g2_nand2_1 _4989_ (.Y(_1787_),
    .A(net725),
    .B(net783));
 sg13g2_nor2_1 _4990_ (.A(_1785_),
    .B(_1787_),
    .Y(_0346_));
 sg13g2_nand2_1 _4991_ (.Y(_1788_),
    .A(\mem[22][0] ),
    .B(\mem[6][1] ));
 sg13g2_a22oi_1 _4992_ (.Y(_1789_),
    .B1(\mem[22][1] ),
    .B2(net725),
    .A2(\mem[6][1] ),
    .A1(\mem[22][0] ));
 sg13g2_nand2_1 _4993_ (.Y(_1790_),
    .A(\mem[6][1] ),
    .B(\mem[22][1] ));
 sg13g2_nor2_1 _4994_ (.A(_1787_),
    .B(_1790_),
    .Y(_1791_));
 sg13g2_nor3_1 _4995_ (.A(_1785_),
    .B(net726),
    .C(_1791_),
    .Y(_0347_));
 sg13g2_and2_1 _4996_ (.A(net725),
    .B(net747),
    .X(_1792_));
 sg13g2_nand2_1 _4997_ (.Y(_1793_),
    .A(\mem[22][0] ),
    .B(net855));
 sg13g2_nor2b_1 _4998_ (.A(_1790_),
    .B_N(_1787_),
    .Y(_1794_));
 sg13g2_xnor2_1 _4999_ (.Y(_1795_),
    .A(_1793_),
    .B(_1794_));
 sg13g2_o21ai_1 _5000_ (.B1(_1786_),
    .Y(_1796_),
    .A1(_1792_),
    .A2(_1795_));
 sg13g2_a21oi_1 _5001_ (.A1(_1792_),
    .A2(_1795_),
    .Y(_0348_),
    .B1(_1796_));
 sg13g2_a22oi_1 _5002_ (.Y(_1797_),
    .B1(_1792_),
    .B2(_1795_),
    .A2(_1791_),
    .A1(_2102_));
 sg13g2_nand2_1 _5003_ (.Y(_1798_),
    .A(\mem[6][1] ),
    .B(\mem[22][2] ));
 sg13g2_a22oi_1 _5004_ (.Y(_1799_),
    .B1(\mem[22][3] ),
    .B2(\mem[6][0] ),
    .A2(\mem[6][3] ),
    .A1(\mem[22][0] ));
 sg13g2_nand4_1 _5005_ (.B(\mem[22][0] ),
    .C(\mem[6][3] ),
    .A(\mem[6][0] ),
    .Y(_1800_),
    .D(\mem[22][3] ));
 sg13g2_nor2b_1 _5006_ (.A(_1799_),
    .B_N(_1800_),
    .Y(_1801_));
 sg13g2_nand2_1 _5007_ (.Y(_1802_),
    .A(\mem[22][1] ),
    .B(\mem[6][2] ));
 sg13g2_nor2b_1 _5008_ (.A(_1802_),
    .B_N(_1788_),
    .Y(_1803_));
 sg13g2_xnor2_1 _5009_ (.Y(_1804_),
    .A(_1801_),
    .B(_1803_));
 sg13g2_nor2_1 _5010_ (.A(_1798_),
    .B(_1804_),
    .Y(_1805_));
 sg13g2_xnor2_1 _5011_ (.Y(_1806_),
    .A(_1798_),
    .B(_1804_));
 sg13g2_and2_1 _5012_ (.A(_1797_),
    .B(_1806_),
    .X(_1807_));
 sg13g2_nor2_1 _5013_ (.A(_1797_),
    .B(_1806_),
    .Y(_1808_));
 sg13g2_nor3_1 _5014_ (.A(_1785_),
    .B(_1807_),
    .C(_1808_),
    .Y(_0349_));
 sg13g2_nor3_1 _5015_ (.A(_1788_),
    .B(_1801_),
    .C(_1802_),
    .Y(_1809_));
 sg13g2_nand2_1 _5016_ (.Y(_1810_),
    .A(\mem[6][2] ),
    .B(\mem[22][2] ));
 sg13g2_a22oi_1 _5017_ (.Y(_1811_),
    .B1(\mem[22][3] ),
    .B2(\mem[6][1] ),
    .A2(\mem[6][3] ),
    .A1(\mem[22][1] ));
 sg13g2_nand4_1 _5018_ (.B(\mem[22][1] ),
    .C(\mem[6][3] ),
    .A(\mem[6][1] ),
    .Y(_1812_),
    .D(\mem[22][3] ));
 sg13g2_nand2b_1 _5019_ (.Y(_1813_),
    .B(_1812_),
    .A_N(_1811_));
 sg13g2_a21oi_1 _5020_ (.A1(_1800_),
    .A2(_1802_),
    .Y(_1814_),
    .B1(_1799_));
 sg13g2_nand2b_1 _5021_ (.Y(_1815_),
    .B(_1814_),
    .A_N(_1813_));
 sg13g2_xor2_1 _5022_ (.B(_1814_),
    .A(_1813_),
    .X(_1816_));
 sg13g2_xor2_1 _5023_ (.B(_1816_),
    .A(_1810_),
    .X(_1817_));
 sg13g2_nor3_1 _5024_ (.A(_1805_),
    .B(_1809_),
    .C(_1817_),
    .Y(_1818_));
 sg13g2_o21ai_1 _5025_ (.B1(_1817_),
    .Y(_1819_),
    .A1(_1805_),
    .A2(_1809_));
 sg13g2_nor2b_1 _5026_ (.A(_1818_),
    .B_N(_1819_),
    .Y(_1820_));
 sg13g2_o21ai_1 _5027_ (.B1(_1786_),
    .Y(_1821_),
    .A1(_1808_),
    .A2(_1820_));
 sg13g2_a21oi_1 _5028_ (.A1(_1808_),
    .A2(_1820_),
    .Y(_0350_),
    .B1(_1821_));
 sg13g2_nand2b_1 _5029_ (.Y(_1822_),
    .B(_1819_),
    .A_N(_1808_));
 sg13g2_nand2b_1 _5030_ (.Y(_1823_),
    .B(_1822_),
    .A_N(_1818_));
 sg13g2_nor2_1 _5031_ (.A(_2102_),
    .B(_1812_),
    .Y(_1824_));
 sg13g2_nand2_1 _5032_ (.Y(_1825_),
    .A(\mem[6][2] ),
    .B(\mem[22][3] ));
 sg13g2_a21o_1 _5033_ (.A2(_1825_),
    .A1(_1812_),
    .B1(_1824_),
    .X(_1826_));
 sg13g2_nand2_1 _5034_ (.Y(_1827_),
    .A(\mem[22][2] ),
    .B(\mem[6][3] ));
 sg13g2_nor2_1 _5035_ (.A(_1826_),
    .B(_1827_),
    .Y(_1828_));
 sg13g2_xor2_1 _5036_ (.B(_1827_),
    .A(_1826_),
    .X(_1829_));
 sg13g2_o21ai_1 _5037_ (.B1(_1815_),
    .Y(_1830_),
    .A1(_1810_),
    .A2(_1816_));
 sg13g2_nand2_1 _5038_ (.Y(_1831_),
    .A(_1829_),
    .B(_1830_));
 sg13g2_or2_1 _5039_ (.X(_1832_),
    .B(_1830_),
    .A(_1829_));
 sg13g2_nand2_1 _5040_ (.Y(_1833_),
    .A(_1831_),
    .B(_1832_));
 sg13g2_xnor2_1 _5041_ (.Y(_1834_),
    .A(_1823_),
    .B(_1833_));
 sg13g2_nor2_1 _5042_ (.A(_1785_),
    .B(_1834_),
    .Y(_0351_));
 sg13g2_nor2_1 _5043_ (.A(_1824_),
    .B(_1828_),
    .Y(_1835_));
 sg13g2_nand3_1 _5044_ (.B(\mem[22][3] ),
    .C(_1835_),
    .A(net752),
    .Y(_1836_));
 sg13g2_nand2_1 _5045_ (.Y(_1837_),
    .A(_1822_),
    .B(_1832_));
 sg13g2_nand2_1 _5046_ (.Y(_1838_),
    .A(_1831_),
    .B(_1837_));
 sg13g2_nand3_1 _5047_ (.B(_1836_),
    .C(_1837_),
    .A(_1831_),
    .Y(_1839_));
 sg13g2_nand2b_1 _5048_ (.Y(_1840_),
    .B(_1838_),
    .A_N(_1836_));
 sg13g2_and3_1 _5049_ (.X(_0352_),
    .A(_1786_),
    .B(_1839_),
    .C(_1840_));
 sg13g2_a21oi_1 _5050_ (.A1(_1835_),
    .A2(_1840_),
    .Y(_0353_),
    .B1(_1785_));
 sg13g2_a21o_2 _5051_ (.A2(_1723_),
    .A1(_1187_),
    .B1(_1725_),
    .X(_1841_));
 sg13g2_inv_1 _5052_ (.Y(_1842_),
    .A(_1841_));
 sg13g2_and3_1 _5053_ (.X(_0354_),
    .A(net409),
    .B(\mem[21][0] ),
    .C(_1842_));
 sg13g2_nand4_1 _5054_ (.B(\mem[21][0] ),
    .C(net820),
    .A(net495),
    .Y(_1843_),
    .D(\mem[21][1] ));
 sg13g2_inv_1 _5055_ (.Y(_1844_),
    .A(_1843_));
 sg13g2_a22oi_1 _5056_ (.Y(_1845_),
    .B1(net815),
    .B2(net495),
    .A2(net494),
    .A1(\mem[21][0] ));
 sg13g2_nor3_1 _5057_ (.A(_1841_),
    .B(_1844_),
    .C(net816),
    .Y(_0355_));
 sg13g2_a22oi_1 _5058_ (.Y(_1846_),
    .B1(\mem[21][2] ),
    .B2(net495),
    .A2(\mem[21][1] ),
    .A1(net494));
 sg13g2_nand4_1 _5059_ (.B(net494),
    .C(\mem[21][1] ),
    .A(net495),
    .Y(_1847_),
    .D(\mem[21][2] ));
 sg13g2_nor2b_1 _5060_ (.A(_1846_),
    .B_N(_1847_),
    .Y(_1848_));
 sg13g2_and3_1 _5061_ (.X(_1849_),
    .A(\mem[21][0] ),
    .B(\mem[5][2] ),
    .C(_1848_));
 sg13g2_a21oi_1 _5062_ (.A1(\mem[21][0] ),
    .A2(\mem[5][2] ),
    .Y(_1850_),
    .B1(_1848_));
 sg13g2_or2_1 _5063_ (.X(_1851_),
    .B(_1850_),
    .A(_1849_));
 sg13g2_and2_1 _5064_ (.A(_1843_),
    .B(_1851_),
    .X(_1852_));
 sg13g2_nor2_2 _5065_ (.A(_1843_),
    .B(_1851_),
    .Y(_1853_));
 sg13g2_nor3_1 _5066_ (.A(_1841_),
    .B(_1852_),
    .C(_1853_),
    .Y(_0356_));
 sg13g2_and2_1 _5067_ (.A(\mem[21][0] ),
    .B(\mem[5][3] ),
    .X(_1854_));
 sg13g2_nand2_1 _5068_ (.Y(_1855_),
    .A(\mem[21][1] ),
    .B(\mem[5][2] ));
 sg13g2_nand2_1 _5069_ (.Y(_1856_),
    .A(net494),
    .B(\mem[21][3] ));
 sg13g2_and4_1 _5070_ (.A(net495),
    .B(net494),
    .C(\mem[21][2] ),
    .D(\mem[21][3] ),
    .X(_1857_));
 sg13g2_a22oi_1 _5071_ (.Y(_1858_),
    .B1(\mem[21][3] ),
    .B2(net495),
    .A2(\mem[21][2] ),
    .A1(net494));
 sg13g2_nor3_1 _5072_ (.A(_1855_),
    .B(_1857_),
    .C(_1858_),
    .Y(_1859_));
 sg13g2_o21ai_1 _5073_ (.B1(_1855_),
    .Y(_1860_),
    .A1(_1857_),
    .A2(_1858_));
 sg13g2_nor2b_1 _5074_ (.A(_1859_),
    .B_N(_1860_),
    .Y(_1861_));
 sg13g2_nor2b_1 _5075_ (.A(_1847_),
    .B_N(_1861_),
    .Y(_1862_));
 sg13g2_xnor2_1 _5076_ (.Y(_1863_),
    .A(_1847_),
    .B(_1861_));
 sg13g2_xor2_1 _5077_ (.B(_1863_),
    .A(_1854_),
    .X(_1864_));
 sg13g2_and2_1 _5078_ (.A(_1849_),
    .B(_1864_),
    .X(_1865_));
 sg13g2_xor2_1 _5079_ (.B(_1864_),
    .A(_1849_),
    .X(_1866_));
 sg13g2_o21ai_1 _5080_ (.B1(_1842_),
    .Y(_1867_),
    .A1(_1853_),
    .A2(_1866_));
 sg13g2_a21oi_1 _5081_ (.A1(_1853_),
    .A2(_1866_),
    .Y(_0357_),
    .B1(_1867_));
 sg13g2_a21o_1 _5082_ (.A2(_1866_),
    .A1(_1853_),
    .B1(_1865_),
    .X(_1868_));
 sg13g2_or2_1 _5083_ (.X(_1869_),
    .B(_1859_),
    .A(_1857_));
 sg13g2_nand2_1 _5084_ (.Y(_1870_),
    .A(\mem[21][1] ),
    .B(\mem[5][3] ));
 sg13g2_nand2_1 _5085_ (.Y(_1871_),
    .A(\mem[5][2] ),
    .B(\mem[21][3] ));
 sg13g2_nand2_2 _5086_ (.Y(_1872_),
    .A(\mem[5][2] ),
    .B(\mem[21][2] ));
 sg13g2_xor2_1 _5087_ (.B(_1872_),
    .A(_1856_),
    .X(_1873_));
 sg13g2_nand2b_1 _5088_ (.Y(_1874_),
    .B(_1873_),
    .A_N(_1870_));
 sg13g2_xnor2_1 _5089_ (.Y(_1875_),
    .A(_1870_),
    .B(_1873_));
 sg13g2_nand2_1 _5090_ (.Y(_1876_),
    .A(_1869_),
    .B(_1875_));
 sg13g2_xor2_1 _5091_ (.B(_1875_),
    .A(_1869_),
    .X(_1877_));
 sg13g2_a21oi_1 _5092_ (.A1(_1854_),
    .A2(_1863_),
    .Y(_1878_),
    .B1(_1862_));
 sg13g2_nand2b_1 _5093_ (.Y(_1879_),
    .B(_1877_),
    .A_N(_1878_));
 sg13g2_xnor2_1 _5094_ (.Y(_1880_),
    .A(_1877_),
    .B(_1878_));
 sg13g2_or2_1 _5095_ (.X(_1881_),
    .B(_1880_),
    .A(_1868_));
 sg13g2_nand2_1 _5096_ (.Y(_1882_),
    .A(_1868_),
    .B(_1880_));
 sg13g2_and3_1 _5097_ (.X(_0358_),
    .A(_1842_),
    .B(_1881_),
    .C(_1882_));
 sg13g2_nor2b_1 _5098_ (.A(_1868_),
    .B_N(_1879_),
    .Y(_1883_));
 sg13g2_nand2_1 _5099_ (.Y(_1884_),
    .A(_1879_),
    .B(_1882_));
 sg13g2_o21ai_1 _5100_ (.B1(_1874_),
    .Y(_1885_),
    .A1(_1856_),
    .A2(_1872_));
 sg13g2_nand2_1 _5101_ (.Y(_1886_),
    .A(\mem[21][2] ),
    .B(\mem[5][3] ));
 sg13g2_nand2_1 _5102_ (.Y(_1887_),
    .A(net805),
    .B(net850));
 sg13g2_xor2_1 _5103_ (.B(_1886_),
    .A(_1871_),
    .X(_1888_));
 sg13g2_nand2_1 _5104_ (.Y(_1889_),
    .A(_1885_),
    .B(_1888_));
 sg13g2_xnor2_1 _5105_ (.Y(_1890_),
    .A(_1885_),
    .B(_1888_));
 sg13g2_xor2_1 _5106_ (.B(_1890_),
    .A(_1876_),
    .X(_1891_));
 sg13g2_xnor2_1 _5107_ (.Y(_1892_),
    .A(_1884_),
    .B(_1891_));
 sg13g2_nor2_1 _5108_ (.A(_1841_),
    .B(_1892_),
    .Y(_0359_));
 sg13g2_a21oi_1 _5109_ (.A1(_1876_),
    .A2(_1883_),
    .Y(_1893_),
    .B1(_1890_));
 sg13g2_nand2b_1 _5110_ (.Y(_1894_),
    .B(_1872_),
    .A_N(_1887_));
 sg13g2_xor2_1 _5111_ (.B(_1894_),
    .A(_1889_),
    .X(_1895_));
 sg13g2_xnor2_1 _5112_ (.Y(_1896_),
    .A(_1893_),
    .B(_1895_));
 sg13g2_nor2_1 _5113_ (.A(_1841_),
    .B(_1896_),
    .Y(_0360_));
 sg13g2_a21oi_1 _5114_ (.A1(_1872_),
    .A2(_1889_),
    .Y(_1897_),
    .B1(_1887_));
 sg13g2_a21oi_1 _5115_ (.A1(_1893_),
    .A2(_1895_),
    .Y(_1898_),
    .B1(_1897_));
 sg13g2_nor2_1 _5116_ (.A(_1841_),
    .B(_1898_),
    .Y(_0361_));
 sg13g2_nand2_1 _5117_ (.Y(_1899_),
    .A(net680),
    .B(net745));
 sg13g2_nor2_1 _5118_ (.A(_1725_),
    .B(net681),
    .Y(_0362_));
 sg13g2_nor3_2 _5119_ (.A(_2099_),
    .B(_2100_),
    .C(_1899_),
    .Y(_1900_));
 sg13g2_a22oi_1 _5120_ (.Y(_1901_),
    .B1(net688),
    .B2(net680),
    .A2(\mem[4][1] ),
    .A1(\mem[20][0] ));
 sg13g2_nor3_1 _5121_ (.A(_1725_),
    .B(_1900_),
    .C(net689),
    .Y(_0363_));
 sg13g2_a22oi_1 _5122_ (.Y(_1902_),
    .B1(\mem[20][2] ),
    .B2(\mem[4][0] ),
    .A2(\mem[20][1] ),
    .A1(\mem[4][1] ));
 sg13g2_nand4_1 _5123_ (.B(\mem[4][1] ),
    .C(\mem[20][1] ),
    .A(\mem[4][0] ),
    .Y(_1903_),
    .D(\mem[20][2] ));
 sg13g2_nor2b_1 _5124_ (.A(_1902_),
    .B_N(_1903_),
    .Y(_1904_));
 sg13g2_and3_1 _5125_ (.X(_1905_),
    .A(\mem[20][0] ),
    .B(\mem[4][2] ),
    .C(_1904_));
 sg13g2_a21oi_1 _5126_ (.A1(net745),
    .A2(\mem[4][2] ),
    .Y(_1906_),
    .B1(_1904_));
 sg13g2_nor2_1 _5127_ (.A(_1905_),
    .B(_1906_),
    .Y(_1907_));
 sg13g2_nor2_1 _5128_ (.A(_1900_),
    .B(_1907_),
    .Y(_1908_));
 sg13g2_nand2_1 _5129_ (.Y(_1909_),
    .A(_1900_),
    .B(_1907_));
 sg13g2_nand2_1 _5130_ (.Y(_1910_),
    .A(_1724_),
    .B(_1909_));
 sg13g2_nor2_1 _5131_ (.A(_1908_),
    .B(_1910_),
    .Y(_0364_));
 sg13g2_and2_1 _5132_ (.A(\mem[20][0] ),
    .B(\mem[4][3] ),
    .X(_1911_));
 sg13g2_nand2_1 _5133_ (.Y(_1912_),
    .A(\mem[20][1] ),
    .B(\mem[4][2] ));
 sg13g2_nand2_2 _5134_ (.Y(_1913_),
    .A(\mem[4][1] ),
    .B(\mem[20][3] ));
 sg13g2_nor3_1 _5135_ (.A(_2096_),
    .B(_2103_),
    .C(_1913_),
    .Y(_1914_));
 sg13g2_a22oi_1 _5136_ (.Y(_1915_),
    .B1(\mem[20][3] ),
    .B2(\mem[4][0] ),
    .A2(\mem[20][2] ),
    .A1(\mem[4][1] ));
 sg13g2_nor3_1 _5137_ (.A(_1912_),
    .B(_1914_),
    .C(_1915_),
    .Y(_1916_));
 sg13g2_o21ai_1 _5138_ (.B1(_1912_),
    .Y(_1917_),
    .A1(_1914_),
    .A2(_1915_));
 sg13g2_nor2b_1 _5139_ (.A(_1916_),
    .B_N(_1917_),
    .Y(_1918_));
 sg13g2_nor2b_1 _5140_ (.A(_1903_),
    .B_N(_1918_),
    .Y(_1919_));
 sg13g2_xnor2_1 _5141_ (.Y(_1920_),
    .A(_1903_),
    .B(_1918_));
 sg13g2_xor2_1 _5142_ (.B(_1920_),
    .A(_1911_),
    .X(_1921_));
 sg13g2_nand2_1 _5143_ (.Y(_1922_),
    .A(_1905_),
    .B(_1921_));
 sg13g2_xnor2_1 _5144_ (.Y(_1923_),
    .A(_1905_),
    .B(_1921_));
 sg13g2_o21ai_1 _5145_ (.B1(_1724_),
    .Y(_1924_),
    .A1(_1909_),
    .A2(_1923_));
 sg13g2_a21oi_1 _5146_ (.A1(_1909_),
    .A2(_1923_),
    .Y(_0365_),
    .B1(_1924_));
 sg13g2_o21ai_1 _5147_ (.B1(_1922_),
    .Y(_1925_),
    .A1(_1909_),
    .A2(_1923_));
 sg13g2_or2_1 _5148_ (.X(_1926_),
    .B(_1916_),
    .A(_1914_));
 sg13g2_nand2_1 _5149_ (.Y(_1927_),
    .A(\mem[20][1] ),
    .B(\mem[4][3] ));
 sg13g2_nand2_1 _5150_ (.Y(_1928_),
    .A(\mem[4][2] ),
    .B(\mem[20][3] ));
 sg13g2_nand2_2 _5151_ (.Y(_1929_),
    .A(\mem[4][2] ),
    .B(\mem[20][2] ));
 sg13g2_xor2_1 _5152_ (.B(_1929_),
    .A(_1913_),
    .X(_1930_));
 sg13g2_nand2b_1 _5153_ (.Y(_1931_),
    .B(_1930_),
    .A_N(_1927_));
 sg13g2_xnor2_1 _5154_ (.Y(_1932_),
    .A(_1927_),
    .B(_1930_));
 sg13g2_nand2_1 _5155_ (.Y(_1933_),
    .A(_1926_),
    .B(_1932_));
 sg13g2_xor2_1 _5156_ (.B(_1932_),
    .A(_1926_),
    .X(_1934_));
 sg13g2_a21oi_1 _5157_ (.A1(_1911_),
    .A2(_1920_),
    .Y(_1935_),
    .B1(_1919_));
 sg13g2_nand2b_1 _5158_ (.Y(_1936_),
    .B(_1934_),
    .A_N(_1935_));
 sg13g2_xnor2_1 _5159_ (.Y(_1937_),
    .A(_1934_),
    .B(_1935_));
 sg13g2_or2_1 _5160_ (.X(_1938_),
    .B(_1937_),
    .A(_1925_));
 sg13g2_nand2_1 _5161_ (.Y(_1939_),
    .A(_1925_),
    .B(_1937_));
 sg13g2_and3_1 _5162_ (.X(_0366_),
    .A(_1724_),
    .B(_1938_),
    .C(_1939_));
 sg13g2_nor2b_1 _5163_ (.A(_1925_),
    .B_N(_1936_),
    .Y(_1940_));
 sg13g2_o21ai_1 _5164_ (.B1(_1931_),
    .Y(_1941_),
    .A1(_1913_),
    .A2(_1929_));
 sg13g2_nand2_1 _5165_ (.Y(_1942_),
    .A(\mem[20][2] ),
    .B(\mem[4][3] ));
 sg13g2_nand2_1 _5166_ (.Y(_1943_),
    .A(net742),
    .B(\mem[20][3] ));
 sg13g2_xor2_1 _5167_ (.B(_1942_),
    .A(_1928_),
    .X(_1944_));
 sg13g2_nand2_1 _5168_ (.Y(_1945_),
    .A(_1941_),
    .B(_1944_));
 sg13g2_xnor2_1 _5169_ (.Y(_1946_),
    .A(_1941_),
    .B(_1944_));
 sg13g2_xnor2_1 _5170_ (.Y(_1947_),
    .A(_1933_),
    .B(_1946_));
 sg13g2_and3_1 _5171_ (.X(_1948_),
    .A(_1936_),
    .B(_1939_),
    .C(_1947_));
 sg13g2_a21oi_1 _5172_ (.A1(_1936_),
    .A2(_1939_),
    .Y(_1949_),
    .B1(_1947_));
 sg13g2_nor3_1 _5173_ (.A(_1725_),
    .B(_1948_),
    .C(_1949_),
    .Y(_0367_));
 sg13g2_a21oi_1 _5174_ (.A1(_1933_),
    .A2(_1940_),
    .Y(_1950_),
    .B1(_1946_));
 sg13g2_nand2b_1 _5175_ (.Y(_1951_),
    .B(_1929_),
    .A_N(_1943_));
 sg13g2_xor2_1 _5176_ (.B(_1951_),
    .A(_1945_),
    .X(_1952_));
 sg13g2_or2_1 _5177_ (.X(_1953_),
    .B(_1952_),
    .A(_1950_));
 sg13g2_nand2_1 _5178_ (.Y(_1954_),
    .A(_1950_),
    .B(_1952_));
 sg13g2_and3_1 _5179_ (.X(_0368_),
    .A(_1724_),
    .B(_1953_),
    .C(_1954_));
 sg13g2_a21o_1 _5180_ (.A2(_1945_),
    .A1(_1929_),
    .B1(_1943_),
    .X(_1955_));
 sg13g2_a21oi_1 _5181_ (.A1(_1954_),
    .A2(_1955_),
    .Y(_0369_),
    .B1(_1725_));
 sg13g2_nor2_2 _5182_ (.A(_1250_),
    .B(_1724_),
    .Y(_1956_));
 sg13g2_inv_1 _5183_ (.Y(_1957_),
    .A(_1956_));
 sg13g2_nand2_1 _5184_ (.Y(_1958_),
    .A(net676),
    .B(\mem[19][0] ));
 sg13g2_nor2_1 _5185_ (.A(_1956_),
    .B(net677),
    .Y(_0370_));
 sg13g2_a22oi_1 _5186_ (.Y(_1959_),
    .B1(net701),
    .B2(net676),
    .A2(\mem[3][1] ),
    .A1(\mem[19][0] ));
 sg13g2_nand2_1 _5187_ (.Y(_1960_),
    .A(\mem[3][1] ),
    .B(\mem[19][1] ));
 sg13g2_or2_1 _5188_ (.X(_1961_),
    .B(_1960_),
    .A(_1958_));
 sg13g2_inv_1 _5189_ (.Y(_1962_),
    .A(_1961_));
 sg13g2_nor3_1 _5190_ (.A(_1956_),
    .B(net702),
    .C(_1962_),
    .Y(_0371_));
 sg13g2_nand2_1 _5191_ (.Y(_1963_),
    .A(net856),
    .B(\mem[19][2] ));
 sg13g2_nand2_2 _5192_ (.Y(_1964_),
    .A(\mem[19][1] ),
    .B(\mem[3][2] ));
 sg13g2_nand2_1 _5193_ (.Y(_1965_),
    .A(\mem[19][0] ),
    .B(\mem[3][2] ));
 sg13g2_or2_1 _5194_ (.X(_1966_),
    .B(_1965_),
    .A(_1960_));
 sg13g2_xnor2_1 _5195_ (.Y(_1967_),
    .A(_1960_),
    .B(_1965_));
 sg13g2_xnor2_1 _5196_ (.Y(_1968_),
    .A(net857),
    .B(_1967_));
 sg13g2_or2_1 _5197_ (.X(_1969_),
    .B(_1968_),
    .A(_1961_));
 sg13g2_nand2_1 _5198_ (.Y(_1970_),
    .A(_1957_),
    .B(_1969_));
 sg13g2_a21oi_1 _5199_ (.A1(_1961_),
    .A2(_1968_),
    .Y(_0372_),
    .B1(_1970_));
 sg13g2_nand2_1 _5200_ (.Y(_1971_),
    .A(\mem[3][0] ),
    .B(\mem[19][3] ));
 sg13g2_o21ai_1 _5201_ (.B1(_1966_),
    .Y(_1972_),
    .A1(_1963_),
    .A2(_1967_));
 sg13g2_nand2_1 _5202_ (.Y(_1973_),
    .A(\mem[3][1] ),
    .B(\mem[19][2] ));
 sg13g2_nand2_1 _5203_ (.Y(_1974_),
    .A(\mem[19][1] ),
    .B(\mem[3][3] ));
 sg13g2_nand2_1 _5204_ (.Y(_1975_),
    .A(\mem[19][0] ),
    .B(\mem[3][3] ));
 sg13g2_xor2_1 _5205_ (.B(_1975_),
    .A(_1964_),
    .X(_1976_));
 sg13g2_nand2b_1 _5206_ (.Y(_1977_),
    .B(_1976_),
    .A_N(_1973_));
 sg13g2_xnor2_1 _5207_ (.Y(_1978_),
    .A(_1973_),
    .B(_1976_));
 sg13g2_nand2_1 _5208_ (.Y(_1979_),
    .A(_1972_),
    .B(_1978_));
 sg13g2_xnor2_1 _5209_ (.Y(_1980_),
    .A(_1972_),
    .B(_1978_));
 sg13g2_xnor2_1 _5210_ (.Y(_1981_),
    .A(_1971_),
    .B(_1980_));
 sg13g2_nor2_1 _5211_ (.A(_1969_),
    .B(_1981_),
    .Y(_1982_));
 sg13g2_a21oi_1 _5212_ (.A1(_1969_),
    .A2(_1981_),
    .Y(_1983_),
    .B1(_1956_));
 sg13g2_nor2b_1 _5213_ (.A(_1982_),
    .B_N(_1983_),
    .Y(_0373_));
 sg13g2_nand2_1 _5214_ (.Y(_1984_),
    .A(\mem[3][1] ),
    .B(\mem[19][3] ));
 sg13g2_o21ai_1 _5215_ (.B1(_1977_),
    .Y(_1985_),
    .A1(_1964_),
    .A2(_1975_));
 sg13g2_nand2_1 _5216_ (.Y(_1986_),
    .A(\mem[3][2] ),
    .B(\mem[19][2] ));
 sg13g2_nand2_1 _5217_ (.Y(_1987_),
    .A(net808),
    .B(net755));
 sg13g2_xor2_1 _5218_ (.B(_1986_),
    .A(_1974_),
    .X(_1988_));
 sg13g2_and2_1 _5219_ (.A(_1985_),
    .B(_1988_),
    .X(_1989_));
 sg13g2_xor2_1 _5220_ (.B(_1988_),
    .A(_1985_),
    .X(_1990_));
 sg13g2_nor2b_1 _5221_ (.A(_1984_),
    .B_N(_1990_),
    .Y(_1991_));
 sg13g2_xnor2_1 _5222_ (.Y(_1992_),
    .A(_1984_),
    .B(_1990_));
 sg13g2_o21ai_1 _5223_ (.B1(_1979_),
    .Y(_1993_),
    .A1(_1971_),
    .A2(_1980_));
 sg13g2_nand2_1 _5224_ (.Y(_1994_),
    .A(_1992_),
    .B(_1993_));
 sg13g2_xor2_1 _5225_ (.B(_1993_),
    .A(_1992_),
    .X(_1995_));
 sg13g2_nand2_1 _5226_ (.Y(_1996_),
    .A(_1982_),
    .B(_1995_));
 sg13g2_o21ai_1 _5227_ (.B1(_1957_),
    .Y(_1997_),
    .A1(_1982_),
    .A2(_1995_));
 sg13g2_nor2b_1 _5228_ (.A(_1997_),
    .B_N(_1996_),
    .Y(_0374_));
 sg13g2_nand2b_1 _5229_ (.Y(_1998_),
    .B(_1964_),
    .A_N(_1987_));
 sg13g2_nand2_1 _5230_ (.Y(_1999_),
    .A(\mem[3][2] ),
    .B(\mem[19][3] ));
 sg13g2_xor2_1 _5231_ (.B(_1999_),
    .A(_1998_),
    .X(_2000_));
 sg13g2_or3_1 _5232_ (.A(_1989_),
    .B(_1991_),
    .C(_2000_),
    .X(_2001_));
 sg13g2_inv_1 _5233_ (.Y(_2002_),
    .A(_2001_));
 sg13g2_o21ai_1 _5234_ (.B1(_2000_),
    .Y(_2003_),
    .A1(_1989_),
    .A2(_1991_));
 sg13g2_nand2_1 _5235_ (.Y(_2004_),
    .A(_2001_),
    .B(_2003_));
 sg13g2_nand2_1 _5236_ (.Y(_2005_),
    .A(_1994_),
    .B(_1996_));
 sg13g2_xor2_1 _5237_ (.B(_2005_),
    .A(_2004_),
    .X(_2006_));
 sg13g2_nor2_1 _5238_ (.A(_1956_),
    .B(_2006_),
    .Y(_0375_));
 sg13g2_a21oi_1 _5239_ (.A1(_1964_),
    .A2(_1999_),
    .Y(_2007_),
    .B1(_1987_));
 sg13g2_nand2_1 _5240_ (.Y(_2008_),
    .A(net755),
    .B(\mem[19][3] ));
 sg13g2_nand2b_1 _5241_ (.Y(_2009_),
    .B(_2007_),
    .A_N(_2008_));
 sg13g2_xnor2_1 _5242_ (.Y(_2010_),
    .A(_2007_),
    .B(_2008_));
 sg13g2_o21ai_1 _5243_ (.B1(_2003_),
    .Y(_2011_),
    .A1(_1994_),
    .A2(_2002_));
 sg13g2_nand2_1 _5244_ (.Y(_2012_),
    .A(_2010_),
    .B(_2011_));
 sg13g2_o21ai_1 _5245_ (.B1(_1957_),
    .Y(_2013_),
    .A1(_2010_),
    .A2(_2011_));
 sg13g2_nor2b_1 _5246_ (.A(_2013_),
    .B_N(_2012_),
    .Y(_0376_));
 sg13g2_a21oi_1 _5247_ (.A1(_2009_),
    .A2(_2012_),
    .Y(_0377_),
    .B1(_1956_));
 sg13g2_nor2_2 _5248_ (.A(_1547_),
    .B(_1666_),
    .Y(_2014_));
 sg13g2_inv_1 _5249_ (.Y(_2015_),
    .A(_2014_));
 sg13g2_and3_1 _5250_ (.X(_0378_),
    .A(net684),
    .B(\mem[18][0] ),
    .C(_2015_));
 sg13g2_a22oi_1 _5251_ (.Y(_2016_),
    .B1(net722),
    .B2(net684),
    .A2(\mem[2][1] ),
    .A1(\mem[18][0] ));
 sg13g2_nand4_1 _5252_ (.B(\mem[18][0] ),
    .C(net749),
    .A(net684),
    .Y(_2017_),
    .D(\mem[18][1] ));
 sg13g2_inv_1 _5253_ (.Y(_2018_),
    .A(_2017_));
 sg13g2_nor3_1 _5254_ (.A(_2014_),
    .B(net723),
    .C(_2018_),
    .Y(_0379_));
 sg13g2_a22oi_1 _5255_ (.Y(_2019_),
    .B1(\mem[18][2] ),
    .B2(\mem[2][0] ),
    .A2(\mem[18][1] ),
    .A1(\mem[2][1] ));
 sg13g2_nand2_1 _5256_ (.Y(_2020_),
    .A(\mem[2][1] ),
    .B(\mem[18][2] ));
 sg13g2_and4_1 _5257_ (.A(\mem[2][0] ),
    .B(\mem[2][1] ),
    .C(\mem[18][1] ),
    .D(\mem[18][2] ),
    .X(_2021_));
 sg13g2_nor2_1 _5258_ (.A(_2019_),
    .B(_2021_),
    .Y(_2022_));
 sg13g2_nand2_1 _5259_ (.Y(_2023_),
    .A(\mem[18][0] ),
    .B(\mem[2][2] ));
 sg13g2_nor3_1 _5260_ (.A(_2019_),
    .B(_2021_),
    .C(_2023_),
    .Y(_2024_));
 sg13g2_xor2_1 _5261_ (.B(_2023_),
    .A(_2022_),
    .X(_2025_));
 sg13g2_and2_1 _5262_ (.A(_2017_),
    .B(_2025_),
    .X(_2026_));
 sg13g2_nor2_1 _5263_ (.A(_2017_),
    .B(_2025_),
    .Y(_2027_));
 sg13g2_nor3_1 _5264_ (.A(_2014_),
    .B(_2026_),
    .C(_2027_),
    .Y(_0380_));
 sg13g2_nand2_1 _5265_ (.Y(_2028_),
    .A(\mem[18][0] ),
    .B(\mem[2][3] ));
 sg13g2_nand2_1 _5266_ (.Y(_2029_),
    .A(\mem[18][1] ),
    .B(\mem[2][2] ));
 sg13g2_nand2_1 _5267_ (.Y(_2030_),
    .A(\mem[2][1] ),
    .B(\mem[18][3] ));
 sg13g2_nand2_1 _5268_ (.Y(_2031_),
    .A(\mem[2][0] ),
    .B(\mem[18][3] ));
 sg13g2_xor2_1 _5269_ (.B(_2031_),
    .A(_2020_),
    .X(_2032_));
 sg13g2_nand2b_1 _5270_ (.Y(_2033_),
    .B(_2032_),
    .A_N(_2029_));
 sg13g2_xnor2_1 _5271_ (.Y(_2034_),
    .A(_2029_),
    .B(_2032_));
 sg13g2_nand2_1 _5272_ (.Y(_2035_),
    .A(_2021_),
    .B(_2034_));
 sg13g2_xor2_1 _5273_ (.B(_2034_),
    .A(_2021_),
    .X(_2036_));
 sg13g2_nand2b_1 _5274_ (.Y(_2037_),
    .B(_2036_),
    .A_N(_2028_));
 sg13g2_xnor2_1 _5275_ (.Y(_2038_),
    .A(_2028_),
    .B(_2036_));
 sg13g2_and2_1 _5276_ (.A(_2024_),
    .B(_2038_),
    .X(_2039_));
 sg13g2_xor2_1 _5277_ (.B(_2038_),
    .A(_2024_),
    .X(_2040_));
 sg13g2_o21ai_1 _5278_ (.B1(_2015_),
    .Y(_2041_),
    .A1(_2027_),
    .A2(_2040_));
 sg13g2_a21oi_1 _5279_ (.A1(_2027_),
    .A2(_2040_),
    .Y(_0381_),
    .B1(_2041_));
 sg13g2_a21oi_1 _5280_ (.A1(_2027_),
    .A2(_2040_),
    .Y(_2042_),
    .B1(_2039_));
 sg13g2_o21ai_1 _5281_ (.B1(_2033_),
    .Y(_2043_),
    .A1(_2020_),
    .A2(_2031_));
 sg13g2_nand2_1 _5282_ (.Y(_2044_),
    .A(\mem[18][1] ),
    .B(\mem[2][3] ));
 sg13g2_nand2_1 _5283_ (.Y(_2045_),
    .A(\mem[2][2] ),
    .B(\mem[18][3] ));
 sg13g2_nand2_2 _5284_ (.Y(_2046_),
    .A(net767),
    .B(\mem[18][2] ));
 sg13g2_xor2_1 _5285_ (.B(_2046_),
    .A(_2030_),
    .X(_2047_));
 sg13g2_nand2b_1 _5286_ (.Y(_2048_),
    .B(_2047_),
    .A_N(_2044_));
 sg13g2_xnor2_1 _5287_ (.Y(_2049_),
    .A(_2044_),
    .B(_2047_));
 sg13g2_nand2_1 _5288_ (.Y(_2050_),
    .A(_2043_),
    .B(_2049_));
 sg13g2_xnor2_1 _5289_ (.Y(_2051_),
    .A(_2043_),
    .B(_2049_));
 sg13g2_a21o_1 _5290_ (.A2(_2037_),
    .A1(_2035_),
    .B1(_2051_),
    .X(_2052_));
 sg13g2_nand3_1 _5291_ (.B(_2037_),
    .C(_2051_),
    .A(_2035_),
    .Y(_2053_));
 sg13g2_nand2_1 _5292_ (.Y(_2054_),
    .A(_2052_),
    .B(_2053_));
 sg13g2_or2_1 _5293_ (.X(_2055_),
    .B(_2054_),
    .A(_2042_));
 sg13g2_nand2_1 _5294_ (.Y(_2056_),
    .A(_2015_),
    .B(_2055_));
 sg13g2_a21oi_1 _5295_ (.A1(_2042_),
    .A2(_2054_),
    .Y(_0382_),
    .B1(_2056_));
 sg13g2_nand2_1 _5296_ (.Y(_2057_),
    .A(_2052_),
    .B(_2055_));
 sg13g2_o21ai_1 _5297_ (.B1(_2048_),
    .Y(_2058_),
    .A1(_2030_),
    .A2(_2046_));
 sg13g2_nand2_1 _5298_ (.Y(_2059_),
    .A(\mem[18][2] ),
    .B(\mem[2][3] ));
 sg13g2_nand2_1 _5299_ (.Y(_2060_),
    .A(net724),
    .B(net786));
 sg13g2_xor2_1 _5300_ (.B(_2059_),
    .A(_2045_),
    .X(_2061_));
 sg13g2_nand2_1 _5301_ (.Y(_2062_),
    .A(_2058_),
    .B(_2061_));
 sg13g2_xnor2_1 _5302_ (.Y(_2063_),
    .A(_2058_),
    .B(_2061_));
 sg13g2_xor2_1 _5303_ (.B(_2063_),
    .A(_2050_),
    .X(_2064_));
 sg13g2_xnor2_1 _5304_ (.Y(_2065_),
    .A(_2057_),
    .B(_2064_));
 sg13g2_nor2_1 _5305_ (.A(_2014_),
    .B(_2065_),
    .Y(_0383_));
 sg13g2_nand2b_1 _5306_ (.Y(_2066_),
    .B(_2046_),
    .A_N(_2060_));
 sg13g2_xor2_1 _5307_ (.B(_2066_),
    .A(_2062_),
    .X(_2067_));
 sg13g2_and2_1 _5308_ (.A(_2050_),
    .B(_2052_),
    .X(_2068_));
 sg13g2_a21oi_1 _5309_ (.A1(_2042_),
    .A2(_2068_),
    .Y(_2069_),
    .B1(_2063_));
 sg13g2_o21ai_1 _5310_ (.B1(_2015_),
    .Y(_2070_),
    .A1(_2067_),
    .A2(_2069_));
 sg13g2_a21oi_1 _5311_ (.A1(_2067_),
    .A2(_2069_),
    .Y(_0384_),
    .B1(_2070_));
 sg13g2_a21oi_1 _5312_ (.A1(_2046_),
    .A2(_2062_),
    .Y(_2071_),
    .B1(_2060_));
 sg13g2_a21oi_1 _5313_ (.A1(_2067_),
    .A2(_2069_),
    .Y(_2072_),
    .B1(_2071_));
 sg13g2_nor2_1 _5314_ (.A(_2014_),
    .B(_2072_),
    .Y(_0385_));
 sg13g2_o21ai_1 _5315_ (.B1(net578),
    .Y(_2073_),
    .A1(uio_out[5]),
    .A2(net733));
 sg13g2_inv_1 _5316_ (.Y(_0386_),
    .A(net734));
 sg13g2_nand2_1 _5317_ (.Y(_2074_),
    .A(net678),
    .B(net579));
 sg13g2_a22oi_1 _5318_ (.Y(_0387_),
    .B1(net484),
    .B2(_2074_),
    .A2(net489),
    .A1(_2089_));
 sg13g2_nand2_1 _5319_ (.Y(_2075_),
    .A(net682),
    .B(net579));
 sg13g2_a22oi_1 _5320_ (.Y(_0388_),
    .B1(net484),
    .B2(_2075_),
    .A2(net489),
    .A1(_2088_));
 sg13g2_nand2_1 _5321_ (.Y(_2076_),
    .A(\prev_acc[2] ),
    .B(net579));
 sg13g2_a22oi_1 _5322_ (.Y(_0389_),
    .B1(net484),
    .B2(_2076_),
    .A2(net489),
    .A1(_2087_));
 sg13g2_nand2_1 _5323_ (.Y(_2077_),
    .A(\prev_acc[3] ),
    .B(net578));
 sg13g2_a22oi_1 _5324_ (.Y(_0390_),
    .B1(net484),
    .B2(_2077_),
    .A2(net489),
    .A1(_2086_));
 sg13g2_nand2_1 _5325_ (.Y(_2078_),
    .A(net709),
    .B(net580));
 sg13g2_a22oi_1 _5326_ (.Y(_0391_),
    .B1(net484),
    .B2(_2078_),
    .A2(net489),
    .A1(_2085_));
 sg13g2_nand2_1 _5327_ (.Y(_2079_),
    .A(net715),
    .B(net578));
 sg13g2_a22oi_1 _5328_ (.Y(_0392_),
    .B1(net484),
    .B2(_2079_),
    .A2(net489),
    .A1(_2084_));
 sg13g2_nand2_1 _5329_ (.Y(_2080_),
    .A(net686),
    .B(net580));
 sg13g2_a22oi_1 _5330_ (.Y(_0393_),
    .B1(net485),
    .B2(_2080_),
    .A2(net489),
    .A1(_2083_));
 sg13g2_nand2_1 _5331_ (.Y(_2081_),
    .A(net695),
    .B(net580));
 sg13g2_a22oi_1 _5332_ (.Y(_0394_),
    .B1(net484),
    .B2(_2081_),
    .A2(_0780_),
    .A1(_2082_));
 sg13g2_dfrbp_1 _5333_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net173),
    .D(_0001_),
    .Q_N(_2663_),
    .Q(\mem[13][0] ));
 sg13g2_dfrbp_1 _5334_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net167),
    .D(_0002_),
    .Q_N(_2662_),
    .Q(\mem[13][1] ));
 sg13g2_dfrbp_1 _5335_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net166),
    .D(_0003_),
    .Q_N(_2661_),
    .Q(\mem[13][2] ));
 sg13g2_dfrbp_1 _5336_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net165),
    .D(_0004_),
    .Q_N(_2660_),
    .Q(\mem[13][3] ));
 sg13g2_dfrbp_1 _5337_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net164),
    .D(_0005_),
    .Q_N(_2659_),
    .Q(\mem[19][0] ));
 sg13g2_dfrbp_1 _5338_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net163),
    .D(_0006_),
    .Q_N(_2658_),
    .Q(\mem[19][1] ));
 sg13g2_dfrbp_1 _5339_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net162),
    .D(_0007_),
    .Q_N(_2657_),
    .Q(\mem[19][2] ));
 sg13g2_dfrbp_1 _5340_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net161),
    .D(_0008_),
    .Q_N(_2656_),
    .Q(\mem[19][3] ));
 sg13g2_dfrbp_1 _5341_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net160),
    .D(_0009_),
    .Q_N(_2655_),
    .Q(\mem[11][0] ));
 sg13g2_dfrbp_1 _5342_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net159),
    .D(_0010_),
    .Q_N(_2654_),
    .Q(\mem[11][1] ));
 sg13g2_dfrbp_1 _5343_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net158),
    .D(_0011_),
    .Q_N(_2653_),
    .Q(\mem[11][2] ));
 sg13g2_dfrbp_1 _5344_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net157),
    .D(_0012_),
    .Q_N(_2652_),
    .Q(\mem[11][3] ));
 sg13g2_dfrbp_1 _5345_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net156),
    .D(_0013_),
    .Q_N(_2651_),
    .Q(\mem[29][0] ));
 sg13g2_dfrbp_1 _5346_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net155),
    .D(_0014_),
    .Q_N(_2650_),
    .Q(\mem[29][1] ));
 sg13g2_dfrbp_1 _5347_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net154),
    .D(_0015_),
    .Q_N(_2649_),
    .Q(\mem[29][2] ));
 sg13g2_dfrbp_1 _5348_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net153),
    .D(_0016_),
    .Q_N(_2648_),
    .Q(\mem[29][3] ));
 sg13g2_dfrbp_1 _5349_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net152),
    .D(_0017_),
    .Q_N(_2647_),
    .Q(\mem[10][0] ));
 sg13g2_dfrbp_1 _5350_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net151),
    .D(_0018_),
    .Q_N(_2646_),
    .Q(\mem[10][1] ));
 sg13g2_dfrbp_1 _5351_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net150),
    .D(_0019_),
    .Q_N(_2645_),
    .Q(\mem[10][2] ));
 sg13g2_dfrbp_1 _5352_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net149),
    .D(_0020_),
    .Q_N(_2644_),
    .Q(\mem[10][3] ));
 sg13g2_dfrbp_1 _5353_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net148),
    .D(_0021_),
    .Q_N(_2643_),
    .Q(\mem[49][0] ));
 sg13g2_dfrbp_1 _5354_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net147),
    .D(_0022_),
    .Q_N(_2642_),
    .Q(\mem[49][1] ));
 sg13g2_dfrbp_1 _5355_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net146),
    .D(_0023_),
    .Q_N(_2641_),
    .Q(\mem[49][2] ));
 sg13g2_dfrbp_1 _5356_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net145),
    .D(_0024_),
    .Q_N(_2640_),
    .Q(\mem[49][3] ));
 sg13g2_dfrbp_1 _5357_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net144),
    .D(_0025_),
    .Q_N(_2639_),
    .Q(\mem[59][0] ));
 sg13g2_dfrbp_1 _5358_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net143),
    .D(_0026_),
    .Q_N(_2638_),
    .Q(\mem[59][1] ));
 sg13g2_dfrbp_1 _5359_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net142),
    .D(_0027_),
    .Q_N(_2637_),
    .Q(\mem[59][2] ));
 sg13g2_dfrbp_1 _5360_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net141),
    .D(_0028_),
    .Q_N(_2636_),
    .Q(\mem[59][3] ));
 sg13g2_dfrbp_1 _5361_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net140),
    .D(_0029_),
    .Q_N(_2635_),
    .Q(\products[0][0] ));
 sg13g2_dfrbp_1 _5362_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net139),
    .D(_0030_),
    .Q_N(_2634_),
    .Q(\products[0][1] ));
 sg13g2_dfrbp_1 _5363_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net138),
    .D(_0031_),
    .Q_N(_2633_),
    .Q(\products[0][2] ));
 sg13g2_dfrbp_1 _5364_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net137),
    .D(_0032_),
    .Q_N(_2632_),
    .Q(\products[0][3] ));
 sg13g2_dfrbp_1 _5365_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net136),
    .D(_0033_),
    .Q_N(_2631_),
    .Q(\products[0][4] ));
 sg13g2_dfrbp_1 _5366_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net135),
    .D(_0034_),
    .Q_N(_2630_),
    .Q(\products[0][5] ));
 sg13g2_dfrbp_1 _5367_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net134),
    .D(_0035_),
    .Q_N(_2629_),
    .Q(\products[0][6] ));
 sg13g2_dfrbp_1 _5368_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net133),
    .D(_0036_),
    .Q_N(_2628_),
    .Q(\products[0][7] ));
 sg13g2_dfrbp_1 _5369_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net132),
    .D(_0037_),
    .Q_N(_2627_),
    .Q(\mem[63][0] ));
 sg13g2_dfrbp_1 _5370_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net131),
    .D(_0038_),
    .Q_N(_2626_),
    .Q(\mem[63][1] ));
 sg13g2_dfrbp_1 _5371_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net130),
    .D(_0039_),
    .Q_N(_2625_),
    .Q(\mem[63][2] ));
 sg13g2_dfrbp_1 _5372_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net129),
    .D(_0040_),
    .Q_N(_2624_),
    .Q(\mem[63][3] ));
 sg13g2_dfrbp_1 _5373_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net128),
    .D(_0041_),
    .Q_N(_2623_),
    .Q(\mem[6][0] ));
 sg13g2_dfrbp_1 _5374_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net127),
    .D(_0042_),
    .Q_N(_2622_),
    .Q(\mem[6][1] ));
 sg13g2_dfrbp_1 _5375_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net126),
    .D(_0043_),
    .Q_N(_2621_),
    .Q(\mem[6][2] ));
 sg13g2_dfrbp_1 _5376_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net125),
    .D(_0044_),
    .Q_N(_2620_),
    .Q(\mem[6][3] ));
 sg13g2_dfrbp_1 _5377_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net124),
    .D(_0045_),
    .Q_N(_2619_),
    .Q(\mem[7][0] ));
 sg13g2_dfrbp_1 _5378_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net123),
    .D(_0046_),
    .Q_N(_2618_),
    .Q(\mem[7][1] ));
 sg13g2_dfrbp_1 _5379_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net122),
    .D(_0047_),
    .Q_N(_2617_),
    .Q(\mem[7][2] ));
 sg13g2_dfrbp_1 _5380_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net121),
    .D(_0048_),
    .Q_N(_2616_),
    .Q(\mem[7][3] ));
 sg13g2_dfrbp_1 _5381_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net120),
    .D(_0049_),
    .Q_N(_2615_),
    .Q(\mem[2][0] ));
 sg13g2_dfrbp_1 _5382_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net119),
    .D(_0050_),
    .Q_N(_2614_),
    .Q(\mem[2][1] ));
 sg13g2_dfrbp_1 _5383_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net118),
    .D(_0051_),
    .Q_N(_2613_),
    .Q(\mem[2][2] ));
 sg13g2_dfrbp_1 _5384_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net117),
    .D(_0052_),
    .Q_N(_2612_),
    .Q(\mem[2][3] ));
 sg13g2_dfrbp_1 _5385_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net116),
    .D(_0053_),
    .Q_N(_2611_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _5386_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net115),
    .D(net704),
    .Q_N(_2610_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _5387_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net114),
    .D(_0055_),
    .Q_N(_2609_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _5388_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net113),
    .D(net773),
    .Q_N(_2608_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _5389_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net112),
    .D(_0057_),
    .Q_N(_2607_),
    .Q(\mem[25][0] ));
 sg13g2_dfrbp_1 _5390_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net111),
    .D(_0058_),
    .Q_N(_2606_),
    .Q(\mem[25][1] ));
 sg13g2_dfrbp_1 _5391_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net110),
    .D(_0059_),
    .Q_N(_2605_),
    .Q(\mem[25][2] ));
 sg13g2_dfrbp_1 _5392_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net109),
    .D(_0060_),
    .Q_N(_2604_),
    .Q(\mem[25][3] ));
 sg13g2_dfrbp_1 _5393_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net108),
    .D(_0061_),
    .Q_N(_2603_),
    .Q(\mem[20][0] ));
 sg13g2_dfrbp_1 _5394_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net107),
    .D(_0062_),
    .Q_N(_2602_),
    .Q(\mem[20][1] ));
 sg13g2_dfrbp_1 _5395_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net106),
    .D(_0063_),
    .Q_N(_2601_),
    .Q(\mem[20][2] ));
 sg13g2_dfrbp_1 _5396_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net105),
    .D(_0064_),
    .Q_N(_2600_),
    .Q(\mem[20][3] ));
 sg13g2_dfrbp_1 _5397_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net104),
    .D(_0065_),
    .Q_N(_2599_),
    .Q(\mem[30][0] ));
 sg13g2_dfrbp_1 _5398_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net103),
    .D(_0066_),
    .Q_N(_2598_),
    .Q(\mem[30][1] ));
 sg13g2_dfrbp_1 _5399_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net102),
    .D(_0067_),
    .Q_N(_2597_),
    .Q(\mem[30][2] ));
 sg13g2_dfrbp_1 _5400_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net101),
    .D(_0068_),
    .Q_N(_2596_),
    .Q(\mem[30][3] ));
 sg13g2_dfrbp_1 _5401_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net100),
    .D(_0069_),
    .Q_N(_2595_),
    .Q(\mem[35][0] ));
 sg13g2_dfrbp_1 _5402_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net99),
    .D(_0070_),
    .Q_N(_2594_),
    .Q(\mem[35][1] ));
 sg13g2_dfrbp_1 _5403_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net98),
    .D(_0071_),
    .Q_N(_2593_),
    .Q(\mem[35][2] ));
 sg13g2_dfrbp_1 _5404_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net97),
    .D(_0072_),
    .Q_N(_2592_),
    .Q(\mem[35][3] ));
 sg13g2_dfrbp_1 _5405_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net96),
    .D(_0073_),
    .Q_N(_2591_),
    .Q(\mem[26][0] ));
 sg13g2_dfrbp_1 _5406_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net95),
    .D(_0074_),
    .Q_N(_2590_),
    .Q(\mem[26][1] ));
 sg13g2_dfrbp_1 _5407_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net94),
    .D(_0075_),
    .Q_N(_2589_),
    .Q(\mem[26][2] ));
 sg13g2_dfrbp_1 _5408_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net93),
    .D(_0076_),
    .Q_N(_2588_),
    .Q(\mem[26][3] ));
 sg13g2_dfrbp_1 _5409_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net92),
    .D(_0077_),
    .Q_N(_2587_),
    .Q(\mem[21][0] ));
 sg13g2_dfrbp_1 _5410_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net91),
    .D(_0078_),
    .Q_N(_2586_),
    .Q(\mem[21][1] ));
 sg13g2_dfrbp_1 _5411_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net90),
    .D(_0079_),
    .Q_N(_2585_),
    .Q(\mem[21][2] ));
 sg13g2_dfrbp_1 _5412_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net89),
    .D(_0080_),
    .Q_N(_2584_),
    .Q(\mem[21][3] ));
 sg13g2_dfrbp_1 _5413_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net88),
    .D(_0081_),
    .Q_N(_2583_),
    .Q(\mem[39][0] ));
 sg13g2_dfrbp_1 _5414_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net87),
    .D(_0082_),
    .Q_N(_2582_),
    .Q(\mem[39][1] ));
 sg13g2_dfrbp_1 _5415_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net86),
    .D(_0083_),
    .Q_N(_2581_),
    .Q(\mem[39][2] ));
 sg13g2_dfrbp_1 _5416_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net85),
    .D(_0084_),
    .Q_N(_2580_),
    .Q(\mem[39][3] ));
 sg13g2_dfrbp_1 _5417_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net84),
    .D(_0085_),
    .Q_N(_2579_),
    .Q(\mem[31][0] ));
 sg13g2_dfrbp_1 _5418_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net83),
    .D(_0086_),
    .Q_N(_2578_),
    .Q(\mem[31][1] ));
 sg13g2_dfrbp_1 _5419_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net82),
    .D(_0087_),
    .Q_N(_2577_),
    .Q(\mem[31][2] ));
 sg13g2_dfrbp_1 _5420_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net81),
    .D(_0088_),
    .Q_N(_2576_),
    .Q(\mem[31][3] ));
 sg13g2_dfrbp_1 _5421_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net80),
    .D(_0089_),
    .Q_N(_2575_),
    .Q(\mem[27][0] ));
 sg13g2_dfrbp_1 _5422_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net79),
    .D(_0090_),
    .Q_N(_2574_),
    .Q(\mem[27][1] ));
 sg13g2_dfrbp_1 _5423_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net78),
    .D(_0091_),
    .Q_N(_2573_),
    .Q(\mem[27][2] ));
 sg13g2_dfrbp_1 _5424_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net77),
    .D(_0092_),
    .Q_N(_2572_),
    .Q(\mem[27][3] ));
 sg13g2_dfrbp_1 _5425_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net76),
    .D(_0093_),
    .Q_N(_2571_),
    .Q(\mem[22][0] ));
 sg13g2_dfrbp_1 _5426_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net75),
    .D(_0094_),
    .Q_N(_2570_),
    .Q(\mem[22][1] ));
 sg13g2_dfrbp_1 _5427_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net74),
    .D(_0095_),
    .Q_N(_2569_),
    .Q(\mem[22][2] ));
 sg13g2_dfrbp_1 _5428_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net73),
    .D(_0096_),
    .Q_N(_2568_),
    .Q(\mem[22][3] ));
 sg13g2_dfrbp_1 _5429_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net72),
    .D(_0097_),
    .Q_N(_2567_),
    .Q(\mem[17][0] ));
 sg13g2_dfrbp_1 _5430_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net71),
    .D(_0098_),
    .Q_N(_2566_),
    .Q(\mem[17][1] ));
 sg13g2_dfrbp_1 _5431_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net70),
    .D(_0099_),
    .Q_N(_2565_),
    .Q(\mem[17][2] ));
 sg13g2_dfrbp_1 _5432_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net69),
    .D(_0100_),
    .Q_N(_2564_),
    .Q(\mem[17][3] ));
 sg13g2_dfrbp_1 _5433_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net68),
    .D(_0101_),
    .Q_N(_2563_),
    .Q(\mem[32][0] ));
 sg13g2_dfrbp_1 _5434_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net67),
    .D(_0102_),
    .Q_N(_2562_),
    .Q(\mem[32][1] ));
 sg13g2_dfrbp_1 _5435_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net66),
    .D(_0103_),
    .Q_N(_2561_),
    .Q(\mem[32][2] ));
 sg13g2_dfrbp_1 _5436_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net65),
    .D(_0104_),
    .Q_N(_2560_),
    .Q(\mem[32][3] ));
 sg13g2_dfrbp_1 _5437_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net64),
    .D(_0105_),
    .Q_N(_2559_),
    .Q(\mem[23][0] ));
 sg13g2_dfrbp_1 _5438_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net63),
    .D(_0106_),
    .Q_N(_2558_),
    .Q(\mem[23][1] ));
 sg13g2_dfrbp_1 _5439_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net62),
    .D(_0107_),
    .Q_N(_2557_),
    .Q(\mem[23][2] ));
 sg13g2_dfrbp_1 _5440_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net61),
    .D(_0108_),
    .Q_N(_2556_),
    .Q(\mem[23][3] ));
 sg13g2_dfrbp_1 _5441_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net60),
    .D(_0109_),
    .Q_N(_2555_),
    .Q(\mem[18][0] ));
 sg13g2_dfrbp_1 _5442_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net59),
    .D(_0110_),
    .Q_N(_2554_),
    .Q(\mem[18][1] ));
 sg13g2_dfrbp_1 _5443_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net58),
    .D(_0111_),
    .Q_N(_2553_),
    .Q(\mem[18][2] ));
 sg13g2_dfrbp_1 _5444_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net57),
    .D(_0112_),
    .Q_N(_2552_),
    .Q(\mem[18][3] ));
 sg13g2_dfrbp_1 _5445_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net56),
    .D(_0113_),
    .Q_N(_2551_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _5446_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net55),
    .D(_0114_),
    .Q_N(_2550_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _5447_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net54),
    .D(_0115_),
    .Q_N(_2549_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _5448_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net53),
    .D(_0116_),
    .Q_N(_2548_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _5449_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net52),
    .D(_0117_),
    .Q_N(_2547_),
    .Q(\mem[28][0] ));
 sg13g2_dfrbp_1 _5450_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net51),
    .D(_0118_),
    .Q_N(_2546_),
    .Q(\mem[28][1] ));
 sg13g2_dfrbp_1 _5451_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net50),
    .D(_0119_),
    .Q_N(_2545_),
    .Q(\mem[28][2] ));
 sg13g2_dfrbp_1 _5452_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net49),
    .D(_0120_),
    .Q_N(_2544_),
    .Q(\mem[28][3] ));
 sg13g2_dfrbp_1 _5453_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net48),
    .D(_0121_),
    .Q_N(_2543_),
    .Q(\mem[24][0] ));
 sg13g2_dfrbp_1 _5454_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net47),
    .D(_0122_),
    .Q_N(_2542_),
    .Q(\mem[24][1] ));
 sg13g2_dfrbp_1 _5455_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net46),
    .D(_0123_),
    .Q_N(_2541_),
    .Q(\mem[24][2] ));
 sg13g2_dfrbp_1 _5456_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net45),
    .D(_0124_),
    .Q_N(_2540_),
    .Q(\mem[24][3] ));
 sg13g2_dfrbp_1 _5457_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net44),
    .D(_0125_),
    .Q_N(_2539_),
    .Q(\mem[1][0] ));
 sg13g2_dfrbp_1 _5458_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net43),
    .D(_0126_),
    .Q_N(_2538_),
    .Q(\mem[1][1] ));
 sg13g2_dfrbp_1 _5459_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net42),
    .D(_0127_),
    .Q_N(_2537_),
    .Q(\mem[1][2] ));
 sg13g2_dfrbp_1 _5460_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net41),
    .D(_0128_),
    .Q_N(_2536_),
    .Q(\mem[1][3] ));
 sg13g2_dfrbp_1 _5461_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net40),
    .D(_0129_),
    .Q_N(_2535_),
    .Q(\mem[40][0] ));
 sg13g2_dfrbp_1 _5462_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net39),
    .D(_0130_),
    .Q_N(_2534_),
    .Q(\mem[40][1] ));
 sg13g2_dfrbp_1 _5463_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net38),
    .D(_0131_),
    .Q_N(_2533_),
    .Q(\mem[40][2] ));
 sg13g2_dfrbp_1 _5464_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net37),
    .D(_0132_),
    .Q_N(_2532_),
    .Q(\mem[40][3] ));
 sg13g2_dfrbp_1 _5465_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net36),
    .D(_0133_),
    .Q_N(_2531_),
    .Q(\mem[3][0] ));
 sg13g2_dfrbp_1 _5466_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net35),
    .D(_0134_),
    .Q_N(_2530_),
    .Q(\mem[3][1] ));
 sg13g2_dfrbp_1 _5467_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net34),
    .D(_0135_),
    .Q_N(_2529_),
    .Q(\mem[3][2] ));
 sg13g2_dfrbp_1 _5468_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net33),
    .D(_0136_),
    .Q_N(_2528_),
    .Q(\mem[3][3] ));
 sg13g2_dfrbp_1 _5469_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net32),
    .D(_0137_),
    .Q_N(_2527_),
    .Q(\mem[38][0] ));
 sg13g2_dfrbp_1 _5470_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net31),
    .D(_0138_),
    .Q_N(_2526_),
    .Q(\mem[38][1] ));
 sg13g2_dfrbp_1 _5471_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net30),
    .D(_0139_),
    .Q_N(_2525_),
    .Q(\mem[38][2] ));
 sg13g2_dfrbp_1 _5472_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net29),
    .D(_0140_),
    .Q_N(_2524_),
    .Q(\mem[38][3] ));
 sg13g2_dfrbp_1 _5473_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net28),
    .D(_0141_),
    .Q_N(_2523_),
    .Q(\mem[37][0] ));
 sg13g2_dfrbp_1 _5474_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net27),
    .D(_0142_),
    .Q_N(_2522_),
    .Q(\mem[37][1] ));
 sg13g2_dfrbp_1 _5475_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net26),
    .D(_0143_),
    .Q_N(_2521_),
    .Q(\mem[37][2] ));
 sg13g2_dfrbp_1 _5476_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net25),
    .D(_0144_),
    .Q_N(_2520_),
    .Q(\mem[37][3] ));
 sg13g2_dfrbp_1 _5477_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net24),
    .D(_0145_),
    .Q_N(_2519_),
    .Q(\mem[36][0] ));
 sg13g2_dfrbp_1 _5478_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net23),
    .D(_0146_),
    .Q_N(_2518_),
    .Q(\mem[36][1] ));
 sg13g2_dfrbp_1 _5479_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net22),
    .D(_0147_),
    .Q_N(_2517_),
    .Q(\mem[36][2] ));
 sg13g2_dfrbp_1 _5480_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net21),
    .D(_0148_),
    .Q_N(_2516_),
    .Q(\mem[36][3] ));
 sg13g2_dfrbp_1 _5481_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net20),
    .D(_0149_),
    .Q_N(_2515_),
    .Q(uio_out[4]));
 sg13g2_dfrbp_1 _5482_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net18),
    .D(_0150_),
    .Q_N(_2514_),
    .Q(\mem[16][0] ));
 sg13g2_dfrbp_1 _5483_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net17),
    .D(_0151_),
    .Q_N(_2513_),
    .Q(\mem[16][1] ));
 sg13g2_dfrbp_1 _5484_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net16),
    .D(_0152_),
    .Q_N(_2512_),
    .Q(\mem[16][2] ));
 sg13g2_dfrbp_1 _5485_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net15),
    .D(_0153_),
    .Q_N(_2511_),
    .Q(\mem[16][3] ));
 sg13g2_dfrbp_1 _5486_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net14),
    .D(_0154_),
    .Q_N(_2510_),
    .Q(\mem[15][0] ));
 sg13g2_dfrbp_1 _5487_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net13),
    .D(_0155_),
    .Q_N(_2509_),
    .Q(\mem[15][1] ));
 sg13g2_dfrbp_1 _5488_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net12),
    .D(_0156_),
    .Q_N(_2508_),
    .Q(\mem[15][2] ));
 sg13g2_dfrbp_1 _5489_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net11),
    .D(_0157_),
    .Q_N(_2507_),
    .Q(\mem[15][3] ));
 sg13g2_dfrbp_1 _5490_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net404),
    .D(_0158_),
    .Q_N(_2506_),
    .Q(\mem[14][0] ));
 sg13g2_dfrbp_1 _5491_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net403),
    .D(_0159_),
    .Q_N(_2505_),
    .Q(\mem[14][1] ));
 sg13g2_dfrbp_1 _5492_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net402),
    .D(_0160_),
    .Q_N(_2504_),
    .Q(\mem[14][2] ));
 sg13g2_dfrbp_1 _5493_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net401),
    .D(_0161_),
    .Q_N(_2503_),
    .Q(\mem[14][3] ));
 sg13g2_dfrbp_1 _5494_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net400),
    .D(_0162_),
    .Q_N(_2502_),
    .Q(\mem[62][0] ));
 sg13g2_dfrbp_1 _5495_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net399),
    .D(_0163_),
    .Q_N(_2501_),
    .Q(\mem[62][1] ));
 sg13g2_dfrbp_1 _5496_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net398),
    .D(_0164_),
    .Q_N(_2500_),
    .Q(\mem[62][2] ));
 sg13g2_dfrbp_1 _5497_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net397),
    .D(_0165_),
    .Q_N(_2499_),
    .Q(\mem[62][3] ));
 sg13g2_dfrbp_1 _5498_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net396),
    .D(_0166_),
    .Q_N(_2498_),
    .Q(\mem[61][0] ));
 sg13g2_dfrbp_1 _5499_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net395),
    .D(_0167_),
    .Q_N(_2497_),
    .Q(\mem[61][1] ));
 sg13g2_dfrbp_1 _5500_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net394),
    .D(_0168_),
    .Q_N(_2496_),
    .Q(\mem[61][2] ));
 sg13g2_dfrbp_1 _5501_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net393),
    .D(_0169_),
    .Q_N(_2495_),
    .Q(\mem[61][3] ));
 sg13g2_dfrbp_1 _5502_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net392),
    .D(_0170_),
    .Q_N(_2494_),
    .Q(\mem[60][0] ));
 sg13g2_dfrbp_1 _5503_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net391),
    .D(_0171_),
    .Q_N(_2493_),
    .Q(\mem[60][1] ));
 sg13g2_dfrbp_1 _5504_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net390),
    .D(_0172_),
    .Q_N(_2492_),
    .Q(\mem[60][2] ));
 sg13g2_dfrbp_1 _5505_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net389),
    .D(_0173_),
    .Q_N(_2491_),
    .Q(\mem[60][3] ));
 sg13g2_dfrbp_1 _5506_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net388),
    .D(_0174_),
    .Q_N(_2490_),
    .Q(\mem[5][0] ));
 sg13g2_dfrbp_1 _5507_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net387),
    .D(_0175_),
    .Q_N(_2489_),
    .Q(\mem[5][1] ));
 sg13g2_dfrbp_1 _5508_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net386),
    .D(_0176_),
    .Q_N(_2488_),
    .Q(\mem[5][2] ));
 sg13g2_dfrbp_1 _5509_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net385),
    .D(_0177_),
    .Q_N(_2487_),
    .Q(\mem[5][3] ));
 sg13g2_dfrbp_1 _5510_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net384),
    .D(_0178_),
    .Q_N(_2486_),
    .Q(\mem[58][0] ));
 sg13g2_dfrbp_1 _5511_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net383),
    .D(_0179_),
    .Q_N(_2485_),
    .Q(\mem[58][1] ));
 sg13g2_dfrbp_1 _5512_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net382),
    .D(_0180_),
    .Q_N(_2484_),
    .Q(\mem[58][2] ));
 sg13g2_dfrbp_1 _5513_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net381),
    .D(_0181_),
    .Q_N(_2483_),
    .Q(\mem[58][3] ));
 sg13g2_dfrbp_1 _5514_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net380),
    .D(_0182_),
    .Q_N(_2482_),
    .Q(\mem[57][0] ));
 sg13g2_dfrbp_1 _5515_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net379),
    .D(_0183_),
    .Q_N(_2481_),
    .Q(\mem[57][1] ));
 sg13g2_dfrbp_1 _5516_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net378),
    .D(_0184_),
    .Q_N(_2480_),
    .Q(\mem[57][2] ));
 sg13g2_dfrbp_1 _5517_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net377),
    .D(_0185_),
    .Q_N(_2479_),
    .Q(\mem[57][3] ));
 sg13g2_dfrbp_1 _5518_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net376),
    .D(_0186_),
    .Q_N(_2478_),
    .Q(\mem[56][0] ));
 sg13g2_dfrbp_1 _5519_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net375),
    .D(_0187_),
    .Q_N(_2477_),
    .Q(\mem[56][1] ));
 sg13g2_dfrbp_1 _5520_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net374),
    .D(_0188_),
    .Q_N(_2476_),
    .Q(\mem[56][2] ));
 sg13g2_dfrbp_1 _5521_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net373),
    .D(_0189_),
    .Q_N(_2475_),
    .Q(\mem[56][3] ));
 sg13g2_dfrbp_1 _5522_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net372),
    .D(_0190_),
    .Q_N(_2474_),
    .Q(\mem[55][0] ));
 sg13g2_dfrbp_1 _5523_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net371),
    .D(_0191_),
    .Q_N(_2473_),
    .Q(\mem[55][1] ));
 sg13g2_dfrbp_1 _5524_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net370),
    .D(_0192_),
    .Q_N(_2472_),
    .Q(\mem[55][2] ));
 sg13g2_dfrbp_1 _5525_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net369),
    .D(_0193_),
    .Q_N(_2471_),
    .Q(\mem[55][3] ));
 sg13g2_dfrbp_1 _5526_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net368),
    .D(_0194_),
    .Q_N(_2470_),
    .Q(\mem[54][0] ));
 sg13g2_dfrbp_1 _5527_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net367),
    .D(_0195_),
    .Q_N(_2469_),
    .Q(\mem[54][1] ));
 sg13g2_dfrbp_1 _5528_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net366),
    .D(_0196_),
    .Q_N(_2468_),
    .Q(\mem[54][2] ));
 sg13g2_dfrbp_1 _5529_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net365),
    .D(_0197_),
    .Q_N(_2467_),
    .Q(\mem[54][3] ));
 sg13g2_dfrbp_1 _5530_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net364),
    .D(_0198_),
    .Q_N(_2466_),
    .Q(\mem[53][0] ));
 sg13g2_dfrbp_1 _5531_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net363),
    .D(_0199_),
    .Q_N(_2465_),
    .Q(\mem[53][1] ));
 sg13g2_dfrbp_1 _5532_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net362),
    .D(_0200_),
    .Q_N(_2464_),
    .Q(\mem[53][2] ));
 sg13g2_dfrbp_1 _5533_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net361),
    .D(_0201_),
    .Q_N(_2463_),
    .Q(\mem[53][3] ));
 sg13g2_dfrbp_1 _5534_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net360),
    .D(_0202_),
    .Q_N(_2462_),
    .Q(\mem[52][0] ));
 sg13g2_dfrbp_1 _5535_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net359),
    .D(_0203_),
    .Q_N(_2461_),
    .Q(\mem[52][1] ));
 sg13g2_dfrbp_1 _5536_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net358),
    .D(_0204_),
    .Q_N(_2460_),
    .Q(\mem[52][2] ));
 sg13g2_dfrbp_1 _5537_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net357),
    .D(_0205_),
    .Q_N(_2459_),
    .Q(\mem[52][3] ));
 sg13g2_dfrbp_1 _5538_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net356),
    .D(_0206_),
    .Q_N(_2458_),
    .Q(\mem[51][0] ));
 sg13g2_dfrbp_1 _5539_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net355),
    .D(_0207_),
    .Q_N(_2457_),
    .Q(\mem[51][1] ));
 sg13g2_dfrbp_1 _5540_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net354),
    .D(_0208_),
    .Q_N(_2456_),
    .Q(\mem[51][2] ));
 sg13g2_dfrbp_1 _5541_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net353),
    .D(_0209_),
    .Q_N(_2455_),
    .Q(\mem[51][3] ));
 sg13g2_dfrbp_1 _5542_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net352),
    .D(_0210_),
    .Q_N(_2454_),
    .Q(\mem[50][0] ));
 sg13g2_dfrbp_1 _5543_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net351),
    .D(_0211_),
    .Q_N(_2453_),
    .Q(\mem[50][1] ));
 sg13g2_dfrbp_1 _5544_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net350),
    .D(_0212_),
    .Q_N(_2452_),
    .Q(\mem[50][2] ));
 sg13g2_dfrbp_1 _5545_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net349),
    .D(_0213_),
    .Q_N(_2451_),
    .Q(\mem[50][3] ));
 sg13g2_dfrbp_1 _5546_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net348),
    .D(_0214_),
    .Q_N(_2450_),
    .Q(\mem[4][0] ));
 sg13g2_dfrbp_1 _5547_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net347),
    .D(_0215_),
    .Q_N(_2449_),
    .Q(\mem[4][1] ));
 sg13g2_dfrbp_1 _5548_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net346),
    .D(_0216_),
    .Q_N(_2448_),
    .Q(\mem[4][2] ));
 sg13g2_dfrbp_1 _5549_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net345),
    .D(_0217_),
    .Q_N(_2447_),
    .Q(\mem[4][3] ));
 sg13g2_dfrbp_1 _5550_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net344),
    .D(_0218_),
    .Q_N(_2446_),
    .Q(\mem[48][0] ));
 sg13g2_dfrbp_1 _5551_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net343),
    .D(_0219_),
    .Q_N(_2445_),
    .Q(\mem[48][1] ));
 sg13g2_dfrbp_1 _5552_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net342),
    .D(_0220_),
    .Q_N(_2444_),
    .Q(\mem[48][2] ));
 sg13g2_dfrbp_1 _5553_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net341),
    .D(_0221_),
    .Q_N(_2443_),
    .Q(\mem[48][3] ));
 sg13g2_dfrbp_1 _5554_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net340),
    .D(_0222_),
    .Q_N(_2442_),
    .Q(\mem[47][0] ));
 sg13g2_dfrbp_1 _5555_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net339),
    .D(_0223_),
    .Q_N(_2441_),
    .Q(\mem[47][1] ));
 sg13g2_dfrbp_1 _5556_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net338),
    .D(_0224_),
    .Q_N(_2440_),
    .Q(\mem[47][2] ));
 sg13g2_dfrbp_1 _5557_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net337),
    .D(_0225_),
    .Q_N(_2439_),
    .Q(\mem[47][3] ));
 sg13g2_dfrbp_1 _5558_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net336),
    .D(_0226_),
    .Q_N(_2438_),
    .Q(\mem[46][0] ));
 sg13g2_dfrbp_1 _5559_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net335),
    .D(_0227_),
    .Q_N(_2437_),
    .Q(\mem[46][1] ));
 sg13g2_dfrbp_1 _5560_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net334),
    .D(_0228_),
    .Q_N(_2436_),
    .Q(\mem[46][2] ));
 sg13g2_dfrbp_1 _5561_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net333),
    .D(_0229_),
    .Q_N(_2435_),
    .Q(\mem[46][3] ));
 sg13g2_dfrbp_1 _5562_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net332),
    .D(_0230_),
    .Q_N(_2434_),
    .Q(\mem[45][0] ));
 sg13g2_dfrbp_1 _5563_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net331),
    .D(_0231_),
    .Q_N(_2433_),
    .Q(\mem[45][1] ));
 sg13g2_dfrbp_1 _5564_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net330),
    .D(_0232_),
    .Q_N(_2432_),
    .Q(\mem[45][2] ));
 sg13g2_dfrbp_1 _5565_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net329),
    .D(_0233_),
    .Q_N(_2431_),
    .Q(\mem[45][3] ));
 sg13g2_dfrbp_1 _5566_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net328),
    .D(_0234_),
    .Q_N(_2430_),
    .Q(\mem[44][0] ));
 sg13g2_dfrbp_1 _5567_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net327),
    .D(_0235_),
    .Q_N(_2429_),
    .Q(\mem[44][1] ));
 sg13g2_dfrbp_1 _5568_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net326),
    .D(_0236_),
    .Q_N(_2428_),
    .Q(\mem[44][2] ));
 sg13g2_dfrbp_1 _5569_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net325),
    .D(_0237_),
    .Q_N(_2427_),
    .Q(\mem[44][3] ));
 sg13g2_dfrbp_1 _5570_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net324),
    .D(_0238_),
    .Q_N(_2426_),
    .Q(\mem[43][0] ));
 sg13g2_dfrbp_1 _5571_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net323),
    .D(_0239_),
    .Q_N(_2425_),
    .Q(\mem[43][1] ));
 sg13g2_dfrbp_1 _5572_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net322),
    .D(_0240_),
    .Q_N(_2424_),
    .Q(\mem[43][2] ));
 sg13g2_dfrbp_1 _5573_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net321),
    .D(_0241_),
    .Q_N(_2423_),
    .Q(\mem[43][3] ));
 sg13g2_dfrbp_1 _5574_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net320),
    .D(_0242_),
    .Q_N(_2422_),
    .Q(\mem[42][0] ));
 sg13g2_dfrbp_1 _5575_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net319),
    .D(_0243_),
    .Q_N(_2421_),
    .Q(\mem[42][1] ));
 sg13g2_dfrbp_1 _5576_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net318),
    .D(_0244_),
    .Q_N(_2420_),
    .Q(\mem[42][2] ));
 sg13g2_dfrbp_1 _5577_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net317),
    .D(_0245_),
    .Q_N(_2419_),
    .Q(\mem[42][3] ));
 sg13g2_dfrbp_1 _5578_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net316),
    .D(_0246_),
    .Q_N(_2418_),
    .Q(\mem[0][0] ));
 sg13g2_dfrbp_1 _5579_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net315),
    .D(_0247_),
    .Q_N(_2417_),
    .Q(\mem[0][1] ));
 sg13g2_dfrbp_1 _5580_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net314),
    .D(_0248_),
    .Q_N(_2416_),
    .Q(\mem[0][2] ));
 sg13g2_dfrbp_1 _5581_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net313),
    .D(_0249_),
    .Q_N(_0000_),
    .Q(\mem[0][3] ));
 sg13g2_dfrbp_1 _5582_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net312),
    .D(_0250_),
    .Q_N(_2415_),
    .Q(\mem[41][0] ));
 sg13g2_dfrbp_1 _5583_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net311),
    .D(_0251_),
    .Q_N(_2414_),
    .Q(\mem[41][1] ));
 sg13g2_dfrbp_1 _5584_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net310),
    .D(_0252_),
    .Q_N(_2413_),
    .Q(\mem[41][2] ));
 sg13g2_dfrbp_1 _5585_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net309),
    .D(_0253_),
    .Q_N(_2412_),
    .Q(\mem[41][3] ));
 sg13g2_dfrbp_1 _5586_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net308),
    .D(_0254_),
    .Q_N(_2411_),
    .Q(\mem[8][0] ));
 sg13g2_dfrbp_1 _5587_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net307),
    .D(_0255_),
    .Q_N(_2410_),
    .Q(\mem[8][1] ));
 sg13g2_dfrbp_1 _5588_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net306),
    .D(_0256_),
    .Q_N(_2409_),
    .Q(\mem[8][2] ));
 sg13g2_dfrbp_1 _5589_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net305),
    .D(_0257_),
    .Q_N(_2408_),
    .Q(\mem[8][3] ));
 sg13g2_dfrbp_1 _5590_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net304),
    .D(_0258_),
    .Q_N(_2407_),
    .Q(\mem[12][0] ));
 sg13g2_dfrbp_1 _5591_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net303),
    .D(_0259_),
    .Q_N(_2406_),
    .Q(\mem[12][1] ));
 sg13g2_dfrbp_1 _5592_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net302),
    .D(_0260_),
    .Q_N(_2405_),
    .Q(\mem[12][2] ));
 sg13g2_dfrbp_1 _5593_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net301),
    .D(_0261_),
    .Q_N(_2404_),
    .Q(\mem[12][3] ));
 sg13g2_dfrbp_1 _5594_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net300),
    .D(_0262_),
    .Q_N(_2403_),
    .Q(\mem[9][0] ));
 sg13g2_dfrbp_1 _5595_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net299),
    .D(_0263_),
    .Q_N(_2402_),
    .Q(\mem[9][1] ));
 sg13g2_dfrbp_1 _5596_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net298),
    .D(_0264_),
    .Q_N(_2401_),
    .Q(\mem[9][2] ));
 sg13g2_dfrbp_1 _5597_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net297),
    .D(_0265_),
    .Q_N(_2400_),
    .Q(\mem[9][3] ));
 sg13g2_dfrbp_1 _5598_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net296),
    .D(_0266_),
    .Q_N(_2399_),
    .Q(\products[15][0] ));
 sg13g2_dfrbp_1 _5599_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net295),
    .D(_0267_),
    .Q_N(_2398_),
    .Q(\products[15][1] ));
 sg13g2_dfrbp_1 _5600_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net294),
    .D(_0268_),
    .Q_N(_2397_),
    .Q(\products[15][2] ));
 sg13g2_dfrbp_1 _5601_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net293),
    .D(_0269_),
    .Q_N(_2396_),
    .Q(\products[15][3] ));
 sg13g2_dfrbp_1 _5602_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net292),
    .D(_0270_),
    .Q_N(_2395_),
    .Q(\products[15][4] ));
 sg13g2_dfrbp_1 _5603_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net291),
    .D(_0271_),
    .Q_N(_2394_),
    .Q(\products[15][5] ));
 sg13g2_dfrbp_1 _5604_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net290),
    .D(_0272_),
    .Q_N(_2393_),
    .Q(\products[15][6] ));
 sg13g2_dfrbp_1 _5605_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net289),
    .D(_0273_),
    .Q_N(_2392_),
    .Q(\products[15][7] ));
 sg13g2_dfrbp_1 _5606_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net288),
    .D(_0274_),
    .Q_N(_2391_),
    .Q(\products[14][0] ));
 sg13g2_dfrbp_1 _5607_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net287),
    .D(_0275_),
    .Q_N(_2390_),
    .Q(\products[14][1] ));
 sg13g2_dfrbp_1 _5608_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net286),
    .D(_0276_),
    .Q_N(_2389_),
    .Q(\products[14][2] ));
 sg13g2_dfrbp_1 _5609_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net285),
    .D(_0277_),
    .Q_N(_2388_),
    .Q(\products[14][3] ));
 sg13g2_dfrbp_1 _5610_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net284),
    .D(_0278_),
    .Q_N(_2387_),
    .Q(\products[14][4] ));
 sg13g2_dfrbp_1 _5611_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net283),
    .D(_0279_),
    .Q_N(_2386_),
    .Q(\products[14][5] ));
 sg13g2_dfrbp_1 _5612_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net282),
    .D(_0280_),
    .Q_N(_2385_),
    .Q(\products[14][6] ));
 sg13g2_dfrbp_1 _5613_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net281),
    .D(_0281_),
    .Q_N(_2384_),
    .Q(\products[14][7] ));
 sg13g2_dfrbp_1 _5614_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net280),
    .D(_0282_),
    .Q_N(_2383_),
    .Q(\products[13][0] ));
 sg13g2_dfrbp_1 _5615_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net279),
    .D(_0283_),
    .Q_N(_2382_),
    .Q(\products[13][1] ));
 sg13g2_dfrbp_1 _5616_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net278),
    .D(_0284_),
    .Q_N(_2381_),
    .Q(\products[13][2] ));
 sg13g2_dfrbp_1 _5617_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net277),
    .D(_0285_),
    .Q_N(_2380_),
    .Q(\products[13][3] ));
 sg13g2_dfrbp_1 _5618_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net276),
    .D(_0286_),
    .Q_N(_2379_),
    .Q(\products[13][4] ));
 sg13g2_dfrbp_1 _5619_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net275),
    .D(_0287_),
    .Q_N(_2378_),
    .Q(\products[13][5] ));
 sg13g2_dfrbp_1 _5620_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net274),
    .D(_0288_),
    .Q_N(_2377_),
    .Q(\products[13][6] ));
 sg13g2_dfrbp_1 _5621_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net273),
    .D(_0289_),
    .Q_N(_2376_),
    .Q(\products[13][7] ));
 sg13g2_dfrbp_1 _5622_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net272),
    .D(net717),
    .Q_N(_2375_),
    .Q(\products[12][0] ));
 sg13g2_dfrbp_1 _5623_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net271),
    .D(_0291_),
    .Q_N(_2374_),
    .Q(\products[12][1] ));
 sg13g2_dfrbp_1 _5624_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net270),
    .D(_0292_),
    .Q_N(_2373_),
    .Q(\products[12][2] ));
 sg13g2_dfrbp_1 _5625_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net269),
    .D(_0293_),
    .Q_N(_2372_),
    .Q(\products[12][3] ));
 sg13g2_dfrbp_1 _5626_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net268),
    .D(_0294_),
    .Q_N(_2371_),
    .Q(\products[12][4] ));
 sg13g2_dfrbp_1 _5627_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net267),
    .D(_0295_),
    .Q_N(_2370_),
    .Q(\products[12][5] ));
 sg13g2_dfrbp_1 _5628_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net266),
    .D(_0296_),
    .Q_N(_2369_),
    .Q(\products[12][6] ));
 sg13g2_dfrbp_1 _5629_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net265),
    .D(_0297_),
    .Q_N(_2368_),
    .Q(\products[12][7] ));
 sg13g2_dfrbp_1 _5630_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net264),
    .D(net675),
    .Q_N(_2367_),
    .Q(\products[11][0] ));
 sg13g2_dfrbp_1 _5631_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net263),
    .D(_0299_),
    .Q_N(_2366_),
    .Q(\products[11][1] ));
 sg13g2_dfrbp_1 _5632_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net262),
    .D(_0300_),
    .Q_N(_2365_),
    .Q(\products[11][2] ));
 sg13g2_dfrbp_1 _5633_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net261),
    .D(_0301_),
    .Q_N(_2364_),
    .Q(\products[11][3] ));
 sg13g2_dfrbp_1 _5634_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net260),
    .D(_0302_),
    .Q_N(_2363_),
    .Q(\products[11][4] ));
 sg13g2_dfrbp_1 _5635_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net259),
    .D(_0303_),
    .Q_N(_2362_),
    .Q(\products[11][5] ));
 sg13g2_dfrbp_1 _5636_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net258),
    .D(_0304_),
    .Q_N(_2361_),
    .Q(\products[11][6] ));
 sg13g2_dfrbp_1 _5637_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net257),
    .D(_0305_),
    .Q_N(_2360_),
    .Q(\products[11][7] ));
 sg13g2_dfrbp_1 _5638_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net256),
    .D(net738),
    .Q_N(_2359_),
    .Q(\products[10][0] ));
 sg13g2_dfrbp_1 _5639_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net255),
    .D(_0307_),
    .Q_N(_2358_),
    .Q(\products[10][1] ));
 sg13g2_dfrbp_1 _5640_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net254),
    .D(_0308_),
    .Q_N(_2357_),
    .Q(\products[10][2] ));
 sg13g2_dfrbp_1 _5641_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net253),
    .D(_0309_),
    .Q_N(_2356_),
    .Q(\products[10][3] ));
 sg13g2_dfrbp_1 _5642_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net252),
    .D(_0310_),
    .Q_N(_2355_),
    .Q(\products[10][4] ));
 sg13g2_dfrbp_1 _5643_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net251),
    .D(_0311_),
    .Q_N(_2354_),
    .Q(\products[10][5] ));
 sg13g2_dfrbp_1 _5644_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net250),
    .D(_0312_),
    .Q_N(_2353_),
    .Q(\products[10][6] ));
 sg13g2_dfrbp_1 _5645_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net249),
    .D(_0313_),
    .Q_N(_2352_),
    .Q(\products[10][7] ));
 sg13g2_dfrbp_1 _5646_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net248),
    .D(_0314_),
    .Q_N(_2351_),
    .Q(\products[9][0] ));
 sg13g2_dfrbp_1 _5647_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net247),
    .D(_0315_),
    .Q_N(_2350_),
    .Q(\products[9][1] ));
 sg13g2_dfrbp_1 _5648_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net246),
    .D(_0316_),
    .Q_N(_2349_),
    .Q(\products[9][2] ));
 sg13g2_dfrbp_1 _5649_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net245),
    .D(_0317_),
    .Q_N(_2348_),
    .Q(\products[9][3] ));
 sg13g2_dfrbp_1 _5650_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net244),
    .D(_0318_),
    .Q_N(_2347_),
    .Q(\products[9][4] ));
 sg13g2_dfrbp_1 _5651_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net243),
    .D(_0319_),
    .Q_N(_2346_),
    .Q(\products[9][5] ));
 sg13g2_dfrbp_1 _5652_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net242),
    .D(_0320_),
    .Q_N(_2345_),
    .Q(\products[9][6] ));
 sg13g2_dfrbp_1 _5653_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net241),
    .D(_0321_),
    .Q_N(_2344_),
    .Q(\products[9][7] ));
 sg13g2_dfrbp_1 _5654_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net240),
    .D(net698),
    .Q_N(_2343_),
    .Q(\products[8][0] ));
 sg13g2_dfrbp_1 _5655_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net239),
    .D(_0323_),
    .Q_N(_2342_),
    .Q(\products[8][1] ));
 sg13g2_dfrbp_1 _5656_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net238),
    .D(_0324_),
    .Q_N(_2341_),
    .Q(\products[8][2] ));
 sg13g2_dfrbp_1 _5657_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net237),
    .D(_0325_),
    .Q_N(_2340_),
    .Q(\products[8][3] ));
 sg13g2_dfrbp_1 _5658_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net236),
    .D(_0326_),
    .Q_N(_2339_),
    .Q(\products[8][4] ));
 sg13g2_dfrbp_1 _5659_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net235),
    .D(_0327_),
    .Q_N(_2338_),
    .Q(\products[8][5] ));
 sg13g2_dfrbp_1 _5660_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net234),
    .D(_0328_),
    .Q_N(_2337_),
    .Q(\products[8][6] ));
 sg13g2_dfrbp_1 _5661_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net233),
    .D(_0329_),
    .Q_N(_2336_),
    .Q(\products[8][7] ));
 sg13g2_dfrbp_1 _5662_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net232),
    .D(net706),
    .Q_N(_2335_),
    .Q(\products[7][0] ));
 sg13g2_dfrbp_1 _5663_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net231),
    .D(_0331_),
    .Q_N(_2334_),
    .Q(\products[7][1] ));
 sg13g2_dfrbp_1 _5664_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net230),
    .D(_0332_),
    .Q_N(_2333_),
    .Q(\products[7][2] ));
 sg13g2_dfrbp_1 _5665_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net229),
    .D(_0333_),
    .Q_N(_2332_),
    .Q(\products[7][3] ));
 sg13g2_dfrbp_1 _5666_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net228),
    .D(_0334_),
    .Q_N(_2331_),
    .Q(\products[7][4] ));
 sg13g2_dfrbp_1 _5667_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net227),
    .D(_0335_),
    .Q_N(_2330_),
    .Q(\products[7][5] ));
 sg13g2_dfrbp_1 _5668_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net226),
    .D(_0336_),
    .Q_N(_2329_),
    .Q(\products[7][6] ));
 sg13g2_dfrbp_1 _5669_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net225),
    .D(net408),
    .Q_N(_2328_),
    .Q(\products[7][7] ));
 sg13g2_dfrbp_1 _5670_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net224),
    .D(net708),
    .Q_N(_2327_),
    .Q(\products[6][0] ));
 sg13g2_dfrbp_1 _5671_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net223),
    .D(_0339_),
    .Q_N(_2326_),
    .Q(\products[6][1] ));
 sg13g2_dfrbp_1 _5672_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net222),
    .D(_0340_),
    .Q_N(_2325_),
    .Q(\products[6][2] ));
 sg13g2_dfrbp_1 _5673_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net221),
    .D(_0341_),
    .Q_N(_2324_),
    .Q(\products[6][3] ));
 sg13g2_dfrbp_1 _5674_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net220),
    .D(_0342_),
    .Q_N(_2323_),
    .Q(\products[6][4] ));
 sg13g2_dfrbp_1 _5675_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net219),
    .D(_0343_),
    .Q_N(_2322_),
    .Q(\products[6][5] ));
 sg13g2_dfrbp_1 _5676_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net218),
    .D(_0344_),
    .Q_N(_2321_),
    .Q(\products[6][6] ));
 sg13g2_dfrbp_1 _5677_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net217),
    .D(_0345_),
    .Q_N(_2320_),
    .Q(\products[6][7] ));
 sg13g2_dfrbp_1 _5678_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net216),
    .D(_0346_),
    .Q_N(_2319_),
    .Q(\products[5][0] ));
 sg13g2_dfrbp_1 _5679_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net215),
    .D(_0347_),
    .Q_N(_2318_),
    .Q(\products[5][1] ));
 sg13g2_dfrbp_1 _5680_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net214),
    .D(_0348_),
    .Q_N(_2317_),
    .Q(\products[5][2] ));
 sg13g2_dfrbp_1 _5681_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net213),
    .D(_0349_),
    .Q_N(_2316_),
    .Q(\products[5][3] ));
 sg13g2_dfrbp_1 _5682_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net212),
    .D(_0350_),
    .Q_N(_2315_),
    .Q(\products[5][4] ));
 sg13g2_dfrbp_1 _5683_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net211),
    .D(_0351_),
    .Q_N(_2314_),
    .Q(\products[5][5] ));
 sg13g2_dfrbp_1 _5684_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net210),
    .D(_0352_),
    .Q_N(_2313_),
    .Q(\products[5][6] ));
 sg13g2_dfrbp_1 _5685_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net209),
    .D(_0353_),
    .Q_N(_2312_),
    .Q(\products[5][7] ));
 sg13g2_dfrbp_1 _5686_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net208),
    .D(net410),
    .Q_N(_2311_),
    .Q(\products[4][0] ));
 sg13g2_dfrbp_1 _5687_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net207),
    .D(net817),
    .Q_N(_2310_),
    .Q(\products[4][1] ));
 sg13g2_dfrbp_1 _5688_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net206),
    .D(_0356_),
    .Q_N(_2309_),
    .Q(\products[4][2] ));
 sg13g2_dfrbp_1 _5689_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net205),
    .D(_0357_),
    .Q_N(_2308_),
    .Q(\products[4][3] ));
 sg13g2_dfrbp_1 _5690_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net204),
    .D(_0358_),
    .Q_N(_2307_),
    .Q(\products[4][4] ));
 sg13g2_dfrbp_1 _5691_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net203),
    .D(_0359_),
    .Q_N(_2306_),
    .Q(\products[4][5] ));
 sg13g2_dfrbp_1 _5692_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net202),
    .D(_0360_),
    .Q_N(_2305_),
    .Q(\products[4][6] ));
 sg13g2_dfrbp_1 _5693_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net201),
    .D(_0361_),
    .Q_N(_2304_),
    .Q(\products[4][7] ));
 sg13g2_dfrbp_1 _5694_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net200),
    .D(_0362_),
    .Q_N(_2303_),
    .Q(\products[3][0] ));
 sg13g2_dfrbp_1 _5695_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net199),
    .D(_0363_),
    .Q_N(_2302_),
    .Q(\products[3][1] ));
 sg13g2_dfrbp_1 _5696_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net198),
    .D(_0364_),
    .Q_N(_2301_),
    .Q(\products[3][2] ));
 sg13g2_dfrbp_1 _5697_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net197),
    .D(_0365_),
    .Q_N(_2300_),
    .Q(\products[3][3] ));
 sg13g2_dfrbp_1 _5698_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net196),
    .D(_0366_),
    .Q_N(_2299_),
    .Q(\products[3][4] ));
 sg13g2_dfrbp_1 _5699_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net195),
    .D(_0367_),
    .Q_N(_2298_),
    .Q(\products[3][5] ));
 sg13g2_dfrbp_1 _5700_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net194),
    .D(_0368_),
    .Q_N(_2297_),
    .Q(\products[3][6] ));
 sg13g2_dfrbp_1 _5701_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net193),
    .D(_0369_),
    .Q_N(_2296_),
    .Q(\products[3][7] ));
 sg13g2_dfrbp_1 _5702_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net192),
    .D(_0370_),
    .Q_N(_2295_),
    .Q(\products[2][0] ));
 sg13g2_dfrbp_1 _5703_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net191),
    .D(_0371_),
    .Q_N(_2294_),
    .Q(\products[2][1] ));
 sg13g2_dfrbp_1 _5704_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net190),
    .D(net858),
    .Q_N(_2293_),
    .Q(\products[2][2] ));
 sg13g2_dfrbp_1 _5705_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net189),
    .D(_0373_),
    .Q_N(_2292_),
    .Q(\products[2][3] ));
 sg13g2_dfrbp_1 _5706_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net188),
    .D(_0374_),
    .Q_N(_2291_),
    .Q(\products[2][4] ));
 sg13g2_dfrbp_1 _5707_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net187),
    .D(_0375_),
    .Q_N(_2290_),
    .Q(\products[2][5] ));
 sg13g2_dfrbp_1 _5708_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net186),
    .D(_0376_),
    .Q_N(_2289_),
    .Q(\products[2][6] ));
 sg13g2_dfrbp_1 _5709_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net185),
    .D(_0377_),
    .Q_N(_2288_),
    .Q(\products[2][7] ));
 sg13g2_dfrbp_1 _5710_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net184),
    .D(net685),
    .Q_N(_2287_),
    .Q(\products[1][0] ));
 sg13g2_dfrbp_1 _5711_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net183),
    .D(_0379_),
    .Q_N(_2286_),
    .Q(\products[1][1] ));
 sg13g2_dfrbp_1 _5712_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net182),
    .D(_0380_),
    .Q_N(_2285_),
    .Q(\products[1][2] ));
 sg13g2_dfrbp_1 _5713_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net181),
    .D(_0381_),
    .Q_N(_2284_),
    .Q(\products[1][3] ));
 sg13g2_dfrbp_1 _5714_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net180),
    .D(_0382_),
    .Q_N(_2283_),
    .Q(\products[1][4] ));
 sg13g2_dfrbp_1 _5715_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net179),
    .D(_0383_),
    .Q_N(_2282_),
    .Q(\products[1][5] ));
 sg13g2_dfrbp_1 _5716_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net178),
    .D(_0384_),
    .Q_N(_2281_),
    .Q(\products[1][6] ));
 sg13g2_dfrbp_1 _5717_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net177),
    .D(_0385_),
    .Q_N(_2280_),
    .Q(\products[1][7] ));
 sg13g2_dfrbp_1 _5718_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net176),
    .D(_0386_),
    .Q_N(_2279_),
    .Q(uio_out[5]));
 sg13g2_dfrbp_1 _5719_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net174),
    .D(net679),
    .Q_N(_2278_),
    .Q(\prev_acc[0] ));
 sg13g2_dfrbp_1 _5720_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net172),
    .D(net683),
    .Q_N(_2277_),
    .Q(\prev_acc[1] ));
 sg13g2_dfrbp_1 _5721_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net170),
    .D(net692),
    .Q_N(_2276_),
    .Q(\prev_acc[2] ));
 sg13g2_dfrbp_1 _5722_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net168),
    .D(net694),
    .Q_N(_2275_),
    .Q(\prev_acc[3] ));
 sg13g2_dfrbp_1 _5723_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net175),
    .D(net710),
    .Q_N(_2274_),
    .Q(\prev_acc[4] ));
 sg13g2_dfrbp_1 _5724_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net171),
    .D(_0392_),
    .Q_N(_2273_),
    .Q(\prev_acc[5] ));
 sg13g2_dfrbp_1 _5725_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net19),
    .D(net687),
    .Q_N(_2272_),
    .Q(\prev_acc[6] ));
 sg13g2_dfrbp_1 _5726_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net169),
    .D(net696),
    .Q_N(_2271_),
    .Q(\prev_acc[7] ));
 sg13g2_tiehi _5488__12 (.L_HI(net12));
 sg13g2_tiehi _5487__13 (.L_HI(net13));
 sg13g2_tiehi _5486__14 (.L_HI(net14));
 sg13g2_tiehi _5485__15 (.L_HI(net15));
 sg13g2_tiehi _5484__16 (.L_HI(net16));
 sg13g2_tiehi _5483__17 (.L_HI(net17));
 sg13g2_tiehi _5482__18 (.L_HI(net18));
 sg13g2_tiehi _5725__19 (.L_HI(net19));
 sg13g2_tiehi _5481__20 (.L_HI(net20));
 sg13g2_tiehi _5480__21 (.L_HI(net21));
 sg13g2_tiehi _5479__22 (.L_HI(net22));
 sg13g2_tiehi _5478__23 (.L_HI(net23));
 sg13g2_tiehi _5477__24 (.L_HI(net24));
 sg13g2_tiehi _5476__25 (.L_HI(net25));
 sg13g2_tiehi _5475__26 (.L_HI(net26));
 sg13g2_tiehi _5474__27 (.L_HI(net27));
 sg13g2_tiehi _5473__28 (.L_HI(net28));
 sg13g2_tiehi _5472__29 (.L_HI(net29));
 sg13g2_tiehi _5471__30 (.L_HI(net30));
 sg13g2_tiehi _5470__31 (.L_HI(net31));
 sg13g2_tiehi _5469__32 (.L_HI(net32));
 sg13g2_tiehi _5468__33 (.L_HI(net33));
 sg13g2_tiehi _5467__34 (.L_HI(net34));
 sg13g2_tiehi _5466__35 (.L_HI(net35));
 sg13g2_tiehi _5465__36 (.L_HI(net36));
 sg13g2_tiehi _5464__37 (.L_HI(net37));
 sg13g2_tiehi _5463__38 (.L_HI(net38));
 sg13g2_tiehi _5462__39 (.L_HI(net39));
 sg13g2_tiehi _5461__40 (.L_HI(net40));
 sg13g2_tiehi _5460__41 (.L_HI(net41));
 sg13g2_tiehi _5459__42 (.L_HI(net42));
 sg13g2_tiehi _5458__43 (.L_HI(net43));
 sg13g2_tiehi _5457__44 (.L_HI(net44));
 sg13g2_tiehi _5456__45 (.L_HI(net45));
 sg13g2_tiehi _5455__46 (.L_HI(net46));
 sg13g2_tiehi _5454__47 (.L_HI(net47));
 sg13g2_tiehi _5453__48 (.L_HI(net48));
 sg13g2_tiehi _5452__49 (.L_HI(net49));
 sg13g2_tiehi _5451__50 (.L_HI(net50));
 sg13g2_tiehi _5450__51 (.L_HI(net51));
 sg13g2_tiehi _5449__52 (.L_HI(net52));
 sg13g2_tiehi _5448__53 (.L_HI(net53));
 sg13g2_tiehi _5447__54 (.L_HI(net54));
 sg13g2_tiehi _5446__55 (.L_HI(net55));
 sg13g2_tiehi _5445__56 (.L_HI(net56));
 sg13g2_tiehi _5444__57 (.L_HI(net57));
 sg13g2_tiehi _5443__58 (.L_HI(net58));
 sg13g2_tiehi _5442__59 (.L_HI(net59));
 sg13g2_tiehi _5441__60 (.L_HI(net60));
 sg13g2_tiehi _5440__61 (.L_HI(net61));
 sg13g2_tiehi _5439__62 (.L_HI(net62));
 sg13g2_tiehi _5438__63 (.L_HI(net63));
 sg13g2_tiehi _5437__64 (.L_HI(net64));
 sg13g2_tiehi _5436__65 (.L_HI(net65));
 sg13g2_tiehi _5435__66 (.L_HI(net66));
 sg13g2_tiehi _5434__67 (.L_HI(net67));
 sg13g2_tiehi _5433__68 (.L_HI(net68));
 sg13g2_tiehi _5432__69 (.L_HI(net69));
 sg13g2_tiehi _5431__70 (.L_HI(net70));
 sg13g2_tiehi _5430__71 (.L_HI(net71));
 sg13g2_tiehi _5429__72 (.L_HI(net72));
 sg13g2_tiehi _5428__73 (.L_HI(net73));
 sg13g2_tiehi _5427__74 (.L_HI(net74));
 sg13g2_tiehi _5426__75 (.L_HI(net75));
 sg13g2_tiehi _5425__76 (.L_HI(net76));
 sg13g2_tiehi _5424__77 (.L_HI(net77));
 sg13g2_tiehi _5423__78 (.L_HI(net78));
 sg13g2_tiehi _5422__79 (.L_HI(net79));
 sg13g2_tiehi _5421__80 (.L_HI(net80));
 sg13g2_tiehi _5420__81 (.L_HI(net81));
 sg13g2_tiehi _5419__82 (.L_HI(net82));
 sg13g2_tiehi _5418__83 (.L_HI(net83));
 sg13g2_tiehi _5417__84 (.L_HI(net84));
 sg13g2_tiehi _5416__85 (.L_HI(net85));
 sg13g2_tiehi _5415__86 (.L_HI(net86));
 sg13g2_tiehi _5414__87 (.L_HI(net87));
 sg13g2_tiehi _5413__88 (.L_HI(net88));
 sg13g2_tiehi _5412__89 (.L_HI(net89));
 sg13g2_tiehi _5411__90 (.L_HI(net90));
 sg13g2_tiehi _5410__91 (.L_HI(net91));
 sg13g2_tiehi _5409__92 (.L_HI(net92));
 sg13g2_tiehi _5408__93 (.L_HI(net93));
 sg13g2_tiehi _5407__94 (.L_HI(net94));
 sg13g2_tiehi _5406__95 (.L_HI(net95));
 sg13g2_tiehi _5405__96 (.L_HI(net96));
 sg13g2_tiehi _5404__97 (.L_HI(net97));
 sg13g2_tiehi _5403__98 (.L_HI(net98));
 sg13g2_tiehi _5402__99 (.L_HI(net99));
 sg13g2_tiehi _5401__100 (.L_HI(net100));
 sg13g2_tiehi _5400__101 (.L_HI(net101));
 sg13g2_tiehi _5399__102 (.L_HI(net102));
 sg13g2_tiehi _5398__103 (.L_HI(net103));
 sg13g2_tiehi _5397__104 (.L_HI(net104));
 sg13g2_tiehi _5396__105 (.L_HI(net105));
 sg13g2_tiehi _5395__106 (.L_HI(net106));
 sg13g2_tiehi _5394__107 (.L_HI(net107));
 sg13g2_tiehi _5393__108 (.L_HI(net108));
 sg13g2_tiehi _5392__109 (.L_HI(net109));
 sg13g2_tiehi _5391__110 (.L_HI(net110));
 sg13g2_tiehi _5390__111 (.L_HI(net111));
 sg13g2_tiehi _5389__112 (.L_HI(net112));
 sg13g2_tiehi _5388__113 (.L_HI(net113));
 sg13g2_tiehi _5387__114 (.L_HI(net114));
 sg13g2_tiehi _5386__115 (.L_HI(net115));
 sg13g2_tiehi _5385__116 (.L_HI(net116));
 sg13g2_tiehi _5384__117 (.L_HI(net117));
 sg13g2_tiehi _5383__118 (.L_HI(net118));
 sg13g2_tiehi _5382__119 (.L_HI(net119));
 sg13g2_tiehi _5381__120 (.L_HI(net120));
 sg13g2_tiehi _5380__121 (.L_HI(net121));
 sg13g2_tiehi _5379__122 (.L_HI(net122));
 sg13g2_tiehi _5378__123 (.L_HI(net123));
 sg13g2_tiehi _5377__124 (.L_HI(net124));
 sg13g2_tiehi _5376__125 (.L_HI(net125));
 sg13g2_tiehi _5375__126 (.L_HI(net126));
 sg13g2_tiehi _5374__127 (.L_HI(net127));
 sg13g2_tiehi _5373__128 (.L_HI(net128));
 sg13g2_tiehi _5372__129 (.L_HI(net129));
 sg13g2_tiehi _5371__130 (.L_HI(net130));
 sg13g2_tiehi _5370__131 (.L_HI(net131));
 sg13g2_tiehi _5369__132 (.L_HI(net132));
 sg13g2_tiehi _5368__133 (.L_HI(net133));
 sg13g2_tiehi _5367__134 (.L_HI(net134));
 sg13g2_tiehi _5366__135 (.L_HI(net135));
 sg13g2_tiehi _5365__136 (.L_HI(net136));
 sg13g2_tiehi _5364__137 (.L_HI(net137));
 sg13g2_tiehi _5363__138 (.L_HI(net138));
 sg13g2_tiehi _5362__139 (.L_HI(net139));
 sg13g2_tiehi _5361__140 (.L_HI(net140));
 sg13g2_tiehi _5360__141 (.L_HI(net141));
 sg13g2_tiehi _5359__142 (.L_HI(net142));
 sg13g2_tiehi _5358__143 (.L_HI(net143));
 sg13g2_tiehi _5357__144 (.L_HI(net144));
 sg13g2_tiehi _5356__145 (.L_HI(net145));
 sg13g2_tiehi _5355__146 (.L_HI(net146));
 sg13g2_tiehi _5354__147 (.L_HI(net147));
 sg13g2_tiehi _5353__148 (.L_HI(net148));
 sg13g2_tiehi _5352__149 (.L_HI(net149));
 sg13g2_tiehi _5351__150 (.L_HI(net150));
 sg13g2_tiehi _5350__151 (.L_HI(net151));
 sg13g2_tiehi _5349__152 (.L_HI(net152));
 sg13g2_tiehi _5348__153 (.L_HI(net153));
 sg13g2_tiehi _5347__154 (.L_HI(net154));
 sg13g2_tiehi _5346__155 (.L_HI(net155));
 sg13g2_tiehi _5345__156 (.L_HI(net156));
 sg13g2_tiehi _5344__157 (.L_HI(net157));
 sg13g2_tiehi _5343__158 (.L_HI(net158));
 sg13g2_tiehi _5342__159 (.L_HI(net159));
 sg13g2_tiehi _5341__160 (.L_HI(net160));
 sg13g2_tiehi _5340__161 (.L_HI(net161));
 sg13g2_tiehi _5339__162 (.L_HI(net162));
 sg13g2_tiehi _5338__163 (.L_HI(net163));
 sg13g2_tiehi _5337__164 (.L_HI(net164));
 sg13g2_tiehi _5336__165 (.L_HI(net165));
 sg13g2_tiehi _5335__166 (.L_HI(net166));
 sg13g2_tiehi _5334__167 (.L_HI(net167));
 sg13g2_tiehi _5722__168 (.L_HI(net168));
 sg13g2_tiehi _5726__169 (.L_HI(net169));
 sg13g2_tiehi _5721__170 (.L_HI(net170));
 sg13g2_tiehi _5724__171 (.L_HI(net171));
 sg13g2_tiehi _5720__172 (.L_HI(net172));
 sg13g2_tiehi _5333__173 (.L_HI(net173));
 sg13g2_tiehi _5719__174 (.L_HI(net174));
 sg13g2_tiehi _5723__175 (.L_HI(net175));
 sg13g2_tiehi _5718__176 (.L_HI(net176));
 sg13g2_tiehi _5717__177 (.L_HI(net177));
 sg13g2_tiehi _5716__178 (.L_HI(net178));
 sg13g2_tiehi _5715__179 (.L_HI(net179));
 sg13g2_tiehi _5714__180 (.L_HI(net180));
 sg13g2_tiehi _5713__181 (.L_HI(net181));
 sg13g2_tiehi _5712__182 (.L_HI(net182));
 sg13g2_tiehi _5711__183 (.L_HI(net183));
 sg13g2_tiehi _5710__184 (.L_HI(net184));
 sg13g2_tiehi _5709__185 (.L_HI(net185));
 sg13g2_tiehi _5708__186 (.L_HI(net186));
 sg13g2_tiehi _5707__187 (.L_HI(net187));
 sg13g2_tiehi _5706__188 (.L_HI(net188));
 sg13g2_tiehi _5705__189 (.L_HI(net189));
 sg13g2_tiehi _5704__190 (.L_HI(net190));
 sg13g2_tiehi _5703__191 (.L_HI(net191));
 sg13g2_tiehi _5702__192 (.L_HI(net192));
 sg13g2_tiehi _5701__193 (.L_HI(net193));
 sg13g2_tiehi _5700__194 (.L_HI(net194));
 sg13g2_tiehi _5699__195 (.L_HI(net195));
 sg13g2_tiehi _5698__196 (.L_HI(net196));
 sg13g2_tiehi _5697__197 (.L_HI(net197));
 sg13g2_tiehi _5696__198 (.L_HI(net198));
 sg13g2_tiehi _5695__199 (.L_HI(net199));
 sg13g2_tiehi _5694__200 (.L_HI(net200));
 sg13g2_tiehi _5693__201 (.L_HI(net201));
 sg13g2_tiehi _5692__202 (.L_HI(net202));
 sg13g2_tiehi _5691__203 (.L_HI(net203));
 sg13g2_tiehi _5690__204 (.L_HI(net204));
 sg13g2_tiehi _5689__205 (.L_HI(net205));
 sg13g2_tiehi _5688__206 (.L_HI(net206));
 sg13g2_tiehi _5687__207 (.L_HI(net207));
 sg13g2_tiehi _5686__208 (.L_HI(net208));
 sg13g2_tiehi _5685__209 (.L_HI(net209));
 sg13g2_tiehi _5684__210 (.L_HI(net210));
 sg13g2_tiehi _5683__211 (.L_HI(net211));
 sg13g2_tiehi _5682__212 (.L_HI(net212));
 sg13g2_tiehi _5681__213 (.L_HI(net213));
 sg13g2_tiehi _5680__214 (.L_HI(net214));
 sg13g2_tiehi _5679__215 (.L_HI(net215));
 sg13g2_tiehi _5678__216 (.L_HI(net216));
 sg13g2_tiehi _5677__217 (.L_HI(net217));
 sg13g2_tiehi _5676__218 (.L_HI(net218));
 sg13g2_tiehi _5675__219 (.L_HI(net219));
 sg13g2_tiehi _5674__220 (.L_HI(net220));
 sg13g2_tiehi _5673__221 (.L_HI(net221));
 sg13g2_tiehi _5672__222 (.L_HI(net222));
 sg13g2_tiehi _5671__223 (.L_HI(net223));
 sg13g2_tiehi _5670__224 (.L_HI(net224));
 sg13g2_tiehi _5669__225 (.L_HI(net225));
 sg13g2_tiehi _5668__226 (.L_HI(net226));
 sg13g2_tiehi _5667__227 (.L_HI(net227));
 sg13g2_tiehi _5666__228 (.L_HI(net228));
 sg13g2_tiehi _5665__229 (.L_HI(net229));
 sg13g2_tiehi _5664__230 (.L_HI(net230));
 sg13g2_tiehi _5663__231 (.L_HI(net231));
 sg13g2_tiehi _5662__232 (.L_HI(net232));
 sg13g2_tiehi _5661__233 (.L_HI(net233));
 sg13g2_tiehi _5660__234 (.L_HI(net234));
 sg13g2_tiehi _5659__235 (.L_HI(net235));
 sg13g2_tiehi _5658__236 (.L_HI(net236));
 sg13g2_tiehi _5657__237 (.L_HI(net237));
 sg13g2_tiehi _5656__238 (.L_HI(net238));
 sg13g2_tiehi _5655__239 (.L_HI(net239));
 sg13g2_tiehi _5654__240 (.L_HI(net240));
 sg13g2_tiehi _5653__241 (.L_HI(net241));
 sg13g2_tiehi _5652__242 (.L_HI(net242));
 sg13g2_tiehi _5651__243 (.L_HI(net243));
 sg13g2_tiehi _5650__244 (.L_HI(net244));
 sg13g2_tiehi _5649__245 (.L_HI(net245));
 sg13g2_tiehi _5648__246 (.L_HI(net246));
 sg13g2_tiehi _5647__247 (.L_HI(net247));
 sg13g2_tiehi _5646__248 (.L_HI(net248));
 sg13g2_tiehi _5645__249 (.L_HI(net249));
 sg13g2_tiehi _5644__250 (.L_HI(net250));
 sg13g2_tiehi _5643__251 (.L_HI(net251));
 sg13g2_tiehi _5642__252 (.L_HI(net252));
 sg13g2_tiehi _5641__253 (.L_HI(net253));
 sg13g2_tiehi _5640__254 (.L_HI(net254));
 sg13g2_tiehi _5639__255 (.L_HI(net255));
 sg13g2_tiehi _5638__256 (.L_HI(net256));
 sg13g2_tiehi _5637__257 (.L_HI(net257));
 sg13g2_tiehi _5636__258 (.L_HI(net258));
 sg13g2_tiehi _5635__259 (.L_HI(net259));
 sg13g2_tiehi _5634__260 (.L_HI(net260));
 sg13g2_tiehi _5633__261 (.L_HI(net261));
 sg13g2_tiehi _5632__262 (.L_HI(net262));
 sg13g2_tiehi _5631__263 (.L_HI(net263));
 sg13g2_tiehi _5630__264 (.L_HI(net264));
 sg13g2_tiehi _5629__265 (.L_HI(net265));
 sg13g2_tiehi _5628__266 (.L_HI(net266));
 sg13g2_tiehi _5627__267 (.L_HI(net267));
 sg13g2_tiehi _5626__268 (.L_HI(net268));
 sg13g2_tiehi _5625__269 (.L_HI(net269));
 sg13g2_tiehi _5624__270 (.L_HI(net270));
 sg13g2_tiehi _5623__271 (.L_HI(net271));
 sg13g2_tiehi _5622__272 (.L_HI(net272));
 sg13g2_tiehi _5621__273 (.L_HI(net273));
 sg13g2_tiehi _5620__274 (.L_HI(net274));
 sg13g2_tiehi _5619__275 (.L_HI(net275));
 sg13g2_tiehi _5618__276 (.L_HI(net276));
 sg13g2_tiehi _5617__277 (.L_HI(net277));
 sg13g2_tiehi _5616__278 (.L_HI(net278));
 sg13g2_tiehi _5615__279 (.L_HI(net279));
 sg13g2_tiehi _5614__280 (.L_HI(net280));
 sg13g2_tiehi _5613__281 (.L_HI(net281));
 sg13g2_tiehi _5612__282 (.L_HI(net282));
 sg13g2_tiehi _5611__283 (.L_HI(net283));
 sg13g2_tiehi _5610__284 (.L_HI(net284));
 sg13g2_tiehi _5609__285 (.L_HI(net285));
 sg13g2_tiehi _5608__286 (.L_HI(net286));
 sg13g2_tiehi _5607__287 (.L_HI(net287));
 sg13g2_tiehi _5606__288 (.L_HI(net288));
 sg13g2_tiehi _5605__289 (.L_HI(net289));
 sg13g2_tiehi _5604__290 (.L_HI(net290));
 sg13g2_tiehi _5603__291 (.L_HI(net291));
 sg13g2_tiehi _5602__292 (.L_HI(net292));
 sg13g2_tiehi _5601__293 (.L_HI(net293));
 sg13g2_tiehi _5600__294 (.L_HI(net294));
 sg13g2_tiehi _5599__295 (.L_HI(net295));
 sg13g2_tiehi _5598__296 (.L_HI(net296));
 sg13g2_tiehi _5597__297 (.L_HI(net297));
 sg13g2_tiehi _5596__298 (.L_HI(net298));
 sg13g2_tiehi _5595__299 (.L_HI(net299));
 sg13g2_tiehi _5594__300 (.L_HI(net300));
 sg13g2_tiehi _5593__301 (.L_HI(net301));
 sg13g2_tiehi _5592__302 (.L_HI(net302));
 sg13g2_tiehi _5591__303 (.L_HI(net303));
 sg13g2_tiehi _5590__304 (.L_HI(net304));
 sg13g2_tiehi _5589__305 (.L_HI(net305));
 sg13g2_tiehi _5588__306 (.L_HI(net306));
 sg13g2_tiehi _5587__307 (.L_HI(net307));
 sg13g2_tiehi _5586__308 (.L_HI(net308));
 sg13g2_tiehi _5585__309 (.L_HI(net309));
 sg13g2_tiehi _5584__310 (.L_HI(net310));
 sg13g2_tiehi _5583__311 (.L_HI(net311));
 sg13g2_tiehi _5582__312 (.L_HI(net312));
 sg13g2_tiehi _5581__313 (.L_HI(net313));
 sg13g2_tiehi _5580__314 (.L_HI(net314));
 sg13g2_tiehi _5579__315 (.L_HI(net315));
 sg13g2_tiehi _5578__316 (.L_HI(net316));
 sg13g2_tiehi _5577__317 (.L_HI(net317));
 sg13g2_tiehi _5576__318 (.L_HI(net318));
 sg13g2_tiehi _5575__319 (.L_HI(net319));
 sg13g2_tiehi _5574__320 (.L_HI(net320));
 sg13g2_tiehi _5573__321 (.L_HI(net321));
 sg13g2_tiehi _5572__322 (.L_HI(net322));
 sg13g2_tiehi _5571__323 (.L_HI(net323));
 sg13g2_tiehi _5570__324 (.L_HI(net324));
 sg13g2_tiehi _5569__325 (.L_HI(net325));
 sg13g2_tiehi _5568__326 (.L_HI(net326));
 sg13g2_tiehi _5567__327 (.L_HI(net327));
 sg13g2_tiehi _5566__328 (.L_HI(net328));
 sg13g2_tiehi _5565__329 (.L_HI(net329));
 sg13g2_tiehi _5564__330 (.L_HI(net330));
 sg13g2_tiehi _5563__331 (.L_HI(net331));
 sg13g2_tiehi _5562__332 (.L_HI(net332));
 sg13g2_tiehi _5561__333 (.L_HI(net333));
 sg13g2_tiehi _5560__334 (.L_HI(net334));
 sg13g2_tiehi _5559__335 (.L_HI(net335));
 sg13g2_tiehi _5558__336 (.L_HI(net336));
 sg13g2_tiehi _5557__337 (.L_HI(net337));
 sg13g2_tiehi _5556__338 (.L_HI(net338));
 sg13g2_tiehi _5555__339 (.L_HI(net339));
 sg13g2_tiehi _5554__340 (.L_HI(net340));
 sg13g2_tiehi _5553__341 (.L_HI(net341));
 sg13g2_tiehi _5552__342 (.L_HI(net342));
 sg13g2_tiehi _5551__343 (.L_HI(net343));
 sg13g2_tiehi _5550__344 (.L_HI(net344));
 sg13g2_tiehi _5549__345 (.L_HI(net345));
 sg13g2_tiehi _5548__346 (.L_HI(net346));
 sg13g2_tiehi _5547__347 (.L_HI(net347));
 sg13g2_tiehi _5546__348 (.L_HI(net348));
 sg13g2_tiehi _5545__349 (.L_HI(net349));
 sg13g2_tiehi _5544__350 (.L_HI(net350));
 sg13g2_tiehi _5543__351 (.L_HI(net351));
 sg13g2_tiehi _5542__352 (.L_HI(net352));
 sg13g2_tiehi _5541__353 (.L_HI(net353));
 sg13g2_tiehi _5540__354 (.L_HI(net354));
 sg13g2_tiehi _5539__355 (.L_HI(net355));
 sg13g2_tiehi _5538__356 (.L_HI(net356));
 sg13g2_tiehi _5537__357 (.L_HI(net357));
 sg13g2_tiehi _5536__358 (.L_HI(net358));
 sg13g2_tiehi _5535__359 (.L_HI(net359));
 sg13g2_tiehi _5534__360 (.L_HI(net360));
 sg13g2_tiehi _5533__361 (.L_HI(net361));
 sg13g2_tiehi _5532__362 (.L_HI(net362));
 sg13g2_tiehi _5531__363 (.L_HI(net363));
 sg13g2_tiehi _5530__364 (.L_HI(net364));
 sg13g2_tiehi _5529__365 (.L_HI(net365));
 sg13g2_tiehi _5528__366 (.L_HI(net366));
 sg13g2_tiehi _5527__367 (.L_HI(net367));
 sg13g2_tiehi _5526__368 (.L_HI(net368));
 sg13g2_tiehi _5525__369 (.L_HI(net369));
 sg13g2_tiehi _5524__370 (.L_HI(net370));
 sg13g2_tiehi _5523__371 (.L_HI(net371));
 sg13g2_tiehi _5522__372 (.L_HI(net372));
 sg13g2_tiehi _5521__373 (.L_HI(net373));
 sg13g2_tiehi _5520__374 (.L_HI(net374));
 sg13g2_tiehi _5519__375 (.L_HI(net375));
 sg13g2_tiehi _5518__376 (.L_HI(net376));
 sg13g2_tiehi _5517__377 (.L_HI(net377));
 sg13g2_tiehi _5516__378 (.L_HI(net378));
 sg13g2_tiehi _5515__379 (.L_HI(net379));
 sg13g2_tiehi _5514__380 (.L_HI(net380));
 sg13g2_tiehi _5513__381 (.L_HI(net381));
 sg13g2_tiehi _5512__382 (.L_HI(net382));
 sg13g2_tiehi _5511__383 (.L_HI(net383));
 sg13g2_tiehi _5510__384 (.L_HI(net384));
 sg13g2_tiehi _5509__385 (.L_HI(net385));
 sg13g2_tiehi _5508__386 (.L_HI(net386));
 sg13g2_tiehi _5507__387 (.L_HI(net387));
 sg13g2_tiehi _5506__388 (.L_HI(net388));
 sg13g2_tiehi _5505__389 (.L_HI(net389));
 sg13g2_tiehi _5504__390 (.L_HI(net390));
 sg13g2_tiehi _5503__391 (.L_HI(net391));
 sg13g2_tiehi _5502__392 (.L_HI(net392));
 sg13g2_tiehi _5501__393 (.L_HI(net393));
 sg13g2_tiehi _5500__394 (.L_HI(net394));
 sg13g2_tiehi _5499__395 (.L_HI(net395));
 sg13g2_tiehi _5498__396 (.L_HI(net396));
 sg13g2_tiehi _5497__397 (.L_HI(net397));
 sg13g2_tiehi _5496__398 (.L_HI(net398));
 sg13g2_tiehi _5495__399 (.L_HI(net399));
 sg13g2_tiehi _5494__400 (.L_HI(net400));
 sg13g2_tiehi _5493__401 (.L_HI(net401));
 sg13g2_tiehi _5492__402 (.L_HI(net402));
 sg13g2_tiehi _5491__403 (.L_HI(net403));
 sg13g2_tiehi _5490__404 (.L_HI(net404));
 sg13g2_tiehi tt_um_jayjaywong12_405 (.L_HI(net405));
 sg13g2_tiehi tt_um_jayjaywong12_406 (.L_HI(net406));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_jayjaywong12_8 (.L_LO(net8));
 sg13g2_tielo tt_um_jayjaywong12_9 (.L_LO(net9));
 sg13g2_tielo tt_um_jayjaywong12_10 (.L_LO(net10));
 sg13g2_tiehi _5489__11 (.L_HI(net11));
 sg13g2_buf_1 _6127_ (.A(read_operation),
    .X(uio_oe[0]));
 sg13g2_buf_1 _6128_ (.A(read_operation),
    .X(uio_oe[1]));
 sg13g2_buf_1 _6129_ (.A(read_operation),
    .X(uio_oe[2]));
 sg13g2_buf_1 _6130_ (.A(read_operation),
    .X(uio_oe[3]));
 sg13g2_buf_2 fanout441 (.A(net442),
    .X(net441));
 sg13g2_buf_4 fanout442 (.X(net442),
    .A(net443));
 sg13g2_buf_2 fanout443 (.A(net450),
    .X(net443));
 sg13g2_buf_4 fanout444 (.X(net444),
    .A(net445));
 sg13g2_buf_4 fanout445 (.X(net445),
    .A(net446));
 sg13g2_buf_2 fanout446 (.A(net450),
    .X(net446));
 sg13g2_buf_4 fanout447 (.X(net447),
    .A(net450));
 sg13g2_buf_4 fanout448 (.X(net448),
    .A(net450));
 sg13g2_buf_4 fanout449 (.X(net449),
    .A(net450));
 sg13g2_buf_4 fanout450 (.X(net450),
    .A(_0755_));
 sg13g2_buf_4 fanout451 (.X(net451),
    .A(net452));
 sg13g2_buf_4 fanout452 (.X(net452),
    .A(net456));
 sg13g2_buf_4 fanout453 (.X(net453),
    .A(net455));
 sg13g2_buf_4 fanout454 (.X(net454),
    .A(net455));
 sg13g2_buf_4 fanout455 (.X(net455),
    .A(net456));
 sg13g2_buf_2 fanout456 (.A(net460),
    .X(net456));
 sg13g2_buf_4 fanout457 (.X(net457),
    .A(net460));
 sg13g2_buf_2 fanout458 (.A(net459),
    .X(net458));
 sg13g2_buf_4 fanout459 (.X(net459),
    .A(net460));
 sg13g2_buf_2 fanout460 (.A(_0687_),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(net462),
    .X(net461));
 sg13g2_buf_4 fanout462 (.X(net462),
    .A(net471));
 sg13g2_buf_4 fanout463 (.X(net463),
    .A(net466));
 sg13g2_buf_2 fanout464 (.A(net466),
    .X(net464));
 sg13g2_buf_4 fanout465 (.X(net465),
    .A(net466));
 sg13g2_buf_2 fanout466 (.A(net471),
    .X(net466));
 sg13g2_buf_4 fanout467 (.X(net467),
    .A(net470));
 sg13g2_buf_2 fanout468 (.A(net470),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(net470),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(net471),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(_0623_),
    .X(net471));
 sg13g2_buf_4 fanout472 (.X(net472),
    .A(net474));
 sg13g2_buf_1 fanout473 (.A(net474),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(net482),
    .X(net474));
 sg13g2_buf_4 fanout475 (.X(net475),
    .A(net478));
 sg13g2_buf_2 fanout476 (.A(net478),
    .X(net476));
 sg13g2_buf_4 fanout477 (.X(net477),
    .A(net478));
 sg13g2_buf_2 fanout478 (.A(net482),
    .X(net478));
 sg13g2_buf_4 fanout479 (.X(net479),
    .A(net482));
 sg13g2_buf_2 fanout480 (.A(net481),
    .X(net480));
 sg13g2_buf_4 fanout481 (.X(net481),
    .A(net482));
 sg13g2_buf_4 fanout482 (.X(net482),
    .A(_0571_));
 sg13g2_buf_2 fanout483 (.A(_1190_),
    .X(net483));
 sg13g2_buf_4 fanout484 (.X(net484),
    .A(net485));
 sg13g2_buf_2 fanout485 (.A(net486),
    .X(net485));
 sg13g2_buf_4 fanout486 (.X(net486),
    .A(_0782_));
 sg13g2_buf_2 fanout487 (.A(net488),
    .X(net487));
 sg13g2_buf_4 fanout488 (.X(net488),
    .A(_0533_));
 sg13g2_buf_2 fanout489 (.A(_0780_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(net412),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(net844),
    .X(net491));
 sg13g2_buf_4 fanout492 (.X(net492),
    .A(net411));
 sg13g2_buf_2 fanout493 (.A(net851),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(net820),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(net409),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(net847),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(net424),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(net658),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(net635),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(net825),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(net784),
    .X(net501));
 sg13g2_buf_4 fanout502 (.X(net502),
    .A(net503));
 sg13g2_buf_2 fanout503 (.A(net504),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(_2095_),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(net509),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(net507),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(net508),
    .X(net507));
 sg13g2_buf_1 fanout508 (.A(net509),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(_2094_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(net511),
    .X(net510));
 sg13g2_buf_4 fanout511 (.X(net511),
    .A(_2094_));
 sg13g2_buf_2 fanout512 (.A(net513),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(_2094_),
    .X(net513));
 sg13g2_buf_4 fanout514 (.X(net514),
    .A(_2093_));
 sg13g2_buf_2 fanout515 (.A(net516),
    .X(net515));
 sg13g2_buf_4 fanout516 (.X(net516),
    .A(net517));
 sg13g2_buf_2 fanout517 (.A(net521),
    .X(net517));
 sg13g2_buf_4 fanout518 (.X(net518),
    .A(net521));
 sg13g2_buf_2 fanout519 (.A(net520),
    .X(net519));
 sg13g2_buf_4 fanout520 (.X(net520),
    .A(net521));
 sg13g2_buf_4 fanout521 (.X(net521),
    .A(_2092_));
 sg13g2_buf_2 fanout522 (.A(net523),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(ui_in[5]),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(net526),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(net526),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(ui_in[4]),
    .X(net526));
 sg13g2_buf_4 fanout527 (.X(net527),
    .A(ui_in[3]));
 sg13g2_buf_2 fanout528 (.A(ui_in[3]),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(net530),
    .X(net529));
 sg13g2_buf_4 fanout530 (.X(net530),
    .A(ui_in[3]));
 sg13g2_buf_4 fanout531 (.X(net531),
    .A(net532));
 sg13g2_buf_4 fanout532 (.X(net532),
    .A(ui_in[2]));
 sg13g2_buf_2 fanout533 (.A(net535),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(net535),
    .X(net534));
 sg13g2_buf_4 fanout535 (.X(net535),
    .A(net536));
 sg13g2_buf_4 fanout536 (.X(net536),
    .A(net550));
 sg13g2_buf_2 fanout537 (.A(net540),
    .X(net537));
 sg13g2_buf_1 fanout538 (.A(net540),
    .X(net538));
 sg13g2_buf_4 fanout539 (.X(net539),
    .A(net540));
 sg13g2_buf_2 fanout540 (.A(net550),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(net542),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(net550),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(net544),
    .X(net543));
 sg13g2_buf_1 fanout544 (.A(net545),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(net550),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(net547),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(net548),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(net549),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(net550),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(ui_in[1]),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(net552),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(net554),
    .X(net552));
 sg13g2_buf_4 fanout553 (.X(net553),
    .A(net554));
 sg13g2_buf_2 fanout554 (.A(net555),
    .X(net554));
 sg13g2_buf_4 fanout555 (.X(net555),
    .A(net577));
 sg13g2_buf_4 fanout556 (.X(net556),
    .A(net557));
 sg13g2_buf_2 fanout557 (.A(net563),
    .X(net557));
 sg13g2_buf_4 fanout558 (.X(net558),
    .A(net563));
 sg13g2_buf_1 fanout559 (.A(net563),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(net562),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(net562),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(net563),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(net577),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(net567),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(net566),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(net567),
    .X(net566));
 sg13g2_buf_1 fanout567 (.A(net568),
    .X(net567));
 sg13g2_buf_4 fanout568 (.X(net568),
    .A(net576));
 sg13g2_buf_2 fanout569 (.A(net573),
    .X(net569));
 sg13g2_buf_1 fanout570 (.A(net573),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(net573),
    .X(net571));
 sg13g2_buf_1 fanout572 (.A(net573),
    .X(net572));
 sg13g2_buf_1 fanout573 (.A(net574),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(net576),
    .X(net574));
 sg13g2_buf_4 fanout575 (.X(net575),
    .A(net576));
 sg13g2_buf_2 fanout576 (.A(net577),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(ui_in[0]),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(net580),
    .X(net578));
 sg13g2_buf_1 fanout579 (.A(net580),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(rst_n),
    .X(net580));
 sg13g2_buf_1 input1 (.A(ui_in[6]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[7]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(uio_in[0]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(uio_in[1]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(uio_in[2]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(uio_in[3]),
    .X(net6));
 sg13g2_tielo tt_um_jayjaywong12_7 (.L_LO(net7));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_4_5_0_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_4_7_0_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_4_9_0_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_4_11_0_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_4_13_0_clk));
 sg13g2_buf_2 clkload6 (.A(clknet_4_15_0_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_4_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_56_clk));
 sg13g2_inv_2 clkload9 (.A(clknet_leaf_7_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_8_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_53_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_55_clk));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_52_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_10_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_11_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_23_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_47_clk));
 sg13g2_inv_4 clkload18 (.A(clknet_leaf_49_clk));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_38_clk));
 sg13g2_inv_2 clkload20 (.A(clknet_leaf_42_clk));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_43_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_45_clk));
 sg13g2_inv_1 clkload23 (.A(clknet_leaf_39_clk));
 sg13g2_inv_1 clkload24 (.A(clknet_leaf_40_clk));
 sg13g2_inv_2 clkload25 (.A(clknet_leaf_24_clk));
 sg13g2_inv_4 clkload26 (.A(clknet_leaf_28_clk));
 sg13g2_inv_4 clkload27 (.A(clknet_leaf_35_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0000_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0337_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold3 (.A(\mem[5][0] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0354_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold5 (.A(\mem[0][3] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold6 (.A(\mem[8][1] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold7 (.A(_1667_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold8 (.A(\mem[38][3] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold9 (.A(\mem[54][0] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold10 (.A(\mem[38][1] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold11 (.A(\mem[46][0] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold12 (.A(\mem[39][3] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold13 (.A(\mem[42][3] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold14 (.A(\mem[38][2] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold15 (.A(\mem[54][3] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold16 (.A(\mem[46][3] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold17 (.A(\mem[57][1] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold18 (.A(\mem[14][0] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold19 (.A(_1312_),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold20 (.A(\mem[39][0] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold21 (.A(\mem[35][0] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold22 (.A(\mem[50][0] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold23 (.A(\mem[42][1] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold24 (.A(\mem[44][0] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold25 (.A(\mem[39][2] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold26 (.A(\mem[42][0] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold27 (.A(\mem[46][1] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold28 (.A(\mem[52][0] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold29 (.A(\mem[56][1] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold30 (.A(\mem[43][0] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold31 (.A(\mem[43][3] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold32 (.A(\mem[50][3] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold33 (.A(\mem[47][1] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold34 (.A(\mem[50][1] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold35 (.A(\mem[57][0] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold36 (.A(\mem[39][1] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold37 (.A(\mem[54][1] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold38 (.A(\mem[54][2] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold39 (.A(\mem[45][1] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold40 (.A(\mem[48][2] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold41 (.A(\mem[43][2] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold42 (.A(\mem[52][2] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold43 (.A(\mem[50][2] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold44 (.A(\mem[52][3] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold45 (.A(\mem[36][0] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold46 (.A(\mem[45][0] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold47 (.A(\mem[44][1] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold48 (.A(\mem[47][3] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold49 (.A(\mem[47][2] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold50 (.A(\mem[48][1] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold51 (.A(\mem[47][0] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold52 (.A(\mem[45][3] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold53 (.A(\mem[42][2] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold54 (.A(\mem[35][1] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold55 (.A(\mem[41][3] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold56 (.A(\mem[36][1] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold57 (.A(\mem[44][2] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold58 (.A(\mem[43][1] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold59 (.A(\mem[57][3] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold60 (.A(\mem[56][2] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold61 (.A(\mem[37][3] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold62 (.A(\mem[49][0] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold63 (.A(\mem[36][2] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold64 (.A(\mem[38][0] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold65 (.A(\mem[56][3] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold66 (.A(\mem[44][3] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold67 (.A(\mem[40][2] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold68 (.A(\mem[48][3] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold69 (.A(\mem[56][0] ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold70 (.A(\mem[35][3] ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold71 (.A(\mem[36][3] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold72 (.A(\mem[49][1] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold73 (.A(\mem[48][0] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold74 (.A(\mem[46][2] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold75 (.A(\mem[45][2] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold76 (.A(\mem[41][1] ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold77 (.A(\mem[41][0] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold78 (.A(\mem[40][1] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold79 (.A(\mem[57][2] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold80 (.A(\mem[35][2] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold81 (.A(\mem[37][0] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold82 (.A(\mem[37][2] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold83 (.A(\mem[49][2] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold84 (.A(\mem[41][2] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold85 (.A(\mem[40][3] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold86 (.A(\mem[52][1] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold87 (.A(\mem[49][3] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold88 (.A(\mem[62][3] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold89 (.A(\mem[15][0] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold90 (.A(\mem[63][2] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold91 (.A(\mem[58][0] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold92 (.A(\mem[63][1] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold93 (.A(\mem[40][0] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold94 (.A(\mem[51][2] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold95 (.A(\mem[59][1] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold96 (.A(\mem[59][2] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold97 (.A(\mem[53][0] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold98 (.A(\mem[51][3] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold99 (.A(\mem[58][1] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold100 (.A(\mem[61][0] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold101 (.A(\mem[58][3] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold102 (.A(\mem[62][2] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold103 (.A(\mem[37][1] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold104 (.A(\mem[62][1] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold105 (.A(\mem[59][3] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold106 (.A(\mem[60][2] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold107 (.A(\mem[63][3] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold108 (.A(\mem[53][3] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold109 (.A(\mem[53][2] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold110 (.A(\mem[55][1] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold111 (.A(\mem[53][1] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold112 (.A(\mem[15][1] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold113 (.A(\mem[55][2] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold114 (.A(\mem[58][2] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold115 (.A(\mem[51][0] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold116 (.A(\mem[61][1] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold117 (.A(\mem[62][0] ),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold118 (.A(\mem[63][0] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold119 (.A(\mem[60][3] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold120 (.A(\mem[55][3] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold121 (.A(\mem[61][3] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold122 (.A(\mem[60][0] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold123 (.A(\mem[51][1] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold124 (.A(\mem[55][0] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold125 (.A(\mem[60][1] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold126 (.A(\mem[61][2] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold127 (.A(\mem[59][0] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold128 (.A(\mem[12][0] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0298_),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold130 (.A(\mem[3][0] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold131 (.A(_1958_),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold132 (.A(\prev_acc[0] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0387_),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold134 (.A(\mem[4][0] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold135 (.A(_1899_),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold136 (.A(\prev_acc[1] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0388_),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold138 (.A(\mem[2][0] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0378_),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold140 (.A(\prev_acc[6] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0393_),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold142 (.A(\mem[20][1] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold143 (.A(_1901_),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold144 (.A(\mem[31][0] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold145 (.A(uo_out[2]),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0389_),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold147 (.A(uo_out[3]),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0390_),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold149 (.A(\prev_acc[7] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0394_),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold151 (.A(\mem[9][0] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0322_),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold153 (.A(\mem[28][0] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold154 (.A(_1430_),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold155 (.A(\mem[19][1] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold156 (.A(_1959_),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold157 (.A(uo_out[5]),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0054_),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold159 (.A(\mem[24][0] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0330_),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold161 (.A(\mem[7][0] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0338_),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold163 (.A(\prev_acc[4] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0391_),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold165 (.A(uo_out[0]),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold166 (.A(\mem[8][3] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold167 (.A(\mem[17][0] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0783_),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold169 (.A(\prev_acc[5] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold170 (.A(\mem[29][0] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0290_),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold172 (.A(\mem[25][3] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold173 (.A(\mem[11][3] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold174 (.A(\mem[9][3] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold175 (.A(uo_out[1]),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold176 (.A(\mem[18][1] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold177 (.A(_2016_),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold178 (.A(\mem[2][3] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold179 (.A(\mem[6][0] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold180 (.A(_1789_),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold181 (.A(\mem[17][1] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0784_),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold183 (.A(\mem[28][3] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold184 (.A(\mem[10][0] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold185 (.A(_1549_),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold186 (.A(\mem[6][2] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold187 (.A(uio_out[4]),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold188 (.A(_2073_),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold189 (.A(\mem[30][0] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold190 (.A(\mem[16][3] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold191 (.A(\mem[27][0] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0306_),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold193 (.A(\mem[15][3] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold194 (.A(\mem[9][2] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold195 (.A(uo_out[6]),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold196 (.A(\mem[4][3] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold197 (.A(\mem[27][3] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold198 (.A(\mem[32][3] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold199 (.A(\mem[20][0] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold200 (.A(\mem[17][3] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold201 (.A(\mem[22][2] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold202 (.A(\mem[3][1] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold203 (.A(\mem[2][1] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold204 (.A(\mem[17][2] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold205 (.A(\mem[24][3] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold206 (.A(\mem[6][3] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold207 (.A(\mem[9][1] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold208 (.A(_1608_),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold209 (.A(\mem[3][3] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold210 (.A(\mem[7][3] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold211 (.A(\mem[1][1] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold212 (.A(\mem[23][3] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold213 (.A(\mem[1][3] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold214 (.A(\mem[26][3] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold215 (.A(\mem[11][2] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold216 (.A(\mem[6][1] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold217 (.A(\mem[7][1] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold218 (.A(_1730_),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold219 (.A(\mem[1][0] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold220 (.A(\mem[7][2] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold221 (.A(\mem[2][2] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold222 (.A(\mem[4][2] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold223 (.A(\mem[11][0] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold224 (.A(_1489_),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold225 (.A(\mem[0][1] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold226 (.A(uo_out[7]),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0056_),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold228 (.A(\mem[14][3] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold229 (.A(\mem[20][3] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold230 (.A(\mem[10][3] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold231 (.A(\mem[31][3] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold232 (.A(\mem[1][2] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold233 (.A(\mem[15][2] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold234 (.A(\mem[31][1] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold235 (.A(\mem[32][0] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold236 (.A(\mem[25][0] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold237 (.A(\mem[22][0] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold238 (.A(\mem[16][0] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold239 (.A(\mem[12][3] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold240 (.A(\mem[18][3] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold241 (.A(\mem[22][1] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold242 (.A(\mem[26][1] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold243 (.A(_1550_),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold244 (.A(\mem[12][1] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold245 (.A(\mem[7][1] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold246 (.A(\mem[24][1] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold247 (.A(\mem[26][2] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold248 (.A(\mem[13][0] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold249 (.A(_1375_),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold250 (.A(\mem[4][1] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold251 (.A(\mem[18][0] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold252 (.A(\mem[11][1] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold253 (.A(\mem[27][1] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold254 (.A(\mem[25][2] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold255 (.A(\mem[8][2] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold256 (.A(\mem[31][0] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold257 (.A(\mem[32][1] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold258 (.A(\mem[0][0] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold259 (.A(\mem[5][3] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold260 (.A(\mem[25][1] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold261 (.A(\mem[23][2] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold262 (.A(\mem[19][2] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold263 (.A(\mem[10][1] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold264 (.A(\mem[29][3] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold265 (.A(\mem[27][2] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold266 (.A(\mem[31][2] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold267 (.A(\mem[24][2] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold268 (.A(\mem[32][2] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold269 (.A(\mem[21][1] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold270 (.A(_1845_),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0355_),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold272 (.A(\mem[19][0] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold273 (.A(\mem[3][2] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold274 (.A(\mem[5][1] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold275 (.A(\mem[19][3] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold276 (.A(uo_out[4]),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold277 (.A(\mem[22][3] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold278 (.A(\mem[28][1] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold279 (.A(\mem[16][1] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold280 (.A(\mem[26][0] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold281 (.A(\mem[30][1] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold282 (.A(\mem[30][3] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold283 (.A(\mem[13][3] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold284 (.A(\mem[14][2] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold285 (.A(\mem[28][2] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold286 (.A(\mem[5][2] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold287 (.A(\mem[10][2] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold288 (.A(\mem[12][2] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold289 (.A(\mem[29][1] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold290 (.A(\mem[23][1] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold291 (.A(\mem[23][0] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold292 (.A(\mem[29][2] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold293 (.A(\mem[16][2] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold294 (.A(\mem[20][2] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold295 (.A(\mem[18][2] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold296 (.A(\mem[13][1] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold297 (.A(\mem[13][2] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold298 (.A(\mem[8][0] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold299 (.A(\mem[21][3] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold300 (.A(\mem[21][0] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold301 (.A(\mem[14][1] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold302 (.A(\mem[21][2] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold303 (.A(\mem[30][2] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold304 (.A(\mem[21][3] ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold305 (.A(\mem[0][2] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold306 (.A(\mem[30][3] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold307 (.A(\mem[12][1] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold308 (.A(uio_out[5]),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold309 (.A(\mem[6][2] ),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold310 (.A(\mem[3][0] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold311 (.A(_1963_),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0372_),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold313 (.A(\mem[7][0] ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold314 (.A(\mem[29][0] ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold315 (.A(\mem[12][2] ),
    .X(net861));
 sg13g2_antennanp ANTENNA_1 (.A(_0269_));
 sg13g2_antennanp ANTENNA_2 (.A(_0272_));
 sg13g2_antennanp ANTENNA_3 (.A(_0272_));
 sg13g2_antennanp ANTENNA_4 (.A(_0331_));
 sg13g2_antennanp ANTENNA_5 (.A(_0272_));
 sg13g2_antennanp ANTENNA_6 (.A(_0272_));
 sg13g2_antennanp ANTENNA_7 (.A(_0273_));
 sg13g2_antennanp ANTENNA_8 (.A(_0273_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_decap_8 FILLER_13_588 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_decap_8 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_637 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_8 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_decap_8 FILLER_13_798 ();
 sg13g2_decap_8 FILLER_13_805 ();
 sg13g2_decap_8 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_833 ();
 sg13g2_decap_8 FILLER_13_840 ();
 sg13g2_decap_8 FILLER_13_847 ();
 sg13g2_decap_8 FILLER_13_854 ();
 sg13g2_fill_1 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_8 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_511 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_574 ();
 sg13g2_decap_8 FILLER_14_581 ();
 sg13g2_decap_8 FILLER_14_588 ();
 sg13g2_decap_8 FILLER_14_595 ();
 sg13g2_decap_8 FILLER_14_602 ();
 sg13g2_decap_8 FILLER_14_609 ();
 sg13g2_decap_8 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_623 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_decap_8 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_decap_8 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_658 ();
 sg13g2_decap_8 FILLER_14_665 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_decap_8 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_decap_8 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_14_840 ();
 sg13g2_decap_8 FILLER_14_847 ();
 sg13g2_decap_8 FILLER_14_854 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_434 ();
 sg13g2_decap_8 FILLER_15_441 ();
 sg13g2_decap_8 FILLER_15_448 ();
 sg13g2_decap_8 FILLER_15_455 ();
 sg13g2_decap_8 FILLER_15_462 ();
 sg13g2_decap_8 FILLER_15_469 ();
 sg13g2_decap_8 FILLER_15_476 ();
 sg13g2_decap_8 FILLER_15_483 ();
 sg13g2_decap_8 FILLER_15_490 ();
 sg13g2_decap_8 FILLER_15_497 ();
 sg13g2_decap_8 FILLER_15_504 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_518 ();
 sg13g2_decap_8 FILLER_15_525 ();
 sg13g2_decap_8 FILLER_15_532 ();
 sg13g2_decap_8 FILLER_15_539 ();
 sg13g2_decap_8 FILLER_15_546 ();
 sg13g2_decap_8 FILLER_15_553 ();
 sg13g2_decap_8 FILLER_15_560 ();
 sg13g2_decap_8 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_574 ();
 sg13g2_decap_8 FILLER_15_581 ();
 sg13g2_decap_8 FILLER_15_588 ();
 sg13g2_decap_8 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_602 ();
 sg13g2_decap_8 FILLER_15_609 ();
 sg13g2_decap_8 FILLER_15_616 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_8 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_644 ();
 sg13g2_decap_8 FILLER_15_651 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_decap_8 FILLER_15_665 ();
 sg13g2_decap_8 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_679 ();
 sg13g2_decap_8 FILLER_15_686 ();
 sg13g2_decap_8 FILLER_15_693 ();
 sg13g2_decap_8 FILLER_15_700 ();
 sg13g2_decap_8 FILLER_15_707 ();
 sg13g2_decap_8 FILLER_15_714 ();
 sg13g2_decap_8 FILLER_15_721 ();
 sg13g2_decap_8 FILLER_15_728 ();
 sg13g2_decap_8 FILLER_15_735 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_decap_8 FILLER_15_749 ();
 sg13g2_decap_8 FILLER_15_756 ();
 sg13g2_decap_8 FILLER_15_763 ();
 sg13g2_decap_8 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_777 ();
 sg13g2_decap_8 FILLER_15_784 ();
 sg13g2_decap_8 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_798 ();
 sg13g2_decap_8 FILLER_15_805 ();
 sg13g2_decap_8 FILLER_15_812 ();
 sg13g2_decap_8 FILLER_15_819 ();
 sg13g2_decap_8 FILLER_15_826 ();
 sg13g2_decap_8 FILLER_15_833 ();
 sg13g2_decap_8 FILLER_15_840 ();
 sg13g2_decap_8 FILLER_15_847 ();
 sg13g2_decap_8 FILLER_15_854 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_8 FILLER_16_455 ();
 sg13g2_decap_8 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_469 ();
 sg13g2_decap_8 FILLER_16_476 ();
 sg13g2_decap_8 FILLER_16_483 ();
 sg13g2_decap_8 FILLER_16_490 ();
 sg13g2_decap_8 FILLER_16_497 ();
 sg13g2_decap_8 FILLER_16_504 ();
 sg13g2_decap_8 FILLER_16_511 ();
 sg13g2_decap_8 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_525 ();
 sg13g2_decap_8 FILLER_16_532 ();
 sg13g2_decap_8 FILLER_16_539 ();
 sg13g2_decap_8 FILLER_16_546 ();
 sg13g2_decap_8 FILLER_16_553 ();
 sg13g2_decap_8 FILLER_16_560 ();
 sg13g2_decap_8 FILLER_16_567 ();
 sg13g2_decap_8 FILLER_16_574 ();
 sg13g2_decap_8 FILLER_16_581 ();
 sg13g2_decap_8 FILLER_16_588 ();
 sg13g2_decap_8 FILLER_16_595 ();
 sg13g2_decap_8 FILLER_16_602 ();
 sg13g2_decap_8 FILLER_16_609 ();
 sg13g2_decap_8 FILLER_16_616 ();
 sg13g2_decap_8 FILLER_16_623 ();
 sg13g2_decap_8 FILLER_16_630 ();
 sg13g2_decap_8 FILLER_16_637 ();
 sg13g2_decap_8 FILLER_16_644 ();
 sg13g2_decap_8 FILLER_16_651 ();
 sg13g2_decap_8 FILLER_16_658 ();
 sg13g2_decap_8 FILLER_16_665 ();
 sg13g2_decap_8 FILLER_16_672 ();
 sg13g2_decap_8 FILLER_16_679 ();
 sg13g2_decap_8 FILLER_16_686 ();
 sg13g2_decap_8 FILLER_16_693 ();
 sg13g2_decap_8 FILLER_16_700 ();
 sg13g2_decap_8 FILLER_16_707 ();
 sg13g2_decap_8 FILLER_16_714 ();
 sg13g2_decap_8 FILLER_16_721 ();
 sg13g2_decap_8 FILLER_16_728 ();
 sg13g2_decap_8 FILLER_16_735 ();
 sg13g2_decap_8 FILLER_16_742 ();
 sg13g2_decap_8 FILLER_16_749 ();
 sg13g2_decap_8 FILLER_16_756 ();
 sg13g2_decap_8 FILLER_16_763 ();
 sg13g2_decap_8 FILLER_16_770 ();
 sg13g2_decap_8 FILLER_16_777 ();
 sg13g2_decap_8 FILLER_16_784 ();
 sg13g2_decap_8 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_798 ();
 sg13g2_decap_8 FILLER_16_805 ();
 sg13g2_decap_8 FILLER_16_812 ();
 sg13g2_decap_8 FILLER_16_819 ();
 sg13g2_decap_8 FILLER_16_826 ();
 sg13g2_decap_8 FILLER_16_833 ();
 sg13g2_decap_8 FILLER_16_840 ();
 sg13g2_decap_8 FILLER_16_847 ();
 sg13g2_decap_8 FILLER_16_854 ();
 sg13g2_fill_1 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_427 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_448 ();
 sg13g2_decap_8 FILLER_17_455 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_497 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_fill_1 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_decap_8 FILLER_18_427 ();
 sg13g2_decap_8 FILLER_18_434 ();
 sg13g2_decap_8 FILLER_18_441 ();
 sg13g2_decap_8 FILLER_18_448 ();
 sg13g2_decap_8 FILLER_18_455 ();
 sg13g2_decap_8 FILLER_18_462 ();
 sg13g2_decap_8 FILLER_18_469 ();
 sg13g2_decap_8 FILLER_18_476 ();
 sg13g2_decap_8 FILLER_18_483 ();
 sg13g2_decap_8 FILLER_18_490 ();
 sg13g2_decap_8 FILLER_18_497 ();
 sg13g2_decap_8 FILLER_18_504 ();
 sg13g2_decap_8 FILLER_18_511 ();
 sg13g2_decap_8 FILLER_18_518 ();
 sg13g2_decap_8 FILLER_18_525 ();
 sg13g2_decap_8 FILLER_18_532 ();
 sg13g2_decap_8 FILLER_18_539 ();
 sg13g2_decap_8 FILLER_18_546 ();
 sg13g2_decap_8 FILLER_18_553 ();
 sg13g2_decap_8 FILLER_18_560 ();
 sg13g2_decap_8 FILLER_18_567 ();
 sg13g2_decap_8 FILLER_18_574 ();
 sg13g2_decap_8 FILLER_18_581 ();
 sg13g2_decap_8 FILLER_18_588 ();
 sg13g2_decap_8 FILLER_18_595 ();
 sg13g2_decap_8 FILLER_18_602 ();
 sg13g2_decap_8 FILLER_18_609 ();
 sg13g2_decap_8 FILLER_18_616 ();
 sg13g2_decap_8 FILLER_18_623 ();
 sg13g2_decap_8 FILLER_18_630 ();
 sg13g2_decap_8 FILLER_18_637 ();
 sg13g2_decap_8 FILLER_18_644 ();
 sg13g2_decap_8 FILLER_18_651 ();
 sg13g2_decap_8 FILLER_18_658 ();
 sg13g2_decap_8 FILLER_18_665 ();
 sg13g2_decap_8 FILLER_18_672 ();
 sg13g2_decap_8 FILLER_18_679 ();
 sg13g2_decap_8 FILLER_18_686 ();
 sg13g2_decap_8 FILLER_18_693 ();
 sg13g2_decap_8 FILLER_18_700 ();
 sg13g2_decap_8 FILLER_18_707 ();
 sg13g2_decap_8 FILLER_18_714 ();
 sg13g2_decap_8 FILLER_18_721 ();
 sg13g2_decap_8 FILLER_18_728 ();
 sg13g2_decap_8 FILLER_18_735 ();
 sg13g2_decap_8 FILLER_18_742 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_decap_8 FILLER_18_756 ();
 sg13g2_decap_8 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_770 ();
 sg13g2_decap_8 FILLER_18_777 ();
 sg13g2_decap_8 FILLER_18_784 ();
 sg13g2_decap_8 FILLER_18_791 ();
 sg13g2_decap_8 FILLER_18_798 ();
 sg13g2_decap_8 FILLER_18_805 ();
 sg13g2_decap_8 FILLER_18_812 ();
 sg13g2_decap_8 FILLER_18_819 ();
 sg13g2_decap_8 FILLER_18_826 ();
 sg13g2_decap_8 FILLER_18_833 ();
 sg13g2_decap_8 FILLER_18_840 ();
 sg13g2_decap_8 FILLER_18_847 ();
 sg13g2_decap_8 FILLER_18_854 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_decap_8 FILLER_19_427 ();
 sg13g2_decap_8 FILLER_19_434 ();
 sg13g2_decap_8 FILLER_19_441 ();
 sg13g2_decap_8 FILLER_19_448 ();
 sg13g2_decap_8 FILLER_19_455 ();
 sg13g2_decap_8 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_490 ();
 sg13g2_decap_8 FILLER_19_497 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_532 ();
 sg13g2_decap_8 FILLER_19_539 ();
 sg13g2_decap_8 FILLER_19_546 ();
 sg13g2_decap_8 FILLER_19_553 ();
 sg13g2_decap_8 FILLER_19_560 ();
 sg13g2_decap_8 FILLER_19_567 ();
 sg13g2_decap_8 FILLER_19_574 ();
 sg13g2_decap_8 FILLER_19_581 ();
 sg13g2_decap_8 FILLER_19_588 ();
 sg13g2_decap_8 FILLER_19_595 ();
 sg13g2_decap_8 FILLER_19_602 ();
 sg13g2_decap_8 FILLER_19_609 ();
 sg13g2_decap_8 FILLER_19_616 ();
 sg13g2_decap_8 FILLER_19_623 ();
 sg13g2_decap_8 FILLER_19_630 ();
 sg13g2_decap_8 FILLER_19_637 ();
 sg13g2_decap_8 FILLER_19_644 ();
 sg13g2_decap_8 FILLER_19_651 ();
 sg13g2_decap_8 FILLER_19_658 ();
 sg13g2_decap_8 FILLER_19_665 ();
 sg13g2_decap_8 FILLER_19_672 ();
 sg13g2_decap_8 FILLER_19_679 ();
 sg13g2_decap_8 FILLER_19_686 ();
 sg13g2_decap_8 FILLER_19_693 ();
 sg13g2_decap_8 FILLER_19_700 ();
 sg13g2_decap_8 FILLER_19_707 ();
 sg13g2_decap_8 FILLER_19_714 ();
 sg13g2_decap_8 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_784 ();
 sg13g2_decap_8 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_798 ();
 sg13g2_decap_8 FILLER_19_805 ();
 sg13g2_decap_8 FILLER_19_812 ();
 sg13g2_decap_8 FILLER_19_819 ();
 sg13g2_decap_8 FILLER_19_826 ();
 sg13g2_decap_8 FILLER_19_833 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_decap_8 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_854 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_decap_8 FILLER_20_427 ();
 sg13g2_decap_8 FILLER_20_434 ();
 sg13g2_decap_8 FILLER_20_441 ();
 sg13g2_decap_8 FILLER_20_448 ();
 sg13g2_decap_8 FILLER_20_455 ();
 sg13g2_decap_8 FILLER_20_462 ();
 sg13g2_decap_8 FILLER_20_469 ();
 sg13g2_decap_8 FILLER_20_476 ();
 sg13g2_decap_8 FILLER_20_483 ();
 sg13g2_decap_8 FILLER_20_490 ();
 sg13g2_decap_8 FILLER_20_497 ();
 sg13g2_decap_8 FILLER_20_504 ();
 sg13g2_decap_8 FILLER_20_511 ();
 sg13g2_decap_8 FILLER_20_518 ();
 sg13g2_decap_8 FILLER_20_525 ();
 sg13g2_decap_8 FILLER_20_532 ();
 sg13g2_decap_8 FILLER_20_539 ();
 sg13g2_decap_8 FILLER_20_546 ();
 sg13g2_decap_8 FILLER_20_553 ();
 sg13g2_decap_8 FILLER_20_560 ();
 sg13g2_decap_8 FILLER_20_567 ();
 sg13g2_decap_8 FILLER_20_574 ();
 sg13g2_decap_8 FILLER_20_581 ();
 sg13g2_decap_8 FILLER_20_588 ();
 sg13g2_decap_8 FILLER_20_595 ();
 sg13g2_decap_8 FILLER_20_602 ();
 sg13g2_decap_8 FILLER_20_609 ();
 sg13g2_decap_8 FILLER_20_616 ();
 sg13g2_decap_8 FILLER_20_623 ();
 sg13g2_decap_8 FILLER_20_630 ();
 sg13g2_decap_8 FILLER_20_637 ();
 sg13g2_decap_8 FILLER_20_644 ();
 sg13g2_decap_8 FILLER_20_651 ();
 sg13g2_decap_8 FILLER_20_658 ();
 sg13g2_decap_8 FILLER_20_665 ();
 sg13g2_decap_8 FILLER_20_672 ();
 sg13g2_decap_8 FILLER_20_679 ();
 sg13g2_decap_8 FILLER_20_686 ();
 sg13g2_decap_8 FILLER_20_693 ();
 sg13g2_decap_8 FILLER_20_700 ();
 sg13g2_decap_8 FILLER_20_707 ();
 sg13g2_decap_8 FILLER_20_714 ();
 sg13g2_decap_8 FILLER_20_721 ();
 sg13g2_decap_8 FILLER_20_728 ();
 sg13g2_decap_8 FILLER_20_735 ();
 sg13g2_decap_8 FILLER_20_742 ();
 sg13g2_decap_8 FILLER_20_749 ();
 sg13g2_decap_8 FILLER_20_756 ();
 sg13g2_decap_8 FILLER_20_763 ();
 sg13g2_decap_8 FILLER_20_770 ();
 sg13g2_decap_8 FILLER_20_777 ();
 sg13g2_decap_8 FILLER_20_784 ();
 sg13g2_decap_8 FILLER_20_791 ();
 sg13g2_decap_8 FILLER_20_798 ();
 sg13g2_decap_8 FILLER_20_805 ();
 sg13g2_decap_8 FILLER_20_812 ();
 sg13g2_decap_8 FILLER_20_819 ();
 sg13g2_decap_8 FILLER_20_826 ();
 sg13g2_decap_8 FILLER_20_833 ();
 sg13g2_decap_8 FILLER_20_840 ();
 sg13g2_decap_8 FILLER_20_847 ();
 sg13g2_decap_8 FILLER_20_854 ();
 sg13g2_fill_1 FILLER_20_861 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_decap_8 FILLER_21_427 ();
 sg13g2_decap_8 FILLER_21_434 ();
 sg13g2_decap_8 FILLER_21_441 ();
 sg13g2_decap_8 FILLER_21_448 ();
 sg13g2_decap_8 FILLER_21_455 ();
 sg13g2_decap_8 FILLER_21_462 ();
 sg13g2_decap_8 FILLER_21_469 ();
 sg13g2_decap_8 FILLER_21_476 ();
 sg13g2_decap_8 FILLER_21_483 ();
 sg13g2_decap_8 FILLER_21_490 ();
 sg13g2_decap_8 FILLER_21_497 ();
 sg13g2_decap_8 FILLER_21_504 ();
 sg13g2_decap_8 FILLER_21_511 ();
 sg13g2_decap_8 FILLER_21_518 ();
 sg13g2_decap_8 FILLER_21_525 ();
 sg13g2_decap_8 FILLER_21_532 ();
 sg13g2_decap_8 FILLER_21_539 ();
 sg13g2_decap_8 FILLER_21_546 ();
 sg13g2_decap_8 FILLER_21_553 ();
 sg13g2_decap_8 FILLER_21_560 ();
 sg13g2_decap_8 FILLER_21_567 ();
 sg13g2_decap_8 FILLER_21_574 ();
 sg13g2_decap_8 FILLER_21_581 ();
 sg13g2_decap_8 FILLER_21_588 ();
 sg13g2_decap_8 FILLER_21_595 ();
 sg13g2_decap_8 FILLER_21_602 ();
 sg13g2_decap_8 FILLER_21_609 ();
 sg13g2_decap_8 FILLER_21_616 ();
 sg13g2_decap_8 FILLER_21_623 ();
 sg13g2_decap_8 FILLER_21_630 ();
 sg13g2_decap_8 FILLER_21_637 ();
 sg13g2_decap_8 FILLER_21_644 ();
 sg13g2_decap_8 FILLER_21_651 ();
 sg13g2_decap_8 FILLER_21_658 ();
 sg13g2_decap_8 FILLER_21_665 ();
 sg13g2_decap_8 FILLER_21_672 ();
 sg13g2_decap_8 FILLER_21_679 ();
 sg13g2_decap_8 FILLER_21_686 ();
 sg13g2_decap_8 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_700 ();
 sg13g2_decap_8 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_714 ();
 sg13g2_decap_8 FILLER_21_721 ();
 sg13g2_decap_8 FILLER_21_728 ();
 sg13g2_decap_8 FILLER_21_735 ();
 sg13g2_decap_8 FILLER_21_742 ();
 sg13g2_decap_8 FILLER_21_749 ();
 sg13g2_decap_8 FILLER_21_756 ();
 sg13g2_decap_8 FILLER_21_763 ();
 sg13g2_decap_8 FILLER_21_770 ();
 sg13g2_decap_8 FILLER_21_777 ();
 sg13g2_decap_8 FILLER_21_784 ();
 sg13g2_decap_8 FILLER_21_791 ();
 sg13g2_decap_8 FILLER_21_798 ();
 sg13g2_decap_8 FILLER_21_805 ();
 sg13g2_decap_8 FILLER_21_812 ();
 sg13g2_decap_8 FILLER_21_819 ();
 sg13g2_decap_8 FILLER_21_826 ();
 sg13g2_decap_8 FILLER_21_833 ();
 sg13g2_decap_8 FILLER_21_840 ();
 sg13g2_decap_8 FILLER_21_847 ();
 sg13g2_decap_8 FILLER_21_854 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_22_406 ();
 sg13g2_decap_8 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_decap_8 FILLER_22_427 ();
 sg13g2_decap_8 FILLER_22_434 ();
 sg13g2_decap_8 FILLER_22_441 ();
 sg13g2_decap_8 FILLER_22_448 ();
 sg13g2_decap_8 FILLER_22_455 ();
 sg13g2_decap_8 FILLER_22_462 ();
 sg13g2_decap_8 FILLER_22_469 ();
 sg13g2_decap_8 FILLER_22_476 ();
 sg13g2_decap_8 FILLER_22_483 ();
 sg13g2_fill_2 FILLER_22_490 ();
 sg13g2_decap_8 FILLER_22_518 ();
 sg13g2_decap_8 FILLER_22_525 ();
 sg13g2_decap_8 FILLER_22_532 ();
 sg13g2_decap_8 FILLER_22_539 ();
 sg13g2_decap_8 FILLER_22_546 ();
 sg13g2_decap_8 FILLER_22_553 ();
 sg13g2_decap_8 FILLER_22_560 ();
 sg13g2_decap_8 FILLER_22_567 ();
 sg13g2_decap_8 FILLER_22_574 ();
 sg13g2_decap_8 FILLER_22_581 ();
 sg13g2_decap_8 FILLER_22_588 ();
 sg13g2_decap_8 FILLER_22_595 ();
 sg13g2_decap_8 FILLER_22_602 ();
 sg13g2_decap_8 FILLER_22_609 ();
 sg13g2_decap_8 FILLER_22_616 ();
 sg13g2_decap_8 FILLER_22_623 ();
 sg13g2_decap_8 FILLER_22_630 ();
 sg13g2_decap_8 FILLER_22_637 ();
 sg13g2_decap_8 FILLER_22_644 ();
 sg13g2_decap_8 FILLER_22_651 ();
 sg13g2_decap_8 FILLER_22_658 ();
 sg13g2_decap_8 FILLER_22_665 ();
 sg13g2_decap_8 FILLER_22_672 ();
 sg13g2_decap_8 FILLER_22_679 ();
 sg13g2_decap_8 FILLER_22_686 ();
 sg13g2_decap_8 FILLER_22_693 ();
 sg13g2_decap_8 FILLER_22_700 ();
 sg13g2_decap_8 FILLER_22_707 ();
 sg13g2_decap_8 FILLER_22_714 ();
 sg13g2_decap_8 FILLER_22_721 ();
 sg13g2_decap_8 FILLER_22_728 ();
 sg13g2_decap_8 FILLER_22_735 ();
 sg13g2_decap_8 FILLER_22_742 ();
 sg13g2_decap_8 FILLER_22_749 ();
 sg13g2_decap_8 FILLER_22_756 ();
 sg13g2_decap_8 FILLER_22_763 ();
 sg13g2_decap_8 FILLER_22_770 ();
 sg13g2_decap_8 FILLER_22_777 ();
 sg13g2_decap_8 FILLER_22_784 ();
 sg13g2_decap_8 FILLER_22_791 ();
 sg13g2_decap_8 FILLER_22_798 ();
 sg13g2_decap_8 FILLER_22_805 ();
 sg13g2_decap_8 FILLER_22_812 ();
 sg13g2_decap_8 FILLER_22_819 ();
 sg13g2_decap_8 FILLER_22_826 ();
 sg13g2_decap_8 FILLER_22_833 ();
 sg13g2_decap_8 FILLER_22_840 ();
 sg13g2_decap_8 FILLER_22_847 ();
 sg13g2_decap_8 FILLER_22_854 ();
 sg13g2_fill_1 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_4 FILLER_23_385 ();
 sg13g2_fill_2 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_decap_4 FILLER_23_408 ();
 sg13g2_fill_1 FILLER_23_412 ();
 sg13g2_decap_4 FILLER_23_423 ();
 sg13g2_fill_2 FILLER_23_427 ();
 sg13g2_decap_8 FILLER_23_442 ();
 sg13g2_fill_2 FILLER_23_449 ();
 sg13g2_fill_1 FILLER_23_451 ();
 sg13g2_fill_2 FILLER_23_456 ();
 sg13g2_fill_2 FILLER_23_474 ();
 sg13g2_fill_1 FILLER_23_476 ();
 sg13g2_fill_1 FILLER_23_512 ();
 sg13g2_decap_8 FILLER_23_539 ();
 sg13g2_decap_8 FILLER_23_546 ();
 sg13g2_decap_8 FILLER_23_553 ();
 sg13g2_decap_8 FILLER_23_560 ();
 sg13g2_decap_8 FILLER_23_567 ();
 sg13g2_decap_8 FILLER_23_574 ();
 sg13g2_decap_8 FILLER_23_581 ();
 sg13g2_decap_8 FILLER_23_588 ();
 sg13g2_decap_8 FILLER_23_595 ();
 sg13g2_decap_8 FILLER_23_602 ();
 sg13g2_decap_8 FILLER_23_609 ();
 sg13g2_decap_8 FILLER_23_616 ();
 sg13g2_decap_8 FILLER_23_623 ();
 sg13g2_decap_8 FILLER_23_630 ();
 sg13g2_decap_8 FILLER_23_637 ();
 sg13g2_decap_8 FILLER_23_644 ();
 sg13g2_decap_8 FILLER_23_651 ();
 sg13g2_decap_8 FILLER_23_658 ();
 sg13g2_decap_8 FILLER_23_665 ();
 sg13g2_decap_8 FILLER_23_672 ();
 sg13g2_decap_8 FILLER_23_679 ();
 sg13g2_decap_8 FILLER_23_686 ();
 sg13g2_decap_8 FILLER_23_693 ();
 sg13g2_decap_8 FILLER_23_700 ();
 sg13g2_decap_8 FILLER_23_707 ();
 sg13g2_decap_8 FILLER_23_714 ();
 sg13g2_decap_8 FILLER_23_721 ();
 sg13g2_decap_8 FILLER_23_728 ();
 sg13g2_decap_8 FILLER_23_735 ();
 sg13g2_decap_8 FILLER_23_742 ();
 sg13g2_decap_8 FILLER_23_749 ();
 sg13g2_decap_8 FILLER_23_756 ();
 sg13g2_decap_8 FILLER_23_763 ();
 sg13g2_decap_8 FILLER_23_770 ();
 sg13g2_decap_8 FILLER_23_777 ();
 sg13g2_decap_8 FILLER_23_784 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_798 ();
 sg13g2_decap_8 FILLER_23_805 ();
 sg13g2_decap_8 FILLER_23_812 ();
 sg13g2_decap_8 FILLER_23_819 ();
 sg13g2_decap_8 FILLER_23_826 ();
 sg13g2_decap_8 FILLER_23_833 ();
 sg13g2_decap_8 FILLER_23_840 ();
 sg13g2_decap_8 FILLER_23_847 ();
 sg13g2_decap_8 FILLER_23_854 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_4 FILLER_24_259 ();
 sg13g2_fill_2 FILLER_24_263 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_4 FILLER_24_357 ();
 sg13g2_fill_2 FILLER_24_387 ();
 sg13g2_decap_4 FILLER_24_467 ();
 sg13g2_fill_2 FILLER_24_518 ();
 sg13g2_fill_1 FILLER_24_520 ();
 sg13g2_fill_2 FILLER_24_534 ();
 sg13g2_fill_1 FILLER_24_536 ();
 sg13g2_decap_8 FILLER_24_549 ();
 sg13g2_fill_1 FILLER_24_556 ();
 sg13g2_decap_8 FILLER_24_562 ();
 sg13g2_fill_2 FILLER_24_569 ();
 sg13g2_fill_1 FILLER_24_571 ();
 sg13g2_decap_8 FILLER_24_598 ();
 sg13g2_decap_8 FILLER_24_605 ();
 sg13g2_decap_8 FILLER_24_612 ();
 sg13g2_decap_8 FILLER_24_619 ();
 sg13g2_decap_8 FILLER_24_652 ();
 sg13g2_decap_8 FILLER_24_659 ();
 sg13g2_decap_8 FILLER_24_666 ();
 sg13g2_decap_8 FILLER_24_673 ();
 sg13g2_decap_8 FILLER_24_680 ();
 sg13g2_decap_8 FILLER_24_687 ();
 sg13g2_decap_8 FILLER_24_694 ();
 sg13g2_decap_8 FILLER_24_701 ();
 sg13g2_decap_8 FILLER_24_708 ();
 sg13g2_decap_8 FILLER_24_715 ();
 sg13g2_decap_8 FILLER_24_722 ();
 sg13g2_decap_8 FILLER_24_729 ();
 sg13g2_decap_8 FILLER_24_736 ();
 sg13g2_decap_8 FILLER_24_743 ();
 sg13g2_decap_8 FILLER_24_750 ();
 sg13g2_decap_8 FILLER_24_757 ();
 sg13g2_decap_8 FILLER_24_764 ();
 sg13g2_decap_8 FILLER_24_771 ();
 sg13g2_decap_8 FILLER_24_778 ();
 sg13g2_decap_8 FILLER_24_785 ();
 sg13g2_decap_8 FILLER_24_792 ();
 sg13g2_decap_8 FILLER_24_799 ();
 sg13g2_decap_8 FILLER_24_806 ();
 sg13g2_decap_8 FILLER_24_813 ();
 sg13g2_decap_8 FILLER_24_820 ();
 sg13g2_decap_8 FILLER_24_827 ();
 sg13g2_decap_8 FILLER_24_834 ();
 sg13g2_decap_8 FILLER_24_841 ();
 sg13g2_decap_8 FILLER_24_848 ();
 sg13g2_decap_8 FILLER_24_855 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_4 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_232 ();
 sg13g2_decap_4 FILLER_25_239 ();
 sg13g2_fill_1 FILLER_25_243 ();
 sg13g2_decap_4 FILLER_25_296 ();
 sg13g2_fill_1 FILLER_25_300 ();
 sg13g2_decap_8 FILLER_25_305 ();
 sg13g2_decap_4 FILLER_25_312 ();
 sg13g2_decap_8 FILLER_25_324 ();
 sg13g2_decap_8 FILLER_25_331 ();
 sg13g2_decap_4 FILLER_25_338 ();
 sg13g2_fill_2 FILLER_25_342 ();
 sg13g2_decap_4 FILLER_25_352 ();
 sg13g2_fill_1 FILLER_25_356 ();
 sg13g2_decap_4 FILLER_25_361 ();
 sg13g2_fill_2 FILLER_25_365 ();
 sg13g2_decap_8 FILLER_25_387 ();
 sg13g2_decap_8 FILLER_25_394 ();
 sg13g2_fill_2 FILLER_25_414 ();
 sg13g2_fill_2 FILLER_25_433 ();
 sg13g2_fill_1 FILLER_25_435 ();
 sg13g2_fill_1 FILLER_25_453 ();
 sg13g2_fill_2 FILLER_25_462 ();
 sg13g2_decap_8 FILLER_25_477 ();
 sg13g2_decap_8 FILLER_25_484 ();
 sg13g2_fill_2 FILLER_25_491 ();
 sg13g2_fill_1 FILLER_25_493 ();
 sg13g2_fill_2 FILLER_25_544 ();
 sg13g2_fill_1 FILLER_25_546 ();
 sg13g2_fill_1 FILLER_25_570 ();
 sg13g2_fill_2 FILLER_25_589 ();
 sg13g2_fill_1 FILLER_25_591 ();
 sg13g2_decap_8 FILLER_25_608 ();
 sg13g2_fill_1 FILLER_25_615 ();
 sg13g2_decap_8 FILLER_25_620 ();
 sg13g2_decap_8 FILLER_25_627 ();
 sg13g2_decap_4 FILLER_25_634 ();
 sg13g2_decap_8 FILLER_25_646 ();
 sg13g2_decap_8 FILLER_25_658 ();
 sg13g2_decap_8 FILLER_25_665 ();
 sg13g2_decap_8 FILLER_25_672 ();
 sg13g2_decap_8 FILLER_25_679 ();
 sg13g2_decap_8 FILLER_25_686 ();
 sg13g2_decap_8 FILLER_25_693 ();
 sg13g2_decap_8 FILLER_25_700 ();
 sg13g2_decap_8 FILLER_25_707 ();
 sg13g2_decap_8 FILLER_25_714 ();
 sg13g2_decap_8 FILLER_25_721 ();
 sg13g2_decap_8 FILLER_25_728 ();
 sg13g2_decap_8 FILLER_25_735 ();
 sg13g2_decap_8 FILLER_25_742 ();
 sg13g2_decap_8 FILLER_25_749 ();
 sg13g2_decap_8 FILLER_25_756 ();
 sg13g2_decap_8 FILLER_25_763 ();
 sg13g2_decap_8 FILLER_25_770 ();
 sg13g2_decap_8 FILLER_25_777 ();
 sg13g2_decap_8 FILLER_25_784 ();
 sg13g2_decap_8 FILLER_25_791 ();
 sg13g2_decap_8 FILLER_25_798 ();
 sg13g2_decap_8 FILLER_25_805 ();
 sg13g2_decap_8 FILLER_25_812 ();
 sg13g2_decap_8 FILLER_25_819 ();
 sg13g2_decap_8 FILLER_25_826 ();
 sg13g2_decap_8 FILLER_25_833 ();
 sg13g2_decap_8 FILLER_25_840 ();
 sg13g2_decap_8 FILLER_25_847 ();
 sg13g2_decap_8 FILLER_25_854 ();
 sg13g2_fill_1 FILLER_25_861 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_fill_2 FILLER_26_210 ();
 sg13g2_fill_1 FILLER_26_212 ();
 sg13g2_fill_1 FILLER_26_261 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_fill_1 FILLER_26_280 ();
 sg13g2_decap_4 FILLER_26_285 ();
 sg13g2_fill_1 FILLER_26_289 ();
 sg13g2_fill_2 FILLER_26_316 ();
 sg13g2_fill_2 FILLER_26_344 ();
 sg13g2_decap_8 FILLER_26_372 ();
 sg13g2_fill_2 FILLER_26_387 ();
 sg13g2_fill_1 FILLER_26_389 ();
 sg13g2_fill_1 FILLER_26_416 ();
 sg13g2_decap_8 FILLER_26_457 ();
 sg13g2_fill_1 FILLER_26_464 ();
 sg13g2_decap_8 FILLER_26_469 ();
 sg13g2_fill_1 FILLER_26_476 ();
 sg13g2_decap_8 FILLER_26_503 ();
 sg13g2_decap_4 FILLER_26_510 ();
 sg13g2_decap_4 FILLER_26_527 ();
 sg13g2_decap_8 FILLER_26_560 ();
 sg13g2_fill_2 FILLER_26_567 ();
 sg13g2_fill_1 FILLER_26_576 ();
 sg13g2_decap_8 FILLER_26_588 ();
 sg13g2_decap_8 FILLER_26_595 ();
 sg13g2_fill_2 FILLER_26_602 ();
 sg13g2_fill_1 FILLER_26_604 ();
 sg13g2_fill_2 FILLER_26_665 ();
 sg13g2_decap_8 FILLER_26_680 ();
 sg13g2_decap_8 FILLER_26_687 ();
 sg13g2_decap_8 FILLER_26_694 ();
 sg13g2_decap_8 FILLER_26_701 ();
 sg13g2_decap_8 FILLER_26_708 ();
 sg13g2_decap_8 FILLER_26_715 ();
 sg13g2_decap_8 FILLER_26_722 ();
 sg13g2_decap_8 FILLER_26_729 ();
 sg13g2_decap_8 FILLER_26_736 ();
 sg13g2_decap_8 FILLER_26_743 ();
 sg13g2_decap_8 FILLER_26_750 ();
 sg13g2_decap_8 FILLER_26_757 ();
 sg13g2_decap_8 FILLER_26_764 ();
 sg13g2_decap_8 FILLER_26_771 ();
 sg13g2_decap_8 FILLER_26_778 ();
 sg13g2_decap_8 FILLER_26_785 ();
 sg13g2_decap_8 FILLER_26_792 ();
 sg13g2_decap_8 FILLER_26_799 ();
 sg13g2_decap_8 FILLER_26_806 ();
 sg13g2_decap_8 FILLER_26_813 ();
 sg13g2_decap_8 FILLER_26_820 ();
 sg13g2_decap_8 FILLER_26_827 ();
 sg13g2_decap_8 FILLER_26_834 ();
 sg13g2_decap_8 FILLER_26_841 ();
 sg13g2_decap_8 FILLER_26_848 ();
 sg13g2_decap_8 FILLER_26_855 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_fill_2 FILLER_27_194 ();
 sg13g2_fill_1 FILLER_27_201 ();
 sg13g2_decap_8 FILLER_27_228 ();
 sg13g2_fill_1 FILLER_27_235 ();
 sg13g2_fill_2 FILLER_27_263 ();
 sg13g2_fill_1 FILLER_27_299 ();
 sg13g2_decap_8 FILLER_27_304 ();
 sg13g2_decap_4 FILLER_27_311 ();
 sg13g2_fill_2 FILLER_27_315 ();
 sg13g2_fill_1 FILLER_27_326 ();
 sg13g2_decap_8 FILLER_27_339 ();
 sg13g2_decap_4 FILLER_27_351 ();
 sg13g2_fill_2 FILLER_27_355 ();
 sg13g2_decap_8 FILLER_27_391 ();
 sg13g2_fill_1 FILLER_27_398 ();
 sg13g2_decap_8 FILLER_27_416 ();
 sg13g2_decap_4 FILLER_27_423 ();
 sg13g2_fill_1 FILLER_27_427 ();
 sg13g2_decap_4 FILLER_27_446 ();
 sg13g2_fill_1 FILLER_27_450 ();
 sg13g2_fill_2 FILLER_27_469 ();
 sg13g2_fill_1 FILLER_27_471 ();
 sg13g2_fill_2 FILLER_27_482 ();
 sg13g2_decap_4 FILLER_27_524 ();
 sg13g2_fill_1 FILLER_27_532 ();
 sg13g2_fill_2 FILLER_27_538 ();
 sg13g2_fill_1 FILLER_27_540 ();
 sg13g2_fill_1 FILLER_27_550 ();
 sg13g2_fill_2 FILLER_27_563 ();
 sg13g2_fill_1 FILLER_27_565 ();
 sg13g2_decap_4 FILLER_27_592 ();
 sg13g2_fill_1 FILLER_27_596 ();
 sg13g2_decap_8 FILLER_27_623 ();
 sg13g2_fill_2 FILLER_27_630 ();
 sg13g2_decap_8 FILLER_27_636 ();
 sg13g2_decap_8 FILLER_27_643 ();
 sg13g2_decap_8 FILLER_27_650 ();
 sg13g2_decap_4 FILLER_27_657 ();
 sg13g2_fill_2 FILLER_27_661 ();
 sg13g2_decap_8 FILLER_27_687 ();
 sg13g2_decap_8 FILLER_27_694 ();
 sg13g2_decap_8 FILLER_27_701 ();
 sg13g2_decap_8 FILLER_27_708 ();
 sg13g2_decap_8 FILLER_27_715 ();
 sg13g2_decap_8 FILLER_27_722 ();
 sg13g2_decap_8 FILLER_27_729 ();
 sg13g2_decap_8 FILLER_27_736 ();
 sg13g2_decap_8 FILLER_27_743 ();
 sg13g2_decap_8 FILLER_27_750 ();
 sg13g2_decap_8 FILLER_27_757 ();
 sg13g2_decap_8 FILLER_27_764 ();
 sg13g2_decap_8 FILLER_27_771 ();
 sg13g2_decap_8 FILLER_27_778 ();
 sg13g2_decap_8 FILLER_27_785 ();
 sg13g2_decap_8 FILLER_27_792 ();
 sg13g2_decap_8 FILLER_27_799 ();
 sg13g2_decap_8 FILLER_27_806 ();
 sg13g2_decap_8 FILLER_27_813 ();
 sg13g2_decap_8 FILLER_27_820 ();
 sg13g2_decap_8 FILLER_27_827 ();
 sg13g2_decap_8 FILLER_27_834 ();
 sg13g2_decap_8 FILLER_27_841 ();
 sg13g2_decap_8 FILLER_27_848 ();
 sg13g2_decap_8 FILLER_27_855 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_4 FILLER_28_182 ();
 sg13g2_fill_2 FILLER_28_194 ();
 sg13g2_decap_8 FILLER_28_216 ();
 sg13g2_decap_4 FILLER_28_223 ();
 sg13g2_fill_1 FILLER_28_227 ();
 sg13g2_fill_1 FILLER_28_253 ();
 sg13g2_fill_2 FILLER_28_272 ();
 sg13g2_fill_1 FILLER_28_274 ();
 sg13g2_decap_4 FILLER_28_279 ();
 sg13g2_fill_2 FILLER_28_283 ();
 sg13g2_decap_4 FILLER_28_299 ();
 sg13g2_fill_1 FILLER_28_334 ();
 sg13g2_decap_4 FILLER_28_378 ();
 sg13g2_fill_1 FILLER_28_382 ();
 sg13g2_fill_1 FILLER_28_432 ();
 sg13g2_fill_1 FILLER_28_457 ();
 sg13g2_fill_2 FILLER_28_463 ();
 sg13g2_fill_2 FILLER_28_486 ();
 sg13g2_fill_1 FILLER_28_488 ();
 sg13g2_decap_8 FILLER_28_498 ();
 sg13g2_fill_2 FILLER_28_505 ();
 sg13g2_fill_1 FILLER_28_507 ();
 sg13g2_fill_2 FILLER_28_521 ();
 sg13g2_fill_1 FILLER_28_523 ();
 sg13g2_fill_2 FILLER_28_557 ();
 sg13g2_decap_4 FILLER_28_571 ();
 sg13g2_fill_2 FILLER_28_575 ();
 sg13g2_decap_8 FILLER_28_595 ();
 sg13g2_fill_1 FILLER_28_602 ();
 sg13g2_fill_1 FILLER_28_607 ();
 sg13g2_decap_8 FILLER_28_612 ();
 sg13g2_fill_2 FILLER_28_619 ();
 sg13g2_fill_2 FILLER_28_678 ();
 sg13g2_decap_8 FILLER_28_700 ();
 sg13g2_decap_8 FILLER_28_707 ();
 sg13g2_decap_8 FILLER_28_714 ();
 sg13g2_decap_8 FILLER_28_721 ();
 sg13g2_decap_8 FILLER_28_728 ();
 sg13g2_decap_8 FILLER_28_735 ();
 sg13g2_decap_8 FILLER_28_742 ();
 sg13g2_decap_8 FILLER_28_749 ();
 sg13g2_decap_8 FILLER_28_756 ();
 sg13g2_decap_8 FILLER_28_763 ();
 sg13g2_decap_8 FILLER_28_770 ();
 sg13g2_decap_8 FILLER_28_777 ();
 sg13g2_decap_8 FILLER_28_784 ();
 sg13g2_decap_8 FILLER_28_791 ();
 sg13g2_decap_8 FILLER_28_798 ();
 sg13g2_decap_8 FILLER_28_805 ();
 sg13g2_decap_8 FILLER_28_812 ();
 sg13g2_decap_8 FILLER_28_819 ();
 sg13g2_decap_8 FILLER_28_826 ();
 sg13g2_decap_8 FILLER_28_833 ();
 sg13g2_decap_8 FILLER_28_840 ();
 sg13g2_decap_8 FILLER_28_847 ();
 sg13g2_decap_8 FILLER_28_854 ();
 sg13g2_fill_1 FILLER_28_861 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_4 FILLER_29_175 ();
 sg13g2_fill_1 FILLER_29_199 ();
 sg13g2_decap_4 FILLER_29_278 ();
 sg13g2_decap_8 FILLER_29_286 ();
 sg13g2_fill_1 FILLER_29_293 ();
 sg13g2_decap_8 FILLER_29_298 ();
 sg13g2_fill_2 FILLER_29_305 ();
 sg13g2_fill_1 FILLER_29_307 ();
 sg13g2_decap_8 FILLER_29_339 ();
 sg13g2_decap_4 FILLER_29_350 ();
 sg13g2_fill_2 FILLER_29_354 ();
 sg13g2_fill_2 FILLER_29_364 ();
 sg13g2_fill_1 FILLER_29_366 ();
 sg13g2_decap_4 FILLER_29_375 ();
 sg13g2_decap_8 FILLER_29_390 ();
 sg13g2_fill_1 FILLER_29_397 ();
 sg13g2_fill_2 FILLER_29_412 ();
 sg13g2_decap_8 FILLER_29_441 ();
 sg13g2_fill_2 FILLER_29_448 ();
 sg13g2_fill_1 FILLER_29_450 ();
 sg13g2_fill_2 FILLER_29_476 ();
 sg13g2_fill_1 FILLER_29_478 ();
 sg13g2_decap_4 FILLER_29_515 ();
 sg13g2_fill_1 FILLER_29_519 ();
 sg13g2_fill_1 FILLER_29_524 ();
 sg13g2_fill_2 FILLER_29_528 ();
 sg13g2_fill_1 FILLER_29_530 ();
 sg13g2_fill_1 FILLER_29_540 ();
 sg13g2_fill_1 FILLER_29_557 ();
 sg13g2_decap_4 FILLER_29_571 ();
 sg13g2_decap_4 FILLER_29_580 ();
 sg13g2_fill_2 FILLER_29_584 ();
 sg13g2_fill_2 FILLER_29_591 ();
 sg13g2_decap_4 FILLER_29_619 ();
 sg13g2_fill_1 FILLER_29_623 ();
 sg13g2_decap_8 FILLER_29_640 ();
 sg13g2_decap_8 FILLER_29_647 ();
 sg13g2_fill_1 FILLER_29_654 ();
 sg13g2_fill_1 FILLER_29_659 ();
 sg13g2_fill_1 FILLER_29_672 ();
 sg13g2_decap_8 FILLER_29_713 ();
 sg13g2_decap_8 FILLER_29_720 ();
 sg13g2_decap_8 FILLER_29_727 ();
 sg13g2_decap_8 FILLER_29_734 ();
 sg13g2_decap_8 FILLER_29_741 ();
 sg13g2_decap_8 FILLER_29_748 ();
 sg13g2_decap_8 FILLER_29_755 ();
 sg13g2_decap_8 FILLER_29_762 ();
 sg13g2_decap_8 FILLER_29_769 ();
 sg13g2_decap_8 FILLER_29_776 ();
 sg13g2_decap_8 FILLER_29_783 ();
 sg13g2_decap_8 FILLER_29_790 ();
 sg13g2_decap_8 FILLER_29_797 ();
 sg13g2_decap_8 FILLER_29_804 ();
 sg13g2_decap_8 FILLER_29_811 ();
 sg13g2_decap_8 FILLER_29_818 ();
 sg13g2_decap_8 FILLER_29_825 ();
 sg13g2_decap_8 FILLER_29_832 ();
 sg13g2_decap_8 FILLER_29_839 ();
 sg13g2_decap_8 FILLER_29_846 ();
 sg13g2_decap_8 FILLER_29_853 ();
 sg13g2_fill_2 FILLER_29_860 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_fill_1 FILLER_30_175 ();
 sg13g2_fill_2 FILLER_30_186 ();
 sg13g2_fill_1 FILLER_30_188 ();
 sg13g2_fill_1 FILLER_30_205 ();
 sg13g2_decap_8 FILLER_30_211 ();
 sg13g2_decap_4 FILLER_30_218 ();
 sg13g2_fill_1 FILLER_30_222 ();
 sg13g2_decap_4 FILLER_30_231 ();
 sg13g2_fill_1 FILLER_30_235 ();
 sg13g2_decap_8 FILLER_30_240 ();
 sg13g2_decap_8 FILLER_30_247 ();
 sg13g2_decap_4 FILLER_30_254 ();
 sg13g2_fill_2 FILLER_30_258 ();
 sg13g2_fill_2 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_310 ();
 sg13g2_decap_4 FILLER_30_317 ();
 sg13g2_decap_8 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_fill_2 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_349 ();
 sg13g2_fill_2 FILLER_30_356 ();
 sg13g2_fill_1 FILLER_30_358 ();
 sg13g2_fill_1 FILLER_30_393 ();
 sg13g2_fill_2 FILLER_30_435 ();
 sg13g2_fill_1 FILLER_30_464 ();
 sg13g2_decap_8 FILLER_30_479 ();
 sg13g2_decap_4 FILLER_30_486 ();
 sg13g2_fill_1 FILLER_30_490 ();
 sg13g2_fill_2 FILLER_30_527 ();
 sg13g2_fill_1 FILLER_30_542 ();
 sg13g2_decap_8 FILLER_30_556 ();
 sg13g2_decap_4 FILLER_30_563 ();
 sg13g2_fill_1 FILLER_30_567 ();
 sg13g2_fill_1 FILLER_30_586 ();
 sg13g2_decap_4 FILLER_30_613 ();
 sg13g2_fill_1 FILLER_30_617 ();
 sg13g2_fill_2 FILLER_30_630 ();
 sg13g2_fill_1 FILLER_30_648 ();
 sg13g2_fill_2 FILLER_30_675 ();
 sg13g2_fill_1 FILLER_30_677 ();
 sg13g2_decap_8 FILLER_30_704 ();
 sg13g2_decap_8 FILLER_30_711 ();
 sg13g2_decap_8 FILLER_30_718 ();
 sg13g2_decap_8 FILLER_30_725 ();
 sg13g2_decap_8 FILLER_30_732 ();
 sg13g2_decap_8 FILLER_30_739 ();
 sg13g2_decap_8 FILLER_30_746 ();
 sg13g2_decap_8 FILLER_30_753 ();
 sg13g2_decap_8 FILLER_30_760 ();
 sg13g2_decap_8 FILLER_30_767 ();
 sg13g2_decap_8 FILLER_30_774 ();
 sg13g2_decap_8 FILLER_30_781 ();
 sg13g2_decap_8 FILLER_30_788 ();
 sg13g2_decap_8 FILLER_30_795 ();
 sg13g2_decap_8 FILLER_30_802 ();
 sg13g2_decap_8 FILLER_30_809 ();
 sg13g2_decap_8 FILLER_30_816 ();
 sg13g2_decap_8 FILLER_30_823 ();
 sg13g2_decap_8 FILLER_30_830 ();
 sg13g2_decap_8 FILLER_30_837 ();
 sg13g2_decap_8 FILLER_30_844 ();
 sg13g2_decap_8 FILLER_30_851 ();
 sg13g2_decap_4 FILLER_30_858 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_fill_2 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_195 ();
 sg13g2_decap_4 FILLER_31_202 ();
 sg13g2_fill_1 FILLER_31_215 ();
 sg13g2_fill_1 FILLER_31_221 ();
 sg13g2_fill_2 FILLER_31_234 ();
 sg13g2_fill_1 FILLER_31_236 ();
 sg13g2_fill_2 FILLER_31_251 ();
 sg13g2_decap_4 FILLER_31_261 ();
 sg13g2_fill_2 FILLER_31_265 ();
 sg13g2_fill_2 FILLER_31_276 ();
 sg13g2_fill_1 FILLER_31_278 ();
 sg13g2_decap_8 FILLER_31_284 ();
 sg13g2_fill_2 FILLER_31_305 ();
 sg13g2_fill_1 FILLER_31_307 ();
 sg13g2_decap_8 FILLER_31_360 ();
 sg13g2_fill_2 FILLER_31_367 ();
 sg13g2_fill_1 FILLER_31_369 ();
 sg13g2_decap_8 FILLER_31_374 ();
 sg13g2_decap_4 FILLER_31_381 ();
 sg13g2_decap_4 FILLER_31_390 ();
 sg13g2_fill_2 FILLER_31_394 ();
 sg13g2_decap_4 FILLER_31_400 ();
 sg13g2_fill_1 FILLER_31_404 ();
 sg13g2_decap_4 FILLER_31_409 ();
 sg13g2_decap_4 FILLER_31_433 ();
 sg13g2_fill_2 FILLER_31_437 ();
 sg13g2_fill_1 FILLER_31_450 ();
 sg13g2_decap_8 FILLER_31_487 ();
 sg13g2_fill_1 FILLER_31_494 ();
 sg13g2_fill_2 FILLER_31_518 ();
 sg13g2_fill_1 FILLER_31_544 ();
 sg13g2_decap_4 FILLER_31_574 ();
 sg13g2_decap_8 FILLER_31_583 ();
 sg13g2_decap_8 FILLER_31_590 ();
 sg13g2_decap_8 FILLER_31_605 ();
 sg13g2_decap_8 FILLER_31_612 ();
 sg13g2_decap_8 FILLER_31_619 ();
 sg13g2_fill_1 FILLER_31_626 ();
 sg13g2_fill_2 FILLER_31_647 ();
 sg13g2_decap_8 FILLER_31_665 ();
 sg13g2_decap_8 FILLER_31_672 ();
 sg13g2_fill_2 FILLER_31_696 ();
 sg13g2_fill_1 FILLER_31_698 ();
 sg13g2_decap_8 FILLER_31_725 ();
 sg13g2_decap_8 FILLER_31_732 ();
 sg13g2_decap_8 FILLER_31_739 ();
 sg13g2_decap_8 FILLER_31_746 ();
 sg13g2_decap_8 FILLER_31_753 ();
 sg13g2_decap_8 FILLER_31_760 ();
 sg13g2_decap_8 FILLER_31_767 ();
 sg13g2_decap_8 FILLER_31_774 ();
 sg13g2_decap_8 FILLER_31_781 ();
 sg13g2_decap_8 FILLER_31_788 ();
 sg13g2_decap_8 FILLER_31_795 ();
 sg13g2_decap_8 FILLER_31_802 ();
 sg13g2_decap_8 FILLER_31_809 ();
 sg13g2_decap_8 FILLER_31_816 ();
 sg13g2_decap_8 FILLER_31_823 ();
 sg13g2_decap_8 FILLER_31_830 ();
 sg13g2_decap_8 FILLER_31_837 ();
 sg13g2_decap_8 FILLER_31_844 ();
 sg13g2_decap_8 FILLER_31_851 ();
 sg13g2_decap_4 FILLER_31_858 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_4 FILLER_32_161 ();
 sg13g2_fill_1 FILLER_32_165 ();
 sg13g2_fill_2 FILLER_32_186 ();
 sg13g2_fill_1 FILLER_32_188 ();
 sg13g2_decap_4 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_229 ();
 sg13g2_decap_4 FILLER_32_236 ();
 sg13g2_fill_1 FILLER_32_265 ();
 sg13g2_fill_2 FILLER_32_281 ();
 sg13g2_fill_1 FILLER_32_291 ();
 sg13g2_decap_4 FILLER_32_298 ();
 sg13g2_fill_1 FILLER_32_302 ();
 sg13g2_decap_8 FILLER_32_310 ();
 sg13g2_decap_8 FILLER_32_317 ();
 sg13g2_decap_4 FILLER_32_324 ();
 sg13g2_fill_2 FILLER_32_342 ();
 sg13g2_fill_2 FILLER_32_351 ();
 sg13g2_fill_1 FILLER_32_353 ();
 sg13g2_decap_8 FILLER_32_363 ();
 sg13g2_fill_1 FILLER_32_370 ();
 sg13g2_decap_4 FILLER_32_384 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_418 ();
 sg13g2_decap_8 FILLER_32_445 ();
 sg13g2_fill_2 FILLER_32_457 ();
 sg13g2_decap_8 FILLER_32_473 ();
 sg13g2_decap_8 FILLER_32_480 ();
 sg13g2_decap_4 FILLER_32_487 ();
 sg13g2_fill_1 FILLER_32_491 ();
 sg13g2_fill_2 FILLER_32_518 ();
 sg13g2_fill_2 FILLER_32_528 ();
 sg13g2_fill_2 FILLER_32_556 ();
 sg13g2_decap_4 FILLER_32_584 ();
 sg13g2_fill_2 FILLER_32_588 ();
 sg13g2_decap_8 FILLER_32_620 ();
 sg13g2_decap_8 FILLER_32_627 ();
 sg13g2_fill_2 FILLER_32_634 ();
 sg13g2_fill_1 FILLER_32_640 ();
 sg13g2_decap_8 FILLER_32_672 ();
 sg13g2_decap_4 FILLER_32_705 ();
 sg13g2_fill_1 FILLER_32_709 ();
 sg13g2_decap_8 FILLER_32_714 ();
 sg13g2_decap_8 FILLER_32_721 ();
 sg13g2_decap_8 FILLER_32_728 ();
 sg13g2_decap_8 FILLER_32_735 ();
 sg13g2_decap_8 FILLER_32_742 ();
 sg13g2_decap_8 FILLER_32_749 ();
 sg13g2_decap_8 FILLER_32_756 ();
 sg13g2_decap_8 FILLER_32_763 ();
 sg13g2_decap_8 FILLER_32_770 ();
 sg13g2_decap_8 FILLER_32_777 ();
 sg13g2_decap_8 FILLER_32_784 ();
 sg13g2_decap_8 FILLER_32_791 ();
 sg13g2_decap_8 FILLER_32_798 ();
 sg13g2_decap_8 FILLER_32_805 ();
 sg13g2_decap_8 FILLER_32_812 ();
 sg13g2_decap_8 FILLER_32_819 ();
 sg13g2_decap_8 FILLER_32_826 ();
 sg13g2_decap_8 FILLER_32_833 ();
 sg13g2_decap_8 FILLER_32_840 ();
 sg13g2_decap_8 FILLER_32_847 ();
 sg13g2_decap_8 FILLER_32_854 ();
 sg13g2_fill_1 FILLER_32_861 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_fill_2 FILLER_33_154 ();
 sg13g2_fill_2 FILLER_33_178 ();
 sg13g2_fill_1 FILLER_33_188 ();
 sg13g2_fill_2 FILLER_33_193 ();
 sg13g2_fill_1 FILLER_33_195 ();
 sg13g2_fill_2 FILLER_33_204 ();
 sg13g2_fill_1 FILLER_33_206 ();
 sg13g2_decap_8 FILLER_33_232 ();
 sg13g2_decap_8 FILLER_33_239 ();
 sg13g2_decap_4 FILLER_33_246 ();
 sg13g2_fill_1 FILLER_33_250 ();
 sg13g2_decap_8 FILLER_33_256 ();
 sg13g2_fill_2 FILLER_33_263 ();
 sg13g2_fill_1 FILLER_33_265 ();
 sg13g2_decap_8 FILLER_33_270 ();
 sg13g2_fill_1 FILLER_33_292 ();
 sg13g2_decap_4 FILLER_33_321 ();
 sg13g2_fill_2 FILLER_33_325 ();
 sg13g2_fill_2 FILLER_33_340 ();
 sg13g2_fill_1 FILLER_33_342 ();
 sg13g2_fill_2 FILLER_33_360 ();
 sg13g2_fill_2 FILLER_33_392 ();
 sg13g2_fill_1 FILLER_33_394 ();
 sg13g2_decap_8 FILLER_33_421 ();
 sg13g2_fill_2 FILLER_33_428 ();
 sg13g2_decap_8 FILLER_33_434 ();
 sg13g2_decap_4 FILLER_33_441 ();
 sg13g2_fill_1 FILLER_33_445 ();
 sg13g2_decap_8 FILLER_33_547 ();
 sg13g2_decap_4 FILLER_33_554 ();
 sg13g2_fill_1 FILLER_33_558 ();
 sg13g2_fill_2 FILLER_33_595 ();
 sg13g2_fill_1 FILLER_33_631 ();
 sg13g2_fill_2 FILLER_33_644 ();
 sg13g2_fill_1 FILLER_33_660 ();
 sg13g2_decap_4 FILLER_33_669 ();
 sg13g2_decap_8 FILLER_33_706 ();
 sg13g2_decap_8 FILLER_33_713 ();
 sg13g2_decap_8 FILLER_33_720 ();
 sg13g2_decap_8 FILLER_33_727 ();
 sg13g2_decap_8 FILLER_33_734 ();
 sg13g2_decap_8 FILLER_33_741 ();
 sg13g2_decap_8 FILLER_33_748 ();
 sg13g2_decap_8 FILLER_33_755 ();
 sg13g2_decap_8 FILLER_33_762 ();
 sg13g2_decap_8 FILLER_33_769 ();
 sg13g2_decap_8 FILLER_33_776 ();
 sg13g2_decap_8 FILLER_33_783 ();
 sg13g2_decap_8 FILLER_33_790 ();
 sg13g2_decap_8 FILLER_33_797 ();
 sg13g2_decap_8 FILLER_33_804 ();
 sg13g2_decap_8 FILLER_33_811 ();
 sg13g2_decap_8 FILLER_33_818 ();
 sg13g2_decap_8 FILLER_33_825 ();
 sg13g2_decap_8 FILLER_33_832 ();
 sg13g2_decap_8 FILLER_33_839 ();
 sg13g2_decap_8 FILLER_33_846 ();
 sg13g2_decap_8 FILLER_33_853 ();
 sg13g2_fill_2 FILLER_33_860 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_fill_1 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_fill_1 FILLER_34_203 ();
 sg13g2_fill_2 FILLER_34_221 ();
 sg13g2_fill_1 FILLER_34_223 ();
 sg13g2_fill_1 FILLER_34_281 ();
 sg13g2_fill_1 FILLER_34_317 ();
 sg13g2_fill_2 FILLER_34_330 ();
 sg13g2_decap_4 FILLER_34_337 ();
 sg13g2_fill_1 FILLER_34_354 ();
 sg13g2_fill_2 FILLER_34_360 ();
 sg13g2_decap_4 FILLER_34_372 ();
 sg13g2_fill_1 FILLER_34_376 ();
 sg13g2_decap_8 FILLER_34_381 ();
 sg13g2_decap_4 FILLER_34_388 ();
 sg13g2_fill_2 FILLER_34_403 ();
 sg13g2_fill_1 FILLER_34_405 ();
 sg13g2_fill_2 FILLER_34_443 ();
 sg13g2_fill_2 FILLER_34_453 ();
 sg13g2_decap_4 FILLER_34_494 ();
 sg13g2_fill_2 FILLER_34_498 ();
 sg13g2_fill_2 FILLER_34_505 ();
 sg13g2_fill_1 FILLER_34_507 ();
 sg13g2_fill_1 FILLER_34_522 ();
 sg13g2_fill_1 FILLER_34_573 ();
 sg13g2_decap_4 FILLER_34_629 ();
 sg13g2_decap_4 FILLER_34_638 ();
 sg13g2_fill_2 FILLER_34_642 ();
 sg13g2_fill_2 FILLER_34_652 ();
 sg13g2_fill_1 FILLER_34_672 ();
 sg13g2_decap_8 FILLER_34_678 ();
 sg13g2_fill_1 FILLER_34_685 ();
 sg13g2_decap_8 FILLER_34_696 ();
 sg13g2_decap_8 FILLER_34_703 ();
 sg13g2_decap_8 FILLER_34_710 ();
 sg13g2_decap_8 FILLER_34_717 ();
 sg13g2_decap_8 FILLER_34_724 ();
 sg13g2_decap_8 FILLER_34_731 ();
 sg13g2_decap_8 FILLER_34_738 ();
 sg13g2_decap_8 FILLER_34_745 ();
 sg13g2_decap_8 FILLER_34_752 ();
 sg13g2_decap_8 FILLER_34_759 ();
 sg13g2_decap_8 FILLER_34_766 ();
 sg13g2_decap_8 FILLER_34_773 ();
 sg13g2_decap_8 FILLER_34_780 ();
 sg13g2_decap_8 FILLER_34_787 ();
 sg13g2_decap_8 FILLER_34_794 ();
 sg13g2_decap_8 FILLER_34_801 ();
 sg13g2_decap_8 FILLER_34_808 ();
 sg13g2_decap_8 FILLER_34_815 ();
 sg13g2_decap_8 FILLER_34_822 ();
 sg13g2_decap_8 FILLER_34_829 ();
 sg13g2_decap_8 FILLER_34_836 ();
 sg13g2_decap_8 FILLER_34_843 ();
 sg13g2_decap_8 FILLER_34_850 ();
 sg13g2_decap_4 FILLER_34_857 ();
 sg13g2_fill_1 FILLER_34_861 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_fill_1 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_184 ();
 sg13g2_fill_2 FILLER_35_191 ();
 sg13g2_fill_1 FILLER_35_193 ();
 sg13g2_fill_2 FILLER_35_198 ();
 sg13g2_fill_2 FILLER_35_230 ();
 sg13g2_fill_1 FILLER_35_242 ();
 sg13g2_fill_2 FILLER_35_259 ();
 sg13g2_fill_2 FILLER_35_300 ();
 sg13g2_fill_1 FILLER_35_302 ();
 sg13g2_decap_8 FILLER_35_320 ();
 sg13g2_fill_1 FILLER_35_327 ();
 sg13g2_decap_8 FILLER_35_348 ();
 sg13g2_fill_1 FILLER_35_355 ();
 sg13g2_fill_1 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_379 ();
 sg13g2_fill_2 FILLER_35_386 ();
 sg13g2_fill_1 FILLER_35_388 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_fill_1 FILLER_35_426 ();
 sg13g2_fill_1 FILLER_35_444 ();
 sg13g2_decap_4 FILLER_35_459 ();
 sg13g2_fill_1 FILLER_35_466 ();
 sg13g2_fill_2 FILLER_35_489 ();
 sg13g2_fill_2 FILLER_35_496 ();
 sg13g2_fill_1 FILLER_35_498 ();
 sg13g2_fill_1 FILLER_35_507 ();
 sg13g2_decap_4 FILLER_35_550 ();
 sg13g2_fill_1 FILLER_35_554 ();
 sg13g2_fill_1 FILLER_35_575 ();
 sg13g2_fill_2 FILLER_35_594 ();
 sg13g2_fill_1 FILLER_35_596 ();
 sg13g2_fill_1 FILLER_35_606 ();
 sg13g2_fill_2 FILLER_35_644 ();
 sg13g2_fill_1 FILLER_35_660 ();
 sg13g2_fill_2 FILLER_35_665 ();
 sg13g2_fill_2 FILLER_35_682 ();
 sg13g2_decap_8 FILLER_35_697 ();
 sg13g2_decap_8 FILLER_35_704 ();
 sg13g2_decap_8 FILLER_35_711 ();
 sg13g2_decap_8 FILLER_35_718 ();
 sg13g2_decap_8 FILLER_35_725 ();
 sg13g2_decap_8 FILLER_35_732 ();
 sg13g2_decap_8 FILLER_35_739 ();
 sg13g2_decap_8 FILLER_35_746 ();
 sg13g2_decap_8 FILLER_35_753 ();
 sg13g2_decap_8 FILLER_35_760 ();
 sg13g2_decap_8 FILLER_35_767 ();
 sg13g2_decap_8 FILLER_35_774 ();
 sg13g2_decap_8 FILLER_35_781 ();
 sg13g2_decap_8 FILLER_35_788 ();
 sg13g2_decap_8 FILLER_35_795 ();
 sg13g2_decap_8 FILLER_35_802 ();
 sg13g2_decap_8 FILLER_35_809 ();
 sg13g2_decap_8 FILLER_35_816 ();
 sg13g2_decap_8 FILLER_35_823 ();
 sg13g2_decap_8 FILLER_35_830 ();
 sg13g2_decap_8 FILLER_35_837 ();
 sg13g2_decap_8 FILLER_35_844 ();
 sg13g2_decap_8 FILLER_35_851 ();
 sg13g2_decap_4 FILLER_35_858 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_fill_2 FILLER_36_140 ();
 sg13g2_fill_1 FILLER_36_142 ();
 sg13g2_decap_4 FILLER_36_169 ();
 sg13g2_fill_1 FILLER_36_228 ();
 sg13g2_fill_1 FILLER_36_242 ();
 sg13g2_fill_1 FILLER_36_257 ();
 sg13g2_fill_2 FILLER_36_273 ();
 sg13g2_fill_1 FILLER_36_275 ();
 sg13g2_fill_2 FILLER_36_317 ();
 sg13g2_fill_1 FILLER_36_319 ();
 sg13g2_fill_2 FILLER_36_325 ();
 sg13g2_fill_1 FILLER_36_327 ();
 sg13g2_fill_2 FILLER_36_340 ();
 sg13g2_fill_1 FILLER_36_342 ();
 sg13g2_decap_8 FILLER_36_370 ();
 sg13g2_decap_4 FILLER_36_479 ();
 sg13g2_fill_1 FILLER_36_483 ();
 sg13g2_fill_1 FILLER_36_509 ();
 sg13g2_decap_8 FILLER_36_536 ();
 sg13g2_fill_2 FILLER_36_543 ();
 sg13g2_fill_1 FILLER_36_545 ();
 sg13g2_fill_2 FILLER_36_572 ();
 sg13g2_fill_1 FILLER_36_574 ();
 sg13g2_fill_1 FILLER_36_579 ();
 sg13g2_fill_2 FILLER_36_632 ();
 sg13g2_fill_1 FILLER_36_634 ();
 sg13g2_fill_1 FILLER_36_666 ();
 sg13g2_decap_8 FILLER_36_675 ();
 sg13g2_fill_2 FILLER_36_682 ();
 sg13g2_decap_8 FILLER_36_705 ();
 sg13g2_decap_8 FILLER_36_712 ();
 sg13g2_decap_8 FILLER_36_719 ();
 sg13g2_decap_8 FILLER_36_726 ();
 sg13g2_decap_8 FILLER_36_733 ();
 sg13g2_decap_8 FILLER_36_740 ();
 sg13g2_decap_8 FILLER_36_747 ();
 sg13g2_decap_8 FILLER_36_754 ();
 sg13g2_decap_8 FILLER_36_761 ();
 sg13g2_decap_8 FILLER_36_768 ();
 sg13g2_decap_8 FILLER_36_775 ();
 sg13g2_decap_8 FILLER_36_782 ();
 sg13g2_decap_8 FILLER_36_789 ();
 sg13g2_decap_8 FILLER_36_796 ();
 sg13g2_decap_8 FILLER_36_803 ();
 sg13g2_decap_8 FILLER_36_810 ();
 sg13g2_decap_8 FILLER_36_817 ();
 sg13g2_decap_8 FILLER_36_824 ();
 sg13g2_decap_8 FILLER_36_831 ();
 sg13g2_decap_8 FILLER_36_838 ();
 sg13g2_decap_8 FILLER_36_845 ();
 sg13g2_decap_8 FILLER_36_852 ();
 sg13g2_fill_2 FILLER_36_859 ();
 sg13g2_fill_1 FILLER_36_861 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_4 FILLER_37_162 ();
 sg13g2_fill_1 FILLER_37_166 ();
 sg13g2_fill_2 FILLER_37_206 ();
 sg13g2_fill_1 FILLER_37_208 ();
 sg13g2_decap_4 FILLER_37_245 ();
 sg13g2_fill_2 FILLER_37_313 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_fill_2 FILLER_37_343 ();
 sg13g2_fill_1 FILLER_37_358 ();
 sg13g2_fill_2 FILLER_37_365 ();
 sg13g2_fill_1 FILLER_37_367 ();
 sg13g2_decap_8 FILLER_37_395 ();
 sg13g2_fill_2 FILLER_37_402 ();
 sg13g2_fill_1 FILLER_37_404 ();
 sg13g2_fill_1 FILLER_37_415 ();
 sg13g2_fill_2 FILLER_37_426 ();
 sg13g2_fill_1 FILLER_37_428 ();
 sg13g2_fill_2 FILLER_37_434 ();
 sg13g2_fill_1 FILLER_37_444 ();
 sg13g2_fill_2 FILLER_37_450 ();
 sg13g2_fill_1 FILLER_37_452 ();
 sg13g2_fill_2 FILLER_37_461 ();
 sg13g2_fill_1 FILLER_37_463 ();
 sg13g2_decap_8 FILLER_37_479 ();
 sg13g2_decap_8 FILLER_37_486 ();
 sg13g2_decap_4 FILLER_37_493 ();
 sg13g2_fill_1 FILLER_37_497 ();
 sg13g2_decap_4 FILLER_37_508 ();
 sg13g2_fill_2 FILLER_37_533 ();
 sg13g2_fill_1 FILLER_37_545 ();
 sg13g2_fill_1 FILLER_37_563 ();
 sg13g2_fill_1 FILLER_37_609 ();
 sg13g2_fill_2 FILLER_37_631 ();
 sg13g2_fill_1 FILLER_37_633 ();
 sg13g2_decap_4 FILLER_37_697 ();
 sg13g2_decap_8 FILLER_37_727 ();
 sg13g2_decap_8 FILLER_37_734 ();
 sg13g2_decap_8 FILLER_37_741 ();
 sg13g2_decap_8 FILLER_37_748 ();
 sg13g2_decap_8 FILLER_37_755 ();
 sg13g2_decap_8 FILLER_37_762 ();
 sg13g2_decap_8 FILLER_37_769 ();
 sg13g2_decap_8 FILLER_37_776 ();
 sg13g2_decap_8 FILLER_37_783 ();
 sg13g2_decap_8 FILLER_37_790 ();
 sg13g2_decap_8 FILLER_37_797 ();
 sg13g2_decap_8 FILLER_37_804 ();
 sg13g2_decap_8 FILLER_37_811 ();
 sg13g2_decap_8 FILLER_37_818 ();
 sg13g2_decap_8 FILLER_37_825 ();
 sg13g2_decap_8 FILLER_37_832 ();
 sg13g2_decap_8 FILLER_37_839 ();
 sg13g2_decap_8 FILLER_37_846 ();
 sg13g2_decap_8 FILLER_37_853 ();
 sg13g2_fill_2 FILLER_37_860 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_4 FILLER_38_119 ();
 sg13g2_fill_2 FILLER_38_123 ();
 sg13g2_fill_2 FILLER_38_151 ();
 sg13g2_fill_2 FILLER_38_164 ();
 sg13g2_fill_1 FILLER_38_166 ();
 sg13g2_fill_2 FILLER_38_177 ();
 sg13g2_fill_1 FILLER_38_214 ();
 sg13g2_decap_4 FILLER_38_237 ();
 sg13g2_fill_2 FILLER_38_262 ();
 sg13g2_fill_1 FILLER_38_264 ();
 sg13g2_decap_4 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_321 ();
 sg13g2_decap_4 FILLER_38_326 ();
 sg13g2_fill_1 FILLER_38_330 ();
 sg13g2_fill_2 FILLER_38_341 ();
 sg13g2_fill_1 FILLER_38_357 ();
 sg13g2_fill_1 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_383 ();
 sg13g2_decap_4 FILLER_38_390 ();
 sg13g2_fill_1 FILLER_38_394 ();
 sg13g2_fill_1 FILLER_38_399 ();
 sg13g2_fill_2 FILLER_38_441 ();
 sg13g2_fill_2 FILLER_38_448 ();
 sg13g2_fill_1 FILLER_38_450 ();
 sg13g2_fill_1 FILLER_38_455 ();
 sg13g2_decap_8 FILLER_38_477 ();
 sg13g2_decap_4 FILLER_38_484 ();
 sg13g2_fill_1 FILLER_38_488 ();
 sg13g2_fill_2 FILLER_38_526 ();
 sg13g2_decap_4 FILLER_38_538 ();
 sg13g2_fill_1 FILLER_38_581 ();
 sg13g2_fill_2 FILLER_38_598 ();
 sg13g2_fill_1 FILLER_38_607 ();
 sg13g2_decap_4 FILLER_38_632 ();
 sg13g2_fill_2 FILLER_38_636 ();
 sg13g2_decap_8 FILLER_38_664 ();
 sg13g2_decap_4 FILLER_38_706 ();
 sg13g2_fill_2 FILLER_38_710 ();
 sg13g2_decap_8 FILLER_38_716 ();
 sg13g2_decap_8 FILLER_38_723 ();
 sg13g2_decap_8 FILLER_38_730 ();
 sg13g2_decap_8 FILLER_38_737 ();
 sg13g2_decap_8 FILLER_38_744 ();
 sg13g2_decap_8 FILLER_38_751 ();
 sg13g2_decap_8 FILLER_38_758 ();
 sg13g2_decap_8 FILLER_38_765 ();
 sg13g2_decap_8 FILLER_38_772 ();
 sg13g2_decap_8 FILLER_38_779 ();
 sg13g2_decap_8 FILLER_38_786 ();
 sg13g2_decap_8 FILLER_38_793 ();
 sg13g2_decap_8 FILLER_38_800 ();
 sg13g2_decap_8 FILLER_38_807 ();
 sg13g2_decap_8 FILLER_38_814 ();
 sg13g2_decap_8 FILLER_38_821 ();
 sg13g2_decap_8 FILLER_38_828 ();
 sg13g2_decap_8 FILLER_38_835 ();
 sg13g2_decap_8 FILLER_38_842 ();
 sg13g2_decap_8 FILLER_38_849 ();
 sg13g2_decap_4 FILLER_38_856 ();
 sg13g2_fill_2 FILLER_38_860 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_fill_2 FILLER_39_126 ();
 sg13g2_fill_1 FILLER_39_142 ();
 sg13g2_fill_2 FILLER_39_193 ();
 sg13g2_decap_8 FILLER_39_240 ();
 sg13g2_decap_8 FILLER_39_247 ();
 sg13g2_decap_4 FILLER_39_284 ();
 sg13g2_fill_2 FILLER_39_288 ();
 sg13g2_fill_2 FILLER_39_332 ();
 sg13g2_fill_1 FILLER_39_334 ();
 sg13g2_fill_2 FILLER_39_361 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_fill_2 FILLER_39_422 ();
 sg13g2_decap_4 FILLER_39_431 ();
 sg13g2_decap_4 FILLER_39_444 ();
 sg13g2_fill_1 FILLER_39_448 ();
 sg13g2_decap_8 FILLER_39_462 ();
 sg13g2_fill_1 FILLER_39_469 ();
 sg13g2_fill_2 FILLER_39_567 ();
 sg13g2_fill_2 FILLER_39_583 ();
 sg13g2_decap_8 FILLER_39_618 ();
 sg13g2_fill_1 FILLER_39_625 ();
 sg13g2_decap_8 FILLER_39_630 ();
 sg13g2_decap_8 FILLER_39_637 ();
 sg13g2_fill_1 FILLER_39_648 ();
 sg13g2_decap_8 FILLER_39_653 ();
 sg13g2_decap_4 FILLER_39_673 ();
 sg13g2_fill_1 FILLER_39_677 ();
 sg13g2_decap_4 FILLER_39_682 ();
 sg13g2_fill_2 FILLER_39_686 ();
 sg13g2_decap_8 FILLER_39_696 ();
 sg13g2_decap_8 FILLER_39_703 ();
 sg13g2_decap_8 FILLER_39_710 ();
 sg13g2_decap_8 FILLER_39_717 ();
 sg13g2_decap_8 FILLER_39_724 ();
 sg13g2_decap_8 FILLER_39_731 ();
 sg13g2_decap_8 FILLER_39_738 ();
 sg13g2_decap_8 FILLER_39_745 ();
 sg13g2_decap_8 FILLER_39_752 ();
 sg13g2_decap_8 FILLER_39_759 ();
 sg13g2_decap_8 FILLER_39_766 ();
 sg13g2_decap_8 FILLER_39_773 ();
 sg13g2_decap_8 FILLER_39_780 ();
 sg13g2_decap_8 FILLER_39_787 ();
 sg13g2_decap_8 FILLER_39_794 ();
 sg13g2_decap_8 FILLER_39_801 ();
 sg13g2_decap_8 FILLER_39_808 ();
 sg13g2_decap_8 FILLER_39_815 ();
 sg13g2_decap_8 FILLER_39_822 ();
 sg13g2_decap_8 FILLER_39_829 ();
 sg13g2_decap_8 FILLER_39_836 ();
 sg13g2_decap_8 FILLER_39_843 ();
 sg13g2_decap_8 FILLER_39_850 ();
 sg13g2_decap_4 FILLER_39_857 ();
 sg13g2_fill_1 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_fill_2 FILLER_40_126 ();
 sg13g2_fill_1 FILLER_40_128 ();
 sg13g2_fill_1 FILLER_40_143 ();
 sg13g2_decap_4 FILLER_40_154 ();
 sg13g2_fill_2 FILLER_40_204 ();
 sg13g2_decap_4 FILLER_40_242 ();
 sg13g2_fill_2 FILLER_40_273 ();
 sg13g2_fill_2 FILLER_40_301 ();
 sg13g2_decap_8 FILLER_40_316 ();
 sg13g2_decap_8 FILLER_40_323 ();
 sg13g2_fill_1 FILLER_40_330 ();
 sg13g2_fill_2 FILLER_40_344 ();
 sg13g2_decap_4 FILLER_40_356 ();
 sg13g2_fill_2 FILLER_40_360 ();
 sg13g2_fill_1 FILLER_40_367 ();
 sg13g2_decap_8 FILLER_40_375 ();
 sg13g2_decap_8 FILLER_40_382 ();
 sg13g2_decap_4 FILLER_40_389 ();
 sg13g2_fill_2 FILLER_40_393 ();
 sg13g2_decap_8 FILLER_40_408 ();
 sg13g2_fill_2 FILLER_40_415 ();
 sg13g2_fill_1 FILLER_40_422 ();
 sg13g2_decap_4 FILLER_40_517 ();
 sg13g2_fill_1 FILLER_40_521 ();
 sg13g2_fill_1 FILLER_40_541 ();
 sg13g2_decap_4 FILLER_40_578 ();
 sg13g2_fill_2 FILLER_40_582 ();
 sg13g2_fill_2 FILLER_40_597 ();
 sg13g2_fill_1 FILLER_40_599 ();
 sg13g2_fill_2 FILLER_40_608 ();
 sg13g2_fill_1 FILLER_40_610 ();
 sg13g2_decap_4 FILLER_40_632 ();
 sg13g2_fill_2 FILLER_40_665 ();
 sg13g2_decap_8 FILLER_40_706 ();
 sg13g2_decap_8 FILLER_40_713 ();
 sg13g2_decap_8 FILLER_40_720 ();
 sg13g2_decap_8 FILLER_40_727 ();
 sg13g2_decap_8 FILLER_40_734 ();
 sg13g2_decap_8 FILLER_40_741 ();
 sg13g2_decap_8 FILLER_40_748 ();
 sg13g2_decap_8 FILLER_40_755 ();
 sg13g2_decap_8 FILLER_40_762 ();
 sg13g2_decap_8 FILLER_40_769 ();
 sg13g2_decap_8 FILLER_40_776 ();
 sg13g2_decap_8 FILLER_40_783 ();
 sg13g2_decap_8 FILLER_40_790 ();
 sg13g2_decap_8 FILLER_40_797 ();
 sg13g2_decap_8 FILLER_40_804 ();
 sg13g2_decap_8 FILLER_40_811 ();
 sg13g2_decap_8 FILLER_40_818 ();
 sg13g2_decap_8 FILLER_40_825 ();
 sg13g2_decap_8 FILLER_40_832 ();
 sg13g2_decap_8 FILLER_40_839 ();
 sg13g2_decap_8 FILLER_40_846 ();
 sg13g2_decap_8 FILLER_40_853 ();
 sg13g2_fill_2 FILLER_40_860 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_fill_2 FILLER_41_77 ();
 sg13g2_fill_1 FILLER_41_105 ();
 sg13g2_fill_2 FILLER_41_115 ();
 sg13g2_fill_1 FILLER_41_117 ();
 sg13g2_decap_4 FILLER_41_144 ();
 sg13g2_fill_2 FILLER_41_148 ();
 sg13g2_decap_8 FILLER_41_176 ();
 sg13g2_fill_1 FILLER_41_219 ();
 sg13g2_fill_1 FILLER_41_225 ();
 sg13g2_fill_1 FILLER_41_235 ();
 sg13g2_fill_1 FILLER_41_246 ();
 sg13g2_decap_4 FILLER_41_277 ();
 sg13g2_decap_4 FILLER_41_294 ();
 sg13g2_decap_8 FILLER_41_410 ();
 sg13g2_decap_8 FILLER_41_417 ();
 sg13g2_decap_8 FILLER_41_424 ();
 sg13g2_fill_2 FILLER_41_431 ();
 sg13g2_fill_2 FILLER_41_448 ();
 sg13g2_fill_1 FILLER_41_450 ();
 sg13g2_fill_2 FILLER_41_471 ();
 sg13g2_decap_8 FILLER_41_539 ();
 sg13g2_decap_4 FILLER_41_546 ();
 sg13g2_decap_4 FILLER_41_575 ();
 sg13g2_fill_2 FILLER_41_579 ();
 sg13g2_decap_4 FILLER_41_601 ();
 sg13g2_fill_1 FILLER_41_605 ();
 sg13g2_decap_4 FILLER_41_619 ();
 sg13g2_fill_2 FILLER_41_623 ();
 sg13g2_decap_4 FILLER_41_629 ();
 sg13g2_decap_8 FILLER_41_676 ();
 sg13g2_decap_4 FILLER_41_683 ();
 sg13g2_decap_4 FILLER_41_692 ();
 sg13g2_decap_8 FILLER_41_704 ();
 sg13g2_decap_8 FILLER_41_711 ();
 sg13g2_decap_8 FILLER_41_718 ();
 sg13g2_decap_8 FILLER_41_725 ();
 sg13g2_decap_8 FILLER_41_732 ();
 sg13g2_decap_8 FILLER_41_739 ();
 sg13g2_decap_8 FILLER_41_746 ();
 sg13g2_decap_8 FILLER_41_753 ();
 sg13g2_decap_8 FILLER_41_760 ();
 sg13g2_decap_8 FILLER_41_767 ();
 sg13g2_decap_8 FILLER_41_774 ();
 sg13g2_decap_8 FILLER_41_781 ();
 sg13g2_decap_8 FILLER_41_788 ();
 sg13g2_decap_8 FILLER_41_795 ();
 sg13g2_decap_8 FILLER_41_802 ();
 sg13g2_decap_8 FILLER_41_809 ();
 sg13g2_decap_8 FILLER_41_816 ();
 sg13g2_decap_8 FILLER_41_823 ();
 sg13g2_decap_8 FILLER_41_830 ();
 sg13g2_decap_8 FILLER_41_837 ();
 sg13g2_decap_8 FILLER_41_844 ();
 sg13g2_decap_8 FILLER_41_851 ();
 sg13g2_decap_4 FILLER_41_858 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_fill_1 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_71 ();
 sg13g2_decap_4 FILLER_42_78 ();
 sg13g2_fill_1 FILLER_42_82 ();
 sg13g2_fill_1 FILLER_42_87 ();
 sg13g2_decap_8 FILLER_42_122 ();
 sg13g2_decap_8 FILLER_42_129 ();
 sg13g2_decap_4 FILLER_42_136 ();
 sg13g2_fill_1 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_150 ();
 sg13g2_decap_8 FILLER_42_157 ();
 sg13g2_fill_1 FILLER_42_164 ();
 sg13g2_decap_4 FILLER_42_170 ();
 sg13g2_fill_1 FILLER_42_182 ();
 sg13g2_fill_2 FILLER_42_188 ();
 sg13g2_fill_1 FILLER_42_190 ();
 sg13g2_fill_2 FILLER_42_236 ();
 sg13g2_fill_2 FILLER_42_269 ();
 sg13g2_fill_1 FILLER_42_271 ();
 sg13g2_fill_2 FILLER_42_309 ();
 sg13g2_fill_1 FILLER_42_311 ();
 sg13g2_decap_8 FILLER_42_343 ();
 sg13g2_decap_4 FILLER_42_350 ();
 sg13g2_fill_2 FILLER_42_366 ();
 sg13g2_fill_2 FILLER_42_385 ();
 sg13g2_decap_4 FILLER_42_391 ();
 sg13g2_decap_4 FILLER_42_420 ();
 sg13g2_fill_2 FILLER_42_424 ();
 sg13g2_fill_2 FILLER_42_434 ();
 sg13g2_fill_1 FILLER_42_436 ();
 sg13g2_decap_8 FILLER_42_479 ();
 sg13g2_decap_8 FILLER_42_486 ();
 sg13g2_fill_1 FILLER_42_493 ();
 sg13g2_decap_8 FILLER_42_498 ();
 sg13g2_decap_4 FILLER_42_505 ();
 sg13g2_fill_1 FILLER_42_509 ();
 sg13g2_fill_2 FILLER_42_519 ();
 sg13g2_decap_8 FILLER_42_537 ();
 sg13g2_fill_2 FILLER_42_544 ();
 sg13g2_decap_8 FILLER_42_566 ();
 sg13g2_decap_8 FILLER_42_573 ();
 sg13g2_fill_2 FILLER_42_580 ();
 sg13g2_fill_1 FILLER_42_589 ();
 sg13g2_fill_2 FILLER_42_607 ();
 sg13g2_fill_1 FILLER_42_609 ();
 sg13g2_fill_1 FILLER_42_622 ();
 sg13g2_fill_2 FILLER_42_653 ();
 sg13g2_fill_1 FILLER_42_655 ();
 sg13g2_fill_2 FILLER_42_688 ();
 sg13g2_fill_1 FILLER_42_690 ();
 sg13g2_decap_8 FILLER_42_717 ();
 sg13g2_decap_8 FILLER_42_724 ();
 sg13g2_decap_8 FILLER_42_731 ();
 sg13g2_decap_8 FILLER_42_738 ();
 sg13g2_decap_8 FILLER_42_745 ();
 sg13g2_decap_8 FILLER_42_752 ();
 sg13g2_decap_8 FILLER_42_759 ();
 sg13g2_decap_8 FILLER_42_766 ();
 sg13g2_decap_8 FILLER_42_773 ();
 sg13g2_decap_8 FILLER_42_780 ();
 sg13g2_decap_8 FILLER_42_787 ();
 sg13g2_decap_8 FILLER_42_794 ();
 sg13g2_decap_8 FILLER_42_801 ();
 sg13g2_decap_8 FILLER_42_808 ();
 sg13g2_decap_8 FILLER_42_815 ();
 sg13g2_decap_8 FILLER_42_822 ();
 sg13g2_decap_8 FILLER_42_829 ();
 sg13g2_decap_8 FILLER_42_836 ();
 sg13g2_decap_8 FILLER_42_843 ();
 sg13g2_decap_8 FILLER_42_850 ();
 sg13g2_decap_4 FILLER_42_857 ();
 sg13g2_fill_1 FILLER_42_861 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_fill_2 FILLER_43_28 ();
 sg13g2_fill_1 FILLER_43_34 ();
 sg13g2_decap_4 FILLER_43_44 ();
 sg13g2_fill_1 FILLER_43_48 ();
 sg13g2_fill_2 FILLER_43_89 ();
 sg13g2_fill_1 FILLER_43_91 ();
 sg13g2_fill_2 FILLER_43_178 ();
 sg13g2_decap_4 FILLER_43_193 ();
 sg13g2_fill_1 FILLER_43_197 ();
 sg13g2_fill_1 FILLER_43_237 ();
 sg13g2_decap_8 FILLER_43_264 ();
 sg13g2_decap_8 FILLER_43_271 ();
 sg13g2_fill_2 FILLER_43_278 ();
 sg13g2_fill_1 FILLER_43_280 ();
 sg13g2_fill_1 FILLER_43_298 ();
 sg13g2_fill_2 FILLER_43_304 ();
 sg13g2_fill_1 FILLER_43_306 ();
 sg13g2_fill_1 FILLER_43_319 ();
 sg13g2_fill_2 FILLER_43_325 ();
 sg13g2_fill_1 FILLER_43_327 ();
 sg13g2_fill_2 FILLER_43_332 ();
 sg13g2_decap_4 FILLER_43_360 ();
 sg13g2_fill_1 FILLER_43_364 ();
 sg13g2_decap_8 FILLER_43_396 ();
 sg13g2_fill_2 FILLER_43_403 ();
 sg13g2_fill_1 FILLER_43_405 ();
 sg13g2_decap_8 FILLER_43_444 ();
 sg13g2_decap_4 FILLER_43_456 ();
 sg13g2_fill_2 FILLER_43_467 ();
 sg13g2_decap_4 FILLER_43_494 ();
 sg13g2_fill_1 FILLER_43_517 ();
 sg13g2_decap_4 FILLER_43_544 ();
 sg13g2_fill_2 FILLER_43_548 ();
 sg13g2_fill_1 FILLER_43_555 ();
 sg13g2_decap_8 FILLER_43_569 ();
 sg13g2_decap_4 FILLER_43_581 ();
 sg13g2_fill_1 FILLER_43_585 ();
 sg13g2_fill_2 FILLER_43_594 ();
 sg13g2_fill_1 FILLER_43_596 ();
 sg13g2_decap_4 FILLER_43_628 ();
 sg13g2_fill_2 FILLER_43_632 ();
 sg13g2_decap_8 FILLER_43_638 ();
 sg13g2_decap_4 FILLER_43_645 ();
 sg13g2_fill_2 FILLER_43_649 ();
 sg13g2_decap_4 FILLER_43_669 ();
 sg13g2_decap_8 FILLER_43_677 ();
 sg13g2_decap_8 FILLER_43_684 ();
 sg13g2_decap_4 FILLER_43_691 ();
 sg13g2_fill_1 FILLER_43_695 ();
 sg13g2_decap_8 FILLER_43_713 ();
 sg13g2_decap_8 FILLER_43_720 ();
 sg13g2_decap_8 FILLER_43_727 ();
 sg13g2_decap_8 FILLER_43_734 ();
 sg13g2_decap_8 FILLER_43_741 ();
 sg13g2_decap_8 FILLER_43_748 ();
 sg13g2_decap_8 FILLER_43_755 ();
 sg13g2_decap_8 FILLER_43_762 ();
 sg13g2_decap_8 FILLER_43_769 ();
 sg13g2_decap_8 FILLER_43_776 ();
 sg13g2_decap_8 FILLER_43_783 ();
 sg13g2_decap_8 FILLER_43_790 ();
 sg13g2_decap_8 FILLER_43_797 ();
 sg13g2_decap_8 FILLER_43_804 ();
 sg13g2_decap_8 FILLER_43_811 ();
 sg13g2_decap_8 FILLER_43_818 ();
 sg13g2_decap_8 FILLER_43_825 ();
 sg13g2_decap_8 FILLER_43_832 ();
 sg13g2_decap_8 FILLER_43_839 ();
 sg13g2_decap_8 FILLER_43_846 ();
 sg13g2_decap_8 FILLER_43_853 ();
 sg13g2_fill_2 FILLER_43_860 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_4 FILLER_44_14 ();
 sg13g2_fill_1 FILLER_44_18 ();
 sg13g2_fill_2 FILLER_44_55 ();
 sg13g2_fill_1 FILLER_44_57 ();
 sg13g2_decap_4 FILLER_44_68 ();
 sg13g2_fill_2 FILLER_44_134 ();
 sg13g2_fill_1 FILLER_44_151 ();
 sg13g2_decap_8 FILLER_44_175 ();
 sg13g2_decap_8 FILLER_44_182 ();
 sg13g2_decap_4 FILLER_44_189 ();
 sg13g2_fill_2 FILLER_44_193 ();
 sg13g2_fill_2 FILLER_44_205 ();
 sg13g2_fill_1 FILLER_44_207 ();
 sg13g2_fill_2 FILLER_44_221 ();
 sg13g2_fill_1 FILLER_44_223 ();
 sg13g2_fill_1 FILLER_44_228 ();
 sg13g2_fill_2 FILLER_44_248 ();
 sg13g2_decap_4 FILLER_44_308 ();
 sg13g2_fill_2 FILLER_44_333 ();
 sg13g2_decap_4 FILLER_44_340 ();
 sg13g2_fill_1 FILLER_44_344 ();
 sg13g2_decap_8 FILLER_44_349 ();
 sg13g2_fill_2 FILLER_44_356 ();
 sg13g2_fill_1 FILLER_44_358 ();
 sg13g2_fill_2 FILLER_44_375 ();
 sg13g2_fill_2 FILLER_44_382 ();
 sg13g2_decap_8 FILLER_44_418 ();
 sg13g2_fill_2 FILLER_44_429 ();
 sg13g2_fill_1 FILLER_44_431 ();
 sg13g2_fill_1 FILLER_44_447 ();
 sg13g2_decap_4 FILLER_44_460 ();
 sg13g2_fill_2 FILLER_44_464 ();
 sg13g2_fill_2 FILLER_44_487 ();
 sg13g2_fill_1 FILLER_44_489 ();
 sg13g2_decap_4 FILLER_44_511 ();
 sg13g2_decap_8 FILLER_44_538 ();
 sg13g2_fill_1 FILLER_44_548 ();
 sg13g2_decap_8 FILLER_44_586 ();
 sg13g2_fill_1 FILLER_44_612 ();
 sg13g2_decap_4 FILLER_44_617 ();
 sg13g2_fill_2 FILLER_44_621 ();
 sg13g2_fill_1 FILLER_44_636 ();
 sg13g2_fill_1 FILLER_44_666 ();
 sg13g2_decap_8 FILLER_44_672 ();
 sg13g2_decap_8 FILLER_44_679 ();
 sg13g2_fill_2 FILLER_44_686 ();
 sg13g2_fill_1 FILLER_44_688 ();
 sg13g2_decap_8 FILLER_44_726 ();
 sg13g2_decap_8 FILLER_44_733 ();
 sg13g2_decap_8 FILLER_44_740 ();
 sg13g2_decap_8 FILLER_44_747 ();
 sg13g2_decap_8 FILLER_44_754 ();
 sg13g2_decap_8 FILLER_44_761 ();
 sg13g2_decap_8 FILLER_44_768 ();
 sg13g2_decap_8 FILLER_44_775 ();
 sg13g2_decap_8 FILLER_44_782 ();
 sg13g2_decap_8 FILLER_44_789 ();
 sg13g2_decap_8 FILLER_44_796 ();
 sg13g2_decap_8 FILLER_44_803 ();
 sg13g2_decap_8 FILLER_44_810 ();
 sg13g2_decap_8 FILLER_44_817 ();
 sg13g2_decap_8 FILLER_44_824 ();
 sg13g2_decap_8 FILLER_44_831 ();
 sg13g2_decap_8 FILLER_44_838 ();
 sg13g2_decap_8 FILLER_44_845 ();
 sg13g2_decap_8 FILLER_44_852 ();
 sg13g2_fill_2 FILLER_44_859 ();
 sg13g2_fill_1 FILLER_44_861 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_fill_2 FILLER_45_54 ();
 sg13g2_fill_1 FILLER_45_56 ();
 sg13g2_fill_2 FILLER_45_88 ();
 sg13g2_fill_2 FILLER_45_100 ();
 sg13g2_fill_2 FILLER_45_125 ();
 sg13g2_fill_1 FILLER_45_127 ();
 sg13g2_fill_2 FILLER_45_226 ();
 sg13g2_fill_1 FILLER_45_228 ();
 sg13g2_fill_2 FILLER_45_270 ();
 sg13g2_decap_8 FILLER_45_277 ();
 sg13g2_fill_2 FILLER_45_284 ();
 sg13g2_fill_1 FILLER_45_286 ();
 sg13g2_fill_2 FILLER_45_318 ();
 sg13g2_fill_1 FILLER_45_329 ();
 sg13g2_fill_1 FILLER_45_348 ();
 sg13g2_decap_8 FILLER_45_389 ();
 sg13g2_fill_1 FILLER_45_396 ();
 sg13g2_fill_2 FILLER_45_405 ();
 sg13g2_fill_2 FILLER_45_415 ();
 sg13g2_fill_1 FILLER_45_417 ();
 sg13g2_fill_2 FILLER_45_438 ();
 sg13g2_fill_1 FILLER_45_440 ();
 sg13g2_decap_4 FILLER_45_446 ();
 sg13g2_fill_1 FILLER_45_450 ();
 sg13g2_decap_8 FILLER_45_455 ();
 sg13g2_fill_2 FILLER_45_462 ();
 sg13g2_fill_1 FILLER_45_464 ();
 sg13g2_decap_8 FILLER_45_486 ();
 sg13g2_fill_1 FILLER_45_498 ();
 sg13g2_decap_4 FILLER_45_510 ();
 sg13g2_decap_8 FILLER_45_538 ();
 sg13g2_fill_1 FILLER_45_584 ();
 sg13g2_decap_8 FILLER_45_603 ();
 sg13g2_decap_8 FILLER_45_610 ();
 sg13g2_decap_8 FILLER_45_617 ();
 sg13g2_decap_8 FILLER_45_637 ();
 sg13g2_fill_2 FILLER_45_644 ();
 sg13g2_decap_8 FILLER_45_655 ();
 sg13g2_decap_8 FILLER_45_678 ();
 sg13g2_fill_2 FILLER_45_685 ();
 sg13g2_fill_1 FILLER_45_695 ();
 sg13g2_fill_1 FILLER_45_712 ();
 sg13g2_decap_8 FILLER_45_733 ();
 sg13g2_decap_8 FILLER_45_740 ();
 sg13g2_decap_8 FILLER_45_747 ();
 sg13g2_decap_8 FILLER_45_754 ();
 sg13g2_decap_8 FILLER_45_761 ();
 sg13g2_decap_8 FILLER_45_768 ();
 sg13g2_decap_8 FILLER_45_775 ();
 sg13g2_decap_8 FILLER_45_782 ();
 sg13g2_decap_8 FILLER_45_789 ();
 sg13g2_decap_8 FILLER_45_796 ();
 sg13g2_decap_8 FILLER_45_803 ();
 sg13g2_decap_8 FILLER_45_810 ();
 sg13g2_decap_8 FILLER_45_817 ();
 sg13g2_decap_8 FILLER_45_824 ();
 sg13g2_decap_8 FILLER_45_831 ();
 sg13g2_decap_8 FILLER_45_838 ();
 sg13g2_decap_8 FILLER_45_845 ();
 sg13g2_decap_8 FILLER_45_852 ();
 sg13g2_fill_2 FILLER_45_859 ();
 sg13g2_fill_1 FILLER_45_861 ();
 sg13g2_fill_2 FILLER_46_26 ();
 sg13g2_fill_1 FILLER_46_28 ();
 sg13g2_fill_2 FILLER_46_48 ();
 sg13g2_fill_2 FILLER_46_55 ();
 sg13g2_fill_1 FILLER_46_67 ();
 sg13g2_fill_1 FILLER_46_72 ();
 sg13g2_fill_1 FILLER_46_82 ();
 sg13g2_fill_1 FILLER_46_105 ();
 sg13g2_fill_1 FILLER_46_115 ();
 sg13g2_fill_2 FILLER_46_152 ();
 sg13g2_fill_2 FILLER_46_160 ();
 sg13g2_decap_4 FILLER_46_172 ();
 sg13g2_fill_2 FILLER_46_205 ();
 sg13g2_fill_2 FILLER_46_249 ();
 sg13g2_fill_1 FILLER_46_270 ();
 sg13g2_decap_4 FILLER_46_277 ();
 sg13g2_fill_2 FILLER_46_286 ();
 sg13g2_fill_2 FILLER_46_303 ();
 sg13g2_fill_2 FILLER_46_357 ();
 sg13g2_fill_1 FILLER_46_359 ();
 sg13g2_decap_8 FILLER_46_364 ();
 sg13g2_fill_1 FILLER_46_371 ();
 sg13g2_fill_2 FILLER_46_395 ();
 sg13g2_fill_1 FILLER_46_397 ();
 sg13g2_decap_4 FILLER_46_408 ();
 sg13g2_fill_2 FILLER_46_445 ();
 sg13g2_fill_1 FILLER_46_487 ();
 sg13g2_decap_8 FILLER_46_514 ();
 sg13g2_fill_2 FILLER_46_521 ();
 sg13g2_fill_1 FILLER_46_523 ();
 sg13g2_fill_2 FILLER_46_537 ();
 sg13g2_fill_1 FILLER_46_539 ();
 sg13g2_decap_4 FILLER_46_543 ();
 sg13g2_decap_4 FILLER_46_552 ();
 sg13g2_decap_8 FILLER_46_560 ();
 sg13g2_decap_8 FILLER_46_567 ();
 sg13g2_fill_1 FILLER_46_574 ();
 sg13g2_fill_2 FILLER_46_579 ();
 sg13g2_fill_1 FILLER_46_594 ();
 sg13g2_fill_2 FILLER_46_603 ();
 sg13g2_fill_1 FILLER_46_605 ();
 sg13g2_decap_8 FILLER_46_658 ();
 sg13g2_decap_4 FILLER_46_670 ();
 sg13g2_fill_2 FILLER_46_674 ();
 sg13g2_decap_8 FILLER_46_689 ();
 sg13g2_decap_8 FILLER_46_696 ();
 sg13g2_decap_8 FILLER_46_724 ();
 sg13g2_decap_8 FILLER_46_731 ();
 sg13g2_decap_8 FILLER_46_738 ();
 sg13g2_decap_8 FILLER_46_745 ();
 sg13g2_decap_8 FILLER_46_752 ();
 sg13g2_decap_8 FILLER_46_759 ();
 sg13g2_decap_8 FILLER_46_766 ();
 sg13g2_decap_8 FILLER_46_773 ();
 sg13g2_decap_8 FILLER_46_780 ();
 sg13g2_decap_8 FILLER_46_787 ();
 sg13g2_decap_8 FILLER_46_794 ();
 sg13g2_decap_8 FILLER_46_801 ();
 sg13g2_decap_8 FILLER_46_808 ();
 sg13g2_decap_8 FILLER_46_815 ();
 sg13g2_decap_8 FILLER_46_822 ();
 sg13g2_decap_8 FILLER_46_829 ();
 sg13g2_decap_8 FILLER_46_836 ();
 sg13g2_decap_8 FILLER_46_843 ();
 sg13g2_decap_8 FILLER_46_850 ();
 sg13g2_decap_4 FILLER_46_857 ();
 sg13g2_fill_1 FILLER_46_861 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_7 ();
 sg13g2_decap_4 FILLER_47_53 ();
 sg13g2_fill_1 FILLER_47_57 ();
 sg13g2_fill_2 FILLER_47_115 ();
 sg13g2_fill_1 FILLER_47_117 ();
 sg13g2_decap_4 FILLER_47_160 ();
 sg13g2_decap_8 FILLER_47_182 ();
 sg13g2_decap_8 FILLER_47_189 ();
 sg13g2_decap_4 FILLER_47_196 ();
 sg13g2_fill_2 FILLER_47_216 ();
 sg13g2_fill_2 FILLER_47_236 ();
 sg13g2_fill_1 FILLER_47_257 ();
 sg13g2_fill_2 FILLER_47_284 ();
 sg13g2_decap_4 FILLER_47_300 ();
 sg13g2_fill_2 FILLER_47_319 ();
 sg13g2_fill_1 FILLER_47_321 ();
 sg13g2_decap_4 FILLER_47_369 ();
 sg13g2_fill_2 FILLER_47_417 ();
 sg13g2_fill_1 FILLER_47_419 ();
 sg13g2_fill_2 FILLER_47_445 ();
 sg13g2_fill_1 FILLER_47_447 ();
 sg13g2_decap_8 FILLER_47_452 ();
 sg13g2_fill_2 FILLER_47_459 ();
 sg13g2_decap_4 FILLER_47_469 ();
 sg13g2_decap_8 FILLER_47_483 ();
 sg13g2_fill_2 FILLER_47_490 ();
 sg13g2_decap_4 FILLER_47_500 ();
 sg13g2_decap_4 FILLER_47_514 ();
 sg13g2_fill_1 FILLER_47_518 ();
 sg13g2_fill_2 FILLER_47_564 ();
 sg13g2_fill_2 FILLER_47_587 ();
 sg13g2_fill_2 FILLER_47_614 ();
 sg13g2_fill_1 FILLER_47_616 ();
 sg13g2_decap_8 FILLER_47_621 ();
 sg13g2_decap_8 FILLER_47_628 ();
 sg13g2_decap_4 FILLER_47_647 ();
 sg13g2_fill_2 FILLER_47_659 ();
 sg13g2_fill_2 FILLER_47_705 ();
 sg13g2_decap_8 FILLER_47_724 ();
 sg13g2_decap_8 FILLER_47_731 ();
 sg13g2_decap_8 FILLER_47_738 ();
 sg13g2_decap_8 FILLER_47_745 ();
 sg13g2_decap_8 FILLER_47_752 ();
 sg13g2_decap_8 FILLER_47_759 ();
 sg13g2_decap_8 FILLER_47_766 ();
 sg13g2_decap_8 FILLER_47_773 ();
 sg13g2_decap_8 FILLER_47_780 ();
 sg13g2_decap_8 FILLER_47_787 ();
 sg13g2_decap_8 FILLER_47_794 ();
 sg13g2_decap_8 FILLER_47_801 ();
 sg13g2_decap_8 FILLER_47_808 ();
 sg13g2_decap_8 FILLER_47_815 ();
 sg13g2_decap_8 FILLER_47_822 ();
 sg13g2_decap_8 FILLER_47_829 ();
 sg13g2_decap_8 FILLER_47_836 ();
 sg13g2_decap_8 FILLER_47_843 ();
 sg13g2_decap_8 FILLER_47_850 ();
 sg13g2_decap_4 FILLER_47_857 ();
 sg13g2_fill_1 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_fill_1 FILLER_48_14 ();
 sg13g2_fill_2 FILLER_48_37 ();
 sg13g2_fill_1 FILLER_48_47 ();
 sg13g2_decap_8 FILLER_48_53 ();
 sg13g2_decap_8 FILLER_48_60 ();
 sg13g2_fill_1 FILLER_48_67 ();
 sg13g2_fill_2 FILLER_48_118 ();
 sg13g2_decap_4 FILLER_48_156 ();
 sg13g2_fill_1 FILLER_48_168 ();
 sg13g2_fill_2 FILLER_48_183 ();
 sg13g2_fill_1 FILLER_48_185 ();
 sg13g2_decap_8 FILLER_48_197 ();
 sg13g2_fill_2 FILLER_48_204 ();
 sg13g2_fill_1 FILLER_48_206 ();
 sg13g2_fill_2 FILLER_48_261 ();
 sg13g2_fill_1 FILLER_48_263 ();
 sg13g2_decap_8 FILLER_48_279 ();
 sg13g2_decap_8 FILLER_48_299 ();
 sg13g2_decap_4 FILLER_48_306 ();
 sg13g2_fill_1 FILLER_48_330 ();
 sg13g2_decap_4 FILLER_48_348 ();
 sg13g2_fill_2 FILLER_48_352 ();
 sg13g2_decap_4 FILLER_48_358 ();
 sg13g2_fill_1 FILLER_48_362 ();
 sg13g2_decap_8 FILLER_48_383 ();
 sg13g2_decap_8 FILLER_48_390 ();
 sg13g2_fill_1 FILLER_48_397 ();
 sg13g2_fill_2 FILLER_48_403 ();
 sg13g2_decap_8 FILLER_48_409 ();
 sg13g2_decap_8 FILLER_48_416 ();
 sg13g2_decap_8 FILLER_48_423 ();
 sg13g2_decap_8 FILLER_48_438 ();
 sg13g2_decap_4 FILLER_48_445 ();
 sg13g2_fill_2 FILLER_48_453 ();
 sg13g2_decap_8 FILLER_48_480 ();
 sg13g2_fill_2 FILLER_48_487 ();
 sg13g2_fill_1 FILLER_48_489 ();
 sg13g2_decap_4 FILLER_48_503 ();
 sg13g2_fill_1 FILLER_48_524 ();
 sg13g2_decap_8 FILLER_48_537 ();
 sg13g2_decap_4 FILLER_48_544 ();
 sg13g2_fill_1 FILLER_48_548 ();
 sg13g2_decap_8 FILLER_48_569 ();
 sg13g2_decap_8 FILLER_48_576 ();
 sg13g2_decap_8 FILLER_48_583 ();
 sg13g2_fill_1 FILLER_48_590 ();
 sg13g2_decap_8 FILLER_48_608 ();
 sg13g2_decap_4 FILLER_48_615 ();
 sg13g2_fill_1 FILLER_48_619 ();
 sg13g2_decap_4 FILLER_48_646 ();
 sg13g2_fill_2 FILLER_48_667 ();
 sg13g2_decap_4 FILLER_48_674 ();
 sg13g2_fill_2 FILLER_48_678 ();
 sg13g2_decap_4 FILLER_48_689 ();
 sg13g2_fill_1 FILLER_48_693 ();
 sg13g2_fill_2 FILLER_48_711 ();
 sg13g2_fill_1 FILLER_48_713 ();
 sg13g2_decap_8 FILLER_48_722 ();
 sg13g2_decap_8 FILLER_48_729 ();
 sg13g2_decap_8 FILLER_48_736 ();
 sg13g2_decap_8 FILLER_48_743 ();
 sg13g2_decap_8 FILLER_48_750 ();
 sg13g2_decap_8 FILLER_48_757 ();
 sg13g2_decap_8 FILLER_48_764 ();
 sg13g2_decap_8 FILLER_48_771 ();
 sg13g2_decap_8 FILLER_48_778 ();
 sg13g2_decap_8 FILLER_48_785 ();
 sg13g2_decap_8 FILLER_48_792 ();
 sg13g2_decap_8 FILLER_48_799 ();
 sg13g2_decap_8 FILLER_48_806 ();
 sg13g2_decap_8 FILLER_48_813 ();
 sg13g2_decap_8 FILLER_48_820 ();
 sg13g2_decap_8 FILLER_48_827 ();
 sg13g2_decap_8 FILLER_48_834 ();
 sg13g2_decap_8 FILLER_48_841 ();
 sg13g2_decap_8 FILLER_48_848 ();
 sg13g2_decap_8 FILLER_48_855 ();
 sg13g2_fill_1 FILLER_49_0 ();
 sg13g2_decap_4 FILLER_49_27 ();
 sg13g2_fill_1 FILLER_49_31 ();
 sg13g2_fill_1 FILLER_49_67 ();
 sg13g2_fill_2 FILLER_49_83 ();
 sg13g2_fill_1 FILLER_49_130 ();
 sg13g2_fill_2 FILLER_49_135 ();
 sg13g2_fill_1 FILLER_49_171 ();
 sg13g2_decap_4 FILLER_49_177 ();
 sg13g2_fill_2 FILLER_49_229 ();
 sg13g2_fill_1 FILLER_49_231 ();
 sg13g2_fill_2 FILLER_49_240 ();
 sg13g2_decap_4 FILLER_49_263 ();
 sg13g2_fill_1 FILLER_49_267 ();
 sg13g2_fill_2 FILLER_49_280 ();
 sg13g2_fill_2 FILLER_49_295 ();
 sg13g2_fill_1 FILLER_49_297 ();
 sg13g2_decap_8 FILLER_49_303 ();
 sg13g2_decap_8 FILLER_49_310 ();
 sg13g2_fill_1 FILLER_49_317 ();
 sg13g2_fill_2 FILLER_49_326 ();
 sg13g2_fill_1 FILLER_49_328 ();
 sg13g2_decap_8 FILLER_49_342 ();
 sg13g2_decap_8 FILLER_49_349 ();
 sg13g2_fill_1 FILLER_49_356 ();
 sg13g2_decap_4 FILLER_49_360 ();
 sg13g2_fill_2 FILLER_49_364 ();
 sg13g2_fill_2 FILLER_49_376 ();
 sg13g2_fill_2 FILLER_49_382 ();
 sg13g2_fill_1 FILLER_49_384 ();
 sg13g2_decap_8 FILLER_49_415 ();
 sg13g2_fill_1 FILLER_49_422 ();
 sg13g2_fill_2 FILLER_49_436 ();
 sg13g2_fill_1 FILLER_49_438 ();
 sg13g2_fill_1 FILLER_49_465 ();
 sg13g2_decap_8 FILLER_49_500 ();
 sg13g2_decap_4 FILLER_49_507 ();
 sg13g2_fill_2 FILLER_49_511 ();
 sg13g2_decap_8 FILLER_49_521 ();
 sg13g2_decap_8 FILLER_49_541 ();
 sg13g2_fill_1 FILLER_49_548 ();
 sg13g2_decap_8 FILLER_49_575 ();
 sg13g2_fill_2 FILLER_49_582 ();
 sg13g2_fill_1 FILLER_49_584 ();
 sg13g2_fill_2 FILLER_49_598 ();
 sg13g2_decap_4 FILLER_49_626 ();
 sg13g2_fill_1 FILLER_49_630 ();
 sg13g2_fill_2 FILLER_49_635 ();
 sg13g2_decap_8 FILLER_49_658 ();
 sg13g2_decap_8 FILLER_49_665 ();
 sg13g2_decap_8 FILLER_49_676 ();
 sg13g2_decap_4 FILLER_49_683 ();
 sg13g2_decap_4 FILLER_49_700 ();
 sg13g2_fill_2 FILLER_49_704 ();
 sg13g2_decap_8 FILLER_49_731 ();
 sg13g2_decap_8 FILLER_49_738 ();
 sg13g2_decap_8 FILLER_49_745 ();
 sg13g2_decap_8 FILLER_49_752 ();
 sg13g2_decap_8 FILLER_49_759 ();
 sg13g2_decap_8 FILLER_49_766 ();
 sg13g2_decap_8 FILLER_49_773 ();
 sg13g2_decap_8 FILLER_49_780 ();
 sg13g2_decap_8 FILLER_49_787 ();
 sg13g2_decap_8 FILLER_49_794 ();
 sg13g2_decap_8 FILLER_49_801 ();
 sg13g2_decap_8 FILLER_49_808 ();
 sg13g2_decap_8 FILLER_49_815 ();
 sg13g2_decap_8 FILLER_49_822 ();
 sg13g2_decap_8 FILLER_49_829 ();
 sg13g2_decap_8 FILLER_49_836 ();
 sg13g2_decap_8 FILLER_49_843 ();
 sg13g2_decap_8 FILLER_49_850 ();
 sg13g2_decap_4 FILLER_49_857 ();
 sg13g2_fill_1 FILLER_49_861 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_4 FILLER_50_7 ();
 sg13g2_decap_4 FILLER_50_34 ();
 sg13g2_fill_1 FILLER_50_38 ();
 sg13g2_fill_2 FILLER_50_100 ();
 sg13g2_decap_8 FILLER_50_157 ();
 sg13g2_fill_1 FILLER_50_164 ();
 sg13g2_decap_8 FILLER_50_182 ();
 sg13g2_fill_1 FILLER_50_198 ();
 sg13g2_decap_8 FILLER_50_217 ();
 sg13g2_decap_8 FILLER_50_224 ();
 sg13g2_fill_2 FILLER_50_231 ();
 sg13g2_fill_1 FILLER_50_233 ();
 sg13g2_fill_2 FILLER_50_258 ();
 sg13g2_fill_1 FILLER_50_260 ();
 sg13g2_fill_2 FILLER_50_287 ();
 sg13g2_fill_1 FILLER_50_289 ();
 sg13g2_fill_1 FILLER_50_300 ();
 sg13g2_decap_8 FILLER_50_312 ();
 sg13g2_fill_1 FILLER_50_319 ();
 sg13g2_decap_8 FILLER_50_327 ();
 sg13g2_decap_8 FILLER_50_334 ();
 sg13g2_fill_1 FILLER_50_341 ();
 sg13g2_fill_2 FILLER_50_364 ();
 sg13g2_fill_1 FILLER_50_375 ();
 sg13g2_fill_2 FILLER_50_395 ();
 sg13g2_fill_1 FILLER_50_397 ();
 sg13g2_decap_4 FILLER_50_416 ();
 sg13g2_fill_1 FILLER_50_420 ();
 sg13g2_decap_8 FILLER_50_456 ();
 sg13g2_decap_8 FILLER_50_463 ();
 sg13g2_decap_8 FILLER_50_470 ();
 sg13g2_decap_4 FILLER_50_481 ();
 sg13g2_decap_8 FILLER_50_503 ();
 sg13g2_decap_8 FILLER_50_510 ();
 sg13g2_fill_1 FILLER_50_517 ();
 sg13g2_decap_8 FILLER_50_548 ();
 sg13g2_fill_2 FILLER_50_555 ();
 sg13g2_fill_1 FILLER_50_557 ();
 sg13g2_fill_1 FILLER_50_570 ();
 sg13g2_decap_4 FILLER_50_586 ();
 sg13g2_decap_4 FILLER_50_606 ();
 sg13g2_fill_1 FILLER_50_610 ();
 sg13g2_fill_2 FILLER_50_615 ();
 sg13g2_fill_2 FILLER_50_625 ();
 sg13g2_fill_1 FILLER_50_627 ();
 sg13g2_fill_2 FILLER_50_640 ();
 sg13g2_fill_2 FILLER_50_658 ();
 sg13g2_fill_1 FILLER_50_660 ();
 sg13g2_decap_4 FILLER_50_705 ();
 sg13g2_fill_1 FILLER_50_709 ();
 sg13g2_decap_8 FILLER_50_723 ();
 sg13g2_decap_8 FILLER_50_730 ();
 sg13g2_decap_8 FILLER_50_737 ();
 sg13g2_decap_8 FILLER_50_744 ();
 sg13g2_decap_8 FILLER_50_751 ();
 sg13g2_decap_8 FILLER_50_758 ();
 sg13g2_decap_8 FILLER_50_765 ();
 sg13g2_decap_8 FILLER_50_772 ();
 sg13g2_decap_8 FILLER_50_779 ();
 sg13g2_decap_8 FILLER_50_786 ();
 sg13g2_decap_8 FILLER_50_793 ();
 sg13g2_decap_8 FILLER_50_800 ();
 sg13g2_decap_8 FILLER_50_807 ();
 sg13g2_decap_8 FILLER_50_814 ();
 sg13g2_decap_8 FILLER_50_821 ();
 sg13g2_decap_8 FILLER_50_828 ();
 sg13g2_decap_8 FILLER_50_835 ();
 sg13g2_decap_8 FILLER_50_842 ();
 sg13g2_decap_8 FILLER_50_849 ();
 sg13g2_decap_4 FILLER_50_856 ();
 sg13g2_fill_2 FILLER_50_860 ();
 sg13g2_fill_1 FILLER_51_0 ();
 sg13g2_decap_4 FILLER_51_50 ();
 sg13g2_fill_1 FILLER_51_54 ();
 sg13g2_fill_2 FILLER_51_85 ();
 sg13g2_fill_2 FILLER_51_111 ();
 sg13g2_fill_2 FILLER_51_126 ();
 sg13g2_fill_1 FILLER_51_145 ();
 sg13g2_decap_8 FILLER_51_159 ();
 sg13g2_fill_2 FILLER_51_166 ();
 sg13g2_fill_1 FILLER_51_168 ();
 sg13g2_fill_1 FILLER_51_211 ();
 sg13g2_decap_4 FILLER_51_242 ();
 sg13g2_fill_1 FILLER_51_246 ();
 sg13g2_decap_4 FILLER_51_257 ();
 sg13g2_decap_8 FILLER_51_268 ();
 sg13g2_decap_8 FILLER_51_275 ();
 sg13g2_decap_8 FILLER_51_282 ();
 sg13g2_fill_2 FILLER_51_289 ();
 sg13g2_fill_1 FILLER_51_291 ();
 sg13g2_fill_1 FILLER_51_305 ();
 sg13g2_fill_2 FILLER_51_339 ();
 sg13g2_fill_1 FILLER_51_341 ();
 sg13g2_decap_4 FILLER_51_348 ();
 sg13g2_fill_2 FILLER_51_378 ();
 sg13g2_fill_1 FILLER_51_389 ();
 sg13g2_fill_2 FILLER_51_400 ();
 sg13g2_fill_1 FILLER_51_421 ();
 sg13g2_decap_4 FILLER_51_433 ();
 sg13g2_fill_1 FILLER_51_437 ();
 sg13g2_decap_4 FILLER_51_454 ();
 sg13g2_decap_8 FILLER_51_510 ();
 sg13g2_decap_4 FILLER_51_517 ();
 sg13g2_fill_1 FILLER_51_521 ();
 sg13g2_fill_1 FILLER_51_534 ();
 sg13g2_decap_4 FILLER_51_543 ();
 sg13g2_decap_8 FILLER_51_586 ();
 sg13g2_fill_1 FILLER_51_593 ();
 sg13g2_decap_8 FILLER_51_606 ();
 sg13g2_fill_1 FILLER_51_613 ();
 sg13g2_decap_8 FILLER_51_629 ();
 sg13g2_decap_4 FILLER_51_636 ();
 sg13g2_fill_2 FILLER_51_649 ();
 sg13g2_decap_8 FILLER_51_664 ();
 sg13g2_decap_8 FILLER_51_671 ();
 sg13g2_decap_4 FILLER_51_678 ();
 sg13g2_fill_1 FILLER_51_682 ();
 sg13g2_fill_2 FILLER_51_708 ();
 sg13g2_fill_2 FILLER_51_723 ();
 sg13g2_decap_8 FILLER_51_737 ();
 sg13g2_decap_8 FILLER_51_744 ();
 sg13g2_decap_8 FILLER_51_751 ();
 sg13g2_decap_8 FILLER_51_758 ();
 sg13g2_decap_8 FILLER_51_765 ();
 sg13g2_decap_8 FILLER_51_772 ();
 sg13g2_decap_8 FILLER_51_779 ();
 sg13g2_decap_8 FILLER_51_786 ();
 sg13g2_decap_8 FILLER_51_793 ();
 sg13g2_decap_8 FILLER_51_800 ();
 sg13g2_decap_8 FILLER_51_807 ();
 sg13g2_decap_8 FILLER_51_814 ();
 sg13g2_decap_8 FILLER_51_821 ();
 sg13g2_decap_8 FILLER_51_828 ();
 sg13g2_decap_8 FILLER_51_835 ();
 sg13g2_decap_8 FILLER_51_842 ();
 sg13g2_decap_8 FILLER_51_849 ();
 sg13g2_decap_4 FILLER_51_856 ();
 sg13g2_fill_2 FILLER_51_860 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_2 ();
 sg13g2_fill_2 FILLER_52_30 ();
 sg13g2_fill_1 FILLER_52_32 ();
 sg13g2_fill_1 FILLER_52_59 ();
 sg13g2_fill_2 FILLER_52_101 ();
 sg13g2_fill_1 FILLER_52_134 ();
 sg13g2_fill_2 FILLER_52_182 ();
 sg13g2_fill_1 FILLER_52_184 ();
 sg13g2_fill_2 FILLER_52_207 ();
 sg13g2_fill_1 FILLER_52_209 ();
 sg13g2_fill_1 FILLER_52_232 ();
 sg13g2_decap_4 FILLER_52_249 ();
 sg13g2_fill_1 FILLER_52_253 ();
 sg13g2_decap_8 FILLER_52_279 ();
 sg13g2_fill_1 FILLER_52_286 ();
 sg13g2_fill_2 FILLER_52_322 ();
 sg13g2_fill_2 FILLER_52_329 ();
 sg13g2_fill_1 FILLER_52_331 ();
 sg13g2_decap_8 FILLER_52_337 ();
 sg13g2_fill_1 FILLER_52_344 ();
 sg13g2_fill_1 FILLER_52_360 ();
 sg13g2_fill_2 FILLER_52_421 ();
 sg13g2_decap_8 FILLER_52_431 ();
 sg13g2_fill_1 FILLER_52_438 ();
 sg13g2_decap_4 FILLER_52_455 ();
 sg13g2_fill_1 FILLER_52_459 ();
 sg13g2_decap_4 FILLER_52_488 ();
 sg13g2_fill_1 FILLER_52_492 ();
 sg13g2_fill_2 FILLER_52_503 ();
 sg13g2_decap_8 FILLER_52_517 ();
 sg13g2_decap_8 FILLER_52_566 ();
 sg13g2_decap_8 FILLER_52_573 ();
 sg13g2_decap_4 FILLER_52_580 ();
 sg13g2_fill_2 FILLER_52_584 ();
 sg13g2_fill_2 FILLER_52_621 ();
 sg13g2_fill_1 FILLER_52_623 ();
 sg13g2_fill_2 FILLER_52_650 ();
 sg13g2_decap_8 FILLER_52_657 ();
 sg13g2_fill_1 FILLER_52_664 ();
 sg13g2_decap_8 FILLER_52_699 ();
 sg13g2_decap_8 FILLER_52_740 ();
 sg13g2_decap_8 FILLER_52_747 ();
 sg13g2_decap_8 FILLER_52_754 ();
 sg13g2_decap_8 FILLER_52_761 ();
 sg13g2_decap_8 FILLER_52_768 ();
 sg13g2_decap_8 FILLER_52_775 ();
 sg13g2_decap_8 FILLER_52_782 ();
 sg13g2_decap_8 FILLER_52_789 ();
 sg13g2_decap_8 FILLER_52_796 ();
 sg13g2_decap_8 FILLER_52_803 ();
 sg13g2_decap_8 FILLER_52_810 ();
 sg13g2_decap_8 FILLER_52_817 ();
 sg13g2_decap_8 FILLER_52_824 ();
 sg13g2_decap_8 FILLER_52_831 ();
 sg13g2_decap_8 FILLER_52_838 ();
 sg13g2_decap_8 FILLER_52_845 ();
 sg13g2_decap_8 FILLER_52_852 ();
 sg13g2_fill_2 FILLER_52_859 ();
 sg13g2_fill_1 FILLER_52_861 ();
 sg13g2_fill_2 FILLER_53_26 ();
 sg13g2_decap_4 FILLER_53_64 ();
 sg13g2_fill_2 FILLER_53_90 ();
 sg13g2_decap_4 FILLER_53_96 ();
 sg13g2_fill_1 FILLER_53_100 ();
 sg13g2_fill_2 FILLER_53_106 ();
 sg13g2_fill_2 FILLER_53_138 ();
 sg13g2_fill_2 FILLER_53_154 ();
 sg13g2_fill_1 FILLER_53_156 ();
 sg13g2_fill_1 FILLER_53_165 ();
 sg13g2_fill_2 FILLER_53_185 ();
 sg13g2_fill_1 FILLER_53_187 ();
 sg13g2_decap_8 FILLER_53_192 ();
 sg13g2_decap_4 FILLER_53_199 ();
 sg13g2_fill_2 FILLER_53_203 ();
 sg13g2_decap_8 FILLER_53_249 ();
 sg13g2_fill_2 FILLER_53_256 ();
 sg13g2_fill_1 FILLER_53_291 ();
 sg13g2_fill_2 FILLER_53_305 ();
 sg13g2_fill_1 FILLER_53_307 ();
 sg13g2_fill_2 FILLER_53_332 ();
 sg13g2_fill_1 FILLER_53_334 ();
 sg13g2_decap_4 FILLER_53_352 ();
 sg13g2_fill_1 FILLER_53_356 ();
 sg13g2_decap_8 FILLER_53_367 ();
 sg13g2_fill_2 FILLER_53_388 ();
 sg13g2_decap_8 FILLER_53_394 ();
 sg13g2_fill_1 FILLER_53_418 ();
 sg13g2_decap_4 FILLER_53_424 ();
 sg13g2_fill_1 FILLER_53_428 ();
 sg13g2_decap_8 FILLER_53_438 ();
 sg13g2_fill_1 FILLER_53_479 ();
 sg13g2_fill_2 FILLER_53_517 ();
 sg13g2_fill_1 FILLER_53_519 ();
 sg13g2_decap_8 FILLER_53_553 ();
 sg13g2_fill_2 FILLER_53_560 ();
 sg13g2_fill_1 FILLER_53_562 ();
 sg13g2_fill_2 FILLER_53_589 ();
 sg13g2_fill_1 FILLER_53_591 ();
 sg13g2_decap_8 FILLER_53_618 ();
 sg13g2_decap_4 FILLER_53_625 ();
 sg13g2_fill_2 FILLER_53_629 ();
 sg13g2_decap_4 FILLER_53_683 ();
 sg13g2_decap_8 FILLER_53_692 ();
 sg13g2_fill_2 FILLER_53_699 ();
 sg13g2_fill_1 FILLER_53_701 ();
 sg13g2_decap_8 FILLER_53_710 ();
 sg13g2_decap_4 FILLER_53_725 ();
 sg13g2_decap_8 FILLER_53_734 ();
 sg13g2_decap_8 FILLER_53_741 ();
 sg13g2_decap_8 FILLER_53_748 ();
 sg13g2_decap_8 FILLER_53_755 ();
 sg13g2_decap_8 FILLER_53_762 ();
 sg13g2_decap_8 FILLER_53_769 ();
 sg13g2_decap_8 FILLER_53_776 ();
 sg13g2_decap_8 FILLER_53_783 ();
 sg13g2_decap_8 FILLER_53_790 ();
 sg13g2_decap_8 FILLER_53_797 ();
 sg13g2_decap_8 FILLER_53_804 ();
 sg13g2_decap_8 FILLER_53_811 ();
 sg13g2_decap_8 FILLER_53_818 ();
 sg13g2_decap_8 FILLER_53_825 ();
 sg13g2_decap_8 FILLER_53_832 ();
 sg13g2_decap_8 FILLER_53_839 ();
 sg13g2_decap_8 FILLER_53_846 ();
 sg13g2_decap_8 FILLER_53_853 ();
 sg13g2_fill_2 FILLER_53_860 ();
 sg13g2_decap_4 FILLER_54_26 ();
 sg13g2_fill_1 FILLER_54_30 ();
 sg13g2_fill_2 FILLER_54_54 ();
 sg13g2_fill_1 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_83 ();
 sg13g2_decap_4 FILLER_54_90 ();
 sg13g2_fill_2 FILLER_54_166 ();
 sg13g2_decap_8 FILLER_54_204 ();
 sg13g2_fill_1 FILLER_54_211 ();
 sg13g2_decap_8 FILLER_54_239 ();
 sg13g2_decap_4 FILLER_54_246 ();
 sg13g2_decap_8 FILLER_54_277 ();
 sg13g2_fill_2 FILLER_54_290 ();
 sg13g2_fill_1 FILLER_54_292 ();
 sg13g2_decap_8 FILLER_54_298 ();
 sg13g2_decap_4 FILLER_54_305 ();
 sg13g2_fill_1 FILLER_54_309 ();
 sg13g2_decap_8 FILLER_54_336 ();
 sg13g2_decap_8 FILLER_54_343 ();
 sg13g2_fill_2 FILLER_54_350 ();
 sg13g2_fill_1 FILLER_54_445 ();
 sg13g2_decap_4 FILLER_54_456 ();
 sg13g2_fill_1 FILLER_54_486 ();
 sg13g2_fill_2 FILLER_54_514 ();
 sg13g2_fill_1 FILLER_54_516 ();
 sg13g2_fill_2 FILLER_54_542 ();
 sg13g2_fill_1 FILLER_54_544 ();
 sg13g2_fill_1 FILLER_54_565 ();
 sg13g2_fill_1 FILLER_54_582 ();
 sg13g2_decap_4 FILLER_54_597 ();
 sg13g2_fill_2 FILLER_54_601 ();
 sg13g2_decap_8 FILLER_54_607 ();
 sg13g2_fill_1 FILLER_54_614 ();
 sg13g2_fill_1 FILLER_54_624 ();
 sg13g2_fill_2 FILLER_54_639 ();
 sg13g2_decap_8 FILLER_54_645 ();
 sg13g2_decap_8 FILLER_54_652 ();
 sg13g2_decap_8 FILLER_54_659 ();
 sg13g2_fill_2 FILLER_54_666 ();
 sg13g2_fill_1 FILLER_54_668 ();
 sg13g2_decap_8 FILLER_54_682 ();
 sg13g2_decap_8 FILLER_54_689 ();
 sg13g2_fill_1 FILLER_54_696 ();
 sg13g2_decap_8 FILLER_54_744 ();
 sg13g2_decap_8 FILLER_54_751 ();
 sg13g2_decap_8 FILLER_54_758 ();
 sg13g2_decap_8 FILLER_54_765 ();
 sg13g2_decap_8 FILLER_54_772 ();
 sg13g2_decap_8 FILLER_54_779 ();
 sg13g2_decap_8 FILLER_54_786 ();
 sg13g2_decap_8 FILLER_54_793 ();
 sg13g2_decap_8 FILLER_54_800 ();
 sg13g2_decap_8 FILLER_54_807 ();
 sg13g2_decap_8 FILLER_54_814 ();
 sg13g2_decap_8 FILLER_54_821 ();
 sg13g2_decap_8 FILLER_54_828 ();
 sg13g2_decap_8 FILLER_54_835 ();
 sg13g2_decap_8 FILLER_54_842 ();
 sg13g2_decap_8 FILLER_54_849 ();
 sg13g2_decap_4 FILLER_54_856 ();
 sg13g2_fill_2 FILLER_54_860 ();
 sg13g2_fill_1 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_67 ();
 sg13g2_decap_8 FILLER_55_108 ();
 sg13g2_fill_2 FILLER_55_115 ();
 sg13g2_fill_1 FILLER_55_127 ();
 sg13g2_decap_4 FILLER_55_143 ();
 sg13g2_fill_2 FILLER_55_147 ();
 sg13g2_decap_4 FILLER_55_164 ();
 sg13g2_fill_2 FILLER_55_168 ();
 sg13g2_fill_2 FILLER_55_212 ();
 sg13g2_fill_1 FILLER_55_214 ();
 sg13g2_decap_8 FILLER_55_246 ();
 sg13g2_decap_8 FILLER_55_253 ();
 sg13g2_fill_1 FILLER_55_260 ();
 sg13g2_fill_2 FILLER_55_273 ();
 sg13g2_fill_1 FILLER_55_275 ();
 sg13g2_fill_2 FILLER_55_295 ();
 sg13g2_fill_2 FILLER_55_310 ();
 sg13g2_decap_8 FILLER_55_328 ();
 sg13g2_decap_4 FILLER_55_335 ();
 sg13g2_decap_4 FILLER_55_357 ();
 sg13g2_fill_1 FILLER_55_361 ();
 sg13g2_fill_2 FILLER_55_366 ();
 sg13g2_decap_4 FILLER_55_387 ();
 sg13g2_fill_2 FILLER_55_391 ();
 sg13g2_decap_4 FILLER_55_407 ();
 sg13g2_fill_2 FILLER_55_411 ();
 sg13g2_fill_2 FILLER_55_426 ();
 sg13g2_fill_1 FILLER_55_428 ();
 sg13g2_decap_8 FILLER_55_433 ();
 sg13g2_fill_1 FILLER_55_440 ();
 sg13g2_fill_2 FILLER_55_477 ();
 sg13g2_fill_1 FILLER_55_502 ();
 sg13g2_fill_2 FILLER_55_528 ();
 sg13g2_fill_1 FILLER_55_530 ();
 sg13g2_fill_1 FILLER_55_535 ();
 sg13g2_decap_8 FILLER_55_549 ();
 sg13g2_decap_4 FILLER_55_556 ();
 sg13g2_fill_2 FILLER_55_569 ();
 sg13g2_fill_2 FILLER_55_579 ();
 sg13g2_fill_1 FILLER_55_581 ();
 sg13g2_decap_8 FILLER_55_601 ();
 sg13g2_fill_1 FILLER_55_608 ();
 sg13g2_fill_2 FILLER_55_621 ();
 sg13g2_fill_1 FILLER_55_623 ();
 sg13g2_decap_4 FILLER_55_639 ();
 sg13g2_decap_8 FILLER_55_669 ();
 sg13g2_fill_2 FILLER_55_706 ();
 sg13g2_fill_1 FILLER_55_708 ();
 sg13g2_decap_8 FILLER_55_735 ();
 sg13g2_decap_8 FILLER_55_742 ();
 sg13g2_decap_8 FILLER_55_749 ();
 sg13g2_decap_8 FILLER_55_756 ();
 sg13g2_decap_8 FILLER_55_763 ();
 sg13g2_decap_8 FILLER_55_770 ();
 sg13g2_decap_8 FILLER_55_777 ();
 sg13g2_decap_8 FILLER_55_784 ();
 sg13g2_decap_8 FILLER_55_791 ();
 sg13g2_decap_8 FILLER_55_798 ();
 sg13g2_decap_8 FILLER_55_805 ();
 sg13g2_decap_8 FILLER_55_812 ();
 sg13g2_decap_8 FILLER_55_819 ();
 sg13g2_decap_8 FILLER_55_826 ();
 sg13g2_decap_8 FILLER_55_833 ();
 sg13g2_decap_8 FILLER_55_840 ();
 sg13g2_decap_8 FILLER_55_847 ();
 sg13g2_decap_8 FILLER_55_854 ();
 sg13g2_fill_1 FILLER_55_861 ();
 sg13g2_decap_4 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_4 ();
 sg13g2_fill_2 FILLER_56_30 ();
 sg13g2_fill_1 FILLER_56_32 ();
 sg13g2_fill_2 FILLER_56_42 ();
 sg13g2_fill_1 FILLER_56_44 ();
 sg13g2_decap_8 FILLER_56_68 ();
 sg13g2_fill_1 FILLER_56_75 ();
 sg13g2_decap_4 FILLER_56_85 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_4 FILLER_56_105 ();
 sg13g2_fill_1 FILLER_56_109 ();
 sg13g2_fill_2 FILLER_56_119 ();
 sg13g2_fill_2 FILLER_56_147 ();
 sg13g2_decap_4 FILLER_56_180 ();
 sg13g2_fill_2 FILLER_56_209 ();
 sg13g2_fill_2 FILLER_56_216 ();
 sg13g2_fill_1 FILLER_56_218 ();
 sg13g2_fill_2 FILLER_56_233 ();
 sg13g2_fill_1 FILLER_56_235 ();
 sg13g2_fill_1 FILLER_56_245 ();
 sg13g2_decap_4 FILLER_56_259 ();
 sg13g2_fill_1 FILLER_56_287 ();
 sg13g2_fill_1 FILLER_56_293 ();
 sg13g2_decap_8 FILLER_56_299 ();
 sg13g2_decap_4 FILLER_56_306 ();
 sg13g2_fill_1 FILLER_56_310 ();
 sg13g2_fill_1 FILLER_56_321 ();
 sg13g2_fill_2 FILLER_56_348 ();
 sg13g2_fill_1 FILLER_56_350 ();
 sg13g2_decap_4 FILLER_56_377 ();
 sg13g2_decap_8 FILLER_56_433 ();
 sg13g2_decap_4 FILLER_56_440 ();
 sg13g2_fill_2 FILLER_56_444 ();
 sg13g2_fill_1 FILLER_56_451 ();
 sg13g2_fill_1 FILLER_56_483 ();
 sg13g2_fill_2 FILLER_56_520 ();
 sg13g2_fill_1 FILLER_56_522 ();
 sg13g2_fill_1 FILLER_56_544 ();
 sg13g2_fill_2 FILLER_56_557 ();
 sg13g2_fill_1 FILLER_56_559 ();
 sg13g2_fill_2 FILLER_56_614 ();
 sg13g2_fill_1 FILLER_56_616 ();
 sg13g2_decap_8 FILLER_56_647 ();
 sg13g2_decap_8 FILLER_56_658 ();
 sg13g2_decap_8 FILLER_56_695 ();
 sg13g2_decap_8 FILLER_56_702 ();
 sg13g2_fill_2 FILLER_56_717 ();
 sg13g2_fill_1 FILLER_56_719 ();
 sg13g2_decap_8 FILLER_56_724 ();
 sg13g2_decap_8 FILLER_56_731 ();
 sg13g2_decap_8 FILLER_56_738 ();
 sg13g2_decap_8 FILLER_56_745 ();
 sg13g2_decap_8 FILLER_56_752 ();
 sg13g2_decap_8 FILLER_56_759 ();
 sg13g2_decap_8 FILLER_56_766 ();
 sg13g2_decap_8 FILLER_56_773 ();
 sg13g2_decap_8 FILLER_56_780 ();
 sg13g2_decap_8 FILLER_56_787 ();
 sg13g2_decap_8 FILLER_56_794 ();
 sg13g2_decap_8 FILLER_56_801 ();
 sg13g2_decap_8 FILLER_56_808 ();
 sg13g2_decap_8 FILLER_56_815 ();
 sg13g2_decap_8 FILLER_56_822 ();
 sg13g2_decap_8 FILLER_56_829 ();
 sg13g2_decap_8 FILLER_56_836 ();
 sg13g2_decap_8 FILLER_56_843 ();
 sg13g2_decap_8 FILLER_56_850 ();
 sg13g2_decap_4 FILLER_56_857 ();
 sg13g2_fill_1 FILLER_56_861 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_4 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_15 ();
 sg13g2_decap_4 FILLER_57_57 ();
 sg13g2_decap_8 FILLER_57_95 ();
 sg13g2_fill_1 FILLER_57_102 ();
 sg13g2_fill_2 FILLER_57_117 ();
 sg13g2_fill_2 FILLER_57_133 ();
 sg13g2_fill_1 FILLER_57_135 ();
 sg13g2_decap_4 FILLER_57_169 ();
 sg13g2_fill_2 FILLER_57_191 ();
 sg13g2_fill_1 FILLER_57_193 ();
 sg13g2_fill_2 FILLER_57_203 ();
 sg13g2_fill_1 FILLER_57_215 ();
 sg13g2_decap_8 FILLER_57_242 ();
 sg13g2_fill_1 FILLER_57_249 ();
 sg13g2_fill_2 FILLER_57_258 ();
 sg13g2_fill_1 FILLER_57_260 ();
 sg13g2_fill_2 FILLER_57_271 ();
 sg13g2_decap_4 FILLER_57_282 ();
 sg13g2_fill_1 FILLER_57_286 ();
 sg13g2_fill_1 FILLER_57_317 ();
 sg13g2_decap_4 FILLER_57_328 ();
 sg13g2_fill_1 FILLER_57_332 ();
 sg13g2_fill_1 FILLER_57_337 ();
 sg13g2_decap_8 FILLER_57_377 ();
 sg13g2_decap_4 FILLER_57_384 ();
 sg13g2_fill_1 FILLER_57_388 ();
 sg13g2_fill_1 FILLER_57_407 ();
 sg13g2_fill_1 FILLER_57_444 ();
 sg13g2_decap_4 FILLER_57_455 ();
 sg13g2_fill_1 FILLER_57_459 ();
 sg13g2_fill_2 FILLER_57_473 ();
 sg13g2_fill_1 FILLER_57_475 ();
 sg13g2_fill_2 FILLER_57_485 ();
 sg13g2_fill_1 FILLER_57_505 ();
 sg13g2_decap_4 FILLER_57_515 ();
 sg13g2_decap_8 FILLER_57_535 ();
 sg13g2_fill_2 FILLER_57_564 ();
 sg13g2_fill_1 FILLER_57_566 ();
 sg13g2_fill_2 FILLER_57_584 ();
 sg13g2_fill_1 FILLER_57_586 ();
 sg13g2_fill_1 FILLER_57_604 ();
 sg13g2_decap_8 FILLER_57_610 ();
 sg13g2_decap_4 FILLER_57_617 ();
 sg13g2_fill_1 FILLER_57_621 ();
 sg13g2_fill_2 FILLER_57_626 ();
 sg13g2_decap_4 FILLER_57_641 ();
 sg13g2_decap_8 FILLER_57_671 ();
 sg13g2_decap_4 FILLER_57_678 ();
 sg13g2_fill_1 FILLER_57_682 ();
 sg13g2_decap_4 FILLER_57_687 ();
 sg13g2_decap_8 FILLER_57_730 ();
 sg13g2_decap_8 FILLER_57_737 ();
 sg13g2_decap_8 FILLER_57_744 ();
 sg13g2_decap_8 FILLER_57_751 ();
 sg13g2_decap_8 FILLER_57_758 ();
 sg13g2_decap_8 FILLER_57_765 ();
 sg13g2_decap_8 FILLER_57_772 ();
 sg13g2_decap_8 FILLER_57_779 ();
 sg13g2_decap_8 FILLER_57_786 ();
 sg13g2_decap_8 FILLER_57_793 ();
 sg13g2_decap_8 FILLER_57_800 ();
 sg13g2_decap_8 FILLER_57_807 ();
 sg13g2_decap_8 FILLER_57_814 ();
 sg13g2_decap_8 FILLER_57_821 ();
 sg13g2_decap_8 FILLER_57_828 ();
 sg13g2_decap_8 FILLER_57_835 ();
 sg13g2_decap_8 FILLER_57_842 ();
 sg13g2_decap_8 FILLER_57_849 ();
 sg13g2_decap_4 FILLER_57_856 ();
 sg13g2_fill_2 FILLER_57_860 ();
 sg13g2_fill_1 FILLER_58_66 ();
 sg13g2_decap_4 FILLER_58_167 ();
 sg13g2_fill_1 FILLER_58_171 ();
 sg13g2_decap_4 FILLER_58_176 ();
 sg13g2_fill_1 FILLER_58_180 ();
 sg13g2_fill_2 FILLER_58_231 ();
 sg13g2_fill_1 FILLER_58_233 ();
 sg13g2_decap_4 FILLER_58_243 ();
 sg13g2_fill_1 FILLER_58_247 ();
 sg13g2_decap_8 FILLER_58_274 ();
 sg13g2_decap_4 FILLER_58_286 ();
 sg13g2_fill_2 FILLER_58_298 ();
 sg13g2_decap_4 FILLER_58_319 ();
 sg13g2_fill_1 FILLER_58_323 ();
 sg13g2_fill_2 FILLER_58_343 ();
 sg13g2_fill_1 FILLER_58_345 ();
 sg13g2_fill_2 FILLER_58_351 ();
 sg13g2_fill_1 FILLER_58_353 ();
 sg13g2_decap_4 FILLER_58_359 ();
 sg13g2_fill_1 FILLER_58_368 ();
 sg13g2_fill_1 FILLER_58_386 ();
 sg13g2_fill_2 FILLER_58_395 ();
 sg13g2_decap_4 FILLER_58_406 ();
 sg13g2_fill_2 FILLER_58_410 ();
 sg13g2_fill_2 FILLER_58_422 ();
 sg13g2_fill_2 FILLER_58_437 ();
 sg13g2_fill_1 FILLER_58_439 ();
 sg13g2_decap_4 FILLER_58_451 ();
 sg13g2_fill_1 FILLER_58_455 ();
 sg13g2_fill_2 FILLER_58_602 ();
 sg13g2_fill_2 FILLER_58_630 ();
 sg13g2_fill_1 FILLER_58_648 ();
 sg13g2_fill_2 FILLER_58_653 ();
 sg13g2_fill_1 FILLER_58_655 ();
 sg13g2_fill_2 FILLER_58_660 ();
 sg13g2_fill_1 FILLER_58_662 ();
 sg13g2_fill_1 FILLER_58_671 ();
 sg13g2_decap_8 FILLER_58_698 ();
 sg13g2_fill_1 FILLER_58_705 ();
 sg13g2_decap_8 FILLER_58_722 ();
 sg13g2_decap_8 FILLER_58_729 ();
 sg13g2_decap_8 FILLER_58_736 ();
 sg13g2_decap_8 FILLER_58_743 ();
 sg13g2_decap_8 FILLER_58_750 ();
 sg13g2_decap_8 FILLER_58_757 ();
 sg13g2_decap_8 FILLER_58_764 ();
 sg13g2_decap_8 FILLER_58_771 ();
 sg13g2_decap_8 FILLER_58_778 ();
 sg13g2_decap_8 FILLER_58_785 ();
 sg13g2_decap_8 FILLER_58_792 ();
 sg13g2_decap_8 FILLER_58_799 ();
 sg13g2_decap_8 FILLER_58_806 ();
 sg13g2_decap_8 FILLER_58_813 ();
 sg13g2_decap_8 FILLER_58_820 ();
 sg13g2_decap_8 FILLER_58_827 ();
 sg13g2_decap_8 FILLER_58_834 ();
 sg13g2_decap_8 FILLER_58_841 ();
 sg13g2_decap_8 FILLER_58_848 ();
 sg13g2_decap_8 FILLER_58_855 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_7 ();
 sg13g2_fill_2 FILLER_59_78 ();
 sg13g2_fill_1 FILLER_59_80 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_fill_1 FILLER_59_151 ();
 sg13g2_decap_4 FILLER_59_157 ();
 sg13g2_fill_1 FILLER_59_161 ();
 sg13g2_fill_2 FILLER_59_172 ();
 sg13g2_decap_8 FILLER_59_188 ();
 sg13g2_decap_8 FILLER_59_195 ();
 sg13g2_decap_4 FILLER_59_202 ();
 sg13g2_fill_2 FILLER_59_206 ();
 sg13g2_fill_2 FILLER_59_218 ();
 sg13g2_fill_1 FILLER_59_220 ();
 sg13g2_decap_4 FILLER_59_234 ();
 sg13g2_fill_1 FILLER_59_238 ();
 sg13g2_decap_8 FILLER_59_249 ();
 sg13g2_fill_2 FILLER_59_256 ();
 sg13g2_decap_8 FILLER_59_271 ();
 sg13g2_fill_2 FILLER_59_278 ();
 sg13g2_decap_4 FILLER_59_294 ();
 sg13g2_fill_1 FILLER_59_298 ();
 sg13g2_fill_2 FILLER_59_314 ();
 sg13g2_fill_2 FILLER_59_341 ();
 sg13g2_fill_1 FILLER_59_348 ();
 sg13g2_fill_2 FILLER_59_353 ();
 sg13g2_fill_1 FILLER_59_355 ();
 sg13g2_fill_1 FILLER_59_361 ();
 sg13g2_fill_1 FILLER_59_367 ();
 sg13g2_fill_2 FILLER_59_378 ();
 sg13g2_decap_4 FILLER_59_391 ();
 sg13g2_fill_2 FILLER_59_405 ();
 sg13g2_decap_8 FILLER_59_422 ();
 sg13g2_decap_8 FILLER_59_429 ();
 sg13g2_fill_2 FILLER_59_436 ();
 sg13g2_fill_1 FILLER_59_438 ();
 sg13g2_fill_2 FILLER_59_448 ();
 sg13g2_fill_2 FILLER_59_474 ();
 sg13g2_fill_1 FILLER_59_476 ();
 sg13g2_decap_8 FILLER_59_513 ();
 sg13g2_fill_1 FILLER_59_520 ();
 sg13g2_fill_2 FILLER_59_525 ();
 sg13g2_fill_2 FILLER_59_537 ();
 sg13g2_fill_1 FILLER_59_539 ();
 sg13g2_decap_4 FILLER_59_566 ();
 sg13g2_fill_2 FILLER_59_570 ();
 sg13g2_fill_2 FILLER_59_580 ();
 sg13g2_fill_1 FILLER_59_582 ();
 sg13g2_fill_1 FILLER_59_590 ();
 sg13g2_decap_8 FILLER_59_603 ();
 sg13g2_decap_8 FILLER_59_610 ();
 sg13g2_decap_8 FILLER_59_617 ();
 sg13g2_decap_8 FILLER_59_624 ();
 sg13g2_fill_2 FILLER_59_636 ();
 sg13g2_fill_2 FILLER_59_664 ();
 sg13g2_fill_1 FILLER_59_674 ();
 sg13g2_decap_4 FILLER_59_679 ();
 sg13g2_fill_1 FILLER_59_688 ();
 sg13g2_decap_4 FILLER_59_693 ();
 sg13g2_fill_2 FILLER_59_697 ();
 sg13g2_fill_1 FILLER_59_703 ();
 sg13g2_decap_8 FILLER_59_720 ();
 sg13g2_decap_8 FILLER_59_727 ();
 sg13g2_decap_8 FILLER_59_734 ();
 sg13g2_decap_8 FILLER_59_741 ();
 sg13g2_decap_8 FILLER_59_748 ();
 sg13g2_decap_8 FILLER_59_755 ();
 sg13g2_decap_8 FILLER_59_762 ();
 sg13g2_decap_8 FILLER_59_769 ();
 sg13g2_decap_8 FILLER_59_776 ();
 sg13g2_decap_8 FILLER_59_783 ();
 sg13g2_decap_8 FILLER_59_790 ();
 sg13g2_decap_8 FILLER_59_797 ();
 sg13g2_decap_8 FILLER_59_804 ();
 sg13g2_decap_8 FILLER_59_811 ();
 sg13g2_decap_8 FILLER_59_818 ();
 sg13g2_decap_8 FILLER_59_825 ();
 sg13g2_decap_8 FILLER_59_832 ();
 sg13g2_decap_8 FILLER_59_839 ();
 sg13g2_decap_8 FILLER_59_846 ();
 sg13g2_decap_8 FILLER_59_853 ();
 sg13g2_fill_2 FILLER_59_860 ();
 sg13g2_fill_2 FILLER_60_26 ();
 sg13g2_fill_1 FILLER_60_28 ();
 sg13g2_fill_2 FILLER_60_60 ();
 sg13g2_fill_1 FILLER_60_62 ();
 sg13g2_fill_2 FILLER_60_115 ();
 sg13g2_fill_1 FILLER_60_117 ();
 sg13g2_decap_8 FILLER_60_154 ();
 sg13g2_fill_1 FILLER_60_161 ();
 sg13g2_fill_2 FILLER_60_173 ();
 sg13g2_fill_1 FILLER_60_175 ();
 sg13g2_fill_2 FILLER_60_201 ();
 sg13g2_fill_1 FILLER_60_203 ();
 sg13g2_fill_2 FILLER_60_223 ();
 sg13g2_fill_1 FILLER_60_225 ();
 sg13g2_fill_1 FILLER_60_274 ();
 sg13g2_fill_1 FILLER_60_288 ();
 sg13g2_fill_1 FILLER_60_331 ();
 sg13g2_fill_2 FILLER_60_348 ();
 sg13g2_fill_1 FILLER_60_350 ();
 sg13g2_decap_8 FILLER_60_368 ();
 sg13g2_fill_1 FILLER_60_375 ();
 sg13g2_fill_2 FILLER_60_386 ();
 sg13g2_fill_1 FILLER_60_388 ();
 sg13g2_fill_2 FILLER_60_394 ();
 sg13g2_fill_1 FILLER_60_402 ();
 sg13g2_decap_8 FILLER_60_425 ();
 sg13g2_fill_2 FILLER_60_432 ();
 sg13g2_decap_8 FILLER_60_440 ();
 sg13g2_fill_2 FILLER_60_447 ();
 sg13g2_decap_8 FILLER_60_467 ();
 sg13g2_fill_1 FILLER_60_474 ();
 sg13g2_decap_8 FILLER_60_485 ();
 sg13g2_fill_1 FILLER_60_492 ();
 sg13g2_fill_2 FILLER_60_506 ();
 sg13g2_decap_4 FILLER_60_518 ();
 sg13g2_fill_1 FILLER_60_522 ();
 sg13g2_decap_8 FILLER_60_533 ();
 sg13g2_fill_2 FILLER_60_540 ();
 sg13g2_fill_1 FILLER_60_542 ();
 sg13g2_decap_4 FILLER_60_593 ();
 sg13g2_fill_1 FILLER_60_597 ();
 sg13g2_fill_1 FILLER_60_603 ();
 sg13g2_decap_8 FILLER_60_646 ();
 sg13g2_fill_2 FILLER_60_653 ();
 sg13g2_fill_1 FILLER_60_655 ();
 sg13g2_decap_4 FILLER_60_660 ();
 sg13g2_fill_1 FILLER_60_664 ();
 sg13g2_decap_8 FILLER_60_712 ();
 sg13g2_decap_8 FILLER_60_719 ();
 sg13g2_decap_4 FILLER_60_726 ();
 sg13g2_decap_8 FILLER_60_738 ();
 sg13g2_decap_8 FILLER_60_745 ();
 sg13g2_decap_8 FILLER_60_752 ();
 sg13g2_decap_8 FILLER_60_759 ();
 sg13g2_decap_8 FILLER_60_766 ();
 sg13g2_decap_8 FILLER_60_773 ();
 sg13g2_decap_8 FILLER_60_780 ();
 sg13g2_decap_8 FILLER_60_787 ();
 sg13g2_decap_8 FILLER_60_794 ();
 sg13g2_decap_8 FILLER_60_801 ();
 sg13g2_decap_8 FILLER_60_808 ();
 sg13g2_decap_8 FILLER_60_815 ();
 sg13g2_decap_8 FILLER_60_822 ();
 sg13g2_decap_8 FILLER_60_829 ();
 sg13g2_decap_8 FILLER_60_836 ();
 sg13g2_decap_8 FILLER_60_843 ();
 sg13g2_decap_8 FILLER_60_850 ();
 sg13g2_decap_4 FILLER_60_857 ();
 sg13g2_fill_1 FILLER_60_861 ();
 sg13g2_decap_4 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_4 ();
 sg13g2_fill_2 FILLER_61_85 ();
 sg13g2_fill_1 FILLER_61_87 ();
 sg13g2_fill_2 FILLER_61_97 ();
 sg13g2_fill_1 FILLER_61_99 ();
 sg13g2_decap_4 FILLER_61_104 ();
 sg13g2_fill_2 FILLER_61_108 ();
 sg13g2_decap_8 FILLER_61_124 ();
 sg13g2_fill_2 FILLER_61_131 ();
 sg13g2_fill_1 FILLER_61_133 ();
 sg13g2_decap_4 FILLER_61_147 ();
 sg13g2_fill_2 FILLER_61_151 ();
 sg13g2_fill_2 FILLER_61_170 ();
 sg13g2_fill_1 FILLER_61_172 ();
 sg13g2_decap_4 FILLER_61_202 ();
 sg13g2_fill_2 FILLER_61_224 ();
 sg13g2_fill_1 FILLER_61_226 ();
 sg13g2_decap_4 FILLER_61_232 ();
 sg13g2_fill_2 FILLER_61_236 ();
 sg13g2_decap_4 FILLER_61_248 ();
 sg13g2_fill_2 FILLER_61_252 ();
 sg13g2_fill_2 FILLER_61_267 ();
 sg13g2_decap_4 FILLER_61_279 ();
 sg13g2_fill_1 FILLER_61_283 ();
 sg13g2_fill_2 FILLER_61_297 ();
 sg13g2_fill_1 FILLER_61_299 ();
 sg13g2_decap_8 FILLER_61_304 ();
 sg13g2_decap_4 FILLER_61_311 ();
 sg13g2_fill_2 FILLER_61_321 ();
 sg13g2_fill_1 FILLER_61_338 ();
 sg13g2_decap_8 FILLER_61_345 ();
 sg13g2_fill_1 FILLER_61_352 ();
 sg13g2_fill_1 FILLER_61_366 ();
 sg13g2_fill_2 FILLER_61_393 ();
 sg13g2_decap_8 FILLER_61_476 ();
 sg13g2_fill_2 FILLER_61_493 ();
 sg13g2_fill_2 FILLER_61_557 ();
 sg13g2_fill_2 FILLER_61_572 ();
 sg13g2_fill_2 FILLER_61_600 ();
 sg13g2_decap_8 FILLER_61_623 ();
 sg13g2_decap_4 FILLER_61_630 ();
 sg13g2_decap_4 FILLER_61_696 ();
 sg13g2_fill_1 FILLER_61_700 ();
 sg13g2_fill_1 FILLER_61_706 ();
 sg13g2_decap_8 FILLER_61_741 ();
 sg13g2_decap_8 FILLER_61_748 ();
 sg13g2_decap_8 FILLER_61_755 ();
 sg13g2_decap_8 FILLER_61_762 ();
 sg13g2_decap_8 FILLER_61_769 ();
 sg13g2_decap_8 FILLER_61_776 ();
 sg13g2_decap_8 FILLER_61_783 ();
 sg13g2_decap_8 FILLER_61_790 ();
 sg13g2_decap_8 FILLER_61_797 ();
 sg13g2_decap_8 FILLER_61_804 ();
 sg13g2_decap_8 FILLER_61_811 ();
 sg13g2_decap_8 FILLER_61_818 ();
 sg13g2_decap_8 FILLER_61_825 ();
 sg13g2_decap_8 FILLER_61_832 ();
 sg13g2_decap_8 FILLER_61_839 ();
 sg13g2_decap_8 FILLER_61_846 ();
 sg13g2_decap_8 FILLER_61_853 ();
 sg13g2_fill_2 FILLER_61_860 ();
 sg13g2_fill_1 FILLER_62_26 ();
 sg13g2_decap_8 FILLER_62_106 ();
 sg13g2_fill_1 FILLER_62_113 ();
 sg13g2_fill_1 FILLER_62_150 ();
 sg13g2_decap_4 FILLER_62_169 ();
 sg13g2_fill_2 FILLER_62_209 ();
 sg13g2_fill_1 FILLER_62_211 ();
 sg13g2_decap_4 FILLER_62_238 ();
 sg13g2_decap_4 FILLER_62_272 ();
 sg13g2_fill_2 FILLER_62_276 ();
 sg13g2_fill_2 FILLER_62_304 ();
 sg13g2_decap_4 FILLER_62_310 ();
 sg13g2_fill_2 FILLER_62_314 ();
 sg13g2_decap_8 FILLER_62_369 ();
 sg13g2_fill_2 FILLER_62_376 ();
 sg13g2_decap_4 FILLER_62_403 ();
 sg13g2_fill_2 FILLER_62_407 ();
 sg13g2_fill_2 FILLER_62_414 ();
 sg13g2_decap_8 FILLER_62_424 ();
 sg13g2_decap_4 FILLER_62_431 ();
 sg13g2_fill_2 FILLER_62_440 ();
 sg13g2_fill_1 FILLER_62_442 ();
 sg13g2_decap_4 FILLER_62_465 ();
 sg13g2_fill_2 FILLER_62_469 ();
 sg13g2_decap_8 FILLER_62_497 ();
 sg13g2_decap_8 FILLER_62_517 ();
 sg13g2_decap_8 FILLER_62_524 ();
 sg13g2_fill_2 FILLER_62_531 ();
 sg13g2_fill_1 FILLER_62_533 ();
 sg13g2_fill_2 FILLER_62_560 ();
 sg13g2_fill_1 FILLER_62_562 ();
 sg13g2_decap_8 FILLER_62_567 ();
 sg13g2_decap_4 FILLER_62_574 ();
 sg13g2_fill_2 FILLER_62_578 ();
 sg13g2_fill_1 FILLER_62_601 ();
 sg13g2_fill_1 FILLER_62_623 ();
 sg13g2_fill_2 FILLER_62_635 ();
 sg13g2_fill_2 FILLER_62_660 ();
 sg13g2_fill_1 FILLER_62_662 ();
 sg13g2_fill_1 FILLER_62_678 ();
 sg13g2_decap_4 FILLER_62_713 ();
 sg13g2_fill_1 FILLER_62_717 ();
 sg13g2_decap_4 FILLER_62_722 ();
 sg13g2_fill_2 FILLER_62_726 ();
 sg13g2_decap_8 FILLER_62_739 ();
 sg13g2_decap_8 FILLER_62_746 ();
 sg13g2_decap_8 FILLER_62_753 ();
 sg13g2_decap_8 FILLER_62_760 ();
 sg13g2_decap_8 FILLER_62_767 ();
 sg13g2_decap_8 FILLER_62_774 ();
 sg13g2_decap_8 FILLER_62_781 ();
 sg13g2_decap_8 FILLER_62_788 ();
 sg13g2_decap_8 FILLER_62_795 ();
 sg13g2_decap_8 FILLER_62_802 ();
 sg13g2_decap_8 FILLER_62_809 ();
 sg13g2_decap_8 FILLER_62_816 ();
 sg13g2_decap_8 FILLER_62_823 ();
 sg13g2_decap_8 FILLER_62_830 ();
 sg13g2_decap_8 FILLER_62_837 ();
 sg13g2_decap_8 FILLER_62_844 ();
 sg13g2_decap_8 FILLER_62_851 ();
 sg13g2_decap_4 FILLER_62_858 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_fill_2 FILLER_63_37 ();
 sg13g2_fill_1 FILLER_63_39 ();
 sg13g2_fill_2 FILLER_63_82 ();
 sg13g2_fill_1 FILLER_63_84 ();
 sg13g2_fill_2 FILLER_63_111 ();
 sg13g2_fill_2 FILLER_63_119 ();
 sg13g2_decap_4 FILLER_63_130 ();
 sg13g2_fill_1 FILLER_63_134 ();
 sg13g2_decap_4 FILLER_63_143 ();
 sg13g2_decap_8 FILLER_63_150 ();
 sg13g2_fill_1 FILLER_63_157 ();
 sg13g2_decap_4 FILLER_63_173 ();
 sg13g2_fill_2 FILLER_63_187 ();
 sg13g2_fill_1 FILLER_63_189 ();
 sg13g2_decap_8 FILLER_63_199 ();
 sg13g2_decap_4 FILLER_63_206 ();
 sg13g2_fill_2 FILLER_63_210 ();
 sg13g2_decap_4 FILLER_63_230 ();
 sg13g2_fill_2 FILLER_63_234 ();
 sg13g2_fill_2 FILLER_63_246 ();
 sg13g2_fill_1 FILLER_63_266 ();
 sg13g2_decap_8 FILLER_63_283 ();
 sg13g2_fill_2 FILLER_63_326 ();
 sg13g2_fill_1 FILLER_63_333 ();
 sg13g2_decap_8 FILLER_63_353 ();
 sg13g2_decap_4 FILLER_63_370 ();
 sg13g2_decap_8 FILLER_63_378 ();
 sg13g2_fill_2 FILLER_63_385 ();
 sg13g2_decap_4 FILLER_63_392 ();
 sg13g2_fill_2 FILLER_63_396 ();
 sg13g2_decap_8 FILLER_63_434 ();
 sg13g2_decap_4 FILLER_63_441 ();
 sg13g2_decap_8 FILLER_63_449 ();
 sg13g2_decap_4 FILLER_63_456 ();
 sg13g2_fill_2 FILLER_63_460 ();
 sg13g2_fill_1 FILLER_63_481 ();
 sg13g2_fill_2 FILLER_63_486 ();
 sg13g2_fill_1 FILLER_63_494 ();
 sg13g2_fill_2 FILLER_63_513 ();
 sg13g2_fill_2 FILLER_63_524 ();
 sg13g2_fill_2 FILLER_63_539 ();
 sg13g2_fill_1 FILLER_63_558 ();
 sg13g2_decap_4 FILLER_63_585 ();
 sg13g2_fill_1 FILLER_63_589 ();
 sg13g2_decap_4 FILLER_63_598 ();
 sg13g2_decap_8 FILLER_63_682 ();
 sg13g2_decap_8 FILLER_63_689 ();
 sg13g2_decap_4 FILLER_63_703 ();
 sg13g2_fill_2 FILLER_63_707 ();
 sg13g2_decap_8 FILLER_63_740 ();
 sg13g2_decap_8 FILLER_63_747 ();
 sg13g2_decap_8 FILLER_63_754 ();
 sg13g2_decap_8 FILLER_63_761 ();
 sg13g2_decap_8 FILLER_63_768 ();
 sg13g2_decap_8 FILLER_63_775 ();
 sg13g2_decap_8 FILLER_63_782 ();
 sg13g2_decap_8 FILLER_63_789 ();
 sg13g2_decap_8 FILLER_63_796 ();
 sg13g2_decap_8 FILLER_63_803 ();
 sg13g2_decap_8 FILLER_63_810 ();
 sg13g2_decap_8 FILLER_63_817 ();
 sg13g2_decap_8 FILLER_63_824 ();
 sg13g2_decap_8 FILLER_63_831 ();
 sg13g2_decap_8 FILLER_63_838 ();
 sg13g2_decap_8 FILLER_63_845 ();
 sg13g2_decap_8 FILLER_63_852 ();
 sg13g2_fill_2 FILLER_63_859 ();
 sg13g2_fill_1 FILLER_63_861 ();
 sg13g2_decap_4 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_27 ();
 sg13g2_decap_4 FILLER_64_64 ();
 sg13g2_fill_2 FILLER_64_91 ();
 sg13g2_decap_4 FILLER_64_103 ();
 sg13g2_fill_1 FILLER_64_107 ();
 sg13g2_fill_2 FILLER_64_112 ();
 sg13g2_fill_2 FILLER_64_120 ();
 sg13g2_fill_1 FILLER_64_122 ();
 sg13g2_decap_4 FILLER_64_175 ();
 sg13g2_fill_1 FILLER_64_179 ();
 sg13g2_decap_8 FILLER_64_185 ();
 sg13g2_fill_1 FILLER_64_192 ();
 sg13g2_fill_2 FILLER_64_210 ();
 sg13g2_fill_1 FILLER_64_223 ();
 sg13g2_decap_8 FILLER_64_229 ();
 sg13g2_decap_4 FILLER_64_236 ();
 sg13g2_fill_2 FILLER_64_240 ();
 sg13g2_decap_4 FILLER_64_313 ();
 sg13g2_fill_1 FILLER_64_332 ();
 sg13g2_decap_4 FILLER_64_359 ();
 sg13g2_decap_4 FILLER_64_389 ();
 sg13g2_fill_2 FILLER_64_393 ();
 sg13g2_fill_1 FILLER_64_405 ();
 sg13g2_fill_2 FILLER_64_432 ();
 sg13g2_fill_1 FILLER_64_536 ();
 sg13g2_fill_1 FILLER_64_551 ();
 sg13g2_fill_2 FILLER_64_565 ();
 sg13g2_fill_2 FILLER_64_611 ();
 sg13g2_decap_8 FILLER_64_617 ();
 sg13g2_fill_2 FILLER_64_624 ();
 sg13g2_decap_8 FILLER_64_630 ();
 sg13g2_decap_4 FILLER_64_637 ();
 sg13g2_fill_2 FILLER_64_641 ();
 sg13g2_fill_2 FILLER_64_655 ();
 sg13g2_fill_1 FILLER_64_677 ();
 sg13g2_fill_2 FILLER_64_686 ();
 sg13g2_decap_8 FILLER_64_710 ();
 sg13g2_fill_2 FILLER_64_717 ();
 sg13g2_decap_8 FILLER_64_727 ();
 sg13g2_decap_8 FILLER_64_734 ();
 sg13g2_decap_8 FILLER_64_741 ();
 sg13g2_decap_8 FILLER_64_748 ();
 sg13g2_decap_8 FILLER_64_755 ();
 sg13g2_decap_8 FILLER_64_762 ();
 sg13g2_decap_8 FILLER_64_769 ();
 sg13g2_decap_8 FILLER_64_776 ();
 sg13g2_decap_8 FILLER_64_783 ();
 sg13g2_decap_8 FILLER_64_790 ();
 sg13g2_decap_8 FILLER_64_797 ();
 sg13g2_decap_8 FILLER_64_804 ();
 sg13g2_decap_8 FILLER_64_811 ();
 sg13g2_decap_8 FILLER_64_818 ();
 sg13g2_decap_8 FILLER_64_825 ();
 sg13g2_decap_8 FILLER_64_832 ();
 sg13g2_decap_8 FILLER_64_839 ();
 sg13g2_decap_8 FILLER_64_846 ();
 sg13g2_decap_8 FILLER_64_853 ();
 sg13g2_fill_2 FILLER_64_860 ();
 sg13g2_decap_4 FILLER_65_26 ();
 sg13g2_fill_2 FILLER_65_30 ();
 sg13g2_fill_1 FILLER_65_64 ();
 sg13g2_fill_2 FILLER_65_91 ();
 sg13g2_fill_1 FILLER_65_123 ();
 sg13g2_fill_1 FILLER_65_132 ();
 sg13g2_fill_1 FILLER_65_138 ();
 sg13g2_fill_2 FILLER_65_164 ();
 sg13g2_fill_1 FILLER_65_166 ();
 sg13g2_decap_8 FILLER_65_215 ();
 sg13g2_decap_4 FILLER_65_222 ();
 sg13g2_fill_2 FILLER_65_231 ();
 sg13g2_decap_8 FILLER_65_246 ();
 sg13g2_fill_1 FILLER_65_253 ();
 sg13g2_fill_2 FILLER_65_271 ();
 sg13g2_decap_4 FILLER_65_318 ();
 sg13g2_decap_4 FILLER_65_340 ();
 sg13g2_fill_2 FILLER_65_348 ();
 sg13g2_fill_1 FILLER_65_350 ();
 sg13g2_decap_8 FILLER_65_387 ();
 sg13g2_fill_2 FILLER_65_394 ();
 sg13g2_fill_1 FILLER_65_396 ();
 sg13g2_decap_4 FILLER_65_428 ();
 sg13g2_fill_2 FILLER_65_455 ();
 sg13g2_fill_2 FILLER_65_476 ();
 sg13g2_fill_2 FILLER_65_495 ();
 sg13g2_fill_1 FILLER_65_506 ();
 sg13g2_fill_2 FILLER_65_515 ();
 sg13g2_fill_1 FILLER_65_517 ();
 sg13g2_fill_2 FILLER_65_526 ();
 sg13g2_fill_2 FILLER_65_541 ();
 sg13g2_fill_1 FILLER_65_543 ();
 sg13g2_fill_2 FILLER_65_550 ();
 sg13g2_decap_4 FILLER_65_578 ();
 sg13g2_fill_1 FILLER_65_582 ();
 sg13g2_decap_8 FILLER_65_601 ();
 sg13g2_fill_1 FILLER_65_608 ();
 sg13g2_fill_2 FILLER_65_613 ();
 sg13g2_decap_4 FILLER_65_641 ();
 sg13g2_fill_2 FILLER_65_645 ();
 sg13g2_fill_1 FILLER_65_651 ();
 sg13g2_decap_4 FILLER_65_668 ();
 sg13g2_fill_1 FILLER_65_672 ();
 sg13g2_fill_1 FILLER_65_686 ();
 sg13g2_fill_1 FILLER_65_696 ();
 sg13g2_decap_8 FILLER_65_704 ();
 sg13g2_fill_1 FILLER_65_711 ();
 sg13g2_decap_8 FILLER_65_738 ();
 sg13g2_decap_8 FILLER_65_745 ();
 sg13g2_decap_8 FILLER_65_752 ();
 sg13g2_decap_8 FILLER_65_759 ();
 sg13g2_decap_8 FILLER_65_766 ();
 sg13g2_decap_8 FILLER_65_773 ();
 sg13g2_decap_8 FILLER_65_780 ();
 sg13g2_decap_8 FILLER_65_787 ();
 sg13g2_decap_8 FILLER_65_794 ();
 sg13g2_decap_8 FILLER_65_801 ();
 sg13g2_decap_8 FILLER_65_808 ();
 sg13g2_decap_8 FILLER_65_815 ();
 sg13g2_decap_8 FILLER_65_822 ();
 sg13g2_decap_8 FILLER_65_829 ();
 sg13g2_decap_8 FILLER_65_836 ();
 sg13g2_decap_8 FILLER_65_843 ();
 sg13g2_decap_8 FILLER_65_850 ();
 sg13g2_decap_4 FILLER_65_857 ();
 sg13g2_fill_1 FILLER_65_861 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_4 FILLER_66_7 ();
 sg13g2_fill_2 FILLER_66_15 ();
 sg13g2_decap_8 FILLER_66_27 ();
 sg13g2_fill_2 FILLER_66_34 ();
 sg13g2_fill_2 FILLER_66_55 ();
 sg13g2_fill_1 FILLER_66_57 ();
 sg13g2_decap_8 FILLER_66_68 ();
 sg13g2_fill_1 FILLER_66_75 ();
 sg13g2_fill_2 FILLER_66_85 ();
 sg13g2_fill_2 FILLER_66_95 ();
 sg13g2_fill_1 FILLER_66_97 ();
 sg13g2_fill_2 FILLER_66_112 ();
 sg13g2_fill_1 FILLER_66_114 ();
 sg13g2_fill_2 FILLER_66_134 ();
 sg13g2_decap_4 FILLER_66_146 ();
 sg13g2_fill_2 FILLER_66_173 ();
 sg13g2_fill_1 FILLER_66_175 ();
 sg13g2_decap_8 FILLER_66_193 ();
 sg13g2_fill_2 FILLER_66_214 ();
 sg13g2_fill_1 FILLER_66_216 ();
 sg13g2_decap_4 FILLER_66_222 ();
 sg13g2_decap_8 FILLER_66_248 ();
 sg13g2_decap_4 FILLER_66_255 ();
 sg13g2_fill_1 FILLER_66_302 ();
 sg13g2_decap_4 FILLER_66_327 ();
 sg13g2_decap_8 FILLER_66_357 ();
 sg13g2_fill_2 FILLER_66_364 ();
 sg13g2_fill_1 FILLER_66_366 ();
 sg13g2_decap_4 FILLER_66_385 ();
 sg13g2_fill_2 FILLER_66_389 ();
 sg13g2_decap_4 FILLER_66_396 ();
 sg13g2_fill_2 FILLER_66_405 ();
 sg13g2_fill_1 FILLER_66_420 ();
 sg13g2_fill_2 FILLER_66_476 ();
 sg13g2_fill_1 FILLER_66_478 ();
 sg13g2_fill_2 FILLER_66_561 ();
 sg13g2_fill_2 FILLER_66_567 ();
 sg13g2_fill_1 FILLER_66_577 ();
 sg13g2_decap_4 FILLER_66_585 ();
 sg13g2_fill_1 FILLER_66_589 ();
 sg13g2_fill_2 FILLER_66_624 ();
 sg13g2_fill_2 FILLER_66_650 ();
 sg13g2_decap_4 FILLER_66_670 ();
 sg13g2_fill_1 FILLER_66_674 ();
 sg13g2_decap_4 FILLER_66_679 ();
 sg13g2_decap_8 FILLER_66_691 ();
 sg13g2_decap_8 FILLER_66_698 ();
 sg13g2_decap_8 FILLER_66_731 ();
 sg13g2_decap_8 FILLER_66_738 ();
 sg13g2_decap_8 FILLER_66_745 ();
 sg13g2_decap_8 FILLER_66_752 ();
 sg13g2_decap_8 FILLER_66_759 ();
 sg13g2_decap_8 FILLER_66_766 ();
 sg13g2_decap_8 FILLER_66_773 ();
 sg13g2_decap_8 FILLER_66_780 ();
 sg13g2_decap_8 FILLER_66_787 ();
 sg13g2_decap_8 FILLER_66_794 ();
 sg13g2_decap_8 FILLER_66_801 ();
 sg13g2_decap_8 FILLER_66_808 ();
 sg13g2_decap_8 FILLER_66_815 ();
 sg13g2_decap_8 FILLER_66_822 ();
 sg13g2_decap_8 FILLER_66_829 ();
 sg13g2_decap_8 FILLER_66_836 ();
 sg13g2_decap_8 FILLER_66_843 ();
 sg13g2_decap_8 FILLER_66_850 ();
 sg13g2_decap_4 FILLER_66_857 ();
 sg13g2_fill_1 FILLER_66_861 ();
 sg13g2_fill_1 FILLER_67_26 ();
 sg13g2_fill_2 FILLER_67_53 ();
 sg13g2_fill_1 FILLER_67_104 ();
 sg13g2_fill_2 FILLER_67_150 ();
 sg13g2_fill_1 FILLER_67_152 ();
 sg13g2_fill_2 FILLER_67_158 ();
 sg13g2_fill_1 FILLER_67_160 ();
 sg13g2_decap_8 FILLER_67_170 ();
 sg13g2_fill_2 FILLER_67_203 ();
 sg13g2_fill_1 FILLER_67_205 ();
 sg13g2_fill_2 FILLER_67_211 ();
 sg13g2_fill_1 FILLER_67_218 ();
 sg13g2_fill_2 FILLER_67_228 ();
 sg13g2_fill_1 FILLER_67_230 ();
 sg13g2_fill_2 FILLER_67_236 ();
 sg13g2_fill_1 FILLER_67_255 ();
 sg13g2_fill_1 FILLER_67_321 ();
 sg13g2_fill_2 FILLER_67_343 ();
 sg13g2_fill_1 FILLER_67_345 ();
 sg13g2_fill_2 FILLER_67_359 ();
 sg13g2_fill_1 FILLER_67_361 ();
 sg13g2_decap_4 FILLER_67_383 ();
 sg13g2_fill_1 FILLER_67_387 ();
 sg13g2_fill_2 FILLER_67_398 ();
 sg13g2_fill_1 FILLER_67_400 ();
 sg13g2_decap_8 FILLER_67_437 ();
 sg13g2_fill_1 FILLER_67_444 ();
 sg13g2_fill_2 FILLER_67_454 ();
 sg13g2_fill_1 FILLER_67_460 ();
 sg13g2_decap_4 FILLER_67_465 ();
 sg13g2_fill_2 FILLER_67_469 ();
 sg13g2_fill_2 FILLER_67_475 ();
 sg13g2_fill_1 FILLER_67_477 ();
 sg13g2_fill_2 FILLER_67_486 ();
 sg13g2_fill_1 FILLER_67_488 ();
 sg13g2_fill_2 FILLER_67_518 ();
 sg13g2_fill_1 FILLER_67_541 ();
 sg13g2_fill_2 FILLER_67_553 ();
 sg13g2_decap_4 FILLER_67_588 ();
 sg13g2_decap_8 FILLER_67_596 ();
 sg13g2_decap_8 FILLER_67_603 ();
 sg13g2_fill_1 FILLER_67_610 ();
 sg13g2_decap_4 FILLER_67_644 ();
 sg13g2_fill_2 FILLER_67_648 ();
 sg13g2_fill_1 FILLER_67_654 ();
 sg13g2_fill_2 FILLER_67_672 ();
 sg13g2_fill_1 FILLER_67_674 ();
 sg13g2_decap_8 FILLER_67_701 ();
 sg13g2_decap_4 FILLER_67_708 ();
 sg13g2_decap_4 FILLER_67_720 ();
 sg13g2_fill_2 FILLER_67_724 ();
 sg13g2_decap_8 FILLER_67_734 ();
 sg13g2_decap_8 FILLER_67_741 ();
 sg13g2_decap_8 FILLER_67_748 ();
 sg13g2_decap_8 FILLER_67_755 ();
 sg13g2_decap_8 FILLER_67_762 ();
 sg13g2_decap_8 FILLER_67_769 ();
 sg13g2_decap_8 FILLER_67_776 ();
 sg13g2_decap_8 FILLER_67_783 ();
 sg13g2_decap_8 FILLER_67_790 ();
 sg13g2_decap_8 FILLER_67_797 ();
 sg13g2_decap_8 FILLER_67_804 ();
 sg13g2_decap_8 FILLER_67_811 ();
 sg13g2_decap_8 FILLER_67_818 ();
 sg13g2_decap_8 FILLER_67_825 ();
 sg13g2_decap_8 FILLER_67_832 ();
 sg13g2_decap_8 FILLER_67_839 ();
 sg13g2_decap_8 FILLER_67_846 ();
 sg13g2_decap_8 FILLER_67_853 ();
 sg13g2_fill_2 FILLER_67_860 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_4 FILLER_68_7 ();
 sg13g2_decap_4 FILLER_68_15 ();
 sg13g2_fill_2 FILLER_68_42 ();
 sg13g2_fill_1 FILLER_68_44 ();
 sg13g2_fill_1 FILLER_68_60 ();
 sg13g2_decap_4 FILLER_68_66 ();
 sg13g2_fill_1 FILLER_68_70 ();
 sg13g2_fill_2 FILLER_68_75 ();
 sg13g2_fill_1 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_114 ();
 sg13g2_decap_4 FILLER_68_121 ();
 sg13g2_fill_2 FILLER_68_147 ();
 sg13g2_fill_1 FILLER_68_149 ();
 sg13g2_fill_2 FILLER_68_163 ();
 sg13g2_fill_1 FILLER_68_165 ();
 sg13g2_fill_1 FILLER_68_210 ();
 sg13g2_decap_8 FILLER_68_254 ();
 sg13g2_fill_2 FILLER_68_285 ();
 sg13g2_fill_2 FILLER_68_296 ();
 sg13g2_fill_1 FILLER_68_298 ();
 sg13g2_decap_8 FILLER_68_318 ();
 sg13g2_decap_8 FILLER_68_325 ();
 sg13g2_fill_2 FILLER_68_332 ();
 sg13g2_decap_8 FILLER_68_402 ();
 sg13g2_fill_2 FILLER_68_409 ();
 sg13g2_fill_1 FILLER_68_434 ();
 sg13g2_decap_4 FILLER_68_471 ();
 sg13g2_fill_1 FILLER_68_475 ();
 sg13g2_fill_2 FILLER_68_497 ();
 sg13g2_fill_1 FILLER_68_499 ();
 sg13g2_fill_2 FILLER_68_512 ();
 sg13g2_fill_1 FILLER_68_514 ();
 sg13g2_fill_2 FILLER_68_614 ();
 sg13g2_decap_8 FILLER_68_642 ();
 sg13g2_decap_8 FILLER_68_649 ();
 sg13g2_decap_8 FILLER_68_660 ();
 sg13g2_decap_8 FILLER_68_667 ();
 sg13g2_decap_8 FILLER_68_674 ();
 sg13g2_decap_4 FILLER_68_681 ();
 sg13g2_fill_1 FILLER_68_685 ();
 sg13g2_fill_1 FILLER_68_690 ();
 sg13g2_fill_2 FILLER_68_699 ();
 sg13g2_decap_8 FILLER_68_743 ();
 sg13g2_decap_8 FILLER_68_750 ();
 sg13g2_decap_8 FILLER_68_757 ();
 sg13g2_decap_8 FILLER_68_764 ();
 sg13g2_decap_8 FILLER_68_771 ();
 sg13g2_decap_8 FILLER_68_778 ();
 sg13g2_decap_8 FILLER_68_785 ();
 sg13g2_decap_8 FILLER_68_792 ();
 sg13g2_decap_8 FILLER_68_799 ();
 sg13g2_decap_8 FILLER_68_806 ();
 sg13g2_decap_8 FILLER_68_813 ();
 sg13g2_decap_8 FILLER_68_820 ();
 sg13g2_decap_8 FILLER_68_827 ();
 sg13g2_decap_8 FILLER_68_834 ();
 sg13g2_decap_8 FILLER_68_841 ();
 sg13g2_decap_8 FILLER_68_848 ();
 sg13g2_decap_8 FILLER_68_855 ();
 sg13g2_decap_4 FILLER_69_41 ();
 sg13g2_fill_1 FILLER_69_55 ();
 sg13g2_decap_8 FILLER_69_65 ();
 sg13g2_fill_2 FILLER_69_72 ();
 sg13g2_fill_1 FILLER_69_78 ();
 sg13g2_fill_2 FILLER_69_93 ();
 sg13g2_decap_8 FILLER_69_127 ();
 sg13g2_fill_2 FILLER_69_147 ();
 sg13g2_fill_1 FILLER_69_149 ();
 sg13g2_fill_2 FILLER_69_158 ();
 sg13g2_fill_1 FILLER_69_160 ();
 sg13g2_decap_8 FILLER_69_191 ();
 sg13g2_decap_4 FILLER_69_198 ();
 sg13g2_fill_2 FILLER_69_202 ();
 sg13g2_fill_1 FILLER_69_219 ();
 sg13g2_fill_2 FILLER_69_233 ();
 sg13g2_decap_4 FILLER_69_261 ();
 sg13g2_fill_2 FILLER_69_265 ();
 sg13g2_decap_8 FILLER_69_313 ();
 sg13g2_decap_8 FILLER_69_355 ();
 sg13g2_decap_4 FILLER_69_362 ();
 sg13g2_fill_1 FILLER_69_366 ();
 sg13g2_fill_2 FILLER_69_377 ();
 sg13g2_fill_1 FILLER_69_379 ();
 sg13g2_fill_2 FILLER_69_403 ();
 sg13g2_fill_1 FILLER_69_405 ();
 sg13g2_decap_4 FILLER_69_420 ();
 sg13g2_decap_8 FILLER_69_529 ();
 sg13g2_fill_1 FILLER_69_536 ();
 sg13g2_fill_1 FILLER_69_542 ();
 sg13g2_decap_8 FILLER_69_547 ();
 sg13g2_fill_1 FILLER_69_554 ();
 sg13g2_fill_2 FILLER_69_563 ();
 sg13g2_fill_2 FILLER_69_569 ();
 sg13g2_decap_8 FILLER_69_583 ();
 sg13g2_decap_8 FILLER_69_590 ();
 sg13g2_decap_8 FILLER_69_602 ();
 sg13g2_decap_8 FILLER_69_627 ();
 sg13g2_decap_8 FILLER_69_634 ();
 sg13g2_decap_4 FILLER_69_641 ();
 sg13g2_fill_1 FILLER_69_671 ();
 sg13g2_decap_4 FILLER_69_712 ();
 sg13g2_fill_1 FILLER_69_716 ();
 sg13g2_decap_4 FILLER_69_721 ();
 sg13g2_fill_1 FILLER_69_725 ();
 sg13g2_decap_8 FILLER_69_734 ();
 sg13g2_decap_8 FILLER_69_741 ();
 sg13g2_decap_8 FILLER_69_748 ();
 sg13g2_decap_8 FILLER_69_755 ();
 sg13g2_decap_8 FILLER_69_762 ();
 sg13g2_decap_8 FILLER_69_769 ();
 sg13g2_decap_8 FILLER_69_776 ();
 sg13g2_decap_8 FILLER_69_783 ();
 sg13g2_decap_8 FILLER_69_790 ();
 sg13g2_decap_8 FILLER_69_797 ();
 sg13g2_decap_8 FILLER_69_804 ();
 sg13g2_decap_8 FILLER_69_811 ();
 sg13g2_decap_8 FILLER_69_818 ();
 sg13g2_decap_8 FILLER_69_825 ();
 sg13g2_decap_8 FILLER_69_832 ();
 sg13g2_decap_8 FILLER_69_839 ();
 sg13g2_decap_8 FILLER_69_846 ();
 sg13g2_decap_8 FILLER_69_853 ();
 sg13g2_fill_2 FILLER_69_860 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_4 FILLER_70_7 ();
 sg13g2_fill_1 FILLER_70_15 ();
 sg13g2_fill_2 FILLER_70_25 ();
 sg13g2_decap_8 FILLER_70_134 ();
 sg13g2_fill_2 FILLER_70_149 ();
 sg13g2_decap_8 FILLER_70_197 ();
 sg13g2_fill_1 FILLER_70_204 ();
 sg13g2_fill_1 FILLER_70_235 ();
 sg13g2_fill_1 FILLER_70_272 ();
 sg13g2_fill_1 FILLER_70_323 ();
 sg13g2_fill_2 FILLER_70_343 ();
 sg13g2_fill_2 FILLER_70_371 ();
 sg13g2_fill_1 FILLER_70_373 ();
 sg13g2_decap_4 FILLER_70_431 ();
 sg13g2_fill_2 FILLER_70_435 ();
 sg13g2_fill_2 FILLER_70_442 ();
 sg13g2_decap_4 FILLER_70_457 ();
 sg13g2_fill_2 FILLER_70_471 ();
 sg13g2_fill_1 FILLER_70_499 ();
 sg13g2_fill_2 FILLER_70_504 ();
 sg13g2_fill_1 FILLER_70_506 ();
 sg13g2_decap_8 FILLER_70_512 ();
 sg13g2_fill_2 FILLER_70_519 ();
 sg13g2_fill_2 FILLER_70_542 ();
 sg13g2_fill_1 FILLER_70_544 ();
 sg13g2_fill_2 FILLER_70_557 ();
 sg13g2_fill_2 FILLER_70_588 ();
 sg13g2_decap_4 FILLER_70_598 ();
 sg13g2_fill_2 FILLER_70_614 ();
 sg13g2_fill_2 FILLER_70_634 ();
 sg13g2_decap_4 FILLER_70_666 ();
 sg13g2_fill_2 FILLER_70_670 ();
 sg13g2_decap_4 FILLER_70_702 ();
 sg13g2_decap_8 FILLER_70_732 ();
 sg13g2_decap_8 FILLER_70_739 ();
 sg13g2_decap_8 FILLER_70_746 ();
 sg13g2_decap_8 FILLER_70_753 ();
 sg13g2_decap_8 FILLER_70_760 ();
 sg13g2_decap_8 FILLER_70_767 ();
 sg13g2_decap_8 FILLER_70_774 ();
 sg13g2_decap_8 FILLER_70_781 ();
 sg13g2_decap_8 FILLER_70_788 ();
 sg13g2_decap_8 FILLER_70_795 ();
 sg13g2_decap_8 FILLER_70_802 ();
 sg13g2_decap_8 FILLER_70_809 ();
 sg13g2_decap_8 FILLER_70_816 ();
 sg13g2_decap_8 FILLER_70_823 ();
 sg13g2_decap_8 FILLER_70_830 ();
 sg13g2_decap_8 FILLER_70_837 ();
 sg13g2_decap_8 FILLER_70_844 ();
 sg13g2_decap_8 FILLER_70_851 ();
 sg13g2_decap_4 FILLER_70_858 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_7 ();
 sg13g2_fill_1 FILLER_71_9 ();
 sg13g2_fill_2 FILLER_71_46 ();
 sg13g2_fill_1 FILLER_71_60 ();
 sg13g2_decap_8 FILLER_71_125 ();
 sg13g2_fill_1 FILLER_71_132 ();
 sg13g2_decap_4 FILLER_71_174 ();
 sg13g2_decap_4 FILLER_71_190 ();
 sg13g2_fill_2 FILLER_71_203 ();
 sg13g2_fill_1 FILLER_71_205 ();
 sg13g2_fill_2 FILLER_71_222 ();
 sg13g2_fill_1 FILLER_71_224 ();
 sg13g2_decap_8 FILLER_71_264 ();
 sg13g2_decap_4 FILLER_71_271 ();
 sg13g2_decap_8 FILLER_71_280 ();
 sg13g2_decap_8 FILLER_71_299 ();
 sg13g2_fill_2 FILLER_71_306 ();
 sg13g2_decap_8 FILLER_71_311 ();
 sg13g2_fill_1 FILLER_71_318 ();
 sg13g2_decap_8 FILLER_71_331 ();
 sg13g2_decap_4 FILLER_71_338 ();
 sg13g2_fill_1 FILLER_71_342 ();
 sg13g2_fill_1 FILLER_71_353 ();
 sg13g2_fill_2 FILLER_71_377 ();
 sg13g2_fill_1 FILLER_71_379 ();
 sg13g2_decap_8 FILLER_71_394 ();
 sg13g2_fill_1 FILLER_71_410 ();
 sg13g2_decap_4 FILLER_71_425 ();
 sg13g2_fill_2 FILLER_71_429 ();
 sg13g2_fill_1 FILLER_71_441 ();
 sg13g2_decap_8 FILLER_71_468 ();
 sg13g2_fill_1 FILLER_71_475 ();
 sg13g2_fill_1 FILLER_71_502 ();
 sg13g2_fill_2 FILLER_71_515 ();
 sg13g2_decap_8 FILLER_71_530 ();
 sg13g2_decap_8 FILLER_71_537 ();
 sg13g2_fill_1 FILLER_71_544 ();
 sg13g2_fill_1 FILLER_71_590 ();
 sg13g2_fill_2 FILLER_71_603 ();
 sg13g2_fill_2 FILLER_71_632 ();
 sg13g2_fill_2 FILLER_71_660 ();
 sg13g2_decap_8 FILLER_71_688 ();
 sg13g2_decap_8 FILLER_71_695 ();
 sg13g2_decap_8 FILLER_71_702 ();
 sg13g2_decap_8 FILLER_71_709 ();
 sg13g2_decap_8 FILLER_71_716 ();
 sg13g2_decap_8 FILLER_71_723 ();
 sg13g2_decap_8 FILLER_71_730 ();
 sg13g2_decap_8 FILLER_71_737 ();
 sg13g2_decap_8 FILLER_71_744 ();
 sg13g2_decap_8 FILLER_71_751 ();
 sg13g2_decap_8 FILLER_71_758 ();
 sg13g2_decap_8 FILLER_71_765 ();
 sg13g2_decap_8 FILLER_71_772 ();
 sg13g2_decap_8 FILLER_71_779 ();
 sg13g2_decap_8 FILLER_71_786 ();
 sg13g2_decap_8 FILLER_71_793 ();
 sg13g2_decap_8 FILLER_71_800 ();
 sg13g2_decap_8 FILLER_71_807 ();
 sg13g2_decap_8 FILLER_71_814 ();
 sg13g2_decap_8 FILLER_71_821 ();
 sg13g2_decap_8 FILLER_71_828 ();
 sg13g2_decap_8 FILLER_71_835 ();
 sg13g2_decap_8 FILLER_71_842 ();
 sg13g2_decap_8 FILLER_71_849 ();
 sg13g2_decap_4 FILLER_71_856 ();
 sg13g2_fill_2 FILLER_71_860 ();
 sg13g2_fill_1 FILLER_72_0 ();
 sg13g2_fill_1 FILLER_72_55 ();
 sg13g2_decap_4 FILLER_72_82 ();
 sg13g2_fill_1 FILLER_72_86 ();
 sg13g2_fill_1 FILLER_72_113 ();
 sg13g2_fill_1 FILLER_72_122 ();
 sg13g2_fill_2 FILLER_72_138 ();
 sg13g2_fill_2 FILLER_72_165 ();
 sg13g2_fill_1 FILLER_72_167 ();
 sg13g2_fill_1 FILLER_72_245 ();
 sg13g2_fill_1 FILLER_72_255 ();
 sg13g2_fill_2 FILLER_72_297 ();
 sg13g2_fill_1 FILLER_72_299 ();
 sg13g2_fill_1 FILLER_72_304 ();
 sg13g2_fill_2 FILLER_72_317 ();
 sg13g2_fill_1 FILLER_72_319 ();
 sg13g2_fill_1 FILLER_72_418 ();
 sg13g2_decap_4 FILLER_72_449 ();
 sg13g2_fill_1 FILLER_72_492 ();
 sg13g2_decap_8 FILLER_72_524 ();
 sg13g2_decap_8 FILLER_72_531 ();
 sg13g2_decap_8 FILLER_72_554 ();
 sg13g2_decap_8 FILLER_72_561 ();
 sg13g2_decap_8 FILLER_72_577 ();
 sg13g2_decap_8 FILLER_72_584 ();
 sg13g2_fill_1 FILLER_72_591 ();
 sg13g2_fill_2 FILLER_72_597 ();
 sg13g2_decap_4 FILLER_72_631 ();
 sg13g2_fill_2 FILLER_72_635 ();
 sg13g2_fill_2 FILLER_72_663 ();
 sg13g2_fill_1 FILLER_72_686 ();
 sg13g2_decap_8 FILLER_72_711 ();
 sg13g2_decap_8 FILLER_72_718 ();
 sg13g2_decap_8 FILLER_72_725 ();
 sg13g2_decap_8 FILLER_72_732 ();
 sg13g2_decap_8 FILLER_72_739 ();
 sg13g2_decap_8 FILLER_72_746 ();
 sg13g2_decap_8 FILLER_72_753 ();
 sg13g2_decap_8 FILLER_72_760 ();
 sg13g2_decap_8 FILLER_72_767 ();
 sg13g2_decap_8 FILLER_72_774 ();
 sg13g2_decap_8 FILLER_72_781 ();
 sg13g2_decap_8 FILLER_72_788 ();
 sg13g2_decap_8 FILLER_72_795 ();
 sg13g2_decap_8 FILLER_72_802 ();
 sg13g2_decap_8 FILLER_72_809 ();
 sg13g2_decap_8 FILLER_72_816 ();
 sg13g2_decap_8 FILLER_72_823 ();
 sg13g2_decap_8 FILLER_72_830 ();
 sg13g2_decap_8 FILLER_72_837 ();
 sg13g2_decap_8 FILLER_72_844 ();
 sg13g2_decap_8 FILLER_72_851 ();
 sg13g2_decap_4 FILLER_72_858 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_4 FILLER_73_7 ();
 sg13g2_decap_4 FILLER_73_15 ();
 sg13g2_fill_1 FILLER_73_19 ();
 sg13g2_decap_4 FILLER_73_40 ();
 sg13g2_fill_2 FILLER_73_65 ();
 sg13g2_decap_4 FILLER_73_71 ();
 sg13g2_decap_8 FILLER_73_110 ();
 sg13g2_decap_8 FILLER_73_117 ();
 sg13g2_fill_2 FILLER_73_124 ();
 sg13g2_fill_1 FILLER_73_126 ();
 sg13g2_decap_4 FILLER_73_153 ();
 sg13g2_fill_2 FILLER_73_172 ();
 sg13g2_fill_1 FILLER_73_174 ();
 sg13g2_fill_2 FILLER_73_193 ();
 sg13g2_fill_1 FILLER_73_195 ();
 sg13g2_decap_8 FILLER_73_200 ();
 sg13g2_fill_1 FILLER_73_207 ();
 sg13g2_fill_2 FILLER_73_237 ();
 sg13g2_fill_2 FILLER_73_329 ();
 sg13g2_fill_1 FILLER_73_331 ();
 sg13g2_decap_8 FILLER_73_367 ();
 sg13g2_decap_4 FILLER_73_374 ();
 sg13g2_fill_2 FILLER_73_378 ();
 sg13g2_fill_2 FILLER_73_384 ();
 sg13g2_fill_1 FILLER_73_386 ();
 sg13g2_fill_1 FILLER_73_401 ();
 sg13g2_fill_2 FILLER_73_417 ();
 sg13g2_fill_1 FILLER_73_419 ();
 sg13g2_decap_8 FILLER_73_457 ();
 sg13g2_decap_4 FILLER_73_464 ();
 sg13g2_fill_2 FILLER_73_502 ();
 sg13g2_fill_2 FILLER_73_561 ();
 sg13g2_decap_4 FILLER_73_567 ();
 sg13g2_fill_1 FILLER_73_571 ();
 sg13g2_fill_2 FILLER_73_577 ();
 sg13g2_fill_1 FILLER_73_579 ();
 sg13g2_decap_8 FILLER_73_600 ();
 sg13g2_decap_8 FILLER_73_607 ();
 sg13g2_fill_2 FILLER_73_614 ();
 sg13g2_fill_1 FILLER_73_634 ();
 sg13g2_fill_2 FILLER_73_643 ();
 sg13g2_decap_8 FILLER_73_653 ();
 sg13g2_decap_8 FILLER_73_660 ();
 sg13g2_decap_4 FILLER_73_667 ();
 sg13g2_decap_8 FILLER_73_692 ();
 sg13g2_decap_8 FILLER_73_699 ();
 sg13g2_decap_8 FILLER_73_706 ();
 sg13g2_decap_8 FILLER_73_713 ();
 sg13g2_decap_8 FILLER_73_720 ();
 sg13g2_decap_8 FILLER_73_727 ();
 sg13g2_decap_8 FILLER_73_734 ();
 sg13g2_decap_8 FILLER_73_741 ();
 sg13g2_decap_8 FILLER_73_748 ();
 sg13g2_decap_8 FILLER_73_755 ();
 sg13g2_decap_8 FILLER_73_762 ();
 sg13g2_decap_8 FILLER_73_769 ();
 sg13g2_decap_8 FILLER_73_776 ();
 sg13g2_decap_8 FILLER_73_783 ();
 sg13g2_decap_8 FILLER_73_790 ();
 sg13g2_decap_8 FILLER_73_797 ();
 sg13g2_decap_8 FILLER_73_804 ();
 sg13g2_decap_8 FILLER_73_811 ();
 sg13g2_decap_8 FILLER_73_818 ();
 sg13g2_decap_8 FILLER_73_825 ();
 sg13g2_decap_8 FILLER_73_832 ();
 sg13g2_decap_8 FILLER_73_839 ();
 sg13g2_decap_8 FILLER_73_846 ();
 sg13g2_decap_8 FILLER_73_853 ();
 sg13g2_fill_2 FILLER_73_860 ();
 sg13g2_fill_2 FILLER_74_26 ();
 sg13g2_fill_2 FILLER_74_90 ();
 sg13g2_decap_4 FILLER_74_159 ();
 sg13g2_decap_4 FILLER_74_207 ();
 sg13g2_fill_2 FILLER_74_321 ();
 sg13g2_fill_1 FILLER_74_323 ();
 sg13g2_decap_4 FILLER_74_344 ();
 sg13g2_fill_1 FILLER_74_361 ();
 sg13g2_fill_1 FILLER_74_398 ();
 sg13g2_fill_1 FILLER_74_407 ();
 sg13g2_fill_2 FILLER_74_445 ();
 sg13g2_fill_2 FILLER_74_473 ();
 sg13g2_fill_1 FILLER_74_481 ();
 sg13g2_decap_8 FILLER_74_503 ();
 sg13g2_fill_1 FILLER_74_523 ();
 sg13g2_decap_8 FILLER_74_529 ();
 sg13g2_fill_2 FILLER_74_536 ();
 sg13g2_fill_1 FILLER_74_538 ();
 sg13g2_decap_4 FILLER_74_548 ();
 sg13g2_decap_4 FILLER_74_594 ();
 sg13g2_fill_1 FILLER_74_602 ();
 sg13g2_fill_1 FILLER_74_611 ();
 sg13g2_decap_4 FILLER_74_638 ();
 sg13g2_fill_2 FILLER_74_642 ();
 sg13g2_decap_8 FILLER_74_698 ();
 sg13g2_decap_8 FILLER_74_705 ();
 sg13g2_decap_8 FILLER_74_712 ();
 sg13g2_decap_8 FILLER_74_719 ();
 sg13g2_decap_8 FILLER_74_726 ();
 sg13g2_decap_8 FILLER_74_733 ();
 sg13g2_decap_8 FILLER_74_740 ();
 sg13g2_decap_8 FILLER_74_747 ();
 sg13g2_decap_8 FILLER_74_754 ();
 sg13g2_decap_8 FILLER_74_761 ();
 sg13g2_decap_8 FILLER_74_768 ();
 sg13g2_decap_8 FILLER_74_775 ();
 sg13g2_decap_8 FILLER_74_782 ();
 sg13g2_decap_8 FILLER_74_789 ();
 sg13g2_decap_8 FILLER_74_796 ();
 sg13g2_decap_8 FILLER_74_803 ();
 sg13g2_decap_8 FILLER_74_810 ();
 sg13g2_decap_8 FILLER_74_817 ();
 sg13g2_decap_8 FILLER_74_824 ();
 sg13g2_decap_8 FILLER_74_831 ();
 sg13g2_decap_8 FILLER_74_838 ();
 sg13g2_decap_8 FILLER_74_845 ();
 sg13g2_decap_8 FILLER_74_852 ();
 sg13g2_fill_2 FILLER_74_859 ();
 sg13g2_fill_1 FILLER_74_861 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_fill_2 FILLER_75_7 ();
 sg13g2_fill_1 FILLER_75_9 ();
 sg13g2_decap_8 FILLER_75_47 ();
 sg13g2_decap_8 FILLER_75_54 ();
 sg13g2_fill_2 FILLER_75_61 ();
 sg13g2_fill_1 FILLER_75_63 ();
 sg13g2_fill_1 FILLER_75_107 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_fill_2 FILLER_75_126 ();
 sg13g2_fill_1 FILLER_75_128 ();
 sg13g2_fill_1 FILLER_75_133 ();
 sg13g2_fill_2 FILLER_75_188 ();
 sg13g2_fill_1 FILLER_75_190 ();
 sg13g2_fill_2 FILLER_75_217 ();
 sg13g2_fill_1 FILLER_75_219 ();
 sg13g2_fill_1 FILLER_75_233 ();
 sg13g2_fill_1 FILLER_75_260 ();
 sg13g2_fill_2 FILLER_75_289 ();
 sg13g2_fill_1 FILLER_75_291 ();
 sg13g2_fill_2 FILLER_75_332 ();
 sg13g2_fill_1 FILLER_75_360 ();
 sg13g2_fill_2 FILLER_75_370 ();
 sg13g2_fill_2 FILLER_75_386 ();
 sg13g2_fill_2 FILLER_75_405 ();
 sg13g2_fill_2 FILLER_75_415 ();
 sg13g2_fill_1 FILLER_75_417 ();
 sg13g2_fill_2 FILLER_75_427 ();
 sg13g2_fill_1 FILLER_75_439 ();
 sg13g2_fill_1 FILLER_75_457 ();
 sg13g2_decap_8 FILLER_75_462 ();
 sg13g2_decap_8 FILLER_75_469 ();
 sg13g2_fill_2 FILLER_75_495 ();
 sg13g2_fill_1 FILLER_75_497 ();
 sg13g2_fill_2 FILLER_75_510 ();
 sg13g2_decap_8 FILLER_75_540 ();
 sg13g2_fill_2 FILLER_75_547 ();
 sg13g2_decap_8 FILLER_75_566 ();
 sg13g2_fill_2 FILLER_75_573 ();
 sg13g2_fill_1 FILLER_75_575 ();
 sg13g2_decap_8 FILLER_75_580 ();
 sg13g2_fill_1 FILLER_75_613 ();
 sg13g2_decap_8 FILLER_75_630 ();
 sg13g2_decap_8 FILLER_75_637 ();
 sg13g2_decap_8 FILLER_75_644 ();
 sg13g2_fill_2 FILLER_75_651 ();
 sg13g2_fill_1 FILLER_75_653 ();
 sg13g2_decap_4 FILLER_75_658 ();
 sg13g2_decap_8 FILLER_75_670 ();
 sg13g2_decap_8 FILLER_75_677 ();
 sg13g2_fill_1 FILLER_75_684 ();
 sg13g2_decap_8 FILLER_75_697 ();
 sg13g2_decap_8 FILLER_75_704 ();
 sg13g2_decap_8 FILLER_75_711 ();
 sg13g2_decap_8 FILLER_75_718 ();
 sg13g2_decap_8 FILLER_75_725 ();
 sg13g2_decap_8 FILLER_75_732 ();
 sg13g2_decap_8 FILLER_75_739 ();
 sg13g2_decap_8 FILLER_75_746 ();
 sg13g2_decap_8 FILLER_75_753 ();
 sg13g2_decap_8 FILLER_75_760 ();
 sg13g2_decap_8 FILLER_75_767 ();
 sg13g2_decap_8 FILLER_75_774 ();
 sg13g2_decap_8 FILLER_75_781 ();
 sg13g2_decap_8 FILLER_75_788 ();
 sg13g2_decap_8 FILLER_75_795 ();
 sg13g2_decap_8 FILLER_75_802 ();
 sg13g2_decap_8 FILLER_75_809 ();
 sg13g2_decap_8 FILLER_75_816 ();
 sg13g2_decap_8 FILLER_75_823 ();
 sg13g2_decap_8 FILLER_75_830 ();
 sg13g2_decap_8 FILLER_75_837 ();
 sg13g2_decap_8 FILLER_75_844 ();
 sg13g2_decap_8 FILLER_75_851 ();
 sg13g2_decap_4 FILLER_75_858 ();
 sg13g2_fill_2 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_2 ();
 sg13g2_decap_4 FILLER_76_86 ();
 sg13g2_fill_2 FILLER_76_90 ();
 sg13g2_decap_8 FILLER_76_128 ();
 sg13g2_decap_4 FILLER_76_135 ();
 sg13g2_fill_2 FILLER_76_154 ();
 sg13g2_fill_2 FILLER_76_171 ();
 sg13g2_fill_1 FILLER_76_173 ();
 sg13g2_fill_2 FILLER_76_183 ();
 sg13g2_fill_2 FILLER_76_190 ();
 sg13g2_fill_1 FILLER_76_192 ();
 sg13g2_decap_8 FILLER_76_215 ();
 sg13g2_fill_1 FILLER_76_222 ();
 sg13g2_fill_1 FILLER_76_249 ();
 sg13g2_fill_1 FILLER_76_268 ();
 sg13g2_fill_1 FILLER_76_275 ();
 sg13g2_fill_2 FILLER_76_310 ();
 sg13g2_fill_2 FILLER_76_318 ();
 sg13g2_fill_1 FILLER_76_320 ();
 sg13g2_fill_2 FILLER_76_339 ();
 sg13g2_fill_2 FILLER_76_377 ();
 sg13g2_decap_8 FILLER_76_405 ();
 sg13g2_fill_2 FILLER_76_417 ();
 sg13g2_fill_1 FILLER_76_444 ();
 sg13g2_decap_8 FILLER_76_455 ();
 sg13g2_decap_8 FILLER_76_462 ();
 sg13g2_fill_2 FILLER_76_469 ();
 sg13g2_fill_1 FILLER_76_471 ();
 sg13g2_fill_2 FILLER_76_481 ();
 sg13g2_fill_1 FILLER_76_483 ();
 sg13g2_fill_2 FILLER_76_488 ();
 sg13g2_fill_1 FILLER_76_490 ();
 sg13g2_decap_8 FILLER_76_504 ();
 sg13g2_decap_8 FILLER_76_511 ();
 sg13g2_decap_4 FILLER_76_518 ();
 sg13g2_decap_4 FILLER_76_530 ();
 sg13g2_fill_2 FILLER_76_534 ();
 sg13g2_decap_4 FILLER_76_562 ();
 sg13g2_decap_8 FILLER_76_592 ();
 sg13g2_decap_4 FILLER_76_599 ();
 sg13g2_fill_1 FILLER_76_603 ();
 sg13g2_decap_8 FILLER_76_609 ();
 sg13g2_fill_2 FILLER_76_616 ();
 sg13g2_fill_1 FILLER_76_618 ();
 sg13g2_fill_1 FILLER_76_627 ();
 sg13g2_decap_4 FILLER_76_648 ();
 sg13g2_fill_2 FILLER_76_652 ();
 sg13g2_decap_8 FILLER_76_659 ();
 sg13g2_decap_8 FILLER_76_666 ();
 sg13g2_fill_2 FILLER_76_673 ();
 sg13g2_fill_1 FILLER_76_675 ();
 sg13g2_decap_8 FILLER_76_689 ();
 sg13g2_decap_8 FILLER_76_696 ();
 sg13g2_decap_8 FILLER_76_703 ();
 sg13g2_decap_8 FILLER_76_710 ();
 sg13g2_decap_8 FILLER_76_717 ();
 sg13g2_decap_8 FILLER_76_724 ();
 sg13g2_decap_8 FILLER_76_731 ();
 sg13g2_decap_8 FILLER_76_738 ();
 sg13g2_decap_8 FILLER_76_745 ();
 sg13g2_decap_8 FILLER_76_752 ();
 sg13g2_decap_8 FILLER_76_759 ();
 sg13g2_decap_8 FILLER_76_766 ();
 sg13g2_decap_8 FILLER_76_773 ();
 sg13g2_decap_8 FILLER_76_780 ();
 sg13g2_decap_8 FILLER_76_787 ();
 sg13g2_decap_8 FILLER_76_794 ();
 sg13g2_decap_8 FILLER_76_801 ();
 sg13g2_decap_8 FILLER_76_808 ();
 sg13g2_decap_8 FILLER_76_815 ();
 sg13g2_decap_8 FILLER_76_822 ();
 sg13g2_decap_8 FILLER_76_829 ();
 sg13g2_decap_8 FILLER_76_836 ();
 sg13g2_decap_8 FILLER_76_843 ();
 sg13g2_decap_8 FILLER_76_850 ();
 sg13g2_decap_4 FILLER_76_857 ();
 sg13g2_fill_1 FILLER_76_861 ();
 sg13g2_decap_4 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_30 ();
 sg13g2_fill_2 FILLER_77_42 ();
 sg13g2_fill_1 FILLER_77_61 ();
 sg13g2_fill_2 FILLER_77_66 ();
 sg13g2_fill_1 FILLER_77_68 ();
 sg13g2_decap_4 FILLER_77_122 ();
 sg13g2_fill_2 FILLER_77_126 ();
 sg13g2_fill_2 FILLER_77_159 ();
 sg13g2_fill_1 FILLER_77_161 ();
 sg13g2_fill_1 FILLER_77_188 ();
 sg13g2_fill_2 FILLER_77_225 ();
 sg13g2_fill_2 FILLER_77_232 ();
 sg13g2_fill_2 FILLER_77_246 ();
 sg13g2_fill_1 FILLER_77_248 ();
 sg13g2_fill_1 FILLER_77_267 ();
 sg13g2_fill_1 FILLER_77_273 ();
 sg13g2_fill_1 FILLER_77_300 ();
 sg13g2_fill_1 FILLER_77_357 ();
 sg13g2_decap_8 FILLER_77_372 ();
 sg13g2_decap_4 FILLER_77_392 ();
 sg13g2_fill_2 FILLER_77_396 ();
 sg13g2_decap_8 FILLER_77_429 ();
 sg13g2_fill_2 FILLER_77_436 ();
 sg13g2_fill_2 FILLER_77_462 ();
 sg13g2_fill_2 FILLER_77_484 ();
 sg13g2_fill_1 FILLER_77_486 ();
 sg13g2_fill_1 FILLER_77_511 ();
 sg13g2_fill_1 FILLER_77_516 ();
 sg13g2_decap_8 FILLER_77_539 ();
 sg13g2_decap_4 FILLER_77_546 ();
 sg13g2_fill_2 FILLER_77_558 ();
 sg13g2_decap_8 FILLER_77_568 ();
 sg13g2_fill_2 FILLER_77_575 ();
 sg13g2_fill_2 FILLER_77_629 ();
 sg13g2_decap_8 FILLER_77_665 ();
 sg13g2_decap_8 FILLER_77_672 ();
 sg13g2_decap_8 FILLER_77_679 ();
 sg13g2_decap_8 FILLER_77_686 ();
 sg13g2_decap_8 FILLER_77_693 ();
 sg13g2_decap_8 FILLER_77_700 ();
 sg13g2_decap_8 FILLER_77_707 ();
 sg13g2_decap_8 FILLER_77_714 ();
 sg13g2_decap_8 FILLER_77_721 ();
 sg13g2_decap_8 FILLER_77_728 ();
 sg13g2_decap_8 FILLER_77_735 ();
 sg13g2_decap_8 FILLER_77_742 ();
 sg13g2_decap_8 FILLER_77_749 ();
 sg13g2_decap_8 FILLER_77_756 ();
 sg13g2_decap_8 FILLER_77_763 ();
 sg13g2_decap_8 FILLER_77_770 ();
 sg13g2_decap_8 FILLER_77_777 ();
 sg13g2_decap_8 FILLER_77_784 ();
 sg13g2_decap_8 FILLER_77_791 ();
 sg13g2_decap_8 FILLER_77_798 ();
 sg13g2_decap_8 FILLER_77_805 ();
 sg13g2_decap_8 FILLER_77_812 ();
 sg13g2_decap_8 FILLER_77_819 ();
 sg13g2_decap_8 FILLER_77_826 ();
 sg13g2_decap_8 FILLER_77_833 ();
 sg13g2_decap_8 FILLER_77_840 ();
 sg13g2_decap_8 FILLER_77_847 ();
 sg13g2_decap_8 FILLER_77_854 ();
 sg13g2_fill_1 FILLER_77_861 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_2 ();
 sg13g2_decap_4 FILLER_78_29 ();
 sg13g2_fill_2 FILLER_78_33 ();
 sg13g2_fill_1 FILLER_78_71 ();
 sg13g2_decap_4 FILLER_78_76 ();
 sg13g2_decap_4 FILLER_78_129 ();
 sg13g2_fill_1 FILLER_78_133 ();
 sg13g2_fill_2 FILLER_78_174 ();
 sg13g2_fill_2 FILLER_78_186 ();
 sg13g2_decap_4 FILLER_78_221 ();
 sg13g2_fill_2 FILLER_78_225 ();
 sg13g2_fill_1 FILLER_78_253 ();
 sg13g2_fill_1 FILLER_78_308 ();
 sg13g2_fill_2 FILLER_78_364 ();
 sg13g2_fill_1 FILLER_78_366 ();
 sg13g2_decap_4 FILLER_78_401 ();
 sg13g2_fill_2 FILLER_78_418 ();
 sg13g2_fill_2 FILLER_78_445 ();
 sg13g2_fill_1 FILLER_78_447 ();
 sg13g2_fill_1 FILLER_78_452 ();
 sg13g2_fill_2 FILLER_78_477 ();
 sg13g2_fill_1 FILLER_78_479 ();
 sg13g2_fill_2 FILLER_78_496 ();
 sg13g2_decap_4 FILLER_78_507 ();
 sg13g2_fill_2 FILLER_78_511 ();
 sg13g2_decap_8 FILLER_78_529 ();
 sg13g2_decap_8 FILLER_78_567 ();
 sg13g2_decap_8 FILLER_78_574 ();
 sg13g2_decap_8 FILLER_78_581 ();
 sg13g2_decap_8 FILLER_78_592 ();
 sg13g2_fill_1 FILLER_78_599 ();
 sg13g2_decap_4 FILLER_78_605 ();
 sg13g2_decap_8 FILLER_78_613 ();
 sg13g2_fill_1 FILLER_78_625 ();
 sg13g2_decap_8 FILLER_78_630 ();
 sg13g2_decap_8 FILLER_78_637 ();
 sg13g2_fill_1 FILLER_78_644 ();
 sg13g2_decap_8 FILLER_78_658 ();
 sg13g2_decap_8 FILLER_78_665 ();
 sg13g2_decap_8 FILLER_78_672 ();
 sg13g2_decap_8 FILLER_78_679 ();
 sg13g2_decap_8 FILLER_78_686 ();
 sg13g2_decap_8 FILLER_78_693 ();
 sg13g2_decap_8 FILLER_78_700 ();
 sg13g2_decap_8 FILLER_78_707 ();
 sg13g2_decap_8 FILLER_78_714 ();
 sg13g2_decap_8 FILLER_78_721 ();
 sg13g2_decap_8 FILLER_78_728 ();
 sg13g2_decap_8 FILLER_78_735 ();
 sg13g2_decap_8 FILLER_78_742 ();
 sg13g2_decap_8 FILLER_78_749 ();
 sg13g2_decap_8 FILLER_78_756 ();
 sg13g2_decap_8 FILLER_78_763 ();
 sg13g2_decap_8 FILLER_78_770 ();
 sg13g2_decap_8 FILLER_78_777 ();
 sg13g2_decap_8 FILLER_78_784 ();
 sg13g2_decap_8 FILLER_78_791 ();
 sg13g2_decap_8 FILLER_78_798 ();
 sg13g2_decap_8 FILLER_78_805 ();
 sg13g2_decap_8 FILLER_78_812 ();
 sg13g2_decap_8 FILLER_78_819 ();
 sg13g2_decap_8 FILLER_78_826 ();
 sg13g2_decap_8 FILLER_78_833 ();
 sg13g2_decap_8 FILLER_78_840 ();
 sg13g2_decap_8 FILLER_78_847 ();
 sg13g2_decap_8 FILLER_78_854 ();
 sg13g2_fill_1 FILLER_78_861 ();
 sg13g2_fill_2 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_2 ();
 sg13g2_fill_2 FILLER_79_49 ();
 sg13g2_fill_1 FILLER_79_78 ();
 sg13g2_fill_1 FILLER_79_100 ();
 sg13g2_fill_2 FILLER_79_342 ();
 sg13g2_fill_2 FILLER_79_362 ();
 sg13g2_fill_1 FILLER_79_364 ();
 sg13g2_fill_1 FILLER_79_375 ();
 sg13g2_decap_4 FILLER_79_397 ();
 sg13g2_fill_1 FILLER_79_427 ();
 sg13g2_fill_1 FILLER_79_440 ();
 sg13g2_fill_1 FILLER_79_446 ();
 sg13g2_fill_1 FILLER_79_464 ();
 sg13g2_fill_2 FILLER_79_494 ();
 sg13g2_decap_4 FILLER_79_512 ();
 sg13g2_decap_8 FILLER_79_539 ();
 sg13g2_fill_1 FILLER_79_546 ();
 sg13g2_decap_8 FILLER_79_556 ();
 sg13g2_decap_4 FILLER_79_563 ();
 sg13g2_fill_1 FILLER_79_567 ();
 sg13g2_decap_8 FILLER_79_602 ();
 sg13g2_decap_4 FILLER_79_609 ();
 sg13g2_fill_2 FILLER_79_613 ();
 sg13g2_decap_8 FILLER_79_641 ();
 sg13g2_decap_8 FILLER_79_648 ();
 sg13g2_decap_8 FILLER_79_655 ();
 sg13g2_decap_8 FILLER_79_662 ();
 sg13g2_decap_8 FILLER_79_669 ();
 sg13g2_decap_8 FILLER_79_676 ();
 sg13g2_decap_8 FILLER_79_683 ();
 sg13g2_decap_8 FILLER_79_690 ();
 sg13g2_decap_8 FILLER_79_697 ();
 sg13g2_decap_8 FILLER_79_704 ();
 sg13g2_decap_8 FILLER_79_711 ();
 sg13g2_decap_8 FILLER_79_718 ();
 sg13g2_decap_8 FILLER_79_725 ();
 sg13g2_decap_8 FILLER_79_732 ();
 sg13g2_decap_8 FILLER_79_739 ();
 sg13g2_decap_8 FILLER_79_746 ();
 sg13g2_decap_8 FILLER_79_753 ();
 sg13g2_decap_8 FILLER_79_760 ();
 sg13g2_decap_8 FILLER_79_767 ();
 sg13g2_decap_8 FILLER_79_774 ();
 sg13g2_decap_8 FILLER_79_781 ();
 sg13g2_decap_8 FILLER_79_788 ();
 sg13g2_decap_8 FILLER_79_795 ();
 sg13g2_decap_8 FILLER_79_802 ();
 sg13g2_decap_8 FILLER_79_809 ();
 sg13g2_decap_8 FILLER_79_816 ();
 sg13g2_decap_8 FILLER_79_823 ();
 sg13g2_decap_8 FILLER_79_830 ();
 sg13g2_decap_8 FILLER_79_837 ();
 sg13g2_decap_8 FILLER_79_844 ();
 sg13g2_decap_8 FILLER_79_851 ();
 sg13g2_decap_4 FILLER_79_858 ();
 sg13g2_fill_2 FILLER_80_0 ();
 sg13g2_fill_2 FILLER_80_34 ();
 sg13g2_fill_2 FILLER_80_106 ();
 sg13g2_fill_1 FILLER_80_108 ();
 sg13g2_fill_1 FILLER_80_135 ();
 sg13g2_fill_1 FILLER_80_149 ();
 sg13g2_fill_1 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_182 ();
 sg13g2_fill_1 FILLER_80_186 ();
 sg13g2_fill_2 FILLER_80_200 ();
 sg13g2_fill_2 FILLER_80_211 ();
 sg13g2_decap_8 FILLER_80_217 ();
 sg13g2_fill_2 FILLER_80_224 ();
 sg13g2_fill_1 FILLER_80_226 ();
 sg13g2_fill_2 FILLER_80_262 ();
 sg13g2_fill_2 FILLER_80_293 ();
 sg13g2_fill_1 FILLER_80_295 ();
 sg13g2_fill_2 FILLER_80_301 ();
 sg13g2_fill_1 FILLER_80_303 ();
 sg13g2_fill_2 FILLER_80_309 ();
 sg13g2_fill_1 FILLER_80_311 ();
 sg13g2_fill_2 FILLER_80_325 ();
 sg13g2_fill_2 FILLER_80_336 ();
 sg13g2_fill_1 FILLER_80_372 ();
 sg13g2_decap_4 FILLER_80_399 ();
 sg13g2_fill_2 FILLER_80_403 ();
 sg13g2_fill_2 FILLER_80_409 ();
 sg13g2_decap_8 FILLER_80_419 ();
 sg13g2_decap_8 FILLER_80_426 ();
 sg13g2_decap_8 FILLER_80_433 ();
 sg13g2_decap_8 FILLER_80_457 ();
 sg13g2_decap_8 FILLER_80_464 ();
 sg13g2_fill_2 FILLER_80_471 ();
 sg13g2_fill_1 FILLER_80_473 ();
 sg13g2_fill_1 FILLER_80_478 ();
 sg13g2_fill_2 FILLER_80_485 ();
 sg13g2_decap_4 FILLER_80_492 ();
 sg13g2_fill_2 FILLER_80_496 ();
 sg13g2_decap_8 FILLER_80_507 ();
 sg13g2_fill_1 FILLER_80_514 ();
 sg13g2_fill_1 FILLER_80_523 ();
 sg13g2_decap_4 FILLER_80_550 ();
 sg13g2_fill_2 FILLER_80_554 ();
 sg13g2_decap_8 FILLER_80_590 ();
 sg13g2_decap_8 FILLER_80_597 ();
 sg13g2_decap_8 FILLER_80_604 ();
 sg13g2_decap_8 FILLER_80_611 ();
 sg13g2_decap_8 FILLER_80_618 ();
 sg13g2_decap_8 FILLER_80_625 ();
 sg13g2_decap_8 FILLER_80_632 ();
 sg13g2_decap_8 FILLER_80_639 ();
 sg13g2_decap_8 FILLER_80_646 ();
 sg13g2_decap_8 FILLER_80_653 ();
 sg13g2_decap_8 FILLER_80_660 ();
 sg13g2_decap_8 FILLER_80_667 ();
 sg13g2_decap_8 FILLER_80_674 ();
 sg13g2_decap_8 FILLER_80_681 ();
 sg13g2_decap_8 FILLER_80_688 ();
 sg13g2_decap_8 FILLER_80_695 ();
 sg13g2_decap_8 FILLER_80_702 ();
 sg13g2_decap_8 FILLER_80_709 ();
 sg13g2_decap_8 FILLER_80_716 ();
 sg13g2_decap_8 FILLER_80_723 ();
 sg13g2_decap_8 FILLER_80_730 ();
 sg13g2_decap_8 FILLER_80_737 ();
 sg13g2_decap_8 FILLER_80_744 ();
 sg13g2_decap_8 FILLER_80_751 ();
 sg13g2_decap_8 FILLER_80_758 ();
 sg13g2_decap_8 FILLER_80_765 ();
 sg13g2_decap_8 FILLER_80_772 ();
 sg13g2_decap_8 FILLER_80_779 ();
 sg13g2_decap_8 FILLER_80_786 ();
 sg13g2_decap_8 FILLER_80_793 ();
 sg13g2_decap_8 FILLER_80_800 ();
 sg13g2_decap_8 FILLER_80_807 ();
 sg13g2_decap_8 FILLER_80_814 ();
 sg13g2_decap_8 FILLER_80_821 ();
 sg13g2_decap_8 FILLER_80_828 ();
 sg13g2_decap_8 FILLER_80_835 ();
 sg13g2_decap_8 FILLER_80_842 ();
 sg13g2_decap_8 FILLER_80_849 ();
 sg13g2_decap_4 FILLER_80_856 ();
 sg13g2_fill_2 FILLER_80_860 ();
 assign uio_oe[4] = net405;
 assign uio_oe[5] = net406;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net8;
 assign uio_out[6] = net9;
 assign uio_out[7] = net10;
endmodule

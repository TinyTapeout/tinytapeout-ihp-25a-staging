module tt_um_cfib_demo (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire hsync;
 wire pwm;
 wire \top_inst.pwm_inst.cntr[0] ;
 wire \top_inst.pwm_inst.cntr[1] ;
 wire \top_inst.pwm_inst.cntr[2] ;
 wire \top_inst.pwm_inst.cntr[3] ;
 wire \top_inst.sample_ena ;
 wire \top_inst.sndgen_inst.bar_counter[0] ;
 wire \top_inst.sndgen_inst.bar_counter[1] ;
 wire \top_inst.sndgen_inst.bar_counter[2] ;
 wire \top_inst.sndgen_inst.bar_counter[3] ;
 wire \top_inst.sndgen_inst.c1[0] ;
 wire \top_inst.sndgen_inst.c1[1] ;
 wire \top_inst.sndgen_inst.c2[0] ;
 wire \top_inst.sndgen_inst.c2[1] ;
 wire \top_inst.sndgen_inst.c2[2] ;
 wire \top_inst.sndgen_inst.c3[0] ;
 wire \top_inst.sndgen_inst.c3[1] ;
 wire \top_inst.sndgen_inst.c3[2] ;
 wire \top_inst.sndgen_inst.c4[2] ;
 wire \top_inst.sndgen_inst.lfsr[0] ;
 wire \top_inst.sndgen_inst.lfsr[1] ;
 wire \top_inst.sndgen_inst.lfsr[2] ;
 wire \top_inst.sndgen_inst.lfsr[3] ;
 wire \top_inst.sndgen_inst.lfsr[4] ;
 wire \top_inst.sndgen_inst.lfsr[5] ;
 wire \top_inst.sndgen_inst.lfsr[6] ;
 wire \top_inst.sndgen_inst.lfsr[7] ;
 wire \top_inst.sndgen_inst.mask_1[0] ;
 wire \top_inst.sndgen_inst.mask_1[1] ;
 wire \top_inst.sndgen_inst.mask_1[2] ;
 wire \top_inst.sndgen_inst.mask_1[3] ;
 wire \top_inst.sndgen_inst.mask_2 ;
 wire \top_inst.sndgen_inst.p_c2[0] ;
 wire \top_inst.sndgen_inst.p_c2[10] ;
 wire \top_inst.sndgen_inst.p_c2[1] ;
 wire \top_inst.sndgen_inst.p_c2[2] ;
 wire \top_inst.sndgen_inst.p_c2[3] ;
 wire \top_inst.sndgen_inst.p_c2[4] ;
 wire \top_inst.sndgen_inst.p_c2[5] ;
 wire \top_inst.sndgen_inst.p_c2[6] ;
 wire \top_inst.sndgen_inst.p_c2[7] ;
 wire \top_inst.sndgen_inst.p_c3[0] ;
 wire \top_inst.sndgen_inst.p_c3[10] ;
 wire \top_inst.sndgen_inst.p_c3[1] ;
 wire \top_inst.sndgen_inst.p_c3[2] ;
 wire \top_inst.sndgen_inst.p_c3[3] ;
 wire \top_inst.sndgen_inst.p_c3[4] ;
 wire \top_inst.sndgen_inst.p_c3[5] ;
 wire \top_inst.sndgen_inst.p_c3[6] ;
 wire \top_inst.sndgen_inst.p_c3[7] ;
 wire \top_inst.sndgen_inst.p_c4[0] ;
 wire \top_inst.sndgen_inst.p_c4[10] ;
 wire \top_inst.sndgen_inst.p_c4[1] ;
 wire \top_inst.sndgen_inst.p_c4[2] ;
 wire \top_inst.sndgen_inst.p_c4[3] ;
 wire \top_inst.sndgen_inst.p_c4[4] ;
 wire \top_inst.sndgen_inst.p_c4[5] ;
 wire \top_inst.sndgen_inst.p_c4[6] ;
 wire \top_inst.sndgen_inst.p_c4[7] ;
 wire \top_inst.sndgen_inst.phacc2[0] ;
 wire \top_inst.sndgen_inst.phacc2[10] ;
 wire \top_inst.sndgen_inst.phacc2[11] ;
 wire \top_inst.sndgen_inst.phacc2[12] ;
 wire \top_inst.sndgen_inst.phacc2[13] ;
 wire \top_inst.sndgen_inst.phacc2[1] ;
 wire \top_inst.sndgen_inst.phacc2[2] ;
 wire \top_inst.sndgen_inst.phacc2[3] ;
 wire \top_inst.sndgen_inst.phacc2[4] ;
 wire \top_inst.sndgen_inst.phacc2[5] ;
 wire \top_inst.sndgen_inst.phacc2[6] ;
 wire \top_inst.sndgen_inst.phacc2[7] ;
 wire \top_inst.sndgen_inst.phacc2[8] ;
 wire \top_inst.sndgen_inst.phacc2[9] ;
 wire \top_inst.sndgen_inst.phacc3[0] ;
 wire \top_inst.sndgen_inst.phacc3[10] ;
 wire \top_inst.sndgen_inst.phacc3[11] ;
 wire \top_inst.sndgen_inst.phacc3[12] ;
 wire \top_inst.sndgen_inst.phacc3[13] ;
 wire \top_inst.sndgen_inst.phacc3[1] ;
 wire \top_inst.sndgen_inst.phacc3[2] ;
 wire \top_inst.sndgen_inst.phacc3[3] ;
 wire \top_inst.sndgen_inst.phacc3[4] ;
 wire \top_inst.sndgen_inst.phacc3[5] ;
 wire \top_inst.sndgen_inst.phacc3[6] ;
 wire \top_inst.sndgen_inst.phacc3[7] ;
 wire \top_inst.sndgen_inst.phacc3[8] ;
 wire \top_inst.sndgen_inst.phacc3[9] ;
 wire \top_inst.sndgen_inst.phacc4[0] ;
 wire \top_inst.sndgen_inst.phacc4[10] ;
 wire \top_inst.sndgen_inst.phacc4[11] ;
 wire \top_inst.sndgen_inst.phacc4[12] ;
 wire \top_inst.sndgen_inst.phacc4[13] ;
 wire \top_inst.sndgen_inst.phacc4[1] ;
 wire \top_inst.sndgen_inst.phacc4[2] ;
 wire \top_inst.sndgen_inst.phacc4[3] ;
 wire \top_inst.sndgen_inst.phacc4[4] ;
 wire \top_inst.sndgen_inst.phacc4[5] ;
 wire \top_inst.sndgen_inst.phacc4[6] ;
 wire \top_inst.sndgen_inst.phacc4[7] ;
 wire \top_inst.sndgen_inst.phacc4[8] ;
 wire \top_inst.sndgen_inst.phacc4[9] ;
 wire \top_inst.sndgen_inst.rom_addr[0] ;
 wire \top_inst.sndgen_inst.rom_addr[1] ;
 wire \top_inst.sndgen_inst.rom_addr[2] ;
 wire \top_inst.sndgen_inst.rom_addr[3] ;
 wire \top_inst.sndgen_inst.sample_ena_delay[0] ;
 wire \top_inst.sndgen_inst.sample_ena_delay[1] ;
 wire \top_inst.sndgen_inst.sample_ena_delay[2] ;
 wire \top_inst.sndgen_inst.slot_counter[0] ;
 wire \top_inst.sndgen_inst.slot_counter[10] ;
 wire \top_inst.sndgen_inst.slot_counter[1] ;
 wire \top_inst.sndgen_inst.slot_counter[2] ;
 wire \top_inst.sndgen_inst.slot_counter[3] ;
 wire \top_inst.sndgen_inst.slot_counter[4] ;
 wire \top_inst.sndgen_inst.slot_counter[5] ;
 wire \top_inst.sndgen_inst.slot_counter[6] ;
 wire \top_inst.sndgen_inst.slot_counter[7] ;
 wire \top_inst.sndgen_inst.slot_counter[8] ;
 wire \top_inst.sndgen_inst.slot_counter[9] ;
 wire \top_inst.sys_presc[0] ;
 wire \top_inst.sys_presc[1] ;
 wire \top_inst.sys_presc[2] ;
 wire \top_inst.sys_presc[3] ;
 wire \top_inst.sys_presc[4] ;
 wire \top_inst.vga_inst.bg[0] ;
 wire \top_inst.vga_inst.bg[1] ;
 wire \top_inst.vga_inst.bg[4] ;
 wire \top_inst.vga_inst.bg[5] ;
 wire \top_inst.vga_inst.sr1[0] ;
 wire \top_inst.vga_inst.sr1[1] ;
 wire \top_inst.vga_inst.sr1[2] ;
 wire \top_inst.vga_inst.sr1[3] ;
 wire \top_inst.vga_inst.sx1[0] ;
 wire \top_inst.vga_inst.sx1[1] ;
 wire \top_inst.vga_inst.sx1[2] ;
 wire \top_inst.vga_inst.sx1[3] ;
 wire \top_inst.vga_inst.vsync ;
 wire \top_inst.vga_inst.x1[0] ;
 wire \top_inst.vga_inst.x1[1] ;
 wire \top_inst.vga_inst.x1[2] ;
 wire \top_inst.vga_inst.x1[3] ;
 wire \top_inst.vga_inst.x1[4] ;
 wire \top_inst.vga_inst.x1[5] ;
 wire \top_inst.vga_inst.x1[6] ;
 wire \top_inst.vga_inst.x1[7] ;
 wire \top_inst.vga_inst.x[0] ;
 wire \top_inst.vga_inst.x[1] ;
 wire \top_inst.vga_inst.x[2] ;
 wire \top_inst.vga_inst.x[3] ;
 wire \top_inst.vga_inst.x[4] ;
 wire \top_inst.vga_inst.x[5] ;
 wire \top_inst.vga_inst.x[6] ;
 wire \top_inst.vga_inst.x[7] ;
 wire \top_inst.vga_inst.x[8] ;
 wire \top_inst.vga_inst.x[9] ;
 wire \top_inst.vga_inst.xmax[0] ;
 wire \top_inst.vga_inst.xmax[1] ;
 wire \top_inst.vga_inst.xmax[2] ;
 wire \top_inst.vga_inst.xmax[3] ;
 wire \top_inst.vga_inst.xmin[0] ;
 wire \top_inst.vga_inst.xmin[1] ;
 wire \top_inst.vga_inst.xmin[2] ;
 wire \top_inst.vga_inst.xmin[3] ;
 wire \top_inst.vga_inst.y[0] ;
 wire \top_inst.vga_inst.y[1] ;
 wire \top_inst.vga_inst.y[2] ;
 wire \top_inst.vga_inst.y[7] ;
 wire \top_inst.vga_inst.y[8] ;
 wire \top_inst.vga_inst.y[9] ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_0_clk;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net1;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;

 sg13g2_inv_1 _0896_ (.Y(_0236_),
    .A(net25));
 sg13g2_inv_1 _0897_ (.Y(_0237_),
    .A(net241));
 sg13g2_inv_1 _0898_ (.Y(_0238_),
    .A(\top_inst.vga_inst.y[0] ));
 sg13g2_inv_1 _0899_ (.Y(_0239_),
    .A(net183));
 sg13g2_inv_2 _0900_ (.Y(_0240_),
    .A(\top_inst.sndgen_inst.slot_counter[1] ));
 sg13g2_inv_1 _0901_ (.Y(_0241_),
    .A(net370));
 sg13g2_inv_1 _0902_ (.Y(_0242_),
    .A(net384));
 sg13g2_inv_1 _0903_ (.Y(_0243_),
    .A(\top_inst.vga_inst.sr1[3] ));
 sg13g2_inv_1 _0904_ (.Y(_0244_),
    .A(\top_inst.vga_inst.sx1[3] ));
 sg13g2_inv_1 _0905_ (.Y(_0245_),
    .A(\top_inst.vga_inst.sx1[2] ));
 sg13g2_inv_1 _0906_ (.Y(_0246_),
    .A(\top_inst.vga_inst.sr1[2] ));
 sg13g2_inv_1 _0907_ (.Y(_0247_),
    .A(\top_inst.vga_inst.x1[4] ));
 sg13g2_inv_1 _0908_ (.Y(_0248_),
    .A(\top_inst.vga_inst.x1[5] ));
 sg13g2_inv_1 _0909_ (.Y(_0249_),
    .A(\top_inst.vga_inst.x1[6] ));
 sg13g2_inv_1 _0910_ (.Y(_0250_),
    .A(net375));
 sg13g2_inv_1 _0911_ (.Y(_0251_),
    .A(\top_inst.sndgen_inst.rom_addr[3] ));
 sg13g2_inv_1 _0912_ (.Y(_0252_),
    .A(\top_inst.sndgen_inst.rom_addr[0] ));
 sg13g2_inv_1 _0913_ (.Y(_0253_),
    .A(net300));
 sg13g2_inv_1 _0914_ (.Y(_0254_),
    .A(net64));
 sg13g2_inv_1 _0915_ (.Y(_0255_),
    .A(\top_inst.sndgen_inst.c4[2] ));
 sg13g2_inv_1 _0916_ (.Y(_0256_),
    .A(_0008_));
 sg13g2_inv_1 _0917_ (.Y(_0257_),
    .A(\top_inst.sndgen_inst.phacc2[13] ));
 sg13g2_inv_1 _0918_ (.Y(_0258_),
    .A(\top_inst.pwm_inst.cntr[3] ));
 sg13g2_inv_1 _0919_ (.Y(_0259_),
    .A(net315));
 sg13g2_inv_1 _0920_ (.Y(_0260_),
    .A(net189));
 sg13g2_inv_1 _0921_ (.Y(_0261_),
    .A(net80));
 sg13g2_inv_1 _0922_ (.Y(_0262_),
    .A(net71));
 sg13g2_inv_1 _0923_ (.Y(_0263_),
    .A(net117));
 sg13g2_inv_1 _0924_ (.Y(_0264_),
    .A(net216));
 sg13g2_inv_1 _0925_ (.Y(_0265_),
    .A(\top_inst.vga_inst.xmax[0] ));
 sg13g2_inv_1 _0926_ (.Y(_0266_),
    .A(net177));
 sg13g2_inv_1 _0927_ (.Y(_0267_),
    .A(net165));
 sg13g2_inv_1 _0928_ (.Y(_0268_),
    .A(_0010_));
 sg13g2_inv_1 _0929_ (.Y(_0269_),
    .A(_0011_));
 sg13g2_inv_1 _0930_ (.Y(_0270_),
    .A(_0000_));
 sg13g2_nor4_2 _0931_ (.A(\top_inst.vga_inst.x[3] ),
    .B(\top_inst.vga_inst.x[2] ),
    .C(\top_inst.vga_inst.x[1] ),
    .Y(_0271_),
    .D(\top_inst.vga_inst.x[0] ));
 sg13g2_nor2_2 _0932_ (.A(\top_inst.vga_inst.x[4] ),
    .B(\top_inst.vga_inst.x[5] ),
    .Y(_0272_));
 sg13g2_and2_2 _0933_ (.A(_0271_),
    .B(_0272_),
    .X(_0273_));
 sg13g2_nand2_1 _0934_ (.Y(_0274_),
    .A(\top_inst.vga_inst.x[7] ),
    .B(\top_inst.vga_inst.x[9] ));
 sg13g2_nor2_2 _0935_ (.A(net258),
    .B(_0274_),
    .Y(_0275_));
 sg13g2_nor3_1 _0936_ (.A(_0237_),
    .B(\top_inst.vga_inst.x[6] ),
    .C(_0001_),
    .Y(_0276_));
 sg13g2_and3_1 _0937_ (.X(\top_inst.sample_ena ),
    .A(_0273_),
    .B(_0275_),
    .C(_0276_));
 sg13g2_and2_1 _0938_ (.A(\top_inst.vga_inst.x[7] ),
    .B(\top_inst.vga_inst.x[6] ),
    .X(_0277_));
 sg13g2_nand2_1 _0939_ (.Y(_0278_),
    .A(\top_inst.vga_inst.x[7] ),
    .B(\top_inst.vga_inst.x[6] ));
 sg13g2_nand2_1 _0940_ (.Y(_0279_),
    .A(\top_inst.vga_inst.x[5] ),
    .B(_0277_));
 sg13g2_nand3_1 _0941_ (.B(\top_inst.vga_inst.x[5] ),
    .C(_0277_),
    .A(net259),
    .Y(_0280_));
 sg13g2_nand2b_1 _0942_ (.Y(_0281_),
    .B(_0272_),
    .A_N(\top_inst.vga_inst.x[6] ));
 sg13g2_nand3_1 _0943_ (.B(_0280_),
    .C(_0281_),
    .A(_0275_),
    .Y(hsync));
 sg13g2_nand2_1 _0944_ (.Y(_0282_),
    .A(\top_inst.vga_inst.y[7] ),
    .B(\top_inst.vga_inst.bg[5] ));
 sg13g2_nor2_1 _0945_ (.A(_0002_),
    .B(_0282_),
    .Y(_0283_));
 sg13g2_a21oi_1 _0946_ (.A1(\top_inst.vga_inst.y[0] ),
    .A2(net394),
    .Y(_0284_),
    .B1(net365));
 sg13g2_nor3_1 _0947_ (.A(_0002_),
    .B(_0282_),
    .C(_0284_),
    .Y(_0285_));
 sg13g2_nand3_1 _0948_ (.B(\top_inst.vga_inst.bg[5] ),
    .C(\top_inst.vga_inst.y[8] ),
    .A(\top_inst.vga_inst.y[7] ),
    .Y(_0286_));
 sg13g2_inv_1 _0949_ (.Y(_0287_),
    .A(_0286_));
 sg13g2_nand2_1 _0950_ (.Y(_0288_),
    .A(_0242_),
    .B(_0287_));
 sg13g2_nor2b_1 _0951_ (.A(\top_inst.vga_inst.bg[1] ),
    .B_N(\top_inst.vga_inst.bg[4] ),
    .Y(_0289_));
 sg13g2_nand2_1 _0952_ (.Y(_0290_),
    .A(\top_inst.vga_inst.bg[0] ),
    .B(_0289_));
 sg13g2_nor4_1 _0953_ (.A(_0241_),
    .B(\top_inst.vga_inst.y[2] ),
    .C(_0288_),
    .D(_0290_),
    .Y(_0291_));
 sg13g2_o21ai_1 _0954_ (.B1(_0291_),
    .Y(\top_inst.vga_inst.vsync ),
    .A1(_0238_),
    .A2(_0285_));
 sg13g2_nor4_2 _0955_ (.A(\top_inst.vga_inst.y[0] ),
    .B(\top_inst.vga_inst.y[1] ),
    .C(\top_inst.vga_inst.bg[0] ),
    .Y(_0292_),
    .D(\top_inst.vga_inst.y[2] ));
 sg13g2_inv_1 _0956_ (.Y(_0293_),
    .A(_0292_));
 sg13g2_and2_1 _0957_ (.A(_0289_),
    .B(_0292_),
    .X(_0294_));
 sg13g2_a221oi_1 _0958_ (.B2(_0294_),
    .C1(\top_inst.vga_inst.y[9] ),
    .B1(_0287_),
    .A1(\top_inst.vga_inst.y[8] ),
    .Y(_0295_),
    .A2(_0283_));
 sg13g2_nor4_1 _0959_ (.A(\top_inst.vga_inst.y[7] ),
    .B(\top_inst.vga_inst.bg[5] ),
    .C(\top_inst.vga_inst.y[8] ),
    .D(\top_inst.vga_inst.y[9] ),
    .Y(_0296_));
 sg13g2_nand3b_1 _0960_ (.B(_0296_),
    .C(_0002_),
    .Y(_0297_),
    .A_N(_0294_));
 sg13g2_nor2_1 _0961_ (.A(_0272_),
    .B(_0278_),
    .Y(_0298_));
 sg13g2_nor3_2 _0962_ (.A(net257),
    .B(net258),
    .C(_0298_),
    .Y(_0299_));
 sg13g2_nand2_1 _0963_ (.Y(_0300_),
    .A(net258),
    .B(_0277_));
 sg13g2_nor2_1 _0964_ (.A(_0272_),
    .B(_0300_),
    .Y(_0301_));
 sg13g2_nor3_1 _0965_ (.A(net257),
    .B(_0299_),
    .C(_0301_),
    .Y(_0302_));
 sg13g2_nand3_1 _0966_ (.B(_0297_),
    .C(_0302_),
    .A(_0295_),
    .Y(_0303_));
 sg13g2_nor2_1 _0967_ (.A(\top_inst.vga_inst.bg[1] ),
    .B(\top_inst.vga_inst.bg[4] ),
    .Y(_0304_));
 sg13g2_a21oi_1 _0968_ (.A1(\top_inst.vga_inst.bg[1] ),
    .A2(_0293_),
    .Y(_0305_),
    .B1(\top_inst.vga_inst.bg[4] ));
 sg13g2_nor2_1 _0969_ (.A(net257),
    .B(\top_inst.vga_inst.y[9] ),
    .Y(_0306_));
 sg13g2_o21ai_1 _0970_ (.B1(_0306_),
    .Y(_0307_),
    .A1(\top_inst.vga_inst.x[8] ),
    .A2(_0277_));
 sg13g2_nor2_1 _0971_ (.A(_0273_),
    .B(_0278_),
    .Y(_0308_));
 sg13g2_a221oi_1 _0972_ (.B2(net258),
    .C1(_0307_),
    .B1(_0308_),
    .A1(_0296_),
    .Y(_0309_),
    .A2(_0304_));
 sg13g2_o21ai_1 _0973_ (.B1(_0309_),
    .Y(_0310_),
    .A1(_0286_),
    .A2(_0305_));
 sg13g2_nand2_1 _0974_ (.Y(_0311_),
    .A(net257),
    .B(net258));
 sg13g2_o21ai_1 _0975_ (.B1(net257),
    .Y(_0312_),
    .A1(\top_inst.vga_inst.x[7] ),
    .A2(net258));
 sg13g2_nand4_1 _0976_ (.B(_0303_),
    .C(_0310_),
    .A(_0295_),
    .Y(_0313_),
    .D(_0312_));
 sg13g2_inv_1 _0977_ (.Y(_0314_),
    .A(_0313_));
 sg13g2_nor2b_1 _0978_ (.A(_0303_),
    .B_N(_0310_),
    .Y(_0315_));
 sg13g2_a22oi_1 _0979_ (.Y(_0316_),
    .B1(_0315_),
    .B2(\top_inst.vga_inst.bg[1] ),
    .A2(_0314_),
    .A1(\top_inst.vga_inst.bg[0] ));
 sg13g2_inv_1 _0980_ (.Y(uo_out[6]),
    .A(_0316_));
 sg13g2_nor2_1 _0981_ (.A(_0003_),
    .B(_0313_),
    .Y(uo_out[2]));
 sg13g2_nand2b_1 _0982_ (.Y(_0317_),
    .B(_0315_),
    .A_N(_0004_));
 sg13g2_o21ai_1 _0983_ (.B1(_0317_),
    .Y(uo_out[4]),
    .A1(_0002_),
    .A2(_0313_));
 sg13g2_nor2_1 _0984_ (.A(_0004_),
    .B(_0313_),
    .Y(uo_out[0]));
 sg13g2_or2_1 _0985_ (.X(_0318_),
    .B(\top_inst.sndgen_inst.mask_2 ),
    .A(\top_inst.sndgen_inst.mask_1[0] ));
 sg13g2_o21ai_1 _0986_ (.B1(_0318_),
    .Y(_0319_),
    .A1(\top_inst.sndgen_inst.c1[1] ),
    .A2(\top_inst.sndgen_inst.c1[0] ));
 sg13g2_and2_2 _0987_ (.A(\top_inst.sndgen_inst.slot_counter[10] ),
    .B(\top_inst.sndgen_inst.slot_counter[9] ),
    .X(_0320_));
 sg13g2_nor3_1 _0988_ (.A(\top_inst.sndgen_inst.slot_counter[5] ),
    .B(\top_inst.sndgen_inst.slot_counter[8] ),
    .C(\top_inst.sndgen_inst.slot_counter[7] ),
    .Y(_0321_));
 sg13g2_nor2_1 _0989_ (.A(\top_inst.sndgen_inst.slot_counter[0] ),
    .B(\top_inst.sndgen_inst.slot_counter[2] ),
    .Y(_0322_));
 sg13g2_nor4_1 _0990_ (.A(\top_inst.sndgen_inst.slot_counter[1] ),
    .B(\top_inst.sndgen_inst.slot_counter[4] ),
    .C(\top_inst.sndgen_inst.slot_counter[3] ),
    .D(\top_inst.sndgen_inst.slot_counter[6] ),
    .Y(_0323_));
 sg13g2_nand3_1 _0991_ (.B(_0322_),
    .C(_0323_),
    .A(_0321_),
    .Y(_0324_));
 sg13g2_nand2b_1 _0992_ (.Y(_0325_),
    .B(\top_inst.sndgen_inst.c1[0] ),
    .A_N(\top_inst.sndgen_inst.c1[1] ));
 sg13g2_a221oi_1 _0993_ (.B2(\top_inst.sndgen_inst.lfsr[7] ),
    .C1(_0319_),
    .B1(_0325_),
    .A1(_0320_),
    .Y(_0326_),
    .A2(_0324_));
 sg13g2_a21oi_2 _0994_ (.B1(_0008_),
    .Y(_0327_),
    .A2(_0324_),
    .A1(_0320_));
 sg13g2_a21oi_1 _0995_ (.A1(_0257_),
    .A2(_0327_),
    .Y(_0328_),
    .B1(_0326_));
 sg13g2_a21o_1 _0996_ (.A2(_0327_),
    .A1(_0257_),
    .B1(_0326_),
    .X(_0329_));
 sg13g2_nand2b_1 _0997_ (.Y(_0330_),
    .B(\top_inst.sndgen_inst.mask_1[2] ),
    .A_N(\top_inst.sndgen_inst.phacc3[13] ));
 sg13g2_nand3_1 _0998_ (.B(_0326_),
    .C(_0327_),
    .A(_0257_),
    .Y(_0331_));
 sg13g2_and3_1 _0999_ (.X(_0332_),
    .A(_0329_),
    .B(_0330_),
    .C(_0331_));
 sg13g2_nor2_1 _1000_ (.A(_0328_),
    .B(_0332_),
    .Y(_0333_));
 sg13g2_nand2_1 _1001_ (.Y(_0334_),
    .A(\top_inst.sndgen_inst.lfsr[5] ),
    .B(_0325_));
 sg13g2_nand3b_1 _1002_ (.B(\top_inst.sndgen_inst.c1[0] ),
    .C(\top_inst.sndgen_inst.lfsr[7] ),
    .Y(_0335_),
    .A_N(\top_inst.sndgen_inst.c1[1] ));
 sg13g2_a221oi_1 _1003_ (.B2(_0335_),
    .C1(_0319_),
    .B1(_0334_),
    .A1(_0320_),
    .Y(_0336_),
    .A2(_0324_));
 sg13g2_mux2_1 _1004_ (.A0(_0327_),
    .A1(_0008_),
    .S(_0336_),
    .X(_0337_));
 sg13g2_a22oi_1 _1005_ (.Y(_0338_),
    .B1(_0337_),
    .B2(\top_inst.sndgen_inst.mask_1[2] ),
    .A2(_0336_),
    .A1(_0256_));
 sg13g2_a21oi_1 _1006_ (.A1(_0329_),
    .A2(_0331_),
    .Y(_0339_),
    .B1(_0330_));
 sg13g2_nor3_1 _1007_ (.A(_0332_),
    .B(_0338_),
    .C(_0339_),
    .Y(_0340_));
 sg13g2_or3_1 _1008_ (.A(_0332_),
    .B(_0338_),
    .C(_0339_),
    .X(_0341_));
 sg13g2_nand2b_1 _1009_ (.Y(_0342_),
    .B(\top_inst.sndgen_inst.mask_1[3] ),
    .A_N(\top_inst.sndgen_inst.phacc4[13] ));
 sg13g2_o21ai_1 _1010_ (.B1(_0338_),
    .Y(_0343_),
    .A1(_0332_),
    .A2(_0339_));
 sg13g2_nand3_1 _1011_ (.B(_0342_),
    .C(_0343_),
    .A(_0341_),
    .Y(_0344_));
 sg13g2_a21oi_1 _1012_ (.A1(_0342_),
    .A2(_0343_),
    .Y(_0345_),
    .B1(_0340_));
 sg13g2_nor2_1 _1013_ (.A(_0333_),
    .B(_0345_),
    .Y(_0346_));
 sg13g2_xnor2_1 _1014_ (.Y(_0347_),
    .A(\top_inst.sndgen_inst.mask_1[2] ),
    .B(_0337_));
 sg13g2_nor2_1 _1015_ (.A(_0009_),
    .B(_0347_),
    .Y(_0348_));
 sg13g2_a21o_1 _1016_ (.A2(_0343_),
    .A1(_0341_),
    .B1(_0342_),
    .X(_0349_));
 sg13g2_nand3_1 _1017_ (.B(_0348_),
    .C(_0349_),
    .A(_0344_),
    .Y(_0350_));
 sg13g2_xnor2_1 _1018_ (.Y(_0351_),
    .A(_0333_),
    .B(_0345_));
 sg13g2_nor2_1 _1019_ (.A(_0350_),
    .B(_0351_),
    .Y(_0352_));
 sg13g2_nor2_1 _1020_ (.A(_0346_),
    .B(_0352_),
    .Y(_0353_));
 sg13g2_or2_1 _1021_ (.X(_0354_),
    .B(_0352_),
    .A(_0346_));
 sg13g2_xnor2_1 _1022_ (.Y(_0355_),
    .A(_0350_),
    .B(_0351_));
 sg13g2_nand2_1 _1023_ (.Y(_0356_),
    .A(\top_inst.pwm_inst.cntr[2] ),
    .B(_0355_));
 sg13g2_xor2_1 _1024_ (.B(_0347_),
    .A(net123),
    .X(_0357_));
 sg13g2_o21ai_1 _1025_ (.B1(_0357_),
    .Y(_0358_),
    .A1(\top_inst.pwm_inst.cntr[0] ),
    .A2(_0017_));
 sg13g2_o21ai_1 _1026_ (.B1(_0358_),
    .Y(_0359_),
    .A1(_0017_),
    .A2(_0357_));
 sg13g2_a21o_1 _1027_ (.A2(_0349_),
    .A1(_0344_),
    .B1(_0348_),
    .X(_0360_));
 sg13g2_nand2_1 _1028_ (.Y(_0361_),
    .A(_0350_),
    .B(_0360_));
 sg13g2_nor2_1 _1029_ (.A(\top_inst.pwm_inst.cntr[1] ),
    .B(_0359_),
    .Y(_0362_));
 sg13g2_a21oi_1 _1030_ (.A1(\top_inst.pwm_inst.cntr[1] ),
    .A2(_0359_),
    .Y(_0363_),
    .B1(_0361_));
 sg13g2_o21ai_1 _1031_ (.B1(_0356_),
    .Y(_0364_),
    .A1(_0362_),
    .A2(_0363_));
 sg13g2_nor2_1 _1032_ (.A(\top_inst.pwm_inst.cntr[2] ),
    .B(_0355_),
    .Y(_0365_));
 sg13g2_a21oi_1 _1033_ (.A1(_0258_),
    .A2(_0354_),
    .Y(_0366_),
    .B1(_0365_));
 sg13g2_a22oi_1 _1034_ (.Y(pwm),
    .B1(_0364_),
    .B2(_0366_),
    .A2(_0353_),
    .A1(\top_inst.pwm_inst.cntr[3] ));
 sg13g2_nand2b_1 _1035_ (.Y(_0367_),
    .B(net259),
    .A_N(\top_inst.vga_inst.x[5] ));
 sg13g2_or3_1 _1036_ (.A(net257),
    .B(net258),
    .C(_0271_),
    .X(_0368_));
 sg13g2_nor3_1 _1037_ (.A(_0278_),
    .B(_0367_),
    .C(_0368_),
    .Y(_0369_));
 sg13g2_nor4_1 _1038_ (.A(net259),
    .B(\top_inst.vga_inst.x[5] ),
    .C(_0278_),
    .D(_0368_),
    .Y(_0370_));
 sg13g2_nand2_1 _1039_ (.Y(_0371_),
    .A(_0247_),
    .B(\top_inst.vga_inst.xmax[0] ));
 sg13g2_o21ai_1 _1040_ (.B1(_0371_),
    .Y(_0372_),
    .A1(\top_inst.vga_inst.x1[2] ),
    .A2(\top_inst.vga_inst.x1[3] ));
 sg13g2_a22oi_1 _1041_ (.Y(_0373_),
    .B1(_0265_),
    .B2(\top_inst.vga_inst.x1[4] ),
    .A2(_0264_),
    .A1(\top_inst.vga_inst.x1[5] ));
 sg13g2_a22oi_1 _1042_ (.Y(_0374_),
    .B1(_0372_),
    .B2(_0373_),
    .A2(\top_inst.vga_inst.xmax[1] ),
    .A1(_0248_));
 sg13g2_nor2_1 _1043_ (.A(_0249_),
    .B(\top_inst.vga_inst.xmax[2] ),
    .Y(_0375_));
 sg13g2_a22oi_1 _1044_ (.Y(_0376_),
    .B1(\top_inst.vga_inst.xmax[2] ),
    .B2(_0249_),
    .A2(\top_inst.vga_inst.xmax[3] ),
    .A1(_0250_));
 sg13g2_o21ai_1 _1045_ (.B1(_0376_),
    .Y(_0377_),
    .A1(_0374_),
    .A2(_0375_));
 sg13g2_nand2_1 _1046_ (.Y(_0378_),
    .A(_0250_),
    .B(\top_inst.vga_inst.xmin[3] ));
 sg13g2_nand2_1 _1047_ (.Y(_0379_),
    .A(\top_inst.vga_inst.x1[7] ),
    .B(_0262_));
 sg13g2_a22oi_1 _1048_ (.Y(_0380_),
    .B1(\top_inst.vga_inst.xmin[1] ),
    .B2(_0248_),
    .A2(\top_inst.vga_inst.xmin[0] ),
    .A1(_0247_));
 sg13g2_a221oi_1 _1049_ (.B2(\top_inst.vga_inst.x1[6] ),
    .C1(_0380_),
    .B1(_0261_),
    .A1(\top_inst.vga_inst.x1[5] ),
    .Y(_0381_),
    .A2(_0259_));
 sg13g2_a21oi_1 _1050_ (.A1(_0249_),
    .A2(\top_inst.vga_inst.xmin[2] ),
    .Y(_0382_),
    .B1(_0381_));
 sg13g2_a21o_1 _1051_ (.A2(_0260_),
    .A1(\top_inst.vga_inst.x1[7] ),
    .B1(_0382_),
    .X(_0383_));
 sg13g2_nand4_1 _1052_ (.B(_0378_),
    .C(_0379_),
    .A(_0377_),
    .Y(_0384_),
    .D(_0383_));
 sg13g2_nor2_1 _1053_ (.A(_0271_),
    .B(_0292_),
    .Y(_0385_));
 sg13g2_inv_1 _1054_ (.Y(_0386_),
    .A(_0385_));
 sg13g2_and2_1 _1055_ (.A(_0384_),
    .B(_0385_),
    .X(_0387_));
 sg13g2_mux2_1 _1056_ (.A0(_0387_),
    .A1(_0319_),
    .S(_0370_),
    .X(_0388_));
 sg13g2_nor3_1 _1057_ (.A(net259),
    .B(_0279_),
    .C(_0368_),
    .Y(_0389_));
 sg13g2_nor3_1 _1058_ (.A(\top_inst.sndgen_inst.c2[0] ),
    .B(\top_inst.sndgen_inst.c2[1] ),
    .C(\top_inst.sndgen_inst.c2[2] ),
    .Y(_0390_));
 sg13g2_nor2_1 _1059_ (.A(_0008_),
    .B(_0390_),
    .Y(_0391_));
 sg13g2_a21oi_1 _1060_ (.A1(_0369_),
    .A2(_0391_),
    .Y(_0392_),
    .B1(_0389_));
 sg13g2_o21ai_1 _1061_ (.B1(_0392_),
    .Y(_0393_),
    .A1(_0369_),
    .A2(_0388_));
 sg13g2_nor2_1 _1062_ (.A(_0271_),
    .B(_0280_),
    .Y(_0394_));
 sg13g2_nor3_2 _1063_ (.A(\top_inst.sndgen_inst.c3[0] ),
    .B(\top_inst.sndgen_inst.c3[1] ),
    .C(\top_inst.sndgen_inst.c3[2] ),
    .Y(_0395_));
 sg13g2_nand2b_1 _1064_ (.Y(_0396_),
    .B(\top_inst.sndgen_inst.mask_1[2] ),
    .A_N(_0395_));
 sg13g2_a21oi_1 _1065_ (.A1(_0389_),
    .A2(_0396_),
    .Y(_0397_),
    .B1(_0394_));
 sg13g2_nand2_1 _1066_ (.Y(_0398_),
    .A(_0393_),
    .B(_0397_));
 sg13g2_or2_1 _1067_ (.X(_0399_),
    .B(_0305_),
    .A(_0297_));
 sg13g2_a21oi_1 _1068_ (.A1(_0255_),
    .A2(_0395_),
    .Y(_0400_),
    .B1(_0009_));
 sg13g2_a21oi_1 _1069_ (.A1(_0394_),
    .A2(_0400_),
    .Y(_0401_),
    .B1(_0399_));
 sg13g2_a221oi_1 _1070_ (.B2(_0398_),
    .C1(_0310_),
    .B1(_0401_),
    .A1(_0387_),
    .Y(uo_out[1]),
    .A2(_0399_));
 sg13g2_a21oi_2 _1071_ (.B1(_0310_),
    .Y(uo_out[5]),
    .A2(_0386_),
    .A1(_0384_));
 sg13g2_or2_1 _1072_ (.X(_0402_),
    .B(\top_inst.sys_presc[1] ),
    .A(net240));
 sg13g2_xor2_1 _1073_ (.B(net122),
    .A(net240),
    .X(_0012_));
 sg13g2_nand3_1 _1074_ (.B(net122),
    .C(net381),
    .A(net240),
    .Y(_0403_));
 sg13g2_a21o_1 _1075_ (.A2(net122),
    .A1(net240),
    .B1(net381),
    .X(_0404_));
 sg13g2_and2_1 _1076_ (.A(_0403_),
    .B(_0404_),
    .X(_0013_));
 sg13g2_nand4_1 _1077_ (.B(\top_inst.sys_presc[1] ),
    .C(\top_inst.sys_presc[3] ),
    .A(net240),
    .Y(_0405_),
    .D(\top_inst.sys_presc[2] ));
 sg13g2_xnor2_1 _1078_ (.Y(_0014_),
    .A(net119),
    .B(_0403_));
 sg13g2_xnor2_1 _1079_ (.Y(_0015_),
    .A(net49),
    .B(_0405_));
 sg13g2_nand4_1 _1080_ (.B(\top_inst.sndgen_inst.rom_addr[1] ),
    .C(\top_inst.sndgen_inst.rom_addr[0] ),
    .A(\top_inst.sndgen_inst.rom_addr[3] ),
    .Y(_0406_),
    .D(_0006_));
 sg13g2_nor2b_2 _1081_ (.A(net152),
    .B_N(\top_inst.sndgen_inst.rom_addr[2] ),
    .Y(_0407_));
 sg13g2_nand2_1 _1082_ (.Y(_0408_),
    .A(_0252_),
    .B(_0407_));
 sg13g2_and2_1 _1083_ (.A(_0406_),
    .B(_0408_),
    .X(_0409_));
 sg13g2_nor2_1 _1084_ (.A(net180),
    .B(net245),
    .Y(_0410_));
 sg13g2_a21oi_1 _1085_ (.A1(net245),
    .A2(_0409_),
    .Y(_0021_),
    .B1(net181));
 sg13g2_nor2_2 _1086_ (.A(net386),
    .B(_0252_),
    .Y(_0411_));
 sg13g2_nand2_1 _1087_ (.Y(_0412_),
    .A(_0251_),
    .B(\top_inst.sndgen_inst.rom_addr[1] ));
 sg13g2_and2_1 _1088_ (.A(_0411_),
    .B(_0412_),
    .X(_0413_));
 sg13g2_o21ai_1 _1089_ (.B1(_0407_),
    .Y(_0414_),
    .A1(\top_inst.sndgen_inst.rom_addr[1] ),
    .A2(_0252_));
 sg13g2_nor2b_1 _1090_ (.A(_0413_),
    .B_N(_0414_),
    .Y(_0415_));
 sg13g2_nor2_1 _1091_ (.A(net147),
    .B(\top_inst.sndgen_inst.sample_ena_delay[2] ),
    .Y(_0416_));
 sg13g2_a21oi_1 _1092_ (.A1(net245),
    .A2(_0415_),
    .Y(_0022_),
    .B1(net148));
 sg13g2_nand2_1 _1093_ (.Y(_0417_),
    .A(_0251_),
    .B(\top_inst.sndgen_inst.rom_addr[0] ));
 sg13g2_o21ai_1 _1094_ (.B1(_0406_),
    .Y(_0418_),
    .A1(\top_inst.sndgen_inst.rom_addr[2] ),
    .A2(_0417_));
 sg13g2_a21oi_2 _1095_ (.B1(_0418_),
    .Y(_0419_),
    .A2(_0407_),
    .A1(\top_inst.sndgen_inst.rom_addr[1] ));
 sg13g2_nor2_1 _1096_ (.A(net186),
    .B(\top_inst.sndgen_inst.sample_ena_delay[2] ),
    .Y(_0420_));
 sg13g2_a21oi_1 _1097_ (.A1(net245),
    .A2(_0419_),
    .Y(_0023_),
    .B1(net187));
 sg13g2_nor2b_2 _1098_ (.A(\top_inst.sndgen_inst.rom_addr[1] ),
    .B_N(_0407_),
    .Y(_0421_));
 sg13g2_nor2_2 _1099_ (.A(_0418_),
    .B(_0421_),
    .Y(_0422_));
 sg13g2_nor2_1 _1100_ (.A(net158),
    .B(net245),
    .Y(_0423_));
 sg13g2_a21oi_1 _1101_ (.A1(net245),
    .A2(_0422_),
    .Y(_0024_),
    .B1(net159));
 sg13g2_a21oi_2 _1102_ (.B1(_0411_),
    .Y(_0424_),
    .A2(net343),
    .A1(net336));
 sg13g2_nor2_1 _1103_ (.A(net261),
    .B(net245),
    .Y(_0425_));
 sg13g2_a21oi_1 _1104_ (.A1(net245),
    .A2(net344),
    .Y(_0025_),
    .B1(net350));
 sg13g2_nand2_1 _1105_ (.Y(_0426_),
    .A(net108),
    .B(\top_inst.sndgen_inst.slot_counter[3] ));
 sg13g2_nand3_1 _1106_ (.B(\top_inst.sndgen_inst.slot_counter[5] ),
    .C(\top_inst.sndgen_inst.slot_counter[8] ),
    .A(\top_inst.sndgen_inst.slot_counter[2] ),
    .Y(_0427_));
 sg13g2_nand2_1 _1107_ (.Y(_0428_),
    .A(\top_inst.sndgen_inst.slot_counter[6] ),
    .B(\top_inst.sndgen_inst.slot_counter[7] ));
 sg13g2_nor3_1 _1108_ (.A(_0426_),
    .B(_0427_),
    .C(_0428_),
    .Y(_0429_));
 sg13g2_and2_1 _1109_ (.A(_0320_),
    .B(_0429_),
    .X(_0430_));
 sg13g2_nor2_1 _1110_ (.A(\top_inst.vga_inst.x[6] ),
    .B(net66),
    .Y(_0431_));
 sg13g2_and4_2 _1111_ (.A(net241),
    .B(_0273_),
    .C(_0275_),
    .D(_0431_),
    .X(_0432_));
 sg13g2_nand4_1 _1112_ (.B(_0273_),
    .C(_0275_),
    .A(net242),
    .Y(_0433_),
    .D(_0431_));
 sg13g2_nor3_2 _1113_ (.A(_0016_),
    .B(_0240_),
    .C(_0433_),
    .Y(_0434_));
 sg13g2_and3_1 _1114_ (.X(_0435_),
    .A(_0273_),
    .B(_0275_),
    .C(_0276_));
 sg13g2_nand3_1 _1115_ (.B(_0275_),
    .C(_0276_),
    .A(_0273_),
    .Y(_0436_));
 sg13g2_nor3_2 _1116_ (.A(_0016_),
    .B(_0240_),
    .C(net229),
    .Y(_0437_));
 sg13g2_nand2_1 _1117_ (.Y(_0438_),
    .A(_0430_),
    .B(net226));
 sg13g2_nand2_1 _1118_ (.Y(_0439_),
    .A(net387),
    .B(\top_inst.sndgen_inst.bar_counter[0] ));
 sg13g2_o21ai_1 _1119_ (.B1(_0439_),
    .Y(_0440_),
    .A1(net304),
    .A2(\top_inst.sndgen_inst.bar_counter[2] ));
 sg13g2_nor2_1 _1120_ (.A(net304),
    .B(\top_inst.sndgen_inst.bar_counter[0] ),
    .Y(_0441_));
 sg13g2_nor3_1 _1121_ (.A(net221),
    .B(_0440_),
    .C(_0441_),
    .Y(_0442_));
 sg13g2_a21o_1 _1122_ (.A2(net221),
    .A1(net332),
    .B1(_0442_),
    .X(_0026_));
 sg13g2_nand2_1 _1123_ (.Y(_0443_),
    .A(net21),
    .B(net221));
 sg13g2_o21ai_1 _1124_ (.B1(_0443_),
    .Y(_0027_),
    .A1(net221),
    .A2(_0441_));
 sg13g2_nor4_2 _1125_ (.A(net341),
    .B(\top_inst.vga_inst.x[6] ),
    .C(_0311_),
    .Y(_0444_),
    .D(_0367_));
 sg13g2_nand3_1 _1126_ (.B(net380),
    .C(net337),
    .A(net240),
    .Y(_0445_));
 sg13g2_nand4_1 _1127_ (.B(\top_inst.vga_inst.x[2] ),
    .C(\top_inst.vga_inst.x[1] ),
    .A(net240),
    .Y(_0446_),
    .D(\top_inst.vga_inst.x[0] ));
 sg13g2_and4_1 _1128_ (.A(\top_inst.vga_inst.x[3] ),
    .B(\top_inst.vga_inst.x[2] ),
    .C(\top_inst.vga_inst.x[1] ),
    .D(\top_inst.vga_inst.x[0] ),
    .X(_0447_));
 sg13g2_and2_2 _1129_ (.A(net241),
    .B(_0447_),
    .X(_0448_));
 sg13g2_and2_2 _1130_ (.A(_0444_),
    .B(_0448_),
    .X(_0449_));
 sg13g2_nand2_2 _1131_ (.Y(_0450_),
    .A(_0444_),
    .B(_0448_));
 sg13g2_nor4_1 _1132_ (.A(\top_inst.vga_inst.y[0] ),
    .B(\top_inst.vga_inst.y[1] ),
    .C(\top_inst.vga_inst.y[8] ),
    .D(_0242_),
    .Y(_0451_));
 sg13g2_nor4_1 _1133_ (.A(\top_inst.vga_inst.y[7] ),
    .B(\top_inst.vga_inst.bg[5] ),
    .C(\top_inst.vga_inst.bg[1] ),
    .D(\top_inst.vga_inst.bg[4] ),
    .Y(_0452_));
 sg13g2_nand4_1 _1134_ (.B(\top_inst.vga_inst.y[2] ),
    .C(_0451_),
    .A(\top_inst.vga_inst.bg[0] ),
    .Y(_0453_),
    .D(_0452_));
 sg13g2_nand2_1 _1135_ (.Y(_0454_),
    .A(_0449_),
    .B(_0453_));
 sg13g2_nand3_1 _1136_ (.B(_0449_),
    .C(_0453_),
    .A(net66),
    .Y(_0455_));
 sg13g2_o21ai_1 _1137_ (.B1(_0455_),
    .Y(_0028_),
    .A1(_0238_),
    .A2(_0449_));
 sg13g2_xor2_1 _1138_ (.B(net370),
    .A(\top_inst.vga_inst.y[0] ),
    .X(_0456_));
 sg13g2_nor2_1 _1139_ (.A(_0450_),
    .B(_0456_),
    .Y(_0457_));
 sg13g2_a21oi_1 _1140_ (.A1(_0241_),
    .A2(_0450_),
    .Y(_0029_),
    .B1(_0457_));
 sg13g2_and3_1 _1141_ (.X(_0458_),
    .A(\top_inst.vga_inst.y[0] ),
    .B(\top_inst.vga_inst.y[1] ),
    .C(\top_inst.vga_inst.y[2] ));
 sg13g2_nor3_1 _1142_ (.A(_0284_),
    .B(_0454_),
    .C(_0458_),
    .Y(_0459_));
 sg13g2_a21o_1 _1143_ (.A2(_0450_),
    .A1(net365),
    .B1(_0459_),
    .X(_0030_));
 sg13g2_and4_1 _1144_ (.A(net241),
    .B(_0444_),
    .C(_0447_),
    .D(_0458_),
    .X(_0460_));
 sg13g2_nor2_1 _1145_ (.A(net372),
    .B(_0460_),
    .Y(_0461_));
 sg13g2_nand3_1 _1146_ (.B(_0449_),
    .C(_0458_),
    .A(\top_inst.vga_inst.bg[0] ),
    .Y(_0462_));
 sg13g2_inv_1 _1147_ (.Y(_0463_),
    .A(_0462_));
 sg13g2_nor2_1 _1148_ (.A(_0450_),
    .B(_0453_),
    .Y(_0464_));
 sg13g2_nor3_1 _1149_ (.A(_0461_),
    .B(_0463_),
    .C(_0464_),
    .Y(_0031_));
 sg13g2_xnor2_1 _1150_ (.Y(_0032_),
    .A(net366),
    .B(_0462_));
 sg13g2_nor2_1 _1151_ (.A(net323),
    .B(_0462_),
    .Y(_0465_));
 sg13g2_xor2_1 _1152_ (.B(_0465_),
    .A(\top_inst.vga_inst.bg[4] ),
    .X(_0033_));
 sg13g2_and4_1 _1153_ (.A(\top_inst.vga_inst.bg[0] ),
    .B(\top_inst.vga_inst.bg[1] ),
    .C(\top_inst.vga_inst.bg[4] ),
    .D(_0460_),
    .X(_0466_));
 sg13g2_xor2_1 _1154_ (.B(_0466_),
    .A(net360),
    .X(_0034_));
 sg13g2_a21oi_1 _1155_ (.A1(\top_inst.vga_inst.bg[5] ),
    .A2(_0466_),
    .Y(_0467_),
    .B1(net327));
 sg13g2_and3_1 _1156_ (.X(_0468_),
    .A(net327),
    .B(\top_inst.vga_inst.bg[5] ),
    .C(_0466_));
 sg13g2_nor2_1 _1157_ (.A(net328),
    .B(_0468_),
    .Y(_0035_));
 sg13g2_nand2_1 _1158_ (.Y(_0469_),
    .A(net355),
    .B(_0468_));
 sg13g2_xor2_1 _1159_ (.B(_0468_),
    .A(net355),
    .X(_0036_));
 sg13g2_xnor2_1 _1160_ (.Y(_0470_),
    .A(_0242_),
    .B(_0469_));
 sg13g2_nor2_1 _1161_ (.A(_0464_),
    .B(_0470_),
    .Y(_0037_));
 sg13g2_xor2_1 _1162_ (.B(net337),
    .A(net241),
    .X(_0038_));
 sg13g2_a21o_1 _1163_ (.A2(net337),
    .A1(net240),
    .B1(net380),
    .X(_0471_));
 sg13g2_and2_1 _1164_ (.A(_0445_),
    .B(_0471_),
    .X(_0039_));
 sg13g2_xnor2_1 _1165_ (.Y(_0040_),
    .A(net191),
    .B(_0445_));
 sg13g2_xnor2_1 _1166_ (.Y(_0041_),
    .A(net78),
    .B(_0446_));
 sg13g2_xor2_1 _1167_ (.B(_0448_),
    .A(net259),
    .X(_0042_));
 sg13g2_a21oi_1 _1168_ (.A1(net259),
    .A2(_0448_),
    .Y(_0472_),
    .B1(net368));
 sg13g2_and3_1 _1169_ (.X(_0473_),
    .A(net259),
    .B(net368),
    .C(_0448_));
 sg13g2_nand3_1 _1170_ (.B(net368),
    .C(_0448_),
    .A(net259),
    .Y(_0474_));
 sg13g2_nor3_1 _1171_ (.A(_0449_),
    .B(net369),
    .C(_0473_),
    .Y(_0043_));
 sg13g2_xnor2_1 _1172_ (.Y(_0044_),
    .A(net373),
    .B(_0474_));
 sg13g2_a21oi_1 _1173_ (.A1(\top_inst.vga_inst.x[6] ),
    .A2(_0473_),
    .Y(_0475_),
    .B1(net341));
 sg13g2_nor2b_1 _1174_ (.A(_0280_),
    .B_N(_0448_),
    .Y(_0476_));
 sg13g2_nor2_1 _1175_ (.A(net342),
    .B(_0476_),
    .Y(_0045_));
 sg13g2_nor2_1 _1176_ (.A(net258),
    .B(_0476_),
    .Y(_0477_));
 sg13g2_nor2_1 _1177_ (.A(_0300_),
    .B(_0474_),
    .Y(_0478_));
 sg13g2_o21ai_1 _1178_ (.B1(_0450_),
    .Y(_0479_),
    .A1(_0300_),
    .A2(_0474_));
 sg13g2_nor2_1 _1179_ (.A(_0477_),
    .B(_0479_),
    .Y(_0046_));
 sg13g2_nor2_1 _1180_ (.A(net257),
    .B(_0478_),
    .Y(_0480_));
 sg13g2_a21oi_1 _1181_ (.A1(net257),
    .A2(_0479_),
    .Y(_0047_),
    .B1(_0480_));
 sg13g2_and2_1 _1182_ (.A(net242),
    .B(_0299_),
    .X(_0481_));
 sg13g2_nand2_1 _1183_ (.Y(_0482_),
    .A(net242),
    .B(_0299_));
 sg13g2_nand2b_1 _1184_ (.Y(_0483_),
    .B(\top_inst.vga_inst.sx1[1] ),
    .A_N(\top_inst.vga_inst.sr1[1] ));
 sg13g2_nand2b_1 _1185_ (.Y(_0484_),
    .B(\top_inst.vga_inst.sr1[1] ),
    .A_N(\top_inst.vga_inst.sx1[1] ));
 sg13g2_nand3b_1 _1186_ (.B(\top_inst.vga_inst.sx1[0] ),
    .C(_0484_),
    .Y(_0485_),
    .A_N(\top_inst.vga_inst.sr1[0] ));
 sg13g2_a22oi_1 _1187_ (.Y(_0486_),
    .B1(_0483_),
    .B2(_0485_),
    .A2(\top_inst.vga_inst.sr1[2] ),
    .A1(_0245_));
 sg13g2_a221oi_1 _1188_ (.B2(_0246_),
    .C1(_0486_),
    .B1(\top_inst.vga_inst.sx1[2] ),
    .A1(_0243_),
    .Y(_0487_),
    .A2(\top_inst.vga_inst.sx1[3] ));
 sg13g2_a21oi_1 _1189_ (.A1(\top_inst.vga_inst.sr1[3] ),
    .A2(_0244_),
    .Y(_0488_),
    .B1(_0487_));
 sg13g2_nand2_1 _1190_ (.Y(_0489_),
    .A(net32),
    .B(net222));
 sg13g2_nor2b_1 _1191_ (.A(\top_inst.vga_inst.sr1[0] ),
    .B_N(net220),
    .Y(_0490_));
 sg13g2_o21ai_1 _1192_ (.B1(net224),
    .Y(_0491_),
    .A1(\top_inst.vga_inst.sx1[0] ),
    .A2(net220));
 sg13g2_o21ai_1 _1193_ (.B1(_0489_),
    .Y(_0048_),
    .A1(_0490_),
    .A2(_0491_));
 sg13g2_nand2b_1 _1194_ (.Y(_0492_),
    .B(\top_inst.vga_inst.sx1[1] ),
    .A_N(net219));
 sg13g2_a21oi_1 _1195_ (.A1(\top_inst.vga_inst.sr1[1] ),
    .A2(net219),
    .Y(_0493_),
    .B1(net222));
 sg13g2_a22oi_1 _1196_ (.Y(_0049_),
    .B1(_0492_),
    .B2(_0493_),
    .A2(net222),
    .A1(_0259_));
 sg13g2_a21oi_1 _1197_ (.A1(_0246_),
    .A2(net219),
    .Y(_0494_),
    .B1(net223));
 sg13g2_o21ai_1 _1198_ (.B1(_0494_),
    .Y(_0495_),
    .A1(\top_inst.vga_inst.sx1[2] ),
    .A2(net219));
 sg13g2_o21ai_1 _1199_ (.B1(_0495_),
    .Y(_0050_),
    .A1(_0261_),
    .A2(net224));
 sg13g2_nand3_1 _1200_ (.B(\top_inst.vga_inst.sx1[3] ),
    .C(net224),
    .A(\top_inst.vga_inst.sr1[3] ),
    .Y(_0496_));
 sg13g2_o21ai_1 _1201_ (.B1(_0496_),
    .Y(_0051_),
    .A1(_0260_),
    .A2(net224));
 sg13g2_mux2_1 _1202_ (.A0(net30),
    .A1(_0007_),
    .S(net233),
    .X(_0052_));
 sg13g2_mux2_1 _1203_ (.A0(\top_inst.sndgen_inst.lfsr[1] ),
    .A1(net17),
    .S(net233),
    .X(_0053_));
 sg13g2_mux2_1 _1204_ (.A0(net111),
    .A1(net193),
    .S(net233),
    .X(_0054_));
 sg13g2_mux2_1 _1205_ (.A0(\top_inst.sndgen_inst.lfsr[3] ),
    .A1(net111),
    .S(net233),
    .X(_0055_));
 sg13g2_nand2_1 _1206_ (.Y(_0497_),
    .A(net55),
    .B(net229));
 sg13g2_xnor2_1 _1207_ (.Y(_0498_),
    .A(net256),
    .B(\top_inst.sndgen_inst.lfsr[3] ));
 sg13g2_o21ai_1 _1208_ (.B1(_0497_),
    .Y(_0056_),
    .A1(net229),
    .A2(_0498_));
 sg13g2_nand2_1 _1209_ (.Y(_0499_),
    .A(net314),
    .B(net229));
 sg13g2_xnor2_1 _1210_ (.Y(_0500_),
    .A(net256),
    .B(net55));
 sg13g2_o21ai_1 _1211_ (.B1(_0499_),
    .Y(_0057_),
    .A1(net229),
    .A2(_0500_));
 sg13g2_nor2_1 _1212_ (.A(net51),
    .B(net233),
    .Y(_0501_));
 sg13g2_nand2b_1 _1213_ (.Y(_0502_),
    .B(net256),
    .A_N(\top_inst.sndgen_inst.lfsr[5] ));
 sg13g2_xnor2_1 _1214_ (.Y(_0503_),
    .A(net256),
    .B(\top_inst.sndgen_inst.lfsr[5] ));
 sg13g2_a21oi_1 _1215_ (.A1(net233),
    .A2(_0503_),
    .Y(_0058_),
    .B1(_0501_));
 sg13g2_mux2_1 _1216_ (.A0(net256),
    .A1(net51),
    .S(net233),
    .X(_0059_));
 sg13g2_nand2b_1 _1217_ (.Y(_0504_),
    .B(net175),
    .A_N(net220));
 sg13g2_a21oi_1 _1218_ (.A1(\top_inst.vga_inst.sx1[0] ),
    .A2(net219),
    .Y(_0505_),
    .B1(net222));
 sg13g2_a22oi_1 _1219_ (.Y(_0060_),
    .B1(_0504_),
    .B2(_0505_),
    .A2(net222),
    .A1(_0265_));
 sg13g2_nand2b_1 _1220_ (.Y(_0506_),
    .B(\top_inst.vga_inst.sr1[1] ),
    .A_N(net220));
 sg13g2_a21oi_1 _1221_ (.A1(\top_inst.vga_inst.sx1[1] ),
    .A2(net219),
    .Y(_0507_),
    .B1(net222));
 sg13g2_a22oi_1 _1222_ (.Y(_0061_),
    .B1(_0506_),
    .B2(_0507_),
    .A2(net222),
    .A1(_0264_));
 sg13g2_a21oi_1 _1223_ (.A1(_0245_),
    .A2(net219),
    .Y(_0508_),
    .B1(net223));
 sg13g2_o21ai_1 _1224_ (.B1(_0508_),
    .Y(_0509_),
    .A1(\top_inst.vga_inst.sr1[2] ),
    .A2(net219));
 sg13g2_o21ai_1 _1225_ (.B1(_0509_),
    .Y(_0062_),
    .A1(_0263_),
    .A2(net224));
 sg13g2_nor3_1 _1226_ (.A(\top_inst.vga_inst.sr1[3] ),
    .B(\top_inst.vga_inst.sx1[3] ),
    .C(net223),
    .Y(_0510_));
 sg13g2_a21oi_1 _1227_ (.A1(_0262_),
    .A2(net223),
    .Y(_0063_),
    .B1(_0510_));
 sg13g2_nor2_1 _1228_ (.A(net310),
    .B(net234),
    .Y(_0511_));
 sg13g2_a21oi_1 _1229_ (.A1(_0357_),
    .A2(net235),
    .Y(_0064_),
    .B1(_0511_));
 sg13g2_nor2_1 _1230_ (.A(net352),
    .B(net238),
    .Y(_0512_));
 sg13g2_a21oi_1 _1231_ (.A1(net238),
    .A2(_0361_),
    .Y(_0065_),
    .B1(_0512_));
 sg13g2_nor2_1 _1232_ (.A(net215),
    .B(net238),
    .Y(_0513_));
 sg13g2_a21oi_1 _1233_ (.A1(net238),
    .A2(_0355_),
    .Y(_0066_),
    .B1(_0513_));
 sg13g2_nor2_1 _1234_ (.A(net339),
    .B(net237),
    .Y(_0514_));
 sg13g2_a21oi_1 _1235_ (.A1(net237),
    .A2(_0353_),
    .Y(_0067_),
    .B1(_0514_));
 sg13g2_o21ai_1 _1236_ (.B1(net223),
    .Y(_0515_),
    .A1(net242),
    .A2(net62));
 sg13g2_a21oi_1 _1237_ (.A1(net242),
    .A2(net62),
    .Y(_0068_),
    .B1(_0515_));
 sg13g2_and3_1 _1238_ (.X(_0516_),
    .A(net242),
    .B(net62),
    .C(net27));
 sg13g2_a21oi_1 _1239_ (.A1(net242),
    .A2(\top_inst.vga_inst.x1[0] ),
    .Y(_0517_),
    .B1(net27));
 sg13g2_nor3_1 _1240_ (.A(net224),
    .B(_0516_),
    .C(net28),
    .Y(_0069_));
 sg13g2_and2_1 _1241_ (.A(net139),
    .B(_0516_),
    .X(_0518_));
 sg13g2_nor2_1 _1242_ (.A(net139),
    .B(_0516_),
    .Y(_0519_));
 sg13g2_nor3_1 _1243_ (.A(_0481_),
    .B(_0518_),
    .C(net140),
    .Y(_0070_));
 sg13g2_nor2_1 _1244_ (.A(net294),
    .B(_0518_),
    .Y(_0520_));
 sg13g2_and2_1 _1245_ (.A(net294),
    .B(_0518_),
    .X(_0521_));
 sg13g2_nor3_1 _1246_ (.A(_0481_),
    .B(_0520_),
    .C(_0521_),
    .Y(_0071_));
 sg13g2_nor2_1 _1247_ (.A(net340),
    .B(_0521_),
    .Y(_0522_));
 sg13g2_and2_1 _1248_ (.A(net340),
    .B(_0521_),
    .X(_0523_));
 sg13g2_nor3_1 _1249_ (.A(net224),
    .B(_0522_),
    .C(_0523_),
    .Y(_0072_));
 sg13g2_and2_1 _1250_ (.A(net364),
    .B(_0523_),
    .X(_0524_));
 sg13g2_o21ai_1 _1251_ (.B1(net223),
    .Y(_0525_),
    .A1(net364),
    .A2(_0523_));
 sg13g2_nor2_1 _1252_ (.A(_0524_),
    .B(_0525_),
    .Y(_0073_));
 sg13g2_nand2_1 _1253_ (.Y(_0526_),
    .A(net357),
    .B(_0524_));
 sg13g2_o21ai_1 _1254_ (.B1(net222),
    .Y(_0527_),
    .A1(net357),
    .A2(_0524_));
 sg13g2_nor2b_1 _1255_ (.A(net358),
    .B_N(_0526_),
    .Y(_0074_));
 sg13g2_xnor2_1 _1256_ (.Y(_0528_),
    .A(_0250_),
    .B(_0526_));
 sg13g2_nor2_1 _1257_ (.A(net224),
    .B(_0528_),
    .Y(_0075_));
 sg13g2_mux2_1 _1258_ (.A0(net175),
    .A1(net310),
    .S(net235),
    .X(_0076_));
 sg13g2_mux2_1 _1259_ (.A0(net352),
    .A1(net363),
    .S(_0436_),
    .X(_0077_));
 sg13g2_nor2_1 _1260_ (.A(net145),
    .B(net234),
    .Y(_0529_));
 sg13g2_a21oi_1 _1261_ (.A1(_0245_),
    .A2(net234),
    .Y(_0078_),
    .B1(_0529_));
 sg13g2_nor2_1 _1262_ (.A(net321),
    .B(net234),
    .Y(_0530_));
 sg13g2_a21oi_1 _1263_ (.A1(_0244_),
    .A2(net234),
    .Y(_0079_),
    .B1(_0530_));
 sg13g2_and2_1 _1264_ (.A(_0406_),
    .B(_0417_),
    .X(_0531_));
 sg13g2_nor2_1 _1265_ (.A(net249),
    .B(net59),
    .Y(_0532_));
 sg13g2_a21oi_1 _1266_ (.A1(net249),
    .A2(_0531_),
    .Y(_0080_),
    .B1(net60));
 sg13g2_nor2_2 _1267_ (.A(_0413_),
    .B(_0421_),
    .Y(_0533_));
 sg13g2_nor2_1 _1268_ (.A(net249),
    .B(net124),
    .Y(_0534_));
 sg13g2_a21oi_1 _1269_ (.A1(net249),
    .A2(_0533_),
    .Y(_0081_),
    .B1(net125));
 sg13g2_nor2_1 _1270_ (.A(_0251_),
    .B(\top_inst.sndgen_inst.rom_addr[1] ),
    .Y(_0535_));
 sg13g2_a21oi_2 _1271_ (.B1(_0421_),
    .Y(_0536_),
    .A2(_0535_),
    .A1(_0411_));
 sg13g2_nor2_1 _1272_ (.A(net249),
    .B(net153),
    .Y(_0537_));
 sg13g2_a21oi_1 _1273_ (.A1(net249),
    .A2(_0536_),
    .Y(_0082_),
    .B1(_0537_));
 sg13g2_xor2_1 _1274_ (.B(\top_inst.sndgen_inst.rom_addr[0] ),
    .A(\top_inst.sndgen_inst.rom_addr[1] ),
    .X(_0538_));
 sg13g2_a21oi_2 _1275_ (.B1(_0411_),
    .Y(_0539_),
    .A2(_0538_),
    .A1(_0407_));
 sg13g2_nor2_1 _1276_ (.A(net249),
    .B(net161),
    .Y(_0540_));
 sg13g2_a21oi_1 _1277_ (.A1(net249),
    .A2(_0539_),
    .Y(_0083_),
    .B1(_0540_));
 sg13g2_nor2_1 _1278_ (.A(net248),
    .B(net169),
    .Y(_0541_));
 sg13g2_a21oi_1 _1279_ (.A1(net248),
    .A2(_0409_),
    .Y(_0084_),
    .B1(_0541_));
 sg13g2_nor2_1 _1280_ (.A(net248),
    .B(net103),
    .Y(_0542_));
 sg13g2_a21oi_1 _1281_ (.A1(net248),
    .A2(_0415_),
    .Y(_0085_),
    .B1(net104));
 sg13g2_nor2_1 _1282_ (.A(net248),
    .B(net74),
    .Y(_0543_));
 sg13g2_a21oi_1 _1283_ (.A1(net248),
    .A2(_0419_),
    .Y(_0086_),
    .B1(net75));
 sg13g2_nor2_1 _1284_ (.A(net247),
    .B(net73),
    .Y(_0544_));
 sg13g2_a21oi_1 _1285_ (.A1(net247),
    .A2(_0422_),
    .Y(_0087_),
    .B1(_0544_));
 sg13g2_nor2_1 _1286_ (.A(net247),
    .B(net255),
    .Y(_0545_));
 sg13g2_a21oi_1 _1287_ (.A1(net247),
    .A2(net344),
    .Y(_0088_),
    .B1(_0545_));
 sg13g2_nor4_2 _1288_ (.A(net119),
    .B(\top_inst.sys_presc[2] ),
    .C(net49),
    .Y(_0546_),
    .D(_0402_));
 sg13g2_mux2_1 _1289_ (.A0(\top_inst.pwm_inst.cntr[0] ),
    .A1(net87),
    .S(_0546_),
    .X(_0089_));
 sg13g2_nand3_1 _1290_ (.B(net377),
    .C(_0546_),
    .A(\top_inst.pwm_inst.cntr[0] ),
    .Y(_0547_));
 sg13g2_a21o_1 _1291_ (.A2(_0546_),
    .A1(\top_inst.pwm_inst.cntr[0] ),
    .B1(net377),
    .X(_0548_));
 sg13g2_and2_1 _1292_ (.A(_0547_),
    .B(net378),
    .X(_0090_));
 sg13g2_nand4_1 _1293_ (.B(\top_inst.pwm_inst.cntr[2] ),
    .C(\top_inst.pwm_inst.cntr[1] ),
    .A(\top_inst.pwm_inst.cntr[0] ),
    .Y(_0549_),
    .D(_0546_));
 sg13g2_xnor2_1 _1294_ (.Y(_0091_),
    .A(net302),
    .B(_0547_));
 sg13g2_xnor2_1 _1295_ (.Y(_0092_),
    .A(net85),
    .B(_0549_));
 sg13g2_nand2_1 _1296_ (.Y(_0550_),
    .A(\top_inst.sndgen_inst.p_c2[0] ),
    .B(net226));
 sg13g2_xnor2_1 _1297_ (.Y(_0093_),
    .A(net40),
    .B(_0550_));
 sg13g2_nor2_1 _1298_ (.A(net155),
    .B(net226),
    .Y(_0551_));
 sg13g2_nand2_1 _1299_ (.Y(_0552_),
    .A(net44),
    .B(net40));
 sg13g2_nand2_1 _1300_ (.Y(_0553_),
    .A(\top_inst.sndgen_inst.p_c2[1] ),
    .B(\top_inst.sndgen_inst.phacc2[1] ));
 sg13g2_xnor2_1 _1301_ (.Y(_0554_),
    .A(net82),
    .B(net155));
 sg13g2_xnor2_1 _1302_ (.Y(_0555_),
    .A(_0552_),
    .B(_0554_));
 sg13g2_a21oi_1 _1303_ (.A1(net226),
    .A2(_0555_),
    .Y(_0094_),
    .B1(net156));
 sg13g2_nor2_1 _1304_ (.A(net134),
    .B(net226),
    .Y(_0556_));
 sg13g2_and2_1 _1305_ (.A(\top_inst.sndgen_inst.p_c2[2] ),
    .B(\top_inst.sndgen_inst.phacc2[2] ),
    .X(_0557_));
 sg13g2_xor2_1 _1306_ (.B(\top_inst.sndgen_inst.phacc2[2] ),
    .A(\top_inst.sndgen_inst.p_c2[2] ),
    .X(_0558_));
 sg13g2_o21ai_1 _1307_ (.B1(_0553_),
    .Y(_0559_),
    .A1(_0552_),
    .A2(_0554_));
 sg13g2_xnor2_1 _1308_ (.Y(_0560_),
    .A(_0558_),
    .B(_0559_));
 sg13g2_a21oi_1 _1309_ (.A1(net226),
    .A2(_0560_),
    .Y(_0095_),
    .B1(net135));
 sg13g2_nor2_1 _1310_ (.A(net179),
    .B(net225),
    .Y(_0561_));
 sg13g2_nand2_1 _1311_ (.Y(_0562_),
    .A(\top_inst.sndgen_inst.p_c2[3] ),
    .B(net392));
 sg13g2_xnor2_1 _1312_ (.Y(_0563_),
    .A(\top_inst.sndgen_inst.p_c2[3] ),
    .B(net179));
 sg13g2_a21oi_2 _1313_ (.B1(_0557_),
    .Y(_0564_),
    .A2(_0559_),
    .A1(_0558_));
 sg13g2_xnor2_1 _1314_ (.Y(_0565_),
    .A(_0563_),
    .B(_0564_));
 sg13g2_a21oi_1 _1315_ (.A1(net225),
    .A2(_0565_),
    .Y(_0096_),
    .B1(_0561_));
 sg13g2_nor2_1 _1316_ (.A(net154),
    .B(net225),
    .Y(_0566_));
 sg13g2_and2_1 _1317_ (.A(\top_inst.sndgen_inst.p_c2[4] ),
    .B(\top_inst.sndgen_inst.phacc2[4] ),
    .X(_0567_));
 sg13g2_xor2_1 _1318_ (.B(net154),
    .A(net97),
    .X(_0568_));
 sg13g2_o21ai_1 _1319_ (.B1(_0562_),
    .Y(_0569_),
    .A1(_0563_),
    .A2(_0564_));
 sg13g2_xnor2_1 _1320_ (.Y(_0570_),
    .A(_0568_),
    .B(_0569_));
 sg13g2_a21oi_1 _1321_ (.A1(net225),
    .A2(_0570_),
    .Y(_0097_),
    .B1(_0566_));
 sg13g2_a21oi_1 _1322_ (.A1(_0568_),
    .A2(_0569_),
    .Y(_0571_),
    .B1(_0567_));
 sg13g2_nor2_1 _1323_ (.A(\top_inst.sndgen_inst.p_c2[5] ),
    .B(\top_inst.sndgen_inst.phacc2[5] ),
    .Y(_0572_));
 sg13g2_xor2_1 _1324_ (.B(\top_inst.sndgen_inst.phacc2[5] ),
    .A(\top_inst.sndgen_inst.p_c2[5] ),
    .X(_0573_));
 sg13g2_xnor2_1 _1325_ (.Y(_0574_),
    .A(_0571_),
    .B(_0573_));
 sg13g2_mux2_1 _1326_ (.A0(net334),
    .A1(_0574_),
    .S(net227),
    .X(_0098_));
 sg13g2_nand2_1 _1327_ (.Y(_0575_),
    .A(net89),
    .B(\top_inst.sndgen_inst.phacc2[6] ));
 sg13g2_xnor2_1 _1328_ (.Y(_0576_),
    .A(net89),
    .B(net177));
 sg13g2_a221oi_1 _1329_ (.B2(_0569_),
    .C1(_0567_),
    .B1(_0568_),
    .A1(\top_inst.sndgen_inst.p_c2[5] ),
    .Y(_0577_),
    .A2(\top_inst.sndgen_inst.phacc2[5] ));
 sg13g2_or3_1 _1330_ (.A(_0572_),
    .B(_0576_),
    .C(_0577_),
    .X(_0578_));
 sg13g2_o21ai_1 _1331_ (.B1(_0576_),
    .Y(_0579_),
    .A1(_0572_),
    .A2(_0577_));
 sg13g2_nand3_1 _1332_ (.B(_0578_),
    .C(_0579_),
    .A(net227),
    .Y(_0580_));
 sg13g2_o21ai_1 _1333_ (.B1(_0580_),
    .Y(_0099_),
    .A1(_0266_),
    .A2(net227));
 sg13g2_nand2_1 _1334_ (.Y(_0581_),
    .A(\top_inst.sndgen_inst.p_c2[7] ),
    .B(\top_inst.sndgen_inst.phacc2[7] ));
 sg13g2_xnor2_1 _1335_ (.Y(_0582_),
    .A(\top_inst.sndgen_inst.p_c2[7] ),
    .B(\top_inst.sndgen_inst.phacc2[7] ));
 sg13g2_a21o_1 _1336_ (.A2(_0578_),
    .A1(_0575_),
    .B1(_0582_),
    .X(_0583_));
 sg13g2_nand3_1 _1337_ (.B(_0578_),
    .C(_0582_),
    .A(_0575_),
    .Y(_0584_));
 sg13g2_nand3_1 _1338_ (.B(_0583_),
    .C(_0584_),
    .A(net225),
    .Y(_0585_));
 sg13g2_o21ai_1 _1339_ (.B1(_0585_),
    .Y(_0100_),
    .A1(_0267_),
    .A2(net225));
 sg13g2_nor2_1 _1340_ (.A(net34),
    .B(net227),
    .Y(_0586_));
 sg13g2_nand2_2 _1341_ (.Y(_0587_),
    .A(_0581_),
    .B(_0583_));
 sg13g2_xnor2_1 _1342_ (.Y(_0588_),
    .A(_0268_),
    .B(_0587_));
 sg13g2_a21oi_1 _1343_ (.A1(net227),
    .A2(_0588_),
    .Y(_0101_),
    .B1(_0586_));
 sg13g2_nand2b_1 _1344_ (.Y(_0589_),
    .B(net213),
    .A_N(net225));
 sg13g2_nand2_1 _1345_ (.Y(_0590_),
    .A(net243),
    .B(\top_inst.sndgen_inst.phacc2[9] ));
 sg13g2_xor2_1 _1346_ (.B(net213),
    .A(net243),
    .X(_0591_));
 sg13g2_a21oi_1 _1347_ (.A1(_0268_),
    .A2(_0587_),
    .Y(_0592_),
    .B1(_0591_));
 sg13g2_and2_1 _1348_ (.A(_0268_),
    .B(_0591_),
    .X(_0593_));
 sg13g2_nand2_1 _1349_ (.Y(_0594_),
    .A(_0587_),
    .B(_0593_));
 sg13g2_nand2_1 _1350_ (.Y(_0595_),
    .A(net227),
    .B(_0594_));
 sg13g2_o21ai_1 _1351_ (.B1(_0589_),
    .Y(_0102_),
    .A1(_0592_),
    .A2(_0595_));
 sg13g2_nor2_1 _1352_ (.A(net338),
    .B(net227),
    .Y(_0596_));
 sg13g2_a22oi_1 _1353_ (.Y(_0597_),
    .B1(_0587_),
    .B2(_0593_),
    .A2(\top_inst.sndgen_inst.phacc2[9] ),
    .A1(net243));
 sg13g2_nand2_1 _1354_ (.Y(_0598_),
    .A(net243),
    .B(\top_inst.sndgen_inst.phacc2[10] ));
 sg13g2_nor2_1 _1355_ (.A(net243),
    .B(\top_inst.sndgen_inst.phacc2[10] ),
    .Y(_0599_));
 sg13g2_xor2_1 _1356_ (.B(\top_inst.sndgen_inst.phacc2[10] ),
    .A(net243),
    .X(_0600_));
 sg13g2_xor2_1 _1357_ (.B(_0600_),
    .A(_0597_),
    .X(_0601_));
 sg13g2_a21oi_1 _1358_ (.A1(net227),
    .A2(_0601_),
    .Y(_0103_),
    .B1(_0596_));
 sg13g2_o21ai_1 _1359_ (.B1(_0598_),
    .Y(_0602_),
    .A1(_0597_),
    .A2(_0599_));
 sg13g2_xor2_1 _1360_ (.B(\top_inst.sndgen_inst.phacc2[11] ),
    .A(net244),
    .X(_0603_));
 sg13g2_xor2_1 _1361_ (.B(_0603_),
    .A(_0602_),
    .X(_0604_));
 sg13g2_mux2_1 _1362_ (.A0(net167),
    .A1(_0604_),
    .S(net225),
    .X(_0104_));
 sg13g2_nor2_1 _1363_ (.A(net142),
    .B(_0434_),
    .Y(_0605_));
 sg13g2_nand2_1 _1364_ (.Y(_0606_),
    .A(net244),
    .B(\top_inst.sndgen_inst.phacc2[12] ));
 sg13g2_xor2_1 _1365_ (.B(\top_inst.sndgen_inst.phacc2[12] ),
    .A(net243),
    .X(_0607_));
 sg13g2_nand3_1 _1366_ (.B(_0600_),
    .C(_0603_),
    .A(_0593_),
    .Y(_0608_));
 sg13g2_a21oi_1 _1367_ (.A1(_0581_),
    .A2(_0583_),
    .Y(_0609_),
    .B1(_0608_));
 sg13g2_o21ai_1 _1368_ (.B1(net243),
    .Y(_0610_),
    .A1(\top_inst.sndgen_inst.phacc2[10] ),
    .A2(\top_inst.sndgen_inst.phacc2[11] ));
 sg13g2_nand2_1 _1369_ (.Y(_0611_),
    .A(_0590_),
    .B(_0610_));
 sg13g2_o21ai_1 _1370_ (.B1(_0607_),
    .Y(_0612_),
    .A1(_0609_),
    .A2(_0611_));
 sg13g2_or3_1 _1371_ (.A(_0607_),
    .B(_0609_),
    .C(_0611_),
    .X(_0613_));
 sg13g2_nand2_1 _1372_ (.Y(_0614_),
    .A(_0612_),
    .B(_0613_));
 sg13g2_a21oi_1 _1373_ (.A1(_0434_),
    .A2(_0614_),
    .Y(_0105_),
    .B1(net143));
 sg13g2_nand2_1 _1374_ (.Y(_0615_),
    .A(_0606_),
    .B(_0612_));
 sg13g2_xnor2_1 _1375_ (.Y(_0616_),
    .A(\top_inst.sndgen_inst.phacc2[13] ),
    .B(net244));
 sg13g2_xnor2_1 _1376_ (.Y(_0617_),
    .A(_0615_),
    .B(_0616_));
 sg13g2_mux2_1 _1377_ (.A0(net330),
    .A1(_0617_),
    .S(_0437_),
    .X(_0106_));
 sg13g2_nor2_1 _1378_ (.A(net250),
    .B(net44),
    .Y(_0618_));
 sg13g2_a21oi_1 _1379_ (.A1(net250),
    .A2(_0531_),
    .Y(_0107_),
    .B1(_0618_));
 sg13g2_nor2_1 _1380_ (.A(net250),
    .B(net82),
    .Y(_0619_));
 sg13g2_a21oi_1 _1381_ (.A1(net250),
    .A2(_0533_),
    .Y(_0108_),
    .B1(_0619_));
 sg13g2_nor2_1 _1382_ (.A(net250),
    .B(net77),
    .Y(_0620_));
 sg13g2_a21oi_1 _1383_ (.A1(net250),
    .A2(_0536_),
    .Y(_0109_),
    .B1(_0620_));
 sg13g2_nor2_1 _1384_ (.A(net251),
    .B(net101),
    .Y(_0621_));
 sg13g2_a21oi_1 _1385_ (.A1(net251),
    .A2(_0539_),
    .Y(_0110_),
    .B1(_0621_));
 sg13g2_nor2_1 _1386_ (.A(net251),
    .B(net97),
    .Y(_0622_));
 sg13g2_a21oi_1 _1387_ (.A1(net251),
    .A2(_0409_),
    .Y(_0111_),
    .B1(_0622_));
 sg13g2_nor2_1 _1388_ (.A(net251),
    .B(net319),
    .Y(_0623_));
 sg13g2_a21oi_1 _1389_ (.A1(net251),
    .A2(_0415_),
    .Y(_0112_),
    .B1(_0623_));
 sg13g2_nor2_1 _1390_ (.A(net252),
    .B(net89),
    .Y(_0624_));
 sg13g2_a21oi_1 _1391_ (.A1(net252),
    .A2(_0419_),
    .Y(_0113_),
    .B1(net90));
 sg13g2_nor2_1 _1392_ (.A(net252),
    .B(net207),
    .Y(_0625_));
 sg13g2_a21oi_1 _1393_ (.A1(net252),
    .A2(_0422_),
    .Y(_0114_),
    .B1(_0625_));
 sg13g2_nor2_1 _1394_ (.A(net251),
    .B(net244),
    .Y(_0626_));
 sg13g2_a21oi_1 _1395_ (.A1(net251),
    .A2(net344),
    .Y(_0115_),
    .B1(_0626_));
 sg13g2_nand2_1 _1396_ (.Y(_0627_),
    .A(\top_inst.sndgen_inst.p_c3[0] ),
    .B(net230));
 sg13g2_xnor2_1 _1397_ (.Y(_0116_),
    .A(net38),
    .B(_0627_));
 sg13g2_nor2_1 _1398_ (.A(net151),
    .B(net230),
    .Y(_0628_));
 sg13g2_nand2_1 _1399_ (.Y(_0629_),
    .A(net59),
    .B(net38));
 sg13g2_nand2_1 _1400_ (.Y(_0630_),
    .A(\top_inst.sndgen_inst.p_c3[1] ),
    .B(\top_inst.sndgen_inst.phacc3[1] ));
 sg13g2_xnor2_1 _1401_ (.Y(_0631_),
    .A(net124),
    .B(net151));
 sg13g2_xnor2_1 _1402_ (.Y(_0632_),
    .A(_0629_),
    .B(_0631_));
 sg13g2_a21oi_1 _1403_ (.A1(net230),
    .A2(_0632_),
    .Y(_0117_),
    .B1(_0628_));
 sg13g2_nor2_1 _1404_ (.A(net198),
    .B(net231),
    .Y(_0633_));
 sg13g2_and2_1 _1405_ (.A(net388),
    .B(\top_inst.sndgen_inst.phacc3[2] ),
    .X(_0634_));
 sg13g2_xor2_1 _1406_ (.B(net198),
    .A(net153),
    .X(_0635_));
 sg13g2_o21ai_1 _1407_ (.B1(_0630_),
    .Y(_0636_),
    .A1(_0629_),
    .A2(_0631_));
 sg13g2_xnor2_1 _1408_ (.Y(_0637_),
    .A(_0635_),
    .B(_0636_));
 sg13g2_a21oi_1 _1409_ (.A1(net231),
    .A2(_0637_),
    .Y(_0118_),
    .B1(_0633_));
 sg13g2_nor2_1 _1410_ (.A(net133),
    .B(net231),
    .Y(_0638_));
 sg13g2_nand2_1 _1411_ (.Y(_0639_),
    .A(\top_inst.sndgen_inst.p_c3[3] ),
    .B(\top_inst.sndgen_inst.phacc3[3] ));
 sg13g2_xnor2_1 _1412_ (.Y(_0640_),
    .A(\top_inst.sndgen_inst.p_c3[3] ),
    .B(net133));
 sg13g2_a21oi_1 _1413_ (.A1(_0635_),
    .A2(_0636_),
    .Y(_0641_),
    .B1(net389));
 sg13g2_xnor2_1 _1414_ (.Y(_0642_),
    .A(_0640_),
    .B(_0641_));
 sg13g2_a21oi_1 _1415_ (.A1(net231),
    .A2(net390),
    .Y(_0119_),
    .B1(_0638_));
 sg13g2_nor2_1 _1416_ (.A(net83),
    .B(net232),
    .Y(_0643_));
 sg13g2_and2_1 _1417_ (.A(\top_inst.sndgen_inst.p_c3[4] ),
    .B(\top_inst.sndgen_inst.phacc3[4] ),
    .X(_0644_));
 sg13g2_xor2_1 _1418_ (.B(net83),
    .A(\top_inst.sndgen_inst.p_c3[4] ),
    .X(_0645_));
 sg13g2_o21ai_1 _1419_ (.B1(_0639_),
    .Y(_0646_),
    .A1(_0640_),
    .A2(_0641_));
 sg13g2_xnor2_1 _1420_ (.Y(_0647_),
    .A(_0645_),
    .B(_0646_));
 sg13g2_a21oi_1 _1421_ (.A1(net232),
    .A2(_0647_),
    .Y(_0120_),
    .B1(_0643_));
 sg13g2_a21oi_2 _1422_ (.B1(_0644_),
    .Y(_0648_),
    .A2(_0646_),
    .A1(_0645_));
 sg13g2_nor2_1 _1423_ (.A(\top_inst.sndgen_inst.p_c3[5] ),
    .B(\top_inst.sndgen_inst.phacc3[5] ),
    .Y(_0649_));
 sg13g2_nand2_1 _1424_ (.Y(_0650_),
    .A(\top_inst.sndgen_inst.p_c3[5] ),
    .B(\top_inst.sndgen_inst.phacc3[5] ));
 sg13g2_nor2b_1 _1425_ (.A(_0649_),
    .B_N(_0650_),
    .Y(_0651_));
 sg13g2_xnor2_1 _1426_ (.Y(_0652_),
    .A(_0648_),
    .B(_0651_));
 sg13g2_mux2_1 _1427_ (.A0(net121),
    .A1(_0652_),
    .S(_0432_),
    .X(_0121_));
 sg13g2_and2_1 _1428_ (.A(\top_inst.sndgen_inst.p_c3[6] ),
    .B(\top_inst.sndgen_inst.phacc3[6] ),
    .X(_0653_));
 sg13g2_xor2_1 _1429_ (.B(\top_inst.sndgen_inst.phacc3[6] ),
    .A(\top_inst.sndgen_inst.p_c3[6] ),
    .X(_0654_));
 sg13g2_o21ai_1 _1430_ (.B1(_0650_),
    .Y(_0655_),
    .A1(_0648_),
    .A2(_0649_));
 sg13g2_o21ai_1 _1431_ (.B1(net236),
    .Y(_0656_),
    .A1(_0654_),
    .A2(_0655_));
 sg13g2_a21oi_1 _1432_ (.A1(_0654_),
    .A2(_0655_),
    .Y(_0657_),
    .B1(_0656_));
 sg13g2_a21o_1 _1433_ (.A2(net229),
    .A1(net185),
    .B1(_0657_),
    .X(_0122_));
 sg13g2_nor2_1 _1434_ (.A(net96),
    .B(net237),
    .Y(_0658_));
 sg13g2_nand2_1 _1435_ (.Y(_0659_),
    .A(\top_inst.sndgen_inst.p_c3[7] ),
    .B(\top_inst.sndgen_inst.phacc3[7] ));
 sg13g2_xnor2_1 _1436_ (.Y(_0660_),
    .A(net73),
    .B(net96));
 sg13g2_a21oi_1 _1437_ (.A1(_0654_),
    .A2(_0655_),
    .Y(_0661_),
    .B1(_0653_));
 sg13g2_xnor2_1 _1438_ (.Y(_0662_),
    .A(_0660_),
    .B(_0661_));
 sg13g2_a21oi_1 _1439_ (.A1(net237),
    .A2(_0662_),
    .Y(_0123_),
    .B1(_0658_));
 sg13g2_o21ai_1 _1440_ (.B1(_0659_),
    .Y(_0663_),
    .A1(_0660_),
    .A2(_0661_));
 sg13g2_and2_1 _1441_ (.A(_0269_),
    .B(_0663_),
    .X(_0664_));
 sg13g2_nand2_1 _1442_ (.Y(_0665_),
    .A(net19),
    .B(net228));
 sg13g2_o21ai_1 _1443_ (.B1(net235),
    .Y(_0666_),
    .A1(_0269_),
    .A2(_0663_));
 sg13g2_o21ai_1 _1444_ (.B1(_0665_),
    .Y(_0124_),
    .A1(_0664_),
    .A2(_0666_));
 sg13g2_nand2_1 _1445_ (.Y(_0667_),
    .A(net113),
    .B(net228));
 sg13g2_nand2_1 _1446_ (.Y(_0668_),
    .A(net255),
    .B(\top_inst.sndgen_inst.phacc3[9] ));
 sg13g2_xor2_1 _1447_ (.B(net113),
    .A(net255),
    .X(_0669_));
 sg13g2_nor2b_1 _1448_ (.A(_0011_),
    .B_N(_0669_),
    .Y(_0670_));
 sg13g2_nand2_1 _1449_ (.Y(_0671_),
    .A(_0663_),
    .B(_0670_));
 sg13g2_o21ai_1 _1450_ (.B1(_0671_),
    .Y(_0672_),
    .A1(_0664_),
    .A2(_0669_));
 sg13g2_o21ai_1 _1451_ (.B1(_0667_),
    .Y(_0125_),
    .A1(net228),
    .A2(_0672_));
 sg13g2_nor2_1 _1452_ (.A(net95),
    .B(net237),
    .Y(_0673_));
 sg13g2_nor2_1 _1453_ (.A(net254),
    .B(\top_inst.sndgen_inst.phacc3[10] ),
    .Y(_0674_));
 sg13g2_nand2_1 _1454_ (.Y(_0675_),
    .A(net254),
    .B(net391));
 sg13g2_nor2b_1 _1455_ (.A(_0674_),
    .B_N(_0675_),
    .Y(_0676_));
 sg13g2_a22oi_1 _1456_ (.Y(_0677_),
    .B1(_0663_),
    .B2(_0670_),
    .A2(net393),
    .A1(net255));
 sg13g2_xor2_1 _1457_ (.B(_0677_),
    .A(_0676_),
    .X(_0678_));
 sg13g2_a21oi_1 _1458_ (.A1(net238),
    .A2(_0678_),
    .Y(_0126_),
    .B1(_0673_));
 sg13g2_o21ai_1 _1459_ (.B1(_0675_),
    .Y(_0679_),
    .A1(_0674_),
    .A2(_0677_));
 sg13g2_xor2_1 _1460_ (.B(net68),
    .A(net254),
    .X(_0680_));
 sg13g2_nand2_1 _1461_ (.Y(_0681_),
    .A(net68),
    .B(_0436_));
 sg13g2_xnor2_1 _1462_ (.Y(_0682_),
    .A(_0679_),
    .B(_0680_));
 sg13g2_o21ai_1 _1463_ (.B1(_0681_),
    .Y(_0127_),
    .A1(_0433_),
    .A2(_0682_));
 sg13g2_nor2_1 _1464_ (.A(net298),
    .B(net237),
    .Y(_0683_));
 sg13g2_and3_1 _1465_ (.X(_0684_),
    .A(_0670_),
    .B(_0676_),
    .C(_0680_));
 sg13g2_nand2_1 _1466_ (.Y(_0685_),
    .A(_0668_),
    .B(_0675_));
 sg13g2_a221oi_1 _1467_ (.B2(_0684_),
    .C1(_0685_),
    .B1(_0663_),
    .A1(net254),
    .Y(_0686_),
    .A2(net68));
 sg13g2_nand2_1 _1468_ (.Y(_0687_),
    .A(net254),
    .B(\top_inst.sndgen_inst.phacc3[12] ));
 sg13g2_nor2_1 _1469_ (.A(net254),
    .B(\top_inst.sndgen_inst.phacc3[12] ),
    .Y(_0688_));
 sg13g2_xnor2_1 _1470_ (.Y(_0689_),
    .A(net254),
    .B(net298));
 sg13g2_xnor2_1 _1471_ (.Y(_0690_),
    .A(_0686_),
    .B(_0689_));
 sg13g2_a21oi_1 _1472_ (.A1(net237),
    .A2(_0690_),
    .Y(_0128_),
    .B1(_0683_));
 sg13g2_o21ai_1 _1473_ (.B1(_0687_),
    .Y(_0691_),
    .A1(_0686_),
    .A2(_0688_));
 sg13g2_xor2_1 _1474_ (.B(net254),
    .A(net311),
    .X(_0692_));
 sg13g2_xnor2_1 _1475_ (.Y(_0693_),
    .A(_0691_),
    .B(_0692_));
 sg13g2_nor2_1 _1476_ (.A(net311),
    .B(net235),
    .Y(_0694_));
 sg13g2_a21oi_1 _1477_ (.A1(net235),
    .A2(_0693_),
    .Y(_0129_),
    .B1(_0694_));
 sg13g2_nand2_1 _1478_ (.Y(_0695_),
    .A(\top_inst.sndgen_inst.p_c4[0] ),
    .B(net230));
 sg13g2_xnor2_1 _1479_ (.Y(_0130_),
    .A(net36),
    .B(_0695_));
 sg13g2_nor2_1 _1480_ (.A(net200),
    .B(net230),
    .Y(_0696_));
 sg13g2_nand2_1 _1481_ (.Y(_0697_),
    .A(net127),
    .B(net36));
 sg13g2_nand2_1 _1482_ (.Y(_0698_),
    .A(\top_inst.sndgen_inst.p_c4[1] ),
    .B(\top_inst.sndgen_inst.phacc4[1] ));
 sg13g2_xnor2_1 _1483_ (.Y(_0699_),
    .A(\top_inst.sndgen_inst.p_c4[1] ),
    .B(net200));
 sg13g2_xnor2_1 _1484_ (.Y(_0700_),
    .A(_0697_),
    .B(_0699_));
 sg13g2_a21oi_1 _1485_ (.A1(net230),
    .A2(_0700_),
    .Y(_0131_),
    .B1(_0696_));
 sg13g2_nor2_1 _1486_ (.A(net99),
    .B(net232),
    .Y(_0701_));
 sg13g2_and2_1 _1487_ (.A(\top_inst.sndgen_inst.p_c4[2] ),
    .B(\top_inst.sndgen_inst.phacc4[2] ),
    .X(_0702_));
 sg13g2_xor2_1 _1488_ (.B(net99),
    .A(\top_inst.sndgen_inst.p_c4[2] ),
    .X(_0703_));
 sg13g2_o21ai_1 _1489_ (.B1(_0698_),
    .Y(_0704_),
    .A1(_0697_),
    .A2(_0699_));
 sg13g2_xnor2_1 _1490_ (.Y(_0705_),
    .A(_0703_),
    .B(_0704_));
 sg13g2_a21oi_1 _1491_ (.A1(net232),
    .A2(_0705_),
    .Y(_0132_),
    .B1(_0701_));
 sg13g2_nor2_1 _1492_ (.A(net209),
    .B(net232),
    .Y(_0706_));
 sg13g2_nand2_1 _1493_ (.Y(_0707_),
    .A(\top_inst.sndgen_inst.p_c4[3] ),
    .B(\top_inst.sndgen_inst.phacc4[3] ));
 sg13g2_xnor2_1 _1494_ (.Y(_0708_),
    .A(\top_inst.sndgen_inst.p_c4[3] ),
    .B(net209));
 sg13g2_a21oi_1 _1495_ (.A1(_0703_),
    .A2(_0704_),
    .Y(_0709_),
    .B1(_0702_));
 sg13g2_xnor2_1 _1496_ (.Y(_0710_),
    .A(_0708_),
    .B(_0709_));
 sg13g2_a21oi_1 _1497_ (.A1(net232),
    .A2(_0710_),
    .Y(_0133_),
    .B1(_0706_));
 sg13g2_nor2_1 _1498_ (.A(net211),
    .B(net236),
    .Y(_0711_));
 sg13g2_and2_1 _1499_ (.A(\top_inst.sndgen_inst.p_c4[4] ),
    .B(\top_inst.sndgen_inst.phacc4[4] ),
    .X(_0712_));
 sg13g2_xor2_1 _1500_ (.B(net211),
    .A(\top_inst.sndgen_inst.p_c4[4] ),
    .X(_0713_));
 sg13g2_o21ai_1 _1501_ (.B1(_0707_),
    .Y(_0714_),
    .A1(_0708_),
    .A2(_0709_));
 sg13g2_xnor2_1 _1502_ (.Y(_0715_),
    .A(_0713_),
    .B(_0714_));
 sg13g2_a21oi_1 _1503_ (.A1(net236),
    .A2(_0715_),
    .Y(_0134_),
    .B1(_0711_));
 sg13g2_a21oi_2 _1504_ (.B1(_0712_),
    .Y(_0716_),
    .A2(_0714_),
    .A1(_0713_));
 sg13g2_nor2_1 _1505_ (.A(\top_inst.sndgen_inst.p_c4[5] ),
    .B(\top_inst.sndgen_inst.phacc4[5] ),
    .Y(_0717_));
 sg13g2_nand2_1 _1506_ (.Y(_0718_),
    .A(\top_inst.sndgen_inst.p_c4[5] ),
    .B(\top_inst.sndgen_inst.phacc4[5] ));
 sg13g2_nor2b_1 _1507_ (.A(_0717_),
    .B_N(_0718_),
    .Y(_0719_));
 sg13g2_xnor2_1 _1508_ (.Y(_0720_),
    .A(_0716_),
    .B(_0719_));
 sg13g2_mux2_1 _1509_ (.A0(net94),
    .A1(_0720_),
    .S(_0432_),
    .X(_0135_));
 sg13g2_and2_1 _1510_ (.A(\top_inst.sndgen_inst.p_c4[6] ),
    .B(\top_inst.sndgen_inst.phacc4[6] ),
    .X(_0721_));
 sg13g2_xor2_1 _1511_ (.B(\top_inst.sndgen_inst.phacc4[6] ),
    .A(\top_inst.sndgen_inst.p_c4[6] ),
    .X(_0722_));
 sg13g2_o21ai_1 _1512_ (.B1(_0718_),
    .Y(_0723_),
    .A1(_0716_),
    .A2(_0717_));
 sg13g2_o21ai_1 _1513_ (.B1(net236),
    .Y(_0724_),
    .A1(_0722_),
    .A2(_0723_));
 sg13g2_a21oi_1 _1514_ (.A1(_0722_),
    .A2(_0723_),
    .Y(_0725_),
    .B1(_0724_));
 sg13g2_a21o_1 _1515_ (.A2(net228),
    .A1(net164),
    .B1(_0725_),
    .X(_0136_));
 sg13g2_nor2_1 _1516_ (.A(net162),
    .B(net239),
    .Y(_0726_));
 sg13g2_nand2_1 _1517_ (.Y(_0727_),
    .A(\top_inst.sndgen_inst.p_c4[7] ),
    .B(\top_inst.sndgen_inst.phacc4[7] ));
 sg13g2_xnor2_1 _1518_ (.Y(_0728_),
    .A(\top_inst.sndgen_inst.p_c4[7] ),
    .B(net162));
 sg13g2_a21oi_2 _1519_ (.B1(_0721_),
    .Y(_0729_),
    .A2(_0723_),
    .A1(_0722_));
 sg13g2_xnor2_1 _1520_ (.Y(_0730_),
    .A(_0728_),
    .B(_0729_));
 sg13g2_a21oi_1 _1521_ (.A1(net239),
    .A2(_0730_),
    .Y(_0137_),
    .B1(_0726_));
 sg13g2_o21ai_1 _1522_ (.B1(_0727_),
    .Y(_0731_),
    .A1(_0728_),
    .A2(_0729_));
 sg13g2_and2_1 _1523_ (.A(_0270_),
    .B(_0731_),
    .X(_0732_));
 sg13g2_nand2_1 _1524_ (.Y(_0733_),
    .A(net23),
    .B(net228));
 sg13g2_o21ai_1 _1525_ (.B1(net234),
    .Y(_0734_),
    .A1(_0270_),
    .A2(_0731_));
 sg13g2_o21ai_1 _1526_ (.B1(_0733_),
    .Y(_0138_),
    .A1(_0732_),
    .A2(_0734_));
 sg13g2_nand2_1 _1527_ (.Y(_0735_),
    .A(net115),
    .B(net228));
 sg13g2_nand2_1 _1528_ (.Y(_0736_),
    .A(net260),
    .B(\top_inst.sndgen_inst.phacc4[9] ));
 sg13g2_xor2_1 _1529_ (.B(net115),
    .A(net261),
    .X(_0737_));
 sg13g2_nor2b_1 _1530_ (.A(_0000_),
    .B_N(_0737_),
    .Y(_0738_));
 sg13g2_nand2_1 _1531_ (.Y(_0739_),
    .A(_0731_),
    .B(_0738_));
 sg13g2_o21ai_1 _1532_ (.B1(_0739_),
    .Y(_0740_),
    .A1(_0732_),
    .A2(_0737_));
 sg13g2_o21ai_1 _1533_ (.B1(_0735_),
    .Y(_0139_),
    .A1(net228),
    .A2(_0740_));
 sg13g2_nor2_1 _1534_ (.A(net69),
    .B(net239),
    .Y(_0741_));
 sg13g2_nor2_1 _1535_ (.A(net260),
    .B(\top_inst.sndgen_inst.phacc4[10] ),
    .Y(_0742_));
 sg13g2_nand2_1 _1536_ (.Y(_0743_),
    .A(net260),
    .B(\top_inst.sndgen_inst.phacc4[10] ));
 sg13g2_nor2b_1 _1537_ (.A(_0742_),
    .B_N(_0743_),
    .Y(_0744_));
 sg13g2_a22oi_1 _1538_ (.Y(_0745_),
    .B1(_0731_),
    .B2(_0738_),
    .A2(\top_inst.sndgen_inst.phacc4[9] ),
    .A1(net260));
 sg13g2_xor2_1 _1539_ (.B(_0745_),
    .A(_0744_),
    .X(_0746_));
 sg13g2_a21oi_1 _1540_ (.A1(net239),
    .A2(_0746_),
    .Y(_0140_),
    .B1(_0741_));
 sg13g2_o21ai_1 _1541_ (.B1(_0743_),
    .Y(_0179_),
    .A1(_0742_),
    .A2(_0745_));
 sg13g2_xor2_1 _1542_ (.B(net57),
    .A(net260),
    .X(_0180_));
 sg13g2_nand2_1 _1543_ (.Y(_0181_),
    .A(net57),
    .B(net228));
 sg13g2_xnor2_1 _1544_ (.Y(_0182_),
    .A(_0179_),
    .B(_0180_));
 sg13g2_o21ai_1 _1545_ (.B1(_0181_),
    .Y(_0141_),
    .A1(_0433_),
    .A2(_0182_));
 sg13g2_nor2_1 _1546_ (.A(net335),
    .B(net239),
    .Y(_0183_));
 sg13g2_and3_1 _1547_ (.X(_0184_),
    .A(_0738_),
    .B(_0744_),
    .C(_0180_));
 sg13g2_nand2_1 _1548_ (.Y(_0185_),
    .A(_0736_),
    .B(_0743_));
 sg13g2_a221oi_1 _1549_ (.B2(_0184_),
    .C1(_0185_),
    .B1(_0731_),
    .A1(net260),
    .Y(_0186_),
    .A2(net57));
 sg13g2_nand2_1 _1550_ (.Y(_0187_),
    .A(net261),
    .B(\top_inst.sndgen_inst.phacc4[12] ));
 sg13g2_nor2_1 _1551_ (.A(net260),
    .B(\top_inst.sndgen_inst.phacc4[12] ),
    .Y(_0188_));
 sg13g2_xnor2_1 _1552_ (.Y(_0189_),
    .A(net260),
    .B(net335));
 sg13g2_xnor2_1 _1553_ (.Y(_0190_),
    .A(_0186_),
    .B(_0189_));
 sg13g2_a21oi_1 _1554_ (.A1(net239),
    .A2(_0190_),
    .Y(_0142_),
    .B1(_0183_));
 sg13g2_nor2_1 _1555_ (.A(net317),
    .B(net234),
    .Y(_0191_));
 sg13g2_o21ai_1 _1556_ (.B1(_0187_),
    .Y(_0192_),
    .A1(_0186_),
    .A2(_0188_));
 sg13g2_xor2_1 _1557_ (.B(net261),
    .A(net317),
    .X(_0193_));
 sg13g2_xnor2_1 _1558_ (.Y(_0194_),
    .A(_0192_),
    .B(_0193_));
 sg13g2_a21oi_1 _1559_ (.A1(net234),
    .A2(_0194_),
    .Y(_0143_),
    .B1(_0191_));
 sg13g2_mux2_1 _1560_ (.A0(net325),
    .A1(_0016_),
    .S(net230),
    .X(_0144_));
 sg13g2_nand3_1 _1561_ (.B(\top_inst.sndgen_inst.slot_counter[1] ),
    .C(_0432_),
    .A(\top_inst.sndgen_inst.slot_counter[0] ),
    .Y(_0195_));
 sg13g2_nand2_1 _1562_ (.Y(_0196_),
    .A(\top_inst.sndgen_inst.slot_counter[0] ),
    .B(net230));
 sg13g2_xnor2_1 _1563_ (.Y(_0145_),
    .A(net202),
    .B(_0196_));
 sg13g2_nor2_1 _1564_ (.A(_0239_),
    .B(_0195_),
    .Y(_0197_));
 sg13g2_nor3_2 _1565_ (.A(_0239_),
    .B(_0240_),
    .C(_0196_),
    .Y(_0198_));
 sg13g2_xnor2_1 _1566_ (.Y(_0146_),
    .A(net183),
    .B(_0195_));
 sg13g2_xor2_1 _1567_ (.B(_0198_),
    .A(net196),
    .X(_0147_));
 sg13g2_a21oi_1 _1568_ (.A1(\top_inst.sndgen_inst.slot_counter[3] ),
    .A2(_0198_),
    .Y(_0199_),
    .B1(net108));
 sg13g2_nor2b_2 _1569_ (.A(_0426_),
    .B_N(_0198_),
    .Y(_0200_));
 sg13g2_nor2_1 _1570_ (.A(net109),
    .B(_0200_),
    .Y(_0148_));
 sg13g2_and4_1 _1571_ (.A(net108),
    .B(net196),
    .C(net173),
    .D(_0197_),
    .X(_0201_));
 sg13g2_xor2_1 _1572_ (.B(_0200_),
    .A(net173),
    .X(_0149_));
 sg13g2_and2_1 _1573_ (.A(net212),
    .B(_0201_),
    .X(_0202_));
 sg13g2_xor2_1 _1574_ (.B(_0201_),
    .A(net212),
    .X(_0150_));
 sg13g2_and4_1 _1575_ (.A(net212),
    .B(net173),
    .C(\top_inst.sndgen_inst.slot_counter[7] ),
    .D(_0200_),
    .X(_0203_));
 sg13g2_xor2_1 _1576_ (.B(_0202_),
    .A(net299),
    .X(_0151_));
 sg13g2_and3_1 _1577_ (.X(_0204_),
    .A(\top_inst.sndgen_inst.slot_counter[8] ),
    .B(\top_inst.sndgen_inst.slot_counter[7] ),
    .C(_0202_));
 sg13g2_xor2_1 _1578_ (.B(_0203_),
    .A(net296),
    .X(_0152_));
 sg13g2_xor2_1 _1579_ (.B(_0204_),
    .A(net92),
    .X(_0153_));
 sg13g2_a21oi_1 _1580_ (.A1(\top_inst.sndgen_inst.slot_counter[9] ),
    .A2(_0204_),
    .Y(_0205_),
    .B1(net46));
 sg13g2_and4_2 _1581_ (.A(net296),
    .B(net46),
    .C(net92),
    .D(_0203_),
    .X(_0206_));
 sg13g2_nor2_1 _1582_ (.A(net47),
    .B(_0206_),
    .Y(_0154_));
 sg13g2_xor2_1 _1583_ (.B(_0206_),
    .A(net354),
    .X(_0155_));
 sg13g2_a21oi_1 _1584_ (.A1(\top_inst.sndgen_inst.bar_counter[0] ),
    .A2(_0206_),
    .Y(_0207_),
    .B1(net304));
 sg13g2_nand3_1 _1585_ (.B(\top_inst.sndgen_inst.bar_counter[0] ),
    .C(_0206_),
    .A(net304),
    .Y(_0208_));
 sg13g2_nor2b_1 _1586_ (.A(net305),
    .B_N(_0208_),
    .Y(_0156_));
 sg13g2_xnor2_1 _1587_ (.Y(_0157_),
    .A(net347),
    .B(_0208_));
 sg13g2_nand4_1 _1588_ (.B(\top_inst.sndgen_inst.bar_counter[0] ),
    .C(\top_inst.sndgen_inst.bar_counter[2] ),
    .A(\top_inst.sndgen_inst.bar_counter[1] ),
    .Y(_0209_),
    .D(_0206_));
 sg13g2_xnor2_1 _1589_ (.Y(_0158_),
    .A(net194),
    .B(_0209_));
 sg13g2_nand2_1 _1590_ (.Y(_0210_),
    .A(net42),
    .B(_0438_));
 sg13g2_o21ai_1 _1591_ (.B1(_0210_),
    .Y(_0159_),
    .A1(_0438_),
    .A2(_0502_));
 sg13g2_nand2_1 _1592_ (.Y(_0211_),
    .A(net137),
    .B(_0438_));
 sg13g2_nand4_1 _1593_ (.B(\top_inst.sndgen_inst.lfsr[5] ),
    .C(_0430_),
    .A(net256),
    .Y(_0212_),
    .D(net226));
 sg13g2_nand2_1 _1594_ (.Y(_0160_),
    .A(_0211_),
    .B(_0212_));
 sg13g2_nor2_2 _1595_ (.A(net221),
    .B(_0439_),
    .Y(_0213_));
 sg13g2_nand3_1 _1596_ (.B(\top_inst.sndgen_inst.bar_counter[3] ),
    .C(_0213_),
    .A(\top_inst.sndgen_inst.bar_counter[2] ),
    .Y(_0214_));
 sg13g2_mux2_1 _1597_ (.A0(\top_inst.sndgen_inst.lfsr[1] ),
    .A1(net131),
    .S(_0214_),
    .X(_0161_));
 sg13g2_mux2_1 _1598_ (.A0(\top_inst.sndgen_inst.lfsr[2] ),
    .A1(net53),
    .S(_0214_),
    .X(_0162_));
 sg13g2_mux2_1 _1599_ (.A0(net362),
    .A1(net359),
    .S(_0214_),
    .X(_0163_));
 sg13g2_mux2_1 _1600_ (.A0(net55),
    .A1(net123),
    .S(_0214_),
    .X(_0164_));
 sg13g2_nor2_1 _1601_ (.A(net253),
    .B(net247),
    .Y(_0215_));
 sg13g2_and2_1 _1602_ (.A(net229),
    .B(_0215_),
    .X(_0216_));
 sg13g2_and2_1 _1603_ (.A(_0432_),
    .B(_0215_),
    .X(_0217_));
 sg13g2_a22oi_1 _1604_ (.Y(_0218_),
    .B1(_0217_),
    .B2(net168),
    .A2(_0216_),
    .A1(\top_inst.sndgen_inst.rom_addr[0] ));
 sg13g2_o21ai_1 _1605_ (.B1(_0218_),
    .Y(_0165_),
    .A1(_0253_),
    .A2(_0215_));
 sg13g2_a22oi_1 _1606_ (.Y(_0219_),
    .B1(_0217_),
    .B2(net171),
    .A2(_0216_),
    .A1(net313));
 sg13g2_o21ai_1 _1607_ (.B1(_0219_),
    .Y(_0166_),
    .A1(_0254_),
    .A2(_0215_));
 sg13g2_nand2b_1 _1608_ (.Y(_0220_),
    .B(net106),
    .A_N(net253));
 sg13g2_nand2_1 _1609_ (.Y(_0221_),
    .A(net250),
    .B(net137));
 sg13g2_a21oi_1 _1610_ (.A1(_0220_),
    .A2(_0221_),
    .Y(_0222_),
    .B1(net247));
 sg13g2_a21oi_1 _1611_ (.A1(net247),
    .A2(net42),
    .Y(_0223_),
    .B1(_0222_));
 sg13g2_nand2_1 _1612_ (.Y(_0224_),
    .A(net336),
    .B(_0216_));
 sg13g2_o21ai_1 _1613_ (.B1(_0224_),
    .Y(_0167_),
    .A1(_0216_),
    .A2(_0223_));
 sg13g2_a22oi_1 _1614_ (.Y(_0225_),
    .B1(_0216_),
    .B2(net152),
    .A2(net137),
    .A1(net247));
 sg13g2_inv_1 _1615_ (.Y(_0168_),
    .A(_0225_));
 sg13g2_nor4_1 _1616_ (.A(\top_inst.sndgen_inst.lfsr[3] ),
    .B(\top_inst.sndgen_inst.lfsr[2] ),
    .C(\top_inst.sndgen_inst.lfsr[1] ),
    .D(_0214_),
    .Y(_0226_));
 sg13g2_a21oi_1 _1617_ (.A1(_0236_),
    .A2(_0214_),
    .Y(_0169_),
    .B1(_0226_));
 sg13g2_mux2_1 _1618_ (.A0(net256),
    .A1(net300),
    .S(net221),
    .X(_0170_));
 sg13g2_nand2_1 _1619_ (.Y(_0227_),
    .A(net64),
    .B(net221));
 sg13g2_nand2b_1 _1620_ (.Y(_0228_),
    .B(_0007_),
    .A_N(\top_inst.sndgen_inst.lfsr[5] ));
 sg13g2_nand3_1 _1621_ (.B(\top_inst.sndgen_inst.lfsr[3] ),
    .C(_0228_),
    .A(net256),
    .Y(_0229_));
 sg13g2_o21ai_1 _1622_ (.B1(_0227_),
    .Y(_0171_),
    .A1(net221),
    .A2(_0229_));
 sg13g2_or2_1 _1623_ (.X(_0172_),
    .B(_0213_),
    .A(net168));
 sg13g2_xnor2_1 _1624_ (.Y(_0230_),
    .A(\top_inst.sndgen_inst.bar_counter[2] ),
    .B(\top_inst.sndgen_inst.bar_counter[3] ));
 sg13g2_nor2_1 _1625_ (.A(net171),
    .B(_0213_),
    .Y(_0231_));
 sg13g2_a21oi_1 _1626_ (.A1(_0213_),
    .A2(_0230_),
    .Y(_0173_),
    .B1(_0231_));
 sg13g2_mux2_1 _1627_ (.A0(net106),
    .A1(\top_inst.sndgen_inst.bar_counter[3] ),
    .S(_0213_),
    .X(_0174_));
 sg13g2_nor2_1 _1628_ (.A(net127),
    .B(net246),
    .Y(_0232_));
 sg13g2_a21oi_1 _1629_ (.A1(net246),
    .A2(_0531_),
    .Y(_0175_),
    .B1(net128));
 sg13g2_nor2_1 _1630_ (.A(net204),
    .B(net246),
    .Y(_0233_));
 sg13g2_a21oi_1 _1631_ (.A1(net246),
    .A2(_0533_),
    .Y(_0176_),
    .B1(net205));
 sg13g2_nor2_1 _1632_ (.A(net218),
    .B(net246),
    .Y(_0234_));
 sg13g2_a21oi_1 _1633_ (.A1(net246),
    .A2(_0536_),
    .Y(_0177_),
    .B1(net292));
 sg13g2_nor2_1 _1634_ (.A(net307),
    .B(net246),
    .Y(_0235_));
 sg13g2_a21oi_1 _1635_ (.A1(net246),
    .A2(_0539_),
    .Y(_0178_),
    .B1(net308));
 sg13g2_dfrbp_1 _1636_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net277),
    .D(net182),
    .Q_N(_0888_),
    .Q(\top_inst.sndgen_inst.p_c4[4] ));
 sg13g2_dfrbp_1 _1637_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net277),
    .D(net149),
    .Q_N(_0887_),
    .Q(\top_inst.sndgen_inst.p_c4[5] ));
 sg13g2_dfrbp_1 _1638_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net280),
    .D(net188),
    .Q_N(_0886_),
    .Q(\top_inst.sndgen_inst.p_c4[6] ));
 sg13g2_dfrbp_1 _1639_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net280),
    .D(net160),
    .Q_N(_0885_),
    .Q(\top_inst.sndgen_inst.p_c4[7] ));
 sg13g2_dfrbp_1 _1640_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net282),
    .D(net351),
    .Q_N(_0884_),
    .Q(\top_inst.sndgen_inst.p_c4[10] ));
 sg13g2_dfrbp_1 _1641_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net271),
    .D(net333),
    .Q_N(_0883_),
    .Q(\top_inst.sndgen_inst.c1[0] ));
 sg13g2_dfrbp_1 _1642_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net271),
    .D(net22),
    .Q_N(\top_inst.sndgen_inst.c1[1] ),
    .Q(_0018_));
 sg13g2_dfrbp_1 _1643_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net275),
    .D(net67),
    .Q_N(_0001_),
    .Q(\top_inst.vga_inst.y[0] ));
 sg13g2_dfrbp_1 _1644_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net275),
    .D(net371),
    .Q_N(_0882_),
    .Q(\top_inst.vga_inst.y[1] ));
 sg13g2_dfrbp_1 _1645_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net275),
    .D(_0030_),
    .Q_N(_0881_),
    .Q(\top_inst.vga_inst.y[2] ));
 sg13g2_dfrbp_1 _1646_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net275),
    .D(_0031_),
    .Q_N(_0880_),
    .Q(\top_inst.vga_inst.bg[0] ));
 sg13g2_dfrbp_1 _1647_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net275),
    .D(net367),
    .Q_N(_0003_),
    .Q(\top_inst.vga_inst.bg[1] ));
 sg13g2_dfrbp_1 _1648_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net274),
    .D(net324),
    .Q_N(_0002_),
    .Q(\top_inst.vga_inst.bg[4] ));
 sg13g2_dfrbp_1 _1649_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net284),
    .D(net361),
    .Q_N(_0004_),
    .Q(\top_inst.vga_inst.bg[5] ));
 sg13g2_dfrbp_1 _1650_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net284),
    .D(net329),
    .Q_N(_0879_),
    .Q(\top_inst.vga_inst.y[7] ));
 sg13g2_dfrbp_1 _1651_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net284),
    .D(net356),
    .Q_N(_0878_),
    .Q(\top_inst.vga_inst.y[8] ));
 sg13g2_dfrbp_1 _1652_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net284),
    .D(_0037_),
    .Q_N(_0877_),
    .Q(\top_inst.vga_inst.y[9] ));
 sg13g2_dfrbp_1 _1653_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net272),
    .D(_0038_),
    .Q_N(_0876_),
    .Q(\top_inst.vga_inst.x[0] ));
 sg13g2_dfrbp_1 _1654_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net272),
    .D(_0039_),
    .Q_N(_0875_),
    .Q(\top_inst.vga_inst.x[1] ));
 sg13g2_dfrbp_1 _1655_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net272),
    .D(net192),
    .Q_N(_0874_),
    .Q(\top_inst.vga_inst.x[2] ));
 sg13g2_dfrbp_1 _1656_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net272),
    .D(net79),
    .Q_N(_0873_),
    .Q(\top_inst.vga_inst.x[3] ));
 sg13g2_dfrbp_1 _1657_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net273),
    .D(_0042_),
    .Q_N(_0872_),
    .Q(\top_inst.vga_inst.x[4] ));
 sg13g2_dfrbp_1 _1658_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net272),
    .D(_0043_),
    .Q_N(_0871_),
    .Q(\top_inst.vga_inst.x[5] ));
 sg13g2_dfrbp_1 _1659_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net275),
    .D(net374),
    .Q_N(_0870_),
    .Q(\top_inst.vga_inst.x[6] ));
 sg13g2_dfrbp_1 _1660_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net275),
    .D(_0045_),
    .Q_N(_0869_),
    .Q(\top_inst.vga_inst.x[7] ));
 sg13g2_dfrbp_1 _1661_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net273),
    .D(_0046_),
    .Q_N(_0868_),
    .Q(\top_inst.vga_inst.x[8] ));
 sg13g2_dfrbp_1 _1662_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net273),
    .D(_0047_),
    .Q_N(_0867_),
    .Q(\top_inst.vga_inst.x[9] ));
 sg13g2_dfrbp_1 _1663_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net288),
    .D(net33),
    .Q_N(_0866_),
    .Q(\top_inst.vga_inst.xmin[0] ));
 sg13g2_dfrbp_1 _1664_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net288),
    .D(net316),
    .Q_N(_0865_),
    .Q(\top_inst.vga_inst.xmin[1] ));
 sg13g2_dfrbp_1 _1665_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net287),
    .D(net81),
    .Q_N(_0864_),
    .Q(\top_inst.vga_inst.xmin[2] ));
 sg13g2_dfrbp_1 _1666_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net285),
    .D(net190),
    .Q_N(_0863_),
    .Q(\top_inst.vga_inst.xmin[3] ));
 sg13g2_dfrbp_1 _1667_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net270),
    .D(net31),
    .Q_N(\top_inst.sndgen_inst.lfsr[0] ),
    .Q(_0019_));
 sg13g2_dfrbp_1 _1668_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net270),
    .D(net18),
    .Q_N(_0862_),
    .Q(\top_inst.sndgen_inst.lfsr[1] ));
 sg13g2_dfrbp_1 _1669_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net271),
    .D(_0054_),
    .Q_N(_0861_),
    .Q(\top_inst.sndgen_inst.lfsr[2] ));
 sg13g2_dfrbp_1 _1670_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net270),
    .D(net112),
    .Q_N(_0860_),
    .Q(\top_inst.sndgen_inst.lfsr[3] ));
 sg13g2_dfrbp_1 _1671_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net274),
    .D(net56),
    .Q_N(_0859_),
    .Q(\top_inst.sndgen_inst.lfsr[4] ));
 sg13g2_dfrbp_1 _1672_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net274),
    .D(_0057_),
    .Q_N(_0858_),
    .Q(\top_inst.sndgen_inst.lfsr[5] ));
 sg13g2_dfrbp_1 _1673_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net271),
    .D(net52),
    .Q_N(_0857_),
    .Q(\top_inst.sndgen_inst.lfsr[6] ));
 sg13g2_dfrbp_1 _1674_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net271),
    .D(_0059_),
    .Q_N(_0007_),
    .Q(\top_inst.sndgen_inst.lfsr[7] ));
 sg13g2_dfrbp_1 _1675_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net288),
    .D(net176),
    .Q_N(_0856_),
    .Q(\top_inst.vga_inst.xmax[0] ));
 sg13g2_dfrbp_1 _1676_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net287),
    .D(net217),
    .Q_N(_0855_),
    .Q(\top_inst.vga_inst.xmax[1] ));
 sg13g2_dfrbp_1 _1677_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net287),
    .D(net118),
    .Q_N(_0854_),
    .Q(\top_inst.vga_inst.xmax[2] ));
 sg13g2_dfrbp_1 _1678_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net285),
    .D(net72),
    .Q_N(_0853_),
    .Q(\top_inst.vga_inst.xmax[3] ));
 sg13g2_dfrbp_1 _1679_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net286),
    .D(_0064_),
    .Q_N(_0852_),
    .Q(\top_inst.vga_inst.sx1[0] ));
 sg13g2_dfrbp_1 _1680_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net286),
    .D(net353),
    .Q_N(_0851_),
    .Q(\top_inst.vga_inst.sx1[1] ));
 sg13g2_dfrbp_1 _1681_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net286),
    .D(_0066_),
    .Q_N(_0850_),
    .Q(\top_inst.vga_inst.sx1[2] ));
 sg13g2_dfrbp_1 _1682_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net284),
    .D(_0067_),
    .Q_N(_0849_),
    .Q(\top_inst.vga_inst.sx1[3] ));
 sg13g2_dfrbp_1 _1683_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net285),
    .D(net63),
    .Q_N(_0848_),
    .Q(\top_inst.vga_inst.x1[0] ));
 sg13g2_dfrbp_1 _1684_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net285),
    .D(net29),
    .Q_N(_0847_),
    .Q(\top_inst.vga_inst.x1[1] ));
 sg13g2_dfrbp_1 _1685_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net287),
    .D(net141),
    .Q_N(_0846_),
    .Q(\top_inst.vga_inst.x1[2] ));
 sg13g2_dfrbp_1 _1686_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net287),
    .D(net295),
    .Q_N(_0845_),
    .Q(\top_inst.vga_inst.x1[3] ));
 sg13g2_dfrbp_1 _1687_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net287),
    .D(_0072_),
    .Q_N(_0844_),
    .Q(\top_inst.vga_inst.x1[4] ));
 sg13g2_dfrbp_1 _1688_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net288),
    .D(_0073_),
    .Q_N(_0843_),
    .Q(\top_inst.vga_inst.x1[5] ));
 sg13g2_dfrbp_1 _1689_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net287),
    .D(_0074_),
    .Q_N(_0842_),
    .Q(\top_inst.vga_inst.x1[6] ));
 sg13g2_dfrbp_1 _1690_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net287),
    .D(_0075_),
    .Q_N(_0841_),
    .Q(\top_inst.vga_inst.x1[7] ));
 sg13g2_dfrbp_1 _1691_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net289),
    .D(_0076_),
    .Q_N(_0840_),
    .Q(\top_inst.vga_inst.sr1[0] ));
 sg13g2_dfrbp_1 _1692_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net289),
    .D(_0077_),
    .Q_N(_0839_),
    .Q(\top_inst.vga_inst.sr1[1] ));
 sg13g2_dfrbp_1 _1693_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net289),
    .D(net146),
    .Q_N(_0838_),
    .Q(\top_inst.vga_inst.sr1[2] ));
 sg13g2_dfrbp_1 _1694_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net285),
    .D(net322),
    .Q_N(_0837_),
    .Q(\top_inst.vga_inst.sr1[3] ));
 sg13g2_dfrbp_1 _1695_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net262),
    .D(net61),
    .Q_N(_0836_),
    .Q(\top_inst.sndgen_inst.p_c3[0] ));
 sg13g2_dfrbp_1 _1696_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net265),
    .D(net126),
    .Q_N(_0835_),
    .Q(\top_inst.sndgen_inst.p_c3[1] ));
 sg13g2_dfrbp_1 _1697_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net265),
    .D(_0082_),
    .Q_N(_0834_),
    .Q(\top_inst.sndgen_inst.p_c3[2] ));
 sg13g2_dfrbp_1 _1698_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net266),
    .D(_0083_),
    .Q_N(_0833_),
    .Q(\top_inst.sndgen_inst.p_c3[3] ));
 sg13g2_dfrbp_1 _1699_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net266),
    .D(net170),
    .Q_N(_0832_),
    .Q(\top_inst.sndgen_inst.p_c3[4] ));
 sg13g2_dfrbp_1 _1700_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net277),
    .D(net105),
    .Q_N(_0831_),
    .Q(\top_inst.sndgen_inst.p_c3[5] ));
 sg13g2_dfrbp_1 _1701_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net279),
    .D(net76),
    .Q_N(_0830_),
    .Q(\top_inst.sndgen_inst.p_c3[6] ));
 sg13g2_dfrbp_1 _1702_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net279),
    .D(_0087_),
    .Q_N(_0829_),
    .Q(\top_inst.sndgen_inst.p_c3[7] ));
 sg13g2_dfrbp_1 _1703_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net279),
    .D(_0088_),
    .Q_N(_0828_),
    .Q(\top_inst.sndgen_inst.p_c3[10] ));
 sg13g2_dfrbp_1 _1704_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net286),
    .D(net88),
    .Q_N(_0017_),
    .Q(\top_inst.pwm_inst.cntr[0] ));
 sg13g2_dfrbp_1 _1705_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net284),
    .D(net379),
    .Q_N(_0827_),
    .Q(\top_inst.pwm_inst.cntr[1] ));
 sg13g2_dfrbp_1 _1706_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net284),
    .D(net303),
    .Q_N(_0826_),
    .Q(\top_inst.pwm_inst.cntr[2] ));
 sg13g2_dfrbp_1 _1707_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net284),
    .D(net86),
    .Q_N(_0889_),
    .Q(\top_inst.pwm_inst.cntr[3] ));
 sg13g2_dfrbp_1 _1708_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net280),
    .D(net237),
    .Q_N(_0890_),
    .Q(\top_inst.sndgen_inst.sample_ena_delay[0] ));
 sg13g2_dfrbp_1 _1709_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net267),
    .D(net250),
    .Q_N(_0891_),
    .Q(\top_inst.sndgen_inst.sample_ena_delay[1] ));
 sg13g2_dfrbp_1 _1710_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net277),
    .D(net248),
    .Q_N(_0825_),
    .Q(\top_inst.sndgen_inst.sample_ena_delay[2] ));
 sg13g2_dfrbp_1 _1711_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net267),
    .D(net41),
    .Q_N(_0824_),
    .Q(\top_inst.sndgen_inst.phacc2[0] ));
 sg13g2_dfrbp_1 _1712_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net267),
    .D(net157),
    .Q_N(_0823_),
    .Q(\top_inst.sndgen_inst.phacc2[1] ));
 sg13g2_dfrbp_1 _1713_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net277),
    .D(net136),
    .Q_N(_0822_),
    .Q(\top_inst.sndgen_inst.phacc2[2] ));
 sg13g2_dfrbp_1 _1714_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net278),
    .D(_0096_),
    .Q_N(_0821_),
    .Q(\top_inst.sndgen_inst.phacc2[3] ));
 sg13g2_dfrbp_1 _1715_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net283),
    .D(_0097_),
    .Q_N(_0820_),
    .Q(\top_inst.sndgen_inst.phacc2[4] ));
 sg13g2_dfrbp_1 _1716_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net283),
    .D(_0098_),
    .Q_N(_0819_),
    .Q(\top_inst.sndgen_inst.phacc2[5] ));
 sg13g2_dfrbp_1 _1717_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net283),
    .D(net178),
    .Q_N(_0818_),
    .Q(\top_inst.sndgen_inst.phacc2[6] ));
 sg13g2_dfrbp_1 _1718_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net282),
    .D(net166),
    .Q_N(_0817_),
    .Q(\top_inst.sndgen_inst.phacc2[7] ));
 sg13g2_dfrbp_1 _1719_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net283),
    .D(net35),
    .Q_N(_0010_),
    .Q(\top_inst.sndgen_inst.phacc2[8] ));
 sg13g2_dfrbp_1 _1720_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net283),
    .D(net214),
    .Q_N(_0816_),
    .Q(\top_inst.sndgen_inst.phacc2[9] ));
 sg13g2_dfrbp_1 _1721_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net283),
    .D(_0103_),
    .Q_N(_0815_),
    .Q(\top_inst.sndgen_inst.phacc2[10] ));
 sg13g2_dfrbp_1 _1722_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net282),
    .D(_0104_),
    .Q_N(_0814_),
    .Q(\top_inst.sndgen_inst.phacc2[11] ));
 sg13g2_dfrbp_1 _1723_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net282),
    .D(net144),
    .Q_N(_0813_),
    .Q(\top_inst.sndgen_inst.phacc2[12] ));
 sg13g2_dfrbp_1 _1724_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net282),
    .D(net331),
    .Q_N(_0812_),
    .Q(\top_inst.sndgen_inst.phacc2[13] ));
 sg13g2_dfrbp_1 _1725_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net266),
    .D(net45),
    .Q_N(_0811_),
    .Q(\top_inst.sndgen_inst.p_c2[0] ));
 sg13g2_dfrbp_1 _1726_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net267),
    .D(_0108_),
    .Q_N(_0810_),
    .Q(\top_inst.sndgen_inst.p_c2[1] ));
 sg13g2_dfrbp_1 _1727_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net267),
    .D(_0109_),
    .Q_N(_0809_),
    .Q(\top_inst.sndgen_inst.p_c2[2] ));
 sg13g2_dfrbp_1 _1728_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net278),
    .D(net102),
    .Q_N(_0808_),
    .Q(\top_inst.sndgen_inst.p_c2[3] ));
 sg13g2_dfrbp_1 _1729_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net278),
    .D(net98),
    .Q_N(_0807_),
    .Q(\top_inst.sndgen_inst.p_c2[4] ));
 sg13g2_dfrbp_1 _1730_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net278),
    .D(net320),
    .Q_N(_0806_),
    .Q(\top_inst.sndgen_inst.p_c2[5] ));
 sg13g2_dfrbp_1 _1731_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net283),
    .D(net91),
    .Q_N(_0805_),
    .Q(\top_inst.sndgen_inst.p_c2[6] ));
 sg13g2_dfrbp_1 _1732_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net282),
    .D(net208),
    .Q_N(_0804_),
    .Q(\top_inst.sndgen_inst.p_c2[7] ));
 sg13g2_dfrbp_1 _1733_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net282),
    .D(net345),
    .Q_N(_0803_),
    .Q(\top_inst.sndgen_inst.p_c2[10] ));
 sg13g2_dfrbp_1 _1734_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net262),
    .D(net39),
    .Q_N(_0802_),
    .Q(\top_inst.sndgen_inst.phacc3[0] ));
 sg13g2_dfrbp_1 _1735_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net262),
    .D(_0117_),
    .Q_N(_0801_),
    .Q(\top_inst.sndgen_inst.phacc3[1] ));
 sg13g2_dfrbp_1 _1736_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net262),
    .D(net199),
    .Q_N(_0800_),
    .Q(\top_inst.sndgen_inst.phacc3[2] ));
 sg13g2_dfrbp_1 _1737_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net264),
    .D(_0119_),
    .Q_N(_0799_),
    .Q(\top_inst.sndgen_inst.phacc3[3] ));
 sg13g2_dfrbp_1 _1738_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net266),
    .D(net84),
    .Q_N(_0798_),
    .Q(\top_inst.sndgen_inst.phacc3[4] ));
 sg13g2_dfrbp_1 _1739_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net277),
    .D(_0121_),
    .Q_N(_0797_),
    .Q(\top_inst.sndgen_inst.phacc3[5] ));
 sg13g2_dfrbp_1 _1740_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net279),
    .D(_0122_),
    .Q_N(_0796_),
    .Q(\top_inst.sndgen_inst.phacc3[6] ));
 sg13g2_dfrbp_1 _1741_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net279),
    .D(_0123_),
    .Q_N(_0795_),
    .Q(\top_inst.sndgen_inst.phacc3[7] ));
 sg13g2_dfrbp_1 _1742_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net279),
    .D(net20),
    .Q_N(_0011_),
    .Q(\top_inst.sndgen_inst.phacc3[8] ));
 sg13g2_dfrbp_1 _1743_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net280),
    .D(net114),
    .Q_N(_0794_),
    .Q(\top_inst.sndgen_inst.phacc3[9] ));
 sg13g2_dfrbp_1 _1744_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net286),
    .D(_0126_),
    .Q_N(_0793_),
    .Q(\top_inst.sndgen_inst.phacc3[10] ));
 sg13g2_dfrbp_1 _1745_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net286),
    .D(_0127_),
    .Q_N(_0792_),
    .Q(\top_inst.sndgen_inst.phacc3[11] ));
 sg13g2_dfrbp_1 _1746_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net286),
    .D(_0128_),
    .Q_N(_0791_),
    .Q(\top_inst.sndgen_inst.phacc3[12] ));
 sg13g2_dfrbp_1 _1747_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net274),
    .D(net312),
    .Q_N(_0790_),
    .Q(\top_inst.sndgen_inst.phacc3[13] ));
 sg13g2_dfrbp_1 _1748_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net262),
    .D(net37),
    .Q_N(_0789_),
    .Q(\top_inst.sndgen_inst.phacc4[0] ));
 sg13g2_dfrbp_1 _1749_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net262),
    .D(net201),
    .Q_N(_0788_),
    .Q(\top_inst.sndgen_inst.phacc4[1] ));
 sg13g2_dfrbp_1 _1750_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net266),
    .D(net100),
    .Q_N(_0787_),
    .Q(\top_inst.sndgen_inst.phacc4[2] ));
 sg13g2_dfrbp_1 _1751_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net266),
    .D(net210),
    .Q_N(_0786_),
    .Q(\top_inst.sndgen_inst.phacc4[3] ));
 sg13g2_dfrbp_1 _1752_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net277),
    .D(_0134_),
    .Q_N(_0785_),
    .Q(\top_inst.sndgen_inst.phacc4[4] ));
 sg13g2_dfrbp_1 _1753_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net277),
    .D(_0135_),
    .Q_N(_0784_),
    .Q(\top_inst.sndgen_inst.phacc4[5] ));
 sg13g2_dfrbp_1 _1754_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net279),
    .D(_0136_),
    .Q_N(_0783_),
    .Q(\top_inst.sndgen_inst.phacc4[6] ));
 sg13g2_dfrbp_1 _1755_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net279),
    .D(net163),
    .Q_N(_0782_),
    .Q(\top_inst.sndgen_inst.phacc4[7] ));
 sg13g2_dfrbp_1 _1756_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net282),
    .D(net24),
    .Q_N(_0000_),
    .Q(\top_inst.sndgen_inst.phacc4[8] ));
 sg13g2_dfrbp_1 _1757_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net289),
    .D(net116),
    .Q_N(_0781_),
    .Q(\top_inst.sndgen_inst.phacc4[9] ));
 sg13g2_dfrbp_1 _1758_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net289),
    .D(net70),
    .Q_N(_0780_),
    .Q(\top_inst.sndgen_inst.phacc4[10] ));
 sg13g2_dfrbp_1 _1759_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net289),
    .D(net58),
    .Q_N(_0779_),
    .Q(\top_inst.sndgen_inst.phacc4[11] ));
 sg13g2_dfrbp_1 _1760_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net289),
    .D(_0142_),
    .Q_N(_0778_),
    .Q(\top_inst.sndgen_inst.phacc4[12] ));
 sg13g2_dfrbp_1 _1761_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net286),
    .D(net318),
    .Q_N(_0777_),
    .Q(\top_inst.sndgen_inst.phacc4[13] ));
 sg13g2_dfrbp_1 _1762_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net264),
    .D(net326),
    .Q_N(_0016_),
    .Q(\top_inst.sndgen_inst.slot_counter[0] ));
 sg13g2_dfrbp_1 _1763_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net263),
    .D(net203),
    .Q_N(_0776_),
    .Q(\top_inst.sndgen_inst.slot_counter[1] ));
 sg13g2_dfrbp_1 _1764_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net263),
    .D(net184),
    .Q_N(_0775_),
    .Q(\top_inst.sndgen_inst.slot_counter[2] ));
 sg13g2_dfrbp_1 _1765_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net263),
    .D(net197),
    .Q_N(_0774_),
    .Q(\top_inst.sndgen_inst.slot_counter[3] ));
 sg13g2_dfrbp_1 _1766_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net263),
    .D(net110),
    .Q_N(_0773_),
    .Q(\top_inst.sndgen_inst.slot_counter[4] ));
 sg13g2_dfrbp_1 _1767_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net263),
    .D(net174),
    .Q_N(_0772_),
    .Q(\top_inst.sndgen_inst.slot_counter[5] ));
 sg13g2_dfrbp_1 _1768_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net263),
    .D(_0150_),
    .Q_N(_0771_),
    .Q(\top_inst.sndgen_inst.slot_counter[6] ));
 sg13g2_dfrbp_1 _1769_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net264),
    .D(_0151_),
    .Q_N(_0770_),
    .Q(\top_inst.sndgen_inst.slot_counter[7] ));
 sg13g2_dfrbp_1 _1770_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net264),
    .D(net297),
    .Q_N(_0769_),
    .Q(\top_inst.sndgen_inst.slot_counter[8] ));
 sg13g2_dfrbp_1 _1771_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net263),
    .D(net93),
    .Q_N(_0768_),
    .Q(\top_inst.sndgen_inst.slot_counter[9] ));
 sg13g2_dfrbp_1 _1772_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net263),
    .D(net48),
    .Q_N(_0767_),
    .Q(\top_inst.sndgen_inst.slot_counter[10] ));
 sg13g2_dfrbp_1 _1773_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net270),
    .D(_0155_),
    .Q_N(_0766_),
    .Q(\top_inst.sndgen_inst.bar_counter[0] ));
 sg13g2_dfrbp_1 _1774_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net270),
    .D(net306),
    .Q_N(_0765_),
    .Q(\top_inst.sndgen_inst.bar_counter[1] ));
 sg13g2_dfrbp_1 _1775_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net270),
    .D(net348),
    .Q_N(_0764_),
    .Q(\top_inst.sndgen_inst.bar_counter[2] ));
 sg13g2_dfrbp_1 _1776_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net264),
    .D(net195),
    .Q_N(_0763_),
    .Q(\top_inst.sndgen_inst.bar_counter[3] ));
 sg13g2_dfrbp_1 _1777_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net274),
    .D(net43),
    .Q_N(_0762_),
    .Q(\top_inst.sndgen_inst.c4[2] ));
 sg13g2_dfrbp_1 _1778_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net268),
    .D(net138),
    .Q_N(_0761_),
    .Q(\top_inst.sndgen_inst.c3[2] ));
 sg13g2_dfrbp_1 _1779_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net271),
    .D(net132),
    .Q_N(_0760_),
    .Q(\top_inst.sndgen_inst.mask_1[0] ));
 sg13g2_dfrbp_1 _1780_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net274),
    .D(net54),
    .Q_N(_0008_),
    .Q(\top_inst.sndgen_inst.mask_1[1] ));
 sg13g2_dfrbp_1 _1781_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net274),
    .D(_0163_),
    .Q_N(_0759_),
    .Q(\top_inst.sndgen_inst.mask_1[2] ));
 sg13g2_dfrbp_1 _1782_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net274),
    .D(_0164_),
    .Q_N(_0009_),
    .Q(\top_inst.sndgen_inst.mask_1[3] ));
 sg13g2_dfrbp_1 _1783_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net268),
    .D(net301),
    .Q_N(_0758_),
    .Q(\top_inst.sndgen_inst.rom_addr[0] ));
 sg13g2_dfrbp_1 _1784_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net269),
    .D(_0166_),
    .Q_N(_0757_),
    .Q(\top_inst.sndgen_inst.rom_addr[1] ));
 sg13g2_dfrbp_1 _1785_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net268),
    .D(_0167_),
    .Q_N(_0006_),
    .Q(\top_inst.sndgen_inst.rom_addr[2] ));
 sg13g2_dfrbp_1 _1786_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net268),
    .D(_0168_),
    .Q_N(_0005_),
    .Q(\top_inst.sndgen_inst.rom_addr[3] ));
 sg13g2_dfrbp_1 _1787_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net271),
    .D(net26),
    .Q_N(\top_inst.sndgen_inst.mask_2 ),
    .Q(_0020_));
 sg13g2_dfrbp_1 _1788_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net268),
    .D(_0170_),
    .Q_N(_0756_),
    .Q(\top_inst.sndgen_inst.c3[0] ));
 sg13g2_dfrbp_1 _1789_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net268),
    .D(net65),
    .Q_N(_0892_),
    .Q(\top_inst.sndgen_inst.c3[1] ));
 sg13g2_dfrbp_1 _1790_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net272),
    .D(net16),
    .Q_N(_0747_),
    .Q(\top_inst.sys_presc[0] ));
 sg13g2_dfrbp_1 _1791_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net272),
    .D(_0012_),
    .Q_N(_0893_),
    .Q(\top_inst.sys_presc[1] ));
 sg13g2_dfrbp_1 _1792_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net272),
    .D(_0013_),
    .Q_N(_0894_),
    .Q(\top_inst.sys_presc[2] ));
 sg13g2_dfrbp_1 _1793_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net270),
    .D(net120),
    .Q_N(_0895_),
    .Q(\top_inst.sys_presc[3] ));
 sg13g2_dfrbp_1 _1794_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net270),
    .D(net50),
    .Q_N(_0755_),
    .Q(\top_inst.sys_presc[4] ));
 sg13g2_dfrbp_1 _1795_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net268),
    .D(_0172_),
    .Q_N(_0754_),
    .Q(\top_inst.sndgen_inst.c2[0] ));
 sg13g2_dfrbp_1 _1796_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net264),
    .D(net172),
    .Q_N(_0753_),
    .Q(\top_inst.sndgen_inst.c2[1] ));
 sg13g2_dfrbp_1 _1797_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net268),
    .D(net107),
    .Q_N(_0752_),
    .Q(\top_inst.sndgen_inst.c2[2] ));
 sg13g2_dfrbp_1 _1798_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net262),
    .D(net129),
    .Q_N(_0751_),
    .Q(\top_inst.sndgen_inst.p_c4[0] ));
 sg13g2_dfrbp_1 _1799_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net262),
    .D(net206),
    .Q_N(_0750_),
    .Q(\top_inst.sndgen_inst.p_c4[1] ));
 sg13g2_dfrbp_1 _1800_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net266),
    .D(net293),
    .Q_N(_0749_),
    .Q(\top_inst.sndgen_inst.p_c4[2] ));
 sg13g2_dfrbp_1 _1801_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net266),
    .D(net309),
    .Q_N(_0748_),
    .Q(\top_inst.sndgen_inst.p_c4[3] ));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_cfib_demo_2 (.L_LO(net2));
 sg13g2_tielo tt_um_cfib_demo_3 (.L_LO(net3));
 sg13g2_tielo tt_um_cfib_demo_4 (.L_LO(net4));
 sg13g2_tielo tt_um_cfib_demo_5 (.L_LO(net5));
 sg13g2_tielo tt_um_cfib_demo_6 (.L_LO(net6));
 sg13g2_tielo tt_um_cfib_demo_7 (.L_LO(net7));
 sg13g2_tielo tt_um_cfib_demo_8 (.L_LO(net8));
 sg13g2_tielo tt_um_cfib_demo_9 (.L_LO(net9));
 sg13g2_tielo tt_um_cfib_demo_10 (.L_LO(net10));
 sg13g2_tielo tt_um_cfib_demo_11 (.L_LO(net11));
 sg13g2_tielo tt_um_cfib_demo_12 (.L_LO(net12));
 sg13g2_tielo tt_um_cfib_demo_13 (.L_LO(net13));
 sg13g2_tielo tt_um_cfib_demo_14 (.L_LO(net14));
 sg13g2_tiehi tt_um_cfib_demo_15 (.L_HI(net15));
 sg13g2_buf_1 _1817_ (.A(pwm),
    .X(uio_out[7]));
 sg13g2_buf_1 _1818_ (.A(\top_inst.vga_inst.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _1819_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout219 (.A(_0488_),
    .X(net219));
 sg13g2_buf_1 fanout220 (.A(_0488_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_0438_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(net223),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_0482_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_0481_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(net226),
    .X(net225));
 sg13g2_buf_4 fanout226 (.X(net226),
    .A(_0437_));
 sg13g2_buf_2 fanout227 (.A(_0434_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(net229),
    .X(net228));
 sg13g2_buf_4 fanout229 (.X(net229),
    .A(_0436_));
 sg13g2_buf_2 fanout230 (.A(net232),
    .X(net230));
 sg13g2_buf_1 fanout231 (.A(net232),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(net233),
    .X(net232));
 sg13g2_buf_4 fanout233 (.X(net233),
    .A(_0435_));
 sg13g2_buf_2 fanout234 (.A(net235),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(net236),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_0435_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(net239),
    .X(net237));
 sg13g2_buf_1 fanout238 (.A(net239),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(\top_inst.sample_ena ),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(net241),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(net242),
    .X(net241));
 sg13g2_buf_4 fanout242 (.X(net242),
    .A(\top_inst.sys_presc[0] ));
 sg13g2_buf_2 fanout243 (.A(net244),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(\top_inst.sndgen_inst.p_c2[10] ),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(\top_inst.sndgen_inst.sample_ena_delay[2] ),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(\top_inst.sndgen_inst.sample_ena_delay[2] ),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(net248),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(net150),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(net150),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(net253),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(net253),
    .X(net251));
 sg13g2_buf_1 fanout252 (.A(net253),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(net383),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(net255),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(net346),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(net130),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(net376),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(net385),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(net382),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(net261),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(net349),
    .X(net261));
 sg13g2_buf_4 fanout262 (.X(net262),
    .A(net265));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(net264));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(net265));
 sg13g2_buf_2 fanout265 (.A(net276),
    .X(net265));
 sg13g2_buf_4 fanout266 (.X(net266),
    .A(net269));
 sg13g2_buf_2 fanout267 (.A(net269),
    .X(net267));
 sg13g2_buf_4 fanout268 (.X(net268),
    .A(net269));
 sg13g2_buf_2 fanout269 (.A(net276),
    .X(net269));
 sg13g2_buf_4 fanout270 (.X(net270),
    .A(net273));
 sg13g2_buf_4 fanout271 (.X(net271),
    .A(net273));
 sg13g2_buf_4 fanout272 (.X(net272),
    .A(net273));
 sg13g2_buf_2 fanout273 (.A(net276),
    .X(net273));
 sg13g2_buf_4 fanout274 (.X(net274),
    .A(net276));
 sg13g2_buf_4 fanout275 (.X(net275),
    .A(net276));
 sg13g2_buf_2 fanout276 (.A(net291),
    .X(net276));
 sg13g2_buf_4 fanout277 (.X(net277),
    .A(net281));
 sg13g2_buf_2 fanout278 (.A(net281),
    .X(net278));
 sg13g2_buf_4 fanout279 (.X(net279),
    .A(net281));
 sg13g2_buf_2 fanout280 (.A(net281),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(net291),
    .X(net281));
 sg13g2_buf_4 fanout282 (.X(net282),
    .A(net283));
 sg13g2_buf_4 fanout283 (.X(net283),
    .A(net291));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(net290));
 sg13g2_buf_2 fanout285 (.A(net290),
    .X(net285));
 sg13g2_buf_4 fanout286 (.X(net286),
    .A(net290));
 sg13g2_buf_4 fanout287 (.X(net287),
    .A(net290));
 sg13g2_buf_2 fanout288 (.A(net289),
    .X(net288));
 sg13g2_buf_4 fanout289 (.X(net289),
    .A(net290));
 sg13g2_buf_2 fanout290 (.A(net291),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(rst_n),
    .X(net291));
 sg13g2_tielo tt_um_cfib_demo_1 (.L_LO(net1));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_25__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0747_),
    .X(net16));
 sg13g2_dlygate4sd3_1 hold2 (.A(\top_inst.sndgen_inst.lfsr[0] ),
    .X(net17));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0053_),
    .X(net18));
 sg13g2_dlygate4sd3_1 hold4 (.A(\top_inst.sndgen_inst.phacc3[8] ),
    .X(net19));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0124_),
    .X(net20));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0018_),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0027_),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold8 (.A(\top_inst.sndgen_inst.phacc4[8] ),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0138_),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0020_),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0169_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold12 (.A(\top_inst.vga_inst.x1[1] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0517_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0069_),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0019_),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0052_),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold17 (.A(\top_inst.vga_inst.xmin[0] ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0048_),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold19 (.A(\top_inst.sndgen_inst.phacc2[8] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0101_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold21 (.A(\top_inst.sndgen_inst.phacc4[0] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0130_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold23 (.A(\top_inst.sndgen_inst.phacc3[0] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0116_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold25 (.A(\top_inst.sndgen_inst.phacc2[0] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0093_),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold27 (.A(\top_inst.sndgen_inst.c4[2] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0159_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold29 (.A(\top_inst.sndgen_inst.p_c2[0] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0107_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold31 (.A(\top_inst.sndgen_inst.slot_counter[10] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0205_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0154_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold34 (.A(\top_inst.sys_presc[4] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0015_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold36 (.A(\top_inst.sndgen_inst.lfsr[6] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0058_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold38 (.A(\top_inst.sndgen_inst.mask_1[1] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0162_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold40 (.A(\top_inst.sndgen_inst.lfsr[4] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0056_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold42 (.A(\top_inst.sndgen_inst.phacc4[11] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0141_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold44 (.A(\top_inst.sndgen_inst.p_c3[0] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0532_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0080_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold47 (.A(\top_inst.vga_inst.x1[0] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0068_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold49 (.A(\top_inst.sndgen_inst.c3[1] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0171_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0001_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0028_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold53 (.A(\top_inst.sndgen_inst.phacc3[11] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold54 (.A(\top_inst.sndgen_inst.phacc4[10] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0140_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold56 (.A(\top_inst.vga_inst.xmax[3] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0063_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold58 (.A(\top_inst.sndgen_inst.p_c3[7] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold59 (.A(\top_inst.sndgen_inst.p_c3[6] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0543_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0086_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold62 (.A(\top_inst.sndgen_inst.p_c2[2] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold63 (.A(\top_inst.vga_inst.x[3] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0041_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold65 (.A(\top_inst.vga_inst.xmin[2] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0050_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold67 (.A(\top_inst.sndgen_inst.p_c2[1] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold68 (.A(\top_inst.sndgen_inst.phacc3[4] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0120_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold70 (.A(\top_inst.pwm_inst.cntr[3] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0092_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0017_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0089_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold74 (.A(\top_inst.sndgen_inst.p_c2[6] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0624_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0113_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold77 (.A(\top_inst.sndgen_inst.slot_counter[9] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0153_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold79 (.A(\top_inst.sndgen_inst.phacc4[5] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold80 (.A(\top_inst.sndgen_inst.phacc3[10] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold81 (.A(\top_inst.sndgen_inst.phacc3[7] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold82 (.A(\top_inst.sndgen_inst.p_c2[4] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0111_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold84 (.A(\top_inst.sndgen_inst.phacc4[2] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0132_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold86 (.A(\top_inst.sndgen_inst.p_c2[3] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0110_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold88 (.A(\top_inst.sndgen_inst.p_c3[5] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0542_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0085_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold91 (.A(\top_inst.sndgen_inst.c2[2] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0174_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold93 (.A(\top_inst.sndgen_inst.slot_counter[4] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0199_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0148_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold96 (.A(\top_inst.sndgen_inst.lfsr[2] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0055_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold98 (.A(\top_inst.sndgen_inst.phacc3[9] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0125_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold100 (.A(\top_inst.sndgen_inst.phacc4[9] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0139_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold102 (.A(\top_inst.vga_inst.xmax[2] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0062_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold104 (.A(\top_inst.sys_presc[3] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0014_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold106 (.A(\top_inst.sndgen_inst.phacc3[5] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold107 (.A(\top_inst.sys_presc[1] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold108 (.A(\top_inst.sndgen_inst.mask_1[3] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold109 (.A(\top_inst.sndgen_inst.p_c3[1] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0534_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0081_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold112 (.A(\top_inst.sndgen_inst.p_c4[0] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0232_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0175_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold115 (.A(\top_inst.sndgen_inst.lfsr[7] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold116 (.A(\top_inst.sndgen_inst.mask_1[0] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0161_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold118 (.A(\top_inst.sndgen_inst.phacc3[3] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold119 (.A(\top_inst.sndgen_inst.phacc2[2] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0556_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0095_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold122 (.A(\top_inst.sndgen_inst.c3[2] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0160_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold124 (.A(\top_inst.vga_inst.x1[2] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0519_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0070_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold127 (.A(\top_inst.sndgen_inst.phacc2[12] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0605_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0105_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold130 (.A(\top_inst.vga_inst.sr1[2] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0078_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold132 (.A(\top_inst.sndgen_inst.p_c4[5] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0416_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0022_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold135 (.A(\top_inst.sndgen_inst.sample_ena_delay[1] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold136 (.A(\top_inst.sndgen_inst.phacc3[1] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold137 (.A(\top_inst.sndgen_inst.rom_addr[3] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold138 (.A(\top_inst.sndgen_inst.p_c3[2] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold139 (.A(\top_inst.sndgen_inst.phacc2[4] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold140 (.A(\top_inst.sndgen_inst.phacc2[1] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0551_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0094_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold143 (.A(\top_inst.sndgen_inst.p_c4[7] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0423_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0024_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold146 (.A(\top_inst.sndgen_inst.p_c3[3] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold147 (.A(\top_inst.sndgen_inst.phacc4[7] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0137_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold149 (.A(\top_inst.sndgen_inst.phacc4[6] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold150 (.A(\top_inst.sndgen_inst.phacc2[7] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0100_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold152 (.A(\top_inst.sndgen_inst.phacc2[11] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold153 (.A(\top_inst.sndgen_inst.c2[0] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold154 (.A(\top_inst.sndgen_inst.p_c3[4] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0084_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold156 (.A(\top_inst.sndgen_inst.c2[1] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0173_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold158 (.A(\top_inst.sndgen_inst.slot_counter[5] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0149_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold160 (.A(\top_inst.vga_inst.sr1[0] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0060_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold162 (.A(\top_inst.sndgen_inst.phacc2[6] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0099_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold164 (.A(\top_inst.sndgen_inst.phacc2[3] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold165 (.A(\top_inst.sndgen_inst.p_c4[4] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0410_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0021_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold168 (.A(\top_inst.sndgen_inst.slot_counter[2] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0146_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold170 (.A(\top_inst.sndgen_inst.phacc3[6] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold171 (.A(\top_inst.sndgen_inst.p_c4[6] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0420_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0023_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold174 (.A(\top_inst.vga_inst.xmin[3] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0051_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold176 (.A(\top_inst.vga_inst.x[2] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0040_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold178 (.A(\top_inst.sndgen_inst.lfsr[1] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold179 (.A(\top_inst.sndgen_inst.bar_counter[3] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0158_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold181 (.A(\top_inst.sndgen_inst.slot_counter[3] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0147_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold183 (.A(\top_inst.sndgen_inst.phacc3[2] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0118_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold185 (.A(\top_inst.sndgen_inst.phacc4[1] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0131_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold187 (.A(\top_inst.sndgen_inst.slot_counter[1] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0145_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold189 (.A(\top_inst.sndgen_inst.p_c4[1] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0233_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0176_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold192 (.A(\top_inst.sndgen_inst.p_c2[7] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0114_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold194 (.A(\top_inst.sndgen_inst.phacc4[3] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0133_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold196 (.A(\top_inst.sndgen_inst.phacc4[4] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold197 (.A(\top_inst.sndgen_inst.slot_counter[6] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold198 (.A(\top_inst.sndgen_inst.phacc2[9] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0102_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold200 (.A(\top_inst.vga_inst.sx1[2] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold201 (.A(\top_inst.vga_inst.xmax[1] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0061_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold203 (.A(\top_inst.sndgen_inst.p_c4[2] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0234_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0177_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold206 (.A(\top_inst.vga_inst.x1[3] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0071_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold208 (.A(\top_inst.sndgen_inst.slot_counter[8] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0152_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold210 (.A(\top_inst.sndgen_inst.phacc3[12] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold211 (.A(\top_inst.sndgen_inst.slot_counter[7] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold212 (.A(\top_inst.sndgen_inst.c3[0] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0165_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold214 (.A(\top_inst.pwm_inst.cntr[2] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0091_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold216 (.A(\top_inst.sndgen_inst.bar_counter[1] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0207_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0156_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold219 (.A(\top_inst.sndgen_inst.p_c4[3] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0235_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0178_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold222 (.A(\top_inst.vga_inst.sx1[0] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold223 (.A(\top_inst.sndgen_inst.phacc3[13] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0129_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold225 (.A(\top_inst.sndgen_inst.rom_addr[1] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold226 (.A(\top_inst.sndgen_inst.lfsr[5] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold227 (.A(\top_inst.vga_inst.xmin[1] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0049_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold229 (.A(\top_inst.sndgen_inst.phacc4[13] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0143_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold231 (.A(\top_inst.sndgen_inst.p_c2[5] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0112_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold233 (.A(\top_inst.vga_inst.sr1[3] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0079_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0003_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0033_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold237 (.A(\top_inst.sndgen_inst.slot_counter[0] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0144_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold239 (.A(\top_inst.vga_inst.y[7] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0467_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0035_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold242 (.A(\top_inst.sndgen_inst.phacc2[13] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0106_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold244 (.A(\top_inst.sndgen_inst.c1[0] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0026_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold246 (.A(\top_inst.sndgen_inst.phacc2[5] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold247 (.A(\top_inst.sndgen_inst.phacc4[12] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold248 (.A(\top_inst.sndgen_inst.rom_addr[2] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold249 (.A(\top_inst.vga_inst.x[0] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold250 (.A(\top_inst.sndgen_inst.phacc2[10] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold251 (.A(\top_inst.vga_inst.sx1[3] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold252 (.A(\top_inst.vga_inst.x1[4] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold253 (.A(\top_inst.vga_inst.x[7] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0475_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0005_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0424_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0115_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold258 (.A(\top_inst.sndgen_inst.p_c3[10] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold259 (.A(\top_inst.sndgen_inst.bar_counter[2] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0157_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold261 (.A(\top_inst.sndgen_inst.p_c4[10] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0425_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0025_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold264 (.A(\top_inst.vga_inst.sx1[1] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold265 (.A(_0065_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold266 (.A(\top_inst.sndgen_inst.bar_counter[0] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold267 (.A(\top_inst.vga_inst.y[8] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0036_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold269 (.A(\top_inst.vga_inst.x1[6] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0527_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold271 (.A(\top_inst.sndgen_inst.mask_1[2] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold272 (.A(\top_inst.vga_inst.bg[5] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0034_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold274 (.A(\top_inst.sndgen_inst.lfsr[3] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold275 (.A(\top_inst.vga_inst.sr1[1] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold276 (.A(\top_inst.vga_inst.x1[5] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold277 (.A(\top_inst.vga_inst.y[2] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold278 (.A(\top_inst.vga_inst.bg[1] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0032_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold280 (.A(\top_inst.vga_inst.x[5] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0472_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold282 (.A(\top_inst.vga_inst.y[1] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0029_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold284 (.A(\top_inst.vga_inst.bg[0] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold285 (.A(\top_inst.vga_inst.x[6] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0044_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold287 (.A(\top_inst.vga_inst.x1[7] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold288 (.A(\top_inst.vga_inst.x[9] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold289 (.A(\top_inst.pwm_inst.cntr[1] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0548_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0090_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold292 (.A(\top_inst.vga_inst.x[1] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold293 (.A(\top_inst.sys_presc[2] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold294 (.A(\top_inst.vga_inst.x[4] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold295 (.A(\top_inst.sndgen_inst.sample_ena_delay[0] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold296 (.A(\top_inst.vga_inst.y[9] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold297 (.A(\top_inst.vga_inst.x[8] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold298 (.A(\top_inst.sndgen_inst.rom_addr[2] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold299 (.A(\top_inst.sndgen_inst.bar_counter[1] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold300 (.A(\top_inst.sndgen_inst.p_c3[2] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0634_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0642_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold303 (.A(\top_inst.sndgen_inst.phacc3[10] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold304 (.A(\top_inst.sndgen_inst.phacc2[3] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold305 (.A(\top_inst.sndgen_inst.phacc3[9] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold306 (.A(\top_inst.vga_inst.y[1] ),
    .X(net394));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_4 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_274 ();
 sg13g2_decap_8 FILLER_1_281 ();
 sg13g2_decap_8 FILLER_1_288 ();
 sg13g2_decap_8 FILLER_1_295 ();
 sg13g2_decap_8 FILLER_1_302 ();
 sg13g2_decap_8 FILLER_1_309 ();
 sg13g2_decap_8 FILLER_1_316 ();
 sg13g2_decap_8 FILLER_1_323 ();
 sg13g2_decap_8 FILLER_1_330 ();
 sg13g2_decap_8 FILLER_1_337 ();
 sg13g2_decap_8 FILLER_1_344 ();
 sg13g2_decap_8 FILLER_1_351 ();
 sg13g2_decap_8 FILLER_1_358 ();
 sg13g2_decap_8 FILLER_1_365 ();
 sg13g2_decap_8 FILLER_1_372 ();
 sg13g2_decap_8 FILLER_1_379 ();
 sg13g2_decap_8 FILLER_1_386 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_4 FILLER_2_49 ();
 sg13g2_fill_1 FILLER_2_53 ();
 sg13g2_fill_2 FILLER_2_66 ();
 sg13g2_fill_2 FILLER_2_73 ();
 sg13g2_fill_1 FILLER_2_75 ();
 sg13g2_fill_1 FILLER_2_93 ();
 sg13g2_fill_1 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_116 ();
 sg13g2_decap_8 FILLER_2_123 ();
 sg13g2_decap_8 FILLER_2_138 ();
 sg13g2_decap_8 FILLER_2_145 ();
 sg13g2_decap_8 FILLER_2_152 ();
 sg13g2_decap_8 FILLER_2_159 ();
 sg13g2_fill_2 FILLER_2_166 ();
 sg13g2_fill_2 FILLER_2_189 ();
 sg13g2_fill_1 FILLER_2_209 ();
 sg13g2_decap_4 FILLER_2_219 ();
 sg13g2_fill_2 FILLER_2_223 ();
 sg13g2_decap_8 FILLER_2_229 ();
 sg13g2_fill_1 FILLER_2_236 ();
 sg13g2_decap_8 FILLER_2_242 ();
 sg13g2_decap_8 FILLER_2_249 ();
 sg13g2_fill_1 FILLER_2_256 ();
 sg13g2_decap_8 FILLER_2_281 ();
 sg13g2_decap_8 FILLER_2_288 ();
 sg13g2_decap_8 FILLER_2_295 ();
 sg13g2_fill_2 FILLER_2_302 ();
 sg13g2_fill_1 FILLER_2_304 ();
 sg13g2_decap_8 FILLER_2_318 ();
 sg13g2_decap_8 FILLER_2_325 ();
 sg13g2_fill_2 FILLER_2_332 ();
 sg13g2_fill_1 FILLER_2_334 ();
 sg13g2_decap_8 FILLER_2_339 ();
 sg13g2_decap_8 FILLER_2_346 ();
 sg13g2_decap_8 FILLER_2_353 ();
 sg13g2_decap_8 FILLER_2_360 ();
 sg13g2_decap_8 FILLER_2_367 ();
 sg13g2_decap_8 FILLER_2_374 ();
 sg13g2_decap_8 FILLER_2_381 ();
 sg13g2_decap_8 FILLER_2_388 ();
 sg13g2_decap_8 FILLER_2_395 ();
 sg13g2_decap_8 FILLER_2_402 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_fill_2 FILLER_3_64 ();
 sg13g2_fill_1 FILLER_3_66 ();
 sg13g2_fill_1 FILLER_3_94 ();
 sg13g2_fill_2 FILLER_3_116 ();
 sg13g2_fill_1 FILLER_3_118 ();
 sg13g2_decap_4 FILLER_3_145 ();
 sg13g2_fill_2 FILLER_3_222 ();
 sg13g2_fill_1 FILLER_3_224 ();
 sg13g2_fill_2 FILLER_3_260 ();
 sg13g2_fill_1 FILLER_3_262 ();
 sg13g2_fill_2 FILLER_3_298 ();
 sg13g2_decap_4 FILLER_3_326 ();
 sg13g2_fill_2 FILLER_3_335 ();
 sg13g2_fill_2 FILLER_3_346 ();
 sg13g2_fill_1 FILLER_3_348 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_361 ();
 sg13g2_decap_8 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_4 FILLER_3_403 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_fill_2 FILLER_4_35 ();
 sg13g2_fill_1 FILLER_4_37 ();
 sg13g2_fill_1 FILLER_4_158 ();
 sg13g2_fill_1 FILLER_4_173 ();
 sg13g2_fill_1 FILLER_4_217 ();
 sg13g2_fill_2 FILLER_4_231 ();
 sg13g2_fill_1 FILLER_4_259 ();
 sg13g2_fill_2 FILLER_4_291 ();
 sg13g2_fill_1 FILLER_4_293 ();
 sg13g2_fill_1 FILLER_4_334 ();
 sg13g2_fill_1 FILLER_4_369 ();
 sg13g2_decap_8 FILLER_4_374 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_fill_2 FILLER_5_72 ();
 sg13g2_fill_1 FILLER_5_88 ();
 sg13g2_fill_1 FILLER_5_121 ();
 sg13g2_fill_1 FILLER_5_216 ();
 sg13g2_fill_1 FILLER_5_226 ();
 sg13g2_fill_2 FILLER_5_235 ();
 sg13g2_fill_2 FILLER_5_281 ();
 sg13g2_fill_1 FILLER_5_320 ();
 sg13g2_fill_2 FILLER_5_354 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_fill_1 FILLER_6_21 ();
 sg13g2_fill_1 FILLER_6_53 ();
 sg13g2_fill_2 FILLER_6_120 ();
 sg13g2_fill_2 FILLER_6_160 ();
 sg13g2_fill_1 FILLER_6_190 ();
 sg13g2_fill_2 FILLER_6_261 ();
 sg13g2_fill_1 FILLER_6_263 ();
 sg13g2_fill_1 FILLER_6_278 ();
 sg13g2_fill_1 FILLER_6_335 ();
 sg13g2_fill_2 FILLER_6_341 ();
 sg13g2_fill_1 FILLER_6_351 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_fill_2 FILLER_7_56 ();
 sg13g2_fill_2 FILLER_7_154 ();
 sg13g2_fill_1 FILLER_7_217 ();
 sg13g2_fill_1 FILLER_7_236 ();
 sg13g2_fill_2 FILLER_7_250 ();
 sg13g2_fill_1 FILLER_7_252 ();
 sg13g2_fill_1 FILLER_7_342 ();
 sg13g2_fill_1 FILLER_7_370 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_fill_2 FILLER_8_67 ();
 sg13g2_fill_1 FILLER_8_172 ();
 sg13g2_fill_1 FILLER_8_203 ();
 sg13g2_fill_1 FILLER_8_223 ();
 sg13g2_fill_2 FILLER_8_255 ();
 sg13g2_fill_1 FILLER_8_257 ();
 sg13g2_fill_1 FILLER_8_319 ();
 sg13g2_fill_1 FILLER_8_354 ();
 sg13g2_fill_2 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_fill_2 FILLER_9_14 ();
 sg13g2_fill_1 FILLER_9_55 ();
 sg13g2_fill_2 FILLER_9_65 ();
 sg13g2_fill_1 FILLER_9_67 ();
 sg13g2_fill_2 FILLER_9_94 ();
 sg13g2_fill_1 FILLER_9_96 ();
 sg13g2_fill_1 FILLER_9_124 ();
 sg13g2_fill_1 FILLER_9_144 ();
 sg13g2_fill_1 FILLER_9_226 ();
 sg13g2_fill_1 FILLER_9_262 ();
 sg13g2_fill_2 FILLER_9_304 ();
 sg13g2_fill_1 FILLER_9_337 ();
 sg13g2_fill_1 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_4 FILLER_10_14 ();
 sg13g2_fill_1 FILLER_10_97 ();
 sg13g2_fill_2 FILLER_10_137 ();
 sg13g2_fill_1 FILLER_10_190 ();
 sg13g2_fill_2 FILLER_10_210 ();
 sg13g2_fill_1 FILLER_10_218 ();
 sg13g2_fill_2 FILLER_10_300 ();
 sg13g2_fill_1 FILLER_10_354 ();
 sg13g2_fill_2 FILLER_10_375 ();
 sg13g2_fill_1 FILLER_10_382 ();
 sg13g2_fill_2 FILLER_10_388 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_7 ();
 sg13g2_fill_1 FILLER_11_53 ();
 sg13g2_fill_1 FILLER_11_71 ();
 sg13g2_fill_2 FILLER_11_96 ();
 sg13g2_fill_2 FILLER_11_111 ();
 sg13g2_fill_1 FILLER_11_122 ();
 sg13g2_fill_1 FILLER_11_131 ();
 sg13g2_fill_1 FILLER_11_168 ();
 sg13g2_fill_1 FILLER_11_219 ();
 sg13g2_fill_2 FILLER_11_248 ();
 sg13g2_fill_2 FILLER_11_260 ();
 sg13g2_fill_1 FILLER_11_262 ();
 sg13g2_fill_1 FILLER_11_299 ();
 sg13g2_fill_1 FILLER_11_366 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_53 ();
 sg13g2_fill_1 FILLER_12_55 ();
 sg13g2_fill_1 FILLER_12_82 ();
 sg13g2_fill_1 FILLER_12_136 ();
 sg13g2_fill_2 FILLER_12_187 ();
 sg13g2_fill_1 FILLER_12_215 ();
 sg13g2_fill_1 FILLER_12_272 ();
 sg13g2_fill_2 FILLER_12_291 ();
 sg13g2_fill_1 FILLER_12_293 ();
 sg13g2_fill_2 FILLER_12_302 ();
 sg13g2_fill_1 FILLER_12_304 ();
 sg13g2_fill_2 FILLER_12_363 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_2 ();
 sg13g2_fill_2 FILLER_13_38 ();
 sg13g2_fill_1 FILLER_13_40 ();
 sg13g2_fill_1 FILLER_13_59 ();
 sg13g2_fill_1 FILLER_13_122 ();
 sg13g2_fill_2 FILLER_13_235 ();
 sg13g2_fill_2 FILLER_13_258 ();
 sg13g2_fill_1 FILLER_13_260 ();
 sg13g2_fill_2 FILLER_13_278 ();
 sg13g2_fill_2 FILLER_13_312 ();
 sg13g2_fill_2 FILLER_13_350 ();
 sg13g2_fill_1 FILLER_13_352 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_28 ();
 sg13g2_fill_1 FILLER_14_30 ();
 sg13g2_fill_2 FILLER_14_56 ();
 sg13g2_fill_1 FILLER_14_58 ();
 sg13g2_fill_1 FILLER_14_100 ();
 sg13g2_fill_2 FILLER_14_168 ();
 sg13g2_fill_1 FILLER_14_192 ();
 sg13g2_decap_8 FILLER_14_200 ();
 sg13g2_decap_8 FILLER_14_207 ();
 sg13g2_fill_2 FILLER_14_214 ();
 sg13g2_fill_2 FILLER_14_225 ();
 sg13g2_fill_1 FILLER_14_227 ();
 sg13g2_fill_1 FILLER_14_262 ();
 sg13g2_fill_2 FILLER_14_296 ();
 sg13g2_fill_1 FILLER_14_298 ();
 sg13g2_fill_2 FILLER_14_390 ();
 sg13g2_fill_1 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_2 ();
 sg13g2_fill_1 FILLER_15_26 ();
 sg13g2_fill_2 FILLER_15_61 ();
 sg13g2_fill_1 FILLER_15_63 ();
 sg13g2_fill_2 FILLER_15_98 ();
 sg13g2_fill_2 FILLER_15_164 ();
 sg13g2_fill_1 FILLER_15_175 ();
 sg13g2_fill_2 FILLER_15_199 ();
 sg13g2_decap_4 FILLER_15_206 ();
 sg13g2_fill_2 FILLER_15_245 ();
 sg13g2_fill_1 FILLER_15_269 ();
 sg13g2_fill_2 FILLER_15_290 ();
 sg13g2_fill_2 FILLER_15_297 ();
 sg13g2_fill_1 FILLER_15_326 ();
 sg13g2_fill_2 FILLER_15_351 ();
 sg13g2_fill_1 FILLER_15_353 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_fill_2 FILLER_16_35 ();
 sg13g2_fill_2 FILLER_16_61 ();
 sg13g2_fill_2 FILLER_16_94 ();
 sg13g2_fill_2 FILLER_16_180 ();
 sg13g2_fill_2 FILLER_16_208 ();
 sg13g2_fill_1 FILLER_16_210 ();
 sg13g2_fill_1 FILLER_16_225 ();
 sg13g2_fill_2 FILLER_16_229 ();
 sg13g2_fill_1 FILLER_16_231 ();
 sg13g2_fill_2 FILLER_16_241 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_4 ();
 sg13g2_fill_1 FILLER_17_58 ();
 sg13g2_fill_2 FILLER_17_120 ();
 sg13g2_fill_1 FILLER_17_122 ();
 sg13g2_fill_1 FILLER_17_175 ();
 sg13g2_fill_2 FILLER_17_251 ();
 sg13g2_fill_1 FILLER_17_253 ();
 sg13g2_fill_2 FILLER_17_276 ();
 sg13g2_fill_1 FILLER_17_292 ();
 sg13g2_fill_2 FILLER_17_346 ();
 sg13g2_decap_8 FILLER_17_383 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_4 FILLER_18_7 ();
 sg13g2_fill_2 FILLER_18_11 ();
 sg13g2_fill_1 FILLER_18_136 ();
 sg13g2_fill_2 FILLER_18_146 ();
 sg13g2_fill_1 FILLER_18_216 ();
 sg13g2_fill_2 FILLER_18_226 ();
 sg13g2_fill_2 FILLER_18_254 ();
 sg13g2_fill_1 FILLER_18_256 ();
 sg13g2_fill_2 FILLER_18_266 ();
 sg13g2_fill_1 FILLER_18_276 ();
 sg13g2_fill_2 FILLER_18_338 ();
 sg13g2_fill_1 FILLER_18_367 ();
 sg13g2_decap_8 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_4 FILLER_19_14 ();
 sg13g2_fill_2 FILLER_19_18 ();
 sg13g2_fill_2 FILLER_19_105 ();
 sg13g2_fill_1 FILLER_19_117 ();
 sg13g2_fill_2 FILLER_19_133 ();
 sg13g2_fill_2 FILLER_19_177 ();
 sg13g2_fill_1 FILLER_19_179 ();
 sg13g2_decap_8 FILLER_19_206 ();
 sg13g2_fill_2 FILLER_19_222 ();
 sg13g2_fill_1 FILLER_19_224 ();
 sg13g2_decap_4 FILLER_19_237 ();
 sg13g2_fill_1 FILLER_19_241 ();
 sg13g2_fill_1 FILLER_19_326 ();
 sg13g2_fill_1 FILLER_19_335 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_fill_2 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_79 ();
 sg13g2_fill_2 FILLER_20_98 ();
 sg13g2_fill_2 FILLER_20_125 ();
 sg13g2_fill_2 FILLER_20_167 ();
 sg13g2_fill_1 FILLER_20_169 ();
 sg13g2_fill_2 FILLER_20_186 ();
 sg13g2_fill_1 FILLER_20_188 ();
 sg13g2_fill_2 FILLER_20_245 ();
 sg13g2_fill_1 FILLER_20_247 ();
 sg13g2_fill_2 FILLER_20_256 ();
 sg13g2_fill_1 FILLER_20_258 ();
 sg13g2_fill_1 FILLER_20_286 ();
 sg13g2_fill_2 FILLER_20_295 ();
 sg13g2_fill_1 FILLER_20_297 ();
 sg13g2_fill_1 FILLER_20_307 ();
 sg13g2_decap_8 FILLER_20_383 ();
 sg13g2_decap_8 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_397 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_4 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_156 ();
 sg13g2_fill_2 FILLER_21_165 ();
 sg13g2_fill_1 FILLER_21_167 ();
 sg13g2_fill_2 FILLER_21_190 ();
 sg13g2_fill_1 FILLER_21_192 ();
 sg13g2_decap_4 FILLER_21_203 ();
 sg13g2_decap_4 FILLER_21_212 ();
 sg13g2_fill_2 FILLER_21_216 ();
 sg13g2_fill_2 FILLER_21_223 ();
 sg13g2_fill_1 FILLER_21_225 ();
 sg13g2_fill_1 FILLER_21_240 ();
 sg13g2_fill_2 FILLER_21_262 ();
 sg13g2_fill_1 FILLER_21_264 ();
 sg13g2_fill_2 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_332 ();
 sg13g2_fill_1 FILLER_21_339 ();
 sg13g2_fill_2 FILLER_21_344 ();
 sg13g2_fill_1 FILLER_21_350 ();
 sg13g2_fill_2 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_397 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_4 FILLER_22_28 ();
 sg13g2_fill_1 FILLER_22_32 ();
 sg13g2_decap_8 FILLER_22_38 ();
 sg13g2_fill_2 FILLER_22_45 ();
 sg13g2_fill_1 FILLER_22_92 ();
 sg13g2_fill_2 FILLER_22_128 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_fill_2 FILLER_22_210 ();
 sg13g2_fill_1 FILLER_22_241 ();
 sg13g2_fill_2 FILLER_22_268 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_fill_1 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_314 ();
 sg13g2_fill_1 FILLER_22_321 ();
 sg13g2_fill_2 FILLER_22_339 ();
 sg13g2_fill_1 FILLER_22_350 ();
 sg13g2_fill_2 FILLER_22_368 ();
 sg13g2_fill_1 FILLER_22_370 ();
 sg13g2_fill_2 FILLER_22_380 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_4 FILLER_23_49 ();
 sg13g2_fill_2 FILLER_23_53 ();
 sg13g2_fill_2 FILLER_23_74 ();
 sg13g2_fill_2 FILLER_23_156 ();
 sg13g2_fill_2 FILLER_23_175 ();
 sg13g2_fill_1 FILLER_23_177 ();
 sg13g2_fill_2 FILLER_23_191 ();
 sg13g2_fill_1 FILLER_23_193 ();
 sg13g2_decap_4 FILLER_23_212 ();
 sg13g2_fill_1 FILLER_23_216 ();
 sg13g2_decap_4 FILLER_23_243 ();
 sg13g2_fill_1 FILLER_23_256 ();
 sg13g2_fill_2 FILLER_23_296 ();
 sg13g2_fill_1 FILLER_23_298 ();
 sg13g2_fill_2 FILLER_23_325 ();
 sg13g2_fill_2 FILLER_23_357 ();
 sg13g2_fill_1 FILLER_23_359 ();
 sg13g2_decap_8 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_4 FILLER_24_49 ();
 sg13g2_fill_1 FILLER_24_53 ();
 sg13g2_fill_1 FILLER_24_80 ();
 sg13g2_fill_2 FILLER_24_106 ();
 sg13g2_fill_1 FILLER_24_184 ();
 sg13g2_fill_2 FILLER_24_190 ();
 sg13g2_decap_8 FILLER_24_213 ();
 sg13g2_fill_1 FILLER_24_246 ();
 sg13g2_fill_1 FILLER_24_256 ();
 sg13g2_fill_2 FILLER_24_262 ();
 sg13g2_fill_1 FILLER_24_264 ();
 sg13g2_fill_1 FILLER_24_270 ();
 sg13g2_fill_2 FILLER_24_294 ();
 sg13g2_fill_1 FILLER_24_296 ();
 sg13g2_fill_2 FILLER_24_327 ();
 sg13g2_fill_2 FILLER_24_339 ();
 sg13g2_fill_1 FILLER_24_341 ();
 sg13g2_fill_2 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_fill_2 FILLER_25_42 ();
 sg13g2_fill_1 FILLER_25_44 ();
 sg13g2_decap_4 FILLER_25_69 ();
 sg13g2_fill_2 FILLER_25_116 ();
 sg13g2_fill_2 FILLER_25_157 ();
 sg13g2_fill_1 FILLER_25_159 ();
 sg13g2_fill_2 FILLER_25_172 ();
 sg13g2_fill_1 FILLER_25_179 ();
 sg13g2_decap_4 FILLER_25_214 ();
 sg13g2_fill_2 FILLER_25_229 ();
 sg13g2_fill_1 FILLER_25_254 ();
 sg13g2_fill_2 FILLER_25_338 ();
 sg13g2_fill_2 FILLER_25_376 ();
 sg13g2_fill_1 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_388 ();
 sg13g2_decap_8 FILLER_25_395 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_fill_2 FILLER_26_35 ();
 sg13g2_fill_1 FILLER_26_89 ();
 sg13g2_fill_1 FILLER_26_112 ();
 sg13g2_fill_1 FILLER_26_164 ();
 sg13g2_fill_2 FILLER_26_177 ();
 sg13g2_fill_1 FILLER_26_179 ();
 sg13g2_fill_2 FILLER_26_214 ();
 sg13g2_fill_1 FILLER_26_216 ();
 sg13g2_fill_2 FILLER_26_227 ();
 sg13g2_fill_2 FILLER_26_234 ();
 sg13g2_fill_1 FILLER_26_236 ();
 sg13g2_fill_1 FILLER_26_242 ();
 sg13g2_fill_1 FILLER_26_252 ();
 sg13g2_decap_4 FILLER_26_291 ();
 sg13g2_fill_2 FILLER_26_295 ();
 sg13g2_fill_2 FILLER_26_305 ();
 sg13g2_fill_2 FILLER_26_349 ();
 sg13g2_fill_2 FILLER_26_365 ();
 sg13g2_fill_1 FILLER_26_367 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_4 FILLER_27_21 ();
 sg13g2_decap_4 FILLER_27_47 ();
 sg13g2_fill_2 FILLER_27_60 ();
 sg13g2_fill_1 FILLER_27_62 ();
 sg13g2_fill_1 FILLER_27_115 ();
 sg13g2_fill_1 FILLER_27_130 ();
 sg13g2_fill_2 FILLER_27_168 ();
 sg13g2_fill_2 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_181 ();
 sg13g2_fill_2 FILLER_27_188 ();
 sg13g2_fill_1 FILLER_27_190 ();
 sg13g2_fill_2 FILLER_27_224 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_fill_1 FILLER_27_245 ();
 sg13g2_fill_1 FILLER_27_256 ();
 sg13g2_fill_2 FILLER_27_267 ();
 sg13g2_fill_1 FILLER_27_269 ();
 sg13g2_fill_2 FILLER_27_296 ();
 sg13g2_fill_2 FILLER_27_320 ();
 sg13g2_fill_1 FILLER_27_359 ();
 sg13g2_decap_8 FILLER_27_395 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_4 FILLER_28_14 ();
 sg13g2_fill_1 FILLER_28_44 ();
 sg13g2_fill_1 FILLER_28_54 ();
 sg13g2_fill_1 FILLER_28_108 ();
 sg13g2_fill_1 FILLER_28_132 ();
 sg13g2_fill_1 FILLER_28_143 ();
 sg13g2_fill_1 FILLER_28_160 ();
 sg13g2_fill_2 FILLER_28_171 ();
 sg13g2_fill_1 FILLER_28_173 ();
 sg13g2_decap_4 FILLER_28_187 ();
 sg13g2_fill_1 FILLER_28_227 ();
 sg13g2_fill_1 FILLER_28_364 ();
 sg13g2_decap_8 FILLER_28_400 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_fill_1 FILLER_29_28 ();
 sg13g2_fill_1 FILLER_29_68 ();
 sg13g2_fill_2 FILLER_29_151 ();
 sg13g2_fill_1 FILLER_29_153 ();
 sg13g2_fill_2 FILLER_29_167 ();
 sg13g2_fill_2 FILLER_29_178 ();
 sg13g2_fill_1 FILLER_29_198 ();
 sg13g2_decap_4 FILLER_29_260 ();
 sg13g2_fill_2 FILLER_29_264 ();
 sg13g2_fill_2 FILLER_29_275 ();
 sg13g2_fill_1 FILLER_29_277 ();
 sg13g2_fill_2 FILLER_29_376 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_4 FILLER_30_28 ();
 sg13g2_fill_2 FILLER_30_32 ();
 sg13g2_fill_2 FILLER_30_102 ();
 sg13g2_fill_1 FILLER_30_144 ();
 sg13g2_fill_2 FILLER_30_158 ();
 sg13g2_decap_4 FILLER_30_164 ();
 sg13g2_decap_4 FILLER_30_172 ();
 sg13g2_fill_2 FILLER_30_176 ();
 sg13g2_fill_1 FILLER_30_192 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_fill_1 FILLER_30_203 ();
 sg13g2_fill_1 FILLER_30_256 ();
 sg13g2_fill_2 FILLER_30_265 ();
 sg13g2_fill_2 FILLER_30_311 ();
 sg13g2_fill_1 FILLER_30_347 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_4 FILLER_31_21 ();
 sg13g2_fill_2 FILLER_31_62 ();
 sg13g2_fill_1 FILLER_31_64 ();
 sg13g2_fill_2 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_79 ();
 sg13g2_fill_1 FILLER_31_120 ();
 sg13g2_fill_1 FILLER_31_170 ();
 sg13g2_fill_1 FILLER_31_187 ();
 sg13g2_decap_8 FILLER_31_240 ();
 sg13g2_decap_8 FILLER_31_247 ();
 sg13g2_decap_8 FILLER_31_254 ();
 sg13g2_fill_1 FILLER_31_261 ();
 sg13g2_fill_1 FILLER_31_297 ();
 sg13g2_fill_1 FILLER_31_311 ();
 sg13g2_fill_1 FILLER_31_344 ();
 sg13g2_fill_2 FILLER_31_378 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_4 FILLER_32_14 ();
 sg13g2_fill_2 FILLER_32_53 ();
 sg13g2_fill_1 FILLER_32_55 ();
 sg13g2_fill_2 FILLER_32_91 ();
 sg13g2_fill_1 FILLER_32_93 ();
 sg13g2_fill_2 FILLER_32_115 ();
 sg13g2_fill_1 FILLER_32_117 ();
 sg13g2_fill_2 FILLER_32_123 ();
 sg13g2_decap_8 FILLER_32_155 ();
 sg13g2_decap_4 FILLER_32_162 ();
 sg13g2_fill_1 FILLER_32_171 ();
 sg13g2_fill_1 FILLER_32_187 ();
 sg13g2_fill_2 FILLER_32_217 ();
 sg13g2_fill_1 FILLER_32_254 ();
 sg13g2_decap_4 FILLER_32_274 ();
 sg13g2_fill_2 FILLER_32_278 ();
 sg13g2_fill_2 FILLER_32_373 ();
 sg13g2_decap_8 FILLER_32_401 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_4 FILLER_33_28 ();
 sg13g2_fill_1 FILLER_33_32 ();
 sg13g2_decap_4 FILLER_33_67 ();
 sg13g2_decap_4 FILLER_33_85 ();
 sg13g2_fill_1 FILLER_33_89 ();
 sg13g2_fill_1 FILLER_33_154 ();
 sg13g2_fill_2 FILLER_33_206 ();
 sg13g2_decap_4 FILLER_33_258 ();
 sg13g2_fill_1 FILLER_33_353 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_4 FILLER_34_35 ();
 sg13g2_fill_2 FILLER_34_39 ();
 sg13g2_fill_1 FILLER_34_50 ();
 sg13g2_fill_1 FILLER_34_60 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_fill_1 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_153 ();
 sg13g2_fill_2 FILLER_34_164 ();
 sg13g2_fill_1 FILLER_34_196 ();
 sg13g2_fill_2 FILLER_34_201 ();
 sg13g2_fill_1 FILLER_34_203 ();
 sg13g2_fill_2 FILLER_34_216 ();
 sg13g2_fill_2 FILLER_34_258 ();
 sg13g2_decap_8 FILLER_34_388 ();
 sg13g2_decap_8 FILLER_34_395 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_fill_2 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_57 ();
 sg13g2_decap_8 FILLER_35_64 ();
 sg13g2_decap_8 FILLER_35_71 ();
 sg13g2_decap_8 FILLER_35_78 ();
 sg13g2_decap_4 FILLER_35_85 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_4 FILLER_35_105 ();
 sg13g2_fill_2 FILLER_35_262 ();
 sg13g2_fill_1 FILLER_35_301 ();
 sg13g2_fill_2 FILLER_35_339 ();
 sg13g2_fill_1 FILLER_35_341 ();
 sg13g2_decap_4 FILLER_35_345 ();
 sg13g2_fill_1 FILLER_35_349 ();
 sg13g2_fill_2 FILLER_35_363 ();
 sg13g2_fill_1 FILLER_35_365 ();
 sg13g2_decap_8 FILLER_35_379 ();
 sg13g2_decap_8 FILLER_35_386 ();
 sg13g2_decap_8 FILLER_35_393 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_fill_2 FILLER_36_119 ();
 sg13g2_fill_2 FILLER_36_137 ();
 sg13g2_fill_1 FILLER_36_139 ();
 sg13g2_fill_2 FILLER_36_161 ();
 sg13g2_fill_2 FILLER_36_183 ();
 sg13g2_fill_1 FILLER_36_185 ();
 sg13g2_fill_2 FILLER_36_208 ();
 sg13g2_decap_8 FILLER_36_219 ();
 sg13g2_fill_2 FILLER_36_226 ();
 sg13g2_fill_1 FILLER_36_228 ();
 sg13g2_decap_8 FILLER_36_256 ();
 sg13g2_decap_8 FILLER_36_263 ();
 sg13g2_fill_1 FILLER_36_270 ();
 sg13g2_decap_4 FILLER_36_276 ();
 sg13g2_fill_1 FILLER_36_280 ();
 sg13g2_fill_2 FILLER_36_286 ();
 sg13g2_fill_1 FILLER_36_288 ();
 sg13g2_decap_4 FILLER_36_298 ();
 sg13g2_fill_2 FILLER_36_311 ();
 sg13g2_fill_1 FILLER_36_313 ();
 sg13g2_decap_8 FILLER_36_328 ();
 sg13g2_decap_8 FILLER_36_335 ();
 sg13g2_decap_8 FILLER_36_342 ();
 sg13g2_decap_8 FILLER_36_349 ();
 sg13g2_decap_8 FILLER_36_356 ();
 sg13g2_decap_8 FILLER_36_363 ();
 sg13g2_decap_8 FILLER_36_370 ();
 sg13g2_decap_8 FILLER_36_377 ();
 sg13g2_decap_8 FILLER_36_384 ();
 sg13g2_decap_8 FILLER_36_391 ();
 sg13g2_decap_8 FILLER_36_398 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_fill_1 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_198 ();
 sg13g2_fill_1 FILLER_37_205 ();
 sg13g2_decap_8 FILLER_37_209 ();
 sg13g2_decap_8 FILLER_37_216 ();
 sg13g2_decap_8 FILLER_37_223 ();
 sg13g2_decap_8 FILLER_37_230 ();
 sg13g2_decap_8 FILLER_37_237 ();
 sg13g2_decap_8 FILLER_37_244 ();
 sg13g2_decap_8 FILLER_37_251 ();
 sg13g2_decap_8 FILLER_37_258 ();
 sg13g2_decap_8 FILLER_37_265 ();
 sg13g2_decap_8 FILLER_37_272 ();
 sg13g2_decap_8 FILLER_37_279 ();
 sg13g2_decap_8 FILLER_37_286 ();
 sg13g2_decap_4 FILLER_37_293 ();
 sg13g2_decap_8 FILLER_37_302 ();
 sg13g2_decap_8 FILLER_37_309 ();
 sg13g2_decap_8 FILLER_37_316 ();
 sg13g2_decap_8 FILLER_37_323 ();
 sg13g2_decap_8 FILLER_37_330 ();
 sg13g2_decap_8 FILLER_37_337 ();
 sg13g2_decap_8 FILLER_37_344 ();
 sg13g2_decap_8 FILLER_37_351 ();
 sg13g2_decap_8 FILLER_37_358 ();
 sg13g2_decap_8 FILLER_37_365 ();
 sg13g2_decap_8 FILLER_37_372 ();
 sg13g2_decap_8 FILLER_37_379 ();
 sg13g2_decap_8 FILLER_37_386 ();
 sg13g2_decap_8 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_fill_2 FILLER_38_174 ();
 sg13g2_decap_8 FILLER_38_193 ();
 sg13g2_decap_8 FILLER_38_200 ();
 sg13g2_decap_8 FILLER_38_207 ();
 sg13g2_decap_8 FILLER_38_214 ();
 sg13g2_decap_8 FILLER_38_221 ();
 sg13g2_decap_8 FILLER_38_228 ();
 sg13g2_decap_8 FILLER_38_235 ();
 sg13g2_decap_8 FILLER_38_242 ();
 sg13g2_decap_8 FILLER_38_249 ();
 sg13g2_decap_8 FILLER_38_256 ();
 sg13g2_decap_8 FILLER_38_263 ();
 sg13g2_decap_8 FILLER_38_270 ();
 sg13g2_decap_8 FILLER_38_277 ();
 sg13g2_decap_8 FILLER_38_284 ();
 sg13g2_decap_8 FILLER_38_291 ();
 sg13g2_decap_8 FILLER_38_298 ();
 sg13g2_decap_8 FILLER_38_305 ();
 sg13g2_decap_8 FILLER_38_312 ();
 sg13g2_decap_8 FILLER_38_319 ();
 sg13g2_decap_8 FILLER_38_326 ();
 sg13g2_decap_8 FILLER_38_333 ();
 sg13g2_decap_8 FILLER_38_340 ();
 sg13g2_decap_8 FILLER_38_347 ();
 sg13g2_decap_8 FILLER_38_354 ();
 sg13g2_decap_8 FILLER_38_361 ();
 sg13g2_decap_8 FILLER_38_368 ();
 sg13g2_decap_8 FILLER_38_375 ();
 sg13g2_decap_8 FILLER_38_382 ();
 sg13g2_decap_8 FILLER_38_389 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net1;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net3;
 assign uio_oe[3] = net4;
 assign uio_oe[4] = net5;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net15;
 assign uio_out[0] = net8;
 assign uio_out[1] = net9;
 assign uio_out[2] = net10;
 assign uio_out[3] = net11;
 assign uio_out[4] = net12;
 assign uio_out[5] = net13;
 assign uio_out[6] = net14;
endmodule

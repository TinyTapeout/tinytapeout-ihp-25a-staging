module tt_um_demosiine_sda (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire audio;
 wire \audio_engine_1.counter[0] ;
 wire \audio_engine_1.counter[10] ;
 wire \audio_engine_1.counter[11] ;
 wire \audio_engine_1.counter[12] ;
 wire \audio_engine_1.counter[13] ;
 wire \audio_engine_1.counter[14] ;
 wire \audio_engine_1.counter[15] ;
 wire \audio_engine_1.counter[16] ;
 wire \audio_engine_1.counter[17] ;
 wire \audio_engine_1.counter[1] ;
 wire \audio_engine_1.counter[2] ;
 wire \audio_engine_1.counter[3] ;
 wire \audio_engine_1.counter[4] ;
 wire \audio_engine_1.counter[5] ;
 wire \audio_engine_1.counter[6] ;
 wire \audio_engine_1.counter[7] ;
 wire \audio_engine_1.counter[8] ;
 wire \audio_engine_1.counter[9] ;
 wire \audio_engine_1.en_seq_clk ;
 wire \audio_engine_1.freq_synth1.audio_reg ;
 wire \audio_engine_1.freq_synth1.en_synth_clk ;
 wire \audio_engine_1.freq_synth1.hp_ctr[0] ;
 wire \audio_engine_1.freq_synth1.hp_ctr[1] ;
 wire \audio_engine_1.freq_synth1.hp_ctr[2] ;
 wire \audio_engine_1.freq_synth1.hp_ctr[3] ;
 wire \audio_engine_1.freq_synth1.hp_ctr[4] ;
 wire \audio_engine_1.freq_synth1.hp_ctr[5] ;
 wire \audio_engine_1.freq_synth1.hp_ctr[6] ;
 wire \audio_engine_1.seq_ctr[0] ;
 wire \audio_engine_1.seq_ctr[1] ;
 wire \audio_engine_1.seq_ctr[2] ;
 wire \audio_engine_1.seq_ctr[3] ;
 wire \audio_engine_1.seq_ctr[4] ;
 wire \audio_engine_1.seq_time[0] ;
 wire \audio_engine_1.seq_time[1] ;
 wire \audio_engine_1.seq_time[2] ;
 wire \audio_engine_1.seq_time[3] ;
 wire \audio_engine_1.seq_time[4] ;
 wire \audio_engine_1.seq_time[5] ;
 wire \audio_engine_1.seq_time[6] ;
 wire \graphics_engine_1.anim_2x[0] ;
 wire \graphics_engine_1.ctr[0] ;
 wire \graphics_engine_1.ctr[1] ;
 wire \graphics_engine_1.ctr[2] ;
 wire \graphics_engine_1.ctr[3] ;
 wire \graphics_engine_1.ctr[4] ;
 wire \graphics_engine_1.ctr[5] ;
 wire \graphics_engine_1.ctr[6] ;
 wire \graphics_engine_1.ctr[7] ;
 wire \graphics_engine_1.ctr[8] ;
 wire \graphics_engine_1.en_v_sync ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_x[0] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_y[0] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_y[1] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.x[1] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.x[2] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.x[4] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.x[5] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.x[6] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.x[7] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.x[8] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.x[9] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.y[0] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.y[1] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.y[2] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.y[5] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.y[6] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.y[7] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.y[8] ;
 wire \graphics_engine_1.v_sync ;
 wire h_sync;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire clknet_0_clk;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire \vga_controller_1.y[9] ;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;

 sg13g2_inv_1 _1710_ (.Y(_0039_),
    .A(net45));
 sg13g2_inv_1 _1711_ (.Y(_0038_),
    .A(net46));
 sg13g2_inv_1 _1712_ (.Y(_0852_),
    .A(net50));
 sg13g2_inv_1 _1713_ (.Y(_0853_),
    .A(\audio_engine_1.seq_ctr[3] ));
 sg13g2_inv_1 _1714_ (.Y(_0854_),
    .A(net476));
 sg13g2_inv_1 _1715_ (.Y(_0855_),
    .A(net471));
 sg13g2_inv_1 _1716_ (.Y(_0856_),
    .A(net469));
 sg13g2_inv_2 _1717_ (.Y(_0857_),
    .A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[8] ));
 sg13g2_inv_2 _1718_ (.Y(_0858_),
    .A(net501));
 sg13g2_inv_2 _1719_ (.Y(_0859_),
    .A(net511));
 sg13g2_inv_1 _1720_ (.Y(_0860_),
    .A(net485));
 sg13g2_inv_4 _1721_ (.A(net482),
    .Y(_0861_));
 sg13g2_inv_2 _1722_ (.Y(_0862_),
    .A(net480));
 sg13g2_inv_1 _1723_ (.Y(_0863_),
    .A(net494));
 sg13g2_inv_1 _1724_ (.Y(_0864_),
    .A(\graphics_engine_1.ctr[0] ));
 sg13g2_inv_2 _1725_ (.Y(_0865_),
    .A(_0028_));
 sg13g2_inv_1 _1726_ (.Y(_0866_),
    .A(net3));
 sg13g2_inv_1 _1727_ (.Y(_0867_),
    .A(net4));
 sg13g2_inv_1 _1728_ (.Y(_0868_),
    .A(\audio_engine_1.freq_synth1.audio_reg ));
 sg13g2_inv_1 _1729_ (.Y(_0869_),
    .A(\audio_engine_1.counter[2] ));
 sg13g2_inv_1 _1730_ (.Y(_0870_),
    .A(net80));
 sg13g2_nand2_2 _1731_ (.Y(_0871_),
    .A(net157),
    .B(net500));
 sg13g2_and2_1 _1732_ (.A(net498),
    .B(net501),
    .X(_0872_));
 sg13g2_nand2_1 _1733_ (.Y(_0873_),
    .A(net499),
    .B(net501));
 sg13g2_nor3_2 _1734_ (.A(_0857_),
    .B(_0858_),
    .C(_0871_),
    .Y(_0874_));
 sg13g2_nor2_2 _1735_ (.A(net507),
    .B(_0859_),
    .Y(_0875_));
 sg13g2_nor2_1 _1736_ (.A(net133),
    .B(net513),
    .Y(_0876_));
 sg13g2_and4_1 _1737_ (.A(net154),
    .B(_0874_),
    .C(_0875_),
    .D(_0876_),
    .X(_0005_));
 sg13g2_nor2_2 _1738_ (.A(net468),
    .B(_0861_),
    .Y(_0877_));
 sg13g2_nand2_2 _1739_ (.Y(_0878_),
    .A(net485),
    .B(net482));
 sg13g2_nor2_1 _1740_ (.A(_0862_),
    .B(_0878_),
    .Y(_0879_));
 sg13g2_nand2_1 _1741_ (.Y(_0880_),
    .A(net478),
    .B(_0879_));
 sg13g2_a21oi_1 _1742_ (.A1(net478),
    .A2(_0879_),
    .Y(_0881_),
    .B1(\graphics_engine_1.overlay_creator1.text_demosiine1.x[8] ));
 sg13g2_nor2_2 _1743_ (.A(net485),
    .B(net482),
    .Y(_0882_));
 sg13g2_nand2_2 _1744_ (.Y(_0883_),
    .A(net468),
    .B(_0861_));
 sg13g2_nor2_1 _1745_ (.A(net480),
    .B(_0883_),
    .Y(_0884_));
 sg13g2_o21ai_1 _1746_ (.B1(net478),
    .Y(_0885_),
    .A1(net480),
    .A2(_0883_));
 sg13g2_nor2b_1 _1747_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[8] ),
    .B_N(_0885_),
    .Y(_0886_));
 sg13g2_o21ai_1 _1748_ (.B1(net120),
    .Y(_0887_),
    .A1(_0015_),
    .A2(_0881_));
 sg13g2_nor2_1 _1749_ (.A(_0886_),
    .B(net121),
    .Y(_0004_));
 sg13g2_nor2_2 _1750_ (.A(net487),
    .B(net491),
    .Y(_0888_));
 sg13g2_nand2_2 _1751_ (.Y(_0889_),
    .A(_0860_),
    .B(net466));
 sg13g2_nor2_1 _1752_ (.A(net495),
    .B(net491),
    .Y(_0890_));
 sg13g2_nor2_1 _1753_ (.A(net495),
    .B(_0889_),
    .Y(_0891_));
 sg13g2_nor3_2 _1754_ (.A(net483),
    .B(net495),
    .C(_0889_),
    .Y(_0892_));
 sg13g2_nand2_1 _1755_ (.Y(_0893_),
    .A(_0862_),
    .B(_0892_));
 sg13g2_xor2_1 _1756_ (.B(_0893_),
    .A(_0017_),
    .X(_0894_));
 sg13g2_inv_1 _1757_ (.Y(_0895_),
    .A(_0894_));
 sg13g2_xnor2_1 _1758_ (.Y(_0896_),
    .A(_0018_),
    .B(_0892_));
 sg13g2_inv_1 _1759_ (.Y(_0897_),
    .A(net452));
 sg13g2_xnor2_1 _1760_ (.Y(_0898_),
    .A(_0023_),
    .B(_0891_));
 sg13g2_xnor2_1 _1761_ (.Y(_0899_),
    .A(net484),
    .B(_0890_));
 sg13g2_xor2_1 _1762_ (.B(_0890_),
    .A(net484),
    .X(_0900_));
 sg13g2_nor2_2 _1763_ (.A(net451),
    .B(_0899_),
    .Y(_0901_));
 sg13g2_nor3_1 _1764_ (.A(net452),
    .B(net451),
    .C(_0899_),
    .Y(_0902_));
 sg13g2_nor2_1 _1765_ (.A(_0895_),
    .B(_0902_),
    .Y(_0903_));
 sg13g2_xnor2_1 _1766_ (.Y(_0904_),
    .A(_0894_),
    .B(_0902_));
 sg13g2_nor2_1 _1767_ (.A(net478),
    .B(_0893_),
    .Y(_0905_));
 sg13g2_xnor2_1 _1768_ (.Y(_0906_),
    .A(_0016_),
    .B(_0905_));
 sg13g2_nor2_1 _1769_ (.A(net509),
    .B(net513),
    .Y(_0907_));
 sg13g2_xor2_1 _1770_ (.B(net512),
    .A(net509),
    .X(_0908_));
 sg13g2_xnor2_1 _1771_ (.Y(_0909_),
    .A(net509),
    .B(net512));
 sg13g2_and2_1 _1772_ (.A(net503),
    .B(_0908_),
    .X(_0910_));
 sg13g2_nand2_2 _1773_ (.Y(_0911_),
    .A(net503),
    .B(_0908_));
 sg13g2_nor2_2 _1774_ (.A(net501),
    .B(net506),
    .Y(_0912_));
 sg13g2_nor2_2 _1775_ (.A(net505),
    .B(net508),
    .Y(_0913_));
 sg13g2_or2_2 _1776_ (.X(_0914_),
    .B(net508),
    .A(net505));
 sg13g2_nor3_2 _1777_ (.A(net506),
    .B(net509),
    .C(net512),
    .Y(_0915_));
 sg13g2_nor4_2 _1778_ (.A(net502),
    .B(net506),
    .C(net509),
    .Y(_0916_),
    .D(net512));
 sg13g2_xnor2_1 _1779_ (.Y(_0917_),
    .A(_0865_),
    .B(_0916_));
 sg13g2_xnor2_1 _1780_ (.Y(_0918_),
    .A(_0028_),
    .B(_0916_));
 sg13g2_nor2_2 _1781_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[7] ),
    .B(net500),
    .Y(_0919_));
 sg13g2_nor2b_1 _1782_ (.A(net499),
    .B_N(_0916_),
    .Y(_0920_));
 sg13g2_nand2_1 _1783_ (.Y(_0921_),
    .A(_0916_),
    .B(_0919_));
 sg13g2_xnor2_1 _1784_ (.Y(_0922_),
    .A(_0022_),
    .B(_0921_));
 sg13g2_xor2_1 _1785_ (.B(_0921_),
    .A(_0022_),
    .X(_0923_));
 sg13g2_xnor2_1 _1786_ (.Y(_0924_),
    .A(net497),
    .B(_0920_));
 sg13g2_xor2_1 _1787_ (.B(_0920_),
    .A(net497),
    .X(_0925_));
 sg13g2_xnor2_1 _1788_ (.Y(_0926_),
    .A(_0021_),
    .B(_0915_));
 sg13g2_xor2_1 _1789_ (.B(_0915_),
    .A(_0021_),
    .X(_0927_));
 sg13g2_nor2_2 _1790_ (.A(_0917_),
    .B(_0927_),
    .Y(_0928_));
 sg13g2_nand2_2 _1791_ (.Y(_0929_),
    .A(_0918_),
    .B(_0926_));
 sg13g2_xnor2_1 _1792_ (.Y(_0930_),
    .A(_0924_),
    .B(_0928_));
 sg13g2_nor4_2 _1793_ (.A(_0911_),
    .B(_0918_),
    .C(net455),
    .Y(_0931_),
    .D(_0925_));
 sg13g2_nor2_1 _1794_ (.A(_0918_),
    .B(_0926_),
    .Y(_0932_));
 sg13g2_nor4_2 _1795_ (.A(_0918_),
    .B(net455),
    .C(_0925_),
    .Y(_0933_),
    .D(_0926_));
 sg13g2_and2_1 _1796_ (.A(_0911_),
    .B(_0933_),
    .X(_0934_));
 sg13g2_or2_2 _1797_ (.X(_0935_),
    .B(_0933_),
    .A(net450));
 sg13g2_nor3_2 _1798_ (.A(net455),
    .B(_0924_),
    .C(_0929_),
    .Y(_0936_));
 sg13g2_or2_1 _1799_ (.X(_0937_),
    .B(_0936_),
    .A(_0935_));
 sg13g2_a21o_1 _1800_ (.A2(_0936_),
    .A1(_0911_),
    .B1(_0935_),
    .X(_0938_));
 sg13g2_xor2_1 _1801_ (.B(net491),
    .A(net495),
    .X(_0939_));
 sg13g2_xnor2_1 _1802_ (.Y(_0940_),
    .A(net495),
    .B(net491));
 sg13g2_nor2_2 _1803_ (.A(net503),
    .B(_0909_),
    .Y(_0941_));
 sg13g2_and2_2 _1804_ (.A(_0933_),
    .B(_0941_),
    .X(_0942_));
 sg13g2_nand2_1 _1805_ (.Y(_0943_),
    .A(net460),
    .B(_0942_));
 sg13g2_xor2_1 _1806_ (.B(_0907_),
    .A(net503),
    .X(_0944_));
 sg13g2_xnor2_1 _1807_ (.Y(_0945_),
    .A(net503),
    .B(_0907_));
 sg13g2_nor2_2 _1808_ (.A(_0908_),
    .B(_0945_),
    .Y(_0946_));
 sg13g2_nand3_1 _1809_ (.B(net461),
    .C(_0946_),
    .A(_0933_),
    .Y(_0947_));
 sg13g2_nand3_1 _1810_ (.B(_0943_),
    .C(_0947_),
    .A(_0938_),
    .Y(_0948_));
 sg13g2_xnor2_1 _1811_ (.Y(_0949_),
    .A(net452),
    .B(_0901_));
 sg13g2_xnor2_1 _1812_ (.Y(_0950_),
    .A(_0897_),
    .B(_0901_));
 sg13g2_nand2_2 _1813_ (.Y(_0951_),
    .A(_0019_),
    .B(net464));
 sg13g2_inv_1 _1814_ (.Y(_0952_),
    .A(_0951_));
 sg13g2_nand2_1 _1815_ (.Y(_0953_),
    .A(_0910_),
    .B(_0932_));
 sg13g2_nor2_1 _1816_ (.A(_0908_),
    .B(_0944_),
    .Y(_0954_));
 sg13g2_a22oi_1 _1817_ (.Y(_0955_),
    .B1(_0933_),
    .B2(_0954_),
    .A2(net450),
    .A1(_0927_));
 sg13g2_o21ai_1 _1818_ (.B1(_0950_),
    .Y(_0956_),
    .A1(_0951_),
    .A2(_0955_));
 sg13g2_nand2_1 _1819_ (.Y(_0957_),
    .A(_0911_),
    .B(_0928_));
 sg13g2_and2_1 _1820_ (.A(_0953_),
    .B(_0957_),
    .X(_0958_));
 sg13g2_nand3_1 _1821_ (.B(_0928_),
    .C(_0944_),
    .A(_0909_),
    .Y(_0959_));
 sg13g2_nor3_1 _1822_ (.A(net455),
    .B(_0930_),
    .C(_0959_),
    .Y(_0960_));
 sg13g2_or3_1 _1823_ (.A(_0931_),
    .B(net461),
    .C(_0960_),
    .X(_0961_));
 sg13g2_nor2_2 _1824_ (.A(net450),
    .B(net463),
    .Y(_0962_));
 sg13g2_o21ai_1 _1825_ (.B1(_0938_),
    .Y(_0963_),
    .A1(_0900_),
    .A2(_0962_));
 sg13g2_a221oi_1 _1826_ (.B2(_0963_),
    .C1(_0956_),
    .B1(_0961_),
    .A1(_0900_),
    .Y(_0964_),
    .A2(_0948_));
 sg13g2_and2_2 _1827_ (.A(net451),
    .B(_0899_),
    .X(_0965_));
 sg13g2_nand2_1 _1828_ (.Y(_0966_),
    .A(net451),
    .B(_0899_));
 sg13g2_nor2_2 _1829_ (.A(_0901_),
    .B(_0965_),
    .Y(_0967_));
 sg13g2_nand2b_1 _1830_ (.Y(_0968_),
    .B(_0966_),
    .A_N(_0901_));
 sg13g2_nor2_1 _1831_ (.A(net484),
    .B(net460),
    .Y(_0969_));
 sg13g2_nand2b_2 _1832_ (.Y(_0970_),
    .B(net465),
    .A_N(net484));
 sg13g2_nand2_1 _1833_ (.Y(_0971_),
    .A(_0900_),
    .B(net460));
 sg13g2_nor2_2 _1834_ (.A(_0900_),
    .B(net463),
    .Y(_0972_));
 sg13g2_nand2_2 _1835_ (.Y(_0973_),
    .A(_0899_),
    .B(net460));
 sg13g2_nand2_1 _1836_ (.Y(_0974_),
    .A(_0951_),
    .B(_0973_));
 sg13g2_nand2_2 _1837_ (.Y(_0975_),
    .A(_0970_),
    .B(_0971_));
 sg13g2_a221oi_1 _1838_ (.B2(net450),
    .C1(_0950_),
    .B1(_0975_),
    .A1(_0934_),
    .Y(_0976_),
    .A2(net463));
 sg13g2_nor2_1 _1839_ (.A(_0934_),
    .B(net463),
    .Y(_0977_));
 sg13g2_o21ai_1 _1840_ (.B1(_0899_),
    .Y(_0978_),
    .A1(net450),
    .A2(net461));
 sg13g2_nor2_1 _1841_ (.A(_0977_),
    .B(_0978_),
    .Y(_0979_));
 sg13g2_nand2_2 _1842_ (.Y(_0980_),
    .A(_0926_),
    .B(_0945_));
 sg13g2_nand2_1 _1843_ (.Y(_0981_),
    .A(_0936_),
    .B(_0945_));
 sg13g2_nand2_1 _1844_ (.Y(_0982_),
    .A(_0926_),
    .B(_0931_));
 sg13g2_a21oi_1 _1845_ (.A1(_0981_),
    .A2(_0982_),
    .Y(_0983_),
    .B1(_0971_));
 sg13g2_nand2_1 _1846_ (.Y(_0984_),
    .A(_0935_),
    .B(_0970_));
 sg13g2_o21ai_1 _1847_ (.B1(_0949_),
    .Y(_0985_),
    .A1(_0979_),
    .A2(_0983_));
 sg13g2_or3_1 _1848_ (.A(_0949_),
    .B(_0962_),
    .C(_0984_),
    .X(_0986_));
 sg13g2_nand3_1 _1849_ (.B(_0985_),
    .C(_0986_),
    .A(_0968_),
    .Y(_0987_));
 sg13g2_o21ai_1 _1850_ (.B1(_0967_),
    .Y(_0988_),
    .A1(_0964_),
    .A2(_0976_));
 sg13g2_nand3_1 _1851_ (.B(_0987_),
    .C(_0988_),
    .A(_0906_),
    .Y(_0989_));
 sg13g2_nand2_1 _1852_ (.Y(_0990_),
    .A(_0904_),
    .B(_0989_));
 sg13g2_or2_1 _1853_ (.X(_0991_),
    .B(_0906_),
    .A(_0903_));
 sg13g2_nor2_2 _1854_ (.A(net479),
    .B(\graphics_engine_1.overlay_creator1.text_demosiine1.x[8] ),
    .Y(_0992_));
 sg13g2_nand3_1 _1855_ (.B(_0892_),
    .C(_0992_),
    .A(_0862_),
    .Y(_0993_));
 sg13g2_xor2_1 _1856_ (.B(_0993_),
    .A(_0015_),
    .X(_0994_));
 sg13g2_inv_1 _1857_ (.Y(_0995_),
    .A(_0994_));
 sg13g2_nand4_1 _1858_ (.B(_0990_),
    .C(_0991_),
    .A(_0937_),
    .Y(_0996_),
    .D(_0995_));
 sg13g2_nand2_1 _1859_ (.Y(_0997_),
    .A(_0903_),
    .B(_0906_));
 sg13g2_a221oi_1 _1860_ (.B2(_0946_),
    .C1(_0942_),
    .B1(_0933_),
    .A1(_0927_),
    .Y(_0998_),
    .A2(net450));
 sg13g2_nand2_1 _1861_ (.Y(_0999_),
    .A(_0981_),
    .B(_0998_));
 sg13g2_nand2_1 _1862_ (.Y(_1000_),
    .A(_0938_),
    .B(_0982_));
 sg13g2_nor3_1 _1863_ (.A(net460),
    .B(_0999_),
    .C(_1000_),
    .Y(_1001_));
 sg13g2_a21oi_1 _1864_ (.A1(net460),
    .A2(_0999_),
    .Y(_1002_),
    .B1(_0900_));
 sg13g2_nand2b_1 _1865_ (.Y(_1003_),
    .B(_1002_),
    .A_N(_1001_));
 sg13g2_nand2_1 _1866_ (.Y(_1004_),
    .A(_0935_),
    .B(net460));
 sg13g2_nand3_1 _1867_ (.B(_0970_),
    .C(_0982_),
    .A(_0938_),
    .Y(_1005_));
 sg13g2_a21oi_1 _1868_ (.A1(_0966_),
    .A2(_1004_),
    .Y(_1006_),
    .B1(_0967_));
 sg13g2_a221oi_1 _1869_ (.B2(_1003_),
    .C1(_0950_),
    .B1(_1006_),
    .A1(_0967_),
    .Y(_1007_),
    .A2(_1005_));
 sg13g2_a221oi_1 _1870_ (.B2(_0935_),
    .C1(_0967_),
    .B1(_0969_),
    .A1(net463),
    .Y(_1008_),
    .A2(_0942_));
 sg13g2_a221oi_1 _1871_ (.B2(net450),
    .C1(_0968_),
    .B1(_0971_),
    .A1(_0899_),
    .Y(_1009_),
    .A2(_0942_));
 sg13g2_a21oi_1 _1872_ (.A1(_0947_),
    .A2(_1008_),
    .Y(_1010_),
    .B1(_1009_));
 sg13g2_nor2_1 _1873_ (.A(_0949_),
    .B(_1010_),
    .Y(_1011_));
 sg13g2_o21ai_1 _1874_ (.B1(_0997_),
    .Y(_1012_),
    .A1(_1007_),
    .A2(_1011_));
 sg13g2_a21oi_1 _1875_ (.A1(net463),
    .A2(_0942_),
    .Y(_1013_),
    .B1(net450));
 sg13g2_nand3_1 _1876_ (.B(_0967_),
    .C(_0973_),
    .A(_0935_),
    .Y(_1014_));
 sg13g2_o21ai_1 _1877_ (.B1(_1014_),
    .Y(_1015_),
    .A1(_0966_),
    .A2(_1013_));
 sg13g2_nand2b_1 _1878_ (.Y(_1016_),
    .B(_0962_),
    .A_N(_0942_));
 sg13g2_nand3_1 _1879_ (.B(_1015_),
    .C(_1016_),
    .A(_0950_),
    .Y(_1017_));
 sg13g2_o21ai_1 _1880_ (.B1(_0967_),
    .Y(_1018_),
    .A1(_0962_),
    .A2(_0984_));
 sg13g2_a21oi_1 _1881_ (.A1(_0965_),
    .A2(_1004_),
    .Y(_1019_),
    .B1(_0950_));
 sg13g2_nand3_1 _1882_ (.B(net463),
    .C(_0946_),
    .A(_0933_),
    .Y(_1020_));
 sg13g2_nand3_1 _1883_ (.B(_0943_),
    .C(_1020_),
    .A(_0901_),
    .Y(_1021_));
 sg13g2_nand3_1 _1884_ (.B(_1019_),
    .C(_1021_),
    .A(_1018_),
    .Y(_1022_));
 sg13g2_nand4_1 _1885_ (.B(_0906_),
    .C(_1017_),
    .A(_0903_),
    .Y(_1023_),
    .D(_1022_));
 sg13g2_a21oi_1 _1886_ (.A1(_1012_),
    .A2(_1023_),
    .Y(_1024_),
    .B1(_0904_));
 sg13g2_or2_1 _1887_ (.X(_1025_),
    .B(_1024_),
    .A(_0996_));
 sg13g2_nor2_1 _1888_ (.A(net451),
    .B(_0972_),
    .Y(_1026_));
 sg13g2_nand2b_1 _1889_ (.Y(_1027_),
    .B(_0973_),
    .A_N(net451));
 sg13g2_a21oi_1 _1890_ (.A1(net453),
    .A2(_1027_),
    .Y(_1028_),
    .B1(_0894_));
 sg13g2_xor2_1 _1891_ (.B(_1028_),
    .A(_0906_),
    .X(_1029_));
 sg13g2_a21oi_2 _1892_ (.B1(_0918_),
    .Y(_1030_),
    .A2(_0945_),
    .A1(_0926_));
 sg13g2_nand2_1 _1893_ (.Y(_1031_),
    .A(_0925_),
    .B(_1030_));
 sg13g2_nand2b_1 _1894_ (.Y(_1032_),
    .B(_0924_),
    .A_N(_1030_));
 sg13g2_xnor2_1 _1895_ (.Y(_1033_),
    .A(_0924_),
    .B(_1030_));
 sg13g2_nand2_2 _1896_ (.Y(_1034_),
    .A(_0923_),
    .B(_1033_));
 sg13g2_a21oi_2 _1897_ (.B1(_0917_),
    .Y(_1035_),
    .A2(_0944_),
    .A1(_0927_));
 sg13g2_and2_1 _1898_ (.A(_0980_),
    .B(_1035_),
    .X(_1036_));
 sg13g2_nand3_1 _1899_ (.B(_0980_),
    .C(_1035_),
    .A(_0941_),
    .Y(_1037_));
 sg13g2_nand4_1 _1900_ (.B(_0941_),
    .C(_1033_),
    .A(net455),
    .Y(_1038_),
    .D(_1036_));
 sg13g2_nor4_2 _1901_ (.A(_0908_),
    .B(_0917_),
    .C(_0926_),
    .Y(_1039_),
    .D(_0944_));
 sg13g2_nand3_1 _1902_ (.B(_1033_),
    .C(_1039_),
    .A(net455),
    .Y(_1040_));
 sg13g2_and2_1 _1903_ (.A(_1038_),
    .B(_1040_),
    .X(_1041_));
 sg13g2_nand2_1 _1904_ (.Y(_1042_),
    .A(_1038_),
    .B(_1040_));
 sg13g2_nand2_1 _1905_ (.Y(_1043_),
    .A(_0928_),
    .B(_0941_));
 sg13g2_nand3_1 _1906_ (.B(_0980_),
    .C(_1035_),
    .A(_0910_),
    .Y(_1044_));
 sg13g2_nand3_1 _1907_ (.B(_1043_),
    .C(_1044_),
    .A(_0959_),
    .Y(_1045_));
 sg13g2_nor2b_1 _1908_ (.A(_1034_),
    .B_N(_1045_),
    .Y(_1046_));
 sg13g2_nor2_1 _1909_ (.A(_1042_),
    .B(_1046_),
    .Y(_1047_));
 sg13g2_nor4_2 _1910_ (.A(_0908_),
    .B(_0929_),
    .C(_0944_),
    .Y(_1048_),
    .D(_1034_));
 sg13g2_nor4_2 _1911_ (.A(_0922_),
    .B(_0924_),
    .C(_1030_),
    .Y(_1049_),
    .D(_1035_));
 sg13g2_nor2b_1 _1912_ (.A(_0941_),
    .B_N(_1049_),
    .Y(_1050_));
 sg13g2_nand2_1 _1913_ (.Y(_1051_),
    .A(_0954_),
    .B(_1049_));
 sg13g2_nand2_1 _1914_ (.Y(_1052_),
    .A(_0944_),
    .B(_1049_));
 sg13g2_nor4_1 _1915_ (.A(_1042_),
    .B(_1046_),
    .C(_1048_),
    .D(_1050_),
    .Y(_1053_));
 sg13g2_xnor2_1 _1916_ (.Y(_1054_),
    .A(_0911_),
    .B(_0926_));
 sg13g2_or2_1 _1917_ (.X(_1055_),
    .B(_1054_),
    .A(net415));
 sg13g2_o21ai_1 _1918_ (.B1(_0952_),
    .Y(_1056_),
    .A1(net415),
    .A2(_1054_));
 sg13g2_and4_2 _1919_ (.A(_0910_),
    .B(net455),
    .C(_1033_),
    .D(_1036_),
    .X(_1057_));
 sg13g2_or2_1 _1920_ (.X(_1058_),
    .B(_1044_),
    .A(_1034_));
 sg13g2_nor2_2 _1921_ (.A(_0908_),
    .B(_1052_),
    .Y(_1059_));
 sg13g2_a21oi_1 _1922_ (.A1(_0946_),
    .A2(_1049_),
    .Y(_1060_),
    .B1(_1057_));
 sg13g2_or2_1 _1923_ (.X(_1061_),
    .B(_1059_),
    .A(_1057_));
 sg13g2_a22oi_1 _1924_ (.Y(_1062_),
    .B1(_1061_),
    .B2(net462),
    .A2(_1056_),
    .A1(_0973_));
 sg13g2_xnor2_1 _1925_ (.Y(_1063_),
    .A(_0898_),
    .B(_0972_));
 sg13g2_o21ai_1 _1926_ (.B1(net449),
    .Y(_1064_),
    .A1(net464),
    .A2(_1058_));
 sg13g2_nand2_1 _1927_ (.Y(_1065_),
    .A(net445),
    .B(_1064_));
 sg13g2_xnor2_1 _1928_ (.Y(_1066_),
    .A(net453),
    .B(_1026_));
 sg13g2_nand2_1 _1929_ (.Y(_1067_),
    .A(net464),
    .B(_1042_));
 sg13g2_nor2_2 _1930_ (.A(net462),
    .B(_1059_),
    .Y(_1068_));
 sg13g2_nand2_1 _1931_ (.Y(_1069_),
    .A(net462),
    .B(_1060_));
 sg13g2_or2_1 _1932_ (.X(_1070_),
    .B(_1069_),
    .A(_1048_));
 sg13g2_a221oi_1 _1933_ (.B2(_1047_),
    .C1(net445),
    .B1(_1068_),
    .A1(_0975_),
    .Y(_1071_),
    .A2(_1067_));
 sg13g2_a21oi_1 _1934_ (.A1(_1070_),
    .A2(_1071_),
    .Y(_1072_),
    .B1(_1066_));
 sg13g2_o21ai_1 _1935_ (.B1(_1072_),
    .Y(_1073_),
    .A1(_1062_),
    .A2(_1065_));
 sg13g2_and2_1 _1936_ (.A(net445),
    .B(_1066_),
    .X(_1074_));
 sg13g2_inv_1 _1937_ (.Y(_1075_),
    .A(_1074_));
 sg13g2_nor2_1 _1938_ (.A(_0958_),
    .B(net415),
    .Y(_1076_));
 sg13g2_nor2_1 _1939_ (.A(net415),
    .B(_1057_),
    .Y(_1077_));
 sg13g2_mux2_1 _1940_ (.A0(net449),
    .A1(net464),
    .S(_1077_),
    .X(_1078_));
 sg13g2_o21ai_1 _1941_ (.B1(_1074_),
    .Y(_1079_),
    .A1(_1076_),
    .A2(_1078_));
 sg13g2_nand3_1 _1942_ (.B(net453),
    .C(_1027_),
    .A(_0894_),
    .Y(_1080_));
 sg13g2_nor2b_1 _1943_ (.A(_1028_),
    .B_N(_1080_),
    .Y(_1081_));
 sg13g2_nand2b_1 _1944_ (.Y(_1082_),
    .B(_1080_),
    .A_N(_1028_));
 sg13g2_nor2_1 _1945_ (.A(net453),
    .B(net445),
    .Y(_1083_));
 sg13g2_inv_1 _1946_ (.Y(_1084_),
    .A(_1083_));
 sg13g2_and2_1 _1947_ (.A(net464),
    .B(_1038_),
    .X(_1085_));
 sg13g2_nor2_1 _1948_ (.A(_0946_),
    .B(_0974_),
    .Y(_1086_));
 sg13g2_nor3_1 _1949_ (.A(_1055_),
    .B(_1085_),
    .C(_1086_),
    .Y(_1087_));
 sg13g2_o21ai_1 _1950_ (.B1(_1082_),
    .Y(_1088_),
    .A1(_1084_),
    .A2(_1087_));
 sg13g2_nor2b_1 _1951_ (.A(_1088_),
    .B_N(_1079_),
    .Y(_1089_));
 sg13g2_nor3_1 _1952_ (.A(net462),
    .B(_1034_),
    .C(_1043_),
    .Y(_1090_));
 sg13g2_nor2_1 _1953_ (.A(_1064_),
    .B(_1090_),
    .Y(_1091_));
 sg13g2_a21o_1 _1954_ (.A2(_1091_),
    .A1(_1067_),
    .B1(_1062_),
    .X(_1092_));
 sg13g2_a21oi_1 _1955_ (.A1(_0910_),
    .A2(_1049_),
    .Y(_1093_),
    .B1(_1057_));
 sg13g2_a21o_1 _1956_ (.A2(_1093_),
    .A1(_1051_),
    .B1(_0970_),
    .X(_1094_));
 sg13g2_nand4_1 _1957_ (.B(_1040_),
    .C(_1051_),
    .A(net464),
    .Y(_1095_),
    .D(_1052_));
 sg13g2_o21ai_1 _1958_ (.B1(_1095_),
    .Y(_1096_),
    .A1(_1053_),
    .A2(_1069_));
 sg13g2_o21ai_1 _1959_ (.B1(_1094_),
    .Y(_1097_),
    .A1(net449),
    .A2(_1096_));
 sg13g2_nand2_1 _1960_ (.Y(_1098_),
    .A(_1085_),
    .B(_1093_));
 sg13g2_a21oi_1 _1961_ (.A1(_1069_),
    .A2(_1098_),
    .Y(_1099_),
    .B1(net415));
 sg13g2_nand4_1 _1962_ (.B(net464),
    .C(_1040_),
    .A(net484),
    .Y(_1100_),
    .D(_1051_));
 sg13g2_and2_1 _1963_ (.A(net461),
    .B(_1038_),
    .X(_1101_));
 sg13g2_nand3_1 _1964_ (.B(_1038_),
    .C(_1052_),
    .A(_0972_),
    .Y(_1102_));
 sg13g2_nand3b_1 _1965_ (.B(_1100_),
    .C(_1102_),
    .Y(_1103_),
    .A_N(net445));
 sg13g2_a21o_1 _1966_ (.A2(_1099_),
    .A1(net449),
    .B1(_1103_),
    .X(_1104_));
 sg13g2_a21oi_1 _1967_ (.A1(_1063_),
    .A2(_1097_),
    .Y(_1105_),
    .B1(_1066_));
 sg13g2_a21oi_1 _1968_ (.A1(net461),
    .A2(_1061_),
    .Y(_1106_),
    .B1(net415));
 sg13g2_o21ai_1 _1969_ (.B1(_1067_),
    .Y(_1107_),
    .A1(net449),
    .A2(_1106_));
 sg13g2_o21ai_1 _1970_ (.B1(_1081_),
    .Y(_1108_),
    .A1(_1084_),
    .A2(_1107_));
 sg13g2_a221oi_1 _1971_ (.B2(_1105_),
    .C1(_1108_),
    .B1(_1104_),
    .A1(_1074_),
    .Y(_1109_),
    .A2(_1092_));
 sg13g2_a21oi_1 _1972_ (.A1(_1073_),
    .A2(_1089_),
    .Y(_1110_),
    .B1(_1109_));
 sg13g2_and2_1 _1973_ (.A(_1029_),
    .B(_1082_),
    .X(_1111_));
 sg13g2_o21ai_1 _1974_ (.B1(net449),
    .Y(_1112_),
    .A1(_1055_),
    .A2(_1085_));
 sg13g2_nor3_1 _1975_ (.A(net445),
    .B(_1068_),
    .C(_1076_),
    .Y(_1113_));
 sg13g2_nor2_1 _1976_ (.A(net461),
    .B(_1057_),
    .Y(_1114_));
 sg13g2_o21ai_1 _1977_ (.B1(net449),
    .Y(_1115_),
    .A1(_1055_),
    .A2(_1114_));
 sg13g2_a22oi_1 _1978_ (.Y(_1116_),
    .B1(_1060_),
    .B2(_0952_),
    .A2(_1041_),
    .A1(_0972_));
 sg13g2_and2_1 _1979_ (.A(net445),
    .B(_1116_),
    .X(_1117_));
 sg13g2_a22oi_1 _1980_ (.Y(_1118_),
    .B1(_1115_),
    .B2(_1117_),
    .A2(_1113_),
    .A1(_1112_));
 sg13g2_o21ai_1 _1981_ (.B1(_0951_),
    .Y(_1119_),
    .A1(_1068_),
    .A2(_1101_));
 sg13g2_nand4_1 _1982_ (.B(_1056_),
    .C(_1083_),
    .A(_0973_),
    .Y(_1120_),
    .D(_1119_));
 sg13g2_o21ai_1 _1983_ (.B1(_1120_),
    .Y(_1121_),
    .A1(_1066_),
    .A2(_1118_));
 sg13g2_o21ai_1 _1984_ (.B1(_1116_),
    .Y(_1122_),
    .A1(_0974_),
    .A2(_1061_));
 sg13g2_nand3_1 _1985_ (.B(_1038_),
    .C(_1060_),
    .A(net449),
    .Y(_1123_));
 sg13g2_a21oi_1 _1986_ (.A1(_1116_),
    .A2(_1123_),
    .Y(_1124_),
    .B1(_1063_));
 sg13g2_nor3_1 _1987_ (.A(net464),
    .B(_1042_),
    .C(_1059_),
    .Y(_1125_));
 sg13g2_o21ai_1 _1988_ (.B1(net445),
    .Y(_1126_),
    .A1(_1114_),
    .A2(_1125_));
 sg13g2_nand3b_1 _1989_ (.B(_1068_),
    .C(_1083_),
    .Y(_1127_),
    .A_N(net415));
 sg13g2_nand2_1 _1990_ (.Y(_1128_),
    .A(_1074_),
    .B(_1122_));
 sg13g2_nand4_1 _1991_ (.B(_0970_),
    .C(_1081_),
    .A(_0906_),
    .Y(_1129_),
    .D(_1128_));
 sg13g2_nand2b_1 _1992_ (.Y(_1130_),
    .B(_0958_),
    .A_N(net415));
 sg13g2_nand3_1 _1993_ (.B(_0967_),
    .C(_1130_),
    .A(net461),
    .Y(_1131_));
 sg13g2_nor2_1 _1994_ (.A(_1066_),
    .B(_1124_),
    .Y(_1132_));
 sg13g2_a22oi_1 _1995_ (.Y(_1133_),
    .B1(_1132_),
    .B2(_1126_),
    .A2(_1131_),
    .A1(_1066_));
 sg13g2_nor2_1 _1996_ (.A(_1129_),
    .B(_1133_),
    .Y(_1134_));
 sg13g2_a22oi_1 _1997_ (.Y(_1135_),
    .B1(_1127_),
    .B2(_1134_),
    .A2(_1121_),
    .A1(_1111_));
 sg13g2_o21ai_1 _1998_ (.B1(_1135_),
    .Y(_1136_),
    .A1(_1029_),
    .A2(_1110_));
 sg13g2_a21oi_1 _1999_ (.A1(_0972_),
    .A2(_0991_),
    .Y(_1137_),
    .B1(_1075_));
 sg13g2_o21ai_1 _2000_ (.B1(_1137_),
    .Y(_1138_),
    .A1(_0972_),
    .A2(_1111_));
 sg13g2_nor3_1 _2001_ (.A(_0894_),
    .B(net452),
    .C(_0906_),
    .Y(_1139_));
 sg13g2_xor2_1 _2002_ (.B(_1139_),
    .A(_0994_),
    .X(_1140_));
 sg13g2_nor3_1 _2003_ (.A(_1030_),
    .B(_1034_),
    .C(_1140_),
    .Y(_1141_));
 sg13g2_nand3_1 _2004_ (.B(_1138_),
    .C(_1141_),
    .A(_1136_),
    .Y(_1142_));
 sg13g2_nor2_2 _2005_ (.A(_0860_),
    .B(net466),
    .Y(_1143_));
 sg13g2_nand2_1 _2006_ (.Y(_1144_),
    .A(net485),
    .B(net489));
 sg13g2_a21oi_2 _2007_ (.B1(_0862_),
    .Y(_1145_),
    .A2(net459),
    .A1(_0861_));
 sg13g2_xor2_1 _2008_ (.B(_1145_),
    .A(_0017_),
    .X(_1146_));
 sg13g2_and2_2 _2009_ (.A(net505),
    .B(net508),
    .X(_1147_));
 sg13g2_nand2_1 _2010_ (.Y(_1148_),
    .A(net506),
    .B(net509));
 sg13g2_and2_2 _2011_ (.A(net501),
    .B(net506),
    .X(_1149_));
 sg13g2_nand2_2 _2012_ (.Y(_1150_),
    .A(net502),
    .B(net506));
 sg13g2_nor2_2 _2013_ (.A(_0912_),
    .B(_1149_),
    .Y(_1151_));
 sg13g2_nand2b_2 _2014_ (.Y(_1152_),
    .B(_1150_),
    .A_N(_0912_));
 sg13g2_nand2_1 _2015_ (.Y(_1153_),
    .A(_0919_),
    .B(_1150_));
 sg13g2_a21o_2 _2016_ (.A2(_1150_),
    .A1(_0919_),
    .B1(_0022_),
    .X(_1154_));
 sg13g2_nand3_1 _2017_ (.B(_0919_),
    .C(_1150_),
    .A(_0022_),
    .Y(_1155_));
 sg13g2_nand3b_1 _2018_ (.B(_1150_),
    .C(_0028_),
    .Y(_1156_),
    .A_N(_0012_));
 sg13g2_o21ai_1 _2019_ (.B1(_0012_),
    .Y(_1157_),
    .A1(_0865_),
    .A2(_1149_));
 sg13g2_and2_1 _2020_ (.A(_1156_),
    .B(_1157_),
    .X(_1158_));
 sg13g2_a22oi_1 _2021_ (.Y(_1159_),
    .B1(_1156_),
    .B2(_1157_),
    .A2(_1155_),
    .A1(_1154_));
 sg13g2_xnor2_1 _2022_ (.Y(_1160_),
    .A(net499),
    .B(_1149_));
 sg13g2_a221oi_1 _2023_ (.B2(_1157_),
    .C1(_1160_),
    .B1(_1156_),
    .A1(_1154_),
    .Y(_1161_),
    .A2(_1155_));
 sg13g2_nand3_1 _2024_ (.B(_1152_),
    .C(_1161_),
    .A(_1147_),
    .Y(_1162_));
 sg13g2_a221oi_1 _2025_ (.B2(_1157_),
    .C1(_0873_),
    .B1(_1156_),
    .A1(_1154_),
    .Y(_1163_),
    .A2(_1155_));
 sg13g2_and2_1 _2026_ (.A(net499),
    .B(_1151_),
    .X(_1164_));
 sg13g2_nand3_1 _2027_ (.B(_1159_),
    .C(_1164_),
    .A(_1147_),
    .Y(_1165_));
 sg13g2_nor2b_2 _2028_ (.A(net508),
    .B_N(net505),
    .Y(_1166_));
 sg13g2_nand3_1 _2029_ (.B(_1164_),
    .C(_1166_),
    .A(_1159_),
    .Y(_1167_));
 sg13g2_nand3_1 _2030_ (.B(_1159_),
    .C(_1164_),
    .A(net505),
    .Y(_1168_));
 sg13g2_nand3_1 _2031_ (.B(_0858_),
    .C(_1159_),
    .A(net499),
    .Y(_1169_));
 sg13g2_nand2_1 _2032_ (.Y(_1170_),
    .A(_1162_),
    .B(_1169_));
 sg13g2_or2_2 _2033_ (.X(_1171_),
    .B(_1170_),
    .A(_1163_));
 sg13g2_nand2_2 _2034_ (.Y(_1172_),
    .A(_0913_),
    .B(_1163_));
 sg13g2_a21oi_2 _2035_ (.B1(net491),
    .Y(_1173_),
    .A2(_1163_),
    .A1(_0913_));
 sg13g2_nand2_1 _2036_ (.Y(_1174_),
    .A(_1171_),
    .B(_1173_));
 sg13g2_nor2_2 _2037_ (.A(_0888_),
    .B(_1143_),
    .Y(_1175_));
 sg13g2_nand2_2 _2038_ (.Y(_1176_),
    .A(_0889_),
    .B(net459));
 sg13g2_nand3_1 _2039_ (.B(_1169_),
    .C(_1172_),
    .A(_1162_),
    .Y(_1177_));
 sg13g2_nand4_1 _2040_ (.B(_1162_),
    .C(_1163_),
    .A(_0914_),
    .Y(_1178_),
    .D(_1169_));
 sg13g2_nor2_1 _2041_ (.A(_0020_),
    .B(_1176_),
    .Y(_1179_));
 sg13g2_nand2_1 _2042_ (.Y(_1180_),
    .A(_0023_),
    .B(net459));
 sg13g2_xnor2_1 _2043_ (.Y(_1181_),
    .A(_0862_),
    .B(_1180_));
 sg13g2_xnor2_1 _2044_ (.Y(_1182_),
    .A(net481),
    .B(_1180_));
 sg13g2_nor2_1 _2045_ (.A(net468),
    .B(net482),
    .Y(_1183_));
 sg13g2_xnor2_1 _2046_ (.Y(_1184_),
    .A(_0861_),
    .B(net459));
 sg13g2_xnor2_1 _2047_ (.Y(_1185_),
    .A(net483),
    .B(net459));
 sg13g2_nor2_1 _2048_ (.A(_1182_),
    .B(_1185_),
    .Y(_1186_));
 sg13g2_or2_1 _2049_ (.X(_1187_),
    .B(_1168_),
    .A(net491));
 sg13g2_a21oi_1 _2050_ (.A1(_1175_),
    .A2(_1187_),
    .Y(_1188_),
    .B1(net456));
 sg13g2_nand3_1 _2051_ (.B(_0912_),
    .C(_1161_),
    .A(net508),
    .Y(_1189_));
 sg13g2_and2_1 _2052_ (.A(_1172_),
    .B(net448),
    .X(_1190_));
 sg13g2_nand3_1 _2053_ (.B(_1147_),
    .C(_1159_),
    .A(_0872_),
    .Y(_1191_));
 sg13g2_nand3_1 _2054_ (.B(_1190_),
    .C(_1191_),
    .A(net491),
    .Y(_1192_));
 sg13g2_nand2_1 _2055_ (.Y(_1193_),
    .A(_1148_),
    .B(_1163_));
 sg13g2_nand4_1 _2056_ (.B(_1168_),
    .C(net448),
    .A(net467),
    .Y(_1194_),
    .D(_1193_));
 sg13g2_nand3_1 _2057_ (.B(_1192_),
    .C(_1194_),
    .A(_1188_),
    .Y(_1195_));
 sg13g2_nand2_1 _2058_ (.Y(_1196_),
    .A(_1187_),
    .B(_1190_));
 sg13g2_o21ai_1 _2059_ (.B1(_1184_),
    .Y(_1197_),
    .A1(_1175_),
    .A2(_1196_));
 sg13g2_o21ai_1 _2060_ (.B1(_1175_),
    .Y(_1198_),
    .A1(_0020_),
    .A2(_1172_));
 sg13g2_nand2b_1 _2061_ (.Y(_1199_),
    .B(_1198_),
    .A_N(_1197_));
 sg13g2_nand3_1 _2062_ (.B(_1195_),
    .C(_1199_),
    .A(_1182_),
    .Y(_1200_));
 sg13g2_nand3_1 _2063_ (.B(_1172_),
    .C(net448),
    .A(_1168_),
    .Y(_1201_));
 sg13g2_inv_1 _2064_ (.Y(_1202_),
    .A(_1201_));
 sg13g2_nand3_1 _2065_ (.B(_1178_),
    .C(_1184_),
    .A(_1174_),
    .Y(_1203_));
 sg13g2_a21oi_1 _2066_ (.A1(net467),
    .A2(_1167_),
    .Y(_1204_),
    .B1(net456));
 sg13g2_nand2_1 _2067_ (.Y(_1205_),
    .A(_1201_),
    .B(_1204_));
 sg13g2_a21oi_1 _2068_ (.A1(_1203_),
    .A2(_1205_),
    .Y(_1206_),
    .B1(_1175_));
 sg13g2_nand3_1 _2069_ (.B(_1170_),
    .C(net456),
    .A(_0873_),
    .Y(_1207_));
 sg13g2_o21ai_1 _2070_ (.B1(_1207_),
    .Y(_1208_),
    .A1(net456),
    .A2(_1189_));
 sg13g2_a21o_1 _2071_ (.A2(_1208_),
    .A1(_1179_),
    .B1(_1182_),
    .X(_1209_));
 sg13g2_o21ai_1 _2072_ (.B1(_1200_),
    .Y(_1210_),
    .A1(_1206_),
    .A2(_1209_));
 sg13g2_nand3_1 _2073_ (.B(_1171_),
    .C(_1190_),
    .A(net491),
    .Y(_1211_));
 sg13g2_nand4_1 _2074_ (.B(_0858_),
    .C(_0859_),
    .A(net499),
    .Y(_1212_),
    .D(_1159_));
 sg13g2_nand3_1 _2075_ (.B(_1173_),
    .C(_1212_),
    .A(_1171_),
    .Y(_1213_));
 sg13g2_a21oi_1 _2076_ (.A1(_1211_),
    .A2(_1213_),
    .Y(_1214_),
    .B1(_1176_));
 sg13g2_and2_1 _2077_ (.A(_1162_),
    .B(_1165_),
    .X(_1215_));
 sg13g2_nand2b_1 _2078_ (.Y(_1216_),
    .B(_1215_),
    .A_N(_1169_));
 sg13g2_a221oi_1 _2079_ (.B2(_1143_),
    .C1(_1214_),
    .B1(_1216_),
    .A1(_0888_),
    .Y(_1217_),
    .A2(_1215_));
 sg13g2_a21oi_1 _2080_ (.A1(_0912_),
    .A2(_1161_),
    .Y(_1218_),
    .B1(net494));
 sg13g2_a21oi_1 _2081_ (.A1(_1215_),
    .A2(_1218_),
    .Y(_1219_),
    .B1(_1175_));
 sg13g2_nor2_2 _2082_ (.A(net468),
    .B(net492),
    .Y(_1220_));
 sg13g2_nand2_1 _2083_ (.Y(_1221_),
    .A(net498),
    .B(_0914_));
 sg13g2_nand3_1 _2084_ (.B(_1220_),
    .C(_1221_),
    .A(_1171_),
    .Y(_1222_));
 sg13g2_a21oi_1 _2085_ (.A1(_1211_),
    .A2(_1219_),
    .Y(_1223_),
    .B1(_1185_));
 sg13g2_a21oi_1 _2086_ (.A1(_1222_),
    .A2(_1223_),
    .Y(_1224_),
    .B1(_1181_));
 sg13g2_o21ai_1 _2087_ (.B1(_1224_),
    .Y(_1225_),
    .A1(net456),
    .A2(_1217_));
 sg13g2_nand3_1 _2088_ (.B(_1159_),
    .C(_1166_),
    .A(_0872_),
    .Y(_1226_));
 sg13g2_nand3_1 _2089_ (.B(_1168_),
    .C(_1226_),
    .A(net467),
    .Y(_1227_));
 sg13g2_nand2_1 _2090_ (.Y(_1228_),
    .A(net468),
    .B(_1172_));
 sg13g2_a21oi_1 _2091_ (.A1(_1227_),
    .A2(_1228_),
    .Y(_1229_),
    .B1(_1176_));
 sg13g2_nand3_1 _2092_ (.B(_1168_),
    .C(_1171_),
    .A(net467),
    .Y(_1230_));
 sg13g2_nand3_1 _2093_ (.B(_1211_),
    .C(_1230_),
    .A(_1188_),
    .Y(_1231_));
 sg13g2_o21ai_1 _2094_ (.B1(_1231_),
    .Y(_1232_),
    .A1(_1197_),
    .A2(_1229_));
 sg13g2_a21oi_1 _2095_ (.A1(_1181_),
    .A2(_1232_),
    .Y(_1233_),
    .B1(_1146_));
 sg13g2_a22oi_1 _2096_ (.Y(_1234_),
    .B1(_1225_),
    .B2(_1233_),
    .A2(_1210_),
    .A1(_1146_));
 sg13g2_nor2_1 _2097_ (.A(net478),
    .B(_1145_),
    .Y(_1235_));
 sg13g2_xnor2_1 _2098_ (.Y(_1236_),
    .A(_0016_),
    .B(_1235_));
 sg13g2_xor2_1 _2099_ (.B(_1235_),
    .A(_0016_),
    .X(_1237_));
 sg13g2_a21oi_1 _2100_ (.A1(net467),
    .A2(net448),
    .Y(_1238_),
    .B1(_1175_));
 sg13g2_o21ai_1 _2101_ (.B1(_1175_),
    .Y(_1239_),
    .A1(_1173_),
    .A2(_1202_));
 sg13g2_a22oi_1 _2102_ (.Y(_1240_),
    .B1(_1190_),
    .B2(_0888_),
    .A2(_1168_),
    .A1(_1143_));
 sg13g2_nor2_1 _2103_ (.A(net487),
    .B(net466),
    .Y(_1241_));
 sg13g2_nand3_1 _2104_ (.B(net459),
    .C(_1181_),
    .A(net483),
    .Y(_1242_));
 sg13g2_a221oi_1 _2105_ (.B2(_1167_),
    .C1(_1242_),
    .B1(_1241_),
    .A1(net448),
    .Y(_1243_),
    .A2(_1220_));
 sg13g2_o21ai_1 _2106_ (.B1(_1243_),
    .Y(_1244_),
    .A1(_0889_),
    .A2(_1201_));
 sg13g2_a21oi_1 _2107_ (.A1(_1239_),
    .A2(_1240_),
    .Y(_1245_),
    .B1(_1185_));
 sg13g2_a221oi_1 _2108_ (.B2(_1178_),
    .C1(net456),
    .B1(_1238_),
    .A1(_1179_),
    .Y(_1246_),
    .A2(_1201_));
 sg13g2_or2_1 _2109_ (.X(_1247_),
    .B(_1246_),
    .A(_1181_));
 sg13g2_o21ai_1 _2110_ (.B1(_1244_),
    .Y(_1248_),
    .A1(_1245_),
    .A2(_1247_));
 sg13g2_a21oi_1 _2111_ (.A1(_1172_),
    .A2(net448),
    .Y(_1249_),
    .B1(net488));
 sg13g2_a21oi_1 _2112_ (.A1(_1167_),
    .A2(_1185_),
    .Y(_1250_),
    .B1(net488));
 sg13g2_nor3_1 _2113_ (.A(_1176_),
    .B(_1249_),
    .C(_1250_),
    .Y(_1251_));
 sg13g2_a21oi_1 _2114_ (.A1(_1168_),
    .A2(net448),
    .Y(_1252_),
    .B1(_0888_));
 sg13g2_o21ai_1 _2115_ (.B1(net456),
    .Y(_1253_),
    .A1(_0889_),
    .A2(_1172_));
 sg13g2_nor2_1 _2116_ (.A(_1252_),
    .B(_1253_),
    .Y(_1254_));
 sg13g2_o21ai_1 _2117_ (.B1(_1240_),
    .Y(_1255_),
    .A1(_1176_),
    .A2(_1249_));
 sg13g2_nor2_1 _2118_ (.A(_1251_),
    .B(_1254_),
    .Y(_1256_));
 sg13g2_o21ai_1 _2119_ (.B1(_1256_),
    .Y(_1257_),
    .A1(net456),
    .A2(_1240_));
 sg13g2_nand3_1 _2120_ (.B(_1171_),
    .C(net448),
    .A(net467),
    .Y(_1258_));
 sg13g2_and2_1 _2121_ (.A(_1143_),
    .B(_1177_),
    .X(_1259_));
 sg13g2_o21ai_1 _2122_ (.B1(_1258_),
    .Y(_1260_),
    .A1(_0888_),
    .A2(_1259_));
 sg13g2_nand2_1 _2123_ (.Y(_1261_),
    .A(_1177_),
    .B(_1179_));
 sg13g2_nand4_1 _2124_ (.B(_1185_),
    .C(_1260_),
    .A(_1181_),
    .Y(_1262_),
    .D(_1261_));
 sg13g2_a221oi_1 _2125_ (.B2(_1182_),
    .C1(_1146_),
    .B1(_1257_),
    .A1(_1186_),
    .Y(_1263_),
    .A2(_1255_));
 sg13g2_a221oi_1 _2126_ (.B2(_1263_),
    .C1(_1237_),
    .B1(_1262_),
    .A1(_1146_),
    .Y(_1264_),
    .A2(_1248_));
 sg13g2_nor2b_1 _2127_ (.A(_1145_),
    .B_N(_0992_),
    .Y(_1265_));
 sg13g2_xnor2_1 _2128_ (.Y(_1266_),
    .A(_0015_),
    .B(_1265_));
 sg13g2_o21ai_1 _2129_ (.B1(_1159_),
    .Y(_1267_),
    .A1(net499),
    .A2(_1149_));
 sg13g2_nor3_1 _2130_ (.A(_1264_),
    .B(_1266_),
    .C(_1267_),
    .Y(_1268_));
 sg13g2_o21ai_1 _2131_ (.B1(_1268_),
    .Y(_1269_),
    .A1(_1234_),
    .A2(_1236_));
 sg13g2_xnor2_1 _2132_ (.Y(_1270_),
    .A(_0016_),
    .B(_0885_));
 sg13g2_inv_1 _2133_ (.Y(_1271_),
    .A(_1270_));
 sg13g2_nor2_1 _2134_ (.A(net498),
    .B(_1152_),
    .Y(_1272_));
 sg13g2_nand3_1 _2135_ (.B(net497),
    .C(_0872_),
    .A(_0857_),
    .Y(_1273_));
 sg13g2_nor4_2 _2136_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[8] ),
    .B(net500),
    .C(net497),
    .Y(_1274_),
    .D(_1152_));
 sg13g2_nand2_1 _2137_ (.Y(_1275_),
    .A(_0913_),
    .B(_1274_));
 sg13g2_inv_1 _2138_ (.Y(_1276_),
    .A(_1275_));
 sg13g2_nand4_1 _2139_ (.B(net497),
    .C(_0872_),
    .A(_0857_),
    .Y(_1277_),
    .D(_0875_));
 sg13g2_nor4_2 _2140_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[8] ),
    .B(net498),
    .C(net501),
    .Y(_1278_),
    .D(net497));
 sg13g2_or4_2 _2141_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[8] ),
    .B(net498),
    .C(net501),
    .D(net497),
    .X(_1279_));
 sg13g2_nand4_1 _2142_ (.B(net505),
    .C(net497),
    .A(_0857_),
    .Y(_1280_),
    .D(_0872_));
 sg13g2_and4_2 _2143_ (.A(_1275_),
    .B(_1277_),
    .C(_1279_),
    .D(_1280_),
    .X(_1281_));
 sg13g2_nor2_2 _2144_ (.A(net498),
    .B(_1281_),
    .Y(_1282_));
 sg13g2_nor2_2 _2145_ (.A(_0877_),
    .B(_0882_),
    .Y(_1283_));
 sg13g2_nand2_2 _2146_ (.Y(_1284_),
    .A(_0878_),
    .B(_0883_));
 sg13g2_nand2_1 _2147_ (.Y(_1285_),
    .A(_1166_),
    .B(_1278_));
 sg13g2_nor2_1 _2148_ (.A(net489),
    .B(_1285_),
    .Y(_1286_));
 sg13g2_nor2_1 _2149_ (.A(_1283_),
    .B(_1286_),
    .Y(_1287_));
 sg13g2_and2_1 _2150_ (.A(_0875_),
    .B(_1278_),
    .X(_1288_));
 sg13g2_nand2_1 _2151_ (.Y(_1289_),
    .A(_0875_),
    .B(_1278_));
 sg13g2_a22oi_1 _2152_ (.Y(_1290_),
    .B1(_1288_),
    .B2(net490),
    .A2(_1282_),
    .A1(_1220_));
 sg13g2_xor2_1 _2153_ (.B(_0884_),
    .A(_0017_),
    .X(_1291_));
 sg13g2_o21ai_1 _2154_ (.B1(_0913_),
    .Y(_1292_),
    .A1(_1274_),
    .A2(_1278_));
 sg13g2_nand2_1 _2155_ (.Y(_1293_),
    .A(_1285_),
    .B(_1292_));
 sg13g2_o21ai_1 _2156_ (.B1(net482),
    .Y(_1294_),
    .A1(net489),
    .A2(_1292_));
 sg13g2_nand2_1 _2157_ (.Y(_1295_),
    .A(_1293_),
    .B(_1294_));
 sg13g2_xor2_1 _2158_ (.B(_0882_),
    .A(_0018_),
    .X(_1296_));
 sg13g2_nand2_1 _2159_ (.Y(_1297_),
    .A(net489),
    .B(_1292_));
 sg13g2_a21oi_1 _2160_ (.A1(net490),
    .A2(_1292_),
    .Y(_1298_),
    .B1(net485));
 sg13g2_nor3_1 _2161_ (.A(net468),
    .B(net488),
    .C(_1292_),
    .Y(_1299_));
 sg13g2_a21oi_1 _2162_ (.A1(_1282_),
    .A2(_1298_),
    .Y(_1300_),
    .B1(_1299_));
 sg13g2_a21oi_1 _2163_ (.A1(_0913_),
    .A2(_1278_),
    .Y(_1301_),
    .B1(net489));
 sg13g2_nand3_1 _2164_ (.B(_1277_),
    .C(_1301_),
    .A(_1275_),
    .Y(_1302_));
 sg13g2_o21ai_1 _2165_ (.B1(_1302_),
    .Y(_1303_),
    .A1(_1281_),
    .A2(_1297_));
 sg13g2_nand2_1 _2166_ (.Y(_1304_),
    .A(_1147_),
    .B(_1278_));
 sg13g2_a21oi_2 _2167_ (.B1(net466),
    .Y(_1305_),
    .A2(_1278_),
    .A1(_1166_));
 sg13g2_a22oi_1 _2168_ (.Y(_1306_),
    .B1(_1305_),
    .B2(_1289_),
    .A2(_1304_),
    .A1(_1301_));
 sg13g2_nor4_1 _2169_ (.A(net485),
    .B(_0861_),
    .C(_1281_),
    .D(_1306_),
    .Y(_1307_));
 sg13g2_o21ai_1 _2170_ (.B1(_1280_),
    .Y(_1308_),
    .A1(_1147_),
    .A2(_1279_));
 sg13g2_nor2_1 _2171_ (.A(_1144_),
    .B(_1308_),
    .Y(_1309_));
 sg13g2_nor3_1 _2172_ (.A(_1276_),
    .B(_1281_),
    .C(_1308_),
    .Y(_1310_));
 sg13g2_nor2b_1 _2173_ (.A(_1310_),
    .B_N(_1220_),
    .Y(_1311_));
 sg13g2_nor3_1 _2174_ (.A(net498),
    .B(net488),
    .C(_1281_),
    .Y(_1312_));
 sg13g2_a221oi_1 _2175_ (.B2(_1274_),
    .C1(_1281_),
    .B1(_0913_),
    .A1(_0861_),
    .Y(_1313_),
    .A2(net488));
 sg13g2_o21ai_1 _2176_ (.B1(_1284_),
    .Y(_1314_),
    .A1(_0877_),
    .A2(_1312_));
 sg13g2_or3_1 _2177_ (.A(_1309_),
    .B(_1311_),
    .C(_1314_),
    .X(_1315_));
 sg13g2_o21ai_1 _2178_ (.B1(_1315_),
    .Y(_1316_),
    .A1(_1284_),
    .A2(_1313_));
 sg13g2_o21ai_1 _2179_ (.B1(net466),
    .Y(_1317_),
    .A1(_0913_),
    .A2(_1279_));
 sg13g2_a22oi_1 _2180_ (.Y(_1318_),
    .B1(_1298_),
    .B2(_1317_),
    .A2(_1282_),
    .A1(_1220_));
 sg13g2_nand2b_1 _2181_ (.Y(_1319_),
    .B(_0882_),
    .A_N(net488));
 sg13g2_a21oi_1 _2182_ (.A1(_1275_),
    .A2(_1280_),
    .Y(_1320_),
    .B1(_1319_));
 sg13g2_nor3_1 _2183_ (.A(net466),
    .B(_0913_),
    .C(_1279_),
    .Y(_1321_));
 sg13g2_nor2_1 _2184_ (.A(net468),
    .B(_1321_),
    .Y(_1322_));
 sg13g2_o21ai_1 _2185_ (.B1(_1322_),
    .Y(_1323_),
    .A1(net490),
    .A2(_1292_));
 sg13g2_o21ai_1 _2186_ (.B1(_1323_),
    .Y(_1324_),
    .A1(_0877_),
    .A2(_1320_));
 sg13g2_a221oi_1 _2187_ (.B2(_1283_),
    .C1(_1296_),
    .B1(_1295_),
    .A1(_1287_),
    .Y(_1325_),
    .A2(_1290_));
 sg13g2_a21oi_1 _2188_ (.A1(_1296_),
    .A2(_1316_),
    .Y(_1326_),
    .B1(_1325_));
 sg13g2_o21ai_1 _2189_ (.B1(_1324_),
    .Y(_1327_),
    .A1(_1284_),
    .A2(_1318_));
 sg13g2_or2_1 _2190_ (.X(_1328_),
    .B(_1307_),
    .A(_1296_));
 sg13g2_a221oi_1 _2191_ (.B2(_1183_),
    .C1(_1328_),
    .B1(_1303_),
    .A1(_1284_),
    .Y(_1329_),
    .A2(_1300_));
 sg13g2_a21oi_1 _2192_ (.A1(_1296_),
    .A2(_1327_),
    .Y(_1330_),
    .B1(_1329_));
 sg13g2_mux2_1 _2193_ (.A0(_1326_),
    .A1(_1330_),
    .S(_1291_),
    .X(_1331_));
 sg13g2_a21o_1 _2194_ (.A2(_1289_),
    .A1(net466),
    .B1(_1305_),
    .X(_1332_));
 sg13g2_o21ai_1 _2195_ (.B1(_1296_),
    .Y(_1333_),
    .A1(_0878_),
    .A2(_1312_));
 sg13g2_a221oi_1 _2196_ (.B2(_0882_),
    .C1(_1333_),
    .B1(_1332_),
    .A1(_1283_),
    .Y(_1334_),
    .A2(_1300_));
 sg13g2_a21oi_1 _2197_ (.A1(net459),
    .A2(_1282_),
    .Y(_1335_),
    .B1(_1284_));
 sg13g2_o21ai_1 _2198_ (.B1(_1292_),
    .Y(_1336_),
    .A1(_1287_),
    .A2(_1305_));
 sg13g2_a21oi_1 _2199_ (.A1(net484),
    .A2(_1284_),
    .Y(_1337_),
    .B1(_1296_));
 sg13g2_nand2_1 _2200_ (.Y(_1338_),
    .A(_1336_),
    .B(_1337_));
 sg13g2_o21ai_1 _2201_ (.B1(_1270_),
    .Y(_1339_),
    .A1(_1335_),
    .A2(_1338_));
 sg13g2_a21oi_1 _2202_ (.A1(_0018_),
    .A2(_0882_),
    .Y(_1340_),
    .B1(_1291_));
 sg13g2_xnor2_1 _2203_ (.Y(_1341_),
    .A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[9] ),
    .B(_0886_));
 sg13g2_o21ai_1 _2204_ (.B1(_1341_),
    .Y(_1342_),
    .A1(_1271_),
    .A2(_1340_));
 sg13g2_a21oi_1 _2205_ (.A1(_1273_),
    .A2(_1281_),
    .Y(_1343_),
    .B1(_1342_));
 sg13g2_o21ai_1 _2206_ (.B1(_1343_),
    .Y(_1344_),
    .A1(_1334_),
    .A2(_1339_));
 sg13g2_a21oi_1 _2207_ (.A1(_1271_),
    .A2(_1331_),
    .Y(_1345_),
    .B1(_1344_));
 sg13g2_xnor2_1 _2208_ (.Y(_1346_),
    .A(net480),
    .B(_0878_));
 sg13g2_xnor2_1 _2209_ (.Y(_1347_),
    .A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[7] ),
    .B(net500));
 sg13g2_xor2_1 _2210_ (.B(net501),
    .A(net498),
    .X(_1348_));
 sg13g2_o21ai_1 _2211_ (.B1(_1221_),
    .Y(_1349_),
    .A1(_0914_),
    .A2(_1348_));
 sg13g2_and4_1 _2212_ (.A(_1154_),
    .B(_1155_),
    .C(_1347_),
    .D(_1349_),
    .X(_1350_));
 sg13g2_nand4_1 _2213_ (.B(_1155_),
    .C(_1347_),
    .A(_1154_),
    .Y(_1351_),
    .D(_1349_));
 sg13g2_nand2_1 _2214_ (.Y(_1352_),
    .A(_0021_),
    .B(_1350_));
 sg13g2_nand3_1 _2215_ (.B(_1147_),
    .C(_1350_),
    .A(_0021_),
    .Y(_1353_));
 sg13g2_nor2_2 _2216_ (.A(_0021_),
    .B(_1351_),
    .Y(_1354_));
 sg13g2_nand2b_1 _2217_ (.Y(_1355_),
    .B(_1350_),
    .A_N(_0021_));
 sg13g2_nand2_1 _2218_ (.Y(_1356_),
    .A(net505),
    .B(_1354_));
 sg13g2_a21o_1 _2219_ (.A2(_1356_),
    .A1(_1353_),
    .B1(net493),
    .X(_1357_));
 sg13g2_nor2_2 _2220_ (.A(_1147_),
    .B(_1355_),
    .Y(_1358_));
 sg13g2_inv_1 _2221_ (.Y(_1359_),
    .A(_1358_));
 sg13g2_a21oi_1 _2222_ (.A1(net493),
    .A2(_1358_),
    .Y(_1360_),
    .B1(net486));
 sg13g2_nand3b_1 _2223_ (.B(net466),
    .C(_1354_),
    .Y(_1361_),
    .A_N(net505));
 sg13g2_o21ai_1 _2224_ (.B1(_1353_),
    .Y(_1362_),
    .A1(_0859_),
    .A2(_1355_));
 sg13g2_or2_1 _2225_ (.X(_1363_),
    .B(_1362_),
    .A(_1361_));
 sg13g2_a21oi_1 _2226_ (.A1(_1361_),
    .A2(_1362_),
    .Y(_1364_),
    .B1(net468));
 sg13g2_a22oi_1 _2227_ (.Y(_1365_),
    .B1(_1363_),
    .B2(_1364_),
    .A2(_1360_),
    .A1(_1357_));
 sg13g2_nor2_1 _2228_ (.A(_1284_),
    .B(_1365_),
    .Y(_1366_));
 sg13g2_nand3_1 _2229_ (.B(_1357_),
    .C(_1361_),
    .A(_0877_),
    .Y(_1367_));
 sg13g2_nor2_1 _2230_ (.A(_0018_),
    .B(_0878_),
    .Y(_1368_));
 sg13g2_xor2_1 _2231_ (.B(_1368_),
    .A(_0017_),
    .X(_1369_));
 sg13g2_o21ai_1 _2232_ (.B1(_0882_),
    .Y(_1370_),
    .A1(net488),
    .A2(_1359_));
 sg13g2_nand3_1 _2233_ (.B(_1369_),
    .C(_1370_),
    .A(_1367_),
    .Y(_1371_));
 sg13g2_o21ai_1 _2234_ (.B1(_1346_),
    .Y(_1372_),
    .A1(_1366_),
    .A2(_1371_));
 sg13g2_nand2_1 _2235_ (.Y(_1373_),
    .A(_0021_),
    .B(_0875_));
 sg13g2_inv_1 _2236_ (.Y(_1374_),
    .A(_1373_));
 sg13g2_nor2_1 _2237_ (.A(_1349_),
    .B(_1373_),
    .Y(_1375_));
 sg13g2_nand4_1 _2238_ (.B(_1155_),
    .C(_1347_),
    .A(_1154_),
    .Y(_1376_),
    .D(_1375_));
 sg13g2_o21ai_1 _2239_ (.B1(_1376_),
    .Y(_1377_),
    .A1(_1351_),
    .A2(_1374_));
 sg13g2_nand2_1 _2240_ (.Y(_1378_),
    .A(_0875_),
    .B(_1354_));
 sg13g2_a21oi_1 _2241_ (.A1(_0875_),
    .A2(_1354_),
    .Y(_1379_),
    .B1(net493));
 sg13g2_o21ai_1 _2242_ (.B1(_1377_),
    .Y(_1380_),
    .A1(net486),
    .A2(_1379_));
 sg13g2_o21ai_1 _2243_ (.B1(_1241_),
    .Y(_1381_),
    .A1(net508),
    .A2(_1352_));
 sg13g2_nand3_1 _2244_ (.B(_1376_),
    .C(_1378_),
    .A(_1353_),
    .Y(_1382_));
 sg13g2_xnor2_1 _2245_ (.Y(_1383_),
    .A(_0021_),
    .B(_0914_));
 sg13g2_a21oi_1 _2246_ (.A1(_1349_),
    .A2(_1383_),
    .Y(_1384_),
    .B1(net459));
 sg13g2_nand2b_1 _2247_ (.Y(_1385_),
    .B(_1283_),
    .A_N(_1384_));
 sg13g2_a221oi_1 _2248_ (.B2(_1220_),
    .C1(_1385_),
    .B1(_1382_),
    .A1(_1380_),
    .Y(_1386_),
    .A2(_1381_));
 sg13g2_o21ai_1 _2249_ (.B1(net493),
    .Y(_1387_),
    .A1(_0875_),
    .A2(_1352_));
 sg13g2_nand2b_1 _2250_ (.Y(_1388_),
    .B(_1387_),
    .A_N(_1379_));
 sg13g2_nand3_1 _2251_ (.B(_1357_),
    .C(_1388_),
    .A(net480),
    .Y(_1389_));
 sg13g2_a21oi_1 _2252_ (.A1(net493),
    .A2(_1358_),
    .Y(_1390_),
    .B1(_0883_));
 sg13g2_nand4_1 _2253_ (.B(_1353_),
    .C(_1373_),
    .A(_1350_),
    .Y(_1391_),
    .D(_1390_));
 sg13g2_nand3b_1 _2254_ (.B(_1389_),
    .C(_1391_),
    .Y(_1392_),
    .A_N(_1386_));
 sg13g2_nand3b_1 _2255_ (.B(_1369_),
    .C(_1392_),
    .Y(_1393_),
    .A_N(_1346_));
 sg13g2_xor2_1 _2256_ (.B(_0880_),
    .A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[8] ),
    .X(_1394_));
 sg13g2_a21oi_1 _2257_ (.A1(_1351_),
    .A2(_1376_),
    .Y(_1395_),
    .B1(_1394_));
 sg13g2_a21o_1 _2258_ (.A2(_1362_),
    .A1(net490),
    .B1(net484),
    .X(_1396_));
 sg13g2_nor3_1 _2259_ (.A(net508),
    .B(net488),
    .C(_1355_),
    .Y(_1397_));
 sg13g2_a22oi_1 _2260_ (.Y(_1398_),
    .B1(_1362_),
    .B2(_0861_),
    .A2(_1358_),
    .A1(_1143_));
 sg13g2_a22oi_1 _2261_ (.Y(_1399_),
    .B1(_1398_),
    .B2(_0878_),
    .A2(_1396_),
    .A1(_1283_));
 sg13g2_o21ai_1 _2262_ (.B1(_1399_),
    .Y(_1400_),
    .A1(_0878_),
    .A2(_1397_));
 sg13g2_nand2b_1 _2263_ (.Y(_1401_),
    .B(_1400_),
    .A_N(_1369_));
 sg13g2_nand4_1 _2264_ (.B(_1393_),
    .C(_1395_),
    .A(_1372_),
    .Y(_1402_),
    .D(_1401_));
 sg13g2_nand2_1 _2265_ (.Y(_1403_),
    .A(_1269_),
    .B(_1402_));
 sg13g2_nor2_2 _2266_ (.A(_1345_),
    .B(_1403_),
    .Y(_1404_));
 sg13g2_xnor2_1 _2267_ (.Y(_1405_),
    .A(_0917_),
    .B(_0922_));
 sg13g2_nor2_2 _2268_ (.A(_1033_),
    .B(_1405_),
    .Y(_1406_));
 sg13g2_a221oi_1 _2269_ (.B2(_0959_),
    .C1(_1405_),
    .B1(_1044_),
    .A1(_1031_),
    .Y(_1407_),
    .A2(_1032_));
 sg13g2_a221oi_1 _2270_ (.B2(_0953_),
    .C1(_1405_),
    .B1(_1037_),
    .A1(_1031_),
    .Y(_1408_),
    .A2(_1032_));
 sg13g2_nor4_2 _2271_ (.A(_0917_),
    .B(net455),
    .C(_0925_),
    .Y(_1409_),
    .D(_0980_));
 sg13g2_or3_1 _2272_ (.A(_1407_),
    .B(_1408_),
    .C(_1409_),
    .X(_1410_));
 sg13g2_nand3_1 _2273_ (.B(_1045_),
    .C(_1406_),
    .A(net460),
    .Y(_1411_));
 sg13g2_and2_1 _2274_ (.A(_0901_),
    .B(_1411_),
    .X(_1412_));
 sg13g2_nor2_1 _2275_ (.A(net465),
    .B(_1408_),
    .Y(_1413_));
 sg13g2_nor3_1 _2276_ (.A(_0959_),
    .B(_1033_),
    .C(_1405_),
    .Y(_1414_));
 sg13g2_nand2b_1 _2277_ (.Y(_1415_),
    .B(net465),
    .A_N(_1414_));
 sg13g2_nor2_1 _2278_ (.A(_1409_),
    .B(_1415_),
    .Y(_1416_));
 sg13g2_or2_1 _2279_ (.X(_1417_),
    .B(_1416_),
    .A(_1413_));
 sg13g2_and2_1 _2280_ (.A(_1039_),
    .B(_1406_),
    .X(_1418_));
 sg13g2_nor2_1 _2281_ (.A(_0897_),
    .B(_1418_),
    .Y(_1419_));
 sg13g2_nand2_1 _2282_ (.Y(_1420_),
    .A(net452),
    .B(_0965_));
 sg13g2_a21oi_1 _2283_ (.A1(_0932_),
    .A2(_0946_),
    .Y(_1421_),
    .B1(_1039_));
 sg13g2_nor3_1 _2284_ (.A(_1033_),
    .B(_1405_),
    .C(_1421_),
    .Y(_1422_));
 sg13g2_or2_1 _2285_ (.X(_1423_),
    .B(_1422_),
    .A(_1410_));
 sg13g2_nor2b_1 _2286_ (.A(_1415_),
    .B_N(_1423_),
    .Y(_1424_));
 sg13g2_o21ai_1 _2287_ (.B1(net451),
    .Y(_1425_),
    .A1(_1413_),
    .A2(_1424_));
 sg13g2_nor2_1 _2288_ (.A(_0917_),
    .B(_1054_),
    .Y(_1426_));
 sg13g2_nor3_1 _2289_ (.A(_0917_),
    .B(_0973_),
    .C(_1054_),
    .Y(_1427_));
 sg13g2_nor3_1 _2290_ (.A(_0970_),
    .B(_1414_),
    .C(_1422_),
    .Y(_1428_));
 sg13g2_o21ai_1 _2291_ (.B1(_1423_),
    .Y(_1429_),
    .A1(_1427_),
    .A2(_1428_));
 sg13g2_a21oi_1 _2292_ (.A1(_1425_),
    .A2(_1429_),
    .Y(_1430_),
    .B1(_0965_));
 sg13g2_xnor2_1 _2293_ (.Y(_1431_),
    .A(_0897_),
    .B(_0965_));
 sg13g2_a221oi_1 _2294_ (.B2(_1419_),
    .C1(_1431_),
    .B1(_1417_),
    .A1(_1410_),
    .Y(_1432_),
    .A2(_1412_));
 sg13g2_nor2b_1 _2295_ (.A(_1430_),
    .B_N(_1432_),
    .Y(_1433_));
 sg13g2_nand3_1 _2296_ (.B(net452),
    .C(_0965_),
    .A(_0894_),
    .Y(_1434_));
 sg13g2_xnor2_1 _2297_ (.Y(_1435_),
    .A(_0894_),
    .B(_1420_));
 sg13g2_o21ai_1 _2298_ (.B1(net465),
    .Y(_1436_),
    .A1(_1409_),
    .A2(_1418_));
 sg13g2_nand3_1 _2299_ (.B(_1411_),
    .C(_1436_),
    .A(_0900_),
    .Y(_1437_));
 sg13g2_nand2_1 _2300_ (.Y(_1438_),
    .A(net463),
    .B(_1407_));
 sg13g2_a21oi_1 _2301_ (.A1(_0909_),
    .A2(_1035_),
    .Y(_1439_),
    .B1(_1438_));
 sg13g2_nand4_1 _2302_ (.B(_1035_),
    .C(_1406_),
    .A(_0909_),
    .Y(_1440_),
    .D(_1438_));
 sg13g2_nand3b_1 _2303_ (.B(_1440_),
    .C(_0899_),
    .Y(_1441_),
    .A_N(_1439_));
 sg13g2_a21oi_1 _2304_ (.A1(_1437_),
    .A2(_1441_),
    .Y(_1442_),
    .B1(_0968_));
 sg13g2_nand2_1 _2305_ (.Y(_1443_),
    .A(_1436_),
    .B(_1438_));
 sg13g2_o21ai_1 _2306_ (.B1(_1431_),
    .Y(_1444_),
    .A1(net452),
    .A2(_1443_));
 sg13g2_nor3_1 _2307_ (.A(_1412_),
    .B(_1442_),
    .C(_1444_),
    .Y(_1445_));
 sg13g2_nor3_1 _2308_ (.A(_1433_),
    .B(_1435_),
    .C(_1445_),
    .Y(_1446_));
 sg13g2_a21oi_1 _2309_ (.A1(_1406_),
    .A2(_1426_),
    .Y(_1447_),
    .B1(_1423_));
 sg13g2_nand4_1 _2310_ (.B(_1026_),
    .C(_1035_),
    .A(_0909_),
    .Y(_1448_),
    .D(_1406_));
 sg13g2_a21oi_1 _2311_ (.A1(_1043_),
    .A2(_1044_),
    .Y(_1449_),
    .B1(_0973_));
 sg13g2_nand2_1 _2312_ (.Y(_1450_),
    .A(_1406_),
    .B(_1449_));
 sg13g2_nand3_1 _2313_ (.B(_1448_),
    .C(_1450_),
    .A(_1435_),
    .Y(_1451_));
 sg13g2_o21ai_1 _2314_ (.B1(_0894_),
    .Y(_1452_),
    .A1(net452),
    .A2(net451));
 sg13g2_nor2b_1 _2315_ (.A(_1452_),
    .B_N(_1420_),
    .Y(_1453_));
 sg13g2_xor2_1 _2316_ (.B(_1434_),
    .A(_0906_),
    .X(_1454_));
 sg13g2_nor4_1 _2317_ (.A(_1446_),
    .B(_1447_),
    .C(_1453_),
    .D(_1454_),
    .Y(_1455_));
 sg13g2_nand2_1 _2318_ (.Y(_1456_),
    .A(_1451_),
    .B(_1455_));
 sg13g2_nand4_1 _2319_ (.B(_1142_),
    .C(_1404_),
    .A(_1025_),
    .Y(_1457_),
    .D(_1456_));
 sg13g2_nor2_1 _2320_ (.A(\graphics_engine_1.anim_2x[0] ),
    .B(\graphics_engine_1.overlay_creator1.text_demosiine1.y[0] ),
    .Y(_1458_));
 sg13g2_and2_1 _2321_ (.A(net479),
    .B(\graphics_engine_1.ctr[7] ),
    .X(_1459_));
 sg13g2_xnor2_1 _2322_ (.Y(_1460_),
    .A(net479),
    .B(\graphics_engine_1.ctr[7] ));
 sg13g2_nand2_1 _2323_ (.Y(_1461_),
    .A(net481),
    .B(\graphics_engine_1.ctr[6] ));
 sg13g2_xnor2_1 _2324_ (.Y(_1462_),
    .A(net480),
    .B(\graphics_engine_1.ctr[6] ));
 sg13g2_inv_1 _2325_ (.Y(_1463_),
    .A(_1462_));
 sg13g2_nor2_2 _2326_ (.A(net493),
    .B(\graphics_engine_1.ctr[3] ),
    .Y(_1464_));
 sg13g2_nand2_1 _2327_ (.Y(_1465_),
    .A(net493),
    .B(\graphics_engine_1.ctr[3] ));
 sg13g2_and2_1 _2328_ (.A(net496),
    .B(\graphics_engine_1.ctr[2] ),
    .X(_1466_));
 sg13g2_nor2_1 _2329_ (.A(net496),
    .B(\graphics_engine_1.ctr[2] ),
    .Y(_1467_));
 sg13g2_nor2_1 _2330_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[1] ),
    .B(\graphics_engine_1.ctr[1] ),
    .Y(_1468_));
 sg13g2_a22oi_1 _2331_ (.Y(_1469_),
    .B1(\graphics_engine_1.ctr[0] ),
    .B2(\graphics_engine_1.anim_2x[0] ),
    .A2(\graphics_engine_1.ctr[1] ),
    .A1(\graphics_engine_1.overlay_creator1.text_demosiine1.x[1] ));
 sg13g2_or2_1 _2332_ (.X(_1470_),
    .B(_1469_),
    .A(_1468_));
 sg13g2_nor4_2 _2333_ (.A(_1466_),
    .B(_1467_),
    .C(_1468_),
    .Y(_1471_),
    .D(_1469_));
 sg13g2_nor2_1 _2334_ (.A(_1466_),
    .B(_1471_),
    .Y(_1472_));
 sg13g2_a221oi_1 _2335_ (.B2(net496),
    .C1(_1471_),
    .B1(\graphics_engine_1.ctr[2] ),
    .A1(net494),
    .Y(_1473_),
    .A2(\graphics_engine_1.ctr[3] ));
 sg13g2_nor2_1 _2336_ (.A(_1464_),
    .B(_1473_),
    .Y(_1474_));
 sg13g2_xnor2_1 _2337_ (.Y(_1475_),
    .A(net482),
    .B(\graphics_engine_1.ctr[5] ));
 sg13g2_nand2_1 _2338_ (.Y(_1476_),
    .A(net486),
    .B(\graphics_engine_1.ctr[4] ));
 sg13g2_xnor2_1 _2339_ (.Y(_1477_),
    .A(net486),
    .B(\graphics_engine_1.ctr[4] ));
 sg13g2_nor4_1 _2340_ (.A(_1464_),
    .B(_1473_),
    .C(_1475_),
    .D(_1477_),
    .Y(_1478_));
 sg13g2_nor2_1 _2341_ (.A(_1475_),
    .B(_1476_),
    .Y(_1479_));
 sg13g2_a21oi_1 _2342_ (.A1(net482),
    .A2(\graphics_engine_1.ctr[5] ),
    .Y(_1480_),
    .B1(_1479_));
 sg13g2_inv_1 _2343_ (.Y(_1481_),
    .A(_1480_));
 sg13g2_nor2_1 _2344_ (.A(_1478_),
    .B(_1481_),
    .Y(_1482_));
 sg13g2_o21ai_1 _2345_ (.B1(_1463_),
    .Y(_1483_),
    .A1(_1478_),
    .A2(_1481_));
 sg13g2_nand2_1 _2346_ (.Y(_1484_),
    .A(_1461_),
    .B(_1483_));
 sg13g2_a21oi_1 _2347_ (.A1(_1461_),
    .A2(_1483_),
    .Y(_1485_),
    .B1(_1460_));
 sg13g2_xor2_1 _2348_ (.B(\graphics_engine_1.ctr[8] ),
    .A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[8] ),
    .X(_1486_));
 sg13g2_o21ai_1 _2349_ (.B1(_1486_),
    .Y(_1487_),
    .A1(_1459_),
    .A2(_1485_));
 sg13g2_or3_2 _2350_ (.A(_1459_),
    .B(_1485_),
    .C(_1486_),
    .X(_1488_));
 sg13g2_nand3_1 _2351_ (.B(_1487_),
    .C(_1488_),
    .A(_1272_),
    .Y(_1489_));
 sg13g2_xor2_1 _2352_ (.B(_1489_),
    .A(_1158_),
    .X(_1490_));
 sg13g2_xnor2_1 _2353_ (.Y(_1491_),
    .A(_1158_),
    .B(_1489_));
 sg13g2_nand3_1 _2354_ (.B(_1487_),
    .C(_1488_),
    .A(_1152_),
    .Y(_1492_));
 sg13g2_xnor2_1 _2355_ (.Y(_1493_),
    .A(_1160_),
    .B(_1492_));
 sg13g2_xor2_1 _2356_ (.B(_1492_),
    .A(_1160_),
    .X(_1494_));
 sg13g2_nand3_1 _2357_ (.B(_1487_),
    .C(_1488_),
    .A(net504),
    .Y(_1495_));
 sg13g2_a21o_1 _2358_ (.A2(_1488_),
    .A1(_1487_),
    .B1(net504),
    .X(_1496_));
 sg13g2_nand3_1 _2359_ (.B(_1495_),
    .C(_1496_),
    .A(_1151_),
    .Y(_1497_));
 sg13g2_nand3_1 _2360_ (.B(net397),
    .C(_1497_),
    .A(_1490_),
    .Y(_1498_));
 sg13g2_nor2_1 _2361_ (.A(_1158_),
    .B(_1272_),
    .Y(_1499_));
 sg13g2_nand3_1 _2362_ (.B(_1488_),
    .C(_1499_),
    .A(_1487_),
    .Y(_1500_));
 sg13g2_xnor2_1 _2363_ (.Y(_1501_),
    .A(_0857_),
    .B(_1153_));
 sg13g2_xnor2_1 _2364_ (.Y(_1502_),
    .A(_1500_),
    .B(_1501_));
 sg13g2_xor2_1 _2365_ (.B(_1501_),
    .A(_1500_),
    .X(_1503_));
 sg13g2_a21oi_2 _2366_ (.B1(_1458_),
    .Y(_1504_),
    .A2(net396),
    .A1(_1498_));
 sg13g2_xnor2_1 _2367_ (.Y(_1505_),
    .A(_1460_),
    .B(_1484_));
 sg13g2_xor2_1 _2368_ (.B(_1484_),
    .A(_1460_),
    .X(_1506_));
 sg13g2_xnor2_1 _2369_ (.Y(_1507_),
    .A(_1463_),
    .B(_1482_));
 sg13g2_xnor2_1 _2370_ (.Y(_1508_),
    .A(_1462_),
    .B(_1482_));
 sg13g2_or3_1 _2371_ (.A(_1464_),
    .B(_1473_),
    .C(_1477_),
    .X(_1509_));
 sg13g2_nand3_1 _2372_ (.B(_1476_),
    .C(_1509_),
    .A(_1475_),
    .Y(_1510_));
 sg13g2_a21o_1 _2373_ (.A2(_1509_),
    .A1(_1476_),
    .B1(_1475_),
    .X(_1511_));
 sg13g2_and2_2 _2374_ (.A(_1510_),
    .B(_1511_),
    .X(_1512_));
 sg13g2_nand2_1 _2375_ (.Y(_1513_),
    .A(_1510_),
    .B(_1511_));
 sg13g2_nor2_2 _2376_ (.A(net433),
    .B(net427),
    .Y(_1514_));
 sg13g2_inv_1 _2377_ (.Y(_1515_),
    .A(_1514_));
 sg13g2_xnor2_1 _2378_ (.Y(_1516_),
    .A(_1474_),
    .B(_1477_));
 sg13g2_xor2_1 _2379_ (.B(_1477_),
    .A(_1474_),
    .X(_1517_));
 sg13g2_nor2b_1 _2380_ (.A(_1464_),
    .B_N(_1465_),
    .Y(_1518_));
 sg13g2_xor2_1 _2381_ (.B(_1518_),
    .A(_1472_),
    .X(_1519_));
 sg13g2_xnor2_1 _2382_ (.Y(_1520_),
    .A(_1472_),
    .B(_1518_));
 sg13g2_nor2_2 _2383_ (.A(_1517_),
    .B(_1519_),
    .Y(_1521_));
 sg13g2_nand2_2 _2384_ (.Y(_1522_),
    .A(net443),
    .B(_1520_));
 sg13g2_nand3_1 _2385_ (.B(_1512_),
    .C(_1522_),
    .A(net429),
    .Y(_1523_));
 sg13g2_nor4_2 _2386_ (.A(net400),
    .B(net398),
    .C(_1497_),
    .Y(_1524_),
    .D(net394));
 sg13g2_nand2b_1 _2387_ (.Y(_1525_),
    .B(_1524_),
    .A_N(_1523_));
 sg13g2_a21o_2 _2388_ (.A2(_1496_),
    .A1(_1495_),
    .B1(_1151_),
    .X(_1526_));
 sg13g2_nor2_2 _2389_ (.A(net396),
    .B(_1526_),
    .Y(_1527_));
 sg13g2_nor4_2 _2390_ (.A(net400),
    .B(net397),
    .C(net394),
    .Y(_1528_),
    .D(_1526_));
 sg13g2_a22oi_1 _2391_ (.Y(_1529_),
    .B1(net443),
    .B2(_1520_),
    .A2(_1511_),
    .A1(_1510_));
 sg13g2_nand3_1 _2392_ (.B(_1511_),
    .C(net443),
    .A(_1510_),
    .Y(_1530_));
 sg13g2_nand2_2 _2393_ (.Y(_1531_),
    .A(net431),
    .B(net428));
 sg13g2_and2_1 _2394_ (.A(net429),
    .B(_1530_),
    .X(_1532_));
 sg13g2_nand2_1 _2395_ (.Y(_1533_),
    .A(net430),
    .B(_1530_));
 sg13g2_nand3b_1 _2396_ (.B(_1532_),
    .C(_1528_),
    .Y(_1534_),
    .A_N(_1529_));
 sg13g2_a21oi_1 _2397_ (.A1(_1525_),
    .A2(_1534_),
    .Y(_1535_),
    .B1(net412));
 sg13g2_a21o_2 _2398_ (.A2(_1496_),
    .A1(_1495_),
    .B1(_1152_),
    .X(_1536_));
 sg13g2_nor4_2 _2399_ (.A(_1491_),
    .B(net397),
    .C(net395),
    .Y(_1537_),
    .D(_1536_));
 sg13g2_nor2_1 _2400_ (.A(net429),
    .B(_1512_),
    .Y(_1538_));
 sg13g2_nand2_1 _2401_ (.Y(_1539_),
    .A(net433),
    .B(net427));
 sg13g2_nor2_1 _2402_ (.A(net443),
    .B(_1520_),
    .Y(_1540_));
 sg13g2_nand2_1 _2403_ (.Y(_1541_),
    .A(_1517_),
    .B(_1519_));
 sg13g2_nor2_1 _2404_ (.A(net429),
    .B(net426),
    .Y(_1542_));
 sg13g2_nand3_1 _2405_ (.B(net427),
    .C(_1541_),
    .A(net434),
    .Y(_1543_));
 sg13g2_nand2_2 _2406_ (.Y(_1544_),
    .A(_1514_),
    .B(_1540_));
 sg13g2_a22oi_1 _2407_ (.Y(_1545_),
    .B1(_1543_),
    .B2(_1544_),
    .A2(_1522_),
    .A1(net411));
 sg13g2_nand3_1 _2408_ (.B(_1495_),
    .C(_1496_),
    .A(_1152_),
    .Y(_1546_));
 sg13g2_nor4_2 _2409_ (.A(net400),
    .B(net397),
    .C(net394),
    .Y(_1547_),
    .D(_1546_));
 sg13g2_nor2_2 _2410_ (.A(_1512_),
    .B(net443),
    .Y(_1548_));
 sg13g2_nor2_2 _2411_ (.A(net427),
    .B(net426),
    .Y(_1549_));
 sg13g2_o21ai_1 _2412_ (.B1(net431),
    .Y(_1550_),
    .A1(net428),
    .A2(net426));
 sg13g2_or2_1 _2413_ (.X(_1551_),
    .B(_1550_),
    .A(_1548_));
 sg13g2_nor2_1 _2414_ (.A(net412),
    .B(_1551_),
    .Y(_1552_));
 sg13g2_a22oi_1 _2415_ (.Y(_1553_),
    .B1(_1547_),
    .B2(_1552_),
    .A2(_1545_),
    .A1(_1537_));
 sg13g2_nor4_2 _2416_ (.A(net399),
    .B(net398),
    .C(net395),
    .Y(_1554_),
    .D(_1536_));
 sg13g2_nand2b_1 _2417_ (.Y(_1555_),
    .B(net432),
    .A_N(_1529_));
 sg13g2_nor2_2 _2418_ (.A(net431),
    .B(net427),
    .Y(_1556_));
 sg13g2_nand2_1 _2419_ (.Y(_1557_),
    .A(net432),
    .B(_1512_));
 sg13g2_nor2_1 _2420_ (.A(_1522_),
    .B(_1539_),
    .Y(_1558_));
 sg13g2_nand2_1 _2421_ (.Y(_1559_),
    .A(_1521_),
    .B(_1538_));
 sg13g2_nand3b_1 _2422_ (.B(_1530_),
    .C(net432),
    .Y(_1560_),
    .A_N(_1529_));
 sg13g2_nand2_2 _2423_ (.Y(_1561_),
    .A(net431),
    .B(_1549_));
 sg13g2_nor2_1 _2424_ (.A(_1523_),
    .B(net426),
    .Y(_1562_));
 sg13g2_nor2_1 _2425_ (.A(net406),
    .B(_1562_),
    .Y(_1563_));
 sg13g2_nor2_1 _2426_ (.A(net430),
    .B(_1530_),
    .Y(_1564_));
 sg13g2_nand2_1 _2427_ (.Y(_1565_),
    .A(net444),
    .B(_1556_));
 sg13g2_nand2_2 _2428_ (.Y(_1566_),
    .A(_1521_),
    .B(_1556_));
 sg13g2_nand2_1 _2429_ (.Y(_1567_),
    .A(net432),
    .B(_1529_));
 sg13g2_a21oi_2 _2430_ (.B1(net410),
    .Y(_1568_),
    .A2(_1542_),
    .A1(_1529_));
 sg13g2_o21ai_1 _2431_ (.B1(net407),
    .Y(_1569_),
    .A1(_1521_),
    .A2(_1543_));
 sg13g2_a22oi_1 _2432_ (.Y(_1570_),
    .B1(_1566_),
    .B2(_1568_),
    .A2(_1563_),
    .A1(_1560_));
 sg13g2_nor4_2 _2433_ (.A(net399),
    .B(net397),
    .C(_1497_),
    .Y(_1571_),
    .D(net396));
 sg13g2_a21oi_2 _2434_ (.B1(net407),
    .Y(_1572_),
    .A2(_1556_),
    .A1(net426));
 sg13g2_nand3_1 _2435_ (.B(net428),
    .C(_1521_),
    .A(net431),
    .Y(_1573_));
 sg13g2_and2_1 _2436_ (.A(net408),
    .B(_1573_),
    .X(_1574_));
 sg13g2_a21oi_1 _2437_ (.A1(_1567_),
    .A2(_1574_),
    .Y(_1575_),
    .B1(_1572_));
 sg13g2_nand2_1 _2438_ (.Y(_1576_),
    .A(_1571_),
    .B(_1575_));
 sg13g2_nor4_2 _2439_ (.A(net400),
    .B(net397),
    .C(net394),
    .Y(_1577_),
    .D(_1536_));
 sg13g2_nor2_1 _2440_ (.A(net414),
    .B(_1531_),
    .Y(_1578_));
 sg13g2_nor3_1 _2441_ (.A(net414),
    .B(_1531_),
    .C(net426),
    .Y(_1579_));
 sg13g2_nor4_2 _2442_ (.A(net399),
    .B(net398),
    .C(_1497_),
    .Y(_1580_),
    .D(net394));
 sg13g2_nor2_2 _2443_ (.A(_1512_),
    .B(_1541_),
    .Y(_1581_));
 sg13g2_nand2_1 _2444_ (.Y(_1582_),
    .A(net433),
    .B(net405));
 sg13g2_nand3_1 _2445_ (.B(net427),
    .C(net426),
    .A(net434),
    .Y(_1583_));
 sg13g2_nand2_2 _2446_ (.Y(_1584_),
    .A(_1512_),
    .B(_1521_));
 sg13g2_o21ai_1 _2447_ (.B1(_1539_),
    .Y(_1585_),
    .A1(net434),
    .A2(_1584_));
 sg13g2_o21ai_1 _2448_ (.B1(_1583_),
    .Y(_1586_),
    .A1(net434),
    .A2(_1584_));
 sg13g2_nand2_2 _2449_ (.Y(_1587_),
    .A(net433),
    .B(_1549_));
 sg13g2_nand2b_1 _2450_ (.Y(_1588_),
    .B(_1587_),
    .A_N(_1586_));
 sg13g2_nor4_2 _2451_ (.A(net399),
    .B(_1494_),
    .C(net395),
    .Y(_1589_),
    .D(_1526_));
 sg13g2_or4_2 _2452_ (.A(net399),
    .B(_1494_),
    .C(net396),
    .D(_1526_),
    .X(_1590_));
 sg13g2_nor2_2 _2453_ (.A(net443),
    .B(_1519_),
    .Y(_1591_));
 sg13g2_nand2_2 _2454_ (.Y(_1592_),
    .A(_1517_),
    .B(_1520_));
 sg13g2_nand2_1 _2455_ (.Y(_1593_),
    .A(net432),
    .B(_1591_));
 sg13g2_nor2_2 _2456_ (.A(_1512_),
    .B(_1592_),
    .Y(_1594_));
 sg13g2_nor2_1 _2457_ (.A(_1512_),
    .B(_1593_),
    .Y(_1595_));
 sg13g2_nand2_1 _2458_ (.Y(_1596_),
    .A(net434),
    .B(_1594_));
 sg13g2_nor2_1 _2459_ (.A(net406),
    .B(_1564_),
    .Y(_1597_));
 sg13g2_nand2_1 _2460_ (.Y(_1598_),
    .A(net412),
    .B(_1565_));
 sg13g2_nor2_2 _2461_ (.A(_1517_),
    .B(_1520_),
    .Y(_1599_));
 sg13g2_nand2b_2 _2462_ (.Y(_1600_),
    .B(net429),
    .A_N(_1530_));
 sg13g2_a21oi_1 _2463_ (.A1(_1514_),
    .A2(_1599_),
    .Y(_1601_),
    .B1(net411));
 sg13g2_o21ai_1 _2464_ (.B1(net406),
    .Y(_1602_),
    .A1(_1520_),
    .A2(_1600_));
 sg13g2_a22oi_1 _2465_ (.Y(_1603_),
    .B1(_1601_),
    .B2(_1560_),
    .A2(_1597_),
    .A1(_1596_));
 sg13g2_nor4_2 _2466_ (.A(_1491_),
    .B(net397),
    .C(net395),
    .Y(_1604_),
    .D(_1546_));
 sg13g2_nand2_2 _2467_ (.Y(_1605_),
    .A(_1538_),
    .B(_1599_));
 sg13g2_nand3_1 _2468_ (.B(_1566_),
    .C(_1605_),
    .A(net409),
    .Y(_1606_));
 sg13g2_nand3b_1 _2469_ (.B(net432),
    .C(_1530_),
    .Y(_1607_),
    .A_N(net405));
 sg13g2_nor2_1 _2470_ (.A(net409),
    .B(_1514_),
    .Y(_1608_));
 sg13g2_nor3_1 _2471_ (.A(net432),
    .B(net427),
    .C(_1592_),
    .Y(_1609_));
 sg13g2_inv_1 _2472_ (.Y(_1610_),
    .A(_1609_));
 sg13g2_nor2_1 _2473_ (.A(net409),
    .B(_1609_),
    .Y(_1611_));
 sg13g2_o21ai_1 _2474_ (.B1(_1611_),
    .Y(_1612_),
    .A1(_1591_),
    .A2(_1607_));
 sg13g2_and2_1 _2475_ (.A(_1606_),
    .B(_1612_),
    .X(_1613_));
 sg13g2_nand3_1 _2476_ (.B(net427),
    .C(_1599_),
    .A(net430),
    .Y(_1614_));
 sg13g2_inv_1 _2477_ (.Y(_1615_),
    .A(_1614_));
 sg13g2_nor2_1 _2478_ (.A(net414),
    .B(_1615_),
    .Y(_1616_));
 sg13g2_nor2_1 _2479_ (.A(_1586_),
    .B(_1595_),
    .Y(_1617_));
 sg13g2_nor4_2 _2480_ (.A(net400),
    .B(net398),
    .C(net394),
    .Y(_1618_),
    .D(_1526_));
 sg13g2_nor2_1 _2481_ (.A(_1557_),
    .B(_1592_),
    .Y(_1619_));
 sg13g2_nor2_1 _2482_ (.A(net406),
    .B(_1619_),
    .Y(_1620_));
 sg13g2_a21oi_1 _2483_ (.A1(_1616_),
    .A2(_1617_),
    .Y(_1621_),
    .B1(_1620_));
 sg13g2_nor2_1 _2484_ (.A(net414),
    .B(_1564_),
    .Y(_1622_));
 sg13g2_nor3_2 _2485_ (.A(net399),
    .B(net398),
    .C(_1622_),
    .Y(_1623_));
 sg13g2_nand2_1 _2486_ (.Y(_1624_),
    .A(net430),
    .B(_1548_));
 sg13g2_nand4_1 _2487_ (.B(_1583_),
    .C(_1600_),
    .A(net412),
    .Y(_1625_),
    .D(_1624_));
 sg13g2_nand3_1 _2488_ (.B(_1623_),
    .C(_1625_),
    .A(_1527_),
    .Y(_1626_));
 sg13g2_nor2_2 _2489_ (.A(net413),
    .B(_1624_),
    .Y(_1627_));
 sg13g2_nor4_2 _2490_ (.A(net399),
    .B(net398),
    .C(_1502_),
    .Y(_1628_),
    .D(_1526_));
 sg13g2_nor4_2 _2491_ (.A(net400),
    .B(_1493_),
    .C(net396),
    .Y(_1629_),
    .D(_1546_));
 sg13g2_nor2_1 _2492_ (.A(net407),
    .B(_1556_),
    .Y(_1630_));
 sg13g2_a21o_1 _2493_ (.A2(_1599_),
    .A1(_1556_),
    .B1(net408),
    .X(_1631_));
 sg13g2_nand2_1 _2494_ (.Y(_1632_),
    .A(net408),
    .B(_1531_));
 sg13g2_a21oi_2 _2495_ (.B1(net412),
    .Y(_1633_),
    .A2(_1594_),
    .A1(net430));
 sg13g2_nand3_1 _2496_ (.B(_1600_),
    .C(_1633_),
    .A(_1583_),
    .Y(_1634_));
 sg13g2_nand3_1 _2497_ (.B(_1631_),
    .C(_1634_),
    .A(_1629_),
    .Y(_1635_));
 sg13g2_nor3_2 _2498_ (.A(net413),
    .B(_1521_),
    .C(_1531_),
    .Y(_1636_));
 sg13g2_nor4_2 _2499_ (.A(net400),
    .B(net397),
    .C(_1497_),
    .Y(_1637_),
    .D(net394));
 sg13g2_nor4_2 _2500_ (.A(net400),
    .B(net398),
    .C(net394),
    .Y(_1638_),
    .D(_1536_));
 sg13g2_nand2_1 _2501_ (.Y(_1639_),
    .A(net430),
    .B(_1581_));
 sg13g2_nand2_1 _2502_ (.Y(_1640_),
    .A(_1561_),
    .B(_1639_));
 sg13g2_nor2_1 _2503_ (.A(net406),
    .B(_1584_),
    .Y(_1641_));
 sg13g2_mux2_1 _2504_ (.A0(_1641_),
    .A1(_1506_),
    .S(_1640_),
    .X(_1642_));
 sg13g2_o21ai_1 _2505_ (.B1(net411),
    .Y(_1643_),
    .A1(net405),
    .A2(_1550_));
 sg13g2_nand2b_1 _2506_ (.Y(_1644_),
    .B(_1543_),
    .A_N(_1643_));
 sg13g2_nor4_2 _2507_ (.A(_1491_),
    .B(_1493_),
    .C(net396),
    .Y(_1645_),
    .D(_1546_));
 sg13g2_nand2_2 _2508_ (.Y(_1646_),
    .A(net406),
    .B(_1560_));
 sg13g2_inv_1 _2509_ (.Y(_1647_),
    .A(_1646_));
 sg13g2_nand3_1 _2510_ (.B(_1645_),
    .C(_1646_),
    .A(_1644_),
    .Y(_1648_));
 sg13g2_nor2_2 _2511_ (.A(net414),
    .B(_1639_),
    .Y(_1649_));
 sg13g2_nor4_2 _2512_ (.A(net399),
    .B(net398),
    .C(_1502_),
    .Y(_1650_),
    .D(_1546_));
 sg13g2_nand4_1 _2513_ (.B(_1626_),
    .C(_1635_),
    .A(_1553_),
    .Y(_1651_),
    .D(_1648_));
 sg13g2_a22oi_1 _2514_ (.Y(_0108_),
    .B1(_1589_),
    .B2(_1603_),
    .A2(_1579_),
    .A1(_1577_));
 sg13g2_a22oi_1 _2515_ (.Y(_0109_),
    .B1(_1627_),
    .B2(_1628_),
    .A2(_1621_),
    .A1(_1618_));
 sg13g2_a22oi_1 _2516_ (.Y(_0110_),
    .B1(_1636_),
    .B2(_1637_),
    .A2(_1570_),
    .A1(_1554_));
 sg13g2_a22oi_1 _2517_ (.Y(_0111_),
    .B1(_1649_),
    .B2(_1650_),
    .A2(_1642_),
    .A1(_1638_));
 sg13g2_nand4_1 _2518_ (.B(_0109_),
    .C(_0110_),
    .A(_0108_),
    .Y(_0112_),
    .D(_0111_));
 sg13g2_a22oi_1 _2519_ (.Y(_0113_),
    .B1(_1604_),
    .B2(_1613_),
    .A2(_1588_),
    .A1(_1580_));
 sg13g2_nand2_1 _2520_ (.Y(_0114_),
    .A(_1576_),
    .B(_0113_));
 sg13g2_or4_1 _2521_ (.A(_1535_),
    .B(_1651_),
    .C(_0112_),
    .D(_0114_),
    .X(_0115_));
 sg13g2_and2_1 _2522_ (.A(_1504_),
    .B(_0115_),
    .X(_0116_));
 sg13g2_nand2_2 _2523_ (.Y(_0117_),
    .A(_1504_),
    .B(_0115_));
 sg13g2_nand3_1 _2524_ (.B(_1528_),
    .C(_1578_),
    .A(_1517_),
    .Y(_0118_));
 sg13g2_nand3_1 _2525_ (.B(_1560_),
    .C(_1605_),
    .A(net409),
    .Y(_0119_));
 sg13g2_nor2_1 _2526_ (.A(net409),
    .B(_1586_),
    .Y(_0120_));
 sg13g2_nand3_1 _2527_ (.B(_1561_),
    .C(_1583_),
    .A(net408),
    .Y(_0121_));
 sg13g2_nand3_1 _2528_ (.B(_0119_),
    .C(_0121_),
    .A(_1604_),
    .Y(_0122_));
 sg13g2_or2_1 _2529_ (.X(_0123_),
    .B(_1581_),
    .A(_1550_));
 sg13g2_nand2_1 _2530_ (.Y(_0124_),
    .A(net408),
    .B(_0123_));
 sg13g2_nand3_1 _2531_ (.B(_1629_),
    .C(_0124_),
    .A(_1598_),
    .Y(_0125_));
 sg13g2_nor2_1 _2532_ (.A(_1556_),
    .B(_1646_),
    .Y(_0126_));
 sg13g2_o21ai_1 _2533_ (.B1(net411),
    .Y(_0127_),
    .A1(net433),
    .A2(net405));
 sg13g2_nor2b_1 _2534_ (.A(_0126_),
    .B_N(_0127_),
    .Y(_0128_));
 sg13g2_a21oi_1 _2535_ (.A1(net410),
    .A2(_1555_),
    .Y(_0129_),
    .B1(_1641_));
 sg13g2_nor2b_1 _2536_ (.A(_1608_),
    .B_N(_0129_),
    .Y(_0130_));
 sg13g2_a22oi_1 _2537_ (.Y(_0131_),
    .B1(_0130_),
    .B2(_1537_),
    .A2(_0128_),
    .A1(_1645_));
 sg13g2_and2_1 _2538_ (.A(_1582_),
    .B(_1600_),
    .X(_0132_));
 sg13g2_a22oi_1 _2539_ (.Y(_0133_),
    .B1(_0132_),
    .B2(_1563_),
    .A2(_1607_),
    .A1(_1568_));
 sg13g2_a221oi_1 _2540_ (.B2(_1617_),
    .C1(_1590_),
    .B1(_1601_),
    .A1(_1543_),
    .Y(_0134_),
    .A2(_1572_));
 sg13g2_nand2_2 _2541_ (.Y(_0135_),
    .A(net412),
    .B(_1566_));
 sg13g2_nand3_1 _2542_ (.B(_1638_),
    .C(_0135_),
    .A(_1632_),
    .Y(_0136_));
 sg13g2_o21ai_1 _2543_ (.B1(_1616_),
    .Y(_0137_),
    .A1(_1529_),
    .A2(_1533_));
 sg13g2_nand2_1 _2544_ (.Y(_0138_),
    .A(net410),
    .B(_1587_));
 sg13g2_nand3_1 _2545_ (.B(_0137_),
    .C(_0138_),
    .A(_1618_),
    .Y(_0139_));
 sg13g2_nand2_1 _2546_ (.Y(_0140_),
    .A(net413),
    .B(_1550_));
 sg13g2_nand3_1 _2547_ (.B(_1623_),
    .C(_0140_),
    .A(_1527_),
    .Y(_0141_));
 sg13g2_and2_1 _2548_ (.A(_1523_),
    .B(_1574_),
    .X(_0142_));
 sg13g2_nor2_1 _2549_ (.A(_1630_),
    .B(_0142_),
    .Y(_0143_));
 sg13g2_a22oi_1 _2550_ (.Y(_0144_),
    .B1(_1649_),
    .B2(_1547_),
    .A2(_1585_),
    .A1(_1580_));
 sg13g2_and4_1 _2551_ (.A(_0131_),
    .B(_0139_),
    .C(_0141_),
    .D(_0144_),
    .X(_0145_));
 sg13g2_and4_1 _2552_ (.A(_0118_),
    .B(_0122_),
    .C(_0125_),
    .D(_0136_),
    .X(_0146_));
 sg13g2_a21oi_1 _2553_ (.A1(_1524_),
    .A2(_1636_),
    .Y(_0147_),
    .B1(_0134_));
 sg13g2_a22oi_1 _2554_ (.Y(_0148_),
    .B1(_0143_),
    .B2(_1571_),
    .A2(_0133_),
    .A1(_1554_));
 sg13g2_nand4_1 _2555_ (.B(_0146_),
    .C(_0147_),
    .A(_0145_),
    .Y(_0149_),
    .D(_0148_));
 sg13g2_o21ai_1 _2556_ (.B1(net408),
    .Y(_0150_),
    .A1(_1533_),
    .A2(_1594_));
 sg13g2_nand3_1 _2557_ (.B(_0135_),
    .C(_0150_),
    .A(_1638_),
    .Y(_0151_));
 sg13g2_nand3_1 _2558_ (.B(_1573_),
    .C(_1633_),
    .A(_1523_),
    .Y(_0152_));
 sg13g2_nand3_1 _2559_ (.B(_1631_),
    .C(_0152_),
    .A(_1629_),
    .Y(_0153_));
 sg13g2_nand4_1 _2560_ (.B(_1523_),
    .C(_1573_),
    .A(net413),
    .Y(_0154_),
    .D(_1624_));
 sg13g2_nand3_1 _2561_ (.B(_1623_),
    .C(_0154_),
    .A(_1527_),
    .Y(_0155_));
 sg13g2_nor2_1 _2562_ (.A(net413),
    .B(_0123_),
    .Y(_0156_));
 sg13g2_a22oi_1 _2563_ (.Y(_0157_),
    .B1(_1568_),
    .B2(_1557_),
    .A2(_1563_),
    .A1(_1539_));
 sg13g2_a22oi_1 _2564_ (.Y(_0158_),
    .B1(_0157_),
    .B2(_1554_),
    .A2(_0156_),
    .A1(_1524_));
 sg13g2_nand4_1 _2565_ (.B(_0153_),
    .C(_0155_),
    .A(_0151_),
    .Y(_0159_),
    .D(_0158_));
 sg13g2_nand2_1 _2566_ (.Y(_0160_),
    .A(_1565_),
    .B(_1572_));
 sg13g2_nand3_1 _2567_ (.B(_1574_),
    .C(_1583_),
    .A(_1561_),
    .Y(_0161_));
 sg13g2_nand3_1 _2568_ (.B(_0160_),
    .C(_0161_),
    .A(_1571_),
    .Y(_0162_));
 sg13g2_nand3_1 _2569_ (.B(_1559_),
    .C(_1587_),
    .A(net409),
    .Y(_0163_));
 sg13g2_nand3_1 _2570_ (.B(_1544_),
    .C(_0132_),
    .A(net406),
    .Y(_0164_));
 sg13g2_nand3_1 _2571_ (.B(_0163_),
    .C(_0164_),
    .A(_1537_),
    .Y(_0165_));
 sg13g2_o21ai_1 _2572_ (.B1(_0129_),
    .Y(_0166_),
    .A1(_1538_),
    .A2(_1602_));
 sg13g2_a21o_1 _2573_ (.A2(_0166_),
    .A1(_1596_),
    .B1(_1590_),
    .X(_0167_));
 sg13g2_nand3_1 _2574_ (.B(_0165_),
    .C(_0167_),
    .A(_0162_),
    .Y(_0168_));
 sg13g2_a22oi_1 _2575_ (.Y(_0169_),
    .B1(_1620_),
    .B2(_1566_),
    .A2(_1614_),
    .A1(_1608_));
 sg13g2_nand2b_1 _2576_ (.Y(_0170_),
    .B(_1607_),
    .A_N(_1586_));
 sg13g2_a22oi_1 _2577_ (.Y(_0171_),
    .B1(_0170_),
    .B2(_1580_),
    .A2(_0169_),
    .A1(_1618_));
 sg13g2_a22oi_1 _2578_ (.Y(_0172_),
    .B1(_1636_),
    .B2(_1547_),
    .A2(_1627_),
    .A1(_1577_));
 sg13g2_a22oi_1 _2579_ (.Y(_0173_),
    .B1(_1637_),
    .B2(_1649_),
    .A2(_1578_),
    .A1(_1528_));
 sg13g2_nor2_1 _2580_ (.A(_1569_),
    .B(_1586_),
    .Y(_0174_));
 sg13g2_a22oi_1 _2581_ (.Y(_0175_),
    .B1(_0174_),
    .B2(_1610_),
    .A2(_1630_),
    .A1(_1605_));
 sg13g2_nor3_1 _2582_ (.A(net432),
    .B(net405),
    .C(_1591_),
    .Y(_0176_));
 sg13g2_nor2_1 _2583_ (.A(_1643_),
    .B(_0176_),
    .Y(_0177_));
 sg13g2_a22oi_1 _2584_ (.Y(_0178_),
    .B1(_0177_),
    .B2(_1582_),
    .A2(_1647_),
    .A1(_1566_));
 sg13g2_a22oi_1 _2585_ (.Y(_0179_),
    .B1(_0178_),
    .B2(_1645_),
    .A2(_0175_),
    .A1(_1604_));
 sg13g2_nand4_1 _2586_ (.B(_0172_),
    .C(_0173_),
    .A(_0171_),
    .Y(_0180_),
    .D(_0179_));
 sg13g2_or3_1 _2587_ (.A(_0159_),
    .B(_0168_),
    .C(_0180_),
    .X(_0181_));
 sg13g2_o21ai_1 _2588_ (.B1(_1504_),
    .Y(_0182_),
    .A1(_0149_),
    .A2(_0181_));
 sg13g2_a21o_2 _2589_ (.A2(_0182_),
    .A1(_0117_),
    .B1(net2),
    .X(_0183_));
 sg13g2_nor3_1 _2590_ (.A(net2),
    .B(_0116_),
    .C(_0182_),
    .Y(_0184_));
 sg13g2_xnor2_1 _2591_ (.Y(_0185_),
    .A(net508),
    .B(net444));
 sg13g2_nand2_1 _2592_ (.Y(_0186_),
    .A(net513),
    .B(_1520_));
 sg13g2_o21ai_1 _2593_ (.B1(_1470_),
    .Y(_0187_),
    .A1(_1466_),
    .A2(_1467_));
 sg13g2_nor2b_1 _2594_ (.A(_1471_),
    .B_N(_0187_),
    .Y(_0188_));
 sg13g2_nand2_1 _2595_ (.Y(_0189_),
    .A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[1] ),
    .B(_0188_));
 sg13g2_nor2_1 _2596_ (.A(net513),
    .B(_1520_),
    .Y(_0190_));
 sg13g2_xnor2_1 _2597_ (.Y(_0191_),
    .A(net513),
    .B(_1519_));
 sg13g2_o21ai_1 _2598_ (.B1(_0186_),
    .Y(_0192_),
    .A1(_0189_),
    .A2(_0190_));
 sg13g2_nor2b_1 _2599_ (.A(_0185_),
    .B_N(_0192_),
    .Y(_0193_));
 sg13g2_xor2_1 _2600_ (.B(_0192_),
    .A(_0185_),
    .X(_0194_));
 sg13g2_nor2_1 _2601_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[1] ),
    .B(_0188_),
    .Y(_0195_));
 sg13g2_xnor2_1 _2602_ (.Y(_0196_),
    .A(_0191_),
    .B(_0195_));
 sg13g2_nand2_1 _2603_ (.Y(_0197_),
    .A(_0194_),
    .B(_0196_));
 sg13g2_xor2_1 _2604_ (.B(_0188_),
    .A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[1] ),
    .X(_0198_));
 sg13g2_xor2_1 _2605_ (.B(_0191_),
    .A(_0189_),
    .X(_0199_));
 sg13g2_nand2_1 _2606_ (.Y(_0200_),
    .A(_0194_),
    .B(_0199_));
 sg13g2_a21oi_1 _2607_ (.A1(net511),
    .A2(net444),
    .Y(_0201_),
    .B1(_0193_));
 sg13g2_xnor2_1 _2608_ (.Y(_0202_),
    .A(net507),
    .B(net428));
 sg13g2_xnor2_1 _2609_ (.Y(_0203_),
    .A(_0201_),
    .B(_0202_));
 sg13g2_xnor2_1 _2610_ (.Y(_0204_),
    .A(_0200_),
    .B(_0203_));
 sg13g2_inv_1 _2611_ (.Y(_0205_),
    .A(_0204_));
 sg13g2_nor2_1 _2612_ (.A(_0198_),
    .B(_0204_),
    .Y(_0206_));
 sg13g2_nor2_1 _2613_ (.A(_0197_),
    .B(_0206_),
    .Y(_0207_));
 sg13g2_a21oi_1 _2614_ (.A1(_0197_),
    .A2(_0205_),
    .Y(_0208_),
    .B1(_0207_));
 sg13g2_and2_1 _2615_ (.A(net481),
    .B(\graphics_engine_1.ctr[5] ),
    .X(_0209_));
 sg13g2_nand2_1 _2616_ (.Y(_0210_),
    .A(net481),
    .B(\graphics_engine_1.ctr[5] ));
 sg13g2_nand2_1 _2617_ (.Y(_0211_),
    .A(net483),
    .B(\graphics_engine_1.ctr[4] ));
 sg13g2_xnor2_1 _2618_ (.Y(_0212_),
    .A(net483),
    .B(\graphics_engine_1.ctr[4] ));
 sg13g2_nor2_1 _2619_ (.A(net487),
    .B(\graphics_engine_1.ctr[3] ),
    .Y(_0213_));
 sg13g2_and2_1 _2620_ (.A(net494),
    .B(\graphics_engine_1.ctr[2] ),
    .X(_0214_));
 sg13g2_nand2_1 _2621_ (.Y(_0215_),
    .A(net496),
    .B(\graphics_engine_1.ctr[1] ));
 sg13g2_xnor2_1 _2622_ (.Y(_0216_),
    .A(net495),
    .B(\graphics_engine_1.ctr[1] ));
 sg13g2_nand2_1 _2623_ (.Y(_0217_),
    .A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[1] ),
    .B(\graphics_engine_1.ctr[0] ));
 sg13g2_o21ai_1 _2624_ (.B1(_0215_),
    .Y(_0218_),
    .A1(_0216_),
    .A2(_0217_));
 sg13g2_xor2_1 _2625_ (.B(\graphics_engine_1.ctr[2] ),
    .A(net493),
    .X(_0219_));
 sg13g2_a21oi_2 _2626_ (.B1(_0214_),
    .Y(_0220_),
    .A2(_0219_),
    .A1(_0218_));
 sg13g2_a221oi_1 _2627_ (.B2(_0219_),
    .C1(_0214_),
    .B1(_0218_),
    .A1(net487),
    .Y(_0221_),
    .A2(\graphics_engine_1.ctr[3] ));
 sg13g2_or3_2 _2628_ (.A(_0212_),
    .B(_0213_),
    .C(_0221_),
    .X(_0222_));
 sg13g2_and2_1 _2629_ (.A(_0211_),
    .B(_0222_),
    .X(_0223_));
 sg13g2_xnor2_1 _2630_ (.Y(_0224_),
    .A(net481),
    .B(\graphics_engine_1.ctr[5] ));
 sg13g2_a21oi_1 _2631_ (.A1(_0211_),
    .A2(_0222_),
    .Y(_0225_),
    .B1(_0224_));
 sg13g2_a21o_1 _2632_ (.A2(_0222_),
    .A1(_0211_),
    .B1(_0224_),
    .X(_0226_));
 sg13g2_xnor2_1 _2633_ (.Y(_0227_),
    .A(net479),
    .B(\graphics_engine_1.ctr[6] ));
 sg13g2_xor2_1 _2634_ (.B(\graphics_engine_1.ctr[6] ),
    .A(net479),
    .X(_0228_));
 sg13g2_a21oi_2 _2635_ (.B1(_0228_),
    .Y(_0229_),
    .A2(_0226_),
    .A1(_0210_));
 sg13g2_o21ai_1 _2636_ (.B1(_0227_),
    .Y(_0230_),
    .A1(_0209_),
    .A2(_0225_));
 sg13g2_nor3_2 _2637_ (.A(_0209_),
    .B(_0225_),
    .C(_0227_),
    .Y(_0231_));
 sg13g2_nand3_1 _2638_ (.B(_0226_),
    .C(_0228_),
    .A(_0210_),
    .Y(_0232_));
 sg13g2_nor3_1 _2639_ (.A(_1152_),
    .B(_0229_),
    .C(_0231_),
    .Y(_0233_));
 sg13g2_a21oi_1 _2640_ (.A1(_0230_),
    .A2(_0232_),
    .Y(_0234_),
    .B1(_0858_));
 sg13g2_or2_1 _2641_ (.X(_0235_),
    .B(_0234_),
    .A(_0233_));
 sg13g2_o21ai_1 _2642_ (.B1(_0865_),
    .Y(_0236_),
    .A1(_0233_),
    .A2(_0234_));
 sg13g2_nor3_1 _2643_ (.A(net510),
    .B(_0229_),
    .C(_0231_),
    .Y(_0237_));
 sg13g2_nand3_1 _2644_ (.B(_0230_),
    .C(_0232_),
    .A(_0859_),
    .Y(_0238_));
 sg13g2_a21oi_1 _2645_ (.A1(_0230_),
    .A2(_0232_),
    .Y(_0239_),
    .B1(_0859_));
 sg13g2_o21ai_1 _2646_ (.B1(net510),
    .Y(_0240_),
    .A1(_0229_),
    .A2(_0231_));
 sg13g2_o21ai_1 _2647_ (.B1(net507),
    .Y(_0241_),
    .A1(_0237_),
    .A2(_0239_));
 sg13g2_o21ai_1 _2648_ (.B1(_0028_),
    .Y(_0242_),
    .A1(net502),
    .A2(net507));
 sg13g2_a21oi_2 _2649_ (.B1(_0242_),
    .Y(_0243_),
    .A2(_0232_),
    .A1(_0230_));
 sg13g2_mux2_1 _2650_ (.A0(\graphics_engine_1.overlay_creator1.text_demosiine1.y[7] ),
    .A1(_1347_),
    .S(_0912_),
    .X(_0244_));
 sg13g2_xor2_1 _2651_ (.B(_0244_),
    .A(_0243_),
    .X(_0245_));
 sg13g2_xnor2_1 _2652_ (.Y(_0246_),
    .A(_0243_),
    .B(_0244_));
 sg13g2_nor3_2 _2653_ (.A(_0236_),
    .B(_0241_),
    .C(net403),
    .Y(_0247_));
 sg13g2_nand3b_1 _2654_ (.B(_0238_),
    .C(_0240_),
    .Y(_0248_),
    .A_N(net504));
 sg13g2_nor3_2 _2655_ (.A(_0236_),
    .B(net402),
    .C(_0248_),
    .Y(_0249_));
 sg13g2_o21ai_1 _2656_ (.B1(_0028_),
    .Y(_0250_),
    .A1(_0233_),
    .A2(_0234_));
 sg13g2_nand3b_1 _2657_ (.B(_0238_),
    .C(_0240_),
    .Y(_0251_),
    .A_N(net507));
 sg13g2_nand2b_1 _2658_ (.Y(_0252_),
    .B(_0246_),
    .A_N(_0251_));
 sg13g2_o21ai_1 _2659_ (.B1(_0252_),
    .Y(_0253_),
    .A1(_0241_),
    .A2(_0250_));
 sg13g2_a21o_1 _2660_ (.A2(_0248_),
    .A1(_0241_),
    .B1(net402),
    .X(_0254_));
 sg13g2_o21ai_1 _2661_ (.B1(net503),
    .Y(_0255_),
    .A1(_0237_),
    .A2(_0239_));
 sg13g2_a22oi_1 _2662_ (.Y(_0256_),
    .B1(_0246_),
    .B2(net503),
    .A2(net404),
    .A1(_0028_));
 sg13g2_a21o_1 _2663_ (.A2(_0255_),
    .A1(_0248_),
    .B1(_0256_),
    .X(_0257_));
 sg13g2_o21ai_1 _2664_ (.B1(_0257_),
    .Y(_0258_),
    .A1(net404),
    .A2(_0254_));
 sg13g2_nor4_2 _2665_ (.A(_0247_),
    .B(_0249_),
    .C(_0253_),
    .Y(_0259_),
    .D(_0258_));
 sg13g2_nand2_1 _2666_ (.Y(_0260_),
    .A(\graphics_engine_1.anim_2x[0] ),
    .B(\graphics_engine_1.overlay_creator1.text_demosiine1.y[0] ));
 sg13g2_nor2_1 _2667_ (.A(_0259_),
    .B(_0260_),
    .Y(_0261_));
 sg13g2_nor3_2 _2668_ (.A(net1),
    .B(_0259_),
    .C(_0260_),
    .Y(_0262_));
 sg13g2_xor2_1 _2669_ (.B(_0224_),
    .A(_0223_),
    .X(_0263_));
 sg13g2_xnor2_1 _2670_ (.Y(_0264_),
    .A(_0223_),
    .B(_0224_));
 sg13g2_xor2_1 _2671_ (.B(_0219_),
    .A(_0218_),
    .X(_0265_));
 sg13g2_xnor2_1 _2672_ (.Y(_0266_),
    .A(_0218_),
    .B(_0219_));
 sg13g2_o21ai_1 _2673_ (.B1(_0212_),
    .Y(_0267_),
    .A1(_0213_),
    .A2(_0221_));
 sg13g2_and2_1 _2674_ (.A(_0222_),
    .B(_0267_),
    .X(_0268_));
 sg13g2_nand2_2 _2675_ (.Y(_0269_),
    .A(_0222_),
    .B(_0267_));
 sg13g2_xor2_1 _2676_ (.B(\graphics_engine_1.ctr[3] ),
    .A(net487),
    .X(_0270_));
 sg13g2_xnor2_1 _2677_ (.Y(_0271_),
    .A(_0220_),
    .B(_0270_));
 sg13g2_xor2_1 _2678_ (.B(_0270_),
    .A(_0220_),
    .X(_0272_));
 sg13g2_nor2_2 _2679_ (.A(net441),
    .B(net447),
    .Y(_0273_));
 sg13g2_nand2_1 _2680_ (.Y(_0274_),
    .A(net438),
    .B(_0272_));
 sg13g2_nor2_1 _2681_ (.A(net454),
    .B(net446),
    .Y(_0275_));
 sg13g2_nand2_2 _2682_ (.Y(_0276_),
    .A(_0266_),
    .B(_0272_));
 sg13g2_nand2_2 _2683_ (.Y(_0277_),
    .A(net438),
    .B(_0275_));
 sg13g2_nor4_2 _2684_ (.A(_0241_),
    .B(_0246_),
    .C(_0250_),
    .Y(_0278_),
    .D(_0277_));
 sg13g2_nor3_2 _2685_ (.A(_0236_),
    .B(net401),
    .C(_0251_),
    .Y(_0279_));
 sg13g2_xor2_1 _2686_ (.B(_0217_),
    .A(_0216_),
    .X(_0280_));
 sg13g2_xnor2_1 _2687_ (.Y(_0281_),
    .A(_0216_),
    .B(_0217_));
 sg13g2_nor2_2 _2688_ (.A(_0266_),
    .B(_0281_),
    .Y(_0282_));
 sg13g2_nand2_2 _2689_ (.Y(_0283_),
    .A(net454),
    .B(_0280_));
 sg13g2_nor2_2 _2690_ (.A(net440),
    .B(_0272_),
    .Y(_0284_));
 sg13g2_nand2_1 _2691_ (.Y(_0285_),
    .A(net438),
    .B(net446));
 sg13g2_nand3_1 _2692_ (.B(_0283_),
    .C(_0284_),
    .A(_0279_),
    .Y(_0286_));
 sg13g2_nand3_1 _2693_ (.B(_0230_),
    .C(_0232_),
    .A(_0912_),
    .Y(_0287_));
 sg13g2_xnor2_1 _2694_ (.Y(_0288_),
    .A(_0028_),
    .B(_0287_));
 sg13g2_xnor2_1 _2695_ (.Y(_0289_),
    .A(_0865_),
    .B(_0287_));
 sg13g2_nor4_2 _2696_ (.A(_0235_),
    .B(_0241_),
    .C(net402),
    .Y(_0290_),
    .D(_0288_));
 sg13g2_nor2_2 _2697_ (.A(_0274_),
    .B(_0283_),
    .Y(_0291_));
 sg13g2_nor2_1 _2698_ (.A(net454),
    .B(_0285_),
    .Y(_0292_));
 sg13g2_nor2_1 _2699_ (.A(net447),
    .B(_0282_),
    .Y(_0293_));
 sg13g2_nand2_2 _2700_ (.Y(_0294_),
    .A(_0272_),
    .B(_0283_));
 sg13g2_nor2_2 _2701_ (.A(_0266_),
    .B(_0272_),
    .Y(_0295_));
 sg13g2_nand2_2 _2702_ (.Y(_0296_),
    .A(_0265_),
    .B(net447));
 sg13g2_nand2_2 _2703_ (.Y(_0297_),
    .A(_0269_),
    .B(_0296_));
 sg13g2_o21ai_1 _2704_ (.B1(_0290_),
    .Y(_0298_),
    .A1(_0291_),
    .A2(_0292_));
 sg13g2_nor4_2 _2705_ (.A(_0235_),
    .B(net402),
    .C(_0255_),
    .Y(_0299_),
    .D(_0288_));
 sg13g2_nor2_2 _2706_ (.A(net454),
    .B(_0280_),
    .Y(_0300_));
 sg13g2_nand2_2 _2707_ (.Y(_0301_),
    .A(_0266_),
    .B(_0281_));
 sg13g2_nand3_1 _2708_ (.B(_0299_),
    .C(_0301_),
    .A(_0273_),
    .Y(_0302_));
 sg13g2_nor4_2 _2709_ (.A(net404),
    .B(net402),
    .C(_0248_),
    .Y(_0303_),
    .D(_0288_));
 sg13g2_nand2_1 _2710_ (.Y(_0304_),
    .A(net439),
    .B(_0276_));
 sg13g2_nand2_2 _2711_ (.Y(_0305_),
    .A(net438),
    .B(_0300_));
 sg13g2_inv_1 _2712_ (.Y(_0306_),
    .A(_0305_));
 sg13g2_nand2_1 _2713_ (.Y(_0307_),
    .A(net417),
    .B(_0305_));
 sg13g2_nand3_1 _2714_ (.B(_0303_),
    .C(_0307_),
    .A(_0276_),
    .Y(_0308_));
 sg13g2_nand4_1 _2715_ (.B(_0298_),
    .C(_0302_),
    .A(_0286_),
    .Y(_0309_),
    .D(_0308_));
 sg13g2_o21ai_1 _2716_ (.B1(net420),
    .Y(_0310_),
    .A1(_0278_),
    .A2(_0309_));
 sg13g2_nor2_1 _2717_ (.A(net446),
    .B(_0301_),
    .Y(_0311_));
 sg13g2_xnor2_1 _2718_ (.Y(_0312_),
    .A(net447),
    .B(_0300_));
 sg13g2_nand2_1 _2719_ (.Y(_0313_),
    .A(net442),
    .B(_0312_));
 sg13g2_nor3_2 _2720_ (.A(net401),
    .B(_0250_),
    .C(_0251_),
    .Y(_0314_));
 sg13g2_nand2_2 _2721_ (.Y(_0315_),
    .A(net446),
    .B(_0282_));
 sg13g2_and2_1 _2722_ (.A(net439),
    .B(_0315_),
    .X(_0316_));
 sg13g2_nand2_2 _2723_ (.Y(_0317_),
    .A(net439),
    .B(_0315_));
 sg13g2_nand3_1 _2724_ (.B(_0314_),
    .C(_0317_),
    .A(_0313_),
    .Y(_0318_));
 sg13g2_nor2_2 _2725_ (.A(_0269_),
    .B(_0272_),
    .Y(_0319_));
 sg13g2_nand2_1 _2726_ (.Y(_0320_),
    .A(net441),
    .B(net447));
 sg13g2_nor2_2 _2727_ (.A(_0266_),
    .B(_0280_),
    .Y(_0321_));
 sg13g2_nand2_1 _2728_ (.Y(_0322_),
    .A(net454),
    .B(_0281_));
 sg13g2_nand2_2 _2729_ (.Y(_0323_),
    .A(net440),
    .B(_0295_));
 sg13g2_a21oi_1 _2730_ (.A1(_0319_),
    .A2(_0321_),
    .Y(_0324_),
    .B1(net420));
 sg13g2_nor4_2 _2731_ (.A(_0236_),
    .B(net403),
    .C(_0248_),
    .Y(_0325_),
    .D(_0324_));
 sg13g2_nor2_2 _2732_ (.A(net439),
    .B(net446),
    .Y(_0326_));
 sg13g2_nand2_2 _2733_ (.Y(_0327_),
    .A(net440),
    .B(_0272_));
 sg13g2_nor2_2 _2734_ (.A(net438),
    .B(_0276_),
    .Y(_0328_));
 sg13g2_inv_1 _2735_ (.Y(_0329_),
    .A(_0328_));
 sg13g2_nor2_1 _2736_ (.A(net454),
    .B(_0281_),
    .Y(_0330_));
 sg13g2_nand2_2 _2737_ (.Y(_0331_),
    .A(_0266_),
    .B(_0280_));
 sg13g2_nor2_1 _2738_ (.A(net447),
    .B(_0331_),
    .Y(_0332_));
 sg13g2_o21ai_1 _2739_ (.B1(net420),
    .Y(_0333_),
    .A1(net417),
    .A2(_0331_));
 sg13g2_nand2_2 _2740_ (.Y(_0334_),
    .A(net441),
    .B(_0301_));
 sg13g2_nand3_1 _2741_ (.B(net416),
    .C(_0334_),
    .A(_0297_),
    .Y(_0335_));
 sg13g2_nand2b_1 _2742_ (.Y(_0336_),
    .B(_0335_),
    .A_N(_0333_));
 sg13g2_nor3_2 _2743_ (.A(net440),
    .B(net446),
    .C(_0322_),
    .Y(_0337_));
 sg13g2_nor2_1 _2744_ (.A(net423),
    .B(_0337_),
    .Y(_0338_));
 sg13g2_and3_2 _2745_ (.X(_0339_),
    .A(_0317_),
    .B(net416),
    .C(_0334_));
 sg13g2_nand3_1 _2746_ (.B(net416),
    .C(_0334_),
    .A(_0317_),
    .Y(_0340_));
 sg13g2_nor2_1 _2747_ (.A(_0328_),
    .B(_0339_),
    .Y(_0341_));
 sg13g2_and2_1 _2748_ (.A(_0338_),
    .B(_0341_),
    .X(_0342_));
 sg13g2_o21ai_1 _2749_ (.B1(net425),
    .Y(_0343_),
    .A1(_0320_),
    .A2(_0331_));
 sg13g2_nand2_1 _2750_ (.Y(_0344_),
    .A(_0247_),
    .B(_0343_));
 sg13g2_nor4_2 _2751_ (.A(net404),
    .B(net401),
    .C(_0255_),
    .Y(_0345_),
    .D(_0289_));
 sg13g2_inv_1 _2752_ (.Y(_0346_),
    .A(_0345_));
 sg13g2_nand2_1 _2753_ (.Y(_0347_),
    .A(_0301_),
    .B(_0326_));
 sg13g2_nand2_1 _2754_ (.Y(_0348_),
    .A(_0284_),
    .B(_0300_));
 sg13g2_a22oi_1 _2755_ (.Y(_0349_),
    .B1(_0347_),
    .B2(_0348_),
    .A2(_0283_),
    .A1(_0263_));
 sg13g2_nand2_1 _2756_ (.Y(_0350_),
    .A(_0345_),
    .B(_0349_));
 sg13g2_nor4_2 _2757_ (.A(net404),
    .B(_0241_),
    .C(net402),
    .Y(_0351_),
    .D(_0289_));
 sg13g2_nand2_2 _2758_ (.Y(_0352_),
    .A(_0282_),
    .B(_0326_));
 sg13g2_nand2_1 _2759_ (.Y(_0353_),
    .A(net442),
    .B(_0294_));
 sg13g2_nand3_1 _2760_ (.B(_0294_),
    .C(_0296_),
    .A(net441),
    .Y(_0354_));
 sg13g2_a21oi_2 _2761_ (.B1(net425),
    .Y(_0355_),
    .A2(_0321_),
    .A1(_0284_));
 sg13g2_nor2_1 _2762_ (.A(_0327_),
    .B(_0331_),
    .Y(_0356_));
 sg13g2_and2_1 _2763_ (.A(net423),
    .B(_0323_),
    .X(_0357_));
 sg13g2_nor2_2 _2764_ (.A(net420),
    .B(_0356_),
    .Y(_0358_));
 sg13g2_a22oi_1 _2765_ (.Y(_0359_),
    .B1(_0358_),
    .B2(_0323_),
    .A2(_0355_),
    .A1(_0354_));
 sg13g2_nor4_2 _2766_ (.A(net404),
    .B(net402),
    .C(_0251_),
    .Y(_0360_),
    .D(_0289_));
 sg13g2_a21oi_2 _2767_ (.B1(net420),
    .Y(_0361_),
    .A2(_0319_),
    .A1(_0300_));
 sg13g2_nand2_1 _2768_ (.Y(_0362_),
    .A(net442),
    .B(_0293_));
 sg13g2_nor2_2 _2769_ (.A(net423),
    .B(_0291_),
    .Y(_0363_));
 sg13g2_a21oi_1 _2770_ (.A1(_0362_),
    .A2(_0363_),
    .Y(_0364_),
    .B1(_0361_));
 sg13g2_and2_1 _2771_ (.A(net418),
    .B(_0323_),
    .X(_0365_));
 sg13g2_nor4_2 _2772_ (.A(_0241_),
    .B(net401),
    .C(_0250_),
    .Y(_0366_),
    .D(_0365_));
 sg13g2_nand2_1 _2773_ (.Y(_0367_),
    .A(net423),
    .B(_0277_));
 sg13g2_a21oi_1 _2774_ (.A1(_0276_),
    .A2(_0296_),
    .Y(_0368_),
    .B1(_0306_));
 sg13g2_a21o_1 _2775_ (.A2(_0368_),
    .A1(_0334_),
    .B1(_0367_),
    .X(_0369_));
 sg13g2_nor3_2 _2776_ (.A(net422),
    .B(net417),
    .C(_0282_),
    .Y(_0370_));
 sg13g2_nor4_2 _2777_ (.A(net404),
    .B(net402),
    .C(_0251_),
    .Y(_0371_),
    .D(_0288_));
 sg13g2_nor4_2 _2778_ (.A(net404),
    .B(net401),
    .C(_0248_),
    .Y(_0372_),
    .D(_0289_));
 sg13g2_nand2_1 _2779_ (.Y(_0373_),
    .A(_0321_),
    .B(_0326_));
 sg13g2_nor2_2 _2780_ (.A(net439),
    .B(_0315_),
    .Y(_0374_));
 sg13g2_nor2_1 _2781_ (.A(net418),
    .B(_0374_),
    .Y(_0375_));
 sg13g2_nor3_2 _2782_ (.A(net438),
    .B(_0275_),
    .C(_0295_),
    .Y(_0376_));
 sg13g2_nor2_1 _2783_ (.A(_0285_),
    .B(_0331_),
    .Y(_0377_));
 sg13g2_a21oi_1 _2784_ (.A1(_0331_),
    .A2(_0376_),
    .Y(_0378_),
    .B1(_0377_));
 sg13g2_a22oi_1 _2785_ (.Y(_0379_),
    .B1(_0378_),
    .B2(net418),
    .A2(_0375_),
    .A1(_0373_));
 sg13g2_nor2_1 _2786_ (.A(net423),
    .B(_0277_),
    .Y(_0380_));
 sg13g2_nor3_2 _2787_ (.A(net422),
    .B(_0277_),
    .C(_0280_),
    .Y(_0381_));
 sg13g2_nor3_1 _2788_ (.A(_0246_),
    .B(_0248_),
    .C(_0250_),
    .Y(_0382_));
 sg13g2_nor3_2 _2789_ (.A(net401),
    .B(_0250_),
    .C(_0255_),
    .Y(_0383_));
 sg13g2_nand2_1 _2790_ (.Y(_0384_),
    .A(_0283_),
    .B(_0301_));
 sg13g2_nor2_2 _2791_ (.A(_0282_),
    .B(_0300_),
    .Y(_0385_));
 sg13g2_o21ai_1 _2792_ (.B1(net421),
    .Y(_0386_),
    .A1(_0327_),
    .A2(_0384_));
 sg13g2_inv_1 _2793_ (.Y(_0387_),
    .A(_0386_));
 sg13g2_nor2_1 _2794_ (.A(_0374_),
    .B(_0386_),
    .Y(_0388_));
 sg13g2_nand2_1 _2795_ (.Y(_0389_),
    .A(_0284_),
    .B(_0385_));
 sg13g2_a21oi_2 _2796_ (.B1(net421),
    .Y(_0390_),
    .A2(_0385_),
    .A1(_0284_));
 sg13g2_a21oi_1 _2797_ (.A1(_0354_),
    .A2(_0390_),
    .Y(_0391_),
    .B1(_0388_));
 sg13g2_nand2_1 _2798_ (.Y(_0392_),
    .A(_0383_),
    .B(_0391_));
 sg13g2_a21oi_1 _2799_ (.A1(_0276_),
    .A2(_0307_),
    .Y(_0393_),
    .B1(net418));
 sg13g2_or3_2 _2800_ (.A(net403),
    .B(_0248_),
    .C(_0250_),
    .X(_0394_));
 sg13g2_a221oi_1 _2801_ (.B2(_0347_),
    .C1(_0394_),
    .B1(_0393_),
    .A1(net419),
    .Y(_0395_),
    .A2(_0354_));
 sg13g2_nor4_2 _2802_ (.A(_0236_),
    .B(net401),
    .C(_0255_),
    .Y(_0396_),
    .D(_0375_));
 sg13g2_o21ai_1 _2803_ (.B1(net420),
    .Y(_0397_),
    .A1(net441),
    .A2(_0312_));
 sg13g2_a221oi_1 _2804_ (.B2(_0379_),
    .C1(_0395_),
    .B1(_0372_),
    .A1(_0370_),
    .Y(_0398_),
    .A2(_0371_));
 sg13g2_a22oi_1 _2805_ (.Y(_0399_),
    .B1(_0396_),
    .B2(_0397_),
    .A2(_0336_),
    .A1(_0325_));
 sg13g2_o21ai_1 _2806_ (.B1(_0399_),
    .Y(_0400_),
    .A1(_0342_),
    .A2(_0344_));
 sg13g2_a22oi_1 _2807_ (.Y(_0401_),
    .B1(_0366_),
    .B2(_0369_),
    .A2(_0359_),
    .A1(_0351_));
 sg13g2_a22oi_1 _2808_ (.Y(_0402_),
    .B1(_0381_),
    .B2(_0382_),
    .A2(_0364_),
    .A1(_0360_));
 sg13g2_nand4_1 _2809_ (.B(_0350_),
    .C(_0401_),
    .A(_0318_),
    .Y(_0403_),
    .D(_0402_));
 sg13g2_nor2_1 _2810_ (.A(_0400_),
    .B(_0403_),
    .Y(_0404_));
 sg13g2_nand4_1 _2811_ (.B(_0392_),
    .C(_0398_),
    .A(_0310_),
    .Y(_0405_),
    .D(_0404_));
 sg13g2_a21oi_2 _2812_ (.B1(net424),
    .Y(_0406_),
    .A2(_0316_),
    .A1(_0294_));
 sg13g2_o21ai_1 _2813_ (.B1(_0406_),
    .Y(_0407_),
    .A1(net417),
    .A2(_0331_));
 sg13g2_o21ai_1 _2814_ (.B1(net420),
    .Y(_0408_),
    .A1(_0297_),
    .A2(_0332_));
 sg13g2_a22oi_1 _2815_ (.Y(_0409_),
    .B1(_0408_),
    .B2(_0396_),
    .A2(_0407_),
    .A1(_0325_));
 sg13g2_nor2_1 _2816_ (.A(_0343_),
    .B(_0374_),
    .Y(_0410_));
 sg13g2_nor3_1 _2817_ (.A(net423),
    .B(_0284_),
    .C(_0337_),
    .Y(_0411_));
 sg13g2_nor2_1 _2818_ (.A(_0410_),
    .B(_0411_),
    .Y(_0412_));
 sg13g2_o21ai_1 _2819_ (.B1(_0314_),
    .Y(_0413_),
    .A1(_0339_),
    .A2(_0376_));
 sg13g2_nand2_1 _2820_ (.Y(_0414_),
    .A(_0273_),
    .B(_0290_));
 sg13g2_nand3_1 _2821_ (.B(_0279_),
    .C(_0312_),
    .A(net439),
    .Y(_0415_));
 sg13g2_a21oi_1 _2822_ (.A1(_0414_),
    .A2(_0415_),
    .Y(_0416_),
    .B1(net425));
 sg13g2_nand3_1 _2823_ (.B(_0294_),
    .C(_0315_),
    .A(net441),
    .Y(_0417_));
 sg13g2_a22oi_1 _2824_ (.Y(_0418_),
    .B1(_0358_),
    .B2(_0417_),
    .A2(_0355_),
    .A1(_0327_));
 sg13g2_a22oi_1 _2825_ (.Y(_0419_),
    .B1(_0418_),
    .B2(_0351_),
    .A2(_0381_),
    .A1(_0371_));
 sg13g2_o21ai_1 _2826_ (.B1(net424),
    .Y(_0420_),
    .A1(_0300_),
    .A2(net416));
 sg13g2_inv_1 _2827_ (.Y(_0421_),
    .A(_0420_));
 sg13g2_a21oi_1 _2828_ (.A1(_0284_),
    .A2(_0300_),
    .Y(_0422_),
    .B1(net424));
 sg13g2_a21oi_1 _2829_ (.A1(net438),
    .A2(_0295_),
    .Y(_0423_),
    .B1(_0328_));
 sg13g2_a22oi_1 _2830_ (.Y(_0424_),
    .B1(_0422_),
    .B2(_0423_),
    .A2(_0421_),
    .A1(_0352_));
 sg13g2_a21o_1 _2831_ (.A2(_0316_),
    .A1(_0294_),
    .B1(_0367_),
    .X(_0425_));
 sg13g2_and2_1 _2832_ (.A(_0340_),
    .B(_0389_),
    .X(_0426_));
 sg13g2_a22oi_1 _2833_ (.Y(_0427_),
    .B1(_0363_),
    .B2(_0426_),
    .A2(_0361_),
    .A1(_0323_));
 sg13g2_a22oi_1 _2834_ (.Y(_0428_),
    .B1(_0390_),
    .B2(_0327_),
    .A2(_0387_),
    .A1(net416));
 sg13g2_nor2_2 _2835_ (.A(net420),
    .B(_0319_),
    .Y(_0429_));
 sg13g2_nor2_1 _2836_ (.A(_0339_),
    .B(_0377_),
    .Y(_0430_));
 sg13g2_a22oi_1 _2837_ (.Y(_0431_),
    .B1(_0430_),
    .B2(_0387_),
    .A2(_0429_),
    .A1(_0373_));
 sg13g2_a22oi_1 _2838_ (.Y(_0432_),
    .B1(_0330_),
    .B2(net446),
    .A2(_0329_),
    .A1(_0304_));
 sg13g2_nor4_1 _2839_ (.A(net422),
    .B(net438),
    .C(_0321_),
    .D(_0432_),
    .Y(_0433_));
 sg13g2_a21oi_1 _2840_ (.A1(net422),
    .A2(_0432_),
    .Y(_0434_),
    .B1(_0433_));
 sg13g2_o21ai_1 _2841_ (.B1(_0413_),
    .Y(_0435_),
    .A1(_0394_),
    .A2(_0434_));
 sg13g2_a22oi_1 _2842_ (.Y(_0436_),
    .B1(_0424_),
    .B2(_0345_),
    .A2(_0370_),
    .A1(_0303_));
 sg13g2_a22oi_1 _2843_ (.Y(_0437_),
    .B1(_0431_),
    .B2(_0372_),
    .A2(_0427_),
    .A1(_0360_));
 sg13g2_nand3_1 _2844_ (.B(_0436_),
    .C(_0437_),
    .A(_0409_),
    .Y(_0438_));
 sg13g2_a22oi_1 _2845_ (.Y(_0439_),
    .B1(_0412_),
    .B2(_0247_),
    .A2(_0380_),
    .A1(_0299_));
 sg13g2_a22oi_1 _2846_ (.Y(_0440_),
    .B1(_0428_),
    .B2(_0383_),
    .A2(_0425_),
    .A1(_0366_));
 sg13g2_nand3_1 _2847_ (.B(_0439_),
    .C(_0440_),
    .A(_0419_),
    .Y(_0441_));
 sg13g2_or4_1 _2848_ (.A(_0416_),
    .B(_0435_),
    .C(_0438_),
    .D(_0441_),
    .X(_0442_));
 sg13g2_a22oi_1 _2849_ (.Y(_0443_),
    .B1(_0337_),
    .B2(_0371_),
    .A2(_0306_),
    .A1(_0303_));
 sg13g2_a21oi_1 _2850_ (.A1(_0276_),
    .A2(_0322_),
    .Y(_0444_),
    .B1(net440));
 sg13g2_a22oi_1 _2851_ (.Y(_0445_),
    .B1(_0444_),
    .B2(_0279_),
    .A2(_0280_),
    .A1(_0278_));
 sg13g2_a21oi_1 _2852_ (.A1(_0276_),
    .A2(_0331_),
    .Y(_0446_),
    .B1(net441));
 sg13g2_a22oi_1 _2853_ (.Y(_0447_),
    .B1(_0446_),
    .B2(_0290_),
    .A2(_0299_),
    .A1(_0291_));
 sg13g2_nand3_1 _2854_ (.B(_0445_),
    .C(_0447_),
    .A(_0443_),
    .Y(_0448_));
 sg13g2_nand2_1 _2855_ (.Y(_0449_),
    .A(net418),
    .B(_0448_));
 sg13g2_o21ai_1 _2856_ (.B1(_0338_),
    .Y(_0450_),
    .A1(_0293_),
    .A2(_0297_));
 sg13g2_or2_1 _2857_ (.X(_0451_),
    .B(_0450_),
    .A(_0356_));
 sg13g2_nand3_1 _2858_ (.B(_0420_),
    .C(_0451_),
    .A(_0247_),
    .Y(_0452_));
 sg13g2_a21oi_1 _2859_ (.A1(_0373_),
    .A2(_0406_),
    .Y(_0453_),
    .B1(_0429_));
 sg13g2_a21oi_2 _2860_ (.B1(_0339_),
    .Y(_0454_),
    .A2(_0330_),
    .A1(net442));
 sg13g2_a22oi_1 _2861_ (.Y(_0455_),
    .B1(_0355_),
    .B2(_0454_),
    .A2(_0313_),
    .A1(net424));
 sg13g2_nand2_1 _2862_ (.Y(_0456_),
    .A(_0351_),
    .B(_0455_));
 sg13g2_nand2_1 _2863_ (.Y(_0457_),
    .A(net424),
    .B(_0417_));
 sg13g2_o21ai_1 _2864_ (.B1(_0457_),
    .Y(_0458_),
    .A1(net424),
    .A2(_0284_));
 sg13g2_nand2_1 _2865_ (.Y(_0459_),
    .A(_0352_),
    .B(_0458_));
 sg13g2_a21o_1 _2866_ (.A2(_0353_),
    .A1(net418),
    .B1(_0394_),
    .X(_0460_));
 sg13g2_nand3_1 _2867_ (.B(_0352_),
    .C(_0393_),
    .A(_0285_),
    .Y(_0461_));
 sg13g2_nor2b_1 _2868_ (.A(_0460_),
    .B_N(_0461_),
    .Y(_0462_));
 sg13g2_nor2_1 _2869_ (.A(_0376_),
    .B(_0386_),
    .Y(_0463_));
 sg13g2_a21oi_1 _2870_ (.A1(_0390_),
    .A2(_0454_),
    .Y(_0464_),
    .B1(_0463_));
 sg13g2_nand2_1 _2871_ (.Y(_0465_),
    .A(net417),
    .B(_0314_));
 sg13g2_a21o_1 _2872_ (.A2(net440),
    .A1(net418),
    .B1(_0429_),
    .X(_0466_));
 sg13g2_or4_1 _2873_ (.A(_0236_),
    .B(net401),
    .C(_0255_),
    .D(_0466_),
    .X(_0467_));
 sg13g2_a22oi_1 _2874_ (.Y(_0468_),
    .B1(_0465_),
    .B2(_0467_),
    .A2(_0283_),
    .A1(net446));
 sg13g2_nor2_1 _2875_ (.A(_0273_),
    .B(_0301_),
    .Y(_0469_));
 sg13g2_a22oi_1 _2876_ (.Y(_0470_),
    .B1(_0469_),
    .B2(net416),
    .A2(_0385_),
    .A1(_0273_));
 sg13g2_a21oi_1 _2877_ (.A1(_0363_),
    .A2(_0470_),
    .Y(_0471_),
    .B1(_0357_));
 sg13g2_nor2_1 _2878_ (.A(net419),
    .B(_0376_),
    .Y(_0472_));
 sg13g2_a21oi_1 _2879_ (.A1(_0317_),
    .A2(_0334_),
    .Y(_0473_),
    .B1(net424));
 sg13g2_a21oi_1 _2880_ (.A1(_0389_),
    .A2(_0473_),
    .Y(_0474_),
    .B1(_0472_));
 sg13g2_nand3_1 _2881_ (.B(net417),
    .C(_0305_),
    .A(net422),
    .Y(_0475_));
 sg13g2_nand2_1 _2882_ (.Y(_0476_),
    .A(_0366_),
    .B(_0475_));
 sg13g2_nand2_1 _2883_ (.Y(_0477_),
    .A(_0452_),
    .B(_0456_));
 sg13g2_a22oi_1 _2884_ (.Y(_0478_),
    .B1(_0475_),
    .B2(_0366_),
    .A2(_0464_),
    .A1(_0383_));
 sg13g2_a22oi_1 _2885_ (.Y(_0479_),
    .B1(_0459_),
    .B2(_0345_),
    .A2(_0366_),
    .A1(_0311_));
 sg13g2_a22oi_1 _2886_ (.Y(_0480_),
    .B1(_0471_),
    .B2(_0249_),
    .A2(_0382_),
    .A1(_0381_));
 sg13g2_a22oi_1 _2887_ (.Y(_0481_),
    .B1(_0474_),
    .B2(_0372_),
    .A2(_0453_),
    .A1(_0360_));
 sg13g2_nand4_1 _2888_ (.B(_0479_),
    .C(_0480_),
    .A(_0478_),
    .Y(_0482_),
    .D(_0481_));
 sg13g2_nor4_2 _2889_ (.A(_0462_),
    .B(_0468_),
    .C(_0477_),
    .Y(_0483_),
    .D(_0482_));
 sg13g2_nand2_1 _2890_ (.Y(_0484_),
    .A(_0449_),
    .B(_0483_));
 sg13g2_nand3b_1 _2891_ (.B(_0449_),
    .C(_0483_),
    .Y(_0485_),
    .A_N(_0442_));
 sg13g2_nand2_1 _2892_ (.Y(_0486_),
    .A(_0261_),
    .B(_0405_));
 sg13g2_o21ai_1 _2893_ (.B1(_0262_),
    .Y(_0487_),
    .A1(_0405_),
    .A2(_0485_));
 sg13g2_nand3_1 _2894_ (.B(\graphics_engine_1.overlay_creator1.text_demosiine1.y[0] ),
    .C(net5),
    .A(\graphics_engine_1.anim_2x[0] ),
    .Y(_0488_));
 sg13g2_nand2b_1 _2895_ (.Y(_0489_),
    .B(_0208_),
    .A_N(_0488_));
 sg13g2_mux2_1 _2896_ (.A0(_0486_),
    .A1(_0489_),
    .S(_0487_),
    .X(_0490_));
 sg13g2_a221oi_1 _2897_ (.B2(_0490_),
    .C1(_0184_),
    .B1(_0183_),
    .A1(net514),
    .Y(_0491_),
    .A2(_1457_));
 sg13g2_nor2_1 _2898_ (.A(_0867_),
    .B(_0208_),
    .Y(_0492_));
 sg13g2_a21oi_1 _2899_ (.A1(_0025_),
    .A2(_0867_),
    .Y(_0493_),
    .B1(_0492_));
 sg13g2_and3_1 _2900_ (.X(_0494_),
    .A(net514),
    .B(net393),
    .C(_0493_));
 sg13g2_o21ai_1 _2901_ (.B1(net515),
    .Y(_0495_),
    .A1(_0491_),
    .A2(_0494_));
 sg13g2_nor2_1 _2902_ (.A(_0015_),
    .B(_0992_),
    .Y(_0496_));
 sg13g2_nor3_2 _2903_ (.A(\vga_controller_1.y[9] ),
    .B(_0874_),
    .C(_0496_),
    .Y(_0497_));
 sg13g2_or3_1 _2904_ (.A(net515),
    .B(_0491_),
    .C(_0494_),
    .X(_0498_));
 sg13g2_and3_1 _2905_ (.X(uo_out[6]),
    .A(_0495_),
    .B(_0497_),
    .C(_0498_));
 sg13g2_or2_1 _2906_ (.X(_0499_),
    .B(_1404_),
    .A(net3));
 sg13g2_a21oi_1 _2907_ (.A1(net4),
    .A2(_0205_),
    .Y(_0500_),
    .B1(_0499_));
 sg13g2_nand2b_1 _2908_ (.Y(_0501_),
    .B(_0204_),
    .A_N(_0488_));
 sg13g2_mux2_1 _2909_ (.A0(_0486_),
    .A1(_0501_),
    .S(_0487_),
    .X(_0502_));
 sg13g2_a221oi_1 _2910_ (.B2(_0502_),
    .C1(_0184_),
    .B1(_0183_),
    .A1(_0866_),
    .Y(_0503_),
    .A2(net393));
 sg13g2_o21ai_1 _2911_ (.B1(net515),
    .Y(_0504_),
    .A1(_0500_),
    .A2(_0503_));
 sg13g2_or3_1 _2912_ (.A(net515),
    .B(_0500_),
    .C(_0503_),
    .X(_0505_));
 sg13g2_and3_1 _2913_ (.X(uo_out[2]),
    .A(_0497_),
    .B(_0504_),
    .C(_0505_));
 sg13g2_nor2_1 _2914_ (.A(_0194_),
    .B(_0199_),
    .Y(_0506_));
 sg13g2_nor2_1 _2915_ (.A(_0203_),
    .B(_0506_),
    .Y(_0507_));
 sg13g2_a21oi_1 _2916_ (.A1(_0198_),
    .A2(_0507_),
    .Y(_0508_),
    .B1(_0206_));
 sg13g2_or2_1 _2917_ (.X(_0509_),
    .B(_0508_),
    .A(_0488_));
 sg13g2_a21oi_1 _2918_ (.A1(_0338_),
    .A2(_0389_),
    .Y(_0510_),
    .B1(_0344_));
 sg13g2_a21o_1 _2919_ (.A2(_0329_),
    .A1(_0304_),
    .B1(_0385_),
    .X(_0511_));
 sg13g2_a221oi_1 _2920_ (.B2(_0511_),
    .C1(_0394_),
    .B1(_0393_),
    .A1(net419),
    .Y(_0512_),
    .A2(_0354_));
 sg13g2_nand2_1 _2921_ (.Y(_0513_),
    .A(_0305_),
    .B(_0363_));
 sg13g2_nand4_1 _2922_ (.B(_0383_),
    .C(_0385_),
    .A(net417),
    .Y(_0514_),
    .D(_0466_));
 sg13g2_o21ai_1 _2923_ (.B1(_0355_),
    .Y(_0515_),
    .A1(_0327_),
    .A2(_0384_));
 sg13g2_o21ai_1 _2924_ (.B1(_0358_),
    .Y(_0516_),
    .A1(_0265_),
    .A2(net416));
 sg13g2_nand3_1 _2925_ (.B(_0515_),
    .C(_0516_),
    .A(_0351_),
    .Y(_0517_));
 sg13g2_o21ai_1 _2926_ (.B1(_0325_),
    .Y(_0518_),
    .A1(_0292_),
    .A2(_0333_));
 sg13g2_and2_1 _2927_ (.A(_0303_),
    .B(_0380_),
    .X(_0519_));
 sg13g2_o21ai_1 _2928_ (.B1(net419),
    .Y(_0520_),
    .A1(_0328_),
    .A2(_0377_));
 sg13g2_nand4_1 _2929_ (.B(net440),
    .C(_0276_),
    .A(net422),
    .Y(_0521_),
    .D(_0385_));
 sg13g2_nand2_1 _2930_ (.Y(_0522_),
    .A(_0520_),
    .B(_0521_));
 sg13g2_nand3_1 _2931_ (.B(_0273_),
    .C(_0279_),
    .A(net454),
    .Y(_0523_));
 sg13g2_nand3_1 _2932_ (.B(_0290_),
    .C(_0385_),
    .A(_0273_),
    .Y(_0524_));
 sg13g2_a21o_1 _2933_ (.A2(_0524_),
    .A1(_0523_),
    .B1(net423),
    .X(_0525_));
 sg13g2_o21ai_1 _2934_ (.B1(net422),
    .Y(_0526_),
    .A1(net454),
    .A2(net440));
 sg13g2_o21ai_1 _2935_ (.B1(_0363_),
    .Y(_0527_),
    .A1(net441),
    .A2(_0296_));
 sg13g2_nand2b_1 _2936_ (.Y(_0528_),
    .B(_0361_),
    .A_N(_0374_));
 sg13g2_nand3_1 _2937_ (.B(_0527_),
    .C(_0528_),
    .A(_0360_),
    .Y(_0529_));
 sg13g2_a22oi_1 _2938_ (.Y(_0530_),
    .B1(_0526_),
    .B2(_0366_),
    .A2(_0522_),
    .A1(_0372_));
 sg13g2_nand4_1 _2939_ (.B(_0314_),
    .C(_0323_),
    .A(_0297_),
    .Y(_0531_),
    .D(_0384_));
 sg13g2_nand3_1 _2940_ (.B(_0530_),
    .C(_0531_),
    .A(_0514_),
    .Y(_0532_));
 sg13g2_a22oi_1 _2941_ (.Y(_0533_),
    .B1(_0396_),
    .B2(_0513_),
    .A2(_0381_),
    .A1(_0299_));
 sg13g2_nand2_1 _2942_ (.Y(_0534_),
    .A(_0518_),
    .B(_0533_));
 sg13g2_a221oi_1 _2943_ (.B2(_0340_),
    .C1(_0346_),
    .B1(_0422_),
    .A1(_0352_),
    .Y(_0535_),
    .A2(_0357_));
 sg13g2_nor4_1 _2944_ (.A(_0510_),
    .B(_0512_),
    .C(_0519_),
    .D(_0535_),
    .Y(_0536_));
 sg13g2_nand4_1 _2945_ (.B(_0525_),
    .C(_0529_),
    .A(_0517_),
    .Y(_0537_),
    .D(_0536_));
 sg13g2_nor3_1 _2946_ (.A(_0532_),
    .B(_0534_),
    .C(_0537_),
    .Y(_0538_));
 sg13g2_mux2_1 _2947_ (.A0(_0538_),
    .A1(_0509_),
    .S(_0487_),
    .X(_0539_));
 sg13g2_o21ai_1 _2948_ (.B1(net412),
    .Y(_0540_),
    .A1(net434),
    .A2(net444));
 sg13g2_nand3_1 _2949_ (.B(_1623_),
    .C(_0540_),
    .A(_1527_),
    .Y(_0541_));
 sg13g2_nand2b_1 _2950_ (.Y(_0542_),
    .B(_1616_),
    .A_N(_1562_));
 sg13g2_nand3b_1 _2951_ (.B(_0542_),
    .C(_1618_),
    .Y(_0543_),
    .A_N(_1620_));
 sg13g2_nor2_1 _2952_ (.A(_1591_),
    .B(_1599_),
    .Y(_0544_));
 sg13g2_o21ai_1 _2953_ (.B1(_1633_),
    .Y(_0545_),
    .A1(_1515_),
    .A2(net443));
 sg13g2_nand3_1 _2954_ (.B(_1631_),
    .C(_0545_),
    .A(_1629_),
    .Y(_0546_));
 sg13g2_nand3_1 _2955_ (.B(_1577_),
    .C(_1627_),
    .A(_1519_),
    .Y(_0547_));
 sg13g2_a21o_1 _2956_ (.A2(_0544_),
    .A1(_1532_),
    .B1(net409),
    .X(_0548_));
 sg13g2_nand3_1 _2957_ (.B(_0135_),
    .C(_0548_),
    .A(_1638_),
    .Y(_0549_));
 sg13g2_or2_1 _2958_ (.X(_0550_),
    .B(_1643_),
    .A(_1586_));
 sg13g2_nand3_1 _2959_ (.B(_1646_),
    .C(_0550_),
    .A(_1645_),
    .Y(_0551_));
 sg13g2_a22oi_1 _2960_ (.Y(_0552_),
    .B1(_1574_),
    .B2(_1600_),
    .A2(_1572_),
    .A1(_1566_));
 sg13g2_nand2_1 _2961_ (.Y(_0553_),
    .A(_1571_),
    .B(_0552_));
 sg13g2_nor2_1 _2962_ (.A(net429),
    .B(_0544_),
    .Y(_0554_));
 sg13g2_nor4_1 _2963_ (.A(net406),
    .B(net429),
    .C(net405),
    .D(_0544_),
    .Y(_0555_));
 sg13g2_a21oi_1 _2964_ (.A1(_1582_),
    .A2(_1610_),
    .Y(_0556_),
    .B1(net409));
 sg13g2_o21ai_1 _2965_ (.B1(_1604_),
    .Y(_0557_),
    .A1(_0555_),
    .A2(_0556_));
 sg13g2_a221oi_1 _2966_ (.B2(net434),
    .C1(net407),
    .B1(_1594_),
    .A1(_1517_),
    .Y(_0558_),
    .A2(_1556_));
 sg13g2_a21oi_1 _2967_ (.A1(_1514_),
    .A2(_1599_),
    .Y(_0559_),
    .B1(_1569_));
 sg13g2_nor3_1 _2968_ (.A(_1590_),
    .B(_0558_),
    .C(_0559_),
    .Y(_0560_));
 sg13g2_nor2_1 _2969_ (.A(_1549_),
    .B(_1555_),
    .Y(_0561_));
 sg13g2_o21ai_1 _2970_ (.B1(_1580_),
    .Y(_0562_),
    .A1(_1586_),
    .A2(_0561_));
 sg13g2_a22oi_1 _2971_ (.Y(_0563_),
    .B1(_0120_),
    .B2(_1544_),
    .A2(_1597_),
    .A1(_1559_));
 sg13g2_nand2_1 _2972_ (.Y(_0564_),
    .A(_1537_),
    .B(_0563_));
 sg13g2_nand3_1 _2973_ (.B(_1522_),
    .C(_1549_),
    .A(net410),
    .Y(_0565_));
 sg13g2_mux2_1 _2974_ (.A0(net429),
    .A1(_0554_),
    .S(_0565_),
    .X(_0566_));
 sg13g2_nand3_1 _2975_ (.B(_1524_),
    .C(_1578_),
    .A(net443),
    .Y(_0567_));
 sg13g2_a221oi_1 _2976_ (.B2(_1554_),
    .C1(_0560_),
    .B1(_0566_),
    .A1(_1547_),
    .Y(_0568_),
    .A2(_1627_));
 sg13g2_nand3_1 _2977_ (.B(_0547_),
    .C(_0551_),
    .A(_0546_),
    .Y(_0569_));
 sg13g2_nand3_1 _2978_ (.B(_1528_),
    .C(_1579_),
    .A(_1522_),
    .Y(_0570_));
 sg13g2_nand4_1 _2979_ (.B(_0557_),
    .C(_0567_),
    .A(_0543_),
    .Y(_0571_),
    .D(_0570_));
 sg13g2_nand4_1 _2980_ (.B(_0553_),
    .C(_0562_),
    .A(_0549_),
    .Y(_0572_),
    .D(_0564_));
 sg13g2_nor3_1 _2981_ (.A(_0569_),
    .B(_0571_),
    .C(_0572_),
    .Y(_0573_));
 sg13g2_nand3_1 _2982_ (.B(_0568_),
    .C(_0573_),
    .A(_0541_),
    .Y(_0574_));
 sg13g2_a221oi_1 _2983_ (.B2(_1504_),
    .C1(net2),
    .B1(_0574_),
    .A1(_0117_),
    .Y(_0575_),
    .A2(_0182_));
 sg13g2_a221oi_1 _2984_ (.B2(_0539_),
    .C1(_0575_),
    .B1(_0183_),
    .A1(net514),
    .Y(_0576_),
    .A2(net393));
 sg13g2_nor2b_1 _2985_ (.A(net4),
    .B_N(_0026_),
    .Y(_0577_));
 sg13g2_a21oi_1 _2986_ (.A1(net4),
    .A2(_0508_),
    .Y(_0578_),
    .B1(_0577_));
 sg13g2_and3_1 _2987_ (.X(_0579_),
    .A(net514),
    .B(net393),
    .C(_0578_));
 sg13g2_o21ai_1 _2988_ (.B1(net515),
    .Y(_0580_),
    .A1(_0576_),
    .A2(_0579_));
 sg13g2_or3_1 _2989_ (.A(net515),
    .B(_0576_),
    .C(_0579_),
    .X(_0581_));
 sg13g2_and3_1 _2990_ (.X(uo_out[5]),
    .A(_0497_),
    .B(_0580_),
    .C(_0581_));
 sg13g2_nor2_1 _2991_ (.A(_0203_),
    .B(_0488_),
    .Y(_0582_));
 sg13g2_a22oi_1 _2992_ (.Y(_0583_),
    .B1(_0487_),
    .B2(_0582_),
    .A2(_0442_),
    .A1(_0262_));
 sg13g2_a221oi_1 _2993_ (.B2(_0117_),
    .C1(net2),
    .B1(_0182_),
    .A1(_1504_),
    .Y(_0584_),
    .A2(_0181_));
 sg13g2_a221oi_1 _2994_ (.B2(_0583_),
    .C1(_0584_),
    .B1(_0183_),
    .A1(net514),
    .Y(_0585_),
    .A2(net393));
 sg13g2_a21oi_1 _2995_ (.A1(net4),
    .A2(_0203_),
    .Y(_0586_),
    .B1(_0499_));
 sg13g2_o21ai_1 _2996_ (.B1(net516),
    .Y(_0587_),
    .A1(_0585_),
    .A2(_0586_));
 sg13g2_or3_1 _2997_ (.A(net516),
    .B(_0585_),
    .C(_0586_),
    .X(_0588_));
 sg13g2_and3_1 _2998_ (.X(uo_out[1]),
    .A(_0497_),
    .B(_0587_),
    .C(_0588_));
 sg13g2_nand2b_1 _2999_ (.Y(_0589_),
    .B(_0196_),
    .A_N(_0194_));
 sg13g2_xnor2_1 _3000_ (.Y(_0590_),
    .A(_0203_),
    .B(_0506_));
 sg13g2_o21ai_1 _3001_ (.B1(_0590_),
    .Y(_0591_),
    .A1(_0198_),
    .A2(_0589_));
 sg13g2_o21ai_1 _3002_ (.B1(_0591_),
    .Y(_0592_),
    .A1(_0589_),
    .A2(_0590_));
 sg13g2_nor2_1 _3003_ (.A(_0488_),
    .B(_0592_),
    .Y(_0593_));
 sg13g2_nand3_1 _3004_ (.B(_0317_),
    .C(net416),
    .A(_0314_),
    .Y(_0594_));
 sg13g2_nand2_1 _3005_ (.Y(_0595_),
    .A(net418),
    .B(net417));
 sg13g2_a22oi_1 _3006_ (.Y(_0596_),
    .B1(_0595_),
    .B2(_0396_),
    .A2(_0519_),
    .A1(_0281_));
 sg13g2_nand3_1 _3007_ (.B(_0420_),
    .C(_0450_),
    .A(_0247_),
    .Y(_0597_));
 sg13g2_a22oi_1 _3008_ (.Y(_0598_),
    .B1(_0341_),
    .B2(_0355_),
    .A2(_0313_),
    .A1(net424));
 sg13g2_nand2_1 _3009_ (.Y(_0599_),
    .A(_0351_),
    .B(_0598_));
 sg13g2_a21oi_1 _3010_ (.A1(net421),
    .A2(_0426_),
    .Y(_0600_),
    .B1(_0472_));
 sg13g2_a21oi_1 _3011_ (.A1(_0390_),
    .A2(_0423_),
    .Y(_0601_),
    .B1(_0463_));
 sg13g2_a22oi_1 _3012_ (.Y(_0602_),
    .B1(_0601_),
    .B2(_0383_),
    .A2(_0600_),
    .A1(_0372_));
 sg13g2_nand3_1 _3013_ (.B(_0599_),
    .C(_0602_),
    .A(_0597_),
    .Y(_0603_));
 sg13g2_nor2_1 _3014_ (.A(_0406_),
    .B(_0429_),
    .Y(_0604_));
 sg13g2_a22oi_1 _3015_ (.Y(_0605_),
    .B1(_0604_),
    .B2(_0360_),
    .A2(_0380_),
    .A1(_0290_));
 sg13g2_a21oi_1 _3016_ (.A1(net439),
    .A2(_0312_),
    .Y(_0606_),
    .B1(net423));
 sg13g2_nor2_1 _3017_ (.A(_0357_),
    .B(_0606_),
    .Y(_0607_));
 sg13g2_a22oi_1 _3018_ (.Y(_0608_),
    .B1(_0607_),
    .B2(_0249_),
    .A2(_0370_),
    .A1(_0279_));
 sg13g2_nand2_1 _3019_ (.Y(_0609_),
    .A(_0605_),
    .B(_0608_));
 sg13g2_a21oi_1 _3020_ (.A1(net422),
    .A2(_0304_),
    .Y(_0610_),
    .B1(_0460_));
 sg13g2_o21ai_1 _3021_ (.B1(_0476_),
    .Y(_0611_),
    .A1(_0346_),
    .A2(_0458_));
 sg13g2_nor4_1 _3022_ (.A(_0603_),
    .B(_0609_),
    .C(_0610_),
    .D(_0611_),
    .Y(_0612_));
 sg13g2_nand3_1 _3023_ (.B(_0596_),
    .C(_0612_),
    .A(_0594_),
    .Y(_0613_));
 sg13g2_a22oi_1 _3024_ (.Y(_0614_),
    .B1(_0613_),
    .B2(_0262_),
    .A2(_0593_),
    .A1(_0487_));
 sg13g2_a221oi_1 _3025_ (.B2(_0117_),
    .C1(net2),
    .B1(_0182_),
    .A1(_1504_),
    .Y(_0615_),
    .A2(_0149_));
 sg13g2_a221oi_1 _3026_ (.B2(_0614_),
    .C1(_0615_),
    .B1(_0183_),
    .A1(net514),
    .Y(_0616_),
    .A2(net393));
 sg13g2_nor2b_1 _3027_ (.A(net4),
    .B_N(_0027_),
    .Y(_0617_));
 sg13g2_a21oi_1 _3028_ (.A1(net4),
    .A2(_0592_),
    .Y(_0618_),
    .B1(_0617_));
 sg13g2_and3_1 _3029_ (.X(_0619_),
    .A(net514),
    .B(net393),
    .C(_0618_));
 sg13g2_o21ai_1 _3030_ (.B1(net515),
    .Y(_0620_),
    .A1(_0616_),
    .A2(_0619_));
 sg13g2_or3_1 _3031_ (.A(net515),
    .B(_0616_),
    .C(_0619_),
    .X(_0621_));
 sg13g2_and3_1 _3032_ (.X(uo_out[4]),
    .A(_0497_),
    .B(_0620_),
    .C(_0621_));
 sg13g2_nor2_1 _3033_ (.A(_0488_),
    .B(_0590_),
    .Y(_0622_));
 sg13g2_a22oi_1 _3034_ (.Y(_0623_),
    .B1(_0487_),
    .B2(_0622_),
    .A2(_0484_),
    .A1(_0262_));
 sg13g2_a22oi_1 _3035_ (.Y(_0624_),
    .B1(_1581_),
    .B2(_1650_),
    .A2(_1547_),
    .A1(net426));
 sg13g2_nand2_1 _3036_ (.Y(_0625_),
    .A(_1594_),
    .B(_1628_));
 sg13g2_o21ai_1 _3037_ (.B1(_1524_),
    .Y(_0626_),
    .A1(net405),
    .A2(_1599_));
 sg13g2_o21ai_1 _3038_ (.B1(_1528_),
    .Y(_0627_),
    .A1(net405),
    .A2(_1591_));
 sg13g2_nand4_1 _3039_ (.B(_0625_),
    .C(_0626_),
    .A(_0624_),
    .Y(_0628_),
    .D(_0627_));
 sg13g2_nor2b_1 _3040_ (.A(_1573_),
    .B_N(_1577_),
    .Y(_0629_));
 sg13g2_a221oi_1 _3041_ (.B2(net430),
    .C1(_0629_),
    .B1(_0628_),
    .A1(_1615_),
    .Y(_0630_),
    .A2(_1637_));
 sg13g2_nand3_1 _3042_ (.B(_1581_),
    .C(_1623_),
    .A(_1527_),
    .Y(_0631_));
 sg13g2_a21o_1 _3043_ (.A2(_1521_),
    .A1(net430),
    .B1(_1632_),
    .X(_0632_));
 sg13g2_nand3_1 _3044_ (.B(_0135_),
    .C(_0632_),
    .A(_1638_),
    .Y(_0633_));
 sg13g2_nand3_1 _3045_ (.B(_1583_),
    .C(_1633_),
    .A(_1551_),
    .Y(_0634_));
 sg13g2_nand3_1 _3046_ (.B(_1629_),
    .C(_0634_),
    .A(_1598_),
    .Y(_0635_));
 sg13g2_nor2_1 _3047_ (.A(_1586_),
    .B(_1602_),
    .Y(_0636_));
 sg13g2_a22oi_1 _3048_ (.Y(_0637_),
    .B1(_1593_),
    .B2(_0636_),
    .A2(_1572_),
    .A1(_1543_));
 sg13g2_o21ai_1 _3049_ (.B1(_1611_),
    .Y(_0638_),
    .A1(_1532_),
    .A2(_1542_));
 sg13g2_nand3_1 _3050_ (.B(_0119_),
    .C(_0638_),
    .A(_1604_),
    .Y(_0639_));
 sg13g2_nand3_1 _3051_ (.B(_1618_),
    .C(_0138_),
    .A(_1595_),
    .Y(_0640_));
 sg13g2_a21oi_1 _3052_ (.A1(_1605_),
    .A2(_0142_),
    .Y(_0641_),
    .B1(_1630_));
 sg13g2_nor3_1 _3053_ (.A(_1514_),
    .B(_1558_),
    .C(_1643_),
    .Y(_0642_));
 sg13g2_nor2_1 _3054_ (.A(_0126_),
    .B(_0642_),
    .Y(_0643_));
 sg13g2_nand2_1 _3055_ (.Y(_0644_),
    .A(_1539_),
    .B(_1584_));
 sg13g2_nand3_1 _3056_ (.B(_0639_),
    .C(_0640_),
    .A(_0633_),
    .Y(_0645_));
 sg13g2_nand4_1 _3057_ (.B(_0141_),
    .C(_0631_),
    .A(_0139_),
    .Y(_0646_),
    .D(_0635_));
 sg13g2_a22oi_1 _3058_ (.Y(_0647_),
    .B1(_0644_),
    .B2(_1580_),
    .A2(_0133_),
    .A1(_1554_));
 sg13g2_a22oi_1 _3059_ (.Y(_0648_),
    .B1(_0641_),
    .B2(_1571_),
    .A2(_0637_),
    .A1(_1589_));
 sg13g2_o21ai_1 _3060_ (.B1(_1537_),
    .Y(_0649_),
    .A1(_1558_),
    .A2(_0130_));
 sg13g2_a22oi_1 _3061_ (.Y(_0650_),
    .B1(_1645_),
    .B2(_0643_),
    .A2(_1619_),
    .A1(_1554_));
 sg13g2_nand4_1 _3062_ (.B(_0648_),
    .C(_0649_),
    .A(_0647_),
    .Y(_0651_),
    .D(_0650_));
 sg13g2_nor3_1 _3063_ (.A(_0645_),
    .B(_0646_),
    .C(_0651_),
    .Y(_0652_));
 sg13g2_o21ai_1 _3064_ (.B1(_0652_),
    .Y(_0653_),
    .A1(net412),
    .A2(_0630_));
 sg13g2_a221oi_1 _3065_ (.B2(_1504_),
    .C1(net2),
    .B1(_0653_),
    .A1(_0117_),
    .Y(_0654_),
    .A2(_0182_));
 sg13g2_a221oi_1 _3066_ (.B2(_0623_),
    .C1(_0654_),
    .B1(_0183_),
    .A1(net514),
    .Y(_0655_),
    .A2(net393));
 sg13g2_a21oi_1 _3067_ (.A1(net4),
    .A2(_0590_),
    .Y(_0656_),
    .B1(_0499_));
 sg13g2_o21ai_1 _3068_ (.B1(net516),
    .Y(_0657_),
    .A1(_0655_),
    .A2(_0656_));
 sg13g2_or3_1 _3069_ (.A(net516),
    .B(_0655_),
    .C(_0656_),
    .X(_0658_));
 sg13g2_and3_1 _3070_ (.X(uo_out[0]),
    .A(_0497_),
    .B(_0657_),
    .C(_0658_));
 sg13g2_a21oi_1 _3071_ (.A1(\audio_engine_1.seq_ctr[1] ),
    .A2(_0006_),
    .Y(_0659_),
    .B1(\audio_engine_1.seq_ctr[2] ));
 sg13g2_nand2_1 _3072_ (.Y(_0660_),
    .A(\audio_engine_1.seq_ctr[1] ),
    .B(net117));
 sg13g2_a21oi_1 _3073_ (.A1(_0659_),
    .A2(_0660_),
    .Y(_0661_),
    .B1(_0853_));
 sg13g2_nor4_1 _3074_ (.A(\audio_engine_1.seq_ctr[4] ),
    .B(_0868_),
    .C(net7),
    .D(_0661_),
    .Y(audio));
 sg13g2_nand2_1 _3075_ (.Y(_0662_),
    .A(_0034_),
    .B(net6));
 sg13g2_o21ai_1 _3076_ (.B1(_0662_),
    .Y(_0040_),
    .A1(net48),
    .A2(net6));
 sg13g2_and3_2 _3077_ (.X(_0663_),
    .A(\graphics_engine_1.anim_2x[0] ),
    .B(\graphics_engine_1.overlay_creator1.text_demosiine1.x[1] ),
    .C(net495));
 sg13g2_nor2_1 _3078_ (.A(net478),
    .B(net480),
    .Y(_0664_));
 sg13g2_and2_2 _3079_ (.A(net489),
    .B(_0663_),
    .X(_0665_));
 sg13g2_nand2_1 _3080_ (.Y(_0666_),
    .A(net489),
    .B(_0663_));
 sg13g2_nand4_1 _3081_ (.B(\graphics_engine_1.overlay_creator1.text_demosiine1.x[8] ),
    .C(_1183_),
    .A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[9] ),
    .Y(_0667_),
    .D(_0664_));
 sg13g2_nor2_2 _3082_ (.A(_0666_),
    .B(_0667_),
    .Y(_0668_));
 sg13g2_nor2b_1 _3083_ (.A(_0668_),
    .B_N(net521),
    .Y(_0669_));
 sg13g2_nand2b_2 _3084_ (.Y(_0670_),
    .B(net525),
    .A_N(_0668_));
 sg13g2_nand2_1 _3085_ (.Y(_0671_),
    .A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[0] ),
    .B(net435));
 sg13g2_nand3_1 _3086_ (.B(net509),
    .C(net512),
    .A(\vga_controller_1.y[9] ),
    .Y(_0672_));
 sg13g2_nor4_1 _3087_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[8] ),
    .B(\graphics_engine_1.overlay_creator1.text_demosiine1.y[1] ),
    .C(\graphics_engine_1.overlay_creator1.text_demosiine1.y[0] ),
    .D(_0672_),
    .Y(_0673_));
 sg13g2_nand3_1 _3088_ (.B(_0919_),
    .C(_0673_),
    .A(_0912_),
    .Y(_0674_));
 sg13g2_and2_1 _3089_ (.A(net525),
    .B(_0674_),
    .X(_0675_));
 sg13g2_nand2_2 _3090_ (.Y(_0676_),
    .A(_0668_),
    .B(_0675_));
 sg13g2_o21ai_1 _3091_ (.B1(_0671_),
    .Y(_0041_),
    .A1(_0852_),
    .A2(_0676_));
 sg13g2_nand2_1 _3092_ (.Y(_0677_),
    .A(net154),
    .B(net435));
 sg13g2_and2_1 _3093_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[1] ),
    .B(\graphics_engine_1.overlay_creator1.text_demosiine1.y[0] ),
    .X(_0678_));
 sg13g2_xnor2_1 _3094_ (.Y(_0679_),
    .A(net154),
    .B(\graphics_engine_1.overlay_creator1.text_demosiine1.y[0] ));
 sg13g2_o21ai_1 _3095_ (.B1(_0677_),
    .Y(_0042_),
    .A1(_0676_),
    .A2(_0679_));
 sg13g2_nor2_2 _3096_ (.A(net435),
    .B(_0675_),
    .Y(_0680_));
 sg13g2_nand2_1 _3097_ (.Y(_0681_),
    .A(net512),
    .B(_0678_));
 sg13g2_nor2_1 _3098_ (.A(net435),
    .B(_0681_),
    .Y(_0682_));
 sg13g2_a21oi_1 _3099_ (.A1(_0670_),
    .A2(_0678_),
    .Y(_0683_),
    .B1(net512));
 sg13g2_nor3_1 _3100_ (.A(_0680_),
    .B(_0682_),
    .C(_0683_),
    .Y(_0043_));
 sg13g2_nor3_1 _3101_ (.A(_0859_),
    .B(_0680_),
    .C(_0682_),
    .Y(_0684_));
 sg13g2_nor3_1 _3102_ (.A(net510),
    .B(_0676_),
    .C(_0681_),
    .Y(_0685_));
 sg13g2_or2_1 _3103_ (.X(_0044_),
    .B(_0685_),
    .A(_0684_));
 sg13g2_nand3_1 _3104_ (.B(net512),
    .C(_0678_),
    .A(net509),
    .Y(_0686_));
 sg13g2_nor2_1 _3105_ (.A(net435),
    .B(_0686_),
    .Y(_0687_));
 sg13g2_xnor2_1 _3106_ (.Y(_0688_),
    .A(net506),
    .B(_0687_));
 sg13g2_nor2_1 _3107_ (.A(_0680_),
    .B(_0688_),
    .Y(_0045_));
 sg13g2_nand2_1 _3108_ (.Y(_0689_),
    .A(net502),
    .B(net435));
 sg13g2_nor2_1 _3109_ (.A(net503),
    .B(_0686_),
    .Y(_0690_));
 sg13g2_xnor2_1 _3110_ (.Y(_0691_),
    .A(net502),
    .B(_0690_));
 sg13g2_o21ai_1 _3111_ (.B1(_0689_),
    .Y(_0046_),
    .A1(_0676_),
    .A2(_0691_));
 sg13g2_nor4_1 _3112_ (.A(_0873_),
    .B(_1148_),
    .C(net436),
    .D(_0681_),
    .Y(_0692_));
 sg13g2_a21oi_1 _3113_ (.A1(_1149_),
    .A2(_0687_),
    .Y(_0693_),
    .B1(net499));
 sg13g2_nor3_1 _3114_ (.A(_0680_),
    .B(_0692_),
    .C(_0693_),
    .Y(_0047_));
 sg13g2_nand2_1 _3115_ (.Y(_0694_),
    .A(net135),
    .B(net436));
 sg13g2_nor3_1 _3116_ (.A(_0028_),
    .B(_1150_),
    .C(_0686_),
    .Y(_0695_));
 sg13g2_xnor2_1 _3117_ (.Y(_0696_),
    .A(net135),
    .B(_0695_));
 sg13g2_o21ai_1 _3118_ (.B1(_0694_),
    .Y(_0048_),
    .A1(_0676_),
    .A2(_0696_));
 sg13g2_nand3_1 _3119_ (.B(_0874_),
    .C(_0687_),
    .A(net506),
    .Y(_0697_));
 sg13g2_nor4_1 _3120_ (.A(_0871_),
    .B(_1150_),
    .C(net436),
    .D(_0686_),
    .Y(_0698_));
 sg13g2_o21ai_1 _3121_ (.B1(_0697_),
    .Y(_0699_),
    .A1(net160),
    .A2(_0698_));
 sg13g2_nor2_1 _3122_ (.A(_0680_),
    .B(_0699_),
    .Y(_0049_));
 sg13g2_nand2_1 _3123_ (.Y(_0700_),
    .A(net133),
    .B(net435));
 sg13g2_nor4_1 _3124_ (.A(_0022_),
    .B(_0871_),
    .C(_1150_),
    .D(_0686_),
    .Y(_0701_));
 sg13g2_xnor2_1 _3125_ (.Y(_0702_),
    .A(net133),
    .B(_0701_));
 sg13g2_o21ai_1 _3126_ (.B1(_0700_),
    .Y(_0050_),
    .A1(_0676_),
    .A2(_0702_));
 sg13g2_nand2_1 _3127_ (.Y(_0703_),
    .A(\audio_engine_1.freq_synth1.en_synth_clk ),
    .B(\audio_engine_1.counter[10] ));
 sg13g2_nand2_1 _3128_ (.Y(_0704_),
    .A(net59),
    .B(net457));
 sg13g2_nor2_1 _3129_ (.A(\audio_engine_1.seq_time[0] ),
    .B(_0854_),
    .Y(_0705_));
 sg13g2_nand2b_1 _3130_ (.Y(_0706_),
    .B(\audio_engine_1.seq_time[1] ),
    .A_N(net477));
 sg13g2_nand2_1 _3131_ (.Y(_0707_),
    .A(net472),
    .B(net471));
 sg13g2_nor2b_2 _3132_ (.A(net476),
    .B_N(net477),
    .Y(_0708_));
 sg13g2_nand2_1 _3133_ (.Y(_0709_),
    .A(net477),
    .B(_0854_));
 sg13g2_nand3_1 _3134_ (.B(_0707_),
    .C(_0708_),
    .A(net474),
    .Y(_0710_));
 sg13g2_o21ai_1 _3135_ (.B1(_0710_),
    .Y(_0711_),
    .A1(net474),
    .A2(_0706_));
 sg13g2_a21oi_2 _3136_ (.B1(net472),
    .Y(_0712_),
    .A2(_0708_),
    .A1(net474));
 sg13g2_nand2b_1 _3137_ (.Y(_0713_),
    .B(_0706_),
    .A_N(net474));
 sg13g2_o21ai_1 _3138_ (.B1(net472),
    .Y(_0714_),
    .A1(_0708_),
    .A2(_0713_));
 sg13g2_a21oi_1 _3139_ (.A1(net475),
    .A2(_0705_),
    .Y(_0715_),
    .B1(_0714_));
 sg13g2_nor3_2 _3140_ (.A(net474),
    .B(net472),
    .C(_0706_),
    .Y(_0716_));
 sg13g2_o21ai_1 _3141_ (.B1(net471),
    .Y(_0717_),
    .A1(_0712_),
    .A2(_0715_));
 sg13g2_nor2_1 _3142_ (.A(_0716_),
    .B(_0717_),
    .Y(_0718_));
 sg13g2_nor2_1 _3143_ (.A(net477),
    .B(net476),
    .Y(_0719_));
 sg13g2_and2_1 _3144_ (.A(net475),
    .B(_0719_),
    .X(_0720_));
 sg13g2_a21oi_1 _3145_ (.A1(net472),
    .A2(_0720_),
    .Y(_0721_),
    .B1(net471));
 sg13g2_nor3_1 _3146_ (.A(net469),
    .B(_0718_),
    .C(_0721_),
    .Y(_0722_));
 sg13g2_a21oi_1 _3147_ (.A1(net469),
    .A2(_0711_),
    .Y(_0723_),
    .B1(_0722_));
 sg13g2_xor2_1 _3148_ (.B(_0723_),
    .A(\audio_engine_1.freq_synth1.hp_ctr[1] ),
    .X(_0724_));
 sg13g2_nand2_1 _3149_ (.Y(_0725_),
    .A(_0007_),
    .B(_0705_));
 sg13g2_and2_2 _3150_ (.A(net477),
    .B(net476),
    .X(_0726_));
 sg13g2_nand2_1 _3151_ (.Y(_0727_),
    .A(net477),
    .B(net476));
 sg13g2_o21ai_1 _3152_ (.B1(net472),
    .Y(_0728_),
    .A1(net475),
    .A2(_0719_));
 sg13g2_nand2b_1 _3153_ (.Y(_0729_),
    .B(_0727_),
    .A_N(_0728_));
 sg13g2_o21ai_1 _3154_ (.B1(_0729_),
    .Y(_0730_),
    .A1(net472),
    .A2(_0725_));
 sg13g2_a21oi_1 _3155_ (.A1(_0712_),
    .A2(_0725_),
    .Y(_0731_),
    .B1(_0855_));
 sg13g2_nor2b_1 _3156_ (.A(_0715_),
    .B_N(_0731_),
    .Y(_0732_));
 sg13g2_a21oi_1 _3157_ (.A1(_0855_),
    .A2(_0730_),
    .Y(_0733_),
    .B1(_0732_));
 sg13g2_nand3_1 _3158_ (.B(_0007_),
    .C(_0726_),
    .A(net470),
    .Y(_0734_));
 sg13g2_o21ai_1 _3159_ (.B1(_0734_),
    .Y(_0735_),
    .A1(net469),
    .A2(_0733_));
 sg13g2_xnor2_1 _3160_ (.Y(_0736_),
    .A(_0014_),
    .B(_0735_));
 sg13g2_nand2_1 _3161_ (.Y(_0737_),
    .A(_0709_),
    .B(_0713_));
 sg13g2_a21oi_1 _3162_ (.A1(net475),
    .A2(_0029_),
    .Y(_0738_),
    .B1(_0714_));
 sg13g2_nor2_1 _3163_ (.A(net471),
    .B(_0716_),
    .Y(_0739_));
 sg13g2_o21ai_1 _3164_ (.B1(_0739_),
    .Y(_0740_),
    .A1(_0712_),
    .A2(_0738_));
 sg13g2_nor2_1 _3165_ (.A(net469),
    .B(_0718_),
    .Y(_0741_));
 sg13g2_a22oi_1 _3166_ (.Y(_0742_),
    .B1(_0740_),
    .B2(_0741_),
    .A2(_0737_),
    .A1(net469));
 sg13g2_xnor2_1 _3167_ (.Y(_0743_),
    .A(_0010_),
    .B(_0742_));
 sg13g2_nor2_1 _3168_ (.A(_0720_),
    .B(_0726_),
    .Y(_0744_));
 sg13g2_a21oi_1 _3169_ (.A1(net473),
    .A2(_0744_),
    .Y(_0745_),
    .B1(_0712_));
 sg13g2_nor2_1 _3170_ (.A(_0007_),
    .B(_0709_),
    .Y(_0746_));
 sg13g2_nand3b_1 _3171_ (.B(\audio_engine_1.seq_time[4] ),
    .C(_0746_),
    .Y(_0747_),
    .A_N(net473));
 sg13g2_o21ai_1 _3172_ (.B1(_0747_),
    .Y(_0748_),
    .A1(\audio_engine_1.seq_time[4] ),
    .A2(_0745_));
 sg13g2_o21ai_1 _3173_ (.B1(net470),
    .Y(_0749_),
    .A1(net474),
    .A2(_0726_));
 sg13g2_nand2b_1 _3174_ (.Y(_0750_),
    .B(_0726_),
    .A_N(_0707_));
 sg13g2_o21ai_1 _3175_ (.B1(_0749_),
    .Y(_0751_),
    .A1(net474),
    .A2(_0750_));
 sg13g2_a21oi_1 _3176_ (.A1(_0856_),
    .A2(_0748_),
    .Y(_0752_),
    .B1(_0751_));
 sg13g2_xor2_1 _3177_ (.B(_0752_),
    .A(_0011_),
    .X(_0753_));
 sg13g2_nand3_1 _3178_ (.B(net472),
    .C(net471),
    .A(net475),
    .Y(_0754_));
 sg13g2_nor2_1 _3179_ (.A(_0029_),
    .B(_0754_),
    .Y(_0755_));
 sg13g2_a21o_1 _3180_ (.A2(_0754_),
    .A1(_0854_),
    .B1(_0856_),
    .X(_0756_));
 sg13g2_nor2b_1 _3181_ (.A(_0716_),
    .B_N(_0728_),
    .Y(_0757_));
 sg13g2_nor2_1 _3182_ (.A(net469),
    .B(_0757_),
    .Y(_0758_));
 sg13g2_a21oi_1 _3183_ (.A1(net471),
    .A2(_0856_),
    .Y(_0759_),
    .B1(_0758_));
 sg13g2_o21ai_1 _3184_ (.B1(_0759_),
    .Y(_0760_),
    .A1(_0755_),
    .A2(_0756_));
 sg13g2_a21oi_1 _3185_ (.A1(net473),
    .A2(net471),
    .Y(_0761_),
    .B1(net476));
 sg13g2_nand3_1 _3186_ (.B(net470),
    .C(_0750_),
    .A(net474),
    .Y(_0762_));
 sg13g2_nand4_1 _3187_ (.B(_0856_),
    .C(_0008_),
    .A(net473),
    .Y(_0763_),
    .D(_0746_));
 sg13g2_o21ai_1 _3188_ (.B1(_0763_),
    .Y(_0764_),
    .A1(_0761_),
    .A2(_0762_));
 sg13g2_xnor2_1 _3189_ (.Y(_0765_),
    .A(_0009_),
    .B(_0764_));
 sg13g2_xor2_1 _3190_ (.B(_0760_),
    .A(\audio_engine_1.freq_synth1.hp_ctr[0] ),
    .X(_0766_));
 sg13g2_nand3_1 _3191_ (.B(net469),
    .C(_0007_),
    .A(net476),
    .Y(_0767_));
 sg13g2_o21ai_1 _3192_ (.B1(_0758_),
    .Y(_0768_),
    .A1(_0007_),
    .A2(_0727_));
 sg13g2_o21ai_1 _3193_ (.B1(_0767_),
    .Y(_0769_),
    .A1(_0718_),
    .A2(_0768_));
 sg13g2_xnor2_1 _3194_ (.Y(_0770_),
    .A(_0013_),
    .B(_0769_));
 sg13g2_nand4_1 _3195_ (.B(_0765_),
    .C(_0766_),
    .A(_0753_),
    .Y(_0771_),
    .D(_0770_));
 sg13g2_nor4_2 _3196_ (.A(_0724_),
    .B(_0736_),
    .C(_0743_),
    .Y(_0772_),
    .D(_0771_));
 sg13g2_nand3_1 _3197_ (.B(net136),
    .C(net114),
    .A(\audio_engine_1.freq_synth1.hp_ctr[0] ),
    .Y(_0773_));
 sg13g2_o21ai_1 _3198_ (.B1(net60),
    .Y(_0051_),
    .A1(_0772_),
    .A2(_0773_));
 sg13g2_nand2b_1 _3199_ (.Y(_0774_),
    .B(_0772_),
    .A_N(net457));
 sg13g2_xnor2_1 _3200_ (.Y(_0775_),
    .A(\audio_engine_1.freq_synth1.hp_ctr[1] ),
    .B(net137));
 sg13g2_and2_1 _3201_ (.A(_0774_),
    .B(net138),
    .X(_0052_));
 sg13g2_nand2_1 _3202_ (.Y(_0776_),
    .A(\audio_engine_1.freq_synth1.hp_ctr[0] ),
    .B(\audio_engine_1.freq_synth1.hp_ctr[1] ));
 sg13g2_nor2_1 _3203_ (.A(_0009_),
    .B(_0776_),
    .Y(_0777_));
 sg13g2_and2_1 _3204_ (.A(_0009_),
    .B(_0776_),
    .X(_0778_));
 sg13g2_nor4_1 _3205_ (.A(net458),
    .B(_0772_),
    .C(_0777_),
    .D(_0778_),
    .Y(_0779_));
 sg13g2_a21o_1 _3206_ (.A2(net458),
    .A1(net106),
    .B1(_0779_),
    .X(_0053_));
 sg13g2_xor2_1 _3207_ (.B(_0777_),
    .A(_0010_),
    .X(_0780_));
 sg13g2_nor3_1 _3208_ (.A(net458),
    .B(_0772_),
    .C(_0780_),
    .Y(_0781_));
 sg13g2_a21o_1 _3209_ (.A2(net458),
    .A1(net98),
    .B1(_0781_),
    .X(_0054_));
 sg13g2_nand4_1 _3210_ (.B(\audio_engine_1.freq_synth1.hp_ctr[1] ),
    .C(\audio_engine_1.freq_synth1.hp_ctr[2] ),
    .A(\audio_engine_1.freq_synth1.hp_ctr[0] ),
    .Y(_0782_),
    .D(\audio_engine_1.freq_synth1.hp_ctr[3] ));
 sg13g2_nor2_1 _3211_ (.A(_0011_),
    .B(_0782_),
    .Y(_0783_));
 sg13g2_and2_1 _3212_ (.A(_0011_),
    .B(_0782_),
    .X(_0784_));
 sg13g2_nor4_1 _3213_ (.A(net457),
    .B(_0772_),
    .C(_0783_),
    .D(_0784_),
    .Y(_0785_));
 sg13g2_a21o_1 _3214_ (.A2(net457),
    .A1(net96),
    .B1(_0785_),
    .X(_0055_));
 sg13g2_xor2_1 _3215_ (.B(_0783_),
    .A(_0013_),
    .X(_0786_));
 sg13g2_nor3_1 _3216_ (.A(net457),
    .B(_0772_),
    .C(_0786_),
    .Y(_0787_));
 sg13g2_a21o_1 _3217_ (.A2(net457),
    .A1(net102),
    .B1(_0787_),
    .X(_0056_));
 sg13g2_nand2_1 _3218_ (.Y(_0788_),
    .A(\audio_engine_1.freq_synth1.hp_ctr[4] ),
    .B(\audio_engine_1.freq_synth1.hp_ctr[5] ));
 sg13g2_nor2_1 _3219_ (.A(_0782_),
    .B(_0788_),
    .Y(_0789_));
 sg13g2_xor2_1 _3220_ (.B(_0789_),
    .A(_0014_),
    .X(_0790_));
 sg13g2_nor3_1 _3221_ (.A(net457),
    .B(_0772_),
    .C(_0790_),
    .Y(_0791_));
 sg13g2_a21o_1 _3222_ (.A2(net457),
    .A1(net83),
    .B1(_0791_),
    .X(_0057_));
 sg13g2_nand3b_1 _3223_ (.B(\graphics_engine_1.v_sync ),
    .C(\graphics_engine_1.en_v_sync ),
    .Y(_0792_),
    .A_N(net6));
 sg13g2_nor2_1 _3224_ (.A(net56),
    .B(_0792_),
    .Y(_0793_));
 sg13g2_a21oi_1 _3225_ (.A1(_0864_),
    .A2(_0792_),
    .Y(_0058_),
    .B1(net57));
 sg13g2_nor2_1 _3226_ (.A(_0864_),
    .B(_0792_),
    .Y(_0794_));
 sg13g2_and2_1 _3227_ (.A(net127),
    .B(_0794_),
    .X(_0795_));
 sg13g2_xor2_1 _3228_ (.B(_0794_),
    .A(net127),
    .X(_0059_));
 sg13g2_and2_1 _3229_ (.A(net131),
    .B(_0795_),
    .X(_0796_));
 sg13g2_xor2_1 _3230_ (.B(_0795_),
    .A(net131),
    .X(_0060_));
 sg13g2_and2_1 _3231_ (.A(\graphics_engine_1.ctr[3] ),
    .B(_0796_),
    .X(_0797_));
 sg13g2_xor2_1 _3232_ (.B(_0796_),
    .A(net144),
    .X(_0061_));
 sg13g2_and2_1 _3233_ (.A(\graphics_engine_1.ctr[4] ),
    .B(_0797_),
    .X(_0798_));
 sg13g2_xor2_1 _3234_ (.B(_0797_),
    .A(net139),
    .X(_0062_));
 sg13g2_nand2_1 _3235_ (.Y(_0799_),
    .A(\graphics_engine_1.ctr[5] ),
    .B(_0798_));
 sg13g2_xor2_1 _3236_ (.B(_0798_),
    .A(net150),
    .X(_0063_));
 sg13g2_xnor2_1 _3237_ (.Y(_0064_),
    .A(net148),
    .B(_0799_));
 sg13g2_nor2_1 _3238_ (.A(net110),
    .B(_0799_),
    .Y(_0800_));
 sg13g2_xor2_1 _3239_ (.B(_0800_),
    .A(\graphics_engine_1.ctr[7] ),
    .X(_0065_));
 sg13g2_nand4_1 _3240_ (.B(\graphics_engine_1.ctr[6] ),
    .C(\graphics_engine_1.ctr[7] ),
    .A(\graphics_engine_1.ctr[5] ),
    .Y(_0801_),
    .D(_0798_));
 sg13g2_xnor2_1 _3241_ (.Y(_0066_),
    .A(net104),
    .B(_0801_));
 sg13g2_and2_1 _3242_ (.A(net47),
    .B(net435),
    .X(_0067_));
 sg13g2_o21ai_1 _3243_ (.B1(net437),
    .Y(_0802_),
    .A1(\graphics_engine_1.anim_2x[0] ),
    .A2(net129));
 sg13g2_a21oi_1 _3244_ (.A1(\graphics_engine_1.anim_2x[0] ),
    .A2(net129),
    .Y(_0068_),
    .B1(_0802_));
 sg13g2_a21oi_1 _3245_ (.A1(\graphics_engine_1.anim_2x[0] ),
    .A2(net129),
    .Y(_0803_),
    .B1(net495));
 sg13g2_nor3_1 _3246_ (.A(_0663_),
    .B(_0670_),
    .C(net143),
    .Y(_0069_));
 sg13g2_o21ai_1 _3247_ (.B1(net521),
    .Y(_0804_),
    .A1(net489),
    .A2(_0663_));
 sg13g2_nor2_1 _3248_ (.A(_0665_),
    .B(_0804_),
    .Y(_0070_));
 sg13g2_o21ai_1 _3249_ (.B1(net437),
    .Y(_0805_),
    .A1(net485),
    .A2(_0665_));
 sg13g2_a21oi_1 _3250_ (.A1(net485),
    .A2(_0665_),
    .Y(_0071_),
    .B1(_0805_));
 sg13g2_nor2_1 _3251_ (.A(net484),
    .B(_0666_),
    .Y(_0806_));
 sg13g2_xnor2_1 _3252_ (.Y(_0807_),
    .A(net482),
    .B(_0806_));
 sg13g2_nor2_1 _3253_ (.A(_0670_),
    .B(_0807_),
    .Y(_0072_));
 sg13g2_a21oi_1 _3254_ (.A1(_0877_),
    .A2(_0665_),
    .Y(_0808_),
    .B1(net480));
 sg13g2_and2_1 _3255_ (.A(_0879_),
    .B(_0665_),
    .X(_0809_));
 sg13g2_nor3_1 _3256_ (.A(_0670_),
    .B(_0808_),
    .C(_0809_),
    .Y(_0073_));
 sg13g2_nand2_1 _3257_ (.Y(_0810_),
    .A(_1368_),
    .B(_0665_));
 sg13g2_xor2_1 _3258_ (.B(_0810_),
    .A(net478),
    .X(_0811_));
 sg13g2_nor2_1 _3259_ (.A(_0670_),
    .B(_0811_),
    .Y(_0074_));
 sg13g2_nand2_1 _3260_ (.Y(_0812_),
    .A(net478),
    .B(_0809_));
 sg13g2_xor2_1 _3261_ (.B(_0812_),
    .A(net159),
    .X(_0813_));
 sg13g2_nor2_1 _3262_ (.A(_0670_),
    .B(_0813_),
    .Y(_0075_));
 sg13g2_nor2_1 _3263_ (.A(net123),
    .B(_0812_),
    .Y(_0814_));
 sg13g2_o21ai_1 _3264_ (.B1(net437),
    .Y(_0815_),
    .A1(net120),
    .A2(_0814_));
 sg13g2_a21oi_1 _3265_ (.A1(net120),
    .A2(_0814_),
    .Y(_0076_),
    .B1(_0815_));
 sg13g2_mux2_1 _3266_ (.A0(net52),
    .A1(\audio_engine_1.counter[0] ),
    .S(net7),
    .X(_0077_));
 sg13g2_nand2b_1 _3267_ (.Y(_0816_),
    .B(\audio_engine_1.counter[0] ),
    .A_N(net7));
 sg13g2_nand3b_1 _3268_ (.B(\audio_engine_1.counter[1] ),
    .C(\audio_engine_1.counter[0] ),
    .Y(_0817_),
    .A_N(net7));
 sg13g2_xnor2_1 _3269_ (.Y(_0078_),
    .A(net87),
    .B(_0816_));
 sg13g2_nor2_2 _3270_ (.A(_0869_),
    .B(_0817_),
    .Y(_0818_));
 sg13g2_xnor2_1 _3271_ (.Y(_0079_),
    .A(net85),
    .B(_0817_));
 sg13g2_and2_1 _3272_ (.A(\audio_engine_1.counter[3] ),
    .B(_0818_),
    .X(_0819_));
 sg13g2_xor2_1 _3273_ (.B(_0818_),
    .A(net69),
    .X(_0080_));
 sg13g2_and2_1 _3274_ (.A(net65),
    .B(_0819_),
    .X(_0820_));
 sg13g2_xor2_1 _3275_ (.B(_0819_),
    .A(net65),
    .X(_0081_));
 sg13g2_and2_1 _3276_ (.A(\audio_engine_1.counter[5] ),
    .B(_0820_),
    .X(_0821_));
 sg13g2_xor2_1 _3277_ (.B(_0820_),
    .A(net76),
    .X(_0082_));
 sg13g2_and2_1 _3278_ (.A(net74),
    .B(_0821_),
    .X(_0822_));
 sg13g2_xor2_1 _3279_ (.B(_0821_),
    .A(net74),
    .X(_0083_));
 sg13g2_xor2_1 _3280_ (.B(_0822_),
    .A(net89),
    .X(_0084_));
 sg13g2_and3_1 _3281_ (.X(_0823_),
    .A(\audio_engine_1.counter[7] ),
    .B(net71),
    .C(_0822_));
 sg13g2_a21oi_1 _3282_ (.A1(\audio_engine_1.counter[7] ),
    .A2(_0822_),
    .Y(_0824_),
    .B1(net71));
 sg13g2_nor2_1 _3283_ (.A(_0823_),
    .B(net72),
    .Y(_0085_));
 sg13g2_and2_1 _3284_ (.A(net78),
    .B(_0823_),
    .X(_0825_));
 sg13g2_xor2_1 _3285_ (.B(_0823_),
    .A(net78),
    .X(_0086_));
 sg13g2_xor2_1 _3286_ (.B(_0825_),
    .A(net114),
    .X(_0087_));
 sg13g2_nand2_1 _3287_ (.Y(_0826_),
    .A(_0038_),
    .B(_0825_));
 sg13g2_xnor2_1 _3288_ (.Y(_0088_),
    .A(net82),
    .B(_0826_));
 sg13g2_nand3_1 _3289_ (.B(net82),
    .C(_0825_),
    .A(\audio_engine_1.counter[10] ),
    .Y(_0827_));
 sg13g2_nor2_1 _3290_ (.A(_0870_),
    .B(_0827_),
    .Y(_0828_));
 sg13g2_xnor2_1 _3291_ (.Y(_0089_),
    .A(net80),
    .B(_0827_));
 sg13g2_xor2_1 _3292_ (.B(_0828_),
    .A(net93),
    .X(_0090_));
 sg13g2_and3_1 _3293_ (.X(_0829_),
    .A(net93),
    .B(net62),
    .C(_0828_));
 sg13g2_a21oi_1 _3294_ (.A1(\audio_engine_1.counter[13] ),
    .A2(_0828_),
    .Y(_0830_),
    .B1(net62));
 sg13g2_nor2_1 _3295_ (.A(_0829_),
    .B(net63),
    .Y(_0091_));
 sg13g2_xor2_1 _3296_ (.B(_0829_),
    .A(net95),
    .X(_0092_));
 sg13g2_nand3_1 _3297_ (.B(net132),
    .C(_0829_),
    .A(net95),
    .Y(_0831_));
 sg13g2_a21o_1 _3298_ (.A2(_0829_),
    .A1(net95),
    .B1(net132),
    .X(_0832_));
 sg13g2_and2_1 _3299_ (.A(_0831_),
    .B(_0832_),
    .X(_0093_));
 sg13g2_xnor2_1 _3300_ (.Y(_0094_),
    .A(net112),
    .B(_0831_));
 sg13g2_nor2_1 _3301_ (.A(net54),
    .B(_0774_),
    .Y(_0833_));
 sg13g2_a21oi_1 _3302_ (.A1(_0868_),
    .A2(_0774_),
    .Y(_0095_),
    .B1(_0833_));
 sg13g2_nand2_2 _3303_ (.Y(_0834_),
    .A(net112),
    .B(net90));
 sg13g2_nand3_1 _3304_ (.B(net90),
    .C(\audio_engine_1.seq_ctr[0] ),
    .A(\audio_engine_1.counter[17] ),
    .Y(_0835_));
 sg13g2_xnor2_1 _3305_ (.Y(_0096_),
    .A(net117),
    .B(_0834_));
 sg13g2_nor2_1 _3306_ (.A(_0660_),
    .B(_0834_),
    .Y(_0836_));
 sg13g2_xnor2_1 _3307_ (.Y(_0097_),
    .A(\audio_engine_1.seq_ctr[1] ),
    .B(net91));
 sg13g2_nand2_1 _3308_ (.Y(_0837_),
    .A(\audio_engine_1.seq_ctr[2] ),
    .B(_0836_));
 sg13g2_nor3_1 _3309_ (.A(net118),
    .B(\audio_engine_1.seq_ctr[2] ),
    .C(net124),
    .Y(_0838_));
 sg13g2_xnor2_1 _3310_ (.Y(_0839_),
    .A(\audio_engine_1.seq_ctr[2] ),
    .B(_0836_));
 sg13g2_nor2_1 _3311_ (.A(net125),
    .B(_0839_),
    .Y(_0098_));
 sg13g2_xnor2_1 _3312_ (.Y(_0099_),
    .A(net118),
    .B(_0837_));
 sg13g2_nand4_1 _3313_ (.B(\audio_engine_1.seq_ctr[0] ),
    .C(\audio_engine_1.seq_ctr[3] ),
    .A(\audio_engine_1.seq_ctr[1] ),
    .Y(_0840_),
    .D(\audio_engine_1.seq_ctr[2] ));
 sg13g2_xnor2_1 _3314_ (.Y(_0841_),
    .A(_0006_),
    .B(_0840_));
 sg13g2_nor2b_1 _3315_ (.A(_0660_),
    .B_N(_0838_),
    .Y(_0842_));
 sg13g2_nor3_1 _3316_ (.A(_0834_),
    .B(_0841_),
    .C(_0842_),
    .Y(_0843_));
 sg13g2_a21o_1 _3317_ (.A2(_0834_),
    .A1(net100),
    .B1(_0843_),
    .X(_0100_));
 sg13g2_nor2b_2 _3318_ (.A(_0834_),
    .B_N(_0842_),
    .Y(_0844_));
 sg13g2_mux2_1 _3319_ (.A0(net477),
    .A1(net108),
    .S(_0844_),
    .X(_0101_));
 sg13g2_nand2_1 _3320_ (.Y(_0845_),
    .A(net477),
    .B(_0844_));
 sg13g2_a22oi_1 _3321_ (.Y(_0846_),
    .B1(_0845_),
    .B2(net476),
    .A2(_0844_),
    .A1(_0708_));
 sg13g2_inv_1 _3322_ (.Y(_0102_),
    .A(net153));
 sg13g2_nand2_2 _3323_ (.Y(_0847_),
    .A(_0726_),
    .B(_0844_));
 sg13g2_xnor2_1 _3324_ (.Y(_0103_),
    .A(net475),
    .B(_0847_));
 sg13g2_nor2_1 _3325_ (.A(net145),
    .B(_0847_),
    .Y(_0848_));
 sg13g2_xor2_1 _3326_ (.B(_0848_),
    .A(net473),
    .X(_0104_));
 sg13g2_nor2_1 _3327_ (.A(_0757_),
    .B(_0847_),
    .Y(_0849_));
 sg13g2_xnor2_1 _3328_ (.Y(_0105_),
    .A(_0855_),
    .B(_0849_));
 sg13g2_nor3_1 _3329_ (.A(_0008_),
    .B(_0757_),
    .C(_0847_),
    .Y(_0850_));
 sg13g2_xor2_1 _3330_ (.B(_0850_),
    .A(net67),
    .X(_0106_));
 sg13g2_nand3_1 _3331_ (.B(net67),
    .C(_0849_),
    .A(net115),
    .Y(_0851_));
 sg13g2_xnor2_1 _3332_ (.Y(_0107_),
    .A(net470),
    .B(_0851_));
 sg13g2_dfrbp_1 _3333_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net22),
    .D(net122),
    .Q_N(_1687_),
    .Q(h_sync));
 sg13g2_dfrbp_1 _3334_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net525),
    .D(net49),
    .Q_N(\graphics_engine_1.en_v_sync ),
    .Q(_0034_));
 sg13g2_dfrbp_1 _3335_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net43),
    .D(net158),
    .Q_N(_0003_),
    .Q(\graphics_engine_1.v_sync ));
 sg13g2_dfrbp_1 _3336_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net42),
    .D(net51),
    .Q_N(_0033_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.y[0] ));
 sg13g2_dfrbp_1 _3337_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net41),
    .D(net155),
    .Q_N(_1686_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.y[1] ));
 sg13g2_dfrbp_1 _3338_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net40),
    .D(_0043_),
    .Q_N(_1685_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.y[2] ));
 sg13g2_dfrbp_1 _3339_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net39),
    .D(_0044_),
    .Q_N(_1684_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_y[0] ));
 sg13g2_dfrbp_1 _3340_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net38),
    .D(_0045_),
    .Q_N(_0024_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_y[1] ));
 sg13g2_dfrbp_1 _3341_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net37),
    .D(_0046_),
    .Q_N(_0021_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.y[5] ));
 sg13g2_dfrbp_1 _3342_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net36),
    .D(_0047_),
    .Q_N(_0028_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.y[6] ));
 sg13g2_dfrbp_1 _3343_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net35),
    .D(_0048_),
    .Q_N(_0012_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.y[7] ));
 sg13g2_dfrbp_1 _3344_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net34),
    .D(_0049_),
    .Q_N(_0022_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.y[8] ));
 sg13g2_dfrbp_1 _3345_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net33),
    .D(net134),
    .Q_N(_1683_),
    .Q(\vga_controller_1.y[9] ));
 sg13g2_dfrbp_1 _3346_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net520),
    .D(net61),
    .Q_N(\audio_engine_1.freq_synth1.hp_ctr[0] ),
    .Q(_0035_));
 sg13g2_dfrbp_1 _3347_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net520),
    .D(_0052_),
    .Q_N(_1682_),
    .Q(\audio_engine_1.freq_synth1.hp_ctr[1] ));
 sg13g2_dfrbp_1 _3348_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net517),
    .D(net107),
    .Q_N(_0009_),
    .Q(\audio_engine_1.freq_synth1.hp_ctr[2] ));
 sg13g2_dfrbp_1 _3349_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net517),
    .D(net99),
    .Q_N(_0010_),
    .Q(\audio_engine_1.freq_synth1.hp_ctr[3] ));
 sg13g2_dfrbp_1 _3350_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net517),
    .D(net97),
    .Q_N(_0011_),
    .Q(\audio_engine_1.freq_synth1.hp_ctr[4] ));
 sg13g2_dfrbp_1 _3351_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net517),
    .D(net103),
    .Q_N(_0013_),
    .Q(\audio_engine_1.freq_synth1.hp_ctr[5] ));
 sg13g2_dfrbp_1 _3352_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net517),
    .D(net84),
    .Q_N(_0014_),
    .Q(\audio_engine_1.freq_synth1.hp_ctr[6] ));
 sg13g2_dfrbp_1 _3353_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net524),
    .D(net58),
    .Q_N(_0032_),
    .Q(\graphics_engine_1.ctr[0] ));
 sg13g2_dfrbp_1 _3354_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net524),
    .D(net128),
    .Q_N(_1681_),
    .Q(\graphics_engine_1.ctr[1] ));
 sg13g2_dfrbp_1 _3355_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net524),
    .D(_0060_),
    .Q_N(_1680_),
    .Q(\graphics_engine_1.ctr[2] ));
 sg13g2_dfrbp_1 _3356_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net524),
    .D(_0061_),
    .Q_N(_1679_),
    .Q(\graphics_engine_1.ctr[3] ));
 sg13g2_dfrbp_1 _3357_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net524),
    .D(net140),
    .Q_N(_1678_),
    .Q(\graphics_engine_1.ctr[4] ));
 sg13g2_dfrbp_1 _3358_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net524),
    .D(net151),
    .Q_N(_0025_),
    .Q(\graphics_engine_1.ctr[5] ));
 sg13g2_dfrbp_1 _3359_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net524),
    .D(net149),
    .Q_N(_0026_),
    .Q(\graphics_engine_1.ctr[6] ));
 sg13g2_dfrbp_1 _3360_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net524),
    .D(net111),
    .Q_N(_0027_),
    .Q(\graphics_engine_1.ctr[7] ));
 sg13g2_dfrbp_1 _3361_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net523),
    .D(net105),
    .Q_N(_1677_),
    .Q(\graphics_engine_1.ctr[8] ));
 sg13g2_dfrbp_1 _3362_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net32),
    .D(_0067_),
    .Q_N(_0031_),
    .Q(\graphics_engine_1.anim_2x[0] ));
 sg13g2_dfrbp_1 _3363_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net31),
    .D(net130),
    .Q_N(_1676_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.x[1] ));
 sg13g2_dfrbp_1 _3364_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net30),
    .D(_0069_),
    .Q_N(_1675_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.x[2] ));
 sg13g2_dfrbp_1 _3365_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net29),
    .D(_0070_),
    .Q_N(_0020_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_x[0] ));
 sg13g2_dfrbp_1 _3366_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net28),
    .D(_0071_),
    .Q_N(_0019_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.x[4] ));
 sg13g2_dfrbp_1 _3367_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net27),
    .D(_0072_),
    .Q_N(_0023_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.x[5] ));
 sg13g2_dfrbp_1 _3368_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net26),
    .D(_0073_),
    .Q_N(_0018_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.x[6] ));
 sg13g2_dfrbp_1 _3369_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net25),
    .D(_0074_),
    .Q_N(_0017_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.x[7] ));
 sg13g2_dfrbp_1 _3370_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net24),
    .D(_0075_),
    .Q_N(_0016_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.x[8] ));
 sg13g2_dfrbp_1 _3371_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net23),
    .D(_0076_),
    .Q_N(_0015_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.x[9] ));
 sg13g2_dfrbp_1 _3372_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net517),
    .D(_0038_),
    .Q_N(\audio_engine_1.freq_synth1.en_synth_clk ),
    .Q(_0036_));
 sg13g2_dfrbp_1 _3373_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net523),
    .D(net53),
    .Q_N(_0030_),
    .Q(\audio_engine_1.counter[0] ));
 sg13g2_dfrbp_1 _3374_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net523),
    .D(net88),
    .Q_N(_1674_),
    .Q(\audio_engine_1.counter[1] ));
 sg13g2_dfrbp_1 _3375_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net522),
    .D(net86),
    .Q_N(_1673_),
    .Q(\audio_engine_1.counter[2] ));
 sg13g2_dfrbp_1 _3376_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net522),
    .D(net70),
    .Q_N(_1672_),
    .Q(\audio_engine_1.counter[3] ));
 sg13g2_dfrbp_1 _3377_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net522),
    .D(net66),
    .Q_N(_1671_),
    .Q(\audio_engine_1.counter[4] ));
 sg13g2_dfrbp_1 _3378_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net522),
    .D(net77),
    .Q_N(_1670_),
    .Q(\audio_engine_1.counter[5] ));
 sg13g2_dfrbp_1 _3379_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net518),
    .D(net75),
    .Q_N(_1669_),
    .Q(\audio_engine_1.counter[6] ));
 sg13g2_dfrbp_1 _3380_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net518),
    .D(_0084_),
    .Q_N(_1668_),
    .Q(\audio_engine_1.counter[7] ));
 sg13g2_dfrbp_1 _3381_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net518),
    .D(net73),
    .Q_N(_1667_),
    .Q(\audio_engine_1.counter[8] ));
 sg13g2_dfrbp_1 _3382_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net518),
    .D(net79),
    .Q_N(_1666_),
    .Q(\audio_engine_1.counter[9] ));
 sg13g2_dfrbp_1 _3383_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net517),
    .D(_0087_),
    .Q_N(_0001_),
    .Q(\audio_engine_1.counter[10] ));
 sg13g2_dfrbp_1 _3384_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net518),
    .D(_0088_),
    .Q_N(_1665_),
    .Q(\audio_engine_1.counter[11] ));
 sg13g2_dfrbp_1 _3385_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net518),
    .D(net81),
    .Q_N(_1664_),
    .Q(\audio_engine_1.counter[12] ));
 sg13g2_dfrbp_1 _3386_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net519),
    .D(net94),
    .Q_N(_1663_),
    .Q(\audio_engine_1.counter[13] ));
 sg13g2_dfrbp_1 _3387_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net518),
    .D(net64),
    .Q_N(_1662_),
    .Q(\audio_engine_1.counter[14] ));
 sg13g2_dfrbp_1 _3388_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net519),
    .D(_0092_),
    .Q_N(_1661_),
    .Q(\audio_engine_1.counter[15] ));
 sg13g2_dfrbp_1 _3389_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net519),
    .D(_0093_),
    .Q_N(_1660_),
    .Q(\audio_engine_1.counter[16] ));
 sg13g2_dfrbp_1 _3390_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net519),
    .D(net113),
    .Q_N(_0000_),
    .Q(\audio_engine_1.counter[17] ));
 sg13g2_dfrbp_1 _3391_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net519),
    .D(net55),
    .Q_N(_0002_),
    .Q(\audio_engine_1.freq_synth1.audio_reg ));
 sg13g2_dfrbp_1 _3392_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net518),
    .D(_0096_),
    .Q_N(_1659_),
    .Q(\audio_engine_1.seq_ctr[0] ));
 sg13g2_dfrbp_1 _3393_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net522),
    .D(net92),
    .Q_N(_1658_),
    .Q(\audio_engine_1.seq_ctr[1] ));
 sg13g2_dfrbp_1 _3394_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net522),
    .D(net126),
    .Q_N(_1657_),
    .Q(\audio_engine_1.seq_ctr[2] ));
 sg13g2_dfrbp_1 _3395_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net522),
    .D(net119),
    .Q_N(_1656_),
    .Q(\audio_engine_1.seq_ctr[3] ));
 sg13g2_dfrbp_1 _3396_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net522),
    .D(net101),
    .Q_N(_0006_),
    .Q(\audio_engine_1.seq_ctr[4] ));
 sg13g2_dfrbp_1 _3397_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net519),
    .D(_0039_),
    .Q_N(\audio_engine_1.en_seq_clk ),
    .Q(_0037_));
 sg13g2_dfrbp_1 _3398_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net517),
    .D(net109),
    .Q_N(_0029_),
    .Q(\audio_engine_1.seq_time[0] ));
 sg13g2_dfrbp_1 _3399_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net521),
    .D(_0102_),
    .Q_N(_1655_),
    .Q(\audio_engine_1.seq_time[1] ));
 sg13g2_dfrbp_1 _3400_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net526),
    .D(_0103_),
    .Q_N(_0007_),
    .Q(\audio_engine_1.seq_time[2] ));
 sg13g2_dfrbp_1 _3401_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net521),
    .D(net146),
    .Q_N(_1654_),
    .Q(\audio_engine_1.seq_time[3] ));
 sg13g2_dfrbp_1 _3402_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net521),
    .D(_0105_),
    .Q_N(_0008_),
    .Q(\audio_engine_1.seq_time[4] ));
 sg13g2_dfrbp_1 _3403_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net521),
    .D(net68),
    .Q_N(_1653_),
    .Q(\audio_engine_1.seq_time[5] ));
 sg13g2_dfrbp_1 _3404_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net521),
    .D(net116),
    .Q_N(_1652_),
    .Q(\audio_engine_1.seq_time[6] ));
 sg13g2_tiehi _3371__23 (.L_HI(net23));
 sg13g2_tiehi _3370__24 (.L_HI(net24));
 sg13g2_tiehi _3369__25 (.L_HI(net25));
 sg13g2_tiehi _3368__26 (.L_HI(net26));
 sg13g2_tiehi _3367__27 (.L_HI(net27));
 sg13g2_tiehi _3366__28 (.L_HI(net28));
 sg13g2_tiehi _3365__29 (.L_HI(net29));
 sg13g2_tiehi _3364__30 (.L_HI(net30));
 sg13g2_tiehi _3363__31 (.L_HI(net31));
 sg13g2_tiehi _3362__32 (.L_HI(net32));
 sg13g2_tiehi _3345__33 (.L_HI(net33));
 sg13g2_tiehi _3344__34 (.L_HI(net34));
 sg13g2_tiehi _3343__35 (.L_HI(net35));
 sg13g2_tiehi _3342__36 (.L_HI(net36));
 sg13g2_tiehi _3341__37 (.L_HI(net37));
 sg13g2_tiehi _3340__38 (.L_HI(net38));
 sg13g2_tiehi _3339__39 (.L_HI(net39));
 sg13g2_tiehi _3338__40 (.L_HI(net40));
 sg13g2_tiehi _3337__41 (.L_HI(net41));
 sg13g2_tiehi _3336__42 (.L_HI(net42));
 sg13g2_tiehi _3335__43 (.L_HI(net43));
 sg13g2_tiehi tt_um_demosiine_sda_44 (.L_HI(net44));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_demosiine_sda_9 (.L_LO(net9));
 sg13g2_tielo tt_um_demosiine_sda_10 (.L_LO(net10));
 sg13g2_tielo tt_um_demosiine_sda_11 (.L_LO(net11));
 sg13g2_tielo tt_um_demosiine_sda_12 (.L_LO(net12));
 sg13g2_tielo tt_um_demosiine_sda_13 (.L_LO(net13));
 sg13g2_tielo tt_um_demosiine_sda_14 (.L_LO(net14));
 sg13g2_tielo tt_um_demosiine_sda_15 (.L_LO(net15));
 sg13g2_tielo tt_um_demosiine_sda_16 (.L_LO(net16));
 sg13g2_tielo tt_um_demosiine_sda_17 (.L_LO(net17));
 sg13g2_tielo tt_um_demosiine_sda_18 (.L_LO(net18));
 sg13g2_tielo tt_um_demosiine_sda_19 (.L_LO(net19));
 sg13g2_tielo tt_um_demosiine_sda_20 (.L_LO(net20));
 sg13g2_tielo tt_um_demosiine_sda_21 (.L_LO(net21));
 sg13g2_tiehi _3333__22 (.L_HI(net22));
 sg13g2_buf_2 _3442_ (.A(audio),
    .X(uio_out[7]));
 sg13g2_buf_1 _3443_ (.A(\graphics_engine_1.v_sync ),
    .X(uo_out[3]));
 sg13g2_buf_2 _3444_ (.A(h_sync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout393 (.A(_1457_),
    .X(net393));
 sg13g2_buf_4 fanout394 (.X(net394),
    .A(net396));
 sg13g2_buf_2 fanout395 (.A(net396),
    .X(net395));
 sg13g2_buf_4 fanout396 (.X(net396),
    .A(_1503_));
 sg13g2_buf_4 fanout397 (.X(net397),
    .A(_1494_));
 sg13g2_buf_4 fanout398 (.X(net398),
    .A(_1493_));
 sg13g2_buf_4 fanout399 (.X(net399),
    .A(_1491_));
 sg13g2_buf_4 fanout400 (.X(net400),
    .A(_1490_));
 sg13g2_buf_4 fanout401 (.X(net401),
    .A(net403));
 sg13g2_buf_4 fanout402 (.X(net402),
    .A(net403));
 sg13g2_buf_2 fanout403 (.A(_0245_),
    .X(net403));
 sg13g2_buf_4 fanout404 (.X(net404),
    .A(_0235_));
 sg13g2_buf_2 fanout405 (.A(_1548_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(net408),
    .X(net406));
 sg13g2_buf_1 fanout407 (.A(net408),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_1506_),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(net411),
    .X(net409));
 sg13g2_buf_1 fanout410 (.A(net411),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(_1505_),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(net414),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(net414),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_1505_),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_1053_),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(_0320_),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(_0274_),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(net421),
    .X(net418));
 sg13g2_buf_1 fanout419 (.A(net421),
    .X(net419));
 sg13g2_buf_4 fanout420 (.X(net420),
    .A(net421));
 sg13g2_buf_2 fanout421 (.A(_0264_),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(_0263_),
    .X(net422));
 sg13g2_buf_2 fanout423 (.A(net425),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(net425),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(_0263_),
    .X(net425));
 sg13g2_buf_4 fanout426 (.X(net426),
    .A(_1540_));
 sg13g2_buf_4 fanout427 (.X(net427),
    .A(net428));
 sg13g2_buf_2 fanout428 (.A(_1513_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(net431),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(net431),
    .X(net430));
 sg13g2_buf_4 fanout431 (.X(net431),
    .A(_1508_));
 sg13g2_buf_2 fanout432 (.A(net433),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(net434),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(_1507_),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(net436),
    .X(net435));
 sg13g2_buf_1 fanout436 (.A(net437),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(_0669_),
    .X(net437));
 sg13g2_buf_2 fanout438 (.A(net439),
    .X(net438));
 sg13g2_buf_4 fanout439 (.X(net439),
    .A(_0269_));
 sg13g2_buf_4 fanout440 (.X(net440),
    .A(net442));
 sg13g2_buf_4 fanout441 (.X(net441),
    .A(net442));
 sg13g2_buf_4 fanout442 (.X(net442),
    .A(_0268_));
 sg13g2_buf_4 fanout443 (.X(net443),
    .A(net444));
 sg13g2_buf_2 fanout444 (.A(_1516_),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(_1063_),
    .X(net445));
 sg13g2_buf_4 fanout446 (.X(net446),
    .A(_0271_));
 sg13g2_buf_2 fanout447 (.A(_0271_),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_1189_),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(_0975_),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(_0931_),
    .X(net450));
 sg13g2_buf_4 fanout451 (.X(net451),
    .A(_0898_));
 sg13g2_buf_2 fanout452 (.A(_0896_),
    .X(net452));
 sg13g2_buf_1 fanout453 (.A(_0896_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_0265_),
    .X(net454));
 sg13g2_buf_4 fanout455 (.X(net455),
    .A(_0923_));
 sg13g2_buf_2 fanout456 (.A(_1184_),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(_0703_),
    .X(net457));
 sg13g2_buf_1 fanout458 (.A(_0703_),
    .X(net458));
 sg13g2_buf_4 fanout459 (.X(net459),
    .A(_1144_));
 sg13g2_buf_2 fanout460 (.A(net461),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(_0940_),
    .X(net461));
 sg13g2_buf_1 fanout462 (.A(_0940_),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(net465),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(net465),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(_0939_),
    .X(net465));
 sg13g2_buf_4 fanout466 (.X(net466),
    .A(_0863_));
 sg13g2_buf_2 fanout467 (.A(_0863_),
    .X(net467));
 sg13g2_buf_4 fanout468 (.X(net468),
    .A(_0860_));
 sg13g2_buf_2 fanout469 (.A(net470),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(\audio_engine_1.seq_time[6] ),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(\audio_engine_1.seq_time[4] ),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(\audio_engine_1.seq_time[3] ),
    .X(net472));
 sg13g2_buf_1 fanout473 (.A(\audio_engine_1.seq_time[3] ),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(net475),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(net141),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(net152),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(\audio_engine_1.seq_time[0] ),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(net161),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[7] ),
    .X(net479));
 sg13g2_buf_4 fanout480 (.X(net480),
    .A(net481));
 sg13g2_buf_4 fanout481 (.X(net481),
    .A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[6] ));
 sg13g2_buf_4 fanout482 (.X(net482),
    .A(net156));
 sg13g2_buf_2 fanout483 (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[5] ),
    .X(net483));
 sg13g2_buf_4 fanout484 (.X(net484),
    .A(_0019_));
 sg13g2_buf_2 fanout485 (.A(net487),
    .X(net485));
 sg13g2_buf_1 fanout486 (.A(net487),
    .X(net486));
 sg13g2_buf_4 fanout487 (.X(net487),
    .A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[4] ));
 sg13g2_buf_2 fanout488 (.A(_0020_),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(net492),
    .X(net489));
 sg13g2_buf_1 fanout490 (.A(net492),
    .X(net490));
 sg13g2_buf_4 fanout491 (.X(net491),
    .A(net492));
 sg13g2_buf_2 fanout492 (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_x[0] ),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_x[0] ),
    .X(net493));
 sg13g2_buf_1 fanout494 (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_x[0] ),
    .X(net494));
 sg13g2_buf_4 fanout495 (.X(net495),
    .A(net142));
 sg13g2_buf_1 fanout496 (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[2] ),
    .X(net496));
 sg13g2_buf_4 fanout497 (.X(net497),
    .A(_0012_));
 sg13g2_buf_2 fanout498 (.A(net500),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(net500),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[6] ),
    .X(net500));
 sg13g2_buf_4 fanout501 (.X(net501),
    .A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[5] ));
 sg13g2_buf_2 fanout502 (.A(net147),
    .X(net502));
 sg13g2_buf_4 fanout503 (.X(net503),
    .A(net504));
 sg13g2_buf_2 fanout504 (.A(_0024_),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(net507),
    .X(net505));
 sg13g2_buf_4 fanout506 (.X(net506),
    .A(net507));
 sg13g2_buf_4 fanout507 (.X(net507),
    .A(\graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_y[1] ));
 sg13g2_buf_4 fanout508 (.X(net508),
    .A(net511));
 sg13g2_buf_4 fanout509 (.X(net509),
    .A(net510));
 sg13g2_buf_2 fanout510 (.A(net511),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_y[0] ),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(net513),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[2] ),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(_0866_),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(ui_in[0]),
    .X(net515));
 sg13g2_buf_1 fanout516 (.A(ui_in[0]),
    .X(net516));
 sg13g2_buf_4 fanout517 (.X(net517),
    .A(net520));
 sg13g2_buf_4 fanout518 (.X(net518),
    .A(net519));
 sg13g2_buf_4 fanout519 (.X(net519),
    .A(net520));
 sg13g2_buf_2 fanout520 (.A(net521),
    .X(net520));
 sg13g2_buf_4 fanout521 (.X(net521),
    .A(net526));
 sg13g2_buf_4 fanout522 (.X(net522),
    .A(net523));
 sg13g2_buf_2 fanout523 (.A(net526),
    .X(net523));
 sg13g2_buf_4 fanout524 (.X(net524),
    .A(net525));
 sg13g2_buf_4 fanout525 (.X(net525),
    .A(net526));
 sg13g2_buf_4 fanout526 (.X(net526),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[4]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[5]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[6]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[7]),
    .X(net7));
 sg13g2_tielo tt_um_demosiine_sda_8 (.L_LO(net8));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0000_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0001_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0031_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0003_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0040_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0033_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0041_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0030_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0077_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0002_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0095_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0032_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0793_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0058_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0035_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0704_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0051_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold18 (.A(\audio_engine_1.counter[14] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0830_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0091_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold21 (.A(\audio_engine_1.counter[4] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0081_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold23 (.A(\audio_engine_1.seq_time[5] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0106_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold25 (.A(\audio_engine_1.counter[3] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0080_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold27 (.A(\audio_engine_1.counter[8] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0824_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0085_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold30 (.A(\audio_engine_1.counter[6] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0083_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold32 (.A(\audio_engine_1.counter[5] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0082_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold34 (.A(\audio_engine_1.counter[9] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0086_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold36 (.A(\audio_engine_1.counter[12] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0089_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold38 (.A(\audio_engine_1.counter[11] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold39 (.A(\audio_engine_1.freq_synth1.hp_ctr[6] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0057_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold41 (.A(\audio_engine_1.counter[2] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0079_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold43 (.A(\audio_engine_1.counter[1] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0078_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold45 (.A(\audio_engine_1.counter[7] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold46 (.A(\audio_engine_1.en_seq_clk ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0835_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0097_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold49 (.A(\audio_engine_1.counter[13] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0090_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold51 (.A(\audio_engine_1.counter[15] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold52 (.A(\audio_engine_1.freq_synth1.hp_ctr[4] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0055_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold54 (.A(\audio_engine_1.freq_synth1.hp_ctr[3] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0054_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold56 (.A(\audio_engine_1.seq_ctr[4] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0100_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold58 (.A(\audio_engine_1.freq_synth1.hp_ctr[5] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0056_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold60 (.A(\graphics_engine_1.ctr[8] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0066_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold62 (.A(\audio_engine_1.freq_synth1.hp_ctr[2] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0053_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0029_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0101_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0026_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0065_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold68 (.A(\audio_engine_1.counter[17] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0094_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold70 (.A(\audio_engine_1.counter[10] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold71 (.A(\audio_engine_1.seq_time[4] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0107_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold73 (.A(\audio_engine_1.seq_ctr[0] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold74 (.A(\audio_engine_1.seq_ctr[3] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0099_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold76 (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[9] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0887_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0004_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0016_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0006_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0838_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0098_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold83 (.A(\graphics_engine_1.ctr[1] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0059_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold85 (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[1] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0068_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold87 (.A(\graphics_engine_1.ctr[2] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold88 (.A(\audio_engine_1.counter[16] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold89 (.A(\vga_controller_1.y[9] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0050_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold91 (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[7] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold92 (.A(\audio_engine_1.freq_synth1.en_synth_clk ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0773_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0775_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold95 (.A(\graphics_engine_1.ctr[4] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0062_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold97 (.A(\audio_engine_1.seq_time[2] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold98 (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[2] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0803_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold100 (.A(\graphics_engine_1.ctr[3] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0007_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0104_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold103 (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[5] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold104 (.A(\graphics_engine_1.ctr[6] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0064_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold106 (.A(\graphics_engine_1.ctr[5] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0063_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold108 (.A(\audio_engine_1.seq_time[1] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0846_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold110 (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[1] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0042_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold112 (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[5] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold113 (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[7] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0005_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold115 (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[8] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold116 (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[8] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold117 (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[7] ),
    .X(net161));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_fill_2 FILLER_0_28 ();
 sg13g2_fill_2 FILLER_0_56 ();
 sg13g2_fill_1 FILLER_0_58 ();
 sg13g2_fill_2 FILLER_0_69 ();
 sg13g2_decap_8 FILLER_0_100 ();
 sg13g2_decap_8 FILLER_0_107 ();
 sg13g2_decap_8 FILLER_0_114 ();
 sg13g2_decap_8 FILLER_0_121 ();
 sg13g2_fill_1 FILLER_0_128 ();
 sg13g2_decap_4 FILLER_0_134 ();
 sg13g2_fill_2 FILLER_0_138 ();
 sg13g2_decap_8 FILLER_0_144 ();
 sg13g2_decap_8 FILLER_0_151 ();
 sg13g2_decap_8 FILLER_0_158 ();
 sg13g2_decap_8 FILLER_0_165 ();
 sg13g2_decap_8 FILLER_0_172 ();
 sg13g2_decap_8 FILLER_0_179 ();
 sg13g2_decap_8 FILLER_0_186 ();
 sg13g2_decap_8 FILLER_0_193 ();
 sg13g2_decap_8 FILLER_0_200 ();
 sg13g2_decap_8 FILLER_0_207 ();
 sg13g2_decap_8 FILLER_0_214 ();
 sg13g2_decap_8 FILLER_0_221 ();
 sg13g2_decap_8 FILLER_0_228 ();
 sg13g2_fill_2 FILLER_0_235 ();
 sg13g2_fill_1 FILLER_0_237 ();
 sg13g2_decap_8 FILLER_0_243 ();
 sg13g2_decap_8 FILLER_0_250 ();
 sg13g2_decap_8 FILLER_0_257 ();
 sg13g2_decap_8 FILLER_0_264 ();
 sg13g2_fill_2 FILLER_0_271 ();
 sg13g2_fill_2 FILLER_0_292 ();
 sg13g2_fill_1 FILLER_0_299 ();
 sg13g2_fill_1 FILLER_0_304 ();
 sg13g2_fill_1 FILLER_0_310 ();
 sg13g2_decap_8 FILLER_0_326 ();
 sg13g2_fill_2 FILLER_0_333 ();
 sg13g2_fill_1 FILLER_0_335 ();
 sg13g2_decap_8 FILLER_0_351 ();
 sg13g2_decap_4 FILLER_0_358 ();
 sg13g2_fill_2 FILLER_0_362 ();
 sg13g2_decap_8 FILLER_0_368 ();
 sg13g2_decap_8 FILLER_0_375 ();
 sg13g2_decap_8 FILLER_0_382 ();
 sg13g2_decap_8 FILLER_0_389 ();
 sg13g2_decap_8 FILLER_0_396 ();
 sg13g2_decap_4 FILLER_0_403 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_fill_2 FILLER_1_7 ();
 sg13g2_decap_4 FILLER_1_13 ();
 sg13g2_fill_2 FILLER_1_33 ();
 sg13g2_fill_1 FILLER_1_44 ();
 sg13g2_fill_1 FILLER_1_105 ();
 sg13g2_fill_1 FILLER_1_149 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_fill_2 FILLER_1_260 ();
 sg13g2_fill_2 FILLER_1_281 ();
 sg13g2_fill_1 FILLER_1_283 ();
 sg13g2_fill_1 FILLER_1_291 ();
 sg13g2_fill_2 FILLER_1_307 ();
 sg13g2_fill_1 FILLER_1_309 ();
 sg13g2_fill_2 FILLER_1_329 ();
 sg13g2_fill_1 FILLER_1_336 ();
 sg13g2_fill_2 FILLER_1_356 ();
 sg13g2_fill_2 FILLER_1_380 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_4 FILLER_2_0 ();
 sg13g2_fill_1 FILLER_2_4 ();
 sg13g2_fill_1 FILLER_2_44 ();
 sg13g2_fill_1 FILLER_2_70 ();
 sg13g2_fill_2 FILLER_2_81 ();
 sg13g2_fill_2 FILLER_2_114 ();
 sg13g2_fill_1 FILLER_2_116 ();
 sg13g2_fill_1 FILLER_2_130 ();
 sg13g2_decap_8 FILLER_2_173 ();
 sg13g2_decap_8 FILLER_2_180 ();
 sg13g2_decap_8 FILLER_2_187 ();
 sg13g2_decap_8 FILLER_2_194 ();
 sg13g2_decap_8 FILLER_2_201 ();
 sg13g2_decap_8 FILLER_2_208 ();
 sg13g2_decap_8 FILLER_2_215 ();
 sg13g2_decap_8 FILLER_2_222 ();
 sg13g2_decap_4 FILLER_2_229 ();
 sg13g2_fill_1 FILLER_2_233 ();
 sg13g2_fill_1 FILLER_2_248 ();
 sg13g2_decap_4 FILLER_2_262 ();
 sg13g2_decap_4 FILLER_2_294 ();
 sg13g2_fill_2 FILLER_2_303 ();
 sg13g2_fill_1 FILLER_2_305 ();
 sg13g2_decap_8 FILLER_2_326 ();
 sg13g2_fill_2 FILLER_2_333 ();
 sg13g2_fill_1 FILLER_2_335 ();
 sg13g2_fill_2 FILLER_2_341 ();
 sg13g2_fill_1 FILLER_2_343 ();
 sg13g2_fill_2 FILLER_2_366 ();
 sg13g2_fill_2 FILLER_2_392 ();
 sg13g2_decap_4 FILLER_2_404 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_fill_1 FILLER_3_71 ();
 sg13g2_fill_1 FILLER_3_82 ();
 sg13g2_fill_1 FILLER_3_111 ();
 sg13g2_fill_1 FILLER_3_138 ();
 sg13g2_fill_2 FILLER_3_153 ();
 sg13g2_fill_1 FILLER_3_155 ();
 sg13g2_decap_8 FILLER_3_191 ();
 sg13g2_decap_8 FILLER_3_198 ();
 sg13g2_decap_8 FILLER_3_205 ();
 sg13g2_decap_8 FILLER_3_212 ();
 sg13g2_decap_8 FILLER_3_219 ();
 sg13g2_decap_4 FILLER_3_226 ();
 sg13g2_fill_1 FILLER_3_230 ();
 sg13g2_fill_1 FILLER_3_242 ();
 sg13g2_decap_8 FILLER_3_249 ();
 sg13g2_decap_4 FILLER_3_256 ();
 sg13g2_fill_1 FILLER_3_260 ();
 sg13g2_fill_1 FILLER_3_275 ();
 sg13g2_fill_2 FILLER_3_285 ();
 sg13g2_fill_1 FILLER_3_315 ();
 sg13g2_fill_1 FILLER_3_329 ();
 sg13g2_fill_2 FILLER_3_338 ();
 sg13g2_fill_2 FILLER_3_351 ();
 sg13g2_fill_1 FILLER_3_353 ();
 sg13g2_fill_2 FILLER_3_387 ();
 sg13g2_fill_1 FILLER_3_389 ();
 sg13g2_decap_4 FILLER_3_405 ();
 sg13g2_fill_2 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_2 ();
 sg13g2_fill_2 FILLER_4_73 ();
 sg13g2_fill_2 FILLER_4_194 ();
 sg13g2_decap_8 FILLER_4_200 ();
 sg13g2_decap_4 FILLER_4_207 ();
 sg13g2_fill_1 FILLER_4_211 ();
 sg13g2_decap_8 FILLER_4_220 ();
 sg13g2_fill_2 FILLER_4_230 ();
 sg13g2_fill_2 FILLER_4_248 ();
 sg13g2_fill_2 FILLER_4_267 ();
 sg13g2_fill_2 FILLER_4_289 ();
 sg13g2_fill_1 FILLER_4_291 ();
 sg13g2_decap_8 FILLER_4_305 ();
 sg13g2_fill_2 FILLER_4_312 ();
 sg13g2_fill_2 FILLER_4_332 ();
 sg13g2_decap_8 FILLER_4_339 ();
 sg13g2_fill_1 FILLER_4_346 ();
 sg13g2_decap_4 FILLER_4_357 ();
 sg13g2_decap_4 FILLER_4_367 ();
 sg13g2_fill_1 FILLER_4_371 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_fill_2 FILLER_5_101 ();
 sg13g2_fill_2 FILLER_5_108 ();
 sg13g2_fill_2 FILLER_5_135 ();
 sg13g2_fill_1 FILLER_5_137 ();
 sg13g2_fill_1 FILLER_5_173 ();
 sg13g2_fill_2 FILLER_5_183 ();
 sg13g2_decap_4 FILLER_5_219 ();
 sg13g2_fill_2 FILLER_5_223 ();
 sg13g2_decap_4 FILLER_5_238 ();
 sg13g2_fill_1 FILLER_5_247 ();
 sg13g2_fill_2 FILLER_5_261 ();
 sg13g2_fill_1 FILLER_5_263 ();
 sg13g2_fill_2 FILLER_5_279 ();
 sg13g2_fill_2 FILLER_5_287 ();
 sg13g2_fill_1 FILLER_5_289 ();
 sg13g2_fill_1 FILLER_5_295 ();
 sg13g2_fill_2 FILLER_5_301 ();
 sg13g2_fill_1 FILLER_5_303 ();
 sg13g2_fill_2 FILLER_5_322 ();
 sg13g2_decap_4 FILLER_5_345 ();
 sg13g2_fill_2 FILLER_5_383 ();
 sg13g2_fill_2 FILLER_6_67 ();
 sg13g2_fill_2 FILLER_6_103 ();
 sg13g2_fill_1 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_125 ();
 sg13g2_fill_1 FILLER_6_132 ();
 sg13g2_fill_1 FILLER_6_137 ();
 sg13g2_fill_2 FILLER_6_150 ();
 sg13g2_fill_1 FILLER_6_152 ();
 sg13g2_fill_2 FILLER_6_184 ();
 sg13g2_decap_4 FILLER_6_198 ();
 sg13g2_fill_1 FILLER_6_237 ();
 sg13g2_fill_2 FILLER_6_280 ();
 sg13g2_fill_1 FILLER_6_310 ();
 sg13g2_fill_2 FILLER_6_337 ();
 sg13g2_fill_1 FILLER_6_339 ();
 sg13g2_fill_2 FILLER_6_355 ();
 sg13g2_fill_2 FILLER_6_373 ();
 sg13g2_fill_1 FILLER_6_375 ();
 sg13g2_fill_2 FILLER_6_380 ();
 sg13g2_decap_4 FILLER_6_386 ();
 sg13g2_decap_4 FILLER_6_404 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_fill_2 FILLER_7_26 ();
 sg13g2_fill_1 FILLER_7_108 ();
 sg13g2_fill_2 FILLER_7_156 ();
 sg13g2_fill_1 FILLER_7_158 ();
 sg13g2_fill_1 FILLER_7_211 ();
 sg13g2_fill_2 FILLER_7_229 ();
 sg13g2_fill_1 FILLER_7_239 ();
 sg13g2_decap_8 FILLER_7_248 ();
 sg13g2_decap_8 FILLER_7_263 ();
 sg13g2_decap_8 FILLER_7_279 ();
 sg13g2_decap_4 FILLER_7_286 ();
 sg13g2_fill_2 FILLER_7_299 ();
 sg13g2_fill_1 FILLER_7_301 ();
 sg13g2_fill_1 FILLER_7_311 ();
 sg13g2_fill_2 FILLER_7_322 ();
 sg13g2_fill_1 FILLER_7_324 ();
 sg13g2_fill_1 FILLER_7_334 ();
 sg13g2_fill_2 FILLER_7_348 ();
 sg13g2_decap_4 FILLER_7_358 ();
 sg13g2_fill_2 FILLER_7_362 ();
 sg13g2_fill_2 FILLER_7_378 ();
 sg13g2_fill_1 FILLER_7_380 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_fill_2 FILLER_8_26 ();
 sg13g2_fill_2 FILLER_8_66 ();
 sg13g2_fill_1 FILLER_8_103 ();
 sg13g2_decap_8 FILLER_8_130 ();
 sg13g2_decap_4 FILLER_8_137 ();
 sg13g2_fill_1 FILLER_8_141 ();
 sg13g2_fill_1 FILLER_8_155 ();
 sg13g2_fill_2 FILLER_8_186 ();
 sg13g2_fill_1 FILLER_8_188 ();
 sg13g2_decap_4 FILLER_8_194 ();
 sg13g2_fill_2 FILLER_8_198 ();
 sg13g2_fill_2 FILLER_8_208 ();
 sg13g2_decap_4 FILLER_8_240 ();
 sg13g2_fill_1 FILLER_8_244 ();
 sg13g2_decap_8 FILLER_8_253 ();
 sg13g2_fill_2 FILLER_8_302 ();
 sg13g2_fill_2 FILLER_8_314 ();
 sg13g2_fill_1 FILLER_8_329 ();
 sg13g2_fill_1 FILLER_8_338 ();
 sg13g2_decap_4 FILLER_8_355 ();
 sg13g2_fill_1 FILLER_8_359 ();
 sg13g2_fill_1 FILLER_8_370 ();
 sg13g2_fill_2 FILLER_8_376 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_97 ();
 sg13g2_decap_4 FILLER_9_138 ();
 sg13g2_decap_8 FILLER_9_188 ();
 sg13g2_fill_2 FILLER_9_216 ();
 sg13g2_fill_2 FILLER_9_223 ();
 sg13g2_decap_8 FILLER_9_241 ();
 sg13g2_decap_4 FILLER_9_261 ();
 sg13g2_fill_1 FILLER_9_265 ();
 sg13g2_fill_1 FILLER_9_283 ();
 sg13g2_fill_2 FILLER_9_306 ();
 sg13g2_fill_2 FILLER_9_345 ();
 sg13g2_decap_4 FILLER_9_353 ();
 sg13g2_fill_2 FILLER_9_372 ();
 sg13g2_fill_1 FILLER_9_374 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_fill_1 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_103 ();
 sg13g2_fill_1 FILLER_10_120 ();
 sg13g2_fill_1 FILLER_10_125 ();
 sg13g2_fill_2 FILLER_10_134 ();
 sg13g2_fill_2 FILLER_10_159 ();
 sg13g2_fill_2 FILLER_10_169 ();
 sg13g2_fill_1 FILLER_10_176 ();
 sg13g2_decap_4 FILLER_10_219 ();
 sg13g2_decap_4 FILLER_10_247 ();
 sg13g2_fill_2 FILLER_10_251 ();
 sg13g2_fill_2 FILLER_10_264 ();
 sg13g2_decap_4 FILLER_10_270 ();
 sg13g2_fill_1 FILLER_10_274 ();
 sg13g2_decap_8 FILLER_10_279 ();
 sg13g2_fill_2 FILLER_10_286 ();
 sg13g2_fill_2 FILLER_10_309 ();
 sg13g2_fill_1 FILLER_10_325 ();
 sg13g2_decap_4 FILLER_10_331 ();
 sg13g2_fill_1 FILLER_10_335 ();
 sg13g2_fill_1 FILLER_10_340 ();
 sg13g2_decap_4 FILLER_10_346 ();
 sg13g2_fill_2 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_363 ();
 sg13g2_fill_2 FILLER_10_370 ();
 sg13g2_fill_1 FILLER_10_372 ();
 sg13g2_fill_1 FILLER_10_387 ();
 sg13g2_decap_8 FILLER_10_394 ();
 sg13g2_decap_8 FILLER_10_401 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_fill_1 FILLER_11_52 ();
 sg13g2_fill_2 FILLER_11_77 ();
 sg13g2_fill_2 FILLER_11_88 ();
 sg13g2_fill_2 FILLER_11_125 ();
 sg13g2_fill_2 FILLER_11_157 ();
 sg13g2_fill_1 FILLER_11_164 ();
 sg13g2_fill_2 FILLER_11_174 ();
 sg13g2_fill_1 FILLER_11_181 ();
 sg13g2_fill_2 FILLER_11_196 ();
 sg13g2_fill_2 FILLER_11_203 ();
 sg13g2_fill_1 FILLER_11_205 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_fill_1 FILLER_11_223 ();
 sg13g2_decap_8 FILLER_11_229 ();
 sg13g2_fill_2 FILLER_11_240 ();
 sg13g2_fill_1 FILLER_11_247 ();
 sg13g2_fill_1 FILLER_11_258 ();
 sg13g2_fill_2 FILLER_11_268 ();
 sg13g2_fill_1 FILLER_11_270 ();
 sg13g2_decap_8 FILLER_11_288 ();
 sg13g2_decap_8 FILLER_11_295 ();
 sg13g2_decap_4 FILLER_11_302 ();
 sg13g2_fill_2 FILLER_11_322 ();
 sg13g2_fill_2 FILLER_11_344 ();
 sg13g2_fill_1 FILLER_11_346 ();
 sg13g2_fill_2 FILLER_11_361 ();
 sg13g2_fill_1 FILLER_11_363 ();
 sg13g2_fill_1 FILLER_11_370 ();
 sg13g2_decap_8 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_395 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_119 ();
 sg13g2_fill_1 FILLER_12_153 ();
 sg13g2_fill_2 FILLER_12_159 ();
 sg13g2_fill_1 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_188 ();
 sg13g2_fill_2 FILLER_12_216 ();
 sg13g2_fill_2 FILLER_12_247 ();
 sg13g2_fill_1 FILLER_12_264 ();
 sg13g2_decap_4 FILLER_12_298 ();
 sg13g2_fill_1 FILLER_12_302 ();
 sg13g2_fill_2 FILLER_12_363 ();
 sg13g2_decap_8 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_388 ();
 sg13g2_decap_8 FILLER_12_395 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_fill_1 FILLER_13_51 ();
 sg13g2_fill_1 FILLER_13_92 ();
 sg13g2_fill_1 FILLER_13_102 ();
 sg13g2_fill_1 FILLER_13_115 ();
 sg13g2_fill_2 FILLER_13_120 ();
 sg13g2_fill_1 FILLER_13_122 ();
 sg13g2_fill_2 FILLER_13_144 ();
 sg13g2_fill_2 FILLER_13_156 ();
 sg13g2_fill_1 FILLER_13_181 ();
 sg13g2_fill_2 FILLER_13_186 ();
 sg13g2_decap_4 FILLER_13_192 ();
 sg13g2_fill_1 FILLER_13_205 ();
 sg13g2_decap_4 FILLER_13_212 ();
 sg13g2_fill_2 FILLER_13_240 ();
 sg13g2_fill_1 FILLER_13_242 ();
 sg13g2_fill_2 FILLER_13_262 ();
 sg13g2_fill_1 FILLER_13_278 ();
 sg13g2_fill_2 FILLER_13_303 ();
 sg13g2_fill_1 FILLER_13_305 ();
 sg13g2_fill_2 FILLER_13_322 ();
 sg13g2_fill_1 FILLER_13_324 ();
 sg13g2_fill_2 FILLER_13_341 ();
 sg13g2_decap_8 FILLER_13_379 ();
 sg13g2_decap_8 FILLER_13_386 ();
 sg13g2_decap_8 FILLER_13_393 ();
 sg13g2_decap_8 FILLER_13_400 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_fill_1 FILLER_14_17 ();
 sg13g2_fill_2 FILLER_14_106 ();
 sg13g2_fill_2 FILLER_14_114 ();
 sg13g2_decap_8 FILLER_14_129 ();
 sg13g2_fill_1 FILLER_14_146 ();
 sg13g2_decap_4 FILLER_14_158 ();
 sg13g2_fill_2 FILLER_14_198 ();
 sg13g2_fill_1 FILLER_14_200 ();
 sg13g2_fill_2 FILLER_14_215 ();
 sg13g2_decap_4 FILLER_14_237 ();
 sg13g2_fill_1 FILLER_14_241 ();
 sg13g2_decap_4 FILLER_14_268 ();
 sg13g2_fill_2 FILLER_14_272 ();
 sg13g2_decap_4 FILLER_14_299 ();
 sg13g2_fill_1 FILLER_14_303 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_fill_2 FILLER_14_343 ();
 sg13g2_fill_1 FILLER_14_345 ();
 sg13g2_decap_4 FILLER_14_355 ();
 sg13g2_fill_2 FILLER_14_359 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_fill_1 FILLER_15_26 ();
 sg13g2_fill_1 FILLER_15_58 ();
 sg13g2_fill_2 FILLER_15_68 ();
 sg13g2_fill_2 FILLER_15_79 ();
 sg13g2_fill_1 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_128 ();
 sg13g2_fill_2 FILLER_15_135 ();
 sg13g2_fill_1 FILLER_15_137 ();
 sg13g2_fill_2 FILLER_15_148 ();
 sg13g2_decap_4 FILLER_15_165 ();
 sg13g2_fill_1 FILLER_15_169 ();
 sg13g2_fill_2 FILLER_15_189 ();
 sg13g2_fill_1 FILLER_15_191 ();
 sg13g2_decap_4 FILLER_15_209 ();
 sg13g2_fill_2 FILLER_15_213 ();
 sg13g2_fill_1 FILLER_15_225 ();
 sg13g2_fill_2 FILLER_15_239 ();
 sg13g2_fill_1 FILLER_15_241 ();
 sg13g2_fill_1 FILLER_15_278 ();
 sg13g2_decap_8 FILLER_15_290 ();
 sg13g2_decap_8 FILLER_15_297 ();
 sg13g2_fill_2 FILLER_15_304 ();
 sg13g2_fill_2 FILLER_15_310 ();
 sg13g2_decap_4 FILLER_15_316 ();
 sg13g2_fill_1 FILLER_15_320 ();
 sg13g2_decap_4 FILLER_15_359 ();
 sg13g2_fill_1 FILLER_15_363 ();
 sg13g2_fill_1 FILLER_15_373 ();
 sg13g2_decap_8 FILLER_15_382 ();
 sg13g2_fill_2 FILLER_15_389 ();
 sg13g2_fill_1 FILLER_15_391 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_fill_2 FILLER_16_17 ();
 sg13g2_fill_1 FILLER_16_19 ();
 sg13g2_fill_2 FILLER_16_138 ();
 sg13g2_fill_2 FILLER_16_206 ();
 sg13g2_fill_1 FILLER_16_208 ();
 sg13g2_fill_1 FILLER_16_222 ();
 sg13g2_decap_4 FILLER_16_233 ();
 sg13g2_decap_4 FILLER_16_242 ();
 sg13g2_fill_1 FILLER_16_251 ();
 sg13g2_fill_1 FILLER_16_257 ();
 sg13g2_decap_4 FILLER_16_263 ();
 sg13g2_fill_1 FILLER_16_273 ();
 sg13g2_decap_4 FILLER_16_289 ();
 sg13g2_fill_2 FILLER_16_293 ();
 sg13g2_decap_4 FILLER_16_326 ();
 sg13g2_fill_2 FILLER_16_330 ();
 sg13g2_fill_2 FILLER_16_336 ();
 sg13g2_fill_1 FILLER_16_338 ();
 sg13g2_decap_4 FILLER_16_344 ();
 sg13g2_fill_1 FILLER_16_382 ();
 sg13g2_fill_1 FILLER_17_26 ();
 sg13g2_fill_1 FILLER_17_53 ();
 sg13g2_fill_1 FILLER_17_124 ();
 sg13g2_fill_2 FILLER_17_131 ();
 sg13g2_fill_1 FILLER_17_133 ();
 sg13g2_fill_2 FILLER_17_145 ();
 sg13g2_fill_1 FILLER_17_150 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_fill_2 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_200 ();
 sg13g2_decap_4 FILLER_17_207 ();
 sg13g2_fill_1 FILLER_17_215 ();
 sg13g2_fill_1 FILLER_17_221 ();
 sg13g2_fill_1 FILLER_17_230 ();
 sg13g2_fill_2 FILLER_17_272 ();
 sg13g2_fill_1 FILLER_17_274 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_fill_2 FILLER_17_351 ();
 sg13g2_fill_1 FILLER_17_353 ();
 sg13g2_fill_1 FILLER_17_371 ();
 sg13g2_fill_2 FILLER_17_390 ();
 sg13g2_fill_2 FILLER_17_397 ();
 sg13g2_fill_1 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_18_34 ();
 sg13g2_fill_2 FILLER_18_107 ();
 sg13g2_fill_2 FILLER_18_125 ();
 sg13g2_fill_2 FILLER_18_152 ();
 sg13g2_decap_4 FILLER_18_159 ();
 sg13g2_fill_1 FILLER_18_163 ();
 sg13g2_fill_2 FILLER_18_169 ();
 sg13g2_fill_1 FILLER_18_184 ();
 sg13g2_fill_1 FILLER_18_215 ();
 sg13g2_fill_1 FILLER_18_230 ();
 sg13g2_fill_2 FILLER_18_264 ();
 sg13g2_fill_1 FILLER_18_287 ();
 sg13g2_fill_2 FILLER_18_314 ();
 sg13g2_fill_2 FILLER_18_333 ();
 sg13g2_fill_1 FILLER_18_345 ();
 sg13g2_fill_2 FILLER_19_35 ();
 sg13g2_fill_1 FILLER_19_108 ();
 sg13g2_fill_1 FILLER_19_116 ();
 sg13g2_fill_2 FILLER_19_166 ();
 sg13g2_fill_1 FILLER_19_168 ();
 sg13g2_decap_4 FILLER_19_198 ();
 sg13g2_fill_2 FILLER_19_207 ();
 sg13g2_fill_2 FILLER_19_213 ();
 sg13g2_fill_1 FILLER_19_245 ();
 sg13g2_fill_1 FILLER_19_251 ();
 sg13g2_decap_8 FILLER_19_264 ();
 sg13g2_fill_1 FILLER_19_271 ();
 sg13g2_decap_4 FILLER_19_280 ();
 sg13g2_fill_2 FILLER_19_284 ();
 sg13g2_fill_2 FILLER_19_311 ();
 sg13g2_fill_1 FILLER_19_313 ();
 sg13g2_fill_2 FILLER_19_320 ();
 sg13g2_fill_1 FILLER_19_328 ();
 sg13g2_fill_1 FILLER_19_340 ();
 sg13g2_fill_1 FILLER_19_381 ();
 sg13g2_decap_4 FILLER_19_386 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_97 ();
 sg13g2_decap_8 FILLER_20_104 ();
 sg13g2_fill_1 FILLER_20_116 ();
 sg13g2_decap_8 FILLER_20_122 ();
 sg13g2_decap_8 FILLER_20_129 ();
 sg13g2_fill_2 FILLER_20_147 ();
 sg13g2_decap_4 FILLER_20_157 ();
 sg13g2_fill_2 FILLER_20_173 ();
 sg13g2_fill_1 FILLER_20_175 ();
 sg13g2_fill_1 FILLER_20_181 ();
 sg13g2_fill_2 FILLER_20_220 ();
 sg13g2_fill_2 FILLER_20_245 ();
 sg13g2_fill_2 FILLER_20_269 ();
 sg13g2_fill_2 FILLER_20_310 ();
 sg13g2_fill_2 FILLER_20_330 ();
 sg13g2_fill_1 FILLER_20_332 ();
 sg13g2_fill_1 FILLER_20_346 ();
 sg13g2_fill_1 FILLER_20_377 ();
 sg13g2_fill_2 FILLER_21_59 ();
 sg13g2_fill_2 FILLER_21_90 ();
 sg13g2_decap_4 FILLER_21_129 ();
 sg13g2_fill_2 FILLER_21_133 ();
 sg13g2_fill_2 FILLER_21_139 ();
 sg13g2_fill_1 FILLER_21_154 ();
 sg13g2_fill_2 FILLER_21_180 ();
 sg13g2_decap_4 FILLER_21_211 ();
 sg13g2_decap_8 FILLER_21_219 ();
 sg13g2_fill_1 FILLER_21_226 ();
 sg13g2_fill_2 FILLER_21_231 ();
 sg13g2_fill_1 FILLER_21_259 ();
 sg13g2_fill_1 FILLER_21_272 ();
 sg13g2_fill_2 FILLER_21_278 ();
 sg13g2_fill_2 FILLER_21_296 ();
 sg13g2_fill_1 FILLER_21_308 ();
 sg13g2_fill_2 FILLER_21_331 ();
 sg13g2_fill_1 FILLER_21_333 ();
 sg13g2_fill_2 FILLER_21_344 ();
 sg13g2_fill_1 FILLER_21_346 ();
 sg13g2_fill_2 FILLER_22_13 ();
 sg13g2_fill_1 FILLER_22_50 ();
 sg13g2_fill_2 FILLER_22_69 ();
 sg13g2_fill_1 FILLER_22_117 ();
 sg13g2_fill_1 FILLER_22_130 ();
 sg13g2_decap_4 FILLER_22_149 ();
 sg13g2_fill_1 FILLER_22_153 ();
 sg13g2_fill_2 FILLER_22_275 ();
 sg13g2_fill_1 FILLER_22_277 ();
 sg13g2_fill_2 FILLER_22_291 ();
 sg13g2_fill_1 FILLER_22_312 ();
 sg13g2_fill_2 FILLER_22_326 ();
 sg13g2_fill_2 FILLER_22_353 ();
 sg13g2_fill_1 FILLER_22_355 ();
 sg13g2_fill_2 FILLER_22_380 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_61 ();
 sg13g2_fill_2 FILLER_23_106 ();
 sg13g2_fill_2 FILLER_23_132 ();
 sg13g2_fill_1 FILLER_23_134 ();
 sg13g2_decap_4 FILLER_23_139 ();
 sg13g2_fill_1 FILLER_23_143 ();
 sg13g2_decap_4 FILLER_23_160 ();
 sg13g2_fill_2 FILLER_23_164 ();
 sg13g2_fill_2 FILLER_23_176 ();
 sg13g2_fill_1 FILLER_23_178 ();
 sg13g2_fill_2 FILLER_23_219 ();
 sg13g2_fill_2 FILLER_23_226 ();
 sg13g2_fill_1 FILLER_23_228 ();
 sg13g2_decap_8 FILLER_23_255 ();
 sg13g2_fill_1 FILLER_23_262 ();
 sg13g2_fill_2 FILLER_23_276 ();
 sg13g2_fill_1 FILLER_23_282 ();
 sg13g2_decap_4 FILLER_23_295 ();
 sg13g2_fill_2 FILLER_23_299 ();
 sg13g2_fill_2 FILLER_23_306 ();
 sg13g2_fill_2 FILLER_23_326 ();
 sg13g2_fill_2 FILLER_23_357 ();
 sg13g2_fill_1 FILLER_23_371 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_46 ();
 sg13g2_fill_2 FILLER_24_73 ();
 sg13g2_fill_1 FILLER_24_107 ();
 sg13g2_fill_1 FILLER_24_133 ();
 sg13g2_decap_4 FILLER_24_150 ();
 sg13g2_fill_1 FILLER_24_162 ();
 sg13g2_fill_1 FILLER_24_179 ();
 sg13g2_fill_2 FILLER_24_198 ();
 sg13g2_fill_1 FILLER_24_200 ();
 sg13g2_fill_1 FILLER_24_210 ();
 sg13g2_fill_2 FILLER_24_232 ();
 sg13g2_fill_1 FILLER_24_234 ();
 sg13g2_decap_4 FILLER_24_282 ();
 sg13g2_fill_2 FILLER_24_286 ();
 sg13g2_decap_8 FILLER_24_298 ();
 sg13g2_decap_4 FILLER_24_305 ();
 sg13g2_decap_4 FILLER_24_322 ();
 sg13g2_fill_1 FILLER_24_326 ();
 sg13g2_decap_8 FILLER_24_339 ();
 sg13g2_fill_1 FILLER_24_346 ();
 sg13g2_decap_4 FILLER_24_359 ();
 sg13g2_fill_2 FILLER_24_363 ();
 sg13g2_fill_1 FILLER_25_44 ();
 sg13g2_fill_2 FILLER_25_84 ();
 sg13g2_fill_1 FILLER_25_86 ();
 sg13g2_fill_2 FILLER_25_95 ();
 sg13g2_fill_1 FILLER_25_97 ();
 sg13g2_fill_1 FILLER_25_110 ();
 sg13g2_decap_4 FILLER_25_115 ();
 sg13g2_fill_2 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_125 ();
 sg13g2_decap_8 FILLER_25_142 ();
 sg13g2_decap_8 FILLER_25_149 ();
 sg13g2_decap_4 FILLER_25_156 ();
 sg13g2_fill_1 FILLER_25_160 ();
 sg13g2_decap_8 FILLER_25_177 ();
 sg13g2_fill_2 FILLER_25_184 ();
 sg13g2_fill_2 FILLER_25_216 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_fill_2 FILLER_25_305 ();
 sg13g2_decap_8 FILLER_25_327 ();
 sg13g2_decap_4 FILLER_25_334 ();
 sg13g2_fill_1 FILLER_25_338 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_fill_2 FILLER_26_19 ();
 sg13g2_fill_2 FILLER_26_74 ();
 sg13g2_fill_1 FILLER_26_76 ();
 sg13g2_fill_1 FILLER_26_88 ();
 sg13g2_decap_4 FILLER_26_132 ();
 sg13g2_fill_1 FILLER_26_160 ();
 sg13g2_decap_4 FILLER_26_185 ();
 sg13g2_fill_1 FILLER_26_189 ();
 sg13g2_fill_2 FILLER_26_198 ();
 sg13g2_fill_2 FILLER_26_233 ();
 sg13g2_decap_8 FILLER_26_260 ();
 sg13g2_fill_1 FILLER_26_267 ();
 sg13g2_decap_4 FILLER_26_284 ();
 sg13g2_fill_1 FILLER_26_288 ();
 sg13g2_decap_4 FILLER_26_302 ();
 sg13g2_decap_8 FILLER_26_323 ();
 sg13g2_decap_8 FILLER_26_330 ();
 sg13g2_decap_8 FILLER_26_337 ();
 sg13g2_decap_4 FILLER_26_353 ();
 sg13g2_decap_8 FILLER_26_379 ();
 sg13g2_decap_8 FILLER_26_395 ();
 sg13g2_decap_8 FILLER_26_402 ();
 sg13g2_fill_1 FILLER_27_25 ();
 sg13g2_fill_2 FILLER_27_36 ();
 sg13g2_fill_1 FILLER_27_38 ();
 sg13g2_fill_2 FILLER_27_45 ();
 sg13g2_fill_1 FILLER_27_57 ();
 sg13g2_fill_2 FILLER_27_65 ();
 sg13g2_fill_2 FILLER_27_84 ();
 sg13g2_fill_2 FILLER_27_92 ();
 sg13g2_fill_1 FILLER_27_94 ();
 sg13g2_fill_1 FILLER_27_105 ();
 sg13g2_fill_1 FILLER_27_110 ();
 sg13g2_fill_2 FILLER_27_117 ();
 sg13g2_decap_4 FILLER_27_134 ();
 sg13g2_decap_4 FILLER_27_150 ();
 sg13g2_decap_4 FILLER_27_166 ();
 sg13g2_fill_1 FILLER_27_170 ();
 sg13g2_decap_4 FILLER_27_188 ();
 sg13g2_fill_1 FILLER_27_219 ();
 sg13g2_fill_2 FILLER_27_235 ();
 sg13g2_fill_1 FILLER_27_237 ();
 sg13g2_fill_1 FILLER_27_244 ();
 sg13g2_fill_2 FILLER_27_253 ();
 sg13g2_fill_2 FILLER_27_260 ();
 sg13g2_fill_1 FILLER_27_262 ();
 sg13g2_fill_2 FILLER_27_279 ();
 sg13g2_decap_4 FILLER_27_305 ();
 sg13g2_decap_4 FILLER_27_317 ();
 sg13g2_fill_2 FILLER_27_333 ();
 sg13g2_fill_2 FILLER_27_356 ();
 sg13g2_fill_1 FILLER_27_358 ();
 sg13g2_fill_2 FILLER_27_381 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_45 ();
 sg13g2_fill_1 FILLER_28_52 ();
 sg13g2_fill_2 FILLER_28_82 ();
 sg13g2_fill_1 FILLER_28_84 ();
 sg13g2_fill_2 FILLER_28_95 ();
 sg13g2_decap_8 FILLER_28_121 ();
 sg13g2_decap_8 FILLER_28_128 ();
 sg13g2_decap_4 FILLER_28_135 ();
 sg13g2_decap_8 FILLER_28_151 ();
 sg13g2_fill_2 FILLER_28_212 ();
 sg13g2_fill_1 FILLER_28_214 ();
 sg13g2_fill_1 FILLER_28_223 ();
 sg13g2_fill_2 FILLER_28_271 ();
 sg13g2_fill_2 FILLER_28_312 ();
 sg13g2_fill_1 FILLER_28_314 ();
 sg13g2_fill_2 FILLER_28_340 ();
 sg13g2_fill_1 FILLER_28_356 ();
 sg13g2_decap_4 FILLER_28_361 ();
 sg13g2_fill_1 FILLER_28_365 ();
 sg13g2_decap_4 FILLER_28_380 ();
 sg13g2_fill_1 FILLER_28_384 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_24 ();
 sg13g2_fill_2 FILLER_29_45 ();
 sg13g2_fill_2 FILLER_29_52 ();
 sg13g2_fill_2 FILLER_29_60 ();
 sg13g2_fill_1 FILLER_29_62 ();
 sg13g2_decap_8 FILLER_29_129 ();
 sg13g2_fill_2 FILLER_29_136 ();
 sg13g2_fill_2 FILLER_29_150 ();
 sg13g2_fill_1 FILLER_29_205 ();
 sg13g2_decap_8 FILLER_29_257 ();
 sg13g2_fill_1 FILLER_29_300 ();
 sg13g2_fill_1 FILLER_29_316 ();
 sg13g2_fill_2 FILLER_29_332 ();
 sg13g2_fill_2 FILLER_29_391 ();
 sg13g2_fill_1 FILLER_29_393 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_26 ();
 sg13g2_fill_1 FILLER_30_28 ();
 sg13g2_fill_1 FILLER_30_52 ();
 sg13g2_fill_1 FILLER_30_67 ();
 sg13g2_fill_1 FILLER_30_80 ();
 sg13g2_fill_1 FILLER_30_90 ();
 sg13g2_fill_2 FILLER_30_101 ();
 sg13g2_fill_2 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_151 ();
 sg13g2_decap_8 FILLER_30_158 ();
 sg13g2_fill_1 FILLER_30_177 ();
 sg13g2_fill_2 FILLER_30_221 ();
 sg13g2_fill_2 FILLER_30_227 ();
 sg13g2_fill_1 FILLER_30_229 ();
 sg13g2_fill_1 FILLER_30_259 ();
 sg13g2_fill_2 FILLER_30_272 ();
 sg13g2_fill_1 FILLER_30_274 ();
 sg13g2_decap_8 FILLER_30_284 ();
 sg13g2_fill_2 FILLER_30_291 ();
 sg13g2_decap_4 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_335 ();
 sg13g2_decap_4 FILLER_30_358 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_fill_2 FILLER_30_388 ();
 sg13g2_fill_1 FILLER_30_390 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_15 ();
 sg13g2_decap_4 FILLER_31_45 ();
 sg13g2_fill_1 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_87 ();
 sg13g2_fill_1 FILLER_31_115 ();
 sg13g2_fill_2 FILLER_31_128 ();
 sg13g2_fill_1 FILLER_31_130 ();
 sg13g2_fill_2 FILLER_31_152 ();
 sg13g2_decap_8 FILLER_31_183 ();
 sg13g2_decap_4 FILLER_31_190 ();
 sg13g2_fill_2 FILLER_31_194 ();
 sg13g2_fill_1 FILLER_31_204 ();
 sg13g2_fill_2 FILLER_31_257 ();
 sg13g2_fill_1 FILLER_31_259 ();
 sg13g2_fill_2 FILLER_31_283 ();
 sg13g2_fill_2 FILLER_31_304 ();
 sg13g2_decap_4 FILLER_31_325 ();
 sg13g2_fill_2 FILLER_31_329 ();
 sg13g2_fill_1 FILLER_31_355 ();
 sg13g2_decap_4 FILLER_31_375 ();
 sg13g2_fill_1 FILLER_31_379 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_50 ();
 sg13g2_fill_1 FILLER_32_52 ();
 sg13g2_fill_2 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_80 ();
 sg13g2_decap_8 FILLER_32_87 ();
 sg13g2_fill_2 FILLER_32_94 ();
 sg13g2_decap_4 FILLER_32_107 ();
 sg13g2_fill_2 FILLER_32_111 ();
 sg13g2_fill_1 FILLER_32_119 ();
 sg13g2_fill_1 FILLER_32_126 ();
 sg13g2_decap_4 FILLER_32_137 ();
 sg13g2_fill_1 FILLER_32_185 ();
 sg13g2_fill_2 FILLER_32_199 ();
 sg13g2_fill_1 FILLER_32_215 ();
 sg13g2_fill_2 FILLER_32_234 ();
 sg13g2_fill_1 FILLER_32_236 ();
 sg13g2_fill_1 FILLER_32_241 ();
 sg13g2_fill_2 FILLER_32_268 ();
 sg13g2_fill_2 FILLER_32_293 ();
 sg13g2_fill_1 FILLER_32_295 ();
 sg13g2_decap_4 FILLER_32_307 ();
 sg13g2_fill_1 FILLER_32_354 ();
 sg13g2_decap_4 FILLER_32_361 ();
 sg13g2_fill_1 FILLER_32_365 ();
 sg13g2_fill_1 FILLER_32_371 ();
 sg13g2_fill_1 FILLER_32_392 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_2 ();
 sg13g2_fill_2 FILLER_33_27 ();
 sg13g2_fill_1 FILLER_33_29 ();
 sg13g2_fill_1 FILLER_33_34 ();
 sg13g2_decap_4 FILLER_33_80 ();
 sg13g2_fill_2 FILLER_33_84 ();
 sg13g2_decap_4 FILLER_33_100 ();
 sg13g2_fill_1 FILLER_33_119 ();
 sg13g2_fill_2 FILLER_33_147 ();
 sg13g2_decap_4 FILLER_33_164 ();
 sg13g2_fill_2 FILLER_33_176 ();
 sg13g2_fill_1 FILLER_33_198 ();
 sg13g2_fill_1 FILLER_33_237 ();
 sg13g2_fill_1 FILLER_33_264 ();
 sg13g2_fill_1 FILLER_33_284 ();
 sg13g2_fill_2 FILLER_33_299 ();
 sg13g2_fill_1 FILLER_33_301 ();
 sg13g2_decap_4 FILLER_33_307 ();
 sg13g2_fill_1 FILLER_33_311 ();
 sg13g2_fill_2 FILLER_33_330 ();
 sg13g2_fill_1 FILLER_33_332 ();
 sg13g2_decap_4 FILLER_33_337 ();
 sg13g2_fill_1 FILLER_33_341 ();
 sg13g2_fill_2 FILLER_33_352 ();
 sg13g2_fill_1 FILLER_33_354 ();
 sg13g2_fill_2 FILLER_33_361 ();
 sg13g2_decap_8 FILLER_33_387 ();
 sg13g2_decap_4 FILLER_33_404 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_fill_2 FILLER_34_19 ();
 sg13g2_fill_1 FILLER_34_46 ();
 sg13g2_fill_1 FILLER_34_56 ();
 sg13g2_fill_2 FILLER_34_75 ();
 sg13g2_fill_1 FILLER_34_88 ();
 sg13g2_fill_2 FILLER_34_109 ();
 sg13g2_fill_1 FILLER_34_111 ();
 sg13g2_decap_8 FILLER_34_117 ();
 sg13g2_decap_4 FILLER_34_124 ();
 sg13g2_fill_2 FILLER_34_128 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_4 FILLER_34_147 ();
 sg13g2_fill_2 FILLER_34_164 ();
 sg13g2_fill_1 FILLER_34_166 ();
 sg13g2_decap_8 FILLER_34_172 ();
 sg13g2_fill_2 FILLER_34_179 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_fill_1 FILLER_34_237 ();
 sg13g2_fill_2 FILLER_34_244 ();
 sg13g2_decap_4 FILLER_34_263 ();
 sg13g2_decap_8 FILLER_34_282 ();
 sg13g2_decap_4 FILLER_34_330 ();
 sg13g2_fill_1 FILLER_34_334 ();
 sg13g2_decap_4 FILLER_34_359 ();
 sg13g2_fill_1 FILLER_34_363 ();
 sg13g2_decap_4 FILLER_34_380 ();
 sg13g2_fill_2 FILLER_34_384 ();
 sg13g2_fill_2 FILLER_34_392 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_fill_2 FILLER_35_23 ();
 sg13g2_fill_1 FILLER_35_25 ();
 sg13g2_fill_1 FILLER_35_44 ();
 sg13g2_fill_1 FILLER_35_105 ();
 sg13g2_fill_2 FILLER_35_124 ();
 sg13g2_fill_1 FILLER_35_143 ();
 sg13g2_fill_2 FILLER_35_174 ();
 sg13g2_fill_1 FILLER_35_176 ();
 sg13g2_fill_1 FILLER_35_193 ();
 sg13g2_fill_2 FILLER_35_220 ();
 sg13g2_decap_4 FILLER_35_232 ();
 sg13g2_fill_2 FILLER_35_248 ();
 sg13g2_fill_1 FILLER_35_250 ();
 sg13g2_decap_8 FILLER_35_262 ();
 sg13g2_fill_1 FILLER_35_269 ();
 sg13g2_fill_1 FILLER_35_291 ();
 sg13g2_fill_2 FILLER_35_360 ();
 sg13g2_fill_1 FILLER_35_362 ();
 sg13g2_fill_2 FILLER_35_388 ();
 sg13g2_fill_1 FILLER_35_390 ();
 sg13g2_fill_1 FILLER_36_31 ();
 sg13g2_fill_1 FILLER_36_92 ();
 sg13g2_fill_1 FILLER_36_114 ();
 sg13g2_fill_2 FILLER_36_120 ();
 sg13g2_decap_8 FILLER_36_142 ();
 sg13g2_fill_2 FILLER_36_149 ();
 sg13g2_fill_1 FILLER_36_151 ();
 sg13g2_decap_8 FILLER_36_170 ();
 sg13g2_fill_2 FILLER_36_196 ();
 sg13g2_fill_1 FILLER_36_198 ();
 sg13g2_fill_2 FILLER_36_206 ();
 sg13g2_decap_8 FILLER_36_220 ();
 sg13g2_decap_4 FILLER_36_227 ();
 sg13g2_fill_2 FILLER_36_231 ();
 sg13g2_decap_4 FILLER_36_259 ();
 sg13g2_fill_2 FILLER_36_263 ();
 sg13g2_fill_1 FILLER_36_289 ();
 sg13g2_fill_1 FILLER_36_316 ();
 sg13g2_decap_4 FILLER_36_327 ();
 sg13g2_fill_2 FILLER_36_331 ();
 sg13g2_decap_8 FILLER_36_353 ();
 sg13g2_fill_2 FILLER_36_367 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_14 ();
 sg13g2_fill_1 FILLER_37_76 ();
 sg13g2_fill_2 FILLER_37_106 ();
 sg13g2_decap_8 FILLER_37_130 ();
 sg13g2_fill_1 FILLER_37_137 ();
 sg13g2_decap_8 FILLER_37_146 ();
 sg13g2_decap_8 FILLER_37_153 ();
 sg13g2_decap_8 FILLER_37_160 ();
 sg13g2_decap_4 FILLER_37_167 ();
 sg13g2_fill_2 FILLER_37_171 ();
 sg13g2_decap_4 FILLER_37_199 ();
 sg13g2_fill_1 FILLER_37_222 ();
 sg13g2_decap_4 FILLER_37_264 ();
 sg13g2_fill_1 FILLER_37_288 ();
 sg13g2_fill_2 FILLER_37_307 ();
 sg13g2_fill_1 FILLER_37_345 ();
 sg13g2_fill_2 FILLER_37_393 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_4 ();
 sg13g2_fill_1 FILLER_38_34 ();
 sg13g2_fill_2 FILLER_38_70 ();
 sg13g2_fill_2 FILLER_38_94 ();
 sg13g2_fill_1 FILLER_38_113 ();
 sg13g2_fill_1 FILLER_38_122 ();
 sg13g2_fill_1 FILLER_38_135 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_8 FILLER_38_193 ();
 sg13g2_decap_4 FILLER_38_200 ();
 sg13g2_fill_1 FILLER_38_204 ();
 sg13g2_fill_1 FILLER_38_212 ();
 sg13g2_decap_8 FILLER_38_220 ();
 sg13g2_decap_4 FILLER_38_227 ();
 sg13g2_fill_2 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_260 ();
 sg13g2_decap_4 FILLER_38_267 ();
 sg13g2_fill_2 FILLER_38_276 ();
 sg13g2_fill_1 FILLER_38_278 ();
 sg13g2_decap_8 FILLER_38_283 ();
 sg13g2_fill_2 FILLER_38_290 ();
 sg13g2_fill_1 FILLER_38_292 ();
 sg13g2_decap_8 FILLER_38_303 ();
 sg13g2_fill_2 FILLER_38_310 ();
 sg13g2_fill_2 FILLER_38_334 ();
 sg13g2_fill_2 FILLER_38_354 ();
 sg13g2_fill_1 FILLER_38_381 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net8;
 assign uio_oe[1] = net9;
 assign uio_oe[2] = net10;
 assign uio_oe[3] = net11;
 assign uio_oe[4] = net12;
 assign uio_oe[5] = net13;
 assign uio_oe[6] = net14;
 assign uio_oe[7] = net44;
 assign uio_out[0] = net15;
 assign uio_out[1] = net16;
 assign uio_out[2] = net17;
 assign uio_out[3] = net18;
 assign uio_out[4] = net19;
 assign uio_out[5] = net20;
 assign uio_out[6] = net21;
endmodule

module tt_um_rebeccargb_universal_decoder (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire _463_;
 wire _464_;
 wire _465_;
 wire _466_;
 wire _467_;
 wire _468_;
 wire _469_;
 wire _470_;
 wire _471_;
 wire _472_;
 wire _473_;
 wire _474_;
 wire _475_;
 wire _476_;
 wire _477_;
 wire _478_;
 wire _479_;
 wire _480_;
 wire _481_;
 wire _482_;
 wire _483_;
 wire _484_;
 wire _485_;
 wire _486_;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 sg13g2_inv_1 _487_ (.Y(_169_),
    .A(net298));
 sg13g2_inv_2 _488_ (.Y(_180_),
    .A(net317));
 sg13g2_inv_1 _489_ (.Y(_191_),
    .A(net319));
 sg13g2_inv_1 _490_ (.Y(_202_),
    .A(net297));
 sg13g2_inv_2 _491_ (.Y(_213_),
    .A(net6));
 sg13g2_inv_2 _492_ (.Y(_224_),
    .A(net309));
 sg13g2_inv_2 _493_ (.Y(_234_),
    .A(net292));
 sg13g2_inv_1 _494_ (.Y(_245_),
    .A(net289));
 sg13g2_nor2b_1 _495_ (.A(net298),
    .B_N(net297),
    .Y(_256_));
 sg13g2_nor2_2 _496_ (.A(net322),
    .B(net326),
    .Y(_267_));
 sg13g2_or2_1 _497_ (.X(_277_),
    .B(net325),
    .A(net324));
 sg13g2_nor2_2 _498_ (.A(net315),
    .B(net1),
    .Y(_288_));
 sg13g2_or2_1 _499_ (.X(_299_),
    .B(net319),
    .A(net315));
 sg13g2_nor2_2 _500_ (.A(net281),
    .B(net279),
    .Y(_310_));
 sg13g2_nand2_1 _501_ (.Y(_320_),
    .A(_256_),
    .B(_310_));
 sg13g2_o21ai_1 _502_ (.B1(net291),
    .Y(_331_),
    .A1(net309),
    .A2(_320_));
 sg13g2_nor2_1 _503_ (.A(_213_),
    .B(_331_),
    .Y(_342_));
 sg13g2_nand2b_1 _504_ (.Y(_353_),
    .B(net302),
    .A_N(net304));
 sg13g2_and2_1 _505_ (.A(net298),
    .B(net297),
    .X(_363_));
 sg13g2_nand2_2 _506_ (.Y(_374_),
    .A(net300),
    .B(net295));
 sg13g2_and2_2 _507_ (.A(net303),
    .B(net309),
    .X(_385_));
 sg13g2_nand2_1 _508_ (.Y(_396_),
    .A(net303),
    .B(net311));
 sg13g2_a21oi_1 _509_ (.A1(net302),
    .A2(net310),
    .Y(_406_),
    .B1(net304));
 sg13g2_a22oi_1 _510_ (.Y(_417_),
    .B1(_363_),
    .B2(_406_),
    .A2(_353_),
    .A1(_256_));
 sg13g2_nand2_1 _511_ (.Y(_428_),
    .A(net6),
    .B(_417_));
 sg13g2_o21ai_1 _512_ (.B1(_234_),
    .Y(_437_),
    .A1(net293),
    .A2(_428_));
 sg13g2_a21oi_1 _513_ (.A1(net293),
    .A2(_428_),
    .Y(_441_),
    .B1(_437_));
 sg13g2_o21ai_1 _514_ (.B1(net290),
    .Y(_442_),
    .A1(_342_),
    .A2(_441_));
 sg13g2_a21oi_1 _515_ (.A1(net6),
    .A2(_320_),
    .Y(_443_),
    .B1(net291));
 sg13g2_nor2_1 _516_ (.A(_180_),
    .B(net284),
    .Y(_444_));
 sg13g2_and2_2 _517_ (.A(net322),
    .B(net326),
    .X(_445_));
 sg13g2_nand2_1 _518_ (.Y(_446_),
    .A(net324),
    .B(net325));
 sg13g2_o21ai_1 _519_ (.B1(_444_),
    .Y(_447_),
    .A1(net318),
    .A2(_445_));
 sg13g2_nand2_1 _520_ (.Y(_448_),
    .A(_224_),
    .B(_310_));
 sg13g2_nand4_1 _521_ (.B(net292),
    .C(_447_),
    .A(net2),
    .Y(_449_),
    .D(_448_));
 sg13g2_nand2b_1 _522_ (.Y(_450_),
    .B(_449_),
    .A_N(_443_));
 sg13g2_o21ai_1 _523_ (.B1(_442_),
    .Y(uo_out[7]),
    .A1(net290),
    .A2(_450_));
 sg13g2_nand2_2 _524_ (.Y(_451_),
    .A(net303),
    .B(net306));
 sg13g2_nand2b_1 _525_ (.Y(_452_),
    .B(net303),
    .A_N(net314));
 sg13g2_inv_1 _526_ (.Y(_453_),
    .A(net275));
 sg13g2_nor2_2 _527_ (.A(net309),
    .B(_451_),
    .Y(_454_));
 sg13g2_nand3b_1 _528_ (.B(net307),
    .C(net2),
    .Y(_455_),
    .A_N(net311));
 sg13g2_nand2b_2 _529_ (.Y(_456_),
    .B(net325),
    .A_N(net317));
 sg13g2_nor2b_2 _530_ (.A(net316),
    .B_N(net318),
    .Y(_457_));
 sg13g2_nand2b_1 _531_ (.Y(_458_),
    .B(net319),
    .A_N(net315));
 sg13g2_nand2b_1 _532_ (.Y(_459_),
    .B(net325),
    .A_N(net324));
 sg13g2_nor2_2 _533_ (.A(net270),
    .B(net267),
    .Y(_460_));
 sg13g2_nor3_2 _534_ (.A(net272),
    .B(net269),
    .C(net267),
    .Y(_461_));
 sg13g2_nor2b_2 _535_ (.A(net325),
    .B_N(net323),
    .Y(_462_));
 sg13g2_nand2b_1 _536_ (.Y(_463_),
    .B(net323),
    .A_N(net326));
 sg13g2_nand2_1 _537_ (.Y(_464_),
    .A(net322),
    .B(_457_));
 sg13g2_nor2_2 _538_ (.A(net271),
    .B(net266),
    .Y(_465_));
 sg13g2_nand2_1 _539_ (.Y(_466_),
    .A(_457_),
    .B(_462_));
 sg13g2_nor2_2 _540_ (.A(net284),
    .B(_451_),
    .Y(_467_));
 sg13g2_nand3_1 _541_ (.B(net311),
    .C(net307),
    .A(net2),
    .Y(_468_));
 sg13g2_nor3_1 _542_ (.A(net269),
    .B(net263),
    .C(_468_),
    .Y(_469_));
 sg13g2_a22oi_1 _543_ (.Y(_470_),
    .B1(_469_),
    .B2(net287),
    .A2(_461_),
    .A1(_374_));
 sg13g2_nor2_1 _544_ (.A(net307),
    .B(_396_),
    .Y(_471_));
 sg13g2_nor2b_2 _545_ (.A(net318),
    .B_N(net316),
    .Y(_472_));
 sg13g2_nand2b_1 _546_ (.Y(_473_),
    .B(net315),
    .A_N(net1));
 sg13g2_nor2_1 _547_ (.A(net322),
    .B(net318),
    .Y(_474_));
 sg13g2_nor2_2 _548_ (.A(net322),
    .B(net262),
    .Y(_475_));
 sg13g2_nand2_1 _549_ (.Y(_476_),
    .A(_267_),
    .B(_472_));
 sg13g2_a22oi_1 _550_ (.Y(_477_),
    .B1(_472_),
    .B2(_267_),
    .A2(_462_),
    .A1(_457_));
 sg13g2_nand2b_1 _551_ (.Y(_478_),
    .B(net251),
    .A_N(_477_));
 sg13g2_nand2b_1 _552_ (.Y(_479_),
    .B(net308),
    .A_N(net303));
 sg13g2_nor2_1 _553_ (.A(_224_),
    .B(net258),
    .Y(_480_));
 sg13g2_nand3b_1 _554_ (.B(net313),
    .C(net308),
    .Y(_481_),
    .A_N(net303));
 sg13g2_nor2_1 _555_ (.A(net321),
    .B(net271),
    .Y(_482_));
 sg13g2_nor3_2 _556_ (.A(net320),
    .B(net271),
    .C(net255),
    .Y(_483_));
 sg13g2_nor2_1 _557_ (.A(_234_),
    .B(_483_),
    .Y(_484_));
 sg13g2_nand3_1 _558_ (.B(_478_),
    .C(_484_),
    .A(_470_),
    .Y(_485_));
 sg13g2_nor2_2 _559_ (.A(net281),
    .B(net271),
    .Y(_486_));
 sg13g2_nor4_2 _560_ (.A(net287),
    .B(net283),
    .C(net269),
    .Y(_000_),
    .D(_468_));
 sg13g2_nand2b_2 _561_ (.Y(_001_),
    .B(net322),
    .A_N(net318));
 sg13g2_nor2_2 _562_ (.A(_456_),
    .B(_001_),
    .Y(_002_));
 sg13g2_nor4_1 _563_ (.A(net287),
    .B(net279),
    .C(net276),
    .D(net272),
    .Y(_003_));
 sg13g2_nor2_2 _564_ (.A(_465_),
    .B(_475_),
    .Y(_004_));
 sg13g2_and2_1 _565_ (.A(net316),
    .B(net318),
    .X(_005_));
 sg13g2_nand2_2 _566_ (.Y(_006_),
    .A(net315),
    .B(net319));
 sg13g2_nand3_1 _567_ (.B(net317),
    .C(net318),
    .A(net326),
    .Y(_007_));
 sg13g2_nor2_1 _568_ (.A(net277),
    .B(_006_),
    .Y(_008_));
 sg13g2_nand4_1 _569_ (.B(net326),
    .C(net315),
    .A(net323),
    .Y(_009_),
    .D(net319));
 sg13g2_nor2_1 _570_ (.A(net255),
    .B(_009_),
    .Y(_010_));
 sg13g2_nor2_2 _571_ (.A(net305),
    .B(net274),
    .Y(_011_));
 sg13g2_nor4_2 _572_ (.A(net320),
    .B(net304),
    .C(net279),
    .Y(_012_),
    .D(net274));
 sg13g2_nor2_2 _573_ (.A(_010_),
    .B(_012_),
    .Y(_013_));
 sg13g2_o21ai_1 _574_ (.B1(_013_),
    .Y(_014_),
    .A1(net255),
    .A2(_004_));
 sg13g2_nor4_1 _575_ (.A(_485_),
    .B(_000_),
    .C(_003_),
    .D(_014_),
    .Y(_015_));
 sg13g2_nor3_2 _576_ (.A(net280),
    .B(_396_),
    .C(net277),
    .Y(_016_));
 sg13g2_nor2_2 _577_ (.A(net276),
    .B(net269),
    .Y(_017_));
 sg13g2_nor3_2 _578_ (.A(net277),
    .B(net273),
    .C(net270),
    .Y(_018_));
 sg13g2_a21oi_1 _579_ (.A1(net300),
    .A2(_018_),
    .Y(_019_),
    .B1(_016_));
 sg13g2_or2_1 _580_ (.X(_020_),
    .B(_019_),
    .A(net295));
 sg13g2_nor2_2 _581_ (.A(net265),
    .B(net261),
    .Y(_021_));
 sg13g2_nor3_2 _582_ (.A(net278),
    .B(net264),
    .C(net260),
    .Y(_022_));
 sg13g2_and2_1 _583_ (.A(net285),
    .B(_022_),
    .X(_023_));
 sg13g2_nor2_2 _584_ (.A(net324),
    .B(net253),
    .Y(_024_));
 sg13g2_or2_1 _585_ (.X(_025_),
    .B(net253),
    .A(net321));
 sg13g2_nor3_2 _586_ (.A(net320),
    .B(net255),
    .C(_007_),
    .Y(_026_));
 sg13g2_nand3_1 _587_ (.B(_288_),
    .C(net250),
    .A(net324),
    .Y(_027_));
 sg13g2_nor2_1 _588_ (.A(net311),
    .B(net258),
    .Y(_028_));
 sg13g2_nand2b_1 _589_ (.Y(_029_),
    .B(_224_),
    .A_N(net258));
 sg13g2_nand3b_1 _590_ (.B(net315),
    .C(net323),
    .Y(_030_),
    .A_N(net319));
 sg13g2_nor3_1 _591_ (.A(net313),
    .B(net257),
    .C(_030_),
    .Y(_031_));
 sg13g2_o21ai_1 _592_ (.B1(_027_),
    .Y(_032_),
    .A1(_029_),
    .A2(_030_));
 sg13g2_nor2_1 _593_ (.A(net300),
    .B(net295),
    .Y(_033_));
 sg13g2_nor2_1 _594_ (.A(net272),
    .B(_009_),
    .Y(_034_));
 sg13g2_nor3_1 _595_ (.A(net273),
    .B(_009_),
    .C(_033_),
    .Y(_035_));
 sg13g2_nor4_2 _596_ (.A(_023_),
    .B(_026_),
    .C(_032_),
    .Y(_036_),
    .D(_035_));
 sg13g2_nor2_2 _597_ (.A(net263),
    .B(net254),
    .Y(_037_));
 sg13g2_nor3_1 _598_ (.A(net310),
    .B(net263),
    .C(net254),
    .Y(_038_));
 sg13g2_nor2_2 _599_ (.A(net279),
    .B(net263),
    .Y(_039_));
 sg13g2_a21oi_2 _600_ (.B1(_038_),
    .Y(_040_),
    .A2(_039_),
    .A1(net310));
 sg13g2_nand3_1 _601_ (.B(net302),
    .C(net304),
    .A(net298),
    .Y(_041_));
 sg13g2_nor3_2 _602_ (.A(net320),
    .B(net272),
    .C(net253),
    .Y(_042_));
 sg13g2_nor3_2 _603_ (.A(net320),
    .B(_468_),
    .C(net253),
    .Y(_043_));
 sg13g2_nor4_1 _604_ (.A(net320),
    .B(net310),
    .C(net257),
    .D(net253),
    .Y(_044_));
 sg13g2_a221oi_1 _605_ (.B2(net298),
    .C1(_043_),
    .B1(_042_),
    .A1(_024_),
    .Y(_045_),
    .A2(net247));
 sg13g2_o21ai_1 _606_ (.B1(_045_),
    .Y(_046_),
    .A1(_040_),
    .A2(_041_));
 sg13g2_nor3_2 _607_ (.A(net281),
    .B(_468_),
    .C(net260),
    .Y(_047_));
 sg13g2_nor3_2 _608_ (.A(net265),
    .B(net256),
    .C(_006_),
    .Y(_048_));
 sg13g2_nor3_1 _609_ (.A(net311),
    .B(net257),
    .C(_009_),
    .Y(_049_));
 sg13g2_nor4_1 _610_ (.A(net311),
    .B(net277),
    .C(net270),
    .D(net258),
    .Y(_050_));
 sg13g2_nor4_1 _611_ (.A(_047_),
    .B(_048_),
    .C(_049_),
    .D(_050_),
    .Y(_051_));
 sg13g2_nor3_1 _612_ (.A(net273),
    .B(net270),
    .C(net264),
    .Y(_052_));
 sg13g2_nor4_1 _613_ (.A(net307),
    .B(net274),
    .C(net269),
    .D(net264),
    .Y(_053_));
 sg13g2_a21oi_1 _614_ (.A1(_374_),
    .A2(_052_),
    .Y(_054_),
    .B1(_053_));
 sg13g2_nor3_1 _615_ (.A(net324),
    .B(net273),
    .C(net260),
    .Y(_055_));
 sg13g2_nor3_2 _616_ (.A(net319),
    .B(net282),
    .C(net273),
    .Y(_056_));
 sg13g2_nor2_2 _617_ (.A(net276),
    .B(net259),
    .Y(_057_));
 sg13g2_nand2_1 _618_ (.Y(_058_),
    .A(_445_),
    .B(_472_));
 sg13g2_nor3_2 _619_ (.A(net276),
    .B(_468_),
    .C(net259),
    .Y(_059_));
 sg13g2_nor4_2 _620_ (.A(net310),
    .B(net269),
    .C(net263),
    .Y(_060_),
    .D(net257));
 sg13g2_nor3_1 _621_ (.A(_056_),
    .B(_059_),
    .C(_060_),
    .Y(_061_));
 sg13g2_nor3_1 _622_ (.A(net320),
    .B(net279),
    .C(net278),
    .Y(_062_));
 sg13g2_nor4_1 _623_ (.A(net305),
    .B(net274),
    .C(net269),
    .D(net267),
    .Y(_063_));
 sg13g2_nor3_2 _624_ (.A(net276),
    .B(net274),
    .C(net259),
    .Y(_064_));
 sg13g2_nor2_2 _625_ (.A(net283),
    .B(net254),
    .Y(_065_));
 sg13g2_nor3_2 _626_ (.A(net283),
    .B(net255),
    .C(net254),
    .Y(_066_));
 sg13g2_nor4_1 _627_ (.A(_062_),
    .B(_063_),
    .C(_064_),
    .D(_066_),
    .Y(_067_));
 sg13g2_nand4_1 _628_ (.B(_054_),
    .C(_061_),
    .A(_051_),
    .Y(_068_),
    .D(_067_));
 sg13g2_o21ai_1 _629_ (.B1(net251),
    .Y(_069_),
    .A1(_024_),
    .A2(net246));
 sg13g2_inv_1 _630_ (.Y(_070_),
    .A(_069_));
 sg13g2_nor3_2 _631_ (.A(net305),
    .B(net274),
    .C(_009_),
    .Y(_071_));
 sg13g2_a21oi_1 _632_ (.A1(_475_),
    .A2(net247),
    .Y(_072_),
    .B1(_071_));
 sg13g2_a21oi_1 _633_ (.A1(_069_),
    .A2(_072_),
    .Y(_073_),
    .B1(net286));
 sg13g2_nor3_1 _634_ (.A(net280),
    .B(_452_),
    .C(net264),
    .Y(_074_));
 sg13g2_nor3_2 _635_ (.A(net281),
    .B(_452_),
    .C(net270),
    .Y(_075_));
 sg13g2_nor2_1 _636_ (.A(net279),
    .B(net267),
    .Y(_076_));
 sg13g2_nor3_2 _637_ (.A(net280),
    .B(net273),
    .C(net267),
    .Y(_077_));
 sg13g2_nor3_1 _638_ (.A(_074_),
    .B(_075_),
    .C(_077_),
    .Y(_078_));
 sg13g2_nand2_1 _639_ (.Y(_079_),
    .A(_385_),
    .B(_065_));
 sg13g2_nor4_1 _640_ (.A(net307),
    .B(net281),
    .C(net278),
    .D(net254),
    .Y(_080_));
 sg13g2_nor4_2 _641_ (.A(net307),
    .B(net281),
    .C(net275),
    .Y(_081_),
    .D(net260));
 sg13g2_nand2_1 _642_ (.Y(_082_),
    .A(net309),
    .B(_017_));
 sg13g2_nor3_1 _643_ (.A(net278),
    .B(net277),
    .C(net270),
    .Y(_083_));
 sg13g2_nor2_2 _644_ (.A(net268),
    .B(net261),
    .Y(_084_));
 sg13g2_nor3_1 _645_ (.A(net278),
    .B(net267),
    .C(net259),
    .Y(_085_));
 sg13g2_nor4_2 _646_ (.A(_080_),
    .B(_081_),
    .C(_083_),
    .Y(_086_),
    .D(_085_));
 sg13g2_nand2_1 _647_ (.Y(_087_),
    .A(_078_),
    .B(_086_));
 sg13g2_nor4_1 _648_ (.A(_046_),
    .B(_068_),
    .C(_073_),
    .D(_087_),
    .Y(_088_));
 sg13g2_nor2_1 _649_ (.A(net288),
    .B(net295),
    .Y(_089_));
 sg13g2_nand4_1 _650_ (.B(_020_),
    .C(_036_),
    .A(_015_),
    .Y(_090_),
    .D(_088_));
 sg13g2_nor4_1 _651_ (.A(net304),
    .B(net278),
    .C(net263),
    .D(net259),
    .Y(_091_));
 sg13g2_nor2_2 _652_ (.A(_039_),
    .B(_066_),
    .Y(_092_));
 sg13g2_nor4_2 _653_ (.A(net308),
    .B(net282),
    .C(net275),
    .Y(_093_),
    .D(net254));
 sg13g2_o21ai_1 _654_ (.B1(_011_),
    .Y(_094_),
    .A1(net246),
    .A2(_065_));
 sg13g2_nor3_2 _655_ (.A(net272),
    .B(net264),
    .C(net259),
    .Y(_095_));
 sg13g2_nor4_2 _656_ (.A(net310),
    .B(net276),
    .C(net261),
    .Y(_096_),
    .D(net257));
 sg13g2_nor3_2 _657_ (.A(net283),
    .B(net272),
    .C(net254),
    .Y(_097_));
 sg13g2_nor4_2 _658_ (.A(net320),
    .B(net305),
    .C(net274),
    .Y(_098_),
    .D(net253));
 sg13g2_nand2_1 _659_ (.Y(_099_),
    .A(net297),
    .B(_234_));
 sg13g2_a22oi_1 _660_ (.Y(_100_),
    .B1(net246),
    .B2(_454_),
    .A2(_037_),
    .A1(_385_));
 sg13g2_nor2_1 _661_ (.A(_468_),
    .B(_009_),
    .Y(_101_));
 sg13g2_a221oi_1 _662_ (.B2(net304),
    .C1(_101_),
    .B1(_064_),
    .A1(_385_),
    .Y(_102_),
    .A2(_037_));
 sg13g2_nand2b_2 _663_ (.Y(_103_),
    .B(net309),
    .A_N(net306));
 sg13g2_nor2_2 _664_ (.A(net303),
    .B(_103_),
    .Y(_104_));
 sg13g2_nor2_1 _665_ (.A(_025_),
    .B(_103_),
    .Y(_105_));
 sg13g2_o21ai_1 _666_ (.B1(_104_),
    .Y(_106_),
    .A1(_024_),
    .A2(_065_));
 sg13g2_or2_1 _667_ (.X(_107_),
    .B(_048_),
    .A(_486_));
 sg13g2_nor2_1 _668_ (.A(_460_),
    .B(_010_),
    .Y(_108_));
 sg13g2_or4_1 _669_ (.A(_460_),
    .B(_002_),
    .C(_010_),
    .D(_026_),
    .X(_109_));
 sg13g2_a22oi_1 _670_ (.Y(_110_),
    .B1(_457_),
    .B2(_267_),
    .A2(_445_),
    .A1(_288_));
 sg13g2_nor3_1 _671_ (.A(_002_),
    .B(_026_),
    .C(_107_),
    .Y(_111_));
 sg13g2_or2_1 _672_ (.X(_112_),
    .B(_109_),
    .A(_107_));
 sg13g2_nor3_2 _673_ (.A(net272),
    .B(net263),
    .C(net254),
    .Y(_113_));
 sg13g2_a21o_1 _674_ (.A2(_022_),
    .A1(net304),
    .B1(_113_),
    .X(_114_));
 sg13g2_or2_1 _675_ (.X(_115_),
    .B(_114_),
    .A(_059_));
 sg13g2_nor4_2 _676_ (.A(_180_),
    .B(net302),
    .C(net266),
    .Y(_116_),
    .D(_103_));
 sg13g2_nor4_2 _677_ (.A(net314),
    .B(net263),
    .C(net261),
    .Y(_117_),
    .D(net257));
 sg13g2_nor2_1 _678_ (.A(_116_),
    .B(_117_),
    .Y(_118_));
 sg13g2_a21oi_1 _679_ (.A1(net246),
    .A2(_104_),
    .Y(_119_),
    .B1(_117_));
 sg13g2_a221oi_1 _680_ (.B2(_104_),
    .C1(_116_),
    .B1(net246),
    .A1(_021_),
    .Y(_120_),
    .A2(net247));
 sg13g2_nor3_1 _681_ (.A(_096_),
    .B(_097_),
    .C(_098_),
    .Y(_121_));
 sg13g2_nor4_1 _682_ (.A(_043_),
    .B(_044_),
    .C(_091_),
    .D(_095_),
    .Y(_122_));
 sg13g2_nand4_1 _683_ (.B(_120_),
    .C(_121_),
    .A(_004_),
    .Y(_123_),
    .D(_122_));
 sg13g2_nand4_1 _684_ (.B(_094_),
    .C(_102_),
    .A(_092_),
    .Y(_124_),
    .D(_106_));
 sg13g2_nor4_1 _685_ (.A(_112_),
    .B(_115_),
    .C(_123_),
    .D(_124_),
    .Y(_125_));
 sg13g2_nand2b_1 _686_ (.Y(_126_),
    .B(_125_),
    .A_N(_099_));
 sg13g2_a21o_1 _687_ (.A2(_126_),
    .A1(_090_),
    .B1(net289),
    .X(_127_));
 sg13g2_nand2_2 _688_ (.Y(_128_),
    .A(_234_),
    .B(net5));
 sg13g2_a21oi_1 _689_ (.A1(net321),
    .A2(net317),
    .Y(_129_),
    .B1(_128_));
 sg13g2_nor2b_1 _690_ (.A(_482_),
    .B_N(_129_),
    .Y(_130_));
 sg13g2_and2_1 _691_ (.A(net253),
    .B(_130_),
    .X(_131_));
 sg13g2_nand2_1 _692_ (.Y(_132_),
    .A(net296),
    .B(net292));
 sg13g2_inv_1 _693_ (.Y(_133_),
    .A(_132_));
 sg13g2_nand2_1 _694_ (.Y(_134_),
    .A(net309),
    .B(net279));
 sg13g2_or2_2 _695_ (.X(_135_),
    .B(_134_),
    .A(net302));
 sg13g2_nand3_1 _696_ (.B(_288_),
    .C(net276),
    .A(net313),
    .Y(_136_));
 sg13g2_o21ai_1 _697_ (.B1(_136_),
    .Y(_137_),
    .A1(net313),
    .A2(_009_));
 sg13g2_a21oi_1 _698_ (.A1(net312),
    .A2(_457_),
    .Y(_138_),
    .B1(_137_));
 sg13g2_nand2_2 _699_ (.Y(_139_),
    .A(net276),
    .B(_005_));
 sg13g2_a21oi_1 _700_ (.A1(_058_),
    .A2(_139_),
    .Y(_140_),
    .B1(net313));
 sg13g2_a21oi_1 _701_ (.A1(net284),
    .A2(_021_),
    .Y(_141_),
    .B1(_140_));
 sg13g2_a22oi_1 _702_ (.Y(_142_),
    .B1(_462_),
    .B2(_005_),
    .A2(_445_),
    .A1(_288_));
 sg13g2_a21oi_2 _703_ (.B1(net284),
    .Y(_143_),
    .A2(_142_),
    .A1(_476_));
 sg13g2_nand3b_1 _704_ (.B(_141_),
    .C(_138_),
    .Y(_144_),
    .A_N(_143_));
 sg13g2_a21oi_1 _705_ (.A1(_135_),
    .A2(_144_),
    .Y(_145_),
    .B1(_132_));
 sg13g2_o21ai_1 _706_ (.B1(net290),
    .Y(_146_),
    .A1(_131_),
    .A2(_145_));
 sg13g2_nand3_1 _707_ (.B(_127_),
    .C(_146_),
    .A(net6),
    .Y(_147_));
 sg13g2_xor2_1 _708_ (.B(_147_),
    .A(net293),
    .X(uo_out[6]));
 sg13g2_o21ai_1 _709_ (.B1(_467_),
    .Y(_148_),
    .A1(_460_),
    .A2(_465_));
 sg13g2_nor2_1 _710_ (.A(_042_),
    .B(_113_),
    .Y(_149_));
 sg13g2_nand2_1 _711_ (.Y(_150_),
    .A(net287),
    .B(_042_));
 sg13g2_a21oi_1 _712_ (.A1(_148_),
    .A2(_149_),
    .Y(_151_),
    .B1(net298));
 sg13g2_a221oi_1 _713_ (.B2(_467_),
    .C1(_064_),
    .B1(_065_),
    .A1(_310_),
    .Y(_152_),
    .A2(net249));
 sg13g2_nand2b_1 _714_ (.Y(_153_),
    .B(_097_),
    .A_N(_089_));
 sg13g2_a21oi_1 _715_ (.A1(_460_),
    .A2(net252),
    .Y(_154_),
    .B1(_074_));
 sg13g2_nand2_2 _716_ (.Y(_155_),
    .A(_153_),
    .B(_154_));
 sg13g2_a21oi_1 _717_ (.A1(net286),
    .A2(_043_),
    .Y(_156_),
    .B1(_000_));
 sg13g2_nand2_1 _718_ (.Y(_157_),
    .A(_152_),
    .B(_156_));
 sg13g2_nor4_2 _719_ (.A(net311),
    .B(net281),
    .C(net270),
    .Y(_158_),
    .D(net258));
 sg13g2_nand2_1 _720_ (.Y(_159_),
    .A(net285),
    .B(_158_));
 sg13g2_nand2_1 _721_ (.Y(_160_),
    .A(_460_),
    .B(net248));
 sg13g2_and2_1 _722_ (.A(_159_),
    .B(_160_),
    .X(_161_));
 sg13g2_nand2_1 _723_ (.Y(_162_),
    .A(net4),
    .B(_017_));
 sg13g2_a21oi_1 _724_ (.A1(_004_),
    .A2(_162_),
    .Y(_163_),
    .B1(net255));
 sg13g2_nor3_1 _725_ (.A(net296),
    .B(_476_),
    .C(_029_),
    .Y(_164_));
 sg13g2_nor2_1 _726_ (.A(_062_),
    .B(_071_),
    .Y(_165_));
 sg13g2_a22oi_1 _727_ (.Y(_166_),
    .B1(_039_),
    .B2(_467_),
    .A2(_002_),
    .A1(_454_));
 sg13g2_nor2_1 _728_ (.A(net301),
    .B(_166_),
    .Y(_167_));
 sg13g2_nor4_1 _729_ (.A(net308),
    .B(_267_),
    .C(net275),
    .D(_139_),
    .Y(_168_));
 sg13g2_a221oi_1 _730_ (.B2(_011_),
    .C1(_098_),
    .B1(_037_),
    .A1(net288),
    .Y(_170_),
    .A2(_034_));
 sg13g2_nor4_2 _731_ (.A(net308),
    .B(net275),
    .C(_456_),
    .Y(_171_),
    .D(_474_));
 sg13g2_a221oi_1 _732_ (.B2(_039_),
    .C1(_171_),
    .B1(net252),
    .A1(_453_),
    .Y(_172_),
    .A2(_465_));
 sg13g2_nand2_1 _733_ (.Y(_173_),
    .A(_170_),
    .B(_172_));
 sg13g2_a22oi_1 _734_ (.Y(_174_),
    .B1(_066_),
    .B2(net295),
    .A2(_461_),
    .A1(_374_));
 sg13g2_nand2_1 _735_ (.Y(_175_),
    .A(_165_),
    .B(_174_));
 sg13g2_nor4_1 _736_ (.A(_164_),
    .B(_167_),
    .C(_173_),
    .D(_175_),
    .Y(_176_));
 sg13g2_nand3_1 _737_ (.B(net252),
    .C(_057_),
    .A(net286),
    .Y(_177_));
 sg13g2_nor4_1 _738_ (.A(_191_),
    .B(net308),
    .C(net278),
    .D(net264),
    .Y(_178_));
 sg13g2_nor4_2 _739_ (.A(net317),
    .B(net313),
    .C(net258),
    .Y(_179_),
    .D(_001_));
 sg13g2_nand2_1 _740_ (.Y(_181_),
    .A(net295),
    .B(_059_));
 sg13g2_nor4_1 _741_ (.A(_016_),
    .B(_093_),
    .C(_178_),
    .D(_179_),
    .Y(_182_));
 sg13g2_nor4_1 _742_ (.A(_483_),
    .B(_012_),
    .C(_018_),
    .D(_060_),
    .Y(_183_));
 sg13g2_and2_1 _743_ (.A(_086_),
    .B(_183_),
    .X(_184_));
 sg13g2_a22oi_1 _744_ (.Y(_185_),
    .B1(_077_),
    .B2(net288),
    .A2(_048_),
    .A1(net285));
 sg13g2_nor3_1 _745_ (.A(_234_),
    .B(_056_),
    .C(_117_),
    .Y(_186_));
 sg13g2_nand4_1 _746_ (.B(_181_),
    .C(_185_),
    .A(_177_),
    .Y(_187_),
    .D(_186_));
 sg13g2_nor2_1 _747_ (.A(_151_),
    .B(_187_),
    .Y(_188_));
 sg13g2_nand4_1 _748_ (.B(_182_),
    .C(_184_),
    .A(_161_),
    .Y(_189_),
    .D(_188_));
 sg13g2_nor3_1 _749_ (.A(_155_),
    .B(_157_),
    .C(_163_),
    .Y(_190_));
 sg13g2_nand2_1 _750_ (.Y(_192_),
    .A(_176_),
    .B(_190_));
 sg13g2_and2_1 _751_ (.A(_037_),
    .B(_104_),
    .X(_193_));
 sg13g2_nand3_1 _752_ (.B(_108_),
    .C(_162_),
    .A(_004_),
    .Y(_194_));
 sg13g2_a21oi_2 _753_ (.B1(_099_),
    .Y(_195_),
    .A2(_310_),
    .A1(net299));
 sg13g2_a21oi_1 _754_ (.A1(net249),
    .A2(_021_),
    .Y(_196_),
    .B1(_096_));
 sg13g2_nand2_1 _755_ (.Y(_197_),
    .A(_195_),
    .B(_196_));
 sg13g2_nor4_1 _756_ (.A(_107_),
    .B(_193_),
    .C(_194_),
    .D(_197_),
    .Y(_198_));
 sg13g2_a21oi_2 _757_ (.B1(_042_),
    .Y(_199_),
    .A2(net246),
    .A1(net251));
 sg13g2_nor4_2 _758_ (.A(_042_),
    .B(_070_),
    .C(_097_),
    .Y(_200_),
    .D(_115_));
 sg13g2_and2_1 _759_ (.A(_079_),
    .B(_102_),
    .X(_201_));
 sg13g2_nand4_1 _760_ (.B(_198_),
    .C(_200_),
    .A(_106_),
    .Y(_203_),
    .D(_201_));
 sg13g2_o21ai_1 _761_ (.B1(_203_),
    .Y(_204_),
    .A1(_189_),
    .A2(_192_));
 sg13g2_nand2_1 _762_ (.Y(_205_),
    .A(net292),
    .B(_135_));
 sg13g2_nor4_2 _763_ (.A(net322),
    .B(_180_),
    .C(_191_),
    .Y(_206_),
    .D(net284));
 sg13g2_nor2_1 _764_ (.A(_267_),
    .B(net271),
    .Y(_207_));
 sg13g2_nor2_1 _765_ (.A(_475_),
    .B(_207_),
    .Y(_208_));
 sg13g2_nor2_1 _766_ (.A(net312),
    .B(_208_),
    .Y(_209_));
 sg13g2_nor3_1 _767_ (.A(_137_),
    .B(_206_),
    .C(_209_),
    .Y(_210_));
 sg13g2_o21ai_1 _768_ (.B1(_142_),
    .Y(_211_),
    .A1(_267_),
    .A2(net261));
 sg13g2_nand2_1 _769_ (.Y(_212_),
    .A(net312),
    .B(_211_));
 sg13g2_a22oi_1 _770_ (.Y(_214_),
    .B1(_474_),
    .B2(net316),
    .A2(_457_),
    .A1(_445_));
 sg13g2_a21oi_1 _771_ (.A1(_466_),
    .A2(_214_),
    .Y(_215_),
    .B1(net313));
 sg13g2_nand3_1 _772_ (.B(_210_),
    .C(_212_),
    .A(_141_),
    .Y(_216_));
 sg13g2_nand2b_1 _773_ (.Y(_217_),
    .B(_216_),
    .A_N(_205_));
 sg13g2_nand2_1 _774_ (.Y(_218_),
    .A(net297),
    .B(net289));
 sg13g2_nor2_1 _775_ (.A(net287),
    .B(net247),
    .Y(_219_));
 sg13g2_nand2_1 _776_ (.Y(_220_),
    .A(net302),
    .B(_103_));
 sg13g2_a221oi_1 _777_ (.B2(_220_),
    .C1(net291),
    .B1(_219_),
    .A1(net287),
    .Y(_221_),
    .A2(net255));
 sg13g2_nor2_1 _778_ (.A(_218_),
    .B(_221_),
    .Y(_222_));
 sg13g2_a221oi_1 _779_ (.B2(_222_),
    .C1(_213_),
    .B1(_217_),
    .A1(_245_),
    .Y(_223_),
    .A2(_204_));
 sg13g2_xnor2_1 _780_ (.Y(uo_out[5]),
    .A(net294),
    .B(_223_));
 sg13g2_nor4_2 _781_ (.A(net307),
    .B(net275),
    .C(net264),
    .Y(_225_),
    .D(net261));
 sg13g2_nor4_1 _782_ (.A(_075_),
    .B(_093_),
    .C(_171_),
    .D(_225_),
    .Y(_226_));
 sg13g2_nand2b_1 _783_ (.Y(_227_),
    .B(net249),
    .A_N(_477_));
 sg13g2_o21ai_1 _784_ (.B1(_454_),
    .Y(_228_),
    .A1(_460_),
    .A2(_002_));
 sg13g2_nand3_1 _785_ (.B(_227_),
    .C(_228_),
    .A(_226_),
    .Y(_229_));
 sg13g2_inv_1 _786_ (.Y(_230_),
    .A(_229_));
 sg13g2_and2_1 _787_ (.A(net247),
    .B(_037_),
    .X(_231_));
 sg13g2_o21ai_1 _788_ (.B1(net284),
    .Y(_232_),
    .A1(net302),
    .A2(net306));
 sg13g2_nor2_1 _789_ (.A(_477_),
    .B(_232_),
    .Y(_233_));
 sg13g2_a221oi_1 _790_ (.B2(net297),
    .C1(_233_),
    .B1(_231_),
    .A1(_310_),
    .Y(_235_),
    .A2(_385_));
 sg13g2_nand3b_1 _791_ (.B(_013_),
    .C(net292),
    .Y(_236_),
    .A_N(_049_));
 sg13g2_nand2_1 _792_ (.Y(_237_),
    .A(net278),
    .B(net255));
 sg13g2_a221oi_1 _793_ (.B2(_039_),
    .C1(_236_),
    .B1(_237_),
    .A1(net285),
    .Y(_238_),
    .A2(_048_));
 sg13g2_a22oi_1 _794_ (.Y(_239_),
    .B1(_002_),
    .B2(net247),
    .A2(_467_),
    .A1(_460_));
 sg13g2_nand2_1 _795_ (.Y(_240_),
    .A(net298),
    .B(_469_));
 sg13g2_nand2_1 _796_ (.Y(_241_),
    .A(net302),
    .B(_038_));
 sg13g2_a22oi_1 _797_ (.Y(_242_),
    .B1(_071_),
    .B2(net286),
    .A2(_042_),
    .A1(net298));
 sg13g2_nand4_1 _798_ (.B(_240_),
    .C(_241_),
    .A(_239_),
    .Y(_243_),
    .D(_242_));
 sg13g2_nand2_1 _799_ (.Y(_244_),
    .A(_417_),
    .B(_034_));
 sg13g2_nor2_1 _800_ (.A(_018_),
    .B(_095_),
    .Y(_246_));
 sg13g2_o21ai_1 _801_ (.B1(net288),
    .Y(_247_),
    .A1(_018_),
    .A2(_095_));
 sg13g2_nand2_1 _802_ (.Y(_248_),
    .A(_374_),
    .B(_077_));
 sg13g2_a22oi_1 _803_ (.Y(_249_),
    .B1(_158_),
    .B2(net296),
    .A2(_077_),
    .A1(_374_));
 sg13g2_a221oi_1 _804_ (.B2(net251),
    .C1(_022_),
    .B1(net246),
    .A1(_385_),
    .Y(_250_),
    .A2(_017_));
 sg13g2_nand4_1 _805_ (.B(_247_),
    .C(_249_),
    .A(_244_),
    .Y(_251_),
    .D(_250_));
 sg13g2_nor4_1 _806_ (.A(_155_),
    .B(_157_),
    .C(_243_),
    .D(_251_),
    .Y(_252_));
 sg13g2_nand4_1 _807_ (.B(_235_),
    .C(_238_),
    .A(_230_),
    .Y(_253_),
    .D(_252_));
 sg13g2_a21oi_1 _808_ (.A1(net249),
    .A2(_021_),
    .Y(_254_),
    .B1(_043_));
 sg13g2_nand3_1 _809_ (.B(_092_),
    .C(_254_),
    .A(_079_),
    .Y(_255_));
 sg13g2_nand4_1 _810_ (.B(_102_),
    .C(_118_),
    .A(_477_),
    .Y(_257_),
    .D(_195_));
 sg13g2_nor2_1 _811_ (.A(_255_),
    .B(_257_),
    .Y(_258_));
 sg13g2_a21oi_1 _812_ (.A1(_200_),
    .A2(_258_),
    .Y(_259_),
    .B1(net289));
 sg13g2_nor4_1 _813_ (.A(net309),
    .B(_486_),
    .C(_037_),
    .D(_084_),
    .Y(_260_));
 sg13g2_a21oi_1 _814_ (.A1(net310),
    .A2(_025_),
    .Y(_261_),
    .B1(_260_));
 sg13g2_o21ai_1 _815_ (.B1(_135_),
    .Y(_262_),
    .A1(_143_),
    .A2(_261_));
 sg13g2_a22oi_1 _816_ (.Y(_263_),
    .B1(_005_),
    .B2(net268),
    .A2(_462_),
    .A1(net315));
 sg13g2_nor2_1 _817_ (.A(_002_),
    .B(_128_),
    .Y(_264_));
 sg13g2_a22oi_1 _818_ (.Y(_265_),
    .B1(_263_),
    .B2(_264_),
    .A2(_262_),
    .A1(_133_));
 sg13g2_a22oi_1 _819_ (.Y(_266_),
    .B1(_265_),
    .B2(net289),
    .A2(_259_),
    .A1(_253_));
 sg13g2_nor2_1 _820_ (.A(_213_),
    .B(_266_),
    .Y(_268_));
 sg13g2_xnor2_1 _821_ (.Y(uo_out[4]),
    .A(net293),
    .B(_268_));
 sg13g2_nand2_1 _822_ (.Y(_269_),
    .A(_077_),
    .B(_089_));
 sg13g2_o21ai_1 _823_ (.B1(net250),
    .Y(_270_),
    .A1(_310_),
    .A2(_460_));
 sg13g2_nand4_1 _824_ (.B(_159_),
    .C(_181_),
    .A(_027_),
    .Y(_271_),
    .D(_270_));
 sg13g2_nor4_1 _825_ (.A(net311),
    .B(net280),
    .C(net267),
    .D(net258),
    .Y(_272_));
 sg13g2_or4_1 _826_ (.A(_022_),
    .B(_083_),
    .C(_085_),
    .D(_272_),
    .X(_273_));
 sg13g2_or2_1 _827_ (.X(_274_),
    .B(_026_),
    .A(_000_));
 sg13g2_o21ai_1 _828_ (.B1(net286),
    .Y(_275_),
    .A1(_231_),
    .A2(_274_));
 sg13g2_nand3_1 _829_ (.B(net249),
    .C(_084_),
    .A(net5),
    .Y(_276_));
 sg13g2_nand2_2 _830_ (.Y(_278_),
    .A(net297),
    .B(_043_));
 sg13g2_and2_1 _831_ (.A(net247),
    .B(_065_),
    .X(_279_));
 sg13g2_o21ai_1 _832_ (.B1(_008_),
    .Y(_280_),
    .A1(_453_),
    .A2(net251));
 sg13g2_nor2_1 _833_ (.A(net256),
    .B(_030_),
    .Y(_281_));
 sg13g2_or2_1 _834_ (.X(_282_),
    .B(_030_),
    .A(net256));
 sg13g2_or3_1 _835_ (.A(_016_),
    .B(_047_),
    .C(_279_),
    .X(_283_));
 sg13g2_nor4_2 _836_ (.A(_229_),
    .B(_271_),
    .C(_273_),
    .Y(_284_),
    .D(_283_));
 sg13g2_nor2_1 _837_ (.A(_060_),
    .B(_098_),
    .Y(_285_));
 sg13g2_nand4_1 _838_ (.B(_069_),
    .C(_150_),
    .A(_478_),
    .Y(_286_),
    .D(_285_));
 sg13g2_nand4_1 _839_ (.B(_269_),
    .C(_276_),
    .A(_246_),
    .Y(_287_),
    .D(_278_));
 sg13g2_a22oi_1 _840_ (.Y(_289_),
    .B1(net247),
    .B2(_475_),
    .A2(_011_),
    .A1(_310_));
 sg13g2_nand4_1 _841_ (.B(_280_),
    .C(_282_),
    .A(_148_),
    .Y(_290_),
    .D(_289_));
 sg13g2_nor4_2 _842_ (.A(_155_),
    .B(_286_),
    .C(_287_),
    .Y(_291_),
    .D(_290_));
 sg13g2_nand4_1 _843_ (.B(_275_),
    .C(_284_),
    .A(net291),
    .Y(_292_),
    .D(_291_));
 sg13g2_a21oi_1 _844_ (.A1(net5),
    .A2(_084_),
    .Y(_293_),
    .B1(_225_));
 sg13g2_nand2_1 _845_ (.Y(_294_),
    .A(_477_),
    .B(_293_));
 sg13g2_and3_1 _846_ (.X(_295_),
    .A(_094_),
    .B(_195_),
    .C(_199_));
 sg13g2_a21oi_1 _847_ (.A1(_024_),
    .A2(_104_),
    .Y(_296_),
    .B1(_059_));
 sg13g2_nand2_1 _848_ (.Y(_297_),
    .A(_100_),
    .B(_296_));
 sg13g2_nand2b_1 _849_ (.Y(_298_),
    .B(_120_),
    .A_N(_109_));
 sg13g2_nor4_1 _850_ (.A(_231_),
    .B(_294_),
    .C(_297_),
    .D(_298_),
    .Y(_300_));
 sg13g2_nand3b_1 _851_ (.B(_295_),
    .C(_300_),
    .Y(_301_),
    .A_N(_255_));
 sg13g2_a21oi_1 _852_ (.A1(_292_),
    .A2(_301_),
    .Y(_302_),
    .B1(net289));
 sg13g2_nor2_2 _853_ (.A(_143_),
    .B(_206_),
    .Y(_303_));
 sg13g2_a21oi_1 _854_ (.A1(net261),
    .A2(net253),
    .Y(_304_),
    .B1(net321));
 sg13g2_nor2_1 _855_ (.A(net312),
    .B(_110_),
    .Y(_305_));
 sg13g2_a21oi_1 _856_ (.A1(net284),
    .A2(_304_),
    .Y(_306_),
    .B1(_305_));
 sg13g2_nand4_1 _857_ (.B(_082_),
    .C(_303_),
    .A(_040_),
    .Y(_307_),
    .D(_306_));
 sg13g2_nor2b_1 _858_ (.A(_205_),
    .B_N(_307_),
    .Y(_308_));
 sg13g2_a22oi_1 _859_ (.Y(_309_),
    .B1(net257),
    .B2(net299),
    .A2(net306),
    .A1(net284));
 sg13g2_nor3_1 _860_ (.A(net291),
    .B(_454_),
    .C(_309_),
    .Y(_311_));
 sg13g2_nor3_1 _861_ (.A(_218_),
    .B(_308_),
    .C(_311_),
    .Y(_312_));
 sg13g2_nor3_1 _862_ (.A(_213_),
    .B(_302_),
    .C(_312_),
    .Y(_313_));
 sg13g2_xnor2_1 _863_ (.Y(uo_out[3]),
    .A(net293),
    .B(_313_));
 sg13g2_a21oi_1 _864_ (.A1(_288_),
    .A2(_462_),
    .Y(_314_),
    .B1(net312));
 sg13g2_nand4_1 _865_ (.B(_139_),
    .C(_214_),
    .A(_110_),
    .Y(_315_),
    .D(_314_));
 sg13g2_a21oi_1 _866_ (.A1(net268),
    .A2(net265),
    .Y(_316_),
    .B1(net280));
 sg13g2_nand3_1 _867_ (.B(_464_),
    .C(_058_),
    .A(net312),
    .Y(_317_));
 sg13g2_o21ai_1 _868_ (.B1(_315_),
    .Y(_318_),
    .A1(_316_),
    .A2(_317_));
 sg13g2_nand3_1 _869_ (.B(_303_),
    .C(_318_),
    .A(_448_),
    .Y(_319_));
 sg13g2_o21ai_1 _870_ (.B1(_135_),
    .Y(_321_),
    .A1(net300),
    .A2(_448_));
 sg13g2_nand2b_1 _871_ (.Y(_322_),
    .B(_319_),
    .A_N(_321_));
 sg13g2_nand3_1 _872_ (.B(net264),
    .C(_001_),
    .A(net317),
    .Y(_323_));
 sg13g2_nor2_1 _873_ (.A(net325),
    .B(_001_),
    .Y(_324_));
 sg13g2_nor2_1 _874_ (.A(_128_),
    .B(_324_),
    .Y(_325_));
 sg13g2_a221oi_1 _875_ (.B2(_325_),
    .C1(_245_),
    .B1(_323_),
    .A1(_133_),
    .Y(_326_),
    .A2(_322_));
 sg13g2_nor3_1 _876_ (.A(net280),
    .B(_462_),
    .C(net256),
    .Y(_327_));
 sg13g2_a21oi_1 _877_ (.A1(net251),
    .A2(_024_),
    .Y(_328_),
    .B1(_064_));
 sg13g2_nor4_2 _878_ (.A(net307),
    .B(net275),
    .C(net267),
    .Y(_329_),
    .D(net259));
 sg13g2_nor2b_1 _879_ (.A(_456_),
    .B_N(_001_),
    .Y(_330_));
 sg13g2_o21ai_1 _880_ (.B1(_011_),
    .Y(_332_),
    .A1(_017_),
    .A2(_076_));
 sg13g2_a21oi_1 _881_ (.A1(_466_),
    .A2(_214_),
    .Y(_333_),
    .B1(net256));
 sg13g2_nor4_1 _882_ (.A(net300),
    .B(net281),
    .C(net270),
    .D(_468_),
    .Y(_334_));
 sg13g2_nor2_1 _883_ (.A(_016_),
    .B(_334_),
    .Y(_335_));
 sg13g2_a22oi_1 _884_ (.Y(_336_),
    .B1(_066_),
    .B2(net285),
    .A2(_482_),
    .A1(net252));
 sg13g2_nand2_1 _885_ (.Y(_337_),
    .A(net285),
    .B(_059_));
 sg13g2_nor4_1 _886_ (.A(_018_),
    .B(_055_),
    .C(_095_),
    .D(_333_),
    .Y(_338_));
 sg13g2_a22oi_1 _887_ (.Y(_339_),
    .B1(_097_),
    .B2(net300),
    .A2(_062_),
    .A1(net325));
 sg13g2_and2_1 _888_ (.A(_328_),
    .B(_339_),
    .X(_340_));
 sg13g2_nor4_1 _889_ (.A(_483_),
    .B(_096_),
    .C(_225_),
    .D(_279_),
    .Y(_341_));
 sg13g2_and4_1 _890_ (.A(_332_),
    .B(_337_),
    .C(_340_),
    .D(_341_),
    .X(_343_));
 sg13g2_nand3_1 _891_ (.B(_335_),
    .C(_336_),
    .A(_244_),
    .Y(_344_));
 sg13g2_a22oi_1 _892_ (.Y(_345_),
    .B1(_084_),
    .B2(net248),
    .A2(_057_),
    .A1(net249));
 sg13g2_nor2_1 _893_ (.A(_327_),
    .B(_329_),
    .Y(_346_));
 sg13g2_nand3_1 _894_ (.B(_345_),
    .C(_346_),
    .A(_078_),
    .Y(_347_));
 sg13g2_nand3_1 _895_ (.B(_159_),
    .C(_160_),
    .A(_086_),
    .Y(_348_));
 sg13g2_nor4_1 _896_ (.A(_243_),
    .B(_344_),
    .C(_347_),
    .D(_348_),
    .Y(_349_));
 sg13g2_and4_1 _897_ (.A(net292),
    .B(_338_),
    .C(_343_),
    .D(_349_),
    .X(_350_));
 sg13g2_nor3_1 _898_ (.A(_465_),
    .B(_475_),
    .C(_059_),
    .Y(_351_));
 sg13g2_nor3_1 _899_ (.A(_017_),
    .B(_076_),
    .C(_097_),
    .Y(_352_));
 sg13g2_a22oi_1 _900_ (.Y(_354_),
    .B1(net246),
    .B2(net249),
    .A2(_022_),
    .A1(net304));
 sg13g2_nand2_1 _901_ (.Y(_355_),
    .A(_352_),
    .B(_354_));
 sg13g2_nand4_1 _902_ (.B(_195_),
    .C(_254_),
    .A(_119_),
    .Y(_356_),
    .D(_351_));
 sg13g2_nor3_1 _903_ (.A(_112_),
    .B(_355_),
    .C(_356_),
    .Y(_357_));
 sg13g2_nor3_1 _904_ (.A(net290),
    .B(_350_),
    .C(_357_),
    .Y(_358_));
 sg13g2_o21ai_1 _905_ (.B1(net6),
    .Y(_359_),
    .A1(_326_),
    .A2(_358_));
 sg13g2_xor2_1 _906_ (.B(_359_),
    .A(net294),
    .X(uo_out[2]));
 sg13g2_and2_1 _907_ (.A(_363_),
    .B(_052_),
    .X(_360_));
 sg13g2_a21oi_1 _908_ (.A1(net325),
    .A2(net295),
    .Y(_361_),
    .B1(net300));
 sg13g2_a21oi_1 _909_ (.A1(net251),
    .A2(_024_),
    .Y(_362_),
    .B1(_329_));
 sg13g2_nand3_1 _910_ (.B(net248),
    .C(_084_),
    .A(net285),
    .Y(_364_));
 sg13g2_nand2b_1 _911_ (.Y(_365_),
    .B(net250),
    .A_N(_214_));
 sg13g2_nand2_1 _912_ (.Y(_366_),
    .A(net296),
    .B(_048_));
 sg13g2_nand4_1 _913_ (.B(_364_),
    .C(_365_),
    .A(_013_),
    .Y(_367_),
    .D(_366_));
 sg13g2_o21ai_1 _914_ (.B1(_089_),
    .Y(_368_),
    .A1(_461_),
    .A2(_097_));
 sg13g2_o21ai_1 _915_ (.B1(_368_),
    .Y(_369_),
    .A1(net296),
    .A2(_362_));
 sg13g2_a21oi_1 _916_ (.A1(net285),
    .A2(_059_),
    .Y(_370_),
    .B1(_334_));
 sg13g2_a221oi_1 _917_ (.B2(_361_),
    .C1(_360_),
    .B1(_055_),
    .A1(net300),
    .Y(_371_),
    .A2(_018_));
 sg13g2_nand4_1 _918_ (.B(_278_),
    .C(_370_),
    .A(_165_),
    .Y(_372_),
    .D(_371_));
 sg13g2_nand3_1 _919_ (.B(_249_),
    .C(_336_),
    .A(_170_),
    .Y(_373_));
 sg13g2_a21o_1 _920_ (.A2(_486_),
    .A1(net250),
    .B1(_225_),
    .X(_375_));
 sg13g2_or4_1 _921_ (.A(_081_),
    .B(_178_),
    .C(_273_),
    .D(_375_),
    .X(_376_));
 sg13g2_a221oi_1 _922_ (.B2(net248),
    .C1(_031_),
    .B1(_008_),
    .A1(_288_),
    .Y(_377_),
    .A2(net249));
 sg13g2_nor4_1 _923_ (.A(_050_),
    .B(_075_),
    .C(_095_),
    .D(_179_),
    .Y(_378_));
 sg13g2_nand2_1 _924_ (.Y(_379_),
    .A(_377_),
    .B(_378_));
 sg13g2_or4_1 _925_ (.A(_369_),
    .B(_373_),
    .C(_376_),
    .D(_379_),
    .X(_380_));
 sg13g2_nor4_2 _926_ (.A(_151_),
    .B(_367_),
    .C(_372_),
    .Y(_381_),
    .D(_380_));
 sg13g2_nand2_1 _927_ (.Y(_382_),
    .A(_092_),
    .B(_196_));
 sg13g2_a21oi_1 _928_ (.A1(_065_),
    .A2(_104_),
    .Y(_383_),
    .B1(_475_));
 sg13g2_nor2_1 _929_ (.A(_043_),
    .B(_113_),
    .Y(_384_));
 sg13g2_nand3_1 _930_ (.B(_383_),
    .C(_384_),
    .A(_111_),
    .Y(_386_));
 sg13g2_nor3_1 _931_ (.A(_355_),
    .B(_382_),
    .C(_386_),
    .Y(_387_));
 sg13g2_a22oi_1 _932_ (.Y(_388_),
    .B1(_387_),
    .B2(_195_),
    .A2(_381_),
    .A1(net291));
 sg13g2_a21oi_1 _933_ (.A1(_303_),
    .A2(_318_),
    .Y(_389_),
    .B1(_205_));
 sg13g2_nand3_1 _934_ (.B(net274),
    .C(net257),
    .A(net299),
    .Y(_390_));
 sg13g2_o21ai_1 _935_ (.B1(_390_),
    .Y(_391_),
    .A1(net299),
    .A2(_385_));
 sg13g2_a21oi_1 _936_ (.A1(_103_),
    .A2(_391_),
    .Y(_392_),
    .B1(net291));
 sg13g2_nor3_1 _937_ (.A(_218_),
    .B(_389_),
    .C(_392_),
    .Y(_393_));
 sg13g2_nor2_1 _938_ (.A(_213_),
    .B(_393_),
    .Y(_394_));
 sg13g2_o21ai_1 _939_ (.B1(_394_),
    .Y(_395_),
    .A1(net289),
    .A2(_388_));
 sg13g2_xor2_1 _940_ (.B(_395_),
    .A(net294),
    .X(uo_out[1]));
 sg13g2_o21ai_1 _941_ (.B1(_030_),
    .Y(_397_),
    .A1(net282),
    .A2(net279));
 sg13g2_o21ai_1 _942_ (.B1(net312),
    .Y(_398_),
    .A1(_207_),
    .A2(_397_));
 sg13g2_nor4_1 _943_ (.A(_140_),
    .B(_215_),
    .C(_305_),
    .D(_316_),
    .Y(_399_));
 sg13g2_nand3_1 _944_ (.B(_398_),
    .C(_399_),
    .A(_303_),
    .Y(_400_));
 sg13g2_a21oi_1 _945_ (.A1(_135_),
    .A2(_400_),
    .Y(_401_),
    .B1(_132_));
 sg13g2_o21ai_1 _946_ (.B1(_139_),
    .Y(_402_),
    .A1(_267_),
    .A2(net261));
 sg13g2_nor3_1 _947_ (.A(_128_),
    .B(_330_),
    .C(_402_),
    .Y(_403_));
 sg13g2_o21ai_1 _948_ (.B1(net295),
    .Y(_404_),
    .A1(_026_),
    .A2(_329_));
 sg13g2_nor4_1 _949_ (.A(net272),
    .B(net268),
    .C(net260),
    .D(_033_),
    .Y(_405_));
 sg13g2_nand2_1 _950_ (.Y(_407_),
    .A(net287),
    .B(_047_));
 sg13g2_a21oi_1 _951_ (.A1(net269),
    .A2(net259),
    .Y(_408_),
    .B1(net283));
 sg13g2_nand2_1 _952_ (.Y(_409_),
    .A(net251),
    .B(_408_));
 sg13g2_nand2_1 _953_ (.Y(_410_),
    .A(net3),
    .B(_465_));
 sg13g2_o21ai_1 _954_ (.B1(_407_),
    .Y(_411_),
    .A1(net256),
    .A2(_410_));
 sg13g2_nor3_1 _955_ (.A(_018_),
    .B(_022_),
    .C(_281_),
    .Y(_412_));
 sg13g2_nand3_1 _956_ (.B(_404_),
    .C(_412_),
    .A(_335_),
    .Y(_413_));
 sg13g2_nand4_1 _957_ (.B(_278_),
    .C(_328_),
    .A(_199_),
    .Y(_414_),
    .D(_409_));
 sg13g2_a221oi_1 _958_ (.B2(net287),
    .C1(_117_),
    .B1(_113_),
    .A1(_385_),
    .Y(_415_),
    .A2(_037_));
 sg13g2_nand3_1 _959_ (.B(_248_),
    .C(_415_),
    .A(_240_),
    .Y(_416_));
 sg13g2_nor3_1 _960_ (.A(_413_),
    .B(_414_),
    .C(_416_),
    .Y(_418_));
 sg13g2_nor4_1 _961_ (.A(_271_),
    .B(_367_),
    .C(_405_),
    .D(_411_),
    .Y(_419_));
 sg13g2_nand4_1 _962_ (.B(_176_),
    .C(_418_),
    .A(net292),
    .Y(_420_),
    .D(_419_));
 sg13g2_nand2_1 _963_ (.Y(_421_),
    .A(_214_),
    .B(_410_));
 sg13g2_nor4_1 _964_ (.A(_093_),
    .B(_114_),
    .C(_168_),
    .D(_279_),
    .Y(_422_));
 sg13g2_nor4_1 _965_ (.A(_105_),
    .B(_109_),
    .C(_382_),
    .D(_421_),
    .Y(_423_));
 sg13g2_nand4_1 _966_ (.B(_201_),
    .C(_422_),
    .A(_195_),
    .Y(_424_),
    .D(_423_));
 sg13g2_a21o_1 _967_ (.A2(_424_),
    .A1(_420_),
    .B1(net8),
    .X(_425_));
 sg13g2_o21ai_1 _968_ (.B1(net289),
    .Y(_426_),
    .A1(_401_),
    .A2(_403_));
 sg13g2_nand3_1 _969_ (.B(_425_),
    .C(_426_),
    .A(net6),
    .Y(_427_));
 sg13g2_xor2_1 _970_ (.B(_427_),
    .A(net294),
    .X(uo_out[0]));
 sg13g2_nand2_1 _971_ (.Y(_429_),
    .A(net297),
    .B(_451_));
 sg13g2_o21ai_1 _972_ (.B1(net6),
    .Y(_430_),
    .A1(_219_),
    .A2(_429_));
 sg13g2_xor2_1 _973_ (.B(_430_),
    .A(net293),
    .X(_431_));
 sg13g2_a21oi_1 _974_ (.A1(net7),
    .A2(_134_),
    .Y(_432_),
    .B1(_245_));
 sg13g2_o21ai_1 _975_ (.B1(_432_),
    .Y(_433_),
    .A1(net291),
    .A2(_431_));
 sg13g2_inv_1 _976_ (.Y(uio_out[1]),
    .A(_433_));
 sg13g2_nand3_1 _977_ (.B(net282),
    .C(_472_),
    .A(net312),
    .Y(_434_));
 sg13g2_nand3_1 _978_ (.B(_303_),
    .C(_434_),
    .A(_138_),
    .Y(_435_));
 sg13g2_a21oi_1 _979_ (.A1(_135_),
    .A2(_435_),
    .Y(_436_),
    .B1(_132_));
 sg13g2_a221oi_1 _980_ (.B2(net317),
    .C1(_128_),
    .B1(net265),
    .A1(net322),
    .Y(_438_),
    .A2(net318));
 sg13g2_or3_1 _981_ (.A(_213_),
    .B(_436_),
    .C(_438_),
    .X(_439_));
 sg13g2_o21ai_1 _982_ (.B1(net290),
    .Y(_440_),
    .A1(net293),
    .A2(_439_));
 sg13g2_a21oi_2 _983_ (.B1(_440_),
    .Y(uio_out[0]),
    .A2(_439_),
    .A1(net293));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_10 (.L_LO(net10));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_11 (.L_LO(net11));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_12 (.L_LO(net12));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_13 (.L_LO(net13));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_14 (.L_LO(net14));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_15 (.L_LO(net15));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_16 (.L_LO(net16));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_17 (.L_LO(net17));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_18 (.L_LO(net18));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_19 (.L_LO(net19));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_20 (.L_LO(net20));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_buf_1 _996_ (.A(net290),
    .X(uio_oe[0]));
 sg13g2_buf_1 _997_ (.A(net290),
    .X(uio_oe[1]));
 sg13g2_buf_4 fanout246 (.X(net246),
    .A(_057_));
 sg13g2_buf_4 fanout247 (.X(net247),
    .A(_028_));
 sg13g2_buf_1 fanout248 (.A(_028_),
    .X(net248));
 sg13g2_buf_4 fanout249 (.X(net249),
    .A(_480_));
 sg13g2_buf_1 fanout250 (.A(_480_),
    .X(net250));
 sg13g2_buf_4 fanout251 (.X(net251),
    .A(_471_));
 sg13g2_buf_1 fanout252 (.A(_471_),
    .X(net252));
 sg13g2_buf_4 fanout253 (.X(net253),
    .A(_007_));
 sg13g2_buf_4 fanout254 (.X(net254),
    .A(_006_));
 sg13g2_buf_4 fanout255 (.X(net255),
    .A(_481_));
 sg13g2_buf_2 fanout256 (.A(_481_),
    .X(net256));
 sg13g2_buf_4 fanout257 (.X(net257),
    .A(_479_));
 sg13g2_buf_2 fanout258 (.A(_479_),
    .X(net258));
 sg13g2_buf_4 fanout259 (.X(net259),
    .A(net262));
 sg13g2_buf_2 fanout260 (.A(net262),
    .X(net260));
 sg13g2_buf_4 fanout261 (.X(net261),
    .A(net262));
 sg13g2_buf_2 fanout262 (.A(_473_),
    .X(net262));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(net266));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(net266));
 sg13g2_buf_2 fanout265 (.A(net266),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_463_),
    .X(net266));
 sg13g2_buf_4 fanout267 (.X(net267),
    .A(_459_));
 sg13g2_buf_2 fanout268 (.A(_459_),
    .X(net268));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(net271));
 sg13g2_buf_4 fanout270 (.X(net270),
    .A(net271));
 sg13g2_buf_4 fanout271 (.X(net271),
    .A(_458_));
 sg13g2_buf_4 fanout272 (.X(net272),
    .A(_455_));
 sg13g2_buf_2 fanout273 (.A(_455_),
    .X(net273));
 sg13g2_buf_4 fanout274 (.X(net274),
    .A(net275));
 sg13g2_buf_4 fanout275 (.X(net275),
    .A(_452_));
 sg13g2_buf_4 fanout276 (.X(net276),
    .A(_446_));
 sg13g2_buf_2 fanout277 (.A(_446_),
    .X(net277));
 sg13g2_buf_4 fanout278 (.X(net278),
    .A(_396_));
 sg13g2_buf_4 fanout279 (.X(net279),
    .A(_299_));
 sg13g2_buf_2 fanout280 (.A(_299_),
    .X(net280));
 sg13g2_buf_4 fanout281 (.X(net281),
    .A(net283));
 sg13g2_buf_2 fanout282 (.A(net283),
    .X(net282));
 sg13g2_buf_4 fanout283 (.X(net283),
    .A(_277_));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(_224_));
 sg13g2_buf_2 fanout285 (.A(net286),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_202_),
    .X(net286));
 sg13g2_buf_4 fanout287 (.X(net287),
    .A(_169_));
 sg13g2_buf_2 fanout288 (.A(_169_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(net290),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(net8),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(net292),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(net7),
    .X(net292));
 sg13g2_buf_4 fanout293 (.X(net293),
    .A(net294));
 sg13g2_buf_2 fanout294 (.A(uio_in[5]),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(net296),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(uio_in[3]),
    .X(net296));
 sg13g2_buf_4 fanout297 (.X(net297),
    .A(uio_in[3]));
 sg13g2_buf_2 fanout298 (.A(net301),
    .X(net298));
 sg13g2_buf_1 fanout299 (.A(net301),
    .X(net299));
 sg13g2_buf_4 fanout300 (.X(net300),
    .A(net301));
 sg13g2_buf_1 fanout301 (.A(ui_in[7]),
    .X(net301));
 sg13g2_buf_4 fanout302 (.X(net302),
    .A(net303));
 sg13g2_buf_4 fanout303 (.X(net303),
    .A(net2));
 sg13g2_buf_2 fanout304 (.A(net306),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(net306),
    .X(net305));
 sg13g2_buf_4 fanout306 (.X(net306),
    .A(ui_in[5]));
 sg13g2_buf_4 fanout307 (.X(net307),
    .A(ui_in[5]));
 sg13g2_buf_2 fanout308 (.A(ui_in[5]),
    .X(net308));
 sg13g2_buf_4 fanout309 (.X(net309),
    .A(net310));
 sg13g2_buf_4 fanout310 (.X(net310),
    .A(ui_in[4]));
 sg13g2_buf_2 fanout311 (.A(net314),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(net313),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(net314),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(ui_in[4]),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(ui_in[3]),
    .X(net315));
 sg13g2_buf_1 fanout316 (.A(net317),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(ui_in[3]),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(net319),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(net1),
    .X(net319));
 sg13g2_buf_4 fanout320 (.X(net320),
    .A(ui_in[1]));
 sg13g2_buf_1 fanout321 (.A(ui_in[1]),
    .X(net321));
 sg13g2_buf_4 fanout322 (.X(net322),
    .A(net324));
 sg13g2_buf_1 fanout323 (.A(net324),
    .X(net323));
 sg13g2_buf_4 fanout324 (.X(net324),
    .A(ui_in[1]));
 sg13g2_buf_4 fanout325 (.X(net325),
    .A(ui_in[0]));
 sg13g2_buf_2 fanout326 (.A(ui_in[0]),
    .X(net326));
 sg13g2_buf_1 input1 (.A(ui_in[2]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[6]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(uio_in[0]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[1]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[2]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(uio_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_rebeccargb_universal_decoder_9 (.L_LO(net9));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_4 FILLER_19_259 ();
 sg13g2_fill_1 FILLER_19_263 ();
 sg13g2_decap_8 FILLER_19_269 ();
 sg13g2_decap_8 FILLER_19_276 ();
 sg13g2_decap_8 FILLER_19_283 ();
 sg13g2_decap_4 FILLER_19_290 ();
 sg13g2_fill_1 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_299 ();
 sg13g2_decap_8 FILLER_19_306 ();
 sg13g2_decap_8 FILLER_19_313 ();
 sg13g2_decap_8 FILLER_19_320 ();
 sg13g2_decap_8 FILLER_19_327 ();
 sg13g2_decap_8 FILLER_19_334 ();
 sg13g2_decap_8 FILLER_19_341 ();
 sg13g2_decap_8 FILLER_19_348 ();
 sg13g2_decap_8 FILLER_19_355 ();
 sg13g2_decap_8 FILLER_19_362 ();
 sg13g2_decap_8 FILLER_19_369 ();
 sg13g2_decap_8 FILLER_19_376 ();
 sg13g2_decap_8 FILLER_19_383 ();
 sg13g2_decap_8 FILLER_19_390 ();
 sg13g2_decap_8 FILLER_19_397 ();
 sg13g2_decap_4 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_fill_2 FILLER_20_189 ();
 sg13g2_fill_1 FILLER_20_191 ();
 sg13g2_decap_8 FILLER_20_201 ();
 sg13g2_fill_2 FILLER_20_208 ();
 sg13g2_fill_1 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_220 ();
 sg13g2_decap_8 FILLER_20_227 ();
 sg13g2_decap_8 FILLER_20_247 ();
 sg13g2_fill_1 FILLER_20_254 ();
 sg13g2_decap_8 FILLER_20_275 ();
 sg13g2_decap_4 FILLER_20_282 ();
 sg13g2_fill_1 FILLER_20_286 ();
 sg13g2_fill_2 FILLER_20_295 ();
 sg13g2_decap_8 FILLER_20_305 ();
 sg13g2_decap_4 FILLER_20_312 ();
 sg13g2_decap_4 FILLER_20_328 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_fill_2 FILLER_20_347 ();
 sg13g2_fill_1 FILLER_20_349 ();
 sg13g2_decap_8 FILLER_20_362 ();
 sg13g2_decap_4 FILLER_20_369 ();
 sg13g2_fill_1 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_fill_1 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_181 ();
 sg13g2_decap_4 FILLER_21_188 ();
 sg13g2_fill_1 FILLER_21_192 ();
 sg13g2_decap_4 FILLER_21_202 ();
 sg13g2_fill_2 FILLER_21_235 ();
 sg13g2_fill_1 FILLER_21_243 ();
 sg13g2_decap_4 FILLER_21_255 ();
 sg13g2_fill_2 FILLER_21_277 ();
 sg13g2_fill_2 FILLER_21_312 ();
 sg13g2_fill_1 FILLER_21_314 ();
 sg13g2_decap_4 FILLER_21_340 ();
 sg13g2_fill_2 FILLER_21_367 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_fill_2 FILLER_22_168 ();
 sg13g2_fill_1 FILLER_22_170 ();
 sg13g2_fill_2 FILLER_22_179 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_fill_2 FILLER_22_203 ();
 sg13g2_decap_4 FILLER_22_224 ();
 sg13g2_fill_2 FILLER_22_228 ();
 sg13g2_fill_1 FILLER_22_235 ();
 sg13g2_fill_2 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_276 ();
 sg13g2_fill_2 FILLER_22_283 ();
 sg13g2_fill_2 FILLER_22_290 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_fill_2 FILLER_22_322 ();
 sg13g2_fill_1 FILLER_22_329 ();
 sg13g2_fill_2 FILLER_22_344 ();
 sg13g2_fill_1 FILLER_22_346 ();
 sg13g2_decap_4 FILLER_22_375 ();
 sg13g2_decap_8 FILLER_22_387 ();
 sg13g2_decap_8 FILLER_22_394 ();
 sg13g2_decap_8 FILLER_22_401 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_4 FILLER_23_161 ();
 sg13g2_fill_1 FILLER_23_165 ();
 sg13g2_fill_2 FILLER_23_177 ();
 sg13g2_fill_1 FILLER_23_179 ();
 sg13g2_fill_2 FILLER_23_185 ();
 sg13g2_fill_1 FILLER_23_187 ();
 sg13g2_fill_1 FILLER_23_209 ();
 sg13g2_fill_2 FILLER_23_229 ();
 sg13g2_fill_2 FILLER_23_262 ();
 sg13g2_fill_1 FILLER_23_264 ();
 sg13g2_fill_2 FILLER_23_269 ();
 sg13g2_fill_1 FILLER_23_271 ();
 sg13g2_decap_4 FILLER_23_293 ();
 sg13g2_fill_1 FILLER_23_312 ();
 sg13g2_fill_1 FILLER_23_323 ();
 sg13g2_decap_8 FILLER_23_340 ();
 sg13g2_fill_1 FILLER_23_352 ();
 sg13g2_decap_8 FILLER_23_367 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_4 FILLER_24_161 ();
 sg13g2_fill_2 FILLER_24_170 ();
 sg13g2_fill_1 FILLER_24_172 ();
 sg13g2_fill_1 FILLER_24_184 ();
 sg13g2_decap_4 FILLER_24_204 ();
 sg13g2_fill_1 FILLER_24_208 ();
 sg13g2_fill_2 FILLER_24_225 ();
 sg13g2_decap_4 FILLER_24_239 ();
 sg13g2_fill_2 FILLER_24_243 ();
 sg13g2_fill_2 FILLER_24_255 ();
 sg13g2_decap_8 FILLER_24_272 ();
 sg13g2_decap_4 FILLER_24_279 ();
 sg13g2_fill_1 FILLER_24_283 ();
 sg13g2_fill_2 FILLER_24_295 ();
 sg13g2_fill_2 FILLER_24_316 ();
 sg13g2_fill_1 FILLER_24_318 ();
 sg13g2_decap_4 FILLER_24_367 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_decap_4 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_4 FILLER_24_403 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_4 FILLER_25_147 ();
 sg13g2_fill_1 FILLER_25_151 ();
 sg13g2_decap_4 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_185 ();
 sg13g2_decap_4 FILLER_25_192 ();
 sg13g2_fill_2 FILLER_25_196 ();
 sg13g2_fill_1 FILLER_25_212 ();
 sg13g2_fill_2 FILLER_25_221 ();
 sg13g2_fill_1 FILLER_25_223 ();
 sg13g2_fill_1 FILLER_25_229 ();
 sg13g2_fill_1 FILLER_25_249 ();
 sg13g2_fill_2 FILLER_25_266 ();
 sg13g2_fill_1 FILLER_25_302 ();
 sg13g2_decap_8 FILLER_25_307 ();
 sg13g2_fill_1 FILLER_25_314 ();
 sg13g2_fill_1 FILLER_25_332 ();
 sg13g2_fill_2 FILLER_25_338 ();
 sg13g2_fill_2 FILLER_25_344 ();
 sg13g2_fill_2 FILLER_25_351 ();
 sg13g2_fill_1 FILLER_25_353 ();
 sg13g2_fill_2 FILLER_25_359 ();
 sg13g2_fill_2 FILLER_25_367 ();
 sg13g2_fill_2 FILLER_25_392 ();
 sg13g2_fill_1 FILLER_25_394 ();
 sg13g2_decap_4 FILLER_25_403 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_4 FILLER_26_154 ();
 sg13g2_fill_1 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_174 ();
 sg13g2_fill_2 FILLER_26_193 ();
 sg13g2_decap_4 FILLER_26_224 ();
 sg13g2_fill_1 FILLER_26_228 ();
 sg13g2_fill_2 FILLER_26_247 ();
 sg13g2_fill_1 FILLER_26_249 ();
 sg13g2_decap_8 FILLER_26_260 ();
 sg13g2_decap_4 FILLER_26_273 ();
 sg13g2_fill_1 FILLER_26_277 ();
 sg13g2_fill_2 FILLER_26_297 ();
 sg13g2_fill_2 FILLER_26_307 ();
 sg13g2_fill_1 FILLER_26_309 ();
 sg13g2_decap_4 FILLER_26_330 ();
 sg13g2_decap_4 FILLER_26_358 ();
 sg13g2_decap_8 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_4 FILLER_27_162 ();
 sg13g2_fill_2 FILLER_27_190 ();
 sg13g2_fill_2 FILLER_27_203 ();
 sg13g2_fill_1 FILLER_27_220 ();
 sg13g2_fill_1 FILLER_27_226 ();
 sg13g2_fill_1 FILLER_27_232 ();
 sg13g2_decap_8 FILLER_27_241 ();
 sg13g2_decap_4 FILLER_27_248 ();
 sg13g2_fill_2 FILLER_27_257 ();
 sg13g2_fill_1 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_269 ();
 sg13g2_fill_2 FILLER_27_297 ();
 sg13g2_fill_1 FILLER_27_311 ();
 sg13g2_decap_8 FILLER_27_323 ();
 sg13g2_fill_2 FILLER_27_330 ();
 sg13g2_fill_2 FILLER_27_341 ();
 sg13g2_fill_1 FILLER_27_343 ();
 sg13g2_fill_2 FILLER_27_350 ();
 sg13g2_fill_2 FILLER_27_359 ();
 sg13g2_fill_1 FILLER_27_361 ();
 sg13g2_decap_8 FILLER_27_382 ();
 sg13g2_fill_2 FILLER_27_389 ();
 sg13g2_fill_1 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_fill_1 FILLER_28_177 ();
 sg13g2_fill_2 FILLER_28_186 ();
 sg13g2_fill_1 FILLER_28_188 ();
 sg13g2_decap_8 FILLER_28_194 ();
 sg13g2_decap_8 FILLER_28_201 ();
 sg13g2_fill_2 FILLER_28_220 ();
 sg13g2_fill_2 FILLER_28_267 ();
 sg13g2_fill_1 FILLER_28_275 ();
 sg13g2_fill_2 FILLER_28_303 ();
 sg13g2_fill_2 FILLER_28_320 ();
 sg13g2_fill_1 FILLER_28_322 ();
 sg13g2_fill_2 FILLER_28_341 ();
 sg13g2_fill_1 FILLER_28_367 ();
 sg13g2_fill_2 FILLER_28_380 ();
 sg13g2_fill_1 FILLER_28_382 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_4 FILLER_29_154 ();
 sg13g2_fill_2 FILLER_29_158 ();
 sg13g2_decap_8 FILLER_29_173 ();
 sg13g2_fill_2 FILLER_29_191 ();
 sg13g2_fill_2 FILLER_29_199 ();
 sg13g2_fill_1 FILLER_29_206 ();
 sg13g2_decap_8 FILLER_29_211 ();
 sg13g2_fill_1 FILLER_29_218 ();
 sg13g2_fill_1 FILLER_29_223 ();
 sg13g2_fill_2 FILLER_29_233 ();
 sg13g2_fill_1 FILLER_29_241 ();
 sg13g2_decap_8 FILLER_29_270 ();
 sg13g2_decap_4 FILLER_29_277 ();
 sg13g2_fill_1 FILLER_29_285 ();
 sg13g2_fill_2 FILLER_29_297 ();
 sg13g2_fill_1 FILLER_29_319 ();
 sg13g2_decap_8 FILLER_29_325 ();
 sg13g2_decap_8 FILLER_29_355 ();
 sg13g2_fill_2 FILLER_29_362 ();
 sg13g2_fill_1 FILLER_29_364 ();
 sg13g2_decap_4 FILLER_29_372 ();
 sg13g2_fill_2 FILLER_29_376 ();
 sg13g2_decap_8 FILLER_29_395 ();
 sg13g2_decap_8 FILLER_29_402 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_fill_2 FILLER_30_147 ();
 sg13g2_fill_1 FILLER_30_149 ();
 sg13g2_fill_1 FILLER_30_170 ();
 sg13g2_fill_1 FILLER_30_182 ();
 sg13g2_fill_1 FILLER_30_189 ();
 sg13g2_fill_2 FILLER_30_210 ();
 sg13g2_fill_1 FILLER_30_212 ();
 sg13g2_fill_1 FILLER_30_229 ();
 sg13g2_fill_2 FILLER_30_248 ();
 sg13g2_fill_2 FILLER_30_256 ();
 sg13g2_fill_1 FILLER_30_258 ();
 sg13g2_decap_4 FILLER_30_298 ();
 sg13g2_decap_4 FILLER_30_311 ();
 sg13g2_fill_2 FILLER_30_315 ();
 sg13g2_fill_1 FILLER_30_327 ();
 sg13g2_fill_2 FILLER_30_342 ();
 sg13g2_fill_1 FILLER_30_344 ();
 sg13g2_fill_1 FILLER_30_359 ();
 sg13g2_decap_4 FILLER_30_373 ();
 sg13g2_fill_1 FILLER_30_377 ();
 sg13g2_decap_8 FILLER_30_383 ();
 sg13g2_fill_2 FILLER_30_390 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_4 FILLER_31_147 ();
 sg13g2_fill_2 FILLER_31_151 ();
 sg13g2_fill_2 FILLER_31_161 ();
 sg13g2_fill_2 FILLER_31_167 ();
 sg13g2_fill_1 FILLER_31_169 ();
 sg13g2_fill_2 FILLER_31_177 ();
 sg13g2_decap_4 FILLER_31_190 ();
 sg13g2_fill_1 FILLER_31_213 ();
 sg13g2_fill_1 FILLER_31_233 ();
 sg13g2_fill_1 FILLER_31_252 ();
 sg13g2_decap_8 FILLER_31_257 ();
 sg13g2_fill_2 FILLER_31_264 ();
 sg13g2_fill_1 FILLER_31_266 ();
 sg13g2_fill_2 FILLER_31_272 ();
 sg13g2_fill_1 FILLER_31_274 ();
 sg13g2_fill_1 FILLER_31_287 ();
 sg13g2_fill_2 FILLER_31_296 ();
 sg13g2_decap_4 FILLER_31_304 ();
 sg13g2_fill_1 FILLER_31_308 ();
 sg13g2_decap_8 FILLER_31_313 ();
 sg13g2_decap_8 FILLER_31_350 ();
 sg13g2_decap_8 FILLER_31_367 ();
 sg13g2_fill_1 FILLER_31_374 ();
 sg13g2_fill_2 FILLER_31_388 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_fill_1 FILLER_32_154 ();
 sg13g2_fill_2 FILLER_32_172 ();
 sg13g2_fill_1 FILLER_32_174 ();
 sg13g2_fill_1 FILLER_32_188 ();
 sg13g2_fill_2 FILLER_32_193 ();
 sg13g2_fill_1 FILLER_32_195 ();
 sg13g2_decap_8 FILLER_32_200 ();
 sg13g2_fill_2 FILLER_32_207 ();
 sg13g2_fill_1 FILLER_32_214 ();
 sg13g2_decap_8 FILLER_32_221 ();
 sg13g2_decap_8 FILLER_32_228 ();
 sg13g2_fill_2 FILLER_32_235 ();
 sg13g2_decap_8 FILLER_32_241 ();
 sg13g2_fill_1 FILLER_32_248 ();
 sg13g2_fill_2 FILLER_32_265 ();
 sg13g2_decap_8 FILLER_32_280 ();
 sg13g2_decap_4 FILLER_32_287 ();
 sg13g2_decap_4 FILLER_32_308 ();
 sg13g2_fill_2 FILLER_32_312 ();
 sg13g2_fill_2 FILLER_32_330 ();
 sg13g2_fill_2 FILLER_32_340 ();
 sg13g2_fill_1 FILLER_32_342 ();
 sg13g2_fill_1 FILLER_32_355 ();
 sg13g2_decap_8 FILLER_32_367 ();
 sg13g2_fill_1 FILLER_32_374 ();
 sg13g2_decap_4 FILLER_32_392 ();
 sg13g2_fill_2 FILLER_32_396 ();
 sg13g2_decap_4 FILLER_32_403 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_fill_2 FILLER_33_147 ();
 sg13g2_fill_2 FILLER_33_163 ();
 sg13g2_fill_1 FILLER_33_165 ();
 sg13g2_fill_1 FILLER_33_172 ();
 sg13g2_fill_2 FILLER_33_178 ();
 sg13g2_fill_1 FILLER_33_180 ();
 sg13g2_fill_1 FILLER_33_186 ();
 sg13g2_fill_2 FILLER_33_210 ();
 sg13g2_fill_1 FILLER_33_224 ();
 sg13g2_decap_4 FILLER_33_244 ();
 sg13g2_decap_4 FILLER_33_260 ();
 sg13g2_fill_1 FILLER_33_264 ();
 sg13g2_fill_1 FILLER_33_281 ();
 sg13g2_decap_4 FILLER_33_286 ();
 sg13g2_fill_2 FILLER_33_321 ();
 sg13g2_fill_1 FILLER_33_323 ();
 sg13g2_fill_1 FILLER_33_328 ();
 sg13g2_decap_4 FILLER_33_334 ();
 sg13g2_decap_4 FILLER_33_343 ();
 sg13g2_fill_1 FILLER_33_347 ();
 sg13g2_decap_4 FILLER_33_358 ();
 sg13g2_fill_2 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_4 FILLER_34_147 ();
 sg13g2_fill_2 FILLER_34_151 ();
 sg13g2_fill_1 FILLER_34_180 ();
 sg13g2_decap_4 FILLER_34_199 ();
 sg13g2_fill_2 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_220 ();
 sg13g2_decap_4 FILLER_34_227 ();
 sg13g2_fill_2 FILLER_34_231 ();
 sg13g2_fill_1 FILLER_34_247 ();
 sg13g2_decap_8 FILLER_34_253 ();
 sg13g2_fill_2 FILLER_34_260 ();
 sg13g2_fill_1 FILLER_34_262 ();
 sg13g2_fill_1 FILLER_34_268 ();
 sg13g2_decap_4 FILLER_34_289 ();
 sg13g2_fill_1 FILLER_34_293 ();
 sg13g2_decap_8 FILLER_34_305 ();
 sg13g2_fill_2 FILLER_34_312 ();
 sg13g2_fill_1 FILLER_34_314 ();
 sg13g2_fill_1 FILLER_34_324 ();
 sg13g2_fill_1 FILLER_34_336 ();
 sg13g2_fill_2 FILLER_34_346 ();
 sg13g2_fill_2 FILLER_34_353 ();
 sg13g2_fill_1 FILLER_34_355 ();
 sg13g2_decap_4 FILLER_34_373 ();
 sg13g2_fill_1 FILLER_34_377 ();
 sg13g2_decap_8 FILLER_34_383 ();
 sg13g2_decap_8 FILLER_34_390 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_fill_2 FILLER_35_161 ();
 sg13g2_fill_1 FILLER_35_181 ();
 sg13g2_fill_2 FILLER_35_200 ();
 sg13g2_fill_1 FILLER_35_216 ();
 sg13g2_fill_2 FILLER_35_222 ();
 sg13g2_fill_1 FILLER_35_229 ();
 sg13g2_fill_2 FILLER_35_245 ();
 sg13g2_decap_4 FILLER_35_294 ();
 sg13g2_fill_2 FILLER_35_312 ();
 sg13g2_fill_1 FILLER_35_314 ();
 sg13g2_fill_1 FILLER_35_338 ();
 sg13g2_fill_1 FILLER_35_345 ();
 sg13g2_fill_2 FILLER_35_380 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_4 FILLER_36_161 ();
 sg13g2_fill_2 FILLER_36_165 ();
 sg13g2_decap_8 FILLER_36_191 ();
 sg13g2_fill_2 FILLER_36_198 ();
 sg13g2_fill_1 FILLER_36_208 ();
 sg13g2_decap_4 FILLER_36_222 ();
 sg13g2_fill_1 FILLER_36_226 ();
 sg13g2_fill_2 FILLER_36_258 ();
 sg13g2_fill_1 FILLER_36_260 ();
 sg13g2_fill_2 FILLER_36_270 ();
 sg13g2_fill_2 FILLER_36_289 ();
 sg13g2_fill_1 FILLER_36_291 ();
 sg13g2_fill_1 FILLER_36_318 ();
 sg13g2_fill_2 FILLER_36_324 ();
 sg13g2_fill_1 FILLER_36_326 ();
 sg13g2_decap_4 FILLER_36_336 ();
 sg13g2_fill_1 FILLER_36_340 ();
 sg13g2_fill_1 FILLER_36_355 ();
 sg13g2_fill_1 FILLER_36_361 ();
 sg13g2_decap_8 FILLER_36_372 ();
 sg13g2_decap_8 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_36_386 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_4 FILLER_37_168 ();
 sg13g2_fill_1 FILLER_37_172 ();
 sg13g2_fill_2 FILLER_37_182 ();
 sg13g2_fill_1 FILLER_37_184 ();
 sg13g2_decap_8 FILLER_37_197 ();
 sg13g2_fill_2 FILLER_37_204 ();
 sg13g2_fill_1 FILLER_37_206 ();
 sg13g2_decap_8 FILLER_37_215 ();
 sg13g2_fill_1 FILLER_37_230 ();
 sg13g2_decap_8 FILLER_37_239 ();
 sg13g2_fill_2 FILLER_37_256 ();
 sg13g2_fill_2 FILLER_37_268 ();
 sg13g2_fill_1 FILLER_37_287 ();
 sg13g2_fill_1 FILLER_37_308 ();
 sg13g2_fill_2 FILLER_37_338 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_8 FILLER_38_100 ();
 sg13g2_decap_8 FILLER_38_107 ();
 sg13g2_decap_4 FILLER_38_114 ();
 sg13g2_fill_2 FILLER_38_118 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_8 FILLER_38_164 ();
 sg13g2_decap_8 FILLER_38_171 ();
 sg13g2_decap_8 FILLER_38_178 ();
 sg13g2_decap_8 FILLER_38_185 ();
 sg13g2_decap_8 FILLER_38_192 ();
 sg13g2_decap_4 FILLER_38_199 ();
 sg13g2_fill_2 FILLER_38_224 ();
 sg13g2_decap_4 FILLER_38_231 ();
 sg13g2_fill_2 FILLER_38_235 ();
 sg13g2_fill_2 FILLER_38_286 ();
 sg13g2_decap_4 FILLER_38_292 ();
 sg13g2_fill_2 FILLER_38_296 ();
 sg13g2_decap_8 FILLER_38_310 ();
 sg13g2_decap_8 FILLER_38_336 ();
 sg13g2_fill_2 FILLER_38_343 ();
 sg13g2_fill_1 FILLER_38_345 ();
 sg13g2_decap_8 FILLER_38_358 ();
 sg13g2_decap_8 FILLER_38_365 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[2] = net9;
 assign uio_oe[3] = net10;
 assign uio_oe[4] = net11;
 assign uio_oe[5] = net12;
 assign uio_oe[6] = net13;
 assign uio_oe[7] = net14;
 assign uio_out[2] = net15;
 assign uio_out[3] = net16;
 assign uio_out[4] = net17;
 assign uio_out[5] = net18;
 assign uio_out[6] = net19;
 assign uio_out[7] = net20;
endmodule

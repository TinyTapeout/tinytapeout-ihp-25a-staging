module tt_um_johshoff_metaballs (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire clknet_0_clk;
 wire h_sync;
 wire \mb.b_0.ball_vx[0] ;
 wire \mb.b_0.ball_vx[1] ;
 wire \mb.b_0.ball_vx[2] ;
 wire \mb.b_0.ball_vx[3] ;
 wire \mb.b_0.ball_vx[4] ;
 wire \mb.b_0.ball_vx[5] ;
 wire \mb.b_0.ball_vx[6] ;
 wire \mb.b_0.ball_vx[7] ;
 wire \mb.b_0.ball_vx[8] ;
 wire \mb.b_0.ball_vx[9] ;
 wire \mb.b_0.ball_vy[0] ;
 wire \mb.b_0.ball_vy[1] ;
 wire \mb.b_0.ball_vy[2] ;
 wire \mb.b_0.ball_vy[3] ;
 wire \mb.b_0.ball_vy[4] ;
 wire \mb.b_0.ball_vy[5] ;
 wire \mb.b_0.ball_vy[6] ;
 wire \mb.b_0.ball_vy[7] ;
 wire \mb.b_0.ball_vy[8] ;
 wire \mb.b_0.ball_vy[9] ;
 wire \mb.b_0.ball_x[0] ;
 wire \mb.b_0.ball_x[1] ;
 wire \mb.b_0.ball_x[2] ;
 wire \mb.b_0.ball_x[3] ;
 wire \mb.b_0.ball_x[4] ;
 wire \mb.b_0.ball_x[5] ;
 wire \mb.b_0.ball_x[6] ;
 wire \mb.b_0.ball_x[7] ;
 wire \mb.b_0.ball_x[8] ;
 wire \mb.b_0.ball_x[9] ;
 wire \mb.b_0.ball_y[0] ;
 wire \mb.b_0.ball_y[1] ;
 wire \mb.b_0.ball_y[2] ;
 wire \mb.b_0.ball_y[3] ;
 wire \mb.b_0.ball_y[4] ;
 wire \mb.b_0.ball_y[5] ;
 wire \mb.b_0.ball_y[6] ;
 wire \mb.b_0.ball_y[7] ;
 wire \mb.b_0.ball_y[8] ;
 wire \mb.b_0.ball_y[9] ;
 wire \mb.b_0.next_x[0] ;
 wire \mb.b_0.next_x[1] ;
 wire \mb.b_0.next_x[2] ;
 wire \mb.b_0.next_x[3] ;
 wire \mb.b_0.next_x[4] ;
 wire \mb.b_0.next_x[5] ;
 wire \mb.b_0.next_x[6] ;
 wire \mb.b_0.next_x[7] ;
 wire \mb.b_0.next_x[8] ;
 wire \mb.b_0.next_x[9] ;
 wire \mb.b_0.next_y[0] ;
 wire \mb.b_0.next_y[1] ;
 wire \mb.b_0.next_y[2] ;
 wire \mb.b_0.next_y[3] ;
 wire \mb.b_0.next_y[4] ;
 wire \mb.b_0.next_y[5] ;
 wire \mb.b_0.next_y[6] ;
 wire \mb.b_0.next_y[7] ;
 wire \mb.b_0.next_y[8] ;
 wire \mb.b_0.next_y[9] ;
 wire \mb.b_0.v_sync ;
 wire \mb.b_0.x[0] ;
 wire \mb.b_0.x[1] ;
 wire \mb.b_0.x[2] ;
 wire \mb.b_0.x[3] ;
 wire \mb.b_0.x[4] ;
 wire \mb.b_0.x[5] ;
 wire \mb.b_0.x[6] ;
 wire \mb.b_0.x[7] ;
 wire \mb.b_0.x[8] ;
 wire \mb.b_0.x[9] ;
 wire \mb.b_0.y[0] ;
 wire \mb.b_0.y[1] ;
 wire \mb.b_0.y[2] ;
 wire \mb.b_0.y[3] ;
 wire \mb.b_0.y[4] ;
 wire \mb.b_0.y[5] ;
 wire \mb.b_0.y[6] ;
 wire \mb.b_0.y[7] ;
 wire \mb.b_0.y[8] ;
 wire \mb.b_0.y[9] ;
 wire \mb.b_1.ball_vx[0] ;
 wire \mb.b_1.ball_vx[1] ;
 wire \mb.b_1.ball_vx[2] ;
 wire \mb.b_1.ball_vx[3] ;
 wire \mb.b_1.ball_vx[4] ;
 wire \mb.b_1.ball_vx[5] ;
 wire \mb.b_1.ball_vx[6] ;
 wire \mb.b_1.ball_vx[7] ;
 wire \mb.b_1.ball_vx[8] ;
 wire \mb.b_1.ball_vx[9] ;
 wire \mb.b_1.ball_vy[0] ;
 wire \mb.b_1.ball_vy[1] ;
 wire \mb.b_1.ball_vy[2] ;
 wire \mb.b_1.ball_vy[3] ;
 wire \mb.b_1.ball_vy[4] ;
 wire \mb.b_1.ball_vy[5] ;
 wire \mb.b_1.ball_vy[6] ;
 wire \mb.b_1.ball_vy[7] ;
 wire \mb.b_1.ball_vy[8] ;
 wire \mb.b_1.ball_vy[9] ;
 wire \mb.b_1.ball_x[0] ;
 wire \mb.b_1.ball_x[1] ;
 wire \mb.b_1.ball_x[2] ;
 wire \mb.b_1.ball_x[3] ;
 wire \mb.b_1.ball_x[4] ;
 wire \mb.b_1.ball_x[5] ;
 wire \mb.b_1.ball_x[6] ;
 wire \mb.b_1.ball_x[7] ;
 wire \mb.b_1.ball_x[8] ;
 wire \mb.b_1.ball_x[9] ;
 wire \mb.b_1.ball_y[0] ;
 wire \mb.b_1.ball_y[1] ;
 wire \mb.b_1.ball_y[2] ;
 wire \mb.b_1.ball_y[3] ;
 wire \mb.b_1.ball_y[4] ;
 wire \mb.b_1.ball_y[5] ;
 wire \mb.b_1.ball_y[6] ;
 wire \mb.b_1.ball_y[7] ;
 wire \mb.b_1.ball_y[8] ;
 wire \mb.b_1.ball_y[9] ;
 wire \mb.b_1.next_x[0] ;
 wire \mb.b_1.next_x[1] ;
 wire \mb.b_1.next_x[2] ;
 wire \mb.b_1.next_x[3] ;
 wire \mb.b_1.next_x[4] ;
 wire \mb.b_1.next_x[5] ;
 wire \mb.b_1.next_x[6] ;
 wire \mb.b_1.next_x[7] ;
 wire \mb.b_1.next_x[8] ;
 wire \mb.b_1.next_x[9] ;
 wire \mb.b_1.next_y[0] ;
 wire \mb.b_1.next_y[1] ;
 wire \mb.b_1.next_y[2] ;
 wire \mb.b_1.next_y[3] ;
 wire \mb.b_1.next_y[4] ;
 wire \mb.b_1.next_y[5] ;
 wire \mb.b_1.next_y[6] ;
 wire \mb.b_1.next_y[7] ;
 wire \mb.b_1.next_y[8] ;
 wire \mb.b_1.next_y[9] ;
 wire \mb.pix ;
 wire \mb.rgb ;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire \v.h_counter[10] ;
 wire \v.h_display ;
 wire \v.v_display ;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net1;
 wire net2;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;

 sg13g2_inv_1 _1278_ (.Y(_0322_),
    .A(\mb.b_0.y[9] ));
 sg13g2_inv_2 _1279_ (.Y(_0323_),
    .A(net149));
 sg13g2_inv_1 _1280_ (.Y(_0324_),
    .A(\mb.b_0.y[7] ));
 sg13g2_inv_1 _1281_ (.Y(_0325_),
    .A(net157));
 sg13g2_inv_1 _1282_ (.Y(_0326_),
    .A(\mb.b_0.y[5] ));
 sg13g2_inv_1 _1283_ (.Y(_0327_),
    .A(net128));
 sg13g2_inv_1 _1284_ (.Y(_0328_),
    .A(net135));
 sg13g2_inv_1 _1285_ (.Y(_0329_),
    .A(\mb.b_0.ball_vx[0] ));
 sg13g2_inv_1 _1286_ (.Y(_0330_),
    .A(\mb.b_0.x[6] ));
 sg13g2_inv_1 _1287_ (.Y(_0331_),
    .A(\mb.b_0.ball_x[3] ));
 sg13g2_inv_1 _1288_ (.Y(_0332_),
    .A(\mb.b_0.ball_y[7] ));
 sg13g2_inv_1 _1289_ (.Y(_0333_),
    .A(\mb.b_0.ball_y[8] ));
 sg13g2_inv_1 _1290_ (.Y(_0334_),
    .A(net324));
 sg13g2_inv_2 _1291_ (.Y(_0335_),
    .A(\mb.b_0.x[9] ));
 sg13g2_inv_1 _1292_ (.Y(_0336_),
    .A(\mb.b_0.x[8] ));
 sg13g2_inv_1 _1293_ (.Y(_0337_),
    .A(\mb.b_1.ball_x[3] ));
 sg13g2_inv_1 _1294_ (.Y(_0338_),
    .A(\mb.b_1.ball_y[7] ));
 sg13g2_inv_1 _1295_ (.Y(_0339_),
    .A(\mb.b_1.ball_y[9] ));
 sg13g2_inv_1 _1296_ (.Y(_0340_),
    .A(\mb.b_1.ball_y[8] ));
 sg13g2_inv_1 _1297_ (.Y(_0341_),
    .A(\mb.b_1.ball_x[9] ));
 sg13g2_inv_1 _1298_ (.Y(_0342_),
    .A(\mb.b_1.ball_x[8] ));
 sg13g2_inv_1 _1299_ (.Y(_0343_),
    .A(\mb.b_1.ball_vx[0] ));
 sg13g2_inv_1 _1300_ (.Y(_0344_),
    .A(\mb.b_1.ball_vx[7] ));
 sg13g2_inv_1 _1301_ (.Y(_0345_),
    .A(\mb.b_0.ball_vx[7] ));
 sg13g2_inv_1 _1302_ (.Y(_0346_),
    .A(\mb.b_0.ball_vx[1] ));
 sg13g2_inv_1 _1303_ (.Y(_0347_),
    .A(\mb.b_1.ball_vx[1] ));
 sg13g2_nand2b_1 _1304_ (.Y(_0348_),
    .B(\mb.b_0.y[6] ),
    .A_N(\mb.b_1.ball_y[6] ));
 sg13g2_xor2_1 _1305_ (.B(\mb.b_1.ball_y[6] ),
    .A(\mb.b_0.y[6] ),
    .X(_0349_));
 sg13g2_nand2_1 _1306_ (.Y(_0350_),
    .A(_0326_),
    .B(\mb.b_1.ball_y[5] ));
 sg13g2_nand2b_1 _1307_ (.Y(_0351_),
    .B(net306),
    .A_N(\mb.b_1.ball_y[4] ));
 sg13g2_nor2b_1 _1308_ (.A(\mb.b_1.ball_y[3] ),
    .B_N(\mb.b_0.y[3] ),
    .Y(_0352_));
 sg13g2_nor2b_1 _1309_ (.A(\mb.b_1.ball_y[2] ),
    .B_N(\mb.b_0.y[2] ),
    .Y(_0353_));
 sg13g2_nand2b_1 _1310_ (.Y(_0354_),
    .B(\mb.b_1.ball_y[2] ),
    .A_N(net308));
 sg13g2_nand2b_1 _1311_ (.Y(_0355_),
    .B(_0354_),
    .A_N(_0353_));
 sg13g2_nor2b_1 _1312_ (.A(net309),
    .B_N(\mb.b_1.ball_y[1] ),
    .Y(_0356_));
 sg13g2_nand2b_1 _1313_ (.Y(_0357_),
    .B(net309),
    .A_N(\mb.b_1.ball_y[1] ));
 sg13g2_nor2b_1 _1314_ (.A(\mb.b_0.y[0] ),
    .B_N(\mb.b_1.ball_y[0] ),
    .Y(_0358_));
 sg13g2_a21oi_2 _1315_ (.B1(_0356_),
    .Y(_0359_),
    .A2(_0358_),
    .A1(_0357_));
 sg13g2_a21o_1 _1316_ (.A2(_0359_),
    .A1(_0354_),
    .B1(_0353_),
    .X(_0360_));
 sg13g2_nand2b_1 _1317_ (.Y(_0361_),
    .B(\mb.b_1.ball_y[3] ),
    .A_N(\mb.b_0.y[3] ));
 sg13g2_nand2b_1 _1318_ (.Y(_0362_),
    .B(_0361_),
    .A_N(_0352_));
 sg13g2_a21oi_1 _1319_ (.A1(_0360_),
    .A2(_0361_),
    .Y(_0363_),
    .B1(_0352_));
 sg13g2_nor2b_1 _1320_ (.A(net306),
    .B_N(\mb.b_1.ball_y[4] ),
    .Y(_0364_));
 sg13g2_xnor2_1 _1321_ (.Y(_0365_),
    .A(net305),
    .B(\mb.b_1.ball_y[4] ));
 sg13g2_o21ai_1 _1322_ (.B1(_0351_),
    .Y(_0366_),
    .A1(_0363_),
    .A2(_0364_));
 sg13g2_nor2_1 _1323_ (.A(_0350_),
    .B(_0366_),
    .Y(_0367_));
 sg13g2_nor2_1 _1324_ (.A(_0326_),
    .B(\mb.b_1.ball_y[5] ),
    .Y(_0368_));
 sg13g2_a21oi_1 _1325_ (.A1(_0366_),
    .A2(_0368_),
    .Y(_0369_),
    .B1(_0367_));
 sg13g2_xnor2_1 _1326_ (.Y(_0370_),
    .A(_0349_),
    .B(_0369_));
 sg13g2_xor2_1 _1327_ (.B(_0369_),
    .A(_0349_),
    .X(_0371_));
 sg13g2_a21oi_2 _1328_ (.B1(_0368_),
    .Y(_0372_),
    .A2(_0366_),
    .A1(_0350_));
 sg13g2_xor2_1 _1329_ (.B(_0372_),
    .A(_0349_),
    .X(_0373_));
 sg13g2_xnor2_1 _1330_ (.Y(_0374_),
    .A(_0349_),
    .B(_0372_));
 sg13g2_xnor2_1 _1331_ (.Y(_0375_),
    .A(_0363_),
    .B(_0365_));
 sg13g2_xnor2_1 _1332_ (.Y(_0376_),
    .A(_0373_),
    .B(_0375_));
 sg13g2_xnor2_1 _1333_ (.Y(_0377_),
    .A(_0374_),
    .B(_0375_));
 sg13g2_xor2_1 _1334_ (.B(\mb.b_1.ball_x[6] ),
    .A(\mb.b_0.x[6] ),
    .X(_0378_));
 sg13g2_nand2b_1 _1335_ (.Y(_0379_),
    .B(\mb.b_1.ball_x[5] ),
    .A_N(\mb.b_0.x[5] ));
 sg13g2_nand2b_1 _1336_ (.Y(_0380_),
    .B(\mb.b_0.x[5] ),
    .A_N(\mb.b_1.ball_x[5] ));
 sg13g2_nor2b_1 _1337_ (.A(\mb.b_1.ball_x[4] ),
    .B_N(net325),
    .Y(_0381_));
 sg13g2_xor2_1 _1338_ (.B(\mb.b_1.ball_x[4] ),
    .A(net325),
    .X(_0382_));
 sg13g2_nor2_1 _1339_ (.A(net326),
    .B(_0337_),
    .Y(_0383_));
 sg13g2_nor2b_1 _1340_ (.A(\mb.b_1.ball_x[2] ),
    .B_N(\mb.b_0.x[2] ),
    .Y(_0384_));
 sg13g2_xnor2_1 _1341_ (.Y(_0385_),
    .A(\mb.b_0.x[2] ),
    .B(\mb.b_1.ball_x[2] ));
 sg13g2_nor2b_1 _1342_ (.A(\mb.b_0.x[1] ),
    .B_N(\mb.b_1.ball_x[1] ),
    .Y(_0386_));
 sg13g2_nand2b_1 _1343_ (.Y(_0387_),
    .B(\mb.b_0.x[1] ),
    .A_N(\mb.b_1.ball_x[1] ));
 sg13g2_nor2b_1 _1344_ (.A(\mb.b_0.x[0] ),
    .B_N(\mb.b_1.ball_x[0] ),
    .Y(_0388_));
 sg13g2_a21oi_2 _1345_ (.B1(_0386_),
    .Y(_0389_),
    .A2(_0388_),
    .A1(_0387_));
 sg13g2_a21oi_1 _1346_ (.A1(_0385_),
    .A2(_0389_),
    .Y(_0390_),
    .B1(_0384_));
 sg13g2_a221oi_1 _1347_ (.B2(_0389_),
    .C1(_0384_),
    .B1(_0385_),
    .A1(net326),
    .Y(_0391_),
    .A2(_0337_));
 sg13g2_nor3_1 _1348_ (.A(_0382_),
    .B(_0383_),
    .C(_0391_),
    .Y(_0392_));
 sg13g2_nor2_1 _1349_ (.A(_0381_),
    .B(_0392_),
    .Y(_0393_));
 sg13g2_o21ai_1 _1350_ (.B1(_0379_),
    .Y(_0394_),
    .A1(_0381_),
    .A2(_0392_));
 sg13g2_a21o_2 _1351_ (.A2(_0394_),
    .A1(_0380_),
    .B1(_0378_),
    .X(_0395_));
 sg13g2_nand3_1 _1352_ (.B(_0380_),
    .C(_0394_),
    .A(_0378_),
    .Y(_0396_));
 sg13g2_nand2_1 _1353_ (.Y(_0397_),
    .A(_0395_),
    .B(_0396_));
 sg13g2_xor2_1 _1354_ (.B(\mb.b_1.ball_x[3] ),
    .A(net326),
    .X(_0398_));
 sg13g2_xnor2_1 _1355_ (.Y(_0399_),
    .A(_0390_),
    .B(_0398_));
 sg13g2_a21o_1 _1356_ (.A2(_0396_),
    .A1(_0395_),
    .B1(_0399_),
    .X(_0400_));
 sg13g2_nand3_1 _1357_ (.B(_0396_),
    .C(_0399_),
    .A(_0395_),
    .Y(_0401_));
 sg13g2_nand2_2 _1358_ (.Y(_0402_),
    .A(_0400_),
    .B(_0401_));
 sg13g2_and2_2 _1359_ (.A(_0400_),
    .B(_0401_),
    .X(_0403_));
 sg13g2_xor2_1 _1360_ (.B(_0389_),
    .A(_0385_),
    .X(_0404_));
 sg13g2_xor2_1 _1361_ (.B(_0404_),
    .A(_0397_),
    .X(_0405_));
 sg13g2_xnor2_1 _1362_ (.Y(_0406_),
    .A(_0397_),
    .B(_0404_));
 sg13g2_nand2_1 _1363_ (.Y(_0407_),
    .A(_0403_),
    .B(net285));
 sg13g2_o21ai_1 _1364_ (.B1(_0382_),
    .Y(_0408_),
    .A1(_0383_),
    .A2(_0391_));
 sg13g2_nand2b_1 _1365_ (.Y(_0409_),
    .B(_0408_),
    .A_N(_0392_));
 sg13g2_a21o_1 _1366_ (.A2(_0396_),
    .A1(_0395_),
    .B1(_0409_),
    .X(_0410_));
 sg13g2_nand3_1 _1367_ (.B(_0396_),
    .C(_0409_),
    .A(_0395_),
    .Y(_0411_));
 sg13g2_and2_1 _1368_ (.A(_0410_),
    .B(_0411_),
    .X(_0412_));
 sg13g2_nand2_1 _1369_ (.Y(_0413_),
    .A(_0410_),
    .B(_0411_));
 sg13g2_nor2_2 _1370_ (.A(_0403_),
    .B(net285),
    .Y(_0414_));
 sg13g2_o21ai_1 _1371_ (.B1(net283),
    .Y(_0415_),
    .A1(_0403_),
    .A2(net285));
 sg13g2_nand2_1 _1372_ (.Y(_0416_),
    .A(_0402_),
    .B(net285));
 sg13g2_xnor2_1 _1373_ (.Y(_0417_),
    .A(_0399_),
    .B(_0404_));
 sg13g2_xor2_1 _1374_ (.B(_0404_),
    .A(_0399_),
    .X(_0418_));
 sg13g2_mux2_1 _1375_ (.A0(_0380_),
    .A1(_0379_),
    .S(_0393_),
    .X(_0419_));
 sg13g2_xor2_1 _1376_ (.B(_0419_),
    .A(_0378_),
    .X(_0420_));
 sg13g2_xnor2_1 _1377_ (.Y(_0421_),
    .A(_0378_),
    .B(_0419_));
 sg13g2_a21oi_1 _1378_ (.A1(net283),
    .A2(_0417_),
    .Y(_0422_),
    .B1(net296));
 sg13g2_nor2_2 _1379_ (.A(_0406_),
    .B(net283),
    .Y(_0423_));
 sg13g2_nand2_1 _1380_ (.Y(_0424_),
    .A(net286),
    .B(_0413_));
 sg13g2_a22oi_1 _1381_ (.Y(_0425_),
    .B1(_0410_),
    .B2(_0411_),
    .A2(_0401_),
    .A1(_0400_));
 sg13g2_nand2_1 _1382_ (.Y(_0426_),
    .A(_0402_),
    .B(net281));
 sg13g2_nand3_1 _1383_ (.B(_0424_),
    .C(net258),
    .A(_0422_),
    .Y(_0427_));
 sg13g2_xnor2_1 _1384_ (.Y(_0428_),
    .A(_0355_),
    .B(_0359_));
 sg13g2_xnor2_1 _1385_ (.Y(_0429_),
    .A(_0373_),
    .B(_0428_));
 sg13g2_xnor2_1 _1386_ (.Y(_0430_),
    .A(_0374_),
    .B(_0428_));
 sg13g2_nor2_2 _1387_ (.A(net284),
    .B(net300),
    .Y(_0431_));
 sg13g2_nand2_2 _1388_ (.Y(_0432_),
    .A(_0402_),
    .B(net283));
 sg13g2_nand2_2 _1389_ (.Y(_0433_),
    .A(net284),
    .B(net281));
 sg13g2_nand2_2 _1390_ (.Y(_0434_),
    .A(net284),
    .B(net283));
 sg13g2_a21oi_2 _1391_ (.B1(net298),
    .Y(_0435_),
    .A2(net282),
    .A1(net284));
 sg13g2_nand2_1 _1392_ (.Y(_0436_),
    .A(_0432_),
    .B(_0435_));
 sg13g2_a21oi_1 _1393_ (.A1(_0431_),
    .A2(_0432_),
    .Y(_0437_),
    .B1(net279));
 sg13g2_xnor2_1 _1394_ (.Y(_0438_),
    .A(_0360_),
    .B(_0362_));
 sg13g2_xnor2_1 _1395_ (.Y(_0439_),
    .A(_0373_),
    .B(_0438_));
 sg13g2_xnor2_1 _1396_ (.Y(_0440_),
    .A(_0374_),
    .B(_0438_));
 sg13g2_nor2_1 _1397_ (.A(net286),
    .B(net258),
    .Y(_0441_));
 sg13g2_o21ai_1 _1398_ (.B1(net279),
    .Y(_0442_),
    .A1(net284),
    .A2(net296));
 sg13g2_o21ai_1 _1399_ (.B1(_0439_),
    .Y(_0443_),
    .A1(_0441_),
    .A2(_0442_));
 sg13g2_a21oi_1 _1400_ (.A1(_0427_),
    .A2(_0437_),
    .Y(_0444_),
    .B1(_0443_));
 sg13g2_nand2_2 _1401_ (.Y(_0445_),
    .A(net279),
    .B(net276));
 sg13g2_inv_1 _1402_ (.Y(_0446_),
    .A(_0445_));
 sg13g2_a21o_1 _1403_ (.A2(_0434_),
    .A1(net258),
    .B1(net296),
    .X(_0447_));
 sg13g2_nor2_1 _1404_ (.A(_0403_),
    .B(net299),
    .Y(_0448_));
 sg13g2_nand2_2 _1405_ (.Y(_0449_),
    .A(_0402_),
    .B(net296));
 sg13g2_o21ai_1 _1406_ (.B1(_0447_),
    .Y(_0450_),
    .A1(_0423_),
    .A2(_0449_));
 sg13g2_nand3_1 _1407_ (.B(net283),
    .C(net300),
    .A(net286),
    .Y(_0451_));
 sg13g2_nand3_1 _1408_ (.B(_0449_),
    .C(_0451_),
    .A(_0433_),
    .Y(_0452_));
 sg13g2_nand2_2 _1409_ (.Y(_0453_),
    .A(net280),
    .B(net276));
 sg13g2_nor2_1 _1410_ (.A(_0441_),
    .B(_0453_),
    .Y(_0454_));
 sg13g2_a221oi_1 _1411_ (.B2(_0454_),
    .C1(_0444_),
    .B1(_0452_),
    .A1(_0446_),
    .Y(_0455_),
    .A2(_0450_));
 sg13g2_nor2_1 _1412_ (.A(net287),
    .B(_0455_),
    .Y(_0456_));
 sg13g2_o21ai_1 _1413_ (.B1(net282),
    .Y(_0457_),
    .A1(_0402_),
    .A2(net285));
 sg13g2_nand2_2 _1414_ (.Y(_0458_),
    .A(net282),
    .B(_0418_));
 sg13g2_nor2_2 _1415_ (.A(net294),
    .B(_0425_),
    .Y(_0459_));
 sg13g2_nand2_1 _1416_ (.Y(_0460_),
    .A(net300),
    .B(_0426_));
 sg13g2_nand2_2 _1417_ (.Y(_0461_),
    .A(_0403_),
    .B(_0423_));
 sg13g2_a221oi_1 _1418_ (.B2(_0435_),
    .C1(net279),
    .B1(_0461_),
    .A1(_0458_),
    .Y(_0462_),
    .A2(_0459_));
 sg13g2_nor2_1 _1419_ (.A(_0402_),
    .B(net282),
    .Y(_0463_));
 sg13g2_nand2_1 _1420_ (.Y(_0464_),
    .A(_0403_),
    .B(net281));
 sg13g2_nand2_1 _1421_ (.Y(_0465_),
    .A(net281),
    .B(_0417_));
 sg13g2_a21oi_1 _1422_ (.A1(_0432_),
    .A2(_0465_),
    .Y(_0466_),
    .B1(net298));
 sg13g2_o21ai_1 _1423_ (.B1(_0458_),
    .Y(_0467_),
    .A1(net282),
    .A2(_0414_));
 sg13g2_or2_1 _1424_ (.X(_0468_),
    .B(_0467_),
    .A(_0466_));
 sg13g2_a21oi_1 _1425_ (.A1(_0466_),
    .A2(_0467_),
    .Y(_0469_),
    .B1(net280));
 sg13g2_a21oi_1 _1426_ (.A1(_0468_),
    .A2(_0469_),
    .Y(_0470_),
    .B1(_0462_));
 sg13g2_nor2_1 _1427_ (.A(_0439_),
    .B(_0470_),
    .Y(_0471_));
 sg13g2_nor2_2 _1428_ (.A(net280),
    .B(net276),
    .Y(_0472_));
 sg13g2_inv_1 _1429_ (.Y(_0473_),
    .A(_0472_));
 sg13g2_a221oi_1 _1430_ (.B2(net298),
    .C1(_0473_),
    .B1(_0457_),
    .A1(_0407_),
    .Y(_0474_),
    .A2(_0435_));
 sg13g2_nor2_1 _1431_ (.A(net279),
    .B(net277),
    .Y(_0475_));
 sg13g2_nor2_2 _1432_ (.A(_0402_),
    .B(net281),
    .Y(_0476_));
 sg13g2_nand2_2 _1433_ (.Y(_0477_),
    .A(_0403_),
    .B(net282));
 sg13g2_nand2_2 _1434_ (.Y(_0478_),
    .A(net285),
    .B(_0476_));
 sg13g2_nand2_1 _1435_ (.Y(_0479_),
    .A(net297),
    .B(_0478_));
 sg13g2_nand3_1 _1436_ (.B(net257),
    .C(_0478_),
    .A(net295),
    .Y(_0480_));
 sg13g2_nand4_1 _1437_ (.B(_0434_),
    .C(_0461_),
    .A(net300),
    .Y(_0481_),
    .D(_0475_));
 sg13g2_nand3_1 _1438_ (.B(_0480_),
    .C(_0481_),
    .A(net287),
    .Y(_0482_));
 sg13g2_nor3_1 _1439_ (.A(_0471_),
    .B(_0474_),
    .C(_0482_),
    .Y(_0483_));
 sg13g2_o21ai_1 _1440_ (.B1(_0370_),
    .Y(_0484_),
    .A1(_0456_),
    .A2(_0483_));
 sg13g2_o21ai_1 _1441_ (.B1(_0395_),
    .Y(_0485_),
    .A1(_0330_),
    .A2(\mb.b_1.ball_x[6] ));
 sg13g2_a21oi_1 _1442_ (.A1(net324),
    .A2(\mb.b_1.ball_x[7] ),
    .Y(_0486_),
    .B1(_0485_));
 sg13g2_nand2_1 _1443_ (.Y(_0487_),
    .A(\mb.b_1.ball_x[7] ),
    .B(\mb.b_1.ball_x[8] ));
 sg13g2_xor2_1 _1444_ (.B(\mb.b_1.ball_x[8] ),
    .A(\mb.b_1.ball_x[7] ),
    .X(_0488_));
 sg13g2_inv_1 _1445_ (.Y(_0489_),
    .A(_0488_));
 sg13g2_xor2_1 _1446_ (.B(_0488_),
    .A(_0041_),
    .X(_0490_));
 sg13g2_o21ai_1 _1447_ (.B1(_0490_),
    .Y(_0491_),
    .A1(net324),
    .A2(\mb.b_1.ball_x[7] ));
 sg13g2_nor2_1 _1448_ (.A(_0486_),
    .B(_0491_),
    .Y(_0492_));
 sg13g2_and2_1 _1449_ (.A(_0043_),
    .B(_0487_),
    .X(_0493_));
 sg13g2_a221oi_1 _1450_ (.B2(\mb.b_0.x[9] ),
    .C1(_0492_),
    .B1(_0493_),
    .A1(\mb.b_0.x[8] ),
    .Y(_0494_),
    .A2(_0489_));
 sg13g2_or2_1 _1451_ (.X(_0495_),
    .B(_0487_),
    .A(_0043_));
 sg13g2_o21ai_1 _1452_ (.B1(_0495_),
    .Y(_0496_),
    .A1(\mb.b_0.x[9] ),
    .A2(_0493_));
 sg13g2_a22oi_1 _1453_ (.Y(_0497_),
    .B1(_0342_),
    .B2(\mb.b_0.x[8] ),
    .A2(_0341_),
    .A1(\mb.b_0.x[9] ));
 sg13g2_nor2_1 _1454_ (.A(_0334_),
    .B(\mb.b_1.ball_x[7] ),
    .Y(_0498_));
 sg13g2_a22oi_1 _1455_ (.Y(_0499_),
    .B1(\mb.b_1.ball_x[8] ),
    .B2(_0336_),
    .A2(\mb.b_1.ball_x[7] ),
    .A1(_0334_));
 sg13g2_o21ai_1 _1456_ (.B1(_0499_),
    .Y(_0500_),
    .A1(_0485_),
    .A2(_0498_));
 sg13g2_a22oi_1 _1457_ (.Y(_0501_),
    .B1(_0497_),
    .B2(_0500_),
    .A2(\mb.b_1.ball_x[9] ),
    .A1(_0335_));
 sg13g2_o21ai_1 _1458_ (.B1(_0501_),
    .Y(_0502_),
    .A1(_0494_),
    .A2(_0496_));
 sg13g2_o21ai_1 _1459_ (.B1(_0348_),
    .Y(_0503_),
    .A1(_0349_),
    .A2(_0372_));
 sg13g2_a21o_1 _1460_ (.A2(\mb.b_1.ball_y[7] ),
    .A1(net304),
    .B1(_0503_),
    .X(_0504_));
 sg13g2_nand2_1 _1461_ (.Y(_0505_),
    .A(\mb.b_1.ball_y[7] ),
    .B(\mb.b_1.ball_y[8] ));
 sg13g2_xor2_1 _1462_ (.B(\mb.b_1.ball_y[8] ),
    .A(\mb.b_1.ball_y[7] ),
    .X(_0506_));
 sg13g2_xnor2_1 _1463_ (.Y(_0507_),
    .A(_0040_),
    .B(_0506_));
 sg13g2_a21oi_1 _1464_ (.A1(_0324_),
    .A2(_0338_),
    .Y(_0508_),
    .B1(_0507_));
 sg13g2_nor2_1 _1465_ (.A(_0323_),
    .B(_0506_),
    .Y(_0509_));
 sg13g2_and2_1 _1466_ (.A(_0044_),
    .B(_0505_),
    .X(_0510_));
 sg13g2_a221oi_1 _1467_ (.B2(\mb.b_0.y[9] ),
    .C1(_0509_),
    .B1(_0510_),
    .A1(_0504_),
    .Y(_0511_),
    .A2(_0508_));
 sg13g2_nor2_1 _1468_ (.A(_0044_),
    .B(_0505_),
    .Y(_0512_));
 sg13g2_nor2_1 _1469_ (.A(\mb.b_0.y[9] ),
    .B(_0510_),
    .Y(_0513_));
 sg13g2_nor3_1 _1470_ (.A(_0511_),
    .B(_0512_),
    .C(_0513_),
    .Y(_0514_));
 sg13g2_o21ai_1 _1471_ (.B1(_0503_),
    .Y(_0515_),
    .A1(net304),
    .A2(_0338_));
 sg13g2_a22oi_1 _1472_ (.Y(_0516_),
    .B1(_0340_),
    .B2(\mb.b_0.y[8] ),
    .A2(_0338_),
    .A1(net304));
 sg13g2_nand2_1 _1473_ (.Y(_0517_),
    .A(_0515_),
    .B(_0516_));
 sg13g2_a22oi_1 _1474_ (.Y(_0518_),
    .B1(\mb.b_1.ball_y[8] ),
    .B2(_0323_),
    .A2(\mb.b_1.ball_y[9] ),
    .A1(_0322_));
 sg13g2_a22oi_1 _1475_ (.Y(_0519_),
    .B1(_0517_),
    .B2(_0518_),
    .A2(_0339_),
    .A1(\mb.b_0.y[9] ));
 sg13g2_or3_2 _1476_ (.A(_0502_),
    .B(_0514_),
    .C(_0519_),
    .X(_0520_));
 sg13g2_nor2_1 _1477_ (.A(_0371_),
    .B(_0520_),
    .Y(_0521_));
 sg13g2_nand2_1 _1478_ (.Y(_0522_),
    .A(net281),
    .B(_0416_));
 sg13g2_nor2_2 _1479_ (.A(net299),
    .B(_0425_),
    .Y(_0523_));
 sg13g2_o21ai_1 _1480_ (.B1(_0523_),
    .Y(_0524_),
    .A1(net285),
    .A2(_0477_));
 sg13g2_a22oi_1 _1481_ (.Y(_0525_),
    .B1(_0522_),
    .B2(_0524_),
    .A2(_0463_),
    .A1(net294));
 sg13g2_nor2b_1 _1482_ (.A(_0525_),
    .B_N(net257),
    .Y(_0526_));
 sg13g2_nand3_1 _1483_ (.B(_0434_),
    .C(_0477_),
    .A(net258),
    .Y(_0527_));
 sg13g2_nor2_1 _1484_ (.A(net296),
    .B(_0527_),
    .Y(_0528_));
 sg13g2_nor3_1 _1485_ (.A(_0431_),
    .B(_0445_),
    .C(_0528_),
    .Y(_0529_));
 sg13g2_nor3_1 _1486_ (.A(net286),
    .B(_0460_),
    .C(_0476_),
    .Y(_0530_));
 sg13g2_nor2_1 _1487_ (.A(net300),
    .B(_0426_),
    .Y(_0531_));
 sg13g2_nor4_1 _1488_ (.A(_0431_),
    .B(_0453_),
    .C(_0530_),
    .D(_0531_),
    .Y(_0532_));
 sg13g2_o21ai_1 _1489_ (.B1(_0449_),
    .Y(_0533_),
    .A1(_0423_),
    .A2(_0425_));
 sg13g2_nand3_1 _1490_ (.B(net297),
    .C(_0464_),
    .A(net284),
    .Y(_0534_));
 sg13g2_nand3_1 _1491_ (.B(_0533_),
    .C(_0534_),
    .A(_0472_),
    .Y(_0535_));
 sg13g2_a21oi_1 _1492_ (.A1(net284),
    .A2(_0425_),
    .Y(_0536_),
    .B1(net294));
 sg13g2_and3_1 _1493_ (.X(_0537_),
    .A(net294),
    .B(_0458_),
    .C(_0464_));
 sg13g2_nor3_1 _1494_ (.A(_0453_),
    .B(_0536_),
    .C(_0537_),
    .Y(_0538_));
 sg13g2_nand2_1 _1495_ (.Y(_0539_),
    .A(net285),
    .B(_0425_));
 sg13g2_nand2_1 _1496_ (.Y(_0540_),
    .A(_0418_),
    .B(_0523_));
 sg13g2_a221oi_1 _1497_ (.B2(net299),
    .C1(_0445_),
    .B1(_0539_),
    .A1(_0418_),
    .Y(_0541_),
    .A2(_0523_));
 sg13g2_nand3_1 _1498_ (.B(net294),
    .C(net257),
    .A(_0415_),
    .Y(_0542_));
 sg13g2_nand2b_2 _1499_ (.Y(_0543_),
    .B(net295),
    .A_N(_0415_));
 sg13g2_a21o_1 _1500_ (.A2(net295),
    .A1(_0415_),
    .B1(net278),
    .X(_0544_));
 sg13g2_o21ai_1 _1501_ (.B1(_0542_),
    .Y(_0545_),
    .A1(_0473_),
    .A2(_0543_));
 sg13g2_nor3_1 _1502_ (.A(_0538_),
    .B(_0541_),
    .C(_0545_),
    .Y(_0546_));
 sg13g2_nand2_1 _1503_ (.Y(_0547_),
    .A(_0377_),
    .B(_0535_));
 sg13g2_nor4_1 _1504_ (.A(_0526_),
    .B(_0529_),
    .C(_0532_),
    .D(_0547_),
    .Y(_0548_));
 sg13g2_o21ai_1 _1505_ (.B1(_0371_),
    .Y(_0549_),
    .A1(net287),
    .A2(_0546_));
 sg13g2_nor2_1 _1506_ (.A(_0548_),
    .B(_0549_),
    .Y(_0550_));
 sg13g2_nor2_1 _1507_ (.A(_0520_),
    .B(_0550_),
    .Y(_0551_));
 sg13g2_o21ai_1 _1508_ (.B1(_0522_),
    .Y(_0552_),
    .A1(net281),
    .A2(_0418_));
 sg13g2_nor2_2 _1509_ (.A(_0417_),
    .B(_0476_),
    .Y(_0553_));
 sg13g2_nor2_1 _1510_ (.A(net298),
    .B(_0553_),
    .Y(_0554_));
 sg13g2_a21oi_1 _1511_ (.A1(_0417_),
    .A2(_0523_),
    .Y(_0555_),
    .B1(net279));
 sg13g2_o21ai_1 _1512_ (.B1(_0555_),
    .Y(_0556_),
    .A1(_0552_),
    .A2(_0554_));
 sg13g2_a21oi_1 _1513_ (.A1(_0431_),
    .A2(_0477_),
    .Y(_0557_),
    .B1(net280));
 sg13g2_a21o_1 _1514_ (.A2(_0458_),
    .A1(_0433_),
    .B1(_0435_),
    .X(_0558_));
 sg13g2_a21oi_1 _1515_ (.A1(_0557_),
    .A2(_0558_),
    .Y(_0559_),
    .B1(net276));
 sg13g2_nor2_1 _1516_ (.A(net280),
    .B(_0459_),
    .Y(_0560_));
 sg13g2_o21ai_1 _1517_ (.B1(_0560_),
    .Y(_0561_),
    .A1(net298),
    .A2(_0552_));
 sg13g2_nand3_1 _1518_ (.B(_0433_),
    .C(_0457_),
    .A(net298),
    .Y(_0562_));
 sg13g2_nand4_1 _1519_ (.B(net280),
    .C(_0431_),
    .A(net258),
    .Y(_0563_),
    .D(_0477_));
 sg13g2_and3_1 _1520_ (.X(_0564_),
    .A(net276),
    .B(_0562_),
    .C(_0563_));
 sg13g2_a221oi_1 _1521_ (.B2(_0564_),
    .C1(_0371_),
    .B1(_0561_),
    .A1(_0556_),
    .Y(_0565_),
    .A2(_0559_));
 sg13g2_nand2_1 _1522_ (.Y(_0566_),
    .A(_0433_),
    .B(_0459_));
 sg13g2_nand2_1 _1523_ (.Y(_0567_),
    .A(_0432_),
    .B(_0461_));
 sg13g2_o21ai_1 _1524_ (.B1(_0566_),
    .Y(_0568_),
    .A1(net299),
    .A2(_0567_));
 sg13g2_nor2_1 _1525_ (.A(net298),
    .B(net280),
    .Y(_0569_));
 sg13g2_nor2_1 _1526_ (.A(net294),
    .B(_0463_),
    .Y(_0570_));
 sg13g2_a21oi_1 _1527_ (.A1(_0407_),
    .A2(_0569_),
    .Y(_0571_),
    .B1(_0570_));
 sg13g2_o21ai_1 _1528_ (.B1(net278),
    .Y(_0572_),
    .A1(_0414_),
    .A2(_0571_));
 sg13g2_a21oi_1 _1529_ (.A1(_0540_),
    .A2(_0571_),
    .Y(_0573_),
    .B1(_0439_));
 sg13g2_nand3_1 _1530_ (.B(_0436_),
    .C(net257),
    .A(net258),
    .Y(_0574_));
 sg13g2_nand2_1 _1531_ (.Y(_0575_),
    .A(_0371_),
    .B(_0574_));
 sg13g2_a221oi_1 _1532_ (.B2(_0573_),
    .C1(_0575_),
    .B1(_0572_),
    .A1(_0472_),
    .Y(_0576_),
    .A2(_0568_));
 sg13g2_nor3_1 _1533_ (.A(_0376_),
    .B(_0565_),
    .C(_0576_),
    .Y(_0577_));
 sg13g2_nand3_1 _1534_ (.B(_0432_),
    .C(_0465_),
    .A(net298),
    .Y(_0578_));
 sg13g2_nand2_1 _1535_ (.Y(_0579_),
    .A(_0458_),
    .B(_0523_));
 sg13g2_a21oi_1 _1536_ (.A1(_0578_),
    .A2(_0579_),
    .Y(_0580_),
    .B1(_0453_));
 sg13g2_nand3_1 _1537_ (.B(net300),
    .C(_0433_),
    .A(_0402_),
    .Y(_0581_));
 sg13g2_a21oi_1 _1538_ (.A1(net284),
    .A2(net296),
    .Y(_0582_),
    .B1(net276));
 sg13g2_a21o_1 _1539_ (.A2(_0582_),
    .A1(_0581_),
    .B1(net257),
    .X(_0583_));
 sg13g2_nor2_1 _1540_ (.A(net295),
    .B(_0553_),
    .Y(_0584_));
 sg13g2_a21oi_1 _1541_ (.A1(net296),
    .A2(_0527_),
    .Y(_0585_),
    .B1(net278));
 sg13g2_nand2b_1 _1542_ (.Y(_0586_),
    .B(_0585_),
    .A_N(_0584_));
 sg13g2_nand2_1 _1543_ (.Y(_0587_),
    .A(_0422_),
    .B(_0433_));
 sg13g2_a21oi_1 _1544_ (.A1(_0436_),
    .A2(_0587_),
    .Y(_0588_),
    .B1(_0445_));
 sg13g2_a21oi_1 _1545_ (.A1(_0583_),
    .A2(_0586_),
    .Y(_0589_),
    .B1(_0580_));
 sg13g2_nor2_1 _1546_ (.A(_0371_),
    .B(_0588_),
    .Y(_0590_));
 sg13g2_a21oi_1 _1547_ (.A1(net300),
    .A2(_0441_),
    .Y(_0591_),
    .B1(_0445_));
 sg13g2_a21oi_1 _1548_ (.A1(_0543_),
    .A2(_0591_),
    .Y(_0592_),
    .B1(_0370_));
 sg13g2_nand2_1 _1549_ (.Y(_0593_),
    .A(_0478_),
    .B(_0523_));
 sg13g2_nand2_1 _1550_ (.Y(_0594_),
    .A(_0415_),
    .B(_0569_));
 sg13g2_a22oi_1 _1551_ (.Y(_0595_),
    .B1(_0594_),
    .B2(_0439_),
    .A2(_0593_),
    .A1(net280));
 sg13g2_a221oi_1 _1552_ (.B2(_0595_),
    .C1(net287),
    .B1(_0592_),
    .A1(_0589_),
    .Y(_0596_),
    .A2(_0590_));
 sg13g2_nor3_2 _1553_ (.A(_0520_),
    .B(_0577_),
    .C(_0596_),
    .Y(_0597_));
 sg13g2_nand2b_1 _1554_ (.Y(_0598_),
    .B(\mb.b_0.y[6] ),
    .A_N(\mb.b_0.ball_y[6] ));
 sg13g2_xor2_1 _1555_ (.B(\mb.b_0.ball_y[6] ),
    .A(\mb.b_0.y[6] ),
    .X(_0599_));
 sg13g2_nand2_1 _1556_ (.Y(_0600_),
    .A(_0326_),
    .B(\mb.b_0.ball_y[5] ));
 sg13g2_nor2_1 _1557_ (.A(_0326_),
    .B(\mb.b_0.ball_y[5] ),
    .Y(_0601_));
 sg13g2_nand2b_1 _1558_ (.Y(_0602_),
    .B(net305),
    .A_N(\mb.b_0.ball_y[4] ));
 sg13g2_nor2b_1 _1559_ (.A(\mb.b_0.ball_y[3] ),
    .B_N(net307),
    .Y(_0603_));
 sg13g2_nor2b_1 _1560_ (.A(\mb.b_0.ball_y[2] ),
    .B_N(net308),
    .Y(_0604_));
 sg13g2_nand2b_1 _1561_ (.Y(_0605_),
    .B(\mb.b_0.ball_y[2] ),
    .A_N(net308));
 sg13g2_nand2b_1 _1562_ (.Y(_0606_),
    .B(_0605_),
    .A_N(_0604_));
 sg13g2_nor2b_1 _1563_ (.A(net309),
    .B_N(\mb.b_0.ball_y[1] ),
    .Y(_0607_));
 sg13g2_nand2b_1 _1564_ (.Y(_0608_),
    .B(net309),
    .A_N(\mb.b_0.ball_y[1] ));
 sg13g2_nor2b_1 _1565_ (.A(\mb.b_0.y[0] ),
    .B_N(\mb.b_0.ball_y[0] ),
    .Y(_0609_));
 sg13g2_a21oi_1 _1566_ (.A1(_0608_),
    .A2(_0609_),
    .Y(_0610_),
    .B1(_0607_));
 sg13g2_a21o_1 _1567_ (.A2(_0610_),
    .A1(_0605_),
    .B1(_0604_),
    .X(_0611_));
 sg13g2_nand2b_1 _1568_ (.Y(_0612_),
    .B(\mb.b_0.ball_y[3] ),
    .A_N(net307));
 sg13g2_nand2b_1 _1569_ (.Y(_0613_),
    .B(_0612_),
    .A_N(_0603_));
 sg13g2_a21oi_1 _1570_ (.A1(_0611_),
    .A2(_0612_),
    .Y(_0614_),
    .B1(_0603_));
 sg13g2_nor2b_1 _1571_ (.A(net306),
    .B_N(\mb.b_0.ball_y[4] ),
    .Y(_0615_));
 sg13g2_xnor2_1 _1572_ (.Y(_0616_),
    .A(net306),
    .B(\mb.b_0.ball_y[4] ));
 sg13g2_o21ai_1 _1573_ (.B1(_0602_),
    .Y(_0617_),
    .A1(_0614_),
    .A2(_0615_));
 sg13g2_a21oi_2 _1574_ (.B1(_0601_),
    .Y(_0618_),
    .A2(_0617_),
    .A1(_0600_));
 sg13g2_o21ai_1 _1575_ (.B1(_0598_),
    .Y(_0619_),
    .A1(_0599_),
    .A2(_0618_));
 sg13g2_a21oi_1 _1576_ (.A1(net304),
    .A2(_0332_),
    .Y(_0620_),
    .B1(_0619_));
 sg13g2_a221oi_1 _1577_ (.B2(_0323_),
    .C1(_0620_),
    .B1(\mb.b_0.ball_y[8] ),
    .A1(_0324_),
    .Y(_0621_),
    .A2(\mb.b_0.ball_y[7] ));
 sg13g2_a21oi_1 _1578_ (.A1(\mb.b_0.y[8] ),
    .A2(_0333_),
    .Y(_0622_),
    .B1(_0621_));
 sg13g2_o21ai_1 _1579_ (.B1(_0622_),
    .Y(_0623_),
    .A1(_0322_),
    .A2(\mb.b_0.ball_y[9] ));
 sg13g2_nor2_1 _1580_ (.A(\mb.b_0.ball_x[6] ),
    .B(_0330_),
    .Y(_0624_));
 sg13g2_xor2_1 _1581_ (.B(\mb.b_0.x[6] ),
    .A(\mb.b_0.ball_x[6] ),
    .X(_0625_));
 sg13g2_nand2b_1 _1582_ (.Y(_0626_),
    .B(\mb.b_0.ball_x[5] ),
    .A_N(\mb.b_0.x[5] ));
 sg13g2_nand2b_1 _1583_ (.Y(_0627_),
    .B(\mb.b_0.x[5] ),
    .A_N(\mb.b_0.ball_x[5] ));
 sg13g2_nor2b_1 _1584_ (.A(\mb.b_0.ball_x[4] ),
    .B_N(\mb.b_0.x[4] ),
    .Y(_0628_));
 sg13g2_xor2_1 _1585_ (.B(net325),
    .A(\mb.b_0.ball_x[4] ),
    .X(_0629_));
 sg13g2_nor2_1 _1586_ (.A(_0331_),
    .B(\mb.b_0.x[3] ),
    .Y(_0630_));
 sg13g2_nor2b_1 _1587_ (.A(\mb.b_0.ball_x[2] ),
    .B_N(\mb.b_0.x[2] ),
    .Y(_0631_));
 sg13g2_xnor2_1 _1588_ (.Y(_0632_),
    .A(\mb.b_0.ball_x[2] ),
    .B(\mb.b_0.x[2] ));
 sg13g2_nor2b_1 _1589_ (.A(\mb.b_0.x[1] ),
    .B_N(\mb.b_0.ball_x[1] ),
    .Y(_0633_));
 sg13g2_nand2b_1 _1590_ (.Y(_0634_),
    .B(\mb.b_0.x[1] ),
    .A_N(\mb.b_0.ball_x[1] ));
 sg13g2_nor2b_1 _1591_ (.A(\mb.b_0.x[0] ),
    .B_N(\mb.b_0.ball_x[0] ),
    .Y(_0635_));
 sg13g2_a21oi_2 _1592_ (.B1(_0633_),
    .Y(_0636_),
    .A2(_0635_),
    .A1(_0634_));
 sg13g2_a21oi_1 _1593_ (.A1(_0632_),
    .A2(_0636_),
    .Y(_0637_),
    .B1(_0631_));
 sg13g2_a221oi_1 _1594_ (.B2(_0636_),
    .C1(_0631_),
    .B1(_0632_),
    .A1(_0331_),
    .Y(_0638_),
    .A2(net326));
 sg13g2_nor3_2 _1595_ (.A(_0629_),
    .B(_0630_),
    .C(_0638_),
    .Y(_0639_));
 sg13g2_nor2_1 _1596_ (.A(_0628_),
    .B(_0639_),
    .Y(_0640_));
 sg13g2_o21ai_1 _1597_ (.B1(_0626_),
    .Y(_0641_),
    .A1(_0628_),
    .A2(_0639_));
 sg13g2_a21oi_2 _1598_ (.B1(_0625_),
    .Y(_0642_),
    .A2(_0641_),
    .A1(_0627_));
 sg13g2_or2_1 _1599_ (.X(_0643_),
    .B(_0642_),
    .A(_0624_));
 sg13g2_nand2b_1 _1600_ (.Y(_0644_),
    .B(net324),
    .A_N(\mb.b_0.ball_x[7] ));
 sg13g2_nand2b_1 _1601_ (.Y(_0645_),
    .B(_0644_),
    .A_N(_0643_));
 sg13g2_nand2b_1 _1602_ (.Y(_0646_),
    .B(\mb.b_0.x[8] ),
    .A_N(\mb.b_0.ball_x[8] ));
 sg13g2_nor2_1 _1603_ (.A(\mb.b_0.ball_x[9] ),
    .B(_0335_),
    .Y(_0647_));
 sg13g2_nand2_1 _1604_ (.Y(_0648_),
    .A(\mb.b_0.ball_x[9] ),
    .B(_0335_));
 sg13g2_a221oi_1 _1605_ (.B2(_0336_),
    .C1(_0647_),
    .B1(\mb.b_0.ball_x[8] ),
    .A1(\mb.b_0.ball_x[7] ),
    .Y(_0649_),
    .A2(_0334_));
 sg13g2_and4_1 _1606_ (.A(_0645_),
    .B(_0646_),
    .C(_0648_),
    .D(_0649_),
    .X(_0650_));
 sg13g2_a21oi_1 _1607_ (.A1(\mb.b_0.ball_x[9] ),
    .A2(_0335_),
    .Y(_0651_),
    .B1(_0646_));
 sg13g2_nor3_1 _1608_ (.A(_0647_),
    .B(_0650_),
    .C(_0651_),
    .Y(_0652_));
 sg13g2_nand2_1 _1609_ (.Y(_0653_),
    .A(\mb.b_0.ball_y[7] ),
    .B(\mb.b_0.ball_y[8] ));
 sg13g2_nand2_1 _1610_ (.Y(_0654_),
    .A(\mb.b_0.y[9] ),
    .B(_0037_));
 sg13g2_nor2b_1 _1611_ (.A(_0654_),
    .B_N(_0653_),
    .Y(_0655_));
 sg13g2_a21oi_1 _1612_ (.A1(\mb.b_0.ball_x[7] ),
    .A2(net324),
    .Y(_0656_),
    .B1(_0643_));
 sg13g2_nand2_1 _1613_ (.Y(_0657_),
    .A(\mb.b_0.ball_x[7] ),
    .B(\mb.b_0.ball_x[8] ));
 sg13g2_xor2_1 _1614_ (.B(\mb.b_0.ball_x[8] ),
    .A(\mb.b_0.ball_x[7] ),
    .X(_0658_));
 sg13g2_nor2_1 _1615_ (.A(\mb.b_0.ball_x[7] ),
    .B(net324),
    .Y(_0659_));
 sg13g2_xnor2_1 _1616_ (.Y(_0660_),
    .A(_0041_),
    .B(_0658_));
 sg13g2_nor3_1 _1617_ (.A(_0656_),
    .B(_0659_),
    .C(_0660_),
    .Y(_0661_));
 sg13g2_nor2_1 _1618_ (.A(_0336_),
    .B(_0658_),
    .Y(_0662_));
 sg13g2_nand2_1 _1619_ (.Y(_0663_),
    .A(_0047_),
    .B(_0657_));
 sg13g2_nor2_1 _1620_ (.A(_0335_),
    .B(_0663_),
    .Y(_0664_));
 sg13g2_nor3_1 _1621_ (.A(_0661_),
    .B(_0662_),
    .C(_0664_),
    .Y(_0665_));
 sg13g2_o21ai_1 _1622_ (.B1(\mb.b_0.x[9] ),
    .Y(_0666_),
    .A1(_0047_),
    .A2(_0657_));
 sg13g2_a21oi_1 _1623_ (.A1(_0663_),
    .A2(_0666_),
    .Y(_0667_),
    .B1(_0665_));
 sg13g2_a21oi_1 _1624_ (.A1(net304),
    .A2(\mb.b_0.ball_y[7] ),
    .Y(_0668_),
    .B1(_0619_));
 sg13g2_xnor2_1 _1625_ (.Y(_0669_),
    .A(\mb.b_0.ball_y[7] ),
    .B(\mb.b_0.ball_y[8] ));
 sg13g2_xor2_1 _1626_ (.B(_0669_),
    .A(_0040_),
    .X(_0670_));
 sg13g2_nor2_1 _1627_ (.A(_0668_),
    .B(_0670_),
    .Y(_0671_));
 sg13g2_o21ai_1 _1628_ (.B1(_0671_),
    .Y(_0672_),
    .A1(net304),
    .A2(\mb.b_0.ball_y[7] ));
 sg13g2_nand2_1 _1629_ (.Y(_0673_),
    .A(\mb.b_0.y[8] ),
    .B(_0669_));
 sg13g2_o21ai_1 _1630_ (.B1(_0653_),
    .Y(_0674_),
    .A1(\mb.b_0.y[9] ),
    .A2(_0037_));
 sg13g2_a22oi_1 _1631_ (.Y(_0675_),
    .B1(_0674_),
    .B2(_0654_),
    .A2(_0673_),
    .A1(_0672_));
 sg13g2_a21oi_1 _1632_ (.A1(_0322_),
    .A2(\mb.b_0.ball_y[9] ),
    .Y(_0676_),
    .B1(_0652_));
 sg13g2_nor3_1 _1633_ (.A(_0655_),
    .B(_0667_),
    .C(_0675_),
    .Y(_0677_));
 sg13g2_nand3_1 _1634_ (.B(_0676_),
    .C(_0677_),
    .A(_0623_),
    .Y(_0678_));
 sg13g2_xor2_1 _1635_ (.B(_0618_),
    .A(_0599_),
    .X(_0679_));
 sg13g2_xnor2_1 _1636_ (.Y(_0680_),
    .A(_0614_),
    .B(_0616_));
 sg13g2_xnor2_1 _1637_ (.Y(_0681_),
    .A(_0679_),
    .B(_0680_));
 sg13g2_inv_1 _1638_ (.Y(_0682_),
    .A(_0681_));
 sg13g2_mux2_1 _1639_ (.A0(_0627_),
    .A1(_0626_),
    .S(_0640_),
    .X(_0683_));
 sg13g2_xor2_1 _1640_ (.B(_0683_),
    .A(_0625_),
    .X(_0684_));
 sg13g2_xnor2_1 _1641_ (.Y(_0685_),
    .A(_0625_),
    .B(_0683_));
 sg13g2_xnor2_1 _1642_ (.Y(_0686_),
    .A(_0606_),
    .B(_0610_));
 sg13g2_xnor2_1 _1643_ (.Y(_0687_),
    .A(_0679_),
    .B(_0686_));
 sg13g2_xor2_1 _1644_ (.B(_0686_),
    .A(_0679_),
    .X(_0688_));
 sg13g2_nor2_1 _1645_ (.A(net292),
    .B(net273),
    .Y(_0689_));
 sg13g2_and3_1 _1646_ (.X(_0690_),
    .A(_0625_),
    .B(_0627_),
    .C(_0641_));
 sg13g2_or2_2 _1647_ (.X(_0691_),
    .B(_0690_),
    .A(_0642_));
 sg13g2_xnor2_1 _1648_ (.Y(_0692_),
    .A(\mb.b_0.ball_x[3] ),
    .B(net326));
 sg13g2_xnor2_1 _1649_ (.Y(_0693_),
    .A(_0637_),
    .B(_0692_));
 sg13g2_o21ai_1 _1650_ (.B1(_0693_),
    .Y(_0694_),
    .A1(_0642_),
    .A2(_0690_));
 sg13g2_or3_1 _1651_ (.A(_0642_),
    .B(_0690_),
    .C(_0693_),
    .X(_0695_));
 sg13g2_nand2_2 _1652_ (.Y(_0696_),
    .A(_0694_),
    .B(_0695_));
 sg13g2_and2_1 _1653_ (.A(_0694_),
    .B(_0695_),
    .X(_0697_));
 sg13g2_xor2_1 _1654_ (.B(_0636_),
    .A(_0632_),
    .X(_0698_));
 sg13g2_xor2_1 _1655_ (.B(_0698_),
    .A(_0691_),
    .X(_0699_));
 sg13g2_xnor2_1 _1656_ (.Y(_0700_),
    .A(_0691_),
    .B(_0698_));
 sg13g2_nand2_2 _1657_ (.Y(_0701_),
    .A(net269),
    .B(net268));
 sg13g2_o21ai_1 _1658_ (.B1(_0629_),
    .Y(_0702_),
    .A1(_0630_),
    .A2(_0638_));
 sg13g2_nor2b_2 _1659_ (.A(_0639_),
    .B_N(_0702_),
    .Y(_0703_));
 sg13g2_xor2_1 _1660_ (.B(_0703_),
    .A(_0691_),
    .X(_0704_));
 sg13g2_xnor2_1 _1661_ (.Y(_0705_),
    .A(_0691_),
    .B(_0703_));
 sg13g2_a21oi_2 _1662_ (.B1(net288),
    .Y(_0706_),
    .A2(net261),
    .A1(net270));
 sg13g2_o21ai_1 _1663_ (.B1(net291),
    .Y(_0707_),
    .A1(net271),
    .A2(net264));
 sg13g2_a21oi_1 _1664_ (.A1(_0689_),
    .A2(_0701_),
    .Y(_0708_),
    .B1(_0706_));
 sg13g2_xnor2_1 _1665_ (.Y(_0709_),
    .A(_0611_),
    .B(_0613_));
 sg13g2_xnor2_1 _1666_ (.Y(_0710_),
    .A(_0679_),
    .B(_0709_));
 sg13g2_xor2_1 _1667_ (.B(_0709_),
    .A(_0679_),
    .X(_0711_));
 sg13g2_nand2_2 _1668_ (.Y(_0712_),
    .A(net274),
    .B(net259));
 sg13g2_nor2_1 _1669_ (.A(net270),
    .B(net268),
    .Y(_0713_));
 sg13g2_nand2_2 _1670_ (.Y(_0714_),
    .A(net271),
    .B(net267));
 sg13g2_xor2_1 _1671_ (.B(_0698_),
    .A(_0693_),
    .X(_0715_));
 sg13g2_xnor2_1 _1672_ (.Y(_0716_),
    .A(_0693_),
    .B(_0698_));
 sg13g2_nor2_2 _1673_ (.A(net269),
    .B(net265),
    .Y(_0717_));
 sg13g2_nand2_2 _1674_ (.Y(_0718_),
    .A(net271),
    .B(net263));
 sg13g2_a21oi_2 _1675_ (.B1(net291),
    .Y(_0719_),
    .A2(net263),
    .A1(net271));
 sg13g2_nand4_1 _1676_ (.B(net259),
    .C(_0716_),
    .A(net274),
    .Y(_0720_),
    .D(_0719_));
 sg13g2_a221oi_1 _1677_ (.B2(_0708_),
    .C1(_0710_),
    .B1(_0720_),
    .A1(net272),
    .Y(_0721_),
    .A2(_0713_));
 sg13g2_nor2_2 _1678_ (.A(net274),
    .B(net259),
    .Y(_0722_));
 sg13g2_nor2_2 _1679_ (.A(_0699_),
    .B(net265),
    .Y(_0723_));
 sg13g2_nand2_2 _1680_ (.Y(_0724_),
    .A(net267),
    .B(net261));
 sg13g2_a21oi_2 _1681_ (.B1(net289),
    .Y(_0725_),
    .A2(net263),
    .A1(net266));
 sg13g2_nor2_1 _1682_ (.A(net289),
    .B(_0717_),
    .Y(_0726_));
 sg13g2_nand2_2 _1683_ (.Y(_0727_),
    .A(net292),
    .B(_0718_));
 sg13g2_nor2_1 _1684_ (.A(net270),
    .B(net263),
    .Y(_0728_));
 sg13g2_nand2_2 _1685_ (.Y(_0729_),
    .A(_0696_),
    .B(net265));
 sg13g2_nand2_1 _1686_ (.Y(_0730_),
    .A(_0699_),
    .B(net262));
 sg13g2_nand3_1 _1687_ (.B(net268),
    .C(net263),
    .A(net270),
    .Y(_0731_));
 sg13g2_xnor2_1 _1688_ (.Y(_0732_),
    .A(_0693_),
    .B(_0703_));
 sg13g2_and2_1 _1689_ (.A(_0729_),
    .B(_0731_),
    .X(_0733_));
 sg13g2_nand2_1 _1690_ (.Y(_0734_),
    .A(net288),
    .B(_0733_));
 sg13g2_o21ai_1 _1691_ (.B1(_0734_),
    .Y(_0735_),
    .A1(_0723_),
    .A2(_0727_));
 sg13g2_nand2_1 _1692_ (.Y(_0736_),
    .A(net266),
    .B(net264));
 sg13g2_a21oi_2 _1693_ (.B1(net292),
    .Y(_0737_),
    .A2(net265),
    .A1(net266));
 sg13g2_nor2_2 _1694_ (.A(net272),
    .B(net259),
    .Y(_0738_));
 sg13g2_nand2_2 _1695_ (.Y(_0739_),
    .A(net274),
    .B(_0710_));
 sg13g2_a21oi_1 _1696_ (.A1(net269),
    .A2(_0737_),
    .Y(_0740_),
    .B1(_0717_));
 sg13g2_a221oi_1 _1697_ (.B2(_0740_),
    .C1(_0721_),
    .B1(_0738_),
    .A1(_0722_),
    .Y(_0741_),
    .A2(_0735_));
 sg13g2_nor2_1 _1698_ (.A(_0600_),
    .B(_0617_),
    .Y(_0742_));
 sg13g2_a21oi_2 _1699_ (.B1(_0742_),
    .Y(_0743_),
    .A2(_0617_),
    .A1(_0601_));
 sg13g2_xnor2_1 _1700_ (.Y(_0744_),
    .A(_0599_),
    .B(_0743_));
 sg13g2_xor2_1 _1701_ (.B(_0743_),
    .A(_0599_),
    .X(_0745_));
 sg13g2_o21ai_1 _1702_ (.B1(net288),
    .Y(_0746_),
    .A1(_0696_),
    .A2(net262));
 sg13g2_nor2_2 _1703_ (.A(net267),
    .B(net261),
    .Y(_0747_));
 sg13g2_nor2_1 _1704_ (.A(_0746_),
    .B(_0747_),
    .Y(_0748_));
 sg13g2_or2_2 _1705_ (.X(_0749_),
    .B(_0747_),
    .A(_0746_));
 sg13g2_nand2_1 _1706_ (.Y(_0750_),
    .A(net290),
    .B(net268));
 sg13g2_nand3_1 _1707_ (.B(net266),
    .C(net263),
    .A(net271),
    .Y(_0751_));
 sg13g2_a22oi_1 _1708_ (.Y(_0752_),
    .B1(_0751_),
    .B2(net292),
    .A2(_0717_),
    .A1(net273));
 sg13g2_a22oi_1 _1709_ (.Y(_0753_),
    .B1(_0752_),
    .B2(net260),
    .A2(_0748_),
    .A1(_0688_));
 sg13g2_nand3_1 _1710_ (.B(net269),
    .C(_0747_),
    .A(net273),
    .Y(_0754_));
 sg13g2_nor2_1 _1711_ (.A(net274),
    .B(_0710_),
    .Y(_0755_));
 sg13g2_nand2_2 _1712_ (.Y(_0756_),
    .A(net272),
    .B(net259));
 sg13g2_o21ai_1 _1713_ (.B1(_0754_),
    .Y(_0757_),
    .A1(_0749_),
    .A2(_0756_));
 sg13g2_o21ai_1 _1714_ (.B1(net275),
    .Y(_0758_),
    .A1(_0753_),
    .A2(_0757_));
 sg13g2_and2_1 _1715_ (.A(_0745_),
    .B(_0758_),
    .X(_0759_));
 sg13g2_o21ai_1 _1716_ (.B1(_0759_),
    .Y(_0760_),
    .A1(net275),
    .A2(_0741_));
 sg13g2_a22oi_1 _1717_ (.Y(_0761_),
    .B1(_0725_),
    .B2(net271),
    .A2(net266),
    .A1(net289));
 sg13g2_nand2_1 _1718_ (.Y(_0762_),
    .A(net264),
    .B(_0715_));
 sg13g2_a22oi_1 _1719_ (.Y(_0763_),
    .B1(_0762_),
    .B2(_0725_),
    .A2(_0737_),
    .A1(_0729_));
 sg13g2_a21oi_1 _1720_ (.A1(net259),
    .A2(_0763_),
    .Y(_0764_),
    .B1(net274));
 sg13g2_o21ai_1 _1721_ (.B1(_0764_),
    .Y(_0765_),
    .A1(net259),
    .A2(_0761_));
 sg13g2_nor2_2 _1722_ (.A(_0715_),
    .B(_0747_),
    .Y(_0766_));
 sg13g2_nor2_1 _1723_ (.A(net288),
    .B(_0766_),
    .Y(_0767_));
 sg13g2_nor2_2 _1724_ (.A(net293),
    .B(net269),
    .Y(_0768_));
 sg13g2_a21oi_2 _1725_ (.B1(net292),
    .Y(_0769_),
    .A2(net261),
    .A1(net269));
 sg13g2_o21ai_1 _1726_ (.B1(net288),
    .Y(_0770_),
    .A1(_0696_),
    .A2(net265));
 sg13g2_o21ai_1 _1727_ (.B1(_0769_),
    .Y(_0771_),
    .A1(net266),
    .A2(_0729_));
 sg13g2_o21ai_1 _1728_ (.B1(_0771_),
    .Y(_0772_),
    .A1(_0685_),
    .A2(_0766_));
 sg13g2_nor2_1 _1729_ (.A(net264),
    .B(_0716_),
    .Y(_0773_));
 sg13g2_o21ai_1 _1730_ (.B1(net290),
    .Y(_0774_),
    .A1(_0728_),
    .A2(_0773_));
 sg13g2_a21oi_1 _1731_ (.A1(_0762_),
    .A2(_0769_),
    .Y(_0775_),
    .B1(_0712_));
 sg13g2_nand2_2 _1732_ (.Y(_0776_),
    .A(net275),
    .B(_0744_));
 sg13g2_a221oi_1 _1733_ (.B2(_0775_),
    .C1(_0776_),
    .B1(_0774_),
    .A1(_0738_),
    .Y(_0777_),
    .A2(_0772_));
 sg13g2_nor2_1 _1734_ (.A(net275),
    .B(_0745_),
    .Y(_0778_));
 sg13g2_nand2_1 _1735_ (.Y(_0779_),
    .A(_0682_),
    .B(_0744_));
 sg13g2_o21ai_1 _1736_ (.B1(net264),
    .Y(_0780_),
    .A1(net271),
    .A2(net268));
 sg13g2_nor2_2 _1737_ (.A(net267),
    .B(_0746_),
    .Y(_0781_));
 sg13g2_a22oi_1 _1738_ (.Y(_0782_),
    .B1(_0781_),
    .B2(_0718_),
    .A2(_0780_),
    .A1(_0725_));
 sg13g2_nor2_1 _1739_ (.A(_0716_),
    .B(_0717_),
    .Y(_0783_));
 sg13g2_nand3_1 _1740_ (.B(net268),
    .C(_0732_),
    .A(net290),
    .Y(_0784_));
 sg13g2_a221oi_1 _1741_ (.B2(_0719_),
    .C1(_0739_),
    .B1(_0715_),
    .A1(net264),
    .Y(_0785_),
    .A2(_0713_));
 sg13g2_a21oi_1 _1742_ (.A1(net269),
    .A2(_0747_),
    .Y(_0786_),
    .B1(net293));
 sg13g2_o21ai_1 _1743_ (.B1(net289),
    .Y(_0787_),
    .A1(_0701_),
    .A2(net263));
 sg13g2_nand2_2 _1744_ (.Y(_0788_),
    .A(net264),
    .B(_0716_));
 sg13g2_nand3_1 _1745_ (.B(net268),
    .C(net263),
    .A(net271),
    .Y(_0789_));
 sg13g2_nand3_1 _1746_ (.B(_0788_),
    .C(_0789_),
    .A(net289),
    .Y(_0790_));
 sg13g2_a22oi_1 _1747_ (.Y(_0791_),
    .B1(_0725_),
    .B2(_0780_),
    .A2(_0717_),
    .A1(net290));
 sg13g2_a21oi_1 _1748_ (.A1(_0790_),
    .A2(_0791_),
    .Y(_0792_),
    .B1(_0756_));
 sg13g2_a21oi_1 _1749_ (.A1(_0724_),
    .A2(_0788_),
    .Y(_0793_),
    .B1(_0737_));
 sg13g2_nor2_1 _1750_ (.A(_0781_),
    .B(_0793_),
    .Y(_0794_));
 sg13g2_a221oi_1 _1751_ (.B2(_0722_),
    .C1(_0792_),
    .B1(_0794_),
    .A1(_0784_),
    .Y(_0795_),
    .A2(_0785_));
 sg13g2_o21ai_1 _1752_ (.B1(_0795_),
    .Y(_0796_),
    .A1(_0712_),
    .A2(_0782_));
 sg13g2_a22oi_1 _1753_ (.Y(_0797_),
    .B1(_0778_),
    .B2(_0796_),
    .A2(_0777_),
    .A1(_0765_));
 sg13g2_a21oi_1 _1754_ (.A1(_0760_),
    .A2(_0797_),
    .Y(_0798_),
    .B1(_0678_));
 sg13g2_nand2_1 _1755_ (.Y(_0799_),
    .A(_0597_),
    .B(_0798_));
 sg13g2_a22oi_1 _1756_ (.Y(_0800_),
    .B1(_0788_),
    .B2(_0726_),
    .A2(_0737_),
    .A1(_0731_));
 sg13g2_nor2_1 _1757_ (.A(net272),
    .B(_0800_),
    .Y(_0801_));
 sg13g2_o21ai_1 _1758_ (.B1(net289),
    .Y(_0802_),
    .A1(_0728_),
    .A2(_0773_));
 sg13g2_o21ai_1 _1759_ (.B1(_0788_),
    .Y(_0803_),
    .A1(net264),
    .A2(_0713_));
 sg13g2_xnor2_1 _1760_ (.Y(_0804_),
    .A(_0802_),
    .B(_0803_));
 sg13g2_nor2_1 _1761_ (.A(net274),
    .B(_0804_),
    .Y(_0805_));
 sg13g2_o21ai_1 _1762_ (.B1(net259),
    .Y(_0806_),
    .A1(_0801_),
    .A2(_0805_));
 sg13g2_nand3_1 _1763_ (.B(_0731_),
    .C(_0736_),
    .A(net291),
    .Y(_0807_));
 sg13g2_nand3_1 _1764_ (.B(_0787_),
    .C(_0807_),
    .A(_0738_),
    .Y(_0808_));
 sg13g2_a22oi_1 _1765_ (.Y(_0809_),
    .B1(_0780_),
    .B2(net291),
    .A2(_0737_),
    .A1(_0701_));
 sg13g2_nand2b_1 _1766_ (.Y(_0810_),
    .B(_0722_),
    .A_N(_0809_));
 sg13g2_nand4_1 _1767_ (.B(_0806_),
    .C(_0808_),
    .A(_0744_),
    .Y(_0811_),
    .D(_0810_));
 sg13g2_nand2_1 _1768_ (.Y(_0812_),
    .A(net290),
    .B(_0732_));
 sg13g2_o21ai_1 _1769_ (.B1(_0812_),
    .Y(_0813_),
    .A1(net290),
    .A2(net268));
 sg13g2_o21ai_1 _1770_ (.B1(_0813_),
    .Y(_0814_),
    .A1(net290),
    .A2(_0718_));
 sg13g2_a21oi_1 _1771_ (.A1(_0750_),
    .A2(_0814_),
    .Y(_0815_),
    .B1(_0712_));
 sg13g2_nand2_1 _1772_ (.Y(_0816_),
    .A(net289),
    .B(_0780_));
 sg13g2_nand2_1 _1773_ (.Y(_0817_),
    .A(_0707_),
    .B(_0816_));
 sg13g2_and2_1 _1774_ (.A(_0738_),
    .B(_0751_),
    .X(_0818_));
 sg13g2_nor3_2 _1775_ (.A(_0723_),
    .B(_0747_),
    .C(_0770_),
    .Y(_0819_));
 sg13g2_nand3_1 _1776_ (.B(_0699_),
    .C(_0717_),
    .A(_0689_),
    .Y(_0820_));
 sg13g2_nand3_1 _1777_ (.B(_0718_),
    .C(_0730_),
    .A(net272),
    .Y(_0821_));
 sg13g2_o21ai_1 _1778_ (.B1(_0820_),
    .Y(_0822_),
    .A1(_0819_),
    .A2(_0821_));
 sg13g2_a221oi_1 _1779_ (.B2(_0710_),
    .C1(_0744_),
    .B1(_0822_),
    .A1(_0817_),
    .Y(_0823_),
    .A2(_0818_));
 sg13g2_nand2b_1 _1780_ (.Y(_0824_),
    .B(_0736_),
    .A_N(_0813_));
 sg13g2_a21oi_1 _1781_ (.A1(_0755_),
    .A2(_0824_),
    .Y(_0825_),
    .B1(_0815_));
 sg13g2_a21oi_1 _1782_ (.A1(_0823_),
    .A2(_0825_),
    .Y(_0826_),
    .B1(net275));
 sg13g2_a21oi_1 _1783_ (.A1(_0724_),
    .A2(_0788_),
    .Y(_0827_),
    .B1(_0727_));
 sg13g2_nor3_1 _1784_ (.A(net291),
    .B(net266),
    .C(_0728_),
    .Y(_0828_));
 sg13g2_nor3_1 _1785_ (.A(_0739_),
    .B(_0827_),
    .C(_0828_),
    .Y(_0829_));
 sg13g2_a21oi_1 _1786_ (.A1(net292),
    .A2(_0747_),
    .Y(_0830_),
    .B1(_0768_));
 sg13g2_nand2_1 _1787_ (.Y(_0831_),
    .A(_0724_),
    .B(_0830_));
 sg13g2_a21oi_1 _1788_ (.A1(_0751_),
    .A2(_0831_),
    .Y(_0832_),
    .B1(_0712_));
 sg13g2_a21oi_1 _1789_ (.A1(_0730_),
    .A2(_0768_),
    .Y(_0833_),
    .B1(_0756_));
 sg13g2_o21ai_1 _1790_ (.B1(_0833_),
    .Y(_0834_),
    .A1(_0707_),
    .A2(_0747_));
 sg13g2_nand3_1 _1791_ (.B(_0750_),
    .C(_0751_),
    .A(_0722_),
    .Y(_0835_));
 sg13g2_nand3_1 _1792_ (.B(_0834_),
    .C(_0835_),
    .A(_0744_),
    .Y(_0836_));
 sg13g2_nor3_1 _1793_ (.A(_0829_),
    .B(_0832_),
    .C(_0836_),
    .Y(_0837_));
 sg13g2_a21oi_1 _1794_ (.A1(net293),
    .A2(_0751_),
    .Y(_0838_),
    .B1(_0712_));
 sg13g2_a221oi_1 _1795_ (.B2(_0788_),
    .C1(_0712_),
    .B1(_0769_),
    .A1(net293),
    .Y(_0839_),
    .A2(_0751_));
 sg13g2_a221oi_1 _1796_ (.B2(net290),
    .C1(_0756_),
    .B1(_0789_),
    .A1(_0716_),
    .Y(_0840_),
    .A2(_0719_));
 sg13g2_nand4_1 _1797_ (.B(net265),
    .C(_0714_),
    .A(net288),
    .Y(_0841_),
    .D(_0722_));
 sg13g2_o21ai_1 _1798_ (.B1(_0841_),
    .Y(_0842_),
    .A1(_0739_),
    .A2(_0749_));
 sg13g2_nor4_1 _1799_ (.A(_0744_),
    .B(_0839_),
    .C(_0840_),
    .D(_0842_),
    .Y(_0843_));
 sg13g2_o21ai_1 _1800_ (.B1(net275),
    .Y(_0844_),
    .A1(_0837_),
    .A2(_0843_));
 sg13g2_a21oi_1 _1801_ (.A1(_0811_),
    .A2(_0826_),
    .Y(_0845_),
    .B1(_0678_));
 sg13g2_a22oi_1 _1802_ (.Y(_0846_),
    .B1(_0844_),
    .B2(_0845_),
    .A2(_0551_),
    .A1(_0484_));
 sg13g2_o21ai_1 _1803_ (.B1(_0722_),
    .Y(_0847_),
    .A1(_0773_),
    .A2(_0816_));
 sg13g2_o21ai_1 _1804_ (.B1(_0769_),
    .Y(_0848_),
    .A1(net269),
    .A2(net267));
 sg13g2_nand3_1 _1805_ (.B(_0701_),
    .C(net261),
    .A(_0689_),
    .Y(_0849_));
 sg13g2_nand3_1 _1806_ (.B(_0848_),
    .C(_0849_),
    .A(net260),
    .Y(_0850_));
 sg13g2_nor3_1 _1807_ (.A(_0726_),
    .B(_0739_),
    .C(_0783_),
    .Y(_0851_));
 sg13g2_a22oi_1 _1808_ (.Y(_0852_),
    .B1(_0847_),
    .B2(_0850_),
    .A2(_0726_),
    .A1(_0724_));
 sg13g2_nor3_1 _1809_ (.A(_0779_),
    .B(_0851_),
    .C(_0852_),
    .Y(_0853_));
 sg13g2_and2_1 _1810_ (.A(_0719_),
    .B(_0722_),
    .X(_0854_));
 sg13g2_a221oi_1 _1811_ (.B2(_0724_),
    .C1(net275),
    .B1(_0854_),
    .A1(_0738_),
    .Y(_0855_),
    .A2(_0786_));
 sg13g2_a21oi_1 _1812_ (.A1(net273),
    .A2(_0749_),
    .Y(_0856_),
    .B1(_0787_));
 sg13g2_a21oi_1 _1813_ (.A1(_0855_),
    .A2(_0856_),
    .Y(_0857_),
    .B1(_0744_));
 sg13g2_a21oi_1 _1814_ (.A1(_0689_),
    .A2(net262),
    .Y(_0858_),
    .B1(net260));
 sg13g2_nor2_1 _1815_ (.A(net273),
    .B(_0768_),
    .Y(_0859_));
 sg13g2_nand2_1 _1816_ (.Y(_0860_),
    .A(net260),
    .B(_0727_));
 sg13g2_nand3_1 _1817_ (.B(_0727_),
    .C(_0859_),
    .A(net260),
    .Y(_0861_));
 sg13g2_nand2b_1 _1818_ (.Y(_0862_),
    .B(_0861_),
    .A_N(_0776_));
 sg13g2_a221oi_1 _1819_ (.B2(_0752_),
    .C1(_0862_),
    .B1(_0858_),
    .A1(_0733_),
    .Y(_0863_),
    .A2(_0838_));
 sg13g2_nor4_2 _1820_ (.A(_0678_),
    .B(_0853_),
    .C(_0857_),
    .Y(_0864_),
    .D(_0863_));
 sg13g2_nand3_1 _1821_ (.B(_0457_),
    .C(_0465_),
    .A(net294),
    .Y(_0865_));
 sg13g2_nand2_1 _1822_ (.Y(_0866_),
    .A(_0472_),
    .B(_0865_));
 sg13g2_nand3_1 _1823_ (.B(net281),
    .C(_0569_),
    .A(_0407_),
    .Y(_0867_));
 sg13g2_nand3_1 _1824_ (.B(net294),
    .C(_0464_),
    .A(_0416_),
    .Y(_0868_));
 sg13g2_nand3_1 _1825_ (.B(_0867_),
    .C(_0868_),
    .A(net277),
    .Y(_0869_));
 sg13g2_a22oi_1 _1826_ (.Y(_0870_),
    .B1(_0866_),
    .B2(_0869_),
    .A2(_0459_),
    .A1(_0433_));
 sg13g2_nand2_1 _1827_ (.Y(_0871_),
    .A(_0460_),
    .B(net257));
 sg13g2_a21oi_1 _1828_ (.A1(_0417_),
    .A2(net258),
    .Y(_0872_),
    .B1(_0871_));
 sg13g2_o21ai_1 _1829_ (.B1(net287),
    .Y(_0873_),
    .A1(_0870_),
    .A2(_0872_));
 sg13g2_nor3_1 _1830_ (.A(_0453_),
    .B(_0536_),
    .C(_0567_),
    .Y(_0874_));
 sg13g2_o21ai_1 _1831_ (.B1(_0472_),
    .Y(_0875_),
    .A1(net282),
    .A2(net299));
 sg13g2_nor3_1 _1832_ (.A(_0445_),
    .B(_0448_),
    .C(_0459_),
    .Y(_0876_));
 sg13g2_a21oi_1 _1833_ (.A1(net257),
    .A2(_0523_),
    .Y(_0877_),
    .B1(_0876_));
 sg13g2_o21ai_1 _1834_ (.B1(_0877_),
    .Y(_0878_),
    .A1(_0536_),
    .A2(_0875_));
 sg13g2_o21ai_1 _1835_ (.B1(_0376_),
    .Y(_0879_),
    .A1(_0874_),
    .A2(_0878_));
 sg13g2_and2_1 _1836_ (.A(_0370_),
    .B(_0873_),
    .X(_0880_));
 sg13g2_nand3_1 _1837_ (.B(_0472_),
    .C(_0523_),
    .A(_0433_),
    .Y(_0881_));
 sg13g2_nand3_1 _1838_ (.B(_0480_),
    .C(_0881_),
    .A(net287),
    .Y(_0882_));
 sg13g2_nand3_1 _1839_ (.B(_0478_),
    .C(_0544_),
    .A(net295),
    .Y(_0883_));
 sg13g2_nor3_1 _1840_ (.A(_0520_),
    .B(_0882_),
    .C(_0883_),
    .Y(_0884_));
 sg13g2_nor2_1 _1841_ (.A(_0521_),
    .B(_0884_),
    .Y(_0885_));
 sg13g2_a21oi_1 _1842_ (.A1(_0879_),
    .A2(_0880_),
    .Y(_0886_),
    .B1(_0885_));
 sg13g2_nor2_1 _1843_ (.A(_0864_),
    .B(_0886_),
    .Y(_0887_));
 sg13g2_o21ai_1 _1844_ (.B1(_0718_),
    .Y(_0888_),
    .A1(_0737_),
    .A2(_0768_));
 sg13g2_nand2_1 _1845_ (.Y(_0889_),
    .A(_0729_),
    .B(_0767_));
 sg13g2_a221oi_1 _1846_ (.B2(_0889_),
    .C1(_0779_),
    .B1(_0888_),
    .A1(net272),
    .Y(_0890_),
    .A2(_0766_));
 sg13g2_o21ai_1 _1847_ (.B1(_0730_),
    .Y(_0891_),
    .A1(_0706_),
    .A2(_0737_));
 sg13g2_nor2_1 _1848_ (.A(net272),
    .B(_0768_),
    .Y(_0892_));
 sg13g2_o21ai_1 _1849_ (.B1(_0706_),
    .Y(_0893_),
    .A1(net261),
    .A2(_0714_));
 sg13g2_nor2_1 _1850_ (.A(_0687_),
    .B(_0781_),
    .Y(_0894_));
 sg13g2_a221oi_1 _1851_ (.B2(_0894_),
    .C1(_0776_),
    .B1(_0893_),
    .A1(_0891_),
    .Y(_0895_),
    .A2(_0892_));
 sg13g2_o21ai_1 _1852_ (.B1(net260),
    .Y(_0896_),
    .A1(_0890_),
    .A2(_0895_));
 sg13g2_a21oi_1 _1853_ (.A1(_0769_),
    .A2(_0788_),
    .Y(_0897_),
    .B1(_0767_));
 sg13g2_nor2_1 _1854_ (.A(net272),
    .B(_0819_),
    .Y(_0898_));
 sg13g2_a221oi_1 _1855_ (.B2(_0893_),
    .C1(_0779_),
    .B1(_0898_),
    .A1(_0688_),
    .Y(_0899_),
    .A2(_0897_));
 sg13g2_nand3_1 _1856_ (.B(net261),
    .C(_0714_),
    .A(net292),
    .Y(_0900_));
 sg13g2_o21ai_1 _1857_ (.B1(_0769_),
    .Y(_0901_),
    .A1(net261),
    .A2(_0714_));
 sg13g2_o21ai_1 _1858_ (.B1(_0901_),
    .Y(_0902_),
    .A1(_0723_),
    .A2(_0727_));
 sg13g2_a22oi_1 _1859_ (.Y(_0903_),
    .B1(_0902_),
    .B2(net273),
    .A2(_0900_),
    .A1(_0859_));
 sg13g2_nor2_1 _1860_ (.A(_0776_),
    .B(_0903_),
    .Y(_0904_));
 sg13g2_o21ai_1 _1861_ (.B1(_0710_),
    .Y(_0905_),
    .A1(_0899_),
    .A2(_0904_));
 sg13g2_a21oi_1 _1862_ (.A1(net266),
    .A2(net265),
    .Y(_0906_),
    .B1(net273));
 sg13g2_a22oi_1 _1863_ (.Y(_0907_),
    .B1(_0906_),
    .B2(_0733_),
    .A2(_0749_),
    .A1(net273));
 sg13g2_o21ai_1 _1864_ (.B1(_0855_),
    .Y(_0908_),
    .A1(_0860_),
    .A2(_0907_));
 sg13g2_a21oi_1 _1865_ (.A1(net288),
    .A2(_0717_),
    .Y(_0909_),
    .B1(_0688_));
 sg13g2_nor3_1 _1866_ (.A(_0710_),
    .B(_0749_),
    .C(_0909_),
    .Y(_0910_));
 sg13g2_o21ai_1 _1867_ (.B1(_0908_),
    .Y(_0911_),
    .A1(_0682_),
    .A2(_0910_));
 sg13g2_a21oi_1 _1868_ (.A1(_0745_),
    .A2(_0911_),
    .Y(_0912_),
    .B1(_0678_));
 sg13g2_nand3_1 _1869_ (.B(_0905_),
    .C(_0912_),
    .A(_0896_),
    .Y(_0913_));
 sg13g2_nand4_1 _1870_ (.B(_0432_),
    .C(_0434_),
    .A(net278),
    .Y(_0914_),
    .D(_0461_));
 sg13g2_a221oi_1 _1871_ (.B2(_0914_),
    .C1(_0439_),
    .B1(_0544_),
    .A1(net300),
    .Y(_0915_),
    .A2(_0426_));
 sg13g2_nor2_1 _1872_ (.A(net278),
    .B(_0531_),
    .Y(_0916_));
 sg13g2_nand3_1 _1873_ (.B(net295),
    .C(net276),
    .A(_0415_),
    .Y(_0917_));
 sg13g2_o21ai_1 _1874_ (.B1(_0376_),
    .Y(_0918_),
    .A1(_0916_),
    .A2(_0917_));
 sg13g2_o21ai_1 _1875_ (.B1(_0918_),
    .Y(_0919_),
    .A1(_0882_),
    .A2(_0915_));
 sg13g2_a21oi_1 _1876_ (.A1(_0371_),
    .A2(_0919_),
    .Y(_0920_),
    .B1(_0520_));
 sg13g2_nand2_1 _1877_ (.Y(_0921_),
    .A(_0432_),
    .B(_0584_));
 sg13g2_a22oi_1 _1878_ (.Y(_0922_),
    .B1(_0921_),
    .B2(_0524_),
    .A2(_0553_),
    .A1(net278));
 sg13g2_o21ai_1 _1879_ (.B1(_0472_),
    .Y(_0923_),
    .A1(_0537_),
    .A2(_0584_));
 sg13g2_o21ai_1 _1880_ (.B1(_0570_),
    .Y(_0924_),
    .A1(net286),
    .A2(_0432_));
 sg13g2_and2_1 _1881_ (.A(_0434_),
    .B(_0539_),
    .X(_0925_));
 sg13g2_o21ai_1 _1882_ (.B1(_0924_),
    .Y(_0926_),
    .A1(net301),
    .A2(_0925_));
 sg13g2_nand2_1 _1883_ (.Y(_0927_),
    .A(_0377_),
    .B(_0923_));
 sg13g2_a221oi_1 _1884_ (.B2(net257),
    .C1(_0927_),
    .B1(_0926_),
    .A1(net277),
    .Y(_0928_),
    .A2(_0922_));
 sg13g2_o21ai_1 _1885_ (.B1(_0424_),
    .Y(_0929_),
    .A1(_0435_),
    .A2(_0570_));
 sg13g2_nand3_1 _1886_ (.B(_0449_),
    .C(_0929_),
    .A(_0429_),
    .Y(_0930_));
 sg13g2_a21oi_1 _1887_ (.A1(_0557_),
    .A2(_0924_),
    .Y(_0931_),
    .B1(_0439_));
 sg13g2_nand3_1 _1888_ (.B(_0566_),
    .C(_0916_),
    .A(_0543_),
    .Y(_0932_));
 sg13g2_nor3_1 _1889_ (.A(net282),
    .B(_0414_),
    .C(net297),
    .Y(_0933_));
 sg13g2_o21ai_1 _1890_ (.B1(net278),
    .Y(_0934_),
    .A1(_0448_),
    .A2(_0933_));
 sg13g2_nand3_1 _1891_ (.B(_0932_),
    .C(_0934_),
    .A(_0439_),
    .Y(_0935_));
 sg13g2_a21oi_1 _1892_ (.A1(_0930_),
    .A2(_0931_),
    .Y(_0936_),
    .B1(net287));
 sg13g2_a21o_1 _1893_ (.A2(_0936_),
    .A1(_0935_),
    .B1(_0371_),
    .X(_0937_));
 sg13g2_o21ai_1 _1894_ (.B1(_0920_),
    .Y(_0938_),
    .A1(_0928_),
    .A2(_0937_));
 sg13g2_or2_1 _1895_ (.X(_0939_),
    .B(_0938_),
    .A(_0913_));
 sg13g2_nor2_1 _1896_ (.A(_0597_),
    .B(_0798_),
    .Y(_0940_));
 sg13g2_a221oi_1 _1897_ (.B2(_0939_),
    .C1(_0940_),
    .B1(_0887_),
    .A1(_0799_),
    .Y(_0941_),
    .A2(_0846_));
 sg13g2_o21ai_1 _1898_ (.B1(_0858_),
    .Y(_0942_),
    .A1(net292),
    .A2(_0718_));
 sg13g2_a21oi_1 _1899_ (.A1(net260),
    .A2(_0746_),
    .Y(_0943_),
    .B1(_0682_));
 sg13g2_nor3_1 _1900_ (.A(_0701_),
    .B(net262),
    .C(net260),
    .Y(_0944_));
 sg13g2_nor2_1 _1901_ (.A(net275),
    .B(_0944_),
    .Y(_0945_));
 sg13g2_a22oi_1 _1902_ (.Y(_0946_),
    .B1(_0945_),
    .B2(net288),
    .A2(_0943_),
    .A1(_0942_));
 sg13g2_nor3_1 _1903_ (.A(_0678_),
    .B(_0745_),
    .C(_0946_),
    .Y(_0947_));
 sg13g2_nor3_1 _1904_ (.A(net301),
    .B(net258),
    .C(_0445_),
    .Y(_0948_));
 sg13g2_nor4_1 _1905_ (.A(net283),
    .B(net301),
    .C(net277),
    .D(_0916_),
    .Y(_0949_));
 sg13g2_nand3_1 _1906_ (.B(net276),
    .C(_0477_),
    .A(net295),
    .Y(_0950_));
 sg13g2_a21oi_1 _1907_ (.A1(_0425_),
    .A2(net278),
    .Y(_0951_),
    .B1(_0950_));
 sg13g2_a21oi_1 _1908_ (.A1(net295),
    .A2(net277),
    .Y(_0952_),
    .B1(_0376_));
 sg13g2_nor4_1 _1909_ (.A(net287),
    .B(_0948_),
    .C(_0949_),
    .D(_0951_),
    .Y(_0953_));
 sg13g2_nand2b_1 _1910_ (.Y(_0954_),
    .B(_0521_),
    .A_N(_0953_));
 sg13g2_a21oi_1 _1911_ (.A1(_0479_),
    .A2(_0952_),
    .Y(_0955_),
    .B1(_0954_));
 sg13g2_and2_1 _1912_ (.A(_0913_),
    .B(_0938_),
    .X(_0956_));
 sg13g2_nand2_1 _1913_ (.Y(_0957_),
    .A(_0864_),
    .B(_0886_));
 sg13g2_a21oi_1 _1914_ (.A1(_0956_),
    .A2(_0957_),
    .Y(_0958_),
    .B1(_0887_));
 sg13g2_or4_1 _1915_ (.A(_0941_),
    .B(_0947_),
    .C(_0955_),
    .D(_0958_),
    .X(_0000_));
 sg13g2_and2_1 _1916_ (.A(\mb.b_1.ball_y[6] ),
    .B(\mb.b_1.ball_vy[8] ),
    .X(_0959_));
 sg13g2_xnor2_1 _1917_ (.Y(_0960_),
    .A(\mb.b_1.ball_y[6] ),
    .B(\mb.b_1.ball_vy[8] ));
 sg13g2_nor2_1 _1918_ (.A(\mb.b_1.ball_y[5] ),
    .B(\mb.b_1.ball_vy[7] ),
    .Y(_0961_));
 sg13g2_and2_1 _1919_ (.A(\mb.b_1.ball_y[4] ),
    .B(\mb.b_1.ball_vy[6] ),
    .X(_0962_));
 sg13g2_nand2_1 _1920_ (.Y(_0963_),
    .A(\mb.b_1.ball_y[3] ),
    .B(\mb.b_1.ball_vy[5] ));
 sg13g2_xor2_1 _1921_ (.B(\mb.b_1.ball_vy[5] ),
    .A(\mb.b_1.ball_y[3] ),
    .X(_0964_));
 sg13g2_inv_1 _1922_ (.Y(_0965_),
    .A(_0964_));
 sg13g2_and2_1 _1923_ (.A(\mb.b_1.ball_y[2] ),
    .B(\mb.b_1.ball_vy[4] ),
    .X(_0966_));
 sg13g2_or2_1 _1924_ (.X(_0967_),
    .B(\mb.b_1.ball_vy[4] ),
    .A(\mb.b_1.ball_y[2] ));
 sg13g2_nand2b_1 _1925_ (.Y(_0968_),
    .B(_0967_),
    .A_N(_0966_));
 sg13g2_nand2_1 _1926_ (.Y(_0969_),
    .A(\mb.b_1.ball_y[1] ),
    .B(\mb.b_1.ball_vy[3] ));
 sg13g2_nand2_1 _1927_ (.Y(_0970_),
    .A(\mb.b_1.ball_y[0] ),
    .B(\mb.b_1.ball_vy[2] ));
 sg13g2_nor2_1 _1928_ (.A(\mb.b_1.ball_y[1] ),
    .B(\mb.b_1.ball_vy[3] ),
    .Y(_0971_));
 sg13g2_xor2_1 _1929_ (.B(\mb.b_1.ball_vy[3] ),
    .A(\mb.b_1.ball_y[1] ),
    .X(_0972_));
 sg13g2_o21ai_1 _1930_ (.B1(_0969_),
    .Y(_0973_),
    .A1(_0970_),
    .A2(_0971_));
 sg13g2_a21oi_1 _1931_ (.A1(_0967_),
    .A2(_0973_),
    .Y(_0974_),
    .B1(_0966_));
 sg13g2_o21ai_1 _1932_ (.B1(_0963_),
    .Y(_0975_),
    .A1(_0965_),
    .A2(_0974_));
 sg13g2_or2_1 _1933_ (.X(_0976_),
    .B(\mb.b_1.ball_vy[6] ),
    .A(\mb.b_1.ball_y[4] ));
 sg13g2_nand2b_1 _1934_ (.Y(_0977_),
    .B(_0976_),
    .A_N(_0962_));
 sg13g2_a21oi_1 _1935_ (.A1(_0975_),
    .A2(_0976_),
    .Y(_0978_),
    .B1(_0962_));
 sg13g2_a221oi_1 _1936_ (.B2(_0976_),
    .C1(_0962_),
    .B1(_0975_),
    .A1(\mb.b_1.ball_y[5] ),
    .Y(_0979_),
    .A2(\mb.b_1.ball_vy[7] ));
 sg13g2_nor3_2 _1937_ (.A(_0960_),
    .B(_0961_),
    .C(_0979_),
    .Y(_0980_));
 sg13g2_o21ai_1 _1938_ (.B1(_0960_),
    .Y(_0981_),
    .A1(_0961_),
    .A2(_0979_));
 sg13g2_nor2b_1 _1939_ (.A(_0980_),
    .B_N(_0981_),
    .Y(\mb.b_1.next_y[6] ));
 sg13g2_nand2_1 _1940_ (.Y(_0982_),
    .A(\mb.b_1.ball_y[7] ),
    .B(\mb.b_1.ball_vy[9] ));
 sg13g2_xor2_1 _1941_ (.B(\mb.b_1.ball_vy[9] ),
    .A(\mb.b_1.ball_y[7] ),
    .X(_0983_));
 sg13g2_o21ai_1 _1942_ (.B1(_0983_),
    .Y(_0984_),
    .A1(_0959_),
    .A2(_0980_));
 sg13g2_or3_1 _1943_ (.A(_0959_),
    .B(_0980_),
    .C(_0983_),
    .X(_0985_));
 sg13g2_and2_1 _1944_ (.A(_0984_),
    .B(_0985_),
    .X(\mb.b_1.next_y[7] ));
 sg13g2_and2_1 _1945_ (.A(\mb.b_1.ball_x[4] ),
    .B(\mb.b_1.ball_vx[6] ),
    .X(_0986_));
 sg13g2_xnor2_1 _1946_ (.Y(_0987_),
    .A(\mb.b_1.ball_x[4] ),
    .B(\mb.b_1.ball_vx[6] ));
 sg13g2_inv_1 _1947_ (.Y(_0988_),
    .A(_0987_));
 sg13g2_and2_1 _1948_ (.A(\mb.b_1.ball_x[3] ),
    .B(\mb.b_1.ball_vx[5] ),
    .X(_0989_));
 sg13g2_or2_1 _1949_ (.X(_0990_),
    .B(\mb.b_1.ball_vx[5] ),
    .A(\mb.b_1.ball_x[3] ));
 sg13g2_nand2b_1 _1950_ (.Y(_0991_),
    .B(_0990_),
    .A_N(_0989_));
 sg13g2_and2_1 _1951_ (.A(\mb.b_1.ball_x[2] ),
    .B(\mb.b_1.ball_vx[4] ),
    .X(_0992_));
 sg13g2_or2_1 _1952_ (.X(_0993_),
    .B(\mb.b_1.ball_vx[4] ),
    .A(\mb.b_1.ball_x[2] ));
 sg13g2_nand2b_1 _1953_ (.Y(_0994_),
    .B(_0993_),
    .A_N(_0992_));
 sg13g2_nand2_1 _1954_ (.Y(_0995_),
    .A(\mb.b_1.ball_x[1] ),
    .B(\mb.b_1.ball_vx[3] ));
 sg13g2_nand2_1 _1955_ (.Y(_0996_),
    .A(\mb.b_1.ball_x[0] ),
    .B(\mb.b_1.ball_vx[2] ));
 sg13g2_nor2_1 _1956_ (.A(\mb.b_1.ball_x[1] ),
    .B(\mb.b_1.ball_vx[3] ),
    .Y(_0997_));
 sg13g2_xor2_1 _1957_ (.B(\mb.b_1.ball_vx[3] ),
    .A(\mb.b_1.ball_x[1] ),
    .X(_0998_));
 sg13g2_o21ai_1 _1958_ (.B1(_0995_),
    .Y(_0999_),
    .A1(_0996_),
    .A2(_0997_));
 sg13g2_a21o_1 _1959_ (.A2(_0999_),
    .A1(_0993_),
    .B1(_0992_),
    .X(_1000_));
 sg13g2_a21o_1 _1960_ (.A2(_1000_),
    .A1(_0990_),
    .B1(_0989_),
    .X(_1001_));
 sg13g2_xnor2_1 _1961_ (.Y(\mb.b_1.next_x[4] ),
    .A(_0987_),
    .B(_1001_));
 sg13g2_and2_1 _1962_ (.A(\mb.b_1.ball_x[6] ),
    .B(\mb.b_1.ball_vx[8] ),
    .X(_1002_));
 sg13g2_xor2_1 _1963_ (.B(\mb.b_1.ball_vx[8] ),
    .A(\mb.b_1.ball_x[6] ),
    .X(_1003_));
 sg13g2_inv_1 _1964_ (.Y(_1004_),
    .A(_1003_));
 sg13g2_nor2_1 _1965_ (.A(\mb.b_1.ball_x[5] ),
    .B(\mb.b_1.ball_vx[7] ),
    .Y(_1005_));
 sg13g2_a21oi_1 _1966_ (.A1(_0988_),
    .A2(_1001_),
    .Y(_1006_),
    .B1(_0986_));
 sg13g2_a221oi_1 _1967_ (.B2(_1001_),
    .C1(_0986_),
    .B1(_0988_),
    .A1(\mb.b_1.ball_x[5] ),
    .Y(_1007_),
    .A2(\mb.b_1.ball_vx[7] ));
 sg13g2_nor3_1 _1968_ (.A(_1004_),
    .B(_1005_),
    .C(_1007_),
    .Y(_1008_));
 sg13g2_o21ai_1 _1969_ (.B1(_1004_),
    .Y(_1009_),
    .A1(_1005_),
    .A2(_1007_));
 sg13g2_nor2b_1 _1970_ (.A(_1008_),
    .B_N(_1009_),
    .Y(\mb.b_1.next_x[6] ));
 sg13g2_nand2_1 _1971_ (.Y(_1010_),
    .A(\mb.b_0.ball_x[0] ),
    .B(\mb.b_0.ball_vx[2] ));
 sg13g2_xor2_1 _1972_ (.B(\mb.b_0.ball_vx[2] ),
    .A(\mb.b_0.ball_x[0] ),
    .X(\mb.b_0.next_x[0] ));
 sg13g2_nand2_1 _1973_ (.Y(_1011_),
    .A(\mb.b_0.ball_x[1] ),
    .B(\mb.b_0.ball_vx[3] ));
 sg13g2_nor2_1 _1974_ (.A(\mb.b_0.ball_x[1] ),
    .B(\mb.b_0.ball_vx[3] ),
    .Y(_1012_));
 sg13g2_xor2_1 _1975_ (.B(\mb.b_0.ball_vx[3] ),
    .A(\mb.b_0.ball_x[1] ),
    .X(_1013_));
 sg13g2_xnor2_1 _1976_ (.Y(\mb.b_0.next_x[1] ),
    .A(_1010_),
    .B(_1013_));
 sg13g2_and2_1 _1977_ (.A(\mb.b_0.ball_x[2] ),
    .B(\mb.b_0.ball_vx[4] ),
    .X(_1014_));
 sg13g2_or2_1 _1978_ (.X(_1015_),
    .B(\mb.b_0.ball_vx[4] ),
    .A(\mb.b_0.ball_x[2] ));
 sg13g2_nand2b_1 _1979_ (.Y(_1016_),
    .B(_1015_),
    .A_N(_1014_));
 sg13g2_o21ai_1 _1980_ (.B1(_1011_),
    .Y(_1017_),
    .A1(_1010_),
    .A2(_1012_));
 sg13g2_xnor2_1 _1981_ (.Y(\mb.b_0.next_x[2] ),
    .A(_1016_),
    .B(_1017_));
 sg13g2_and2_1 _1982_ (.A(\mb.b_0.ball_x[3] ),
    .B(\mb.b_0.ball_vx[5] ),
    .X(_1018_));
 sg13g2_or2_1 _1983_ (.X(_1019_),
    .B(\mb.b_0.ball_vx[5] ),
    .A(\mb.b_0.ball_x[3] ));
 sg13g2_nand2b_1 _1984_ (.Y(_1020_),
    .B(_1019_),
    .A_N(_1018_));
 sg13g2_a21o_1 _1985_ (.A2(_1017_),
    .A1(_1015_),
    .B1(_1014_),
    .X(_1021_));
 sg13g2_xnor2_1 _1986_ (.Y(\mb.b_0.next_x[3] ),
    .A(_1020_),
    .B(_1021_));
 sg13g2_and2_1 _1987_ (.A(\mb.b_0.ball_x[4] ),
    .B(\mb.b_0.ball_vx[6] ),
    .X(_1022_));
 sg13g2_xnor2_1 _1988_ (.Y(_1023_),
    .A(\mb.b_0.ball_x[4] ),
    .B(\mb.b_0.ball_vx[6] ));
 sg13g2_inv_1 _1989_ (.Y(_1024_),
    .A(_1023_));
 sg13g2_a21o_1 _1990_ (.A2(_1021_),
    .A1(_1019_),
    .B1(_1018_),
    .X(_1025_));
 sg13g2_xnor2_1 _1991_ (.Y(\mb.b_0.next_x[4] ),
    .A(_1023_),
    .B(_1025_));
 sg13g2_a21oi_1 _1992_ (.A1(_1024_),
    .A2(_1025_),
    .Y(_1026_),
    .B1(_1022_));
 sg13g2_nor2_1 _1993_ (.A(\mb.b_0.ball_x[5] ),
    .B(\mb.b_0.ball_vx[7] ),
    .Y(_1027_));
 sg13g2_xor2_1 _1994_ (.B(\mb.b_0.ball_vx[7] ),
    .A(\mb.b_0.ball_x[5] ),
    .X(_1028_));
 sg13g2_xnor2_1 _1995_ (.Y(\mb.b_0.next_x[5] ),
    .A(_1026_),
    .B(_1028_));
 sg13g2_and2_1 _1996_ (.A(\mb.b_0.ball_x[6] ),
    .B(\mb.b_0.ball_vx[8] ),
    .X(_1029_));
 sg13g2_xnor2_1 _1997_ (.Y(_1030_),
    .A(\mb.b_0.ball_x[6] ),
    .B(\mb.b_0.ball_vx[8] ));
 sg13g2_a221oi_1 _1998_ (.B2(_1025_),
    .C1(_1022_),
    .B1(_1024_),
    .A1(\mb.b_0.ball_x[5] ),
    .Y(_1031_),
    .A2(\mb.b_0.ball_vx[7] ));
 sg13g2_nor3_1 _1999_ (.A(_1027_),
    .B(_1030_),
    .C(_1031_),
    .Y(_1032_));
 sg13g2_o21ai_1 _2000_ (.B1(_1030_),
    .Y(_1033_),
    .A1(_1027_),
    .A2(_1031_));
 sg13g2_nor2b_1 _2001_ (.A(_1032_),
    .B_N(_1033_),
    .Y(\mb.b_0.next_x[6] ));
 sg13g2_nand2_1 _2002_ (.Y(_1034_),
    .A(\mb.b_0.ball_x[7] ),
    .B(\mb.b_0.ball_vx[9] ));
 sg13g2_xor2_1 _2003_ (.B(\mb.b_0.ball_vx[9] ),
    .A(\mb.b_0.ball_x[7] ),
    .X(_1035_));
 sg13g2_o21ai_1 _2004_ (.B1(_1035_),
    .Y(_1036_),
    .A1(_1029_),
    .A2(_1032_));
 sg13g2_or3_1 _2005_ (.A(_1029_),
    .B(_1032_),
    .C(_1035_),
    .X(_1037_));
 sg13g2_and2_1 _2006_ (.A(_1036_),
    .B(_1037_),
    .X(\mb.b_0.next_x[7] ));
 sg13g2_nand2_1 _2007_ (.Y(_1038_),
    .A(\mb.b_0.ball_x[8] ),
    .B(\mb.b_0.ball_vx[9] ));
 sg13g2_xnor2_1 _2008_ (.Y(_1039_),
    .A(\mb.b_0.ball_x[8] ),
    .B(\mb.b_0.ball_vx[9] ));
 sg13g2_a21oi_1 _2009_ (.A1(_1034_),
    .A2(_1036_),
    .Y(_1040_),
    .B1(_1039_));
 sg13g2_a21o_1 _2010_ (.A2(_1036_),
    .A1(_1034_),
    .B1(_1039_),
    .X(_1041_));
 sg13g2_and3_1 _2011_ (.X(_1042_),
    .A(_1034_),
    .B(_1036_),
    .C(_1039_));
 sg13g2_nor2_1 _2012_ (.A(_1040_),
    .B(_1042_),
    .Y(\mb.b_0.next_x[8] ));
 sg13g2_xnor2_1 _2013_ (.Y(_1043_),
    .A(\mb.b_0.ball_x[9] ),
    .B(\mb.b_0.ball_vx[9] ));
 sg13g2_inv_1 _2014_ (.Y(_1044_),
    .A(_1043_));
 sg13g2_a21oi_1 _2015_ (.A1(_1038_),
    .A2(_1041_),
    .Y(_1045_),
    .B1(_1044_));
 sg13g2_and3_1 _2016_ (.X(_1046_),
    .A(_1038_),
    .B(_1041_),
    .C(_1044_));
 sg13g2_or2_1 _2017_ (.X(\mb.b_0.next_x[9] ),
    .B(_1046_),
    .A(_1045_));
 sg13g2_nand2_1 _2018_ (.Y(_1047_),
    .A(\mb.b_0.ball_y[0] ),
    .B(\mb.b_0.ball_vy[2] ));
 sg13g2_xor2_1 _2019_ (.B(\mb.b_0.ball_vy[2] ),
    .A(\mb.b_0.ball_y[0] ),
    .X(\mb.b_0.next_y[0] ));
 sg13g2_nand2_1 _2020_ (.Y(_1048_),
    .A(\mb.b_0.ball_y[1] ),
    .B(\mb.b_0.ball_vy[3] ));
 sg13g2_nor2_1 _2021_ (.A(\mb.b_0.ball_y[1] ),
    .B(\mb.b_0.ball_vy[3] ),
    .Y(_1049_));
 sg13g2_xor2_1 _2022_ (.B(\mb.b_0.ball_vy[3] ),
    .A(\mb.b_0.ball_y[1] ),
    .X(_1050_));
 sg13g2_xnor2_1 _2023_ (.Y(\mb.b_0.next_y[1] ),
    .A(_1047_),
    .B(_1050_));
 sg13g2_and2_1 _2024_ (.A(\mb.b_0.ball_y[2] ),
    .B(\mb.b_0.ball_vy[4] ),
    .X(_1051_));
 sg13g2_or2_1 _2025_ (.X(_1052_),
    .B(\mb.b_0.ball_vy[4] ),
    .A(\mb.b_0.ball_y[2] ));
 sg13g2_nand2b_1 _2026_ (.Y(_1053_),
    .B(_1052_),
    .A_N(_1051_));
 sg13g2_o21ai_1 _2027_ (.B1(_1048_),
    .Y(_1054_),
    .A1(_1047_),
    .A2(_1049_));
 sg13g2_xnor2_1 _2028_ (.Y(\mb.b_0.next_y[2] ),
    .A(_1053_),
    .B(_1054_));
 sg13g2_a21o_1 _2029_ (.A2(_1054_),
    .A1(_1052_),
    .B1(_1051_),
    .X(_1055_));
 sg13g2_and2_1 _2030_ (.A(\mb.b_0.ball_y[3] ),
    .B(\mb.b_0.ball_vy[5] ),
    .X(_1056_));
 sg13g2_or2_1 _2031_ (.X(_1057_),
    .B(\mb.b_0.ball_vy[5] ),
    .A(\mb.b_0.ball_y[3] ));
 sg13g2_nand2b_1 _2032_ (.Y(_1058_),
    .B(_1057_),
    .A_N(_1056_));
 sg13g2_xnor2_1 _2033_ (.Y(\mb.b_0.next_y[3] ),
    .A(_1055_),
    .B(_1058_));
 sg13g2_and2_1 _2034_ (.A(\mb.b_0.ball_y[4] ),
    .B(\mb.b_0.ball_vy[6] ),
    .X(_1059_));
 sg13g2_or2_1 _2035_ (.X(_1060_),
    .B(\mb.b_0.ball_vy[6] ),
    .A(\mb.b_0.ball_y[4] ));
 sg13g2_nand2b_1 _2036_ (.Y(_1061_),
    .B(_1060_),
    .A_N(_1059_));
 sg13g2_a21o_1 _2037_ (.A2(_1057_),
    .A1(_1055_),
    .B1(_1056_),
    .X(_1062_));
 sg13g2_xnor2_1 _2038_ (.Y(\mb.b_0.next_y[4] ),
    .A(_1061_),
    .B(_1062_));
 sg13g2_a21o_1 _2039_ (.A2(_1062_),
    .A1(_1060_),
    .B1(_1059_),
    .X(_1063_));
 sg13g2_nor2_1 _2040_ (.A(\mb.b_0.ball_y[5] ),
    .B(\mb.b_0.ball_vy[7] ),
    .Y(_1064_));
 sg13g2_xnor2_1 _2041_ (.Y(_1065_),
    .A(\mb.b_0.ball_y[5] ),
    .B(\mb.b_0.ball_vy[7] ));
 sg13g2_xnor2_1 _2042_ (.Y(\mb.b_0.next_y[5] ),
    .A(_1063_),
    .B(_1065_));
 sg13g2_and2_1 _2043_ (.A(\mb.b_0.ball_y[6] ),
    .B(\mb.b_0.ball_vy[8] ),
    .X(_1066_));
 sg13g2_xnor2_1 _2044_ (.Y(_1067_),
    .A(\mb.b_0.ball_y[6] ),
    .B(\mb.b_0.ball_vy[8] ));
 sg13g2_a221oi_1 _2045_ (.B2(_1062_),
    .C1(_1059_),
    .B1(_1060_),
    .A1(\mb.b_0.ball_y[5] ),
    .Y(_1068_),
    .A2(\mb.b_0.ball_vy[7] ));
 sg13g2_nor3_1 _2046_ (.A(_1064_),
    .B(_1067_),
    .C(_1068_),
    .Y(_1069_));
 sg13g2_o21ai_1 _2047_ (.B1(_1067_),
    .Y(_1070_),
    .A1(_1064_),
    .A2(_1068_));
 sg13g2_nor2b_1 _2048_ (.A(_1069_),
    .B_N(_1070_),
    .Y(\mb.b_0.next_y[6] ));
 sg13g2_nand2_1 _2049_ (.Y(_1071_),
    .A(\mb.b_0.ball_y[7] ),
    .B(\mb.b_0.ball_vy[9] ));
 sg13g2_xor2_1 _2050_ (.B(\mb.b_0.ball_vy[9] ),
    .A(\mb.b_0.ball_y[7] ),
    .X(_1072_));
 sg13g2_o21ai_1 _2051_ (.B1(_1072_),
    .Y(_1073_),
    .A1(_1066_),
    .A2(_1069_));
 sg13g2_or3_1 _2052_ (.A(_1066_),
    .B(_1069_),
    .C(_1072_),
    .X(_1074_));
 sg13g2_and2_1 _2053_ (.A(_1073_),
    .B(_1074_),
    .X(\mb.b_0.next_y[7] ));
 sg13g2_and2_1 _2054_ (.A(\mb.b_0.ball_y[8] ),
    .B(\mb.b_0.ball_vy[9] ),
    .X(_1075_));
 sg13g2_xnor2_1 _2055_ (.Y(_1076_),
    .A(\mb.b_0.ball_y[8] ),
    .B(\mb.b_0.ball_vy[9] ));
 sg13g2_a21oi_1 _2056_ (.A1(_1071_),
    .A2(_1073_),
    .Y(_0073_),
    .B1(_1076_));
 sg13g2_a21o_1 _2057_ (.A2(_1073_),
    .A1(_1071_),
    .B1(_1076_),
    .X(_0074_));
 sg13g2_nand3_1 _2058_ (.B(_1073_),
    .C(_1076_),
    .A(_1071_),
    .Y(_0075_));
 sg13g2_and2_1 _2059_ (.A(_0074_),
    .B(_0075_),
    .X(\mb.b_0.next_y[8] ));
 sg13g2_xnor2_1 _2060_ (.Y(_0076_),
    .A(\mb.b_0.ball_y[9] ),
    .B(\mb.b_0.ball_vy[9] ));
 sg13g2_o21ai_1 _2061_ (.B1(_0076_),
    .Y(_0077_),
    .A1(_1075_),
    .A2(_0073_));
 sg13g2_or3_1 _2062_ (.A(_1075_),
    .B(_0073_),
    .C(_0076_),
    .X(_0078_));
 sg13g2_nand2_1 _2063_ (.Y(\mb.b_0.next_y[9] ),
    .A(_0077_),
    .B(_0078_));
 sg13g2_xor2_1 _2064_ (.B(\mb.b_1.ball_vy[2] ),
    .A(\mb.b_1.ball_y[0] ),
    .X(\mb.b_1.next_y[0] ));
 sg13g2_xnor2_1 _2065_ (.Y(\mb.b_1.next_y[1] ),
    .A(_0970_),
    .B(_0972_));
 sg13g2_xnor2_1 _2066_ (.Y(\mb.b_1.next_y[2] ),
    .A(_0968_),
    .B(_0973_));
 sg13g2_xnor2_1 _2067_ (.Y(\mb.b_1.next_y[3] ),
    .A(_0964_),
    .B(_0974_));
 sg13g2_xnor2_1 _2068_ (.Y(\mb.b_1.next_y[4] ),
    .A(_0975_),
    .B(_0977_));
 sg13g2_xor2_1 _2069_ (.B(\mb.b_1.ball_vy[7] ),
    .A(\mb.b_1.ball_y[5] ),
    .X(_0079_));
 sg13g2_xnor2_1 _2070_ (.Y(\mb.b_1.next_y[5] ),
    .A(_0978_),
    .B(_0079_));
 sg13g2_and2_1 _2071_ (.A(\mb.b_1.ball_y[8] ),
    .B(\mb.b_1.ball_vy[9] ),
    .X(_0080_));
 sg13g2_xnor2_1 _2072_ (.Y(_0081_),
    .A(\mb.b_1.ball_y[8] ),
    .B(\mb.b_1.ball_vy[9] ));
 sg13g2_a21oi_1 _2073_ (.A1(_0982_),
    .A2(_0984_),
    .Y(_0082_),
    .B1(_0081_));
 sg13g2_a21o_1 _2074_ (.A2(_0984_),
    .A1(_0982_),
    .B1(_0081_),
    .X(_0083_));
 sg13g2_nand3_1 _2075_ (.B(_0984_),
    .C(_0081_),
    .A(_0982_),
    .Y(_0084_));
 sg13g2_and2_1 _2076_ (.A(_0083_),
    .B(_0084_),
    .X(\mb.b_1.next_y[8] ));
 sg13g2_xnor2_1 _2077_ (.Y(_0085_),
    .A(\mb.b_1.ball_y[9] ),
    .B(\mb.b_1.ball_vy[9] ));
 sg13g2_o21ai_1 _2078_ (.B1(_0085_),
    .Y(_0086_),
    .A1(_0080_),
    .A2(_0082_));
 sg13g2_or3_1 _2079_ (.A(_0080_),
    .B(_0082_),
    .C(_0085_),
    .X(_0087_));
 sg13g2_nand2_1 _2080_ (.Y(\mb.b_1.next_y[9] ),
    .A(_0086_),
    .B(_0087_));
 sg13g2_xor2_1 _2081_ (.B(\mb.b_1.ball_vx[2] ),
    .A(\mb.b_1.ball_x[0] ),
    .X(\mb.b_1.next_x[0] ));
 sg13g2_xnor2_1 _2082_ (.Y(\mb.b_1.next_x[1] ),
    .A(_0996_),
    .B(_0998_));
 sg13g2_xnor2_1 _2083_ (.Y(\mb.b_1.next_x[2] ),
    .A(_0994_),
    .B(_0999_));
 sg13g2_xnor2_1 _2084_ (.Y(\mb.b_1.next_x[3] ),
    .A(_0991_),
    .B(_1000_));
 sg13g2_xor2_1 _2085_ (.B(\mb.b_1.ball_vx[7] ),
    .A(\mb.b_1.ball_x[5] ),
    .X(_0088_));
 sg13g2_xnor2_1 _2086_ (.Y(\mb.b_1.next_x[5] ),
    .A(_1006_),
    .B(_0088_));
 sg13g2_nand2_1 _2087_ (.Y(_0089_),
    .A(\mb.b_1.ball_x[7] ),
    .B(\mb.b_1.ball_vx[9] ));
 sg13g2_xor2_1 _2088_ (.B(\mb.b_1.ball_vx[9] ),
    .A(\mb.b_1.ball_x[7] ),
    .X(_0090_));
 sg13g2_o21ai_1 _2089_ (.B1(_0090_),
    .Y(_0091_),
    .A1(_1002_),
    .A2(_1008_));
 sg13g2_or3_1 _2090_ (.A(_1002_),
    .B(_1008_),
    .C(_0090_),
    .X(_0092_));
 sg13g2_and2_1 _2091_ (.A(_0091_),
    .B(_0092_),
    .X(\mb.b_1.next_x[7] ));
 sg13g2_and2_1 _2092_ (.A(\mb.b_1.ball_x[8] ),
    .B(\mb.b_1.ball_vx[9] ),
    .X(_0093_));
 sg13g2_xnor2_1 _2093_ (.Y(_0094_),
    .A(\mb.b_1.ball_x[8] ),
    .B(\mb.b_1.ball_vx[9] ));
 sg13g2_a21oi_2 _2094_ (.B1(_0094_),
    .Y(_0095_),
    .A2(_0091_),
    .A1(_0089_));
 sg13g2_and3_1 _2095_ (.X(_0096_),
    .A(_0089_),
    .B(_0091_),
    .C(_0094_));
 sg13g2_nor2_1 _2096_ (.A(_0095_),
    .B(_0096_),
    .Y(\mb.b_1.next_x[8] ));
 sg13g2_xnor2_1 _2097_ (.Y(_0097_),
    .A(\mb.b_1.ball_x[9] ),
    .B(\mb.b_1.ball_vx[9] ));
 sg13g2_inv_1 _2098_ (.Y(_0098_),
    .A(_0097_));
 sg13g2_o21ai_1 _2099_ (.B1(_0098_),
    .Y(_0099_),
    .A1(_0093_),
    .A2(_0095_));
 sg13g2_or3_1 _2100_ (.A(_0093_),
    .B(_0095_),
    .C(_0098_),
    .X(_0100_));
 sg13g2_and2_1 _2101_ (.A(_0099_),
    .B(_0100_),
    .X(\mb.b_1.next_x[9] ));
 sg13g2_and3_1 _2102_ (.X(\mb.rgb ),
    .A(\v.h_display ),
    .B(\v.v_display ),
    .C(\mb.pix ));
 sg13g2_a21o_1 _2103_ (.A2(\mb.b_0.next_y[3] ),
    .A1(\mb.b_0.next_y[2] ),
    .B1(\mb.b_0.next_y[4] ),
    .X(_0101_));
 sg13g2_and3_1 _2104_ (.X(_0102_),
    .A(\mb.b_0.next_y[5] ),
    .B(\mb.b_0.next_y[6] ),
    .C(_0101_));
 sg13g2_a22oi_1 _2105_ (.Y(_0103_),
    .B1(_0102_),
    .B2(\mb.b_0.next_y[7] ),
    .A2(_0075_),
    .A1(_0074_));
 sg13g2_nand3_1 _2106_ (.B(_0078_),
    .C(_0103_),
    .A(_0077_),
    .Y(_0104_));
 sg13g2_nand2_1 _2107_ (.Y(_0105_),
    .A(\mb.b_0.ball_vy[1] ),
    .B(net254));
 sg13g2_xor2_1 _2108_ (.B(net254),
    .A(\mb.b_0.ball_vy[1] ),
    .X(_0106_));
 sg13g2_xnor2_1 _2109_ (.Y(_0010_),
    .A(_0039_),
    .B(_0106_));
 sg13g2_and2_1 _2110_ (.A(\mb.b_0.ball_vy[2] ),
    .B(net255),
    .X(_0107_));
 sg13g2_xnor2_1 _2111_ (.Y(_0108_),
    .A(\mb.b_0.ball_vy[2] ),
    .B(net255));
 sg13g2_o21ai_1 _2112_ (.B1(\mb.b_0.ball_vy[0] ),
    .Y(_0109_),
    .A1(\mb.b_0.ball_vy[1] ),
    .A2(net254));
 sg13g2_a21oi_1 _2113_ (.A1(_0105_),
    .A2(_0109_),
    .Y(_0110_),
    .B1(_0108_));
 sg13g2_nand3_1 _2114_ (.B(_0108_),
    .C(_0109_),
    .A(_0105_),
    .Y(_0111_));
 sg13g2_nor2b_1 _2115_ (.A(_0110_),
    .B_N(_0111_),
    .Y(_0011_));
 sg13g2_or2_1 _2116_ (.X(_0112_),
    .B(net255),
    .A(\mb.b_0.ball_vy[3] ));
 sg13g2_nand2_1 _2117_ (.Y(_0113_),
    .A(\mb.b_0.ball_vy[3] ),
    .B(net254));
 sg13g2_and2_1 _2118_ (.A(_0112_),
    .B(_0113_),
    .X(_0114_));
 sg13g2_nor2_1 _2119_ (.A(_0107_),
    .B(_0110_),
    .Y(_0115_));
 sg13g2_xnor2_1 _2120_ (.Y(_0012_),
    .A(_0114_),
    .B(_0115_));
 sg13g2_xor2_1 _2121_ (.B(net255),
    .A(\mb.b_0.ball_vy[4] ),
    .X(_0116_));
 sg13g2_inv_1 _2122_ (.Y(_0117_),
    .A(_0116_));
 sg13g2_o21ai_1 _2123_ (.B1(_0112_),
    .Y(_0118_),
    .A1(_0107_),
    .A2(_0110_));
 sg13g2_a21oi_1 _2124_ (.A1(_0113_),
    .A2(_0118_),
    .Y(_0119_),
    .B1(_0117_));
 sg13g2_nand3_1 _2125_ (.B(_0117_),
    .C(_0118_),
    .A(_0113_),
    .Y(_0120_));
 sg13g2_nor2b_1 _2126_ (.A(_0119_),
    .B_N(_0120_),
    .Y(_0013_));
 sg13g2_and2_1 _2127_ (.A(\mb.b_0.ball_vy[5] ),
    .B(net254),
    .X(_0121_));
 sg13g2_xor2_1 _2128_ (.B(net254),
    .A(\mb.b_0.ball_vy[5] ),
    .X(_0122_));
 sg13g2_a21oi_1 _2129_ (.A1(\mb.b_0.ball_vy[4] ),
    .A2(net254),
    .Y(_0123_),
    .B1(_0119_));
 sg13g2_xnor2_1 _2130_ (.Y(_0014_),
    .A(_0122_),
    .B(_0123_));
 sg13g2_xor2_1 _2131_ (.B(_0104_),
    .A(\mb.b_0.ball_vy[6] ),
    .X(_0124_));
 sg13g2_inv_1 _2132_ (.Y(_0125_),
    .A(_0124_));
 sg13g2_a221oi_1 _2133_ (.B2(_0122_),
    .C1(_0121_),
    .B1(_0119_),
    .A1(\mb.b_0.ball_vy[4] ),
    .Y(_0126_),
    .A2(net254));
 sg13g2_nor2_1 _2134_ (.A(_0125_),
    .B(_0126_),
    .Y(_0127_));
 sg13g2_xnor2_1 _2135_ (.Y(_0015_),
    .A(_0124_),
    .B(_0126_));
 sg13g2_xor2_1 _2136_ (.B(net256),
    .A(\mb.b_0.ball_vy[7] ),
    .X(_0128_));
 sg13g2_a21oi_1 _2137_ (.A1(\mb.b_0.ball_vy[6] ),
    .A2(net256),
    .Y(_0129_),
    .B1(_0127_));
 sg13g2_xnor2_1 _2138_ (.Y(_0016_),
    .A(_0128_),
    .B(_0129_));
 sg13g2_and2_1 _2139_ (.A(\mb.b_0.ball_vy[8] ),
    .B(net256),
    .X(_0130_));
 sg13g2_xor2_1 _2140_ (.B(net256),
    .A(\mb.b_0.ball_vy[8] ),
    .X(_0131_));
 sg13g2_nand2_1 _2141_ (.Y(_0132_),
    .A(_0124_),
    .B(_0128_));
 sg13g2_o21ai_1 _2142_ (.B1(net256),
    .Y(_0133_),
    .A1(\mb.b_0.ball_vy[6] ),
    .A2(\mb.b_0.ball_vy[7] ));
 sg13g2_o21ai_1 _2143_ (.B1(_0133_),
    .Y(_0134_),
    .A1(_0126_),
    .A2(_0132_));
 sg13g2_xor2_1 _2144_ (.B(_0134_),
    .A(_0131_),
    .X(_0017_));
 sg13g2_a21oi_1 _2145_ (.A1(_0131_),
    .A2(_0134_),
    .Y(_0135_),
    .B1(_0130_));
 sg13g2_xor2_1 _2146_ (.B(net256),
    .A(\mb.b_0.ball_vy[9] ),
    .X(_0136_));
 sg13g2_xnor2_1 _2147_ (.Y(_0018_),
    .A(_0135_),
    .B(_0136_));
 sg13g2_or2_1 _2148_ (.X(_0137_),
    .B(\mb.b_0.next_x[5] ),
    .A(\mb.b_0.next_x[4] ));
 sg13g2_a22oi_1 _2149_ (.Y(_0138_),
    .B1(_0137_),
    .B2(\mb.b_0.next_x[6] ),
    .A2(_1037_),
    .A1(_1036_));
 sg13g2_nor3_1 _2150_ (.A(_1040_),
    .B(_1042_),
    .C(_0138_),
    .Y(_0139_));
 sg13g2_nor3_1 _2151_ (.A(_1045_),
    .B(_1046_),
    .C(_0139_),
    .Y(_0140_));
 sg13g2_nand2_1 _2152_ (.Y(_0141_),
    .A(_0346_),
    .B(net253));
 sg13g2_xnor2_1 _2153_ (.Y(_0142_),
    .A(\mb.b_0.ball_vx[1] ),
    .B(net253));
 sg13g2_xnor2_1 _2154_ (.Y(_0001_),
    .A(_0038_),
    .B(_0142_));
 sg13g2_nor2b_1 _2155_ (.A(net253),
    .B_N(\mb.b_0.ball_vx[2] ),
    .Y(_0143_));
 sg13g2_xnor2_1 _2156_ (.Y(_0144_),
    .A(\mb.b_0.ball_vx[2] ),
    .B(net253));
 sg13g2_o21ai_1 _2157_ (.B1(_0329_),
    .Y(_0145_),
    .A1(_0346_),
    .A2(net253));
 sg13g2_and3_1 _2158_ (.X(_0146_),
    .A(_0141_),
    .B(_0144_),
    .C(_0145_));
 sg13g2_a21oi_1 _2159_ (.A1(_0141_),
    .A2(_0145_),
    .Y(_0147_),
    .B1(_0144_));
 sg13g2_nor2_1 _2160_ (.A(_0146_),
    .B(_0147_),
    .Y(_0002_));
 sg13g2_nor2b_1 _2161_ (.A(\mb.b_0.ball_vx[3] ),
    .B_N(net251),
    .Y(_0148_));
 sg13g2_nor2b_1 _2162_ (.A(net251),
    .B_N(\mb.b_0.ball_vx[3] ),
    .Y(_0149_));
 sg13g2_nor2_1 _2163_ (.A(_0148_),
    .B(_0149_),
    .Y(_0150_));
 sg13g2_nor2_1 _2164_ (.A(_0143_),
    .B(_0146_),
    .Y(_0151_));
 sg13g2_xnor2_1 _2165_ (.Y(_0003_),
    .A(_0150_),
    .B(_0151_));
 sg13g2_nand2b_1 _2166_ (.Y(_0152_),
    .B(\mb.b_0.ball_vx[4] ),
    .A_N(net252));
 sg13g2_inv_1 _2167_ (.Y(_0153_),
    .A(_0152_));
 sg13g2_xor2_1 _2168_ (.B(net251),
    .A(\mb.b_0.ball_vx[4] ),
    .X(_0154_));
 sg13g2_nor3_1 _2169_ (.A(_0143_),
    .B(_0146_),
    .C(_0149_),
    .Y(_0155_));
 sg13g2_nor2_1 _2170_ (.A(_0148_),
    .B(_0155_),
    .Y(_0156_));
 sg13g2_nand2b_1 _2171_ (.Y(_0157_),
    .B(_0156_),
    .A_N(_0154_));
 sg13g2_xnor2_1 _2172_ (.Y(_0004_),
    .A(_0154_),
    .B(_0156_));
 sg13g2_nor2b_1 _2173_ (.A(net251),
    .B_N(\mb.b_0.ball_vx[5] ),
    .Y(_0158_));
 sg13g2_xor2_1 _2174_ (.B(net251),
    .A(\mb.b_0.ball_vx[5] ),
    .X(_0159_));
 sg13g2_and2_1 _2175_ (.A(_0152_),
    .B(_0157_),
    .X(_0160_));
 sg13g2_xor2_1 _2176_ (.B(_0160_),
    .A(_0159_),
    .X(_0005_));
 sg13g2_nand2b_1 _2177_ (.Y(_0161_),
    .B(\mb.b_0.ball_vx[6] ),
    .A_N(net251));
 sg13g2_xnor2_1 _2178_ (.Y(_0162_),
    .A(\mb.b_0.ball_vx[6] ),
    .B(net251));
 sg13g2_nor4_1 _2179_ (.A(_0148_),
    .B(_0154_),
    .C(_0155_),
    .D(_0159_),
    .Y(_0163_));
 sg13g2_or3_1 _2180_ (.A(_0153_),
    .B(_0158_),
    .C(_0163_),
    .X(_0164_));
 sg13g2_nand2_1 _2181_ (.Y(_0165_),
    .A(_0162_),
    .B(_0164_));
 sg13g2_xor2_1 _2182_ (.B(_0164_),
    .A(_0162_),
    .X(_0006_));
 sg13g2_xnor2_1 _2183_ (.Y(_0166_),
    .A(\mb.b_0.ball_vx[7] ),
    .B(net252));
 sg13g2_nand2_1 _2184_ (.Y(_0167_),
    .A(_0161_),
    .B(_0165_));
 sg13g2_xor2_1 _2185_ (.B(_0167_),
    .A(_0166_),
    .X(_0007_));
 sg13g2_nor2b_1 _2186_ (.A(net252),
    .B_N(\mb.b_0.ball_vx[8] ),
    .Y(_0168_));
 sg13g2_xnor2_1 _2187_ (.Y(_0169_),
    .A(\mb.b_0.ball_vx[8] ),
    .B(net252));
 sg13g2_and2_1 _2188_ (.A(_0162_),
    .B(_0166_),
    .X(_0170_));
 sg13g2_o21ai_1 _2189_ (.B1(_0161_),
    .Y(_0171_),
    .A1(_0345_),
    .A2(net251));
 sg13g2_a21o_1 _2190_ (.A2(_0170_),
    .A1(_0164_),
    .B1(_0171_),
    .X(_0172_));
 sg13g2_xor2_1 _2191_ (.B(_0172_),
    .A(_0169_),
    .X(_0008_));
 sg13g2_a21oi_1 _2192_ (.A1(_0169_),
    .A2(_0172_),
    .Y(_0173_),
    .B1(_0168_));
 sg13g2_xnor2_1 _2193_ (.Y(_0174_),
    .A(\mb.b_0.ball_vx[9] ),
    .B(net252));
 sg13g2_xnor2_1 _2194_ (.Y(_0009_),
    .A(_0173_),
    .B(_0174_));
 sg13g2_a21o_1 _2195_ (.A2(\mb.b_1.next_y[3] ),
    .A1(\mb.b_1.next_y[2] ),
    .B1(\mb.b_1.next_y[4] ),
    .X(_0175_));
 sg13g2_and3_1 _2196_ (.X(_0176_),
    .A(\mb.b_1.next_y[6] ),
    .B(\mb.b_1.next_y[5] ),
    .C(_0175_));
 sg13g2_a22oi_1 _2197_ (.Y(_0177_),
    .B1(_0176_),
    .B2(\mb.b_1.next_y[7] ),
    .A2(_0084_),
    .A1(_0083_));
 sg13g2_nand3_1 _2198_ (.B(_0087_),
    .C(_0177_),
    .A(_0086_),
    .Y(_0178_));
 sg13g2_nand2_1 _2199_ (.Y(_0179_),
    .A(\mb.b_1.ball_vy[1] ),
    .B(net250));
 sg13g2_xor2_1 _2200_ (.B(net250),
    .A(\mb.b_1.ball_vy[1] ),
    .X(_0180_));
 sg13g2_xnor2_1 _2201_ (.Y(_0028_),
    .A(_0046_),
    .B(_0180_));
 sg13g2_and2_1 _2202_ (.A(\mb.b_1.ball_vy[2] ),
    .B(net250),
    .X(_0181_));
 sg13g2_xnor2_1 _2203_ (.Y(_0182_),
    .A(\mb.b_1.ball_vy[2] ),
    .B(net250));
 sg13g2_o21ai_1 _2204_ (.B1(\mb.b_1.ball_vy[0] ),
    .Y(_0183_),
    .A1(\mb.b_1.ball_vy[1] ),
    .A2(net250));
 sg13g2_a21oi_2 _2205_ (.B1(_0182_),
    .Y(_0184_),
    .A2(_0183_),
    .A1(_0179_));
 sg13g2_nand3_1 _2206_ (.B(_0182_),
    .C(_0183_),
    .A(_0179_),
    .Y(_0185_));
 sg13g2_nor2b_1 _2207_ (.A(_0184_),
    .B_N(_0185_),
    .Y(_0029_));
 sg13g2_nor2_1 _2208_ (.A(\mb.b_1.ball_vy[3] ),
    .B(net249),
    .Y(_0186_));
 sg13g2_and2_1 _2209_ (.A(\mb.b_1.ball_vy[3] ),
    .B(net249),
    .X(_0187_));
 sg13g2_nor2_1 _2210_ (.A(_0186_),
    .B(_0187_),
    .Y(_0188_));
 sg13g2_nor2_1 _2211_ (.A(_0181_),
    .B(_0184_),
    .Y(_0189_));
 sg13g2_xnor2_1 _2212_ (.Y(_0030_),
    .A(_0188_),
    .B(_0189_));
 sg13g2_and2_1 _2213_ (.A(\mb.b_1.ball_vy[4] ),
    .B(net249),
    .X(_0190_));
 sg13g2_xor2_1 _2214_ (.B(net249),
    .A(\mb.b_1.ball_vy[4] ),
    .X(_0191_));
 sg13g2_inv_1 _2215_ (.Y(_0192_),
    .A(_0191_));
 sg13g2_nor3_1 _2216_ (.A(_0181_),
    .B(_0184_),
    .C(_0187_),
    .Y(_0193_));
 sg13g2_nor2_1 _2217_ (.A(_0186_),
    .B(_0193_),
    .Y(_0194_));
 sg13g2_xnor2_1 _2218_ (.Y(_0031_),
    .A(_0192_),
    .B(_0194_));
 sg13g2_and2_1 _2219_ (.A(\mb.b_1.ball_vy[5] ),
    .B(_0178_),
    .X(_0195_));
 sg13g2_xnor2_1 _2220_ (.Y(_0196_),
    .A(\mb.b_1.ball_vy[5] ),
    .B(_0178_));
 sg13g2_a21oi_1 _2221_ (.A1(_0191_),
    .A2(_0194_),
    .Y(_0197_),
    .B1(_0190_));
 sg13g2_xor2_1 _2222_ (.B(_0197_),
    .A(_0196_),
    .X(_0032_));
 sg13g2_nand2_1 _2223_ (.Y(_0198_),
    .A(\mb.b_1.ball_vy[6] ),
    .B(net249));
 sg13g2_xor2_1 _2224_ (.B(net249),
    .A(\mb.b_1.ball_vy[6] ),
    .X(_0199_));
 sg13g2_inv_1 _2225_ (.Y(_0200_),
    .A(_0199_));
 sg13g2_nor4_1 _2226_ (.A(_0186_),
    .B(_0192_),
    .C(_0193_),
    .D(_0196_),
    .Y(_0201_));
 sg13g2_nor3_2 _2227_ (.A(_0190_),
    .B(_0195_),
    .C(_0201_),
    .Y(_0202_));
 sg13g2_xnor2_1 _2228_ (.Y(_0033_),
    .A(_0199_),
    .B(_0202_));
 sg13g2_xor2_1 _2229_ (.B(net249),
    .A(\mb.b_1.ball_vy[7] ),
    .X(_0203_));
 sg13g2_o21ai_1 _2230_ (.B1(_0198_),
    .Y(_0204_),
    .A1(_0200_),
    .A2(_0202_));
 sg13g2_xor2_1 _2231_ (.B(_0204_),
    .A(_0203_),
    .X(_0034_));
 sg13g2_and2_1 _2232_ (.A(\mb.b_1.ball_vy[8] ),
    .B(net250),
    .X(_0205_));
 sg13g2_xor2_1 _2233_ (.B(net250),
    .A(\mb.b_1.ball_vy[8] ),
    .X(_0206_));
 sg13g2_nand2_1 _2234_ (.Y(_0207_),
    .A(_0199_),
    .B(_0203_));
 sg13g2_o21ai_1 _2235_ (.B1(net249),
    .Y(_0208_),
    .A1(\mb.b_1.ball_vy[7] ),
    .A2(\mb.b_1.ball_vy[6] ));
 sg13g2_o21ai_1 _2236_ (.B1(_0208_),
    .Y(_0209_),
    .A1(_0202_),
    .A2(_0207_));
 sg13g2_xor2_1 _2237_ (.B(_0209_),
    .A(_0206_),
    .X(_0035_));
 sg13g2_a21oi_1 _2238_ (.A1(_0206_),
    .A2(_0209_),
    .Y(_0210_),
    .B1(_0205_));
 sg13g2_xor2_1 _2239_ (.B(net250),
    .A(\mb.b_1.ball_vy[9] ),
    .X(_0211_));
 sg13g2_xnor2_1 _2240_ (.Y(_0036_),
    .A(_0210_),
    .B(_0211_));
 sg13g2_or2_1 _2241_ (.X(_0212_),
    .B(\mb.b_1.next_x[5] ),
    .A(\mb.b_1.next_x[4] ));
 sg13g2_a22oi_1 _2242_ (.Y(_0213_),
    .B1(_0212_),
    .B2(\mb.b_1.next_x[6] ),
    .A2(_0092_),
    .A1(_0091_));
 sg13g2_nor3_1 _2243_ (.A(_0095_),
    .B(_0096_),
    .C(_0213_),
    .Y(_0214_));
 sg13g2_a21oi_2 _2244_ (.B1(_0214_),
    .Y(_0215_),
    .A2(_0100_),
    .A1(_0099_));
 sg13g2_nand2_1 _2245_ (.Y(_0216_),
    .A(_0347_),
    .B(net248));
 sg13g2_xnor2_1 _2246_ (.Y(_0217_),
    .A(\mb.b_1.ball_vx[1] ),
    .B(net248));
 sg13g2_xnor2_1 _2247_ (.Y(_0019_),
    .A(_0045_),
    .B(_0217_));
 sg13g2_nor2b_1 _2248_ (.A(net247),
    .B_N(\mb.b_1.ball_vx[2] ),
    .Y(_0218_));
 sg13g2_xnor2_1 _2249_ (.Y(_0219_),
    .A(\mb.b_1.ball_vx[2] ),
    .B(net247));
 sg13g2_o21ai_1 _2250_ (.B1(_0343_),
    .Y(_0220_),
    .A1(_0347_),
    .A2(net248));
 sg13g2_and3_1 _2251_ (.X(_0221_),
    .A(_0216_),
    .B(_0219_),
    .C(_0220_));
 sg13g2_a21oi_1 _2252_ (.A1(_0216_),
    .A2(_0220_),
    .Y(_0222_),
    .B1(_0219_));
 sg13g2_nor2_1 _2253_ (.A(_0221_),
    .B(_0222_),
    .Y(_0020_));
 sg13g2_nor2b_1 _2254_ (.A(\mb.b_1.ball_vx[3] ),
    .B_N(net247),
    .Y(_0223_));
 sg13g2_nor2b_1 _2255_ (.A(net247),
    .B_N(\mb.b_1.ball_vx[3] ),
    .Y(_0224_));
 sg13g2_nor2_1 _2256_ (.A(_0223_),
    .B(_0224_),
    .Y(_0225_));
 sg13g2_nor2_1 _2257_ (.A(_0218_),
    .B(_0221_),
    .Y(_0226_));
 sg13g2_xnor2_1 _2258_ (.Y(_0021_),
    .A(_0225_),
    .B(_0226_));
 sg13g2_nand2b_1 _2259_ (.Y(_0227_),
    .B(\mb.b_1.ball_vx[4] ),
    .A_N(net247));
 sg13g2_inv_1 _2260_ (.Y(_0228_),
    .A(_0227_));
 sg13g2_xor2_1 _2261_ (.B(net247),
    .A(\mb.b_1.ball_vx[4] ),
    .X(_0229_));
 sg13g2_nor3_1 _2262_ (.A(_0218_),
    .B(_0221_),
    .C(_0224_),
    .Y(_0230_));
 sg13g2_nor2_1 _2263_ (.A(_0223_),
    .B(_0230_),
    .Y(_0231_));
 sg13g2_nand2b_1 _2264_ (.Y(_0232_),
    .B(_0231_),
    .A_N(_0229_));
 sg13g2_xnor2_1 _2265_ (.Y(_0022_),
    .A(_0229_),
    .B(_0231_));
 sg13g2_nor2b_1 _2266_ (.A(net247),
    .B_N(\mb.b_1.ball_vx[5] ),
    .Y(_0233_));
 sg13g2_xor2_1 _2267_ (.B(net247),
    .A(\mb.b_1.ball_vx[5] ),
    .X(_0234_));
 sg13g2_and2_1 _2268_ (.A(_0227_),
    .B(_0232_),
    .X(_0235_));
 sg13g2_xor2_1 _2269_ (.B(_0235_),
    .A(_0234_),
    .X(_0023_));
 sg13g2_nand2b_1 _2270_ (.Y(_0236_),
    .B(\mb.b_1.ball_vx[6] ),
    .A_N(_0215_));
 sg13g2_xnor2_1 _2271_ (.Y(_0237_),
    .A(\mb.b_1.ball_vx[6] ),
    .B(_0215_));
 sg13g2_nor4_1 _2272_ (.A(_0223_),
    .B(_0229_),
    .C(_0230_),
    .D(_0234_),
    .Y(_0238_));
 sg13g2_or3_1 _2273_ (.A(_0228_),
    .B(_0233_),
    .C(_0238_),
    .X(_0239_));
 sg13g2_nand2_1 _2274_ (.Y(_0240_),
    .A(_0237_),
    .B(_0239_));
 sg13g2_xor2_1 _2275_ (.B(_0239_),
    .A(_0237_),
    .X(_0024_));
 sg13g2_xnor2_1 _2276_ (.Y(_0241_),
    .A(\mb.b_1.ball_vx[7] ),
    .B(net248));
 sg13g2_nand2_1 _2277_ (.Y(_0242_),
    .A(_0236_),
    .B(_0240_));
 sg13g2_xor2_1 _2278_ (.B(_0242_),
    .A(_0241_),
    .X(_0025_));
 sg13g2_nor2b_1 _2279_ (.A(net248),
    .B_N(\mb.b_1.ball_vx[8] ),
    .Y(_0243_));
 sg13g2_xnor2_1 _2280_ (.Y(_0244_),
    .A(\mb.b_1.ball_vx[8] ),
    .B(net248));
 sg13g2_and2_1 _2281_ (.A(_0237_),
    .B(_0241_),
    .X(_0245_));
 sg13g2_o21ai_1 _2282_ (.B1(_0236_),
    .Y(_0246_),
    .A1(_0344_),
    .A2(net248));
 sg13g2_a21o_1 _2283_ (.A2(_0245_),
    .A1(_0239_),
    .B1(_0246_),
    .X(_0247_));
 sg13g2_xor2_1 _2284_ (.B(_0247_),
    .A(_0244_),
    .X(_0026_));
 sg13g2_a21oi_1 _2285_ (.A1(_0244_),
    .A2(_0247_),
    .Y(_0248_),
    .B1(_0243_));
 sg13g2_xnor2_1 _2286_ (.Y(_0249_),
    .A(\mb.b_1.ball_vx[9] ),
    .B(net248));
 sg13g2_xnor2_1 _2287_ (.Y(_0027_),
    .A(_0248_),
    .B(_0249_));
 sg13g2_and3_1 _2288_ (.X(_0250_),
    .A(\mb.b_0.x[2] ),
    .B(\mb.b_0.x[1] ),
    .C(\mb.b_0.x[0] ));
 sg13g2_and2_2 _2289_ (.A(net326),
    .B(_0250_),
    .X(_0251_));
 sg13g2_nor2_1 _2290_ (.A(\mb.b_0.x[5] ),
    .B(net325),
    .Y(_0252_));
 sg13g2_and2_1 _2291_ (.A(_0251_),
    .B(_0252_),
    .X(_0253_));
 sg13g2_nor2_1 _2292_ (.A(\mb.b_0.x[6] ),
    .B(\mb.b_0.x[7] ),
    .Y(_0254_));
 sg13g2_nor2_1 _2293_ (.A(\mb.b_0.x[9] ),
    .B(\mb.b_0.x[8] ),
    .Y(_0255_));
 sg13g2_and4_1 _2294_ (.A(\v.h_counter[10] ),
    .B(_0253_),
    .C(_0254_),
    .D(_0255_),
    .X(_0256_));
 sg13g2_nor2b_2 _2295_ (.A(net303),
    .B_N(net328),
    .Y(_0257_));
 sg13g2_nand2b_2 _2296_ (.Y(_0258_),
    .B(net327),
    .A_N(net303));
 sg13g2_and2_1 _2297_ (.A(net124),
    .B(_0257_),
    .X(_0048_));
 sg13g2_xnor2_1 _2298_ (.Y(_0259_),
    .A(net147),
    .B(\mb.b_0.x[0] ));
 sg13g2_nor2_1 _2299_ (.A(_0258_),
    .B(net148),
    .Y(_0049_));
 sg13g2_a21oi_1 _2300_ (.A1(\mb.b_0.x[1] ),
    .A2(\mb.b_0.x[0] ),
    .Y(_0260_),
    .B1(net139));
 sg13g2_nor3_1 _2301_ (.A(_0250_),
    .B(_0258_),
    .C(net140),
    .Y(_0050_));
 sg13g2_o21ai_1 _2302_ (.B1(net1),
    .Y(_0261_),
    .A1(net326),
    .A2(_0250_));
 sg13g2_nor2_1 _2303_ (.A(_0251_),
    .B(_0261_),
    .Y(_0051_));
 sg13g2_xnor2_1 _2304_ (.Y(_0262_),
    .A(net325),
    .B(_0251_));
 sg13g2_nor2_1 _2305_ (.A(net302),
    .B(_0262_),
    .Y(_0052_));
 sg13g2_and3_1 _2306_ (.X(_0263_),
    .A(\mb.b_0.x[5] ),
    .B(net325),
    .C(_0251_));
 sg13g2_a21oi_1 _2307_ (.A1(net325),
    .A2(_0251_),
    .Y(_0264_),
    .B1(net141));
 sg13g2_nor3_1 _2308_ (.A(net302),
    .B(_0263_),
    .C(net142),
    .Y(_0053_));
 sg13g2_xnor2_1 _2309_ (.Y(_0265_),
    .A(net158),
    .B(_0263_));
 sg13g2_nor2_1 _2310_ (.A(net302),
    .B(_0265_),
    .Y(_0054_));
 sg13g2_a21oi_1 _2311_ (.A1(\mb.b_0.x[6] ),
    .A2(_0263_),
    .Y(_0266_),
    .B1(net130));
 sg13g2_and3_2 _2312_ (.X(_0267_),
    .A(\mb.b_0.x[6] ),
    .B(net130),
    .C(_0263_));
 sg13g2_nor3_1 _2313_ (.A(net302),
    .B(net131),
    .C(_0267_),
    .Y(_0055_));
 sg13g2_xor2_1 _2314_ (.B(_0267_),
    .A(net143),
    .X(_0268_));
 sg13g2_nor2_1 _2315_ (.A(net302),
    .B(_0268_),
    .Y(_0056_));
 sg13g2_a21oi_1 _2316_ (.A1(net144),
    .A2(_0267_),
    .Y(_0269_),
    .B1(\mb.b_0.x[9] ));
 sg13g2_nand3_1 _2317_ (.B(\mb.b_0.x[8] ),
    .C(_0267_),
    .A(\mb.b_0.x[9] ),
    .Y(_0270_));
 sg13g2_nand2_1 _2318_ (.Y(_0271_),
    .A(_0257_),
    .B(_0270_));
 sg13g2_nor2_1 _2319_ (.A(net145),
    .B(_0271_),
    .Y(_0057_));
 sg13g2_xor2_1 _2320_ (.B(_0270_),
    .A(net137),
    .X(_0272_));
 sg13g2_nor2_1 _2321_ (.A(net302),
    .B(net138),
    .Y(_0058_));
 sg13g2_nand2_1 _2322_ (.Y(_0273_),
    .A(\mb.b_0.y[9] ),
    .B(_0323_));
 sg13g2_nor3_1 _2323_ (.A(_0324_),
    .B(\mb.b_0.y[6] ),
    .C(_0273_),
    .Y(_0274_));
 sg13g2_nand2_1 _2324_ (.Y(_0275_),
    .A(_0326_),
    .B(net305));
 sg13g2_nand2_1 _2325_ (.Y(_0276_),
    .A(net307),
    .B(\mb.b_0.y[0] ));
 sg13g2_nor4_1 _2326_ (.A(net308),
    .B(\mb.b_0.y[1] ),
    .C(_0275_),
    .D(_0276_),
    .Y(_0277_));
 sg13g2_nand2_1 _2327_ (.Y(_0278_),
    .A(_0274_),
    .B(_0277_));
 sg13g2_a21oi_2 _2328_ (.B1(_0257_),
    .Y(_0279_),
    .A2(_0278_),
    .A1(net327));
 sg13g2_inv_1 _2329_ (.Y(_0280_),
    .A(_0279_));
 sg13g2_nand2b_1 _2330_ (.Y(_0281_),
    .B(net328),
    .A_N(net307));
 sg13g2_nand2_1 _2331_ (.Y(_0282_),
    .A(_0324_),
    .B(\mb.b_0.y[6] ));
 sg13g2_nor4_1 _2332_ (.A(_0273_),
    .B(_0275_),
    .C(_0281_),
    .D(_0282_),
    .Y(_0283_));
 sg13g2_and2_1 _2333_ (.A(net154),
    .B(net303),
    .X(_0284_));
 sg13g2_and2_1 _2334_ (.A(net152),
    .B(_0284_),
    .X(_0285_));
 sg13g2_and2_1 _2335_ (.A(net308),
    .B(_0285_),
    .X(_0286_));
 sg13g2_a22oi_1 _2336_ (.Y(_0059_),
    .B1(_0283_),
    .B2(_0286_),
    .A2(_0280_),
    .A1(_0328_));
 sg13g2_nor3_2 _2337_ (.A(_0335_),
    .B(_0336_),
    .C(\v.h_counter[10] ),
    .Y(_0287_));
 sg13g2_nor2b_1 _2338_ (.A(\mb.b_0.x[5] ),
    .B_N(net325),
    .Y(_0288_));
 sg13g2_and4_1 _2339_ (.A(net328),
    .B(_0254_),
    .C(_0287_),
    .D(_0288_),
    .X(_0289_));
 sg13g2_a22oi_1 _2340_ (.Y(_0060_),
    .B1(_0289_),
    .B2(_0251_),
    .A2(_0257_),
    .A1(_0327_));
 sg13g2_nor4_1 _2341_ (.A(net309),
    .B(\mb.b_0.y[0] ),
    .C(_0273_),
    .D(_0282_),
    .Y(_0290_));
 sg13g2_and4_1 _2342_ (.A(net126),
    .B(net305),
    .C(net307),
    .D(net308),
    .X(_0291_));
 sg13g2_nand3_1 _2343_ (.B(_0290_),
    .C(_0291_),
    .A(net303),
    .Y(_0292_));
 sg13g2_nand2_1 _2344_ (.Y(_0293_),
    .A(net321),
    .B(_0292_));
 sg13g2_nor2_1 _2345_ (.A(net307),
    .B(net308),
    .Y(_0294_));
 sg13g2_nand2_1 _2346_ (.Y(_0295_),
    .A(net309),
    .B(_0294_));
 sg13g2_nor4_1 _2347_ (.A(net126),
    .B(net305),
    .C(net155),
    .D(_0295_),
    .Y(_0296_));
 sg13g2_nand3_1 _2348_ (.B(_0274_),
    .C(_0296_),
    .A(net303),
    .Y(_0297_));
 sg13g2_nand3_1 _2349_ (.B(_0293_),
    .C(net156),
    .A(net328),
    .Y(_0061_));
 sg13g2_nand4_1 _2350_ (.B(net324),
    .C(_0253_),
    .A(\mb.b_0.x[6] ),
    .Y(_0298_),
    .D(_0287_));
 sg13g2_nor3_1 _2351_ (.A(_0330_),
    .B(net326),
    .C(net324),
    .Y(_0299_));
 sg13g2_nand4_1 _2352_ (.B(_0287_),
    .C(_0288_),
    .A(_0250_),
    .Y(_0300_),
    .D(_0299_));
 sg13g2_nand2_1 _2353_ (.Y(_0301_),
    .A(net132),
    .B(_0300_));
 sg13g2_nand3_1 _2354_ (.B(_0298_),
    .C(net133),
    .A(net1),
    .Y(_0062_));
 sg13g2_o21ai_1 _2355_ (.B1(net327),
    .Y(_0302_),
    .A1(net154),
    .A2(net303));
 sg13g2_nor2_1 _2356_ (.A(_0284_),
    .B(_0302_),
    .Y(_0063_));
 sg13g2_nor2_1 _2357_ (.A(net309),
    .B(_0284_),
    .Y(_0303_));
 sg13g2_nor3_1 _2358_ (.A(_0279_),
    .B(_0285_),
    .C(_0303_),
    .Y(_0064_));
 sg13g2_o21ai_1 _2359_ (.B1(net327),
    .Y(_0304_),
    .A1(net308),
    .A2(_0285_));
 sg13g2_nor2_1 _2360_ (.A(_0286_),
    .B(_0304_),
    .Y(_0065_));
 sg13g2_nor2_1 _2361_ (.A(net307),
    .B(_0286_),
    .Y(_0305_));
 sg13g2_and2_1 _2362_ (.A(net307),
    .B(_0286_),
    .X(_0306_));
 sg13g2_nor3_1 _2363_ (.A(_0279_),
    .B(_0305_),
    .C(_0306_),
    .Y(_0066_));
 sg13g2_o21ai_1 _2364_ (.B1(_0280_),
    .Y(_0307_),
    .A1(net305),
    .A2(_0306_));
 sg13g2_a21oi_1 _2365_ (.A1(net305),
    .A2(_0306_),
    .Y(_0067_),
    .B1(_0307_));
 sg13g2_a21oi_1 _2366_ (.A1(net305),
    .A2(_0306_),
    .Y(_0308_),
    .B1(net126));
 sg13g2_nand2_1 _2367_ (.Y(_0309_),
    .A(_0285_),
    .B(_0291_));
 sg13g2_nand2_1 _2368_ (.Y(_0310_),
    .A(net327),
    .B(_0309_));
 sg13g2_nor2_1 _2369_ (.A(net127),
    .B(_0310_),
    .Y(_0068_));
 sg13g2_and4_1 _2370_ (.A(\mb.b_0.y[6] ),
    .B(net309),
    .C(\mb.b_0.y[0] ),
    .D(_0291_),
    .X(_0311_));
 sg13g2_nand2b_1 _2371_ (.Y(_0312_),
    .B(net327),
    .A_N(_0311_));
 sg13g2_a22oi_1 _2372_ (.Y(_0069_),
    .B1(_0312_),
    .B2(net302),
    .A2(_0309_),
    .A1(_0325_));
 sg13g2_nand2b_1 _2373_ (.Y(_0313_),
    .B(net125),
    .A_N(_0256_));
 sg13g2_and2_1 _2374_ (.A(net303),
    .B(_0278_),
    .X(_0314_));
 sg13g2_and2_1 _2375_ (.A(net304),
    .B(_0311_),
    .X(_0315_));
 sg13g2_nand2b_1 _2376_ (.Y(_0316_),
    .B(_0314_),
    .A_N(_0315_));
 sg13g2_o21ai_1 _2377_ (.B1(net327),
    .Y(_0317_),
    .A1(net304),
    .A2(_0311_));
 sg13g2_a21oi_1 _2378_ (.A1(_0313_),
    .A2(_0316_),
    .Y(_0070_),
    .B1(_0317_));
 sg13g2_xnor2_1 _2379_ (.Y(_0318_),
    .A(_0040_),
    .B(_0315_));
 sg13g2_nand3_1 _2380_ (.B(_0314_),
    .C(_0318_),
    .A(net327),
    .Y(_0319_));
 sg13g2_o21ai_1 _2381_ (.B1(_0319_),
    .Y(_0071_),
    .A1(_0323_),
    .A2(net302));
 sg13g2_nand3_1 _2382_ (.B(net303),
    .C(_0315_),
    .A(net149),
    .Y(_0320_));
 sg13g2_xnor2_1 _2383_ (.Y(_0321_),
    .A(_0322_),
    .B(_0320_));
 sg13g2_nor2_1 _2384_ (.A(_0279_),
    .B(_0321_),
    .Y(_0072_));
 sg13g2_dfrbp_1 _2385_ (.CLK(net313),
    .RESET_B(net20),
    .D(\mb.b_1.next_x[0] ),
    .Q_N(_1125_),
    .Q(\mb.b_1.ball_x[0] ));
 sg13g2_dfrbp_1 _2386_ (.CLK(net313),
    .RESET_B(net21),
    .D(\mb.b_1.next_x[1] ),
    .Q_N(_1126_),
    .Q(\mb.b_1.ball_x[1] ));
 sg13g2_dfrbp_1 _2387_ (.CLK(net317),
    .RESET_B(net22),
    .D(\mb.b_1.next_x[2] ),
    .Q_N(_1127_),
    .Q(\mb.b_1.ball_x[2] ));
 sg13g2_dfrbp_1 _2388_ (.CLK(net315),
    .RESET_B(net23),
    .D(\mb.b_1.next_x[3] ),
    .Q_N(_1128_),
    .Q(\mb.b_1.ball_x[3] ));
 sg13g2_dfrbp_1 _2389_ (.CLK(net315),
    .RESET_B(net24),
    .D(\mb.b_1.next_x[4] ),
    .Q_N(_1129_),
    .Q(\mb.b_1.ball_x[4] ));
 sg13g2_dfrbp_1 _2390_ (.CLK(net315),
    .RESET_B(net25),
    .D(\mb.b_1.next_x[5] ),
    .Q_N(_1130_),
    .Q(\mb.b_1.ball_x[5] ));
 sg13g2_dfrbp_1 _2391_ (.CLK(net315),
    .RESET_B(net26),
    .D(\mb.b_1.next_x[6] ),
    .Q_N(_1131_),
    .Q(\mb.b_1.ball_x[6] ));
 sg13g2_dfrbp_1 _2392_ (.CLK(net315),
    .RESET_B(net27),
    .D(\mb.b_1.next_x[7] ),
    .Q_N(_1132_),
    .Q(\mb.b_1.ball_x[7] ));
 sg13g2_dfrbp_1 _2393_ (.CLK(net312),
    .RESET_B(net28),
    .D(\mb.b_1.next_x[8] ),
    .Q_N(_1133_),
    .Q(\mb.b_1.ball_x[8] ));
 sg13g2_dfrbp_1 _2394_ (.CLK(net315),
    .RESET_B(net29),
    .D(\mb.b_1.next_x[9] ),
    .Q_N(_0043_),
    .Q(\mb.b_1.ball_x[9] ));
 sg13g2_dfrbp_1 _2395_ (.CLK(net319),
    .RESET_B(net30),
    .D(\mb.b_1.next_y[0] ),
    .Q_N(_1134_),
    .Q(\mb.b_1.ball_y[0] ));
 sg13g2_dfrbp_1 _2396_ (.CLK(net320),
    .RESET_B(net31),
    .D(\mb.b_1.next_y[1] ),
    .Q_N(_1135_),
    .Q(\mb.b_1.ball_y[1] ));
 sg13g2_dfrbp_1 _2397_ (.CLK(net320),
    .RESET_B(net32),
    .D(\mb.b_1.next_y[2] ),
    .Q_N(_1136_),
    .Q(\mb.b_1.ball_y[2] ));
 sg13g2_dfrbp_1 _2398_ (.CLK(net320),
    .RESET_B(net33),
    .D(\mb.b_1.next_y[3] ),
    .Q_N(_1137_),
    .Q(\mb.b_1.ball_y[3] ));
 sg13g2_dfrbp_1 _2399_ (.CLK(net320),
    .RESET_B(net34),
    .D(\mb.b_1.next_y[4] ),
    .Q_N(_1138_),
    .Q(\mb.b_1.ball_y[4] ));
 sg13g2_dfrbp_1 _2400_ (.CLK(net320),
    .RESET_B(net35),
    .D(\mb.b_1.next_y[5] ),
    .Q_N(_1139_),
    .Q(\mb.b_1.ball_y[5] ));
 sg13g2_dfrbp_1 _2401_ (.CLK(net320),
    .RESET_B(net36),
    .D(\mb.b_1.next_y[6] ),
    .Q_N(_1140_),
    .Q(\mb.b_1.ball_y[6] ));
 sg13g2_dfrbp_1 _2402_ (.CLK(net318),
    .RESET_B(net37),
    .D(\mb.b_1.next_y[7] ),
    .Q_N(_1141_),
    .Q(\mb.b_1.ball_y[7] ));
 sg13g2_dfrbp_1 _2403_ (.CLK(net318),
    .RESET_B(net38),
    .D(\mb.b_1.next_y[8] ),
    .Q_N(_1142_),
    .Q(\mb.b_1.ball_y[8] ));
 sg13g2_dfrbp_1 _2404_ (.CLK(net319),
    .RESET_B(net39),
    .D(\mb.b_1.next_y[9] ),
    .Q_N(_0044_),
    .Q(\mb.b_1.ball_y[9] ));
 sg13g2_dfrbp_1 _2405_ (.CLK(net314),
    .RESET_B(net40),
    .D(_0045_),
    .Q_N(_0045_),
    .Q(\mb.b_1.ball_vx[0] ));
 sg13g2_dfrbp_1 _2406_ (.CLK(net314),
    .RESET_B(net41),
    .D(_0019_),
    .Q_N(_1143_),
    .Q(\mb.b_1.ball_vx[1] ));
 sg13g2_dfrbp_1 _2407_ (.CLK(net314),
    .RESET_B(net42),
    .D(_0020_),
    .Q_N(_1144_),
    .Q(\mb.b_1.ball_vx[2] ));
 sg13g2_dfrbp_1 _2408_ (.CLK(net313),
    .RESET_B(net43),
    .D(_0021_),
    .Q_N(_1145_),
    .Q(\mb.b_1.ball_vx[3] ));
 sg13g2_dfrbp_1 _2409_ (.CLK(net313),
    .RESET_B(net44),
    .D(_0022_),
    .Q_N(_1146_),
    .Q(\mb.b_1.ball_vx[4] ));
 sg13g2_dfrbp_1 _2410_ (.CLK(net314),
    .RESET_B(net45),
    .D(_0023_),
    .Q_N(_1147_),
    .Q(\mb.b_1.ball_vx[5] ));
 sg13g2_dfrbp_1 _2411_ (.CLK(net314),
    .RESET_B(net46),
    .D(_0024_),
    .Q_N(_1148_),
    .Q(\mb.b_1.ball_vx[6] ));
 sg13g2_dfrbp_1 _2412_ (.CLK(net314),
    .RESET_B(net47),
    .D(_0025_),
    .Q_N(_1149_),
    .Q(\mb.b_1.ball_vx[7] ));
 sg13g2_dfrbp_1 _2413_ (.CLK(net314),
    .RESET_B(net48),
    .D(_0026_),
    .Q_N(_1150_),
    .Q(\mb.b_1.ball_vx[8] ));
 sg13g2_dfrbp_1 _2414_ (.CLK(net312),
    .RESET_B(net49),
    .D(_0027_),
    .Q_N(_1151_),
    .Q(\mb.b_1.ball_vx[9] ));
 sg13g2_dfrbp_1 _2415_ (.CLK(net318),
    .RESET_B(net50),
    .D(_0046_),
    .Q_N(_0046_),
    .Q(\mb.b_1.ball_vy[0] ));
 sg13g2_dfrbp_1 _2416_ (.CLK(net318),
    .RESET_B(net51),
    .D(_0028_),
    .Q_N(_1152_),
    .Q(\mb.b_1.ball_vy[1] ));
 sg13g2_dfrbp_1 _2417_ (.CLK(net319),
    .RESET_B(net52),
    .D(_0029_),
    .Q_N(_1153_),
    .Q(\mb.b_1.ball_vy[2] ));
 sg13g2_dfrbp_1 _2418_ (.CLK(net320),
    .RESET_B(net53),
    .D(_0030_),
    .Q_N(_1154_),
    .Q(\mb.b_1.ball_vy[3] ));
 sg13g2_dfrbp_1 _2419_ (.CLK(net321),
    .RESET_B(net54),
    .D(_0031_),
    .Q_N(_1155_),
    .Q(\mb.b_1.ball_vy[4] ));
 sg13g2_dfrbp_1 _2420_ (.CLK(net321),
    .RESET_B(net55),
    .D(_0032_),
    .Q_N(_1156_),
    .Q(\mb.b_1.ball_vy[5] ));
 sg13g2_dfrbp_1 _2421_ (.CLK(net321),
    .RESET_B(net56),
    .D(_0033_),
    .Q_N(_1157_),
    .Q(\mb.b_1.ball_vy[6] ));
 sg13g2_dfrbp_1 _2422_ (.CLK(net320),
    .RESET_B(net57),
    .D(_0034_),
    .Q_N(_1158_),
    .Q(\mb.b_1.ball_vy[7] ));
 sg13g2_dfrbp_1 _2423_ (.CLK(net318),
    .RESET_B(net58),
    .D(_0035_),
    .Q_N(_1159_),
    .Q(\mb.b_1.ball_vy[8] ));
 sg13g2_dfrbp_1 _2424_ (.CLK(net318),
    .RESET_B(net59),
    .D(_0036_),
    .Q_N(_1160_),
    .Q(\mb.b_1.ball_vy[9] ));
 sg13g2_dfrbp_1 _2425_ (.CLK(net313),
    .RESET_B(net60),
    .D(\mb.b_0.next_x[0] ),
    .Q_N(_1161_),
    .Q(\mb.b_0.ball_x[0] ));
 sg13g2_dfrbp_1 _2426_ (.CLK(net317),
    .RESET_B(net61),
    .D(\mb.b_0.next_x[1] ),
    .Q_N(_1162_),
    .Q(\mb.b_0.ball_x[1] ));
 sg13g2_dfrbp_1 _2427_ (.CLK(net322),
    .RESET_B(net62),
    .D(\mb.b_0.next_x[2] ),
    .Q_N(_1163_),
    .Q(\mb.b_0.ball_x[2] ));
 sg13g2_dfrbp_1 _2428_ (.CLK(net322),
    .RESET_B(net63),
    .D(\mb.b_0.next_x[3] ),
    .Q_N(_1164_),
    .Q(\mb.b_0.ball_x[3] ));
 sg13g2_dfrbp_1 _2429_ (.CLK(net322),
    .RESET_B(net64),
    .D(\mb.b_0.next_x[4] ),
    .Q_N(_1165_),
    .Q(\mb.b_0.ball_x[4] ));
 sg13g2_dfrbp_1 _2430_ (.CLK(net322),
    .RESET_B(net65),
    .D(\mb.b_0.next_x[5] ),
    .Q_N(_1166_),
    .Q(\mb.b_0.ball_x[5] ));
 sg13g2_dfrbp_1 _2431_ (.CLK(net322),
    .RESET_B(net66),
    .D(\mb.b_0.next_x[6] ),
    .Q_N(_1167_),
    .Q(\mb.b_0.ball_x[6] ));
 sg13g2_dfrbp_1 _2432_ (.CLK(net315),
    .RESET_B(net67),
    .D(\mb.b_0.next_x[7] ),
    .Q_N(_1168_),
    .Q(\mb.b_0.ball_x[7] ));
 sg13g2_dfrbp_1 _2433_ (.CLK(net315),
    .RESET_B(net68),
    .D(\mb.b_0.next_x[8] ),
    .Q_N(_1169_),
    .Q(\mb.b_0.ball_x[8] ));
 sg13g2_dfrbp_1 _2434_ (.CLK(net316),
    .RESET_B(net69),
    .D(\mb.b_0.next_x[9] ),
    .Q_N(_0047_),
    .Q(\mb.b_0.ball_x[9] ));
 sg13g2_dfrbp_1 _2435_ (.CLK(net318),
    .RESET_B(net70),
    .D(\mb.b_0.next_y[0] ),
    .Q_N(_1170_),
    .Q(\mb.b_0.ball_y[0] ));
 sg13g2_dfrbp_1 _2436_ (.CLK(net318),
    .RESET_B(net71),
    .D(\mb.b_0.next_y[1] ),
    .Q_N(_1171_),
    .Q(\mb.b_0.ball_y[1] ));
 sg13g2_dfrbp_1 _2437_ (.CLK(net310),
    .RESET_B(net72),
    .D(\mb.b_0.next_y[2] ),
    .Q_N(_1077_),
    .Q(\mb.b_0.ball_y[2] ));
 sg13g2_dfrbp_1 _2438_ (.CLK(net310),
    .RESET_B(net73),
    .D(\mb.b_0.next_y[3] ),
    .Q_N(_1078_),
    .Q(\mb.b_0.ball_y[3] ));
 sg13g2_dfrbp_1 _2439_ (.CLK(net311),
    .RESET_B(net74),
    .D(\mb.b_0.next_y[4] ),
    .Q_N(_1079_),
    .Q(\mb.b_0.ball_y[4] ));
 sg13g2_dfrbp_1 _2440_ (.CLK(net311),
    .RESET_B(net75),
    .D(\mb.b_0.next_y[5] ),
    .Q_N(_1080_),
    .Q(\mb.b_0.ball_y[5] ));
 sg13g2_dfrbp_1 _2441_ (.CLK(net310),
    .RESET_B(net76),
    .D(\mb.b_0.next_y[6] ),
    .Q_N(_1081_),
    .Q(\mb.b_0.ball_y[6] ));
 sg13g2_dfrbp_1 _2442_ (.CLK(net311),
    .RESET_B(net77),
    .D(\mb.b_0.next_y[7] ),
    .Q_N(_1082_),
    .Q(\mb.b_0.ball_y[7] ));
 sg13g2_dfrbp_1 _2443_ (.CLK(net311),
    .RESET_B(net78),
    .D(\mb.b_0.next_y[8] ),
    .Q_N(_1083_),
    .Q(\mb.b_0.ball_y[8] ));
 sg13g2_dfrbp_1 _2444_ (.CLK(net311),
    .RESET_B(net79),
    .D(\mb.b_0.next_y[9] ),
    .Q_N(_0037_),
    .Q(\mb.b_0.ball_y[9] ));
 sg13g2_dfrbp_1 _2445_ (.CLK(net313),
    .RESET_B(net80),
    .D(_0038_),
    .Q_N(_0038_),
    .Q(\mb.b_0.ball_vx[0] ));
 sg13g2_dfrbp_1 _2446_ (.CLK(net313),
    .RESET_B(net81),
    .D(_0001_),
    .Q_N(_1084_),
    .Q(\mb.b_0.ball_vx[1] ));
 sg13g2_dfrbp_1 _2447_ (.CLK(net317),
    .RESET_B(net82),
    .D(_0002_),
    .Q_N(_1085_),
    .Q(\mb.b_0.ball_vx[2] ));
 sg13g2_dfrbp_1 _2448_ (.CLK(net313),
    .RESET_B(net83),
    .D(_0003_),
    .Q_N(_1086_),
    .Q(\mb.b_0.ball_vx[3] ));
 sg13g2_dfrbp_1 _2449_ (.CLK(net316),
    .RESET_B(net84),
    .D(_0004_),
    .Q_N(_1087_),
    .Q(\mb.b_0.ball_vx[4] ));
 sg13g2_dfrbp_1 _2450_ (.CLK(net316),
    .RESET_B(net85),
    .D(_0005_),
    .Q_N(_1088_),
    .Q(\mb.b_0.ball_vx[5] ));
 sg13g2_dfrbp_1 _2451_ (.CLK(net316),
    .RESET_B(net86),
    .D(_0006_),
    .Q_N(_1089_),
    .Q(\mb.b_0.ball_vx[6] ));
 sg13g2_dfrbp_1 _2452_ (.CLK(net316),
    .RESET_B(net87),
    .D(_0007_),
    .Q_N(_1090_),
    .Q(\mb.b_0.ball_vx[7] ));
 sg13g2_dfrbp_1 _2453_ (.CLK(net316),
    .RESET_B(net88),
    .D(_0008_),
    .Q_N(_1091_),
    .Q(\mb.b_0.ball_vx[8] ));
 sg13g2_dfrbp_1 _2454_ (.CLK(net316),
    .RESET_B(net89),
    .D(_0009_),
    .Q_N(_1092_),
    .Q(\mb.b_0.ball_vx[9] ));
 sg13g2_dfrbp_1 _2455_ (.CLK(net310),
    .RESET_B(net90),
    .D(_0039_),
    .Q_N(_0039_),
    .Q(\mb.b_0.ball_vy[0] ));
 sg13g2_dfrbp_1 _2456_ (.CLK(net310),
    .RESET_B(net91),
    .D(_0010_),
    .Q_N(_1093_),
    .Q(\mb.b_0.ball_vy[1] ));
 sg13g2_dfrbp_1 _2457_ (.CLK(net310),
    .RESET_B(net92),
    .D(_0011_),
    .Q_N(_1094_),
    .Q(\mb.b_0.ball_vy[2] ));
 sg13g2_dfrbp_1 _2458_ (.CLK(net310),
    .RESET_B(net93),
    .D(_0012_),
    .Q_N(_1095_),
    .Q(\mb.b_0.ball_vy[3] ));
 sg13g2_dfrbp_1 _2459_ (.CLK(net310),
    .RESET_B(net94),
    .D(_0013_),
    .Q_N(_1096_),
    .Q(\mb.b_0.ball_vy[4] ));
 sg13g2_dfrbp_1 _2460_ (.CLK(net312),
    .RESET_B(net95),
    .D(_0014_),
    .Q_N(_1097_),
    .Q(\mb.b_0.ball_vy[5] ));
 sg13g2_dfrbp_1 _2461_ (.CLK(net312),
    .RESET_B(net96),
    .D(_0015_),
    .Q_N(_1098_),
    .Q(\mb.b_0.ball_vy[6] ));
 sg13g2_dfrbp_1 _2462_ (.CLK(net312),
    .RESET_B(net97),
    .D(_0016_),
    .Q_N(_1099_),
    .Q(\mb.b_0.ball_vy[7] ));
 sg13g2_dfrbp_1 _2463_ (.CLK(net312),
    .RESET_B(net98),
    .D(_0017_),
    .Q_N(_1100_),
    .Q(\mb.b_0.ball_vy[8] ));
 sg13g2_dfrbp_1 _2464_ (.CLK(net312),
    .RESET_B(net99),
    .D(_0018_),
    .Q_N(_1101_),
    .Q(\mb.b_0.ball_vy[9] ));
 sg13g2_dfrbp_1 _2465_ (.CLK(\mb.b_0.x[0] ),
    .RESET_B(net19),
    .D(_0000_),
    .Q_N(_1124_),
    .Q(\mb.pix ));
 sg13g2_dfrbp_1 _2466_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net123),
    .D(_0048_),
    .Q_N(_0042_),
    .Q(\mb.b_0.x[0] ));
 sg13g2_dfrbp_1 _2467_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net122),
    .D(_0049_),
    .Q_N(_1123_),
    .Q(\mb.b_0.x[1] ));
 sg13g2_dfrbp_1 _2468_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net121),
    .D(_0050_),
    .Q_N(_1122_),
    .Q(\mb.b_0.x[2] ));
 sg13g2_dfrbp_1 _2469_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net120),
    .D(_0051_),
    .Q_N(_1121_),
    .Q(\mb.b_0.x[3] ));
 sg13g2_dfrbp_1 _2470_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net119),
    .D(_0052_),
    .Q_N(_1120_),
    .Q(\mb.b_0.x[4] ));
 sg13g2_dfrbp_1 _2471_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net118),
    .D(_0053_),
    .Q_N(_1119_),
    .Q(\mb.b_0.x[5] ));
 sg13g2_dfrbp_1 _2472_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net117),
    .D(_0054_),
    .Q_N(_1118_),
    .Q(\mb.b_0.x[6] ));
 sg13g2_dfrbp_1 _2473_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net116),
    .D(_0055_),
    .Q_N(_1117_),
    .Q(\mb.b_0.x[7] ));
 sg13g2_dfrbp_1 _2474_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net115),
    .D(_0056_),
    .Q_N(_0041_),
    .Q(\mb.b_0.x[8] ));
 sg13g2_dfrbp_1 _2475_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net114),
    .D(net146),
    .Q_N(_1116_),
    .Q(\mb.b_0.x[9] ));
 sg13g2_dfrbp_1 _2476_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net113),
    .D(_0058_),
    .Q_N(_1115_),
    .Q(\v.h_counter[10] ));
 sg13g2_dfrbp_1 _2477_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net112),
    .D(net136),
    .Q_N(_1114_),
    .Q(\v.v_display ));
 sg13g2_dfrbp_1 _2478_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net110),
    .D(net129),
    .Q_N(_1113_),
    .Q(\v.h_display ));
 sg13g2_dfrbp_1 _2479_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net108),
    .D(_0061_),
    .Q_N(_1112_),
    .Q(\mb.b_0.v_sync ));
 sg13g2_dfrbp_1 _2480_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net106),
    .D(net134),
    .Q_N(_1111_),
    .Q(h_sync));
 sg13g2_dfrbp_1 _2481_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net104),
    .D(_0063_),
    .Q_N(_1110_),
    .Q(\mb.b_0.y[0] ));
 sg13g2_dfrbp_1 _2482_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net102),
    .D(net153),
    .Q_N(_1109_),
    .Q(\mb.b_0.y[1] ));
 sg13g2_dfrbp_1 _2483_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net100),
    .D(_0065_),
    .Q_N(_1108_),
    .Q(\mb.b_0.y[2] ));
 sg13g2_dfrbp_1 _2484_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net18),
    .D(_0066_),
    .Q_N(_1107_),
    .Q(\mb.b_0.y[3] ));
 sg13g2_dfrbp_1 _2485_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net109),
    .D(_0067_),
    .Q_N(_1106_),
    .Q(\mb.b_0.y[4] ));
 sg13g2_dfrbp_1 _2486_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net105),
    .D(_0068_),
    .Q_N(_1105_),
    .Q(\mb.b_0.y[5] ));
 sg13g2_dfrbp_1 _2487_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net101),
    .D(_0069_),
    .Q_N(_1104_),
    .Q(\mb.b_0.y[6] ));
 sg13g2_dfrbp_1 _2488_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net111),
    .D(_0070_),
    .Q_N(_1103_),
    .Q(\mb.b_0.y[7] ));
 sg13g2_dfrbp_1 _2489_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net103),
    .D(net150),
    .Q_N(_0040_),
    .Q(\mb.b_0.y[8] ));
 sg13g2_dfrbp_1 _2490_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net107),
    .D(_0072_),
    .Q_N(_1102_),
    .Q(\mb.b_0.y[9] ));
 sg13g2_tiehi _2465__19 (.L_HI(net19));
 sg13g2_tiehi _2385__20 (.L_HI(net20));
 sg13g2_tiehi _2386__21 (.L_HI(net21));
 sg13g2_tiehi _2387__22 (.L_HI(net22));
 sg13g2_tiehi _2388__23 (.L_HI(net23));
 sg13g2_tiehi _2389__24 (.L_HI(net24));
 sg13g2_tiehi _2390__25 (.L_HI(net25));
 sg13g2_tiehi _2391__26 (.L_HI(net26));
 sg13g2_tiehi _2392__27 (.L_HI(net27));
 sg13g2_tiehi _2393__28 (.L_HI(net28));
 sg13g2_tiehi _2394__29 (.L_HI(net29));
 sg13g2_tiehi _2395__30 (.L_HI(net30));
 sg13g2_tiehi _2396__31 (.L_HI(net31));
 sg13g2_tiehi _2397__32 (.L_HI(net32));
 sg13g2_tiehi _2398__33 (.L_HI(net33));
 sg13g2_tiehi _2399__34 (.L_HI(net34));
 sg13g2_tiehi _2400__35 (.L_HI(net35));
 sg13g2_tiehi _2401__36 (.L_HI(net36));
 sg13g2_tiehi _2402__37 (.L_HI(net37));
 sg13g2_tiehi _2403__38 (.L_HI(net38));
 sg13g2_tiehi _2404__39 (.L_HI(net39));
 sg13g2_tiehi _2405__40 (.L_HI(net40));
 sg13g2_tiehi _2406__41 (.L_HI(net41));
 sg13g2_tiehi _2407__42 (.L_HI(net42));
 sg13g2_tiehi _2408__43 (.L_HI(net43));
 sg13g2_tiehi _2409__44 (.L_HI(net44));
 sg13g2_tiehi _2410__45 (.L_HI(net45));
 sg13g2_tiehi _2411__46 (.L_HI(net46));
 sg13g2_tiehi _2412__47 (.L_HI(net47));
 sg13g2_tiehi _2413__48 (.L_HI(net48));
 sg13g2_tiehi _2414__49 (.L_HI(net49));
 sg13g2_tiehi _2415__50 (.L_HI(net50));
 sg13g2_tiehi _2416__51 (.L_HI(net51));
 sg13g2_tiehi _2417__52 (.L_HI(net52));
 sg13g2_tiehi _2418__53 (.L_HI(net53));
 sg13g2_tiehi _2419__54 (.L_HI(net54));
 sg13g2_tiehi _2420__55 (.L_HI(net55));
 sg13g2_tiehi _2421__56 (.L_HI(net56));
 sg13g2_tiehi _2422__57 (.L_HI(net57));
 sg13g2_tiehi _2423__58 (.L_HI(net58));
 sg13g2_tiehi _2424__59 (.L_HI(net59));
 sg13g2_tiehi _2425__60 (.L_HI(net60));
 sg13g2_tiehi _2426__61 (.L_HI(net61));
 sg13g2_tiehi _2427__62 (.L_HI(net62));
 sg13g2_tiehi _2428__63 (.L_HI(net63));
 sg13g2_tiehi _2429__64 (.L_HI(net64));
 sg13g2_tiehi _2430__65 (.L_HI(net65));
 sg13g2_tiehi _2431__66 (.L_HI(net66));
 sg13g2_tiehi _2432__67 (.L_HI(net67));
 sg13g2_tiehi _2433__68 (.L_HI(net68));
 sg13g2_tiehi _2434__69 (.L_HI(net69));
 sg13g2_tiehi _2435__70 (.L_HI(net70));
 sg13g2_tiehi _2436__71 (.L_HI(net71));
 sg13g2_tiehi _2437__72 (.L_HI(net72));
 sg13g2_tiehi _2438__73 (.L_HI(net73));
 sg13g2_tiehi _2439__74 (.L_HI(net74));
 sg13g2_tiehi _2440__75 (.L_HI(net75));
 sg13g2_tiehi _2441__76 (.L_HI(net76));
 sg13g2_tiehi _2442__77 (.L_HI(net77));
 sg13g2_tiehi _2443__78 (.L_HI(net78));
 sg13g2_tiehi _2444__79 (.L_HI(net79));
 sg13g2_tiehi _2445__80 (.L_HI(net80));
 sg13g2_tiehi _2446__81 (.L_HI(net81));
 sg13g2_tiehi _2447__82 (.L_HI(net82));
 sg13g2_tiehi _2448__83 (.L_HI(net83));
 sg13g2_tiehi _2449__84 (.L_HI(net84));
 sg13g2_tiehi _2450__85 (.L_HI(net85));
 sg13g2_tiehi _2451__86 (.L_HI(net86));
 sg13g2_tiehi _2452__87 (.L_HI(net87));
 sg13g2_tiehi _2453__88 (.L_HI(net88));
 sg13g2_tiehi _2454__89 (.L_HI(net89));
 sg13g2_tiehi _2455__90 (.L_HI(net90));
 sg13g2_tiehi _2456__91 (.L_HI(net91));
 sg13g2_tiehi _2457__92 (.L_HI(net92));
 sg13g2_tiehi _2458__93 (.L_HI(net93));
 sg13g2_tiehi _2459__94 (.L_HI(net94));
 sg13g2_tiehi _2460__95 (.L_HI(net95));
 sg13g2_tiehi _2461__96 (.L_HI(net96));
 sg13g2_tiehi _2462__97 (.L_HI(net97));
 sg13g2_tiehi _2463__98 (.L_HI(net98));
 sg13g2_tiehi _2464__99 (.L_HI(net99));
 sg13g2_tiehi _2483__100 (.L_HI(net100));
 sg13g2_tiehi _2487__101 (.L_HI(net101));
 sg13g2_tiehi _2482__102 (.L_HI(net102));
 sg13g2_tiehi _2489__103 (.L_HI(net103));
 sg13g2_tiehi _2481__104 (.L_HI(net104));
 sg13g2_tiehi _2486__105 (.L_HI(net105));
 sg13g2_tiehi _2480__106 (.L_HI(net106));
 sg13g2_tiehi _2490__107 (.L_HI(net107));
 sg13g2_tiehi _2479__108 (.L_HI(net108));
 sg13g2_tiehi _2485__109 (.L_HI(net109));
 sg13g2_tiehi _2478__110 (.L_HI(net110));
 sg13g2_tiehi _2488__111 (.L_HI(net111));
 sg13g2_tiehi _2477__112 (.L_HI(net112));
 sg13g2_tiehi _2476__113 (.L_HI(net113));
 sg13g2_tiehi _2475__114 (.L_HI(net114));
 sg13g2_tiehi _2474__115 (.L_HI(net115));
 sg13g2_tiehi _2473__116 (.L_HI(net116));
 sg13g2_tiehi _2472__117 (.L_HI(net117));
 sg13g2_tiehi _2471__118 (.L_HI(net118));
 sg13g2_tiehi _2470__119 (.L_HI(net119));
 sg13g2_tiehi _2469__120 (.L_HI(net120));
 sg13g2_tiehi _2468__121 (.L_HI(net121));
 sg13g2_tiehi _2467__122 (.L_HI(net122));
 sg13g2_tiehi _2466__123 (.L_HI(net123));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_johshoff_metaballs_3 (.L_LO(net3));
 sg13g2_tielo tt_um_johshoff_metaballs_4 (.L_LO(net4));
 sg13g2_tielo tt_um_johshoff_metaballs_5 (.L_LO(net5));
 sg13g2_tielo tt_um_johshoff_metaballs_6 (.L_LO(net6));
 sg13g2_tielo tt_um_johshoff_metaballs_7 (.L_LO(net7));
 sg13g2_tielo tt_um_johshoff_metaballs_8 (.L_LO(net8));
 sg13g2_tielo tt_um_johshoff_metaballs_9 (.L_LO(net9));
 sg13g2_tielo tt_um_johshoff_metaballs_10 (.L_LO(net10));
 sg13g2_tielo tt_um_johshoff_metaballs_11 (.L_LO(net11));
 sg13g2_tielo tt_um_johshoff_metaballs_12 (.L_LO(net12));
 sg13g2_tielo tt_um_johshoff_metaballs_13 (.L_LO(net13));
 sg13g2_tielo tt_um_johshoff_metaballs_14 (.L_LO(net14));
 sg13g2_tielo tt_um_johshoff_metaballs_15 (.L_LO(net15));
 sg13g2_tielo tt_um_johshoff_metaballs_16 (.L_LO(net16));
 sg13g2_tielo tt_um_johshoff_metaballs_17 (.L_LO(net17));
 sg13g2_tiehi _2484__18 (.L_HI(net18));
 sg13g2_buf_2 _2613_ (.A(\mb.rgb ),
    .X(uo_out[0]));
 sg13g2_buf_2 _2614_ (.A(\mb.rgb ),
    .X(uo_out[1]));
 sg13g2_buf_2 _2615_ (.A(\mb.rgb ),
    .X(uo_out[2]));
 sg13g2_buf_1 _2616_ (.A(net322),
    .X(uo_out[3]));
 sg13g2_buf_2 _2617_ (.A(\mb.rgb ),
    .X(uo_out[4]));
 sg13g2_buf_2 _2618_ (.A(\mb.rgb ),
    .X(uo_out[5]));
 sg13g2_buf_2 _2619_ (.A(\mb.rgb ),
    .X(uo_out[6]));
 sg13g2_buf_1 _2620_ (.A(h_sync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout247 (.A(_0215_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_0215_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_0178_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_0178_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(net252),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(net253),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_0140_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(net256),
    .X(net254));
 sg13g2_buf_1 fanout255 (.A(net256),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_0104_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_0475_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_0426_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_0711_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_0711_),
    .X(net260));
 sg13g2_buf_4 fanout261 (.X(net261),
    .A(net262));
 sg13g2_buf_1 fanout262 (.A(_0705_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_0705_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_0704_),
    .X(net264));
 sg13g2_buf_4 fanout265 (.X(net265),
    .A(_0704_));
 sg13g2_buf_2 fanout266 (.A(_0700_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_0700_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_0699_),
    .X(net268));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(net270));
 sg13g2_buf_2 fanout270 (.A(_0697_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_0696_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_0688_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(net274),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_0687_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_0681_),
    .X(net275));
 sg13g2_buf_4 fanout276 (.X(net276),
    .A(_0440_));
 sg13g2_buf_2 fanout277 (.A(_0440_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(net279),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_0430_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_0429_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_0413_),
    .X(net281));
 sg13g2_buf_4 fanout282 (.X(net282),
    .A(_0412_));
 sg13g2_buf_4 fanout283 (.X(net283),
    .A(_0412_));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(_0406_));
 sg13g2_buf_4 fanout285 (.X(net285),
    .A(_0405_));
 sg13g2_buf_2 fanout286 (.A(_0405_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_0377_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(net289),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_0685_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_0684_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_0684_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(net293),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_0684_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(net297),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(net296),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(net297),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_0421_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(net301),
    .X(net298));
 sg13g2_buf_1 fanout299 (.A(net301),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(net301),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_0420_),
    .X(net301));
 sg13g2_buf_4 fanout302 (.X(net302),
    .A(_0258_));
 sg13g2_buf_2 fanout303 (.A(_0256_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(net125),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(net151),
    .X(net305));
 sg13g2_buf_1 fanout306 (.A(\mb.b_0.y[4] ),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(net159),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(net160),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(net152),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(net323),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(net312),
    .X(net311));
 sg13g2_buf_4 fanout312 (.X(net312),
    .A(net323));
 sg13g2_buf_2 fanout313 (.A(net314),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(net317),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(net316),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(net317),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(net323),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(net319),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(net322),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(net321),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(net322),
    .X(net321));
 sg13g2_buf_4 fanout322 (.X(net322),
    .A(net323));
 sg13g2_buf_2 fanout323 (.A(\mb.b_0.v_sync ),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(net130),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(net162),
    .X(net325));
 sg13g2_buf_4 fanout326 (.X(net326),
    .A(net161));
 sg13g2_buf_4 fanout327 (.X(net327),
    .A(net328));
 sg13g2_buf_2 fanout328 (.A(net1),
    .X(net328));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_tielo tt_um_johshoff_metaballs_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_2_2__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0042_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold2 (.A(\mb.b_0.y[7] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold3 (.A(\mb.b_0.y[5] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0308_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold5 (.A(\v.h_display ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0060_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold7 (.A(\mb.b_0.x[7] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0266_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold9 (.A(h_sync),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0301_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0062_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold12 (.A(\v.v_display ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0059_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold14 (.A(\v.h_counter[10] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0272_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold16 (.A(\mb.b_0.x[2] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0260_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold18 (.A(\mb.b_0.x[5] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0264_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0041_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold21 (.A(\mb.b_0.x[8] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0269_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0057_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold24 (.A(\mb.b_0.x[1] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0259_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold26 (.A(\mb.b_0.y[8] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0071_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold28 (.A(\mb.b_0.y[4] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold29 (.A(\mb.b_0.y[1] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0064_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold31 (.A(\mb.b_0.y[0] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold32 (.A(\mb.b_0.y[0] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0297_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold34 (.A(\mb.b_0.y[6] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold35 (.A(\mb.b_0.x[6] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold36 (.A(\mb.b_0.y[3] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold37 (.A(\mb.b_0.y[2] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold38 (.A(\mb.b_0.x[3] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold39 (.A(\mb.b_0.x[4] ),
    .X(net162));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_4 FILLER_0_210 ();
 sg13g2_fill_1 FILLER_0_214 ();
 sg13g2_decap_4 FILLER_0_224 ();
 sg13g2_decap_4 FILLER_0_232 ();
 sg13g2_fill_2 FILLER_0_236 ();
 sg13g2_decap_4 FILLER_0_247 ();
 sg13g2_fill_2 FILLER_0_251 ();
 sg13g2_decap_4 FILLER_0_265 ();
 sg13g2_decap_8 FILLER_0_295 ();
 sg13g2_decap_8 FILLER_0_302 ();
 sg13g2_decap_8 FILLER_0_309 ();
 sg13g2_decap_8 FILLER_0_316 ();
 sg13g2_decap_8 FILLER_0_323 ();
 sg13g2_decap_8 FILLER_0_330 ();
 sg13g2_decap_8 FILLER_0_337 ();
 sg13g2_decap_8 FILLER_0_344 ();
 sg13g2_decap_8 FILLER_0_351 ();
 sg13g2_decap_8 FILLER_0_358 ();
 sg13g2_decap_8 FILLER_0_365 ();
 sg13g2_decap_8 FILLER_0_372 ();
 sg13g2_decap_8 FILLER_0_379 ();
 sg13g2_decap_8 FILLER_0_386 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_decap_8 FILLER_0_400 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_fill_2 FILLER_1_203 ();
 sg13g2_fill_1 FILLER_1_243 ();
 sg13g2_decap_4 FILLER_1_276 ();
 sg13g2_decap_8 FILLER_1_284 ();
 sg13g2_fill_1 FILLER_1_291 ();
 sg13g2_decap_8 FILLER_1_307 ();
 sg13g2_decap_8 FILLER_1_314 ();
 sg13g2_fill_1 FILLER_1_321 ();
 sg13g2_decap_8 FILLER_1_326 ();
 sg13g2_decap_8 FILLER_1_333 ();
 sg13g2_decap_8 FILLER_1_340 ();
 sg13g2_decap_8 FILLER_1_347 ();
 sg13g2_decap_8 FILLER_1_354 ();
 sg13g2_decap_8 FILLER_1_361 ();
 sg13g2_decap_8 FILLER_1_368 ();
 sg13g2_decap_8 FILLER_1_375 ();
 sg13g2_decap_8 FILLER_1_382 ();
 sg13g2_decap_8 FILLER_1_389 ();
 sg13g2_decap_8 FILLER_1_396 ();
 sg13g2_decap_4 FILLER_1_403 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_4 FILLER_2_154 ();
 sg13g2_fill_1 FILLER_2_163 ();
 sg13g2_decap_4 FILLER_2_174 ();
 sg13g2_fill_2 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_192 ();
 sg13g2_decap_4 FILLER_2_199 ();
 sg13g2_fill_2 FILLER_2_203 ();
 sg13g2_fill_2 FILLER_2_213 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_4 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_248 ();
 sg13g2_fill_2 FILLER_2_293 ();
 sg13g2_fill_2 FILLER_2_308 ();
 sg13g2_fill_1 FILLER_2_310 ();
 sg13g2_decap_8 FILLER_2_337 ();
 sg13g2_decap_8 FILLER_2_344 ();
 sg13g2_decap_8 FILLER_2_351 ();
 sg13g2_decap_8 FILLER_2_358 ();
 sg13g2_decap_8 FILLER_2_365 ();
 sg13g2_decap_8 FILLER_2_372 ();
 sg13g2_decap_8 FILLER_2_379 ();
 sg13g2_decap_8 FILLER_2_386 ();
 sg13g2_decap_8 FILLER_2_393 ();
 sg13g2_decap_8 FILLER_2_400 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_fill_2 FILLER_3_119 ();
 sg13g2_decap_4 FILLER_3_147 ();
 sg13g2_fill_1 FILLER_3_220 ();
 sg13g2_decap_8 FILLER_3_237 ();
 sg13g2_decap_4 FILLER_3_244 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_4 FILLER_3_273 ();
 sg13g2_fill_1 FILLER_3_277 ();
 sg13g2_decap_8 FILLER_3_282 ();
 sg13g2_decap_8 FILLER_3_339 ();
 sg13g2_decap_8 FILLER_3_346 ();
 sg13g2_decap_8 FILLER_3_353 ();
 sg13g2_decap_8 FILLER_3_360 ();
 sg13g2_decap_8 FILLER_3_367 ();
 sg13g2_decap_8 FILLER_3_374 ();
 sg13g2_decap_8 FILLER_3_381 ();
 sg13g2_decap_8 FILLER_3_388 ();
 sg13g2_decap_8 FILLER_3_395 ();
 sg13g2_decap_8 FILLER_3_402 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_fill_2 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_170 ();
 sg13g2_decap_8 FILLER_4_177 ();
 sg13g2_fill_2 FILLER_4_197 ();
 sg13g2_fill_1 FILLER_4_199 ();
 sg13g2_decap_8 FILLER_4_209 ();
 sg13g2_fill_2 FILLER_4_216 ();
 sg13g2_fill_1 FILLER_4_218 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_fill_2 FILLER_4_252 ();
 sg13g2_fill_1 FILLER_4_254 ();
 sg13g2_decap_4 FILLER_4_289 ();
 sg13g2_fill_1 FILLER_4_293 ();
 sg13g2_fill_1 FILLER_4_303 ();
 sg13g2_decap_8 FILLER_4_311 ();
 sg13g2_decap_4 FILLER_4_318 ();
 sg13g2_decap_8 FILLER_4_330 ();
 sg13g2_decap_8 FILLER_4_337 ();
 sg13g2_decap_8 FILLER_4_344 ();
 sg13g2_decap_8 FILLER_4_351 ();
 sg13g2_decap_8 FILLER_4_358 ();
 sg13g2_decap_8 FILLER_4_365 ();
 sg13g2_decap_8 FILLER_4_372 ();
 sg13g2_decap_8 FILLER_4_379 ();
 sg13g2_decap_8 FILLER_4_386 ();
 sg13g2_decap_8 FILLER_4_393 ();
 sg13g2_decap_8 FILLER_4_400 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_fill_1 FILLER_5_54 ();
 sg13g2_decap_8 FILLER_5_74 ();
 sg13g2_decap_4 FILLER_5_81 ();
 sg13g2_fill_1 FILLER_5_85 ();
 sg13g2_decap_8 FILLER_5_90 ();
 sg13g2_decap_8 FILLER_5_97 ();
 sg13g2_decap_8 FILLER_5_104 ();
 sg13g2_decap_8 FILLER_5_111 ();
 sg13g2_decap_8 FILLER_5_118 ();
 sg13g2_fill_2 FILLER_5_125 ();
 sg13g2_fill_1 FILLER_5_131 ();
 sg13g2_decap_8 FILLER_5_136 ();
 sg13g2_decap_4 FILLER_5_143 ();
 sg13g2_decap_8 FILLER_5_151 ();
 sg13g2_decap_4 FILLER_5_158 ();
 sg13g2_fill_2 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_214 ();
 sg13g2_decap_4 FILLER_5_225 ();
 sg13g2_fill_1 FILLER_5_229 ();
 sg13g2_decap_8 FILLER_5_234 ();
 sg13g2_fill_2 FILLER_5_241 ();
 sg13g2_fill_1 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_278 ();
 sg13g2_fill_2 FILLER_5_285 ();
 sg13g2_decap_4 FILLER_5_305 ();
 sg13g2_fill_2 FILLER_5_309 ();
 sg13g2_decap_8 FILLER_5_337 ();
 sg13g2_decap_8 FILLER_5_344 ();
 sg13g2_decap_8 FILLER_5_351 ();
 sg13g2_decap_8 FILLER_5_358 ();
 sg13g2_decap_8 FILLER_5_365 ();
 sg13g2_decap_8 FILLER_5_372 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_4 FILLER_6_21 ();
 sg13g2_fill_2 FILLER_6_33 ();
 sg13g2_fill_1 FILLER_6_35 ();
 sg13g2_decap_4 FILLER_6_44 ();
 sg13g2_fill_2 FILLER_6_48 ();
 sg13g2_decap_4 FILLER_6_71 ();
 sg13g2_decap_8 FILLER_6_101 ();
 sg13g2_decap_8 FILLER_6_142 ();
 sg13g2_decap_4 FILLER_6_149 ();
 sg13g2_fill_2 FILLER_6_153 ();
 sg13g2_decap_8 FILLER_6_164 ();
 sg13g2_fill_2 FILLER_6_171 ();
 sg13g2_decap_8 FILLER_6_177 ();
 sg13g2_decap_8 FILLER_6_194 ();
 sg13g2_fill_1 FILLER_6_201 ();
 sg13g2_decap_4 FILLER_6_207 ();
 sg13g2_decap_8 FILLER_6_237 ();
 sg13g2_decap_8 FILLER_6_268 ();
 sg13g2_decap_4 FILLER_6_275 ();
 sg13g2_fill_2 FILLER_6_279 ();
 sg13g2_fill_2 FILLER_6_286 ();
 sg13g2_fill_1 FILLER_6_288 ();
 sg13g2_fill_2 FILLER_6_310 ();
 sg13g2_decap_8 FILLER_6_338 ();
 sg13g2_decap_8 FILLER_6_345 ();
 sg13g2_decap_8 FILLER_6_352 ();
 sg13g2_decap_8 FILLER_6_359 ();
 sg13g2_decap_8 FILLER_6_366 ();
 sg13g2_decap_8 FILLER_6_373 ();
 sg13g2_decap_8 FILLER_6_380 ();
 sg13g2_decap_8 FILLER_6_387 ();
 sg13g2_decap_8 FILLER_6_394 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_4 FILLER_7_21 ();
 sg13g2_fill_2 FILLER_7_51 ();
 sg13g2_fill_1 FILLER_7_53 ();
 sg13g2_fill_1 FILLER_7_59 ();
 sg13g2_fill_1 FILLER_7_65 ();
 sg13g2_decap_8 FILLER_7_76 ();
 sg13g2_decap_8 FILLER_7_83 ();
 sg13g2_decap_8 FILLER_7_90 ();
 sg13g2_fill_2 FILLER_7_97 ();
 sg13g2_fill_1 FILLER_7_99 ();
 sg13g2_fill_2 FILLER_7_116 ();
 sg13g2_decap_4 FILLER_7_170 ();
 sg13g2_fill_1 FILLER_7_174 ();
 sg13g2_fill_2 FILLER_7_195 ();
 sg13g2_fill_2 FILLER_7_214 ();
 sg13g2_decap_8 FILLER_7_221 ();
 sg13g2_fill_1 FILLER_7_228 ();
 sg13g2_decap_8 FILLER_7_242 ();
 sg13g2_decap_4 FILLER_7_249 ();
 sg13g2_fill_2 FILLER_7_288 ();
 sg13g2_decap_4 FILLER_7_298 ();
 sg13g2_fill_1 FILLER_7_302 ();
 sg13g2_decap_8 FILLER_7_333 ();
 sg13g2_decap_8 FILLER_7_340 ();
 sg13g2_decap_8 FILLER_7_347 ();
 sg13g2_decap_8 FILLER_7_354 ();
 sg13g2_decap_8 FILLER_7_361 ();
 sg13g2_decap_8 FILLER_7_368 ();
 sg13g2_decap_8 FILLER_7_375 ();
 sg13g2_decap_8 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_7_389 ();
 sg13g2_decap_8 FILLER_7_396 ();
 sg13g2_decap_4 FILLER_7_403 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_4 FILLER_8_21 ();
 sg13g2_fill_2 FILLER_8_25 ();
 sg13g2_fill_2 FILLER_8_127 ();
 sg13g2_fill_1 FILLER_8_129 ();
 sg13g2_decap_8 FILLER_8_134 ();
 sg13g2_fill_2 FILLER_8_141 ();
 sg13g2_fill_1 FILLER_8_143 ();
 sg13g2_fill_2 FILLER_8_170 ();
 sg13g2_fill_1 FILLER_8_172 ();
 sg13g2_fill_2 FILLER_8_181 ();
 sg13g2_decap_8 FILLER_8_193 ();
 sg13g2_decap_8 FILLER_8_200 ();
 sg13g2_decap_4 FILLER_8_207 ();
 sg13g2_fill_2 FILLER_8_226 ();
 sg13g2_fill_1 FILLER_8_233 ();
 sg13g2_decap_4 FILLER_8_252 ();
 sg13g2_fill_1 FILLER_8_256 ();
 sg13g2_decap_8 FILLER_8_261 ();
 sg13g2_decap_8 FILLER_8_268 ();
 sg13g2_fill_1 FILLER_8_275 ();
 sg13g2_fill_2 FILLER_8_280 ();
 sg13g2_fill_1 FILLER_8_282 ();
 sg13g2_fill_1 FILLER_8_288 ();
 sg13g2_decap_8 FILLER_8_325 ();
 sg13g2_decap_8 FILLER_8_332 ();
 sg13g2_decap_8 FILLER_8_339 ();
 sg13g2_decap_8 FILLER_8_346 ();
 sg13g2_decap_8 FILLER_8_353 ();
 sg13g2_decap_8 FILLER_8_360 ();
 sg13g2_decap_8 FILLER_8_367 ();
 sg13g2_decap_8 FILLER_8_374 ();
 sg13g2_decap_8 FILLER_8_381 ();
 sg13g2_decap_8 FILLER_8_388 ();
 sg13g2_decap_8 FILLER_8_395 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_fill_2 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_41 ();
 sg13g2_fill_2 FILLER_9_48 ();
 sg13g2_fill_1 FILLER_9_50 ();
 sg13g2_fill_2 FILLER_9_67 ();
 sg13g2_fill_1 FILLER_9_69 ();
 sg13g2_decap_8 FILLER_9_78 ();
 sg13g2_decap_4 FILLER_9_85 ();
 sg13g2_fill_2 FILLER_9_93 ();
 sg13g2_fill_2 FILLER_9_100 ();
 sg13g2_decap_4 FILLER_9_120 ();
 sg13g2_decap_4 FILLER_9_150 ();
 sg13g2_fill_1 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_159 ();
 sg13g2_decap_4 FILLER_9_166 ();
 sg13g2_fill_1 FILLER_9_170 ();
 sg13g2_fill_2 FILLER_9_197 ();
 sg13g2_decap_4 FILLER_9_225 ();
 sg13g2_fill_2 FILLER_9_263 ();
 sg13g2_fill_1 FILLER_9_265 ();
 sg13g2_fill_1 FILLER_9_292 ();
 sg13g2_fill_2 FILLER_9_307 ();
 sg13g2_fill_1 FILLER_9_309 ();
 sg13g2_decap_8 FILLER_9_325 ();
 sg13g2_decap_8 FILLER_9_342 ();
 sg13g2_decap_8 FILLER_9_349 ();
 sg13g2_decap_8 FILLER_9_356 ();
 sg13g2_decap_8 FILLER_9_363 ();
 sg13g2_decap_8 FILLER_9_370 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_384 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_fill_2 FILLER_10_42 ();
 sg13g2_fill_2 FILLER_10_65 ();
 sg13g2_decap_8 FILLER_10_118 ();
 sg13g2_decap_8 FILLER_10_125 ();
 sg13g2_decap_4 FILLER_10_132 ();
 sg13g2_fill_1 FILLER_10_136 ();
 sg13g2_decap_8 FILLER_10_145 ();
 sg13g2_decap_8 FILLER_10_186 ();
 sg13g2_fill_2 FILLER_10_193 ();
 sg13g2_fill_2 FILLER_10_208 ();
 sg13g2_fill_1 FILLER_10_210 ();
 sg13g2_fill_1 FILLER_10_251 ();
 sg13g2_fill_1 FILLER_10_261 ();
 sg13g2_fill_1 FILLER_10_301 ();
 sg13g2_fill_1 FILLER_10_325 ();
 sg13g2_decap_8 FILLER_10_349 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_decap_8 FILLER_10_363 ();
 sg13g2_decap_8 FILLER_10_370 ();
 sg13g2_decap_8 FILLER_10_377 ();
 sg13g2_decap_8 FILLER_10_384 ();
 sg13g2_decap_8 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_398 ();
 sg13g2_decap_4 FILLER_10_405 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_fill_2 FILLER_11_49 ();
 sg13g2_fill_1 FILLER_11_51 ();
 sg13g2_fill_2 FILLER_11_57 ();
 sg13g2_decap_8 FILLER_11_68 ();
 sg13g2_fill_2 FILLER_11_75 ();
 sg13g2_fill_1 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_82 ();
 sg13g2_fill_2 FILLER_11_89 ();
 sg13g2_fill_1 FILLER_11_91 ();
 sg13g2_fill_1 FILLER_11_104 ();
 sg13g2_decap_4 FILLER_11_110 ();
 sg13g2_fill_1 FILLER_11_114 ();
 sg13g2_decap_4 FILLER_11_122 ();
 sg13g2_decap_8 FILLER_11_152 ();
 sg13g2_decap_4 FILLER_11_159 ();
 sg13g2_fill_1 FILLER_11_167 ();
 sg13g2_decap_4 FILLER_11_181 ();
 sg13g2_fill_2 FILLER_11_190 ();
 sg13g2_decap_4 FILLER_11_201 ();
 sg13g2_fill_2 FILLER_11_210 ();
 sg13g2_fill_1 FILLER_11_212 ();
 sg13g2_fill_1 FILLER_11_231 ();
 sg13g2_fill_2 FILLER_11_255 ();
 sg13g2_decap_4 FILLER_11_283 ();
 sg13g2_fill_1 FILLER_11_287 ();
 sg13g2_fill_2 FILLER_11_297 ();
 sg13g2_decap_8 FILLER_11_309 ();
 sg13g2_decap_4 FILLER_11_316 ();
 sg13g2_fill_2 FILLER_11_320 ();
 sg13g2_decap_8 FILLER_11_348 ();
 sg13g2_decap_8 FILLER_11_355 ();
 sg13g2_decap_8 FILLER_11_362 ();
 sg13g2_decap_8 FILLER_11_369 ();
 sg13g2_decap_8 FILLER_11_376 ();
 sg13g2_decap_8 FILLER_11_383 ();
 sg13g2_decap_8 FILLER_11_390 ();
 sg13g2_decap_8 FILLER_11_397 ();
 sg13g2_decap_4 FILLER_11_404 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_4 FILLER_12_28 ();
 sg13g2_fill_1 FILLER_12_32 ();
 sg13g2_decap_8 FILLER_12_37 ();
 sg13g2_fill_2 FILLER_12_44 ();
 sg13g2_decap_4 FILLER_12_105 ();
 sg13g2_fill_2 FILLER_12_117 ();
 sg13g2_fill_2 FILLER_12_124 ();
 sg13g2_decap_8 FILLER_12_152 ();
 sg13g2_decap_4 FILLER_12_159 ();
 sg13g2_decap_4 FILLER_12_180 ();
 sg13g2_fill_1 FILLER_12_184 ();
 sg13g2_decap_8 FILLER_12_211 ();
 sg13g2_fill_2 FILLER_12_237 ();
 sg13g2_fill_1 FILLER_12_255 ();
 sg13g2_fill_2 FILLER_12_321 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_fill_2 FILLER_12_343 ();
 sg13g2_fill_1 FILLER_12_345 ();
 sg13g2_fill_2 FILLER_12_362 ();
 sg13g2_fill_1 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_388 ();
 sg13g2_decap_8 FILLER_12_395 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_fill_1 FILLER_13_21 ();
 sg13g2_fill_2 FILLER_13_48 ();
 sg13g2_fill_1 FILLER_13_76 ();
 sg13g2_decap_8 FILLER_13_81 ();
 sg13g2_fill_2 FILLER_13_93 ();
 sg13g2_decap_8 FILLER_13_118 ();
 sg13g2_fill_2 FILLER_13_125 ();
 sg13g2_fill_2 FILLER_13_153 ();
 sg13g2_fill_1 FILLER_13_155 ();
 sg13g2_fill_1 FILLER_13_168 ();
 sg13g2_fill_1 FILLER_13_174 ();
 sg13g2_decap_8 FILLER_13_188 ();
 sg13g2_fill_1 FILLER_13_257 ();
 sg13g2_fill_1 FILLER_13_263 ();
 sg13g2_fill_1 FILLER_13_273 ();
 sg13g2_fill_1 FILLER_13_290 ();
 sg13g2_fill_1 FILLER_13_299 ();
 sg13g2_decap_4 FILLER_13_305 ();
 sg13g2_fill_1 FILLER_13_309 ();
 sg13g2_decap_8 FILLER_13_328 ();
 sg13g2_decap_4 FILLER_13_335 ();
 sg13g2_fill_1 FILLER_13_339 ();
 sg13g2_fill_2 FILLER_13_356 ();
 sg13g2_decap_4 FILLER_13_374 ();
 sg13g2_decap_8 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_67 ();
 sg13g2_decap_8 FILLER_14_74 ();
 sg13g2_fill_2 FILLER_14_81 ();
 sg13g2_fill_1 FILLER_14_83 ();
 sg13g2_fill_2 FILLER_14_136 ();
 sg13g2_decap_8 FILLER_14_146 ();
 sg13g2_fill_2 FILLER_14_153 ();
 sg13g2_fill_2 FILLER_14_188 ();
 sg13g2_fill_2 FILLER_14_203 ();
 sg13g2_fill_1 FILLER_14_205 ();
 sg13g2_fill_1 FILLER_14_219 ();
 sg13g2_decap_8 FILLER_14_229 ();
 sg13g2_fill_1 FILLER_14_236 ();
 sg13g2_fill_2 FILLER_14_245 ();
 sg13g2_fill_2 FILLER_14_258 ();
 sg13g2_fill_2 FILLER_14_286 ();
 sg13g2_fill_2 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_318 ();
 sg13g2_fill_2 FILLER_14_325 ();
 sg13g2_fill_1 FILLER_14_327 ();
 sg13g2_decap_4 FILLER_14_355 ();
 sg13g2_fill_1 FILLER_14_369 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_4 FILLER_14_382 ();
 sg13g2_fill_1 FILLER_14_386 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_fill_1 FILLER_15_28 ();
 sg13g2_fill_1 FILLER_15_55 ();
 sg13g2_fill_1 FILLER_15_64 ();
 sg13g2_decap_4 FILLER_15_70 ();
 sg13g2_fill_1 FILLER_15_87 ();
 sg13g2_decap_4 FILLER_15_95 ();
 sg13g2_decap_8 FILLER_15_104 ();
 sg13g2_decap_8 FILLER_15_111 ();
 sg13g2_fill_1 FILLER_15_127 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_fill_2 FILLER_15_161 ();
 sg13g2_fill_1 FILLER_15_166 ();
 sg13g2_fill_2 FILLER_15_172 ();
 sg13g2_fill_2 FILLER_15_179 ();
 sg13g2_fill_1 FILLER_15_188 ();
 sg13g2_fill_2 FILLER_15_193 ();
 sg13g2_fill_2 FILLER_15_208 ();
 sg13g2_fill_1 FILLER_15_210 ();
 sg13g2_fill_1 FILLER_15_221 ();
 sg13g2_fill_1 FILLER_15_253 ();
 sg13g2_decap_4 FILLER_15_278 ();
 sg13g2_decap_4 FILLER_15_285 ();
 sg13g2_fill_2 FILLER_15_289 ();
 sg13g2_fill_1 FILLER_15_296 ();
 sg13g2_decap_8 FILLER_15_312 ();
 sg13g2_fill_2 FILLER_15_319 ();
 sg13g2_fill_2 FILLER_15_325 ();
 sg13g2_fill_1 FILLER_15_327 ();
 sg13g2_fill_2 FILLER_15_339 ();
 sg13g2_decap_8 FILLER_15_346 ();
 sg13g2_fill_1 FILLER_15_353 ();
 sg13g2_decap_4 FILLER_15_370 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_4 FILLER_16_35 ();
 sg13g2_decap_4 FILLER_16_43 ();
 sg13g2_decap_8 FILLER_16_68 ();
 sg13g2_decap_4 FILLER_16_75 ();
 sg13g2_fill_2 FILLER_16_79 ();
 sg13g2_fill_2 FILLER_16_89 ();
 sg13g2_fill_2 FILLER_16_103 ();
 sg13g2_decap_8 FILLER_16_111 ();
 sg13g2_decap_8 FILLER_16_118 ();
 sg13g2_fill_1 FILLER_16_125 ();
 sg13g2_decap_8 FILLER_16_130 ();
 sg13g2_fill_2 FILLER_16_137 ();
 sg13g2_decap_8 FILLER_16_143 ();
 sg13g2_fill_2 FILLER_16_166 ();
 sg13g2_fill_2 FILLER_16_195 ();
 sg13g2_fill_1 FILLER_16_220 ();
 sg13g2_decap_4 FILLER_16_228 ();
 sg13g2_fill_1 FILLER_16_232 ();
 sg13g2_decap_4 FILLER_16_246 ();
 sg13g2_fill_2 FILLER_16_250 ();
 sg13g2_fill_2 FILLER_16_300 ();
 sg13g2_fill_2 FILLER_16_332 ();
 sg13g2_fill_1 FILLER_16_334 ();
 sg13g2_decap_4 FILLER_16_348 ();
 sg13g2_fill_2 FILLER_16_352 ();
 sg13g2_fill_1 FILLER_16_368 ();
 sg13g2_decap_4 FILLER_16_378 ();
 sg13g2_fill_1 FILLER_16_382 ();
 sg13g2_decap_4 FILLER_16_404 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_fill_1 FILLER_17_82 ();
 sg13g2_fill_1 FILLER_17_95 ();
 sg13g2_fill_1 FILLER_17_101 ();
 sg13g2_fill_1 FILLER_17_107 ();
 sg13g2_fill_2 FILLER_17_113 ();
 sg13g2_decap_8 FILLER_17_141 ();
 sg13g2_fill_2 FILLER_17_148 ();
 sg13g2_fill_1 FILLER_17_158 ();
 sg13g2_fill_2 FILLER_17_168 ();
 sg13g2_fill_1 FILLER_17_170 ();
 sg13g2_fill_2 FILLER_17_179 ();
 sg13g2_fill_2 FILLER_17_207 ();
 sg13g2_fill_1 FILLER_17_214 ();
 sg13g2_decap_8 FILLER_17_267 ();
 sg13g2_decap_8 FILLER_17_274 ();
 sg13g2_decap_4 FILLER_17_281 ();
 sg13g2_fill_1 FILLER_17_285 ();
 sg13g2_decap_8 FILLER_17_290 ();
 sg13g2_fill_2 FILLER_17_297 ();
 sg13g2_fill_2 FILLER_17_316 ();
 sg13g2_fill_1 FILLER_17_318 ();
 sg13g2_fill_2 FILLER_17_351 ();
 sg13g2_fill_1 FILLER_17_363 ();
 sg13g2_fill_2 FILLER_17_369 ();
 sg13g2_fill_2 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_4 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_71 ();
 sg13g2_decap_8 FILLER_18_78 ();
 sg13g2_fill_2 FILLER_18_85 ();
 sg13g2_decap_4 FILLER_18_116 ();
 sg13g2_fill_1 FILLER_18_120 ();
 sg13g2_fill_2 FILLER_18_147 ();
 sg13g2_fill_2 FILLER_18_165 ();
 sg13g2_fill_1 FILLER_18_167 ();
 sg13g2_decap_8 FILLER_18_173 ();
 sg13g2_fill_2 FILLER_18_180 ();
 sg13g2_fill_1 FILLER_18_190 ();
 sg13g2_fill_1 FILLER_18_195 ();
 sg13g2_fill_2 FILLER_18_205 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_4 FILLER_18_275 ();
 sg13g2_fill_2 FILLER_18_279 ();
 sg13g2_fill_1 FILLER_18_302 ();
 sg13g2_fill_2 FILLER_18_308 ();
 sg13g2_fill_1 FILLER_18_310 ();
 sg13g2_fill_1 FILLER_18_320 ();
 sg13g2_fill_1 FILLER_18_331 ();
 sg13g2_fill_2 FILLER_18_345 ();
 sg13g2_fill_2 FILLER_18_351 ();
 sg13g2_fill_2 FILLER_18_363 ();
 sg13g2_decap_4 FILLER_18_379 ();
 sg13g2_decap_4 FILLER_18_404 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_fill_2 FILLER_19_56 ();
 sg13g2_fill_1 FILLER_19_58 ();
 sg13g2_decap_4 FILLER_19_85 ();
 sg13g2_fill_2 FILLER_19_89 ();
 sg13g2_fill_1 FILLER_19_96 ();
 sg13g2_decap_8 FILLER_19_102 ();
 sg13g2_fill_2 FILLER_19_109 ();
 sg13g2_fill_1 FILLER_19_111 ();
 sg13g2_decap_8 FILLER_19_125 ();
 sg13g2_decap_4 FILLER_19_141 ();
 sg13g2_fill_2 FILLER_19_155 ();
 sg13g2_fill_1 FILLER_19_172 ();
 sg13g2_fill_1 FILLER_19_181 ();
 sg13g2_fill_2 FILLER_19_216 ();
 sg13g2_fill_2 FILLER_19_230 ();
 sg13g2_fill_1 FILLER_19_261 ();
 sg13g2_fill_2 FILLER_19_289 ();
 sg13g2_fill_1 FILLER_19_291 ();
 sg13g2_fill_2 FILLER_19_297 ();
 sg13g2_fill_2 FILLER_19_304 ();
 sg13g2_decap_8 FILLER_19_335 ();
 sg13g2_fill_2 FILLER_19_351 ();
 sg13g2_fill_1 FILLER_19_353 ();
 sg13g2_fill_2 FILLER_19_378 ();
 sg13g2_fill_1 FILLER_19_380 ();
 sg13g2_fill_1 FILLER_19_393 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_fill_2 FILLER_20_35 ();
 sg13g2_decap_4 FILLER_20_63 ();
 sg13g2_fill_1 FILLER_20_67 ();
 sg13g2_fill_2 FILLER_20_80 ();
 sg13g2_fill_1 FILLER_20_82 ();
 sg13g2_fill_2 FILLER_20_103 ();
 sg13g2_fill_1 FILLER_20_131 ();
 sg13g2_fill_2 FILLER_20_163 ();
 sg13g2_fill_1 FILLER_20_165 ();
 sg13g2_fill_2 FILLER_20_178 ();
 sg13g2_fill_1 FILLER_20_193 ();
 sg13g2_fill_1 FILLER_20_208 ();
 sg13g2_fill_2 FILLER_20_223 ();
 sg13g2_fill_1 FILLER_20_225 ();
 sg13g2_decap_4 FILLER_20_253 ();
 sg13g2_fill_2 FILLER_20_257 ();
 sg13g2_fill_1 FILLER_20_268 ();
 sg13g2_fill_1 FILLER_20_277 ();
 sg13g2_fill_2 FILLER_20_297 ();
 sg13g2_fill_1 FILLER_20_312 ();
 sg13g2_fill_1 FILLER_20_317 ();
 sg13g2_fill_2 FILLER_20_325 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_fill_2 FILLER_20_347 ();
 sg13g2_fill_1 FILLER_20_349 ();
 sg13g2_decap_4 FILLER_20_355 ();
 sg13g2_fill_1 FILLER_20_359 ();
 sg13g2_decap_4 FILLER_20_364 ();
 sg13g2_fill_2 FILLER_20_385 ();
 sg13g2_fill_1 FILLER_20_387 ();
 sg13g2_fill_1 FILLER_20_392 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_4 FILLER_21_21 ();
 sg13g2_fill_2 FILLER_21_25 ();
 sg13g2_decap_4 FILLER_21_43 ();
 sg13g2_fill_1 FILLER_21_47 ();
 sg13g2_decap_8 FILLER_21_52 ();
 sg13g2_fill_2 FILLER_21_59 ();
 sg13g2_fill_1 FILLER_21_61 ();
 sg13g2_fill_1 FILLER_21_85 ();
 sg13g2_decap_8 FILLER_21_102 ();
 sg13g2_decap_8 FILLER_21_109 ();
 sg13g2_fill_2 FILLER_21_124 ();
 sg13g2_decap_8 FILLER_21_138 ();
 sg13g2_fill_1 FILLER_21_145 ();
 sg13g2_decap_8 FILLER_21_157 ();
 sg13g2_fill_2 FILLER_21_164 ();
 sg13g2_decap_4 FILLER_21_262 ();
 sg13g2_fill_1 FILLER_21_266 ();
 sg13g2_fill_2 FILLER_21_295 ();
 sg13g2_fill_1 FILLER_21_319 ();
 sg13g2_fill_1 FILLER_21_325 ();
 sg13g2_fill_2 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_382 ();
 sg13g2_fill_1 FILLER_21_389 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_fill_2 FILLER_22_21 ();
 sg13g2_fill_1 FILLER_22_23 ();
 sg13g2_decap_8 FILLER_22_68 ();
 sg13g2_decap_4 FILLER_22_75 ();
 sg13g2_fill_1 FILLER_22_79 ();
 sg13g2_decap_4 FILLER_22_93 ();
 sg13g2_fill_2 FILLER_22_102 ();
 sg13g2_fill_1 FILLER_22_104 ();
 sg13g2_decap_4 FILLER_22_131 ();
 sg13g2_decap_4 FILLER_22_164 ();
 sg13g2_fill_1 FILLER_22_168 ();
 sg13g2_fill_2 FILLER_22_173 ();
 sg13g2_decap_8 FILLER_22_179 ();
 sg13g2_decap_8 FILLER_22_186 ();
 sg13g2_fill_1 FILLER_22_193 ();
 sg13g2_fill_2 FILLER_22_243 ();
 sg13g2_fill_1 FILLER_22_245 ();
 sg13g2_fill_2 FILLER_22_267 ();
 sg13g2_fill_1 FILLER_22_269 ();
 sg13g2_decap_8 FILLER_22_286 ();
 sg13g2_decap_4 FILLER_22_293 ();
 sg13g2_fill_1 FILLER_22_297 ();
 sg13g2_decap_4 FILLER_22_314 ();
 sg13g2_fill_2 FILLER_22_318 ();
 sg13g2_decap_8 FILLER_22_334 ();
 sg13g2_decap_4 FILLER_22_341 ();
 sg13g2_fill_2 FILLER_22_345 ();
 sg13g2_fill_2 FILLER_22_356 ();
 sg13g2_fill_2 FILLER_22_368 ();
 sg13g2_fill_1 FILLER_22_370 ();
 sg13g2_decap_4 FILLER_22_380 ();
 sg13g2_fill_1 FILLER_22_384 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_4 ();
 sg13g2_fill_2 FILLER_23_13 ();
 sg13g2_decap_4 FILLER_23_23 ();
 sg13g2_fill_2 FILLER_23_27 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_4 FILLER_23_49 ();
 sg13g2_fill_1 FILLER_23_53 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_fill_2 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_132 ();
 sg13g2_decap_4 FILLER_23_139 ();
 sg13g2_fill_2 FILLER_23_143 ();
 sg13g2_fill_1 FILLER_23_171 ();
 sg13g2_fill_1 FILLER_23_177 ();
 sg13g2_fill_2 FILLER_23_208 ();
 sg13g2_fill_2 FILLER_23_261 ();
 sg13g2_decap_4 FILLER_23_304 ();
 sg13g2_fill_1 FILLER_23_308 ();
 sg13g2_decap_4 FILLER_23_315 ();
 sg13g2_fill_2 FILLER_23_319 ();
 sg13g2_fill_2 FILLER_23_344 ();
 sg13g2_fill_2 FILLER_23_378 ();
 sg13g2_fill_1 FILLER_23_390 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_26 ();
 sg13g2_fill_1 FILLER_24_33 ();
 sg13g2_fill_1 FILLER_24_42 ();
 sg13g2_fill_2 FILLER_24_51 ();
 sg13g2_fill_1 FILLER_24_79 ();
 sg13g2_decap_8 FILLER_24_102 ();
 sg13g2_decap_8 FILLER_24_109 ();
 sg13g2_fill_1 FILLER_24_116 ();
 sg13g2_decap_8 FILLER_24_125 ();
 sg13g2_decap_4 FILLER_24_132 ();
 sg13g2_fill_2 FILLER_24_161 ();
 sg13g2_decap_4 FILLER_24_167 ();
 sg13g2_fill_2 FILLER_24_188 ();
 sg13g2_fill_1 FILLER_24_190 ();
 sg13g2_fill_2 FILLER_24_208 ();
 sg13g2_fill_1 FILLER_24_210 ();
 sg13g2_fill_1 FILLER_24_231 ();
 sg13g2_fill_1 FILLER_24_250 ();
 sg13g2_fill_1 FILLER_24_268 ();
 sg13g2_fill_1 FILLER_24_281 ();
 sg13g2_fill_1 FILLER_24_287 ();
 sg13g2_fill_2 FILLER_24_304 ();
 sg13g2_fill_1 FILLER_24_306 ();
 sg13g2_fill_2 FILLER_24_317 ();
 sg13g2_fill_2 FILLER_24_339 ();
 sg13g2_fill_1 FILLER_24_341 ();
 sg13g2_fill_2 FILLER_24_356 ();
 sg13g2_fill_2 FILLER_24_363 ();
 sg13g2_fill_1 FILLER_24_378 ();
 sg13g2_fill_1 FILLER_24_391 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_decap_4 FILLER_25_15 ();
 sg13g2_fill_2 FILLER_25_26 ();
 sg13g2_fill_1 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_57 ();
 sg13g2_decap_8 FILLER_25_68 ();
 sg13g2_decap_8 FILLER_25_75 ();
 sg13g2_fill_1 FILLER_25_82 ();
 sg13g2_decap_4 FILLER_25_104 ();
 sg13g2_fill_1 FILLER_25_108 ();
 sg13g2_decap_8 FILLER_25_135 ();
 sg13g2_decap_4 FILLER_25_142 ();
 sg13g2_fill_2 FILLER_25_146 ();
 sg13g2_decap_8 FILLER_25_153 ();
 sg13g2_fill_1 FILLER_25_260 ();
 sg13g2_decap_8 FILLER_25_275 ();
 sg13g2_decap_8 FILLER_25_282 ();
 sg13g2_decap_4 FILLER_25_289 ();
 sg13g2_decap_4 FILLER_25_314 ();
 sg13g2_decap_4 FILLER_25_322 ();
 sg13g2_fill_1 FILLER_25_326 ();
 sg13g2_fill_2 FILLER_25_342 ();
 sg13g2_fill_2 FILLER_25_356 ();
 sg13g2_fill_1 FILLER_25_358 ();
 sg13g2_decap_4 FILLER_25_364 ();
 sg13g2_fill_1 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_25_374 ();
 sg13g2_fill_2 FILLER_25_386 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_fill_1 FILLER_26_50 ();
 sg13g2_fill_2 FILLER_26_77 ();
 sg13g2_fill_2 FILLER_26_129 ();
 sg13g2_fill_1 FILLER_26_131 ();
 sg13g2_decap_4 FILLER_26_158 ();
 sg13g2_decap_8 FILLER_26_166 ();
 sg13g2_decap_8 FILLER_26_173 ();
 sg13g2_decap_4 FILLER_26_180 ();
 sg13g2_fill_2 FILLER_26_184 ();
 sg13g2_fill_1 FILLER_26_190 ();
 sg13g2_fill_1 FILLER_26_287 ();
 sg13g2_decap_4 FILLER_26_296 ();
 sg13g2_fill_2 FILLER_26_300 ();
 sg13g2_decap_8 FILLER_26_307 ();
 sg13g2_decap_4 FILLER_26_314 ();
 sg13g2_decap_8 FILLER_26_334 ();
 sg13g2_decap_4 FILLER_26_341 ();
 sg13g2_decap_4 FILLER_26_353 ();
 sg13g2_fill_1 FILLER_26_357 ();
 sg13g2_fill_1 FILLER_26_362 ();
 sg13g2_decap_8 FILLER_26_372 ();
 sg13g2_fill_1 FILLER_26_387 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_fill_1 FILLER_27_15 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_4 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_52 ();
 sg13g2_fill_2 FILLER_27_59 ();
 sg13g2_fill_1 FILLER_27_61 ();
 sg13g2_decap_8 FILLER_27_66 ();
 sg13g2_decap_8 FILLER_27_73 ();
 sg13g2_fill_1 FILLER_27_80 ();
 sg13g2_fill_2 FILLER_27_86 ();
 sg13g2_fill_1 FILLER_27_88 ();
 sg13g2_decap_8 FILLER_27_94 ();
 sg13g2_decap_4 FILLER_27_101 ();
 sg13g2_fill_1 FILLER_27_105 ();
 sg13g2_fill_2 FILLER_27_111 ();
 sg13g2_fill_1 FILLER_27_113 ();
 sg13g2_fill_2 FILLER_27_123 ();
 sg13g2_fill_1 FILLER_27_125 ();
 sg13g2_fill_1 FILLER_27_134 ();
 sg13g2_decap_4 FILLER_27_147 ();
 sg13g2_fill_1 FILLER_27_151 ();
 sg13g2_fill_2 FILLER_27_231 ();
 sg13g2_fill_1 FILLER_27_233 ();
 sg13g2_fill_1 FILLER_27_247 ();
 sg13g2_fill_2 FILLER_27_269 ();
 sg13g2_fill_2 FILLER_27_297 ();
 sg13g2_fill_2 FILLER_27_323 ();
 sg13g2_fill_1 FILLER_27_325 ();
 sg13g2_decap_4 FILLER_27_331 ();
 sg13g2_fill_2 FILLER_27_357 ();
 sg13g2_fill_1 FILLER_27_359 ();
 sg13g2_decap_8 FILLER_27_383 ();
 sg13g2_fill_2 FILLER_27_390 ();
 sg13g2_fill_1 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_397 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_15 ();
 sg13g2_decap_8 FILLER_28_24 ();
 sg13g2_fill_2 FILLER_28_51 ();
 sg13g2_decap_4 FILLER_28_79 ();
 sg13g2_fill_2 FILLER_28_98 ();
 sg13g2_decap_4 FILLER_28_126 ();
 sg13g2_fill_1 FILLER_28_149 ();
 sg13g2_decap_4 FILLER_28_158 ();
 sg13g2_fill_1 FILLER_28_162 ();
 sg13g2_decap_4 FILLER_28_189 ();
 sg13g2_decap_4 FILLER_28_197 ();
 sg13g2_fill_1 FILLER_28_201 ();
 sg13g2_fill_2 FILLER_28_215 ();
 sg13g2_fill_1 FILLER_28_259 ();
 sg13g2_decap_4 FILLER_28_276 ();
 sg13g2_fill_2 FILLER_28_280 ();
 sg13g2_fill_2 FILLER_28_307 ();
 sg13g2_fill_2 FILLER_28_314 ();
 sg13g2_fill_2 FILLER_28_321 ();
 sg13g2_fill_1 FILLER_28_323 ();
 sg13g2_fill_2 FILLER_28_337 ();
 sg13g2_decap_4 FILLER_28_354 ();
 sg13g2_fill_2 FILLER_28_386 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_fill_2 FILLER_29_26 ();
 sg13g2_fill_1 FILLER_29_28 ();
 sg13g2_decap_4 FILLER_29_40 ();
 sg13g2_decap_8 FILLER_29_57 ();
 sg13g2_decap_8 FILLER_29_68 ();
 sg13g2_fill_2 FILLER_29_75 ();
 sg13g2_fill_2 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_100 ();
 sg13g2_decap_4 FILLER_29_107 ();
 sg13g2_decap_8 FILLER_29_115 ();
 sg13g2_decap_4 FILLER_29_122 ();
 sg13g2_fill_2 FILLER_29_136 ();
 sg13g2_fill_1 FILLER_29_138 ();
 sg13g2_fill_1 FILLER_29_163 ();
 sg13g2_decap_4 FILLER_29_169 ();
 sg13g2_fill_1 FILLER_29_173 ();
 sg13g2_decap_8 FILLER_29_178 ();
 sg13g2_decap_8 FILLER_29_185 ();
 sg13g2_fill_1 FILLER_29_251 ();
 sg13g2_fill_1 FILLER_29_290 ();
 sg13g2_decap_8 FILLER_29_307 ();
 sg13g2_decap_4 FILLER_29_324 ();
 sg13g2_fill_2 FILLER_29_328 ();
 sg13g2_fill_2 FILLER_29_335 ();
 sg13g2_fill_1 FILLER_29_337 ();
 sg13g2_decap_8 FILLER_29_342 ();
 sg13g2_fill_1 FILLER_29_349 ();
 sg13g2_fill_1 FILLER_29_368 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_2 ();
 sg13g2_fill_1 FILLER_30_16 ();
 sg13g2_fill_2 FILLER_30_27 ();
 sg13g2_fill_2 FILLER_30_45 ();
 sg13g2_fill_1 FILLER_30_47 ();
 sg13g2_fill_2 FILLER_30_74 ();
 sg13g2_fill_1 FILLER_30_76 ();
 sg13g2_decap_8 FILLER_30_111 ();
 sg13g2_fill_2 FILLER_30_118 ();
 sg13g2_fill_1 FILLER_30_120 ();
 sg13g2_decap_8 FILLER_30_137 ();
 sg13g2_fill_2 FILLER_30_144 ();
 sg13g2_fill_1 FILLER_30_146 ();
 sg13g2_fill_2 FILLER_30_155 ();
 sg13g2_fill_2 FILLER_30_175 ();
 sg13g2_decap_4 FILLER_30_210 ();
 sg13g2_fill_2 FILLER_30_214 ();
 sg13g2_fill_2 FILLER_30_238 ();
 sg13g2_fill_2 FILLER_30_245 ();
 sg13g2_fill_1 FILLER_30_247 ();
 sg13g2_decap_8 FILLER_30_274 ();
 sg13g2_fill_2 FILLER_30_281 ();
 sg13g2_fill_2 FILLER_30_303 ();
 sg13g2_decap_4 FILLER_30_342 ();
 sg13g2_fill_1 FILLER_30_356 ();
 sg13g2_fill_1 FILLER_30_367 ();
 sg13g2_decap_4 FILLER_30_377 ();
 sg13g2_fill_1 FILLER_30_390 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_4 ();
 sg13g2_decap_4 FILLER_31_13 ();
 sg13g2_fill_1 FILLER_31_31 ();
 sg13g2_fill_2 FILLER_31_36 ();
 sg13g2_decap_8 FILLER_31_43 ();
 sg13g2_decap_4 FILLER_31_50 ();
 sg13g2_fill_2 FILLER_31_54 ();
 sg13g2_decap_8 FILLER_31_65 ();
 sg13g2_fill_2 FILLER_31_72 ();
 sg13g2_decap_8 FILLER_31_89 ();
 sg13g2_fill_1 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_180 ();
 sg13g2_fill_1 FILLER_31_187 ();
 sg13g2_decap_8 FILLER_31_192 ();
 sg13g2_fill_1 FILLER_31_199 ();
 sg13g2_fill_1 FILLER_31_213 ();
 sg13g2_fill_1 FILLER_31_219 ();
 sg13g2_decap_4 FILLER_31_254 ();
 sg13g2_decap_8 FILLER_31_262 ();
 sg13g2_decap_8 FILLER_31_269 ();
 sg13g2_decap_8 FILLER_31_276 ();
 sg13g2_fill_2 FILLER_31_306 ();
 sg13g2_fill_2 FILLER_31_337 ();
 sg13g2_fill_2 FILLER_31_360 ();
 sg13g2_fill_1 FILLER_31_362 ();
 sg13g2_fill_2 FILLER_31_371 ();
 sg13g2_fill_2 FILLER_31_384 ();
 sg13g2_fill_1 FILLER_31_386 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_44 ();
 sg13g2_fill_1 FILLER_32_46 ();
 sg13g2_fill_2 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_4 FILLER_32_98 ();
 sg13g2_fill_1 FILLER_32_106 ();
 sg13g2_decap_8 FILLER_32_111 ();
 sg13g2_decap_4 FILLER_32_118 ();
 sg13g2_fill_1 FILLER_32_122 ();
 sg13g2_decap_8 FILLER_32_136 ();
 sg13g2_fill_2 FILLER_32_143 ();
 sg13g2_fill_1 FILLER_32_145 ();
 sg13g2_decap_8 FILLER_32_150 ();
 sg13g2_decap_4 FILLER_32_157 ();
 sg13g2_fill_2 FILLER_32_179 ();
 sg13g2_decap_8 FILLER_32_190 ();
 sg13g2_decap_8 FILLER_32_201 ();
 sg13g2_fill_2 FILLER_32_208 ();
 sg13g2_fill_1 FILLER_32_210 ();
 sg13g2_decap_4 FILLER_32_255 ();
 sg13g2_fill_2 FILLER_32_259 ();
 sg13g2_fill_1 FILLER_32_282 ();
 sg13g2_fill_2 FILLER_32_287 ();
 sg13g2_fill_1 FILLER_32_289 ();
 sg13g2_decap_4 FILLER_32_298 ();
 sg13g2_fill_2 FILLER_32_302 ();
 sg13g2_decap_8 FILLER_32_324 ();
 sg13g2_decap_8 FILLER_32_331 ();
 sg13g2_decap_4 FILLER_32_353 ();
 sg13g2_fill_1 FILLER_32_357 ();
 sg13g2_decap_4 FILLER_32_374 ();
 sg13g2_fill_2 FILLER_32_387 ();
 sg13g2_fill_1 FILLER_32_389 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_11 ();
 sg13g2_decap_8 FILLER_33_16 ();
 sg13g2_decap_4 FILLER_33_23 ();
 sg13g2_fill_2 FILLER_33_27 ();
 sg13g2_decap_4 FILLER_33_63 ();
 sg13g2_fill_1 FILLER_33_67 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_fill_2 FILLER_33_117 ();
 sg13g2_fill_1 FILLER_33_119 ();
 sg13g2_fill_2 FILLER_33_136 ();
 sg13g2_decap_4 FILLER_33_164 ();
 sg13g2_fill_2 FILLER_33_184 ();
 sg13g2_fill_2 FILLER_33_212 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_fill_2 FILLER_33_266 ();
 sg13g2_fill_1 FILLER_33_268 ();
 sg13g2_decap_8 FILLER_33_274 ();
 sg13g2_fill_1 FILLER_33_281 ();
 sg13g2_fill_2 FILLER_33_287 ();
 sg13g2_decap_8 FILLER_33_307 ();
 sg13g2_fill_1 FILLER_33_314 ();
 sg13g2_fill_1 FILLER_33_320 ();
 sg13g2_fill_2 FILLER_33_326 ();
 sg13g2_fill_2 FILLER_33_341 ();
 sg13g2_fill_1 FILLER_33_343 ();
 sg13g2_decap_8 FILLER_33_358 ();
 sg13g2_decap_4 FILLER_33_365 ();
 sg13g2_decap_8 FILLER_33_374 ();
 sg13g2_decap_4 FILLER_33_381 ();
 sg13g2_fill_1 FILLER_33_389 ();
 sg13g2_decap_4 FILLER_33_404 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_30 ();
 sg13g2_fill_2 FILLER_34_35 ();
 sg13g2_fill_1 FILLER_34_37 ();
 sg13g2_fill_1 FILLER_34_42 ();
 sg13g2_decap_4 FILLER_34_107 ();
 sg13g2_fill_2 FILLER_34_116 ();
 sg13g2_fill_1 FILLER_34_118 ();
 sg13g2_fill_2 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_153 ();
 sg13g2_decap_4 FILLER_34_160 ();
 sg13g2_fill_2 FILLER_34_164 ();
 sg13g2_fill_1 FILLER_34_187 ();
 sg13g2_decap_4 FILLER_34_214 ();
 sg13g2_fill_2 FILLER_34_231 ();
 sg13g2_fill_2 FILLER_34_241 ();
 sg13g2_decap_8 FILLER_34_248 ();
 sg13g2_decap_4 FILLER_34_255 ();
 sg13g2_fill_1 FILLER_34_259 ();
 sg13g2_fill_2 FILLER_34_273 ();
 sg13g2_fill_1 FILLER_34_275 ();
 sg13g2_fill_2 FILLER_34_291 ();
 sg13g2_fill_2 FILLER_34_301 ();
 sg13g2_fill_1 FILLER_34_303 ();
 sg13g2_fill_2 FILLER_34_323 ();
 sg13g2_fill_2 FILLER_34_330 ();
 sg13g2_decap_4 FILLER_34_342 ();
 sg13g2_fill_1 FILLER_34_346 ();
 sg13g2_decap_4 FILLER_34_358 ();
 sg13g2_fill_2 FILLER_34_392 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_4 ();
 sg13g2_fill_2 FILLER_35_13 ();
 sg13g2_decap_8 FILLER_35_19 ();
 sg13g2_fill_1 FILLER_35_26 ();
 sg13g2_fill_2 FILLER_35_35 ();
 sg13g2_fill_2 FILLER_35_42 ();
 sg13g2_fill_1 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_62 ();
 sg13g2_fill_2 FILLER_35_69 ();
 sg13g2_fill_1 FILLER_35_71 ();
 sg13g2_fill_2 FILLER_35_77 ();
 sg13g2_decap_4 FILLER_35_83 ();
 sg13g2_fill_2 FILLER_35_87 ();
 sg13g2_fill_2 FILLER_35_106 ();
 sg13g2_fill_1 FILLER_35_118 ();
 sg13g2_fill_1 FILLER_35_132 ();
 sg13g2_fill_1 FILLER_35_141 ();
 sg13g2_fill_2 FILLER_35_168 ();
 sg13g2_fill_2 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_185 ();
 sg13g2_decap_8 FILLER_35_192 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_4 FILLER_35_210 ();
 sg13g2_fill_1 FILLER_35_227 ();
 sg13g2_fill_2 FILLER_35_256 ();
 sg13g2_decap_4 FILLER_35_335 ();
 sg13g2_decap_4 FILLER_35_359 ();
 sg13g2_decap_4 FILLER_35_377 ();
 sg13g2_fill_1 FILLER_35_381 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_4 ();
 sg13g2_fill_2 FILLER_36_31 ();
 sg13g2_decap_8 FILLER_36_36 ();
 sg13g2_fill_1 FILLER_36_43 ();
 sg13g2_decap_8 FILLER_36_55 ();
 sg13g2_fill_2 FILLER_36_62 ();
 sg13g2_fill_1 FILLER_36_64 ();
 sg13g2_fill_1 FILLER_36_77 ();
 sg13g2_decap_4 FILLER_36_87 ();
 sg13g2_fill_2 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_103 ();
 sg13g2_fill_1 FILLER_36_110 ();
 sg13g2_fill_1 FILLER_36_125 ();
 sg13g2_decap_8 FILLER_36_141 ();
 sg13g2_decap_4 FILLER_36_148 ();
 sg13g2_fill_1 FILLER_36_152 ();
 sg13g2_decap_8 FILLER_36_157 ();
 sg13g2_fill_2 FILLER_36_164 ();
 sg13g2_fill_2 FILLER_36_186 ();
 sg13g2_fill_1 FILLER_36_188 ();
 sg13g2_decap_8 FILLER_36_215 ();
 sg13g2_fill_2 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_245 ();
 sg13g2_fill_2 FILLER_36_252 ();
 sg13g2_fill_1 FILLER_36_254 ();
 sg13g2_fill_2 FILLER_36_261 ();
 sg13g2_fill_2 FILLER_36_268 ();
 sg13g2_fill_1 FILLER_36_270 ();
 sg13g2_decap_4 FILLER_36_275 ();
 sg13g2_fill_1 FILLER_36_279 ();
 sg13g2_decap_4 FILLER_36_284 ();
 sg13g2_fill_1 FILLER_36_288 ();
 sg13g2_decap_4 FILLER_36_293 ();
 sg13g2_decap_8 FILLER_36_302 ();
 sg13g2_decap_4 FILLER_36_309 ();
 sg13g2_fill_2 FILLER_36_334 ();
 sg13g2_fill_2 FILLER_36_341 ();
 sg13g2_fill_1 FILLER_36_343 ();
 sg13g2_decap_4 FILLER_36_349 ();
 sg13g2_fill_2 FILLER_36_353 ();
 sg13g2_fill_1 FILLER_36_374 ();
 sg13g2_fill_1 FILLER_36_383 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_fill_2 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_20 ();
 sg13g2_decap_8 FILLER_37_27 ();
 sg13g2_decap_8 FILLER_37_34 ();
 sg13g2_decap_8 FILLER_37_41 ();
 sg13g2_decap_8 FILLER_37_48 ();
 sg13g2_decap_8 FILLER_37_55 ();
 sg13g2_decap_4 FILLER_37_62 ();
 sg13g2_decap_4 FILLER_37_168 ();
 sg13g2_fill_2 FILLER_37_189 ();
 sg13g2_decap_4 FILLER_37_195 ();
 sg13g2_fill_1 FILLER_37_199 ();
 sg13g2_decap_8 FILLER_37_208 ();
 sg13g2_decap_8 FILLER_37_215 ();
 sg13g2_fill_2 FILLER_37_222 ();
 sg13g2_fill_2 FILLER_37_240 ();
 sg13g2_fill_1 FILLER_37_242 ();
 sg13g2_fill_2 FILLER_37_287 ();
 sg13g2_fill_2 FILLER_37_308 ();
 sg13g2_fill_2 FILLER_37_325 ();
 sg13g2_fill_1 FILLER_37_327 ();
 sg13g2_fill_2 FILLER_37_338 ();
 sg13g2_decap_8 FILLER_37_352 ();
 sg13g2_fill_2 FILLER_37_359 ();
 sg13g2_fill_1 FILLER_37_361 ();
 sg13g2_fill_2 FILLER_37_380 ();
 sg13g2_decap_4 FILLER_37_405 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_fill_2 FILLER_38_125 ();
 sg13g2_fill_2 FILLER_38_141 ();
 sg13g2_fill_1 FILLER_38_143 ();
 sg13g2_fill_1 FILLER_38_148 ();
 sg13g2_fill_2 FILLER_38_157 ();
 sg13g2_fill_2 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_decap_8 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_decap_4 FILLER_38_273 ();
 sg13g2_decap_8 FILLER_38_303 ();
 sg13g2_decap_8 FILLER_38_327 ();
 sg13g2_fill_2 FILLER_38_357 ();
 sg13g2_fill_1 FILLER_38_359 ();
 sg13g2_fill_2 FILLER_38_382 ();
 sg13g2_fill_1 FILLER_38_384 ();
 sg13g2_decap_4 FILLER_38_391 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
endmodule
